module dtc_split5_bm26 (
	input  wire [15-1:0] inp,
	output wire [15-1:0] outp
);

	wire [15-1:0] node1;
	wire [15-1:0] node2;
	wire [15-1:0] node3;
	wire [15-1:0] node4;
	wire [15-1:0] node5;
	wire [15-1:0] node6;
	wire [15-1:0] node7;
	wire [15-1:0] node8;
	wire [15-1:0] node9;
	wire [15-1:0] node10;
	wire [15-1:0] node11;
	wire [15-1:0] node12;
	wire [15-1:0] node15;
	wire [15-1:0] node18;
	wire [15-1:0] node19;
	wire [15-1:0] node22;
	wire [15-1:0] node25;
	wire [15-1:0] node26;
	wire [15-1:0] node27;
	wire [15-1:0] node30;
	wire [15-1:0] node33;
	wire [15-1:0] node34;
	wire [15-1:0] node37;
	wire [15-1:0] node40;
	wire [15-1:0] node41;
	wire [15-1:0] node42;
	wire [15-1:0] node43;
	wire [15-1:0] node46;
	wire [15-1:0] node49;
	wire [15-1:0] node50;
	wire [15-1:0] node53;
	wire [15-1:0] node56;
	wire [15-1:0] node57;
	wire [15-1:0] node58;
	wire [15-1:0] node61;
	wire [15-1:0] node64;
	wire [15-1:0] node65;
	wire [15-1:0] node69;
	wire [15-1:0] node70;
	wire [15-1:0] node71;
	wire [15-1:0] node72;
	wire [15-1:0] node74;
	wire [15-1:0] node77;
	wire [15-1:0] node78;
	wire [15-1:0] node81;
	wire [15-1:0] node84;
	wire [15-1:0] node85;
	wire [15-1:0] node86;
	wire [15-1:0] node89;
	wire [15-1:0] node92;
	wire [15-1:0] node93;
	wire [15-1:0] node96;
	wire [15-1:0] node99;
	wire [15-1:0] node100;
	wire [15-1:0] node101;
	wire [15-1:0] node102;
	wire [15-1:0] node105;
	wire [15-1:0] node108;
	wire [15-1:0] node109;
	wire [15-1:0] node112;
	wire [15-1:0] node115;
	wire [15-1:0] node116;
	wire [15-1:0] node117;
	wire [15-1:0] node120;
	wire [15-1:0] node123;
	wire [15-1:0] node124;
	wire [15-1:0] node127;
	wire [15-1:0] node130;
	wire [15-1:0] node131;
	wire [15-1:0] node132;
	wire [15-1:0] node133;
	wire [15-1:0] node134;
	wire [15-1:0] node135;
	wire [15-1:0] node138;
	wire [15-1:0] node141;
	wire [15-1:0] node142;
	wire [15-1:0] node145;
	wire [15-1:0] node148;
	wire [15-1:0] node149;
	wire [15-1:0] node150;
	wire [15-1:0] node153;
	wire [15-1:0] node156;
	wire [15-1:0] node157;
	wire [15-1:0] node160;
	wire [15-1:0] node163;
	wire [15-1:0] node164;
	wire [15-1:0] node165;
	wire [15-1:0] node166;
	wire [15-1:0] node169;
	wire [15-1:0] node172;
	wire [15-1:0] node173;
	wire [15-1:0] node176;
	wire [15-1:0] node179;
	wire [15-1:0] node180;
	wire [15-1:0] node181;
	wire [15-1:0] node184;
	wire [15-1:0] node187;
	wire [15-1:0] node188;
	wire [15-1:0] node192;
	wire [15-1:0] node193;
	wire [15-1:0] node194;
	wire [15-1:0] node195;
	wire [15-1:0] node196;
	wire [15-1:0] node199;
	wire [15-1:0] node202;
	wire [15-1:0] node203;
	wire [15-1:0] node206;
	wire [15-1:0] node209;
	wire [15-1:0] node210;
	wire [15-1:0] node211;
	wire [15-1:0] node214;
	wire [15-1:0] node217;
	wire [15-1:0] node218;
	wire [15-1:0] node221;
	wire [15-1:0] node224;
	wire [15-1:0] node225;
	wire [15-1:0] node226;
	wire [15-1:0] node227;
	wire [15-1:0] node230;
	wire [15-1:0] node233;
	wire [15-1:0] node234;
	wire [15-1:0] node237;
	wire [15-1:0] node240;
	wire [15-1:0] node241;
	wire [15-1:0] node243;
	wire [15-1:0] node246;
	wire [15-1:0] node248;
	wire [15-1:0] node251;
	wire [15-1:0] node252;
	wire [15-1:0] node253;
	wire [15-1:0] node254;
	wire [15-1:0] node255;
	wire [15-1:0] node256;
	wire [15-1:0] node257;
	wire [15-1:0] node260;
	wire [15-1:0] node263;
	wire [15-1:0] node264;
	wire [15-1:0] node267;
	wire [15-1:0] node270;
	wire [15-1:0] node271;
	wire [15-1:0] node272;
	wire [15-1:0] node275;
	wire [15-1:0] node278;
	wire [15-1:0] node279;
	wire [15-1:0] node282;
	wire [15-1:0] node285;
	wire [15-1:0] node286;
	wire [15-1:0] node287;
	wire [15-1:0] node288;
	wire [15-1:0] node291;
	wire [15-1:0] node294;
	wire [15-1:0] node295;
	wire [15-1:0] node299;
	wire [15-1:0] node300;
	wire [15-1:0] node301;
	wire [15-1:0] node304;
	wire [15-1:0] node307;
	wire [15-1:0] node308;
	wire [15-1:0] node311;
	wire [15-1:0] node314;
	wire [15-1:0] node315;
	wire [15-1:0] node316;
	wire [15-1:0] node317;
	wire [15-1:0] node318;
	wire [15-1:0] node321;
	wire [15-1:0] node324;
	wire [15-1:0] node325;
	wire [15-1:0] node328;
	wire [15-1:0] node331;
	wire [15-1:0] node332;
	wire [15-1:0] node333;
	wire [15-1:0] node336;
	wire [15-1:0] node339;
	wire [15-1:0] node340;
	wire [15-1:0] node343;
	wire [15-1:0] node346;
	wire [15-1:0] node347;
	wire [15-1:0] node348;
	wire [15-1:0] node349;
	wire [15-1:0] node352;
	wire [15-1:0] node355;
	wire [15-1:0] node356;
	wire [15-1:0] node359;
	wire [15-1:0] node362;
	wire [15-1:0] node363;
	wire [15-1:0] node364;
	wire [15-1:0] node367;
	wire [15-1:0] node370;
	wire [15-1:0] node371;
	wire [15-1:0] node374;
	wire [15-1:0] node377;
	wire [15-1:0] node378;
	wire [15-1:0] node379;
	wire [15-1:0] node380;
	wire [15-1:0] node381;
	wire [15-1:0] node382;
	wire [15-1:0] node385;
	wire [15-1:0] node388;
	wire [15-1:0] node389;
	wire [15-1:0] node392;
	wire [15-1:0] node395;
	wire [15-1:0] node396;
	wire [15-1:0] node397;
	wire [15-1:0] node400;
	wire [15-1:0] node403;
	wire [15-1:0] node404;
	wire [15-1:0] node407;
	wire [15-1:0] node410;
	wire [15-1:0] node411;
	wire [15-1:0] node412;
	wire [15-1:0] node413;
	wire [15-1:0] node416;
	wire [15-1:0] node419;
	wire [15-1:0] node420;
	wire [15-1:0] node423;
	wire [15-1:0] node426;
	wire [15-1:0] node427;
	wire [15-1:0] node428;
	wire [15-1:0] node431;
	wire [15-1:0] node434;
	wire [15-1:0] node435;
	wire [15-1:0] node438;
	wire [15-1:0] node441;
	wire [15-1:0] node442;
	wire [15-1:0] node443;
	wire [15-1:0] node444;
	wire [15-1:0] node445;
	wire [15-1:0] node449;
	wire [15-1:0] node450;
	wire [15-1:0] node453;
	wire [15-1:0] node456;
	wire [15-1:0] node457;
	wire [15-1:0] node458;
	wire [15-1:0] node461;
	wire [15-1:0] node464;
	wire [15-1:0] node465;
	wire [15-1:0] node468;
	wire [15-1:0] node471;
	wire [15-1:0] node472;
	wire [15-1:0] node473;
	wire [15-1:0] node474;
	wire [15-1:0] node477;
	wire [15-1:0] node480;
	wire [15-1:0] node481;
	wire [15-1:0] node484;
	wire [15-1:0] node487;
	wire [15-1:0] node488;
	wire [15-1:0] node489;
	wire [15-1:0] node492;
	wire [15-1:0] node495;
	wire [15-1:0] node497;
	wire [15-1:0] node500;
	wire [15-1:0] node501;
	wire [15-1:0] node502;
	wire [15-1:0] node503;
	wire [15-1:0] node504;
	wire [15-1:0] node505;
	wire [15-1:0] node506;
	wire [15-1:0] node507;
	wire [15-1:0] node510;
	wire [15-1:0] node513;
	wire [15-1:0] node514;
	wire [15-1:0] node517;
	wire [15-1:0] node520;
	wire [15-1:0] node521;
	wire [15-1:0] node522;
	wire [15-1:0] node525;
	wire [15-1:0] node528;
	wire [15-1:0] node529;
	wire [15-1:0] node532;
	wire [15-1:0] node535;
	wire [15-1:0] node536;
	wire [15-1:0] node537;
	wire [15-1:0] node538;
	wire [15-1:0] node541;
	wire [15-1:0] node544;
	wire [15-1:0] node545;
	wire [15-1:0] node548;
	wire [15-1:0] node551;
	wire [15-1:0] node552;
	wire [15-1:0] node553;
	wire [15-1:0] node556;
	wire [15-1:0] node560;
	wire [15-1:0] node561;
	wire [15-1:0] node562;
	wire [15-1:0] node563;
	wire [15-1:0] node564;
	wire [15-1:0] node567;
	wire [15-1:0] node570;
	wire [15-1:0] node571;
	wire [15-1:0] node574;
	wire [15-1:0] node577;
	wire [15-1:0] node578;
	wire [15-1:0] node579;
	wire [15-1:0] node582;
	wire [15-1:0] node585;
	wire [15-1:0] node586;
	wire [15-1:0] node589;
	wire [15-1:0] node592;
	wire [15-1:0] node593;
	wire [15-1:0] node594;
	wire [15-1:0] node595;
	wire [15-1:0] node598;
	wire [15-1:0] node601;
	wire [15-1:0] node602;
	wire [15-1:0] node606;
	wire [15-1:0] node607;
	wire [15-1:0] node608;
	wire [15-1:0] node611;
	wire [15-1:0] node614;
	wire [15-1:0] node615;
	wire [15-1:0] node618;
	wire [15-1:0] node621;
	wire [15-1:0] node622;
	wire [15-1:0] node623;
	wire [15-1:0] node624;
	wire [15-1:0] node625;
	wire [15-1:0] node626;
	wire [15-1:0] node629;
	wire [15-1:0] node632;
	wire [15-1:0] node633;
	wire [15-1:0] node636;
	wire [15-1:0] node639;
	wire [15-1:0] node640;
	wire [15-1:0] node641;
	wire [15-1:0] node645;
	wire [15-1:0] node646;
	wire [15-1:0] node649;
	wire [15-1:0] node652;
	wire [15-1:0] node653;
	wire [15-1:0] node654;
	wire [15-1:0] node655;
	wire [15-1:0] node658;
	wire [15-1:0] node661;
	wire [15-1:0] node662;
	wire [15-1:0] node665;
	wire [15-1:0] node668;
	wire [15-1:0] node669;
	wire [15-1:0] node670;
	wire [15-1:0] node673;
	wire [15-1:0] node676;
	wire [15-1:0] node677;
	wire [15-1:0] node680;
	wire [15-1:0] node683;
	wire [15-1:0] node684;
	wire [15-1:0] node685;
	wire [15-1:0] node686;
	wire [15-1:0] node687;
	wire [15-1:0] node691;
	wire [15-1:0] node692;
	wire [15-1:0] node695;
	wire [15-1:0] node698;
	wire [15-1:0] node699;
	wire [15-1:0] node700;
	wire [15-1:0] node703;
	wire [15-1:0] node706;
	wire [15-1:0] node707;
	wire [15-1:0] node710;
	wire [15-1:0] node713;
	wire [15-1:0] node714;
	wire [15-1:0] node715;
	wire [15-1:0] node716;
	wire [15-1:0] node719;
	wire [15-1:0] node722;
	wire [15-1:0] node723;
	wire [15-1:0] node726;
	wire [15-1:0] node729;
	wire [15-1:0] node730;
	wire [15-1:0] node732;
	wire [15-1:0] node735;
	wire [15-1:0] node736;
	wire [15-1:0] node739;
	wire [15-1:0] node742;
	wire [15-1:0] node743;
	wire [15-1:0] node744;
	wire [15-1:0] node745;
	wire [15-1:0] node746;
	wire [15-1:0] node747;
	wire [15-1:0] node748;
	wire [15-1:0] node751;
	wire [15-1:0] node754;
	wire [15-1:0] node755;
	wire [15-1:0] node758;
	wire [15-1:0] node761;
	wire [15-1:0] node762;
	wire [15-1:0] node763;
	wire [15-1:0] node766;
	wire [15-1:0] node769;
	wire [15-1:0] node770;
	wire [15-1:0] node773;
	wire [15-1:0] node776;
	wire [15-1:0] node777;
	wire [15-1:0] node778;
	wire [15-1:0] node779;
	wire [15-1:0] node782;
	wire [15-1:0] node785;
	wire [15-1:0] node786;
	wire [15-1:0] node789;
	wire [15-1:0] node792;
	wire [15-1:0] node793;
	wire [15-1:0] node794;
	wire [15-1:0] node798;
	wire [15-1:0] node799;
	wire [15-1:0] node802;
	wire [15-1:0] node805;
	wire [15-1:0] node806;
	wire [15-1:0] node807;
	wire [15-1:0] node808;
	wire [15-1:0] node809;
	wire [15-1:0] node812;
	wire [15-1:0] node815;
	wire [15-1:0] node816;
	wire [15-1:0] node819;
	wire [15-1:0] node822;
	wire [15-1:0] node823;
	wire [15-1:0] node824;
	wire [15-1:0] node827;
	wire [15-1:0] node830;
	wire [15-1:0] node831;
	wire [15-1:0] node834;
	wire [15-1:0] node837;
	wire [15-1:0] node838;
	wire [15-1:0] node839;
	wire [15-1:0] node840;
	wire [15-1:0] node843;
	wire [15-1:0] node846;
	wire [15-1:0] node847;
	wire [15-1:0] node850;
	wire [15-1:0] node853;
	wire [15-1:0] node854;
	wire [15-1:0] node855;
	wire [15-1:0] node858;
	wire [15-1:0] node861;
	wire [15-1:0] node862;
	wire [15-1:0] node865;
	wire [15-1:0] node868;
	wire [15-1:0] node869;
	wire [15-1:0] node870;
	wire [15-1:0] node871;
	wire [15-1:0] node872;
	wire [15-1:0] node873;
	wire [15-1:0] node876;
	wire [15-1:0] node879;
	wire [15-1:0] node880;
	wire [15-1:0] node883;
	wire [15-1:0] node886;
	wire [15-1:0] node887;
	wire [15-1:0] node888;
	wire [15-1:0] node891;
	wire [15-1:0] node894;
	wire [15-1:0] node895;
	wire [15-1:0] node898;
	wire [15-1:0] node901;
	wire [15-1:0] node902;
	wire [15-1:0] node903;
	wire [15-1:0] node904;
	wire [15-1:0] node907;
	wire [15-1:0] node910;
	wire [15-1:0] node911;
	wire [15-1:0] node914;
	wire [15-1:0] node917;
	wire [15-1:0] node918;
	wire [15-1:0] node919;
	wire [15-1:0] node922;
	wire [15-1:0] node925;
	wire [15-1:0] node926;
	wire [15-1:0] node929;
	wire [15-1:0] node932;
	wire [15-1:0] node933;
	wire [15-1:0] node934;
	wire [15-1:0] node935;
	wire [15-1:0] node936;
	wire [15-1:0] node939;
	wire [15-1:0] node942;
	wire [15-1:0] node943;
	wire [15-1:0] node946;
	wire [15-1:0] node949;
	wire [15-1:0] node950;
	wire [15-1:0] node951;
	wire [15-1:0] node954;
	wire [15-1:0] node957;
	wire [15-1:0] node958;
	wire [15-1:0] node961;
	wire [15-1:0] node964;
	wire [15-1:0] node965;
	wire [15-1:0] node966;
	wire [15-1:0] node967;
	wire [15-1:0] node970;
	wire [15-1:0] node973;
	wire [15-1:0] node974;
	wire [15-1:0] node977;
	wire [15-1:0] node980;
	wire [15-1:0] node981;
	wire [15-1:0] node982;
	wire [15-1:0] node985;
	wire [15-1:0] node988;
	wire [15-1:0] node989;
	wire [15-1:0] node992;
	wire [15-1:0] node995;
	wire [15-1:0] node996;
	wire [15-1:0] node997;
	wire [15-1:0] node998;
	wire [15-1:0] node999;
	wire [15-1:0] node1000;
	wire [15-1:0] node1001;
	wire [15-1:0] node1002;
	wire [15-1:0] node1003;
	wire [15-1:0] node1006;
	wire [15-1:0] node1009;
	wire [15-1:0] node1010;
	wire [15-1:0] node1014;
	wire [15-1:0] node1015;
	wire [15-1:0] node1016;
	wire [15-1:0] node1019;
	wire [15-1:0] node1022;
	wire [15-1:0] node1023;
	wire [15-1:0] node1026;
	wire [15-1:0] node1029;
	wire [15-1:0] node1030;
	wire [15-1:0] node1031;
	wire [15-1:0] node1033;
	wire [15-1:0] node1036;
	wire [15-1:0] node1037;
	wire [15-1:0] node1040;
	wire [15-1:0] node1043;
	wire [15-1:0] node1044;
	wire [15-1:0] node1045;
	wire [15-1:0] node1048;
	wire [15-1:0] node1051;
	wire [15-1:0] node1052;
	wire [15-1:0] node1055;
	wire [15-1:0] node1058;
	wire [15-1:0] node1059;
	wire [15-1:0] node1060;
	wire [15-1:0] node1061;
	wire [15-1:0] node1062;
	wire [15-1:0] node1065;
	wire [15-1:0] node1068;
	wire [15-1:0] node1069;
	wire [15-1:0] node1072;
	wire [15-1:0] node1075;
	wire [15-1:0] node1076;
	wire [15-1:0] node1077;
	wire [15-1:0] node1080;
	wire [15-1:0] node1083;
	wire [15-1:0] node1084;
	wire [15-1:0] node1087;
	wire [15-1:0] node1090;
	wire [15-1:0] node1091;
	wire [15-1:0] node1092;
	wire [15-1:0] node1093;
	wire [15-1:0] node1096;
	wire [15-1:0] node1099;
	wire [15-1:0] node1100;
	wire [15-1:0] node1103;
	wire [15-1:0] node1106;
	wire [15-1:0] node1107;
	wire [15-1:0] node1108;
	wire [15-1:0] node1111;
	wire [15-1:0] node1114;
	wire [15-1:0] node1115;
	wire [15-1:0] node1119;
	wire [15-1:0] node1120;
	wire [15-1:0] node1121;
	wire [15-1:0] node1122;
	wire [15-1:0] node1123;
	wire [15-1:0] node1124;
	wire [15-1:0] node1127;
	wire [15-1:0] node1130;
	wire [15-1:0] node1131;
	wire [15-1:0] node1134;
	wire [15-1:0] node1137;
	wire [15-1:0] node1138;
	wire [15-1:0] node1139;
	wire [15-1:0] node1142;
	wire [15-1:0] node1145;
	wire [15-1:0] node1146;
	wire [15-1:0] node1149;
	wire [15-1:0] node1152;
	wire [15-1:0] node1153;
	wire [15-1:0] node1154;
	wire [15-1:0] node1155;
	wire [15-1:0] node1158;
	wire [15-1:0] node1161;
	wire [15-1:0] node1162;
	wire [15-1:0] node1165;
	wire [15-1:0] node1168;
	wire [15-1:0] node1169;
	wire [15-1:0] node1170;
	wire [15-1:0] node1173;
	wire [15-1:0] node1176;
	wire [15-1:0] node1177;
	wire [15-1:0] node1180;
	wire [15-1:0] node1183;
	wire [15-1:0] node1184;
	wire [15-1:0] node1185;
	wire [15-1:0] node1186;
	wire [15-1:0] node1189;
	wire [15-1:0] node1190;
	wire [15-1:0] node1193;
	wire [15-1:0] node1196;
	wire [15-1:0] node1197;
	wire [15-1:0] node1199;
	wire [15-1:0] node1202;
	wire [15-1:0] node1203;
	wire [15-1:0] node1206;
	wire [15-1:0] node1209;
	wire [15-1:0] node1210;
	wire [15-1:0] node1211;
	wire [15-1:0] node1212;
	wire [15-1:0] node1215;
	wire [15-1:0] node1218;
	wire [15-1:0] node1219;
	wire [15-1:0] node1222;
	wire [15-1:0] node1225;
	wire [15-1:0] node1226;
	wire [15-1:0] node1228;
	wire [15-1:0] node1231;
	wire [15-1:0] node1232;
	wire [15-1:0] node1235;
	wire [15-1:0] node1238;
	wire [15-1:0] node1239;
	wire [15-1:0] node1240;
	wire [15-1:0] node1241;
	wire [15-1:0] node1242;
	wire [15-1:0] node1243;
	wire [15-1:0] node1244;
	wire [15-1:0] node1247;
	wire [15-1:0] node1250;
	wire [15-1:0] node1251;
	wire [15-1:0] node1254;
	wire [15-1:0] node1257;
	wire [15-1:0] node1258;
	wire [15-1:0] node1259;
	wire [15-1:0] node1262;
	wire [15-1:0] node1265;
	wire [15-1:0] node1266;
	wire [15-1:0] node1269;
	wire [15-1:0] node1272;
	wire [15-1:0] node1273;
	wire [15-1:0] node1274;
	wire [15-1:0] node1275;
	wire [15-1:0] node1279;
	wire [15-1:0] node1280;
	wire [15-1:0] node1283;
	wire [15-1:0] node1286;
	wire [15-1:0] node1287;
	wire [15-1:0] node1288;
	wire [15-1:0] node1291;
	wire [15-1:0] node1294;
	wire [15-1:0] node1295;
	wire [15-1:0] node1299;
	wire [15-1:0] node1300;
	wire [15-1:0] node1301;
	wire [15-1:0] node1302;
	wire [15-1:0] node1303;
	wire [15-1:0] node1306;
	wire [15-1:0] node1309;
	wire [15-1:0] node1310;
	wire [15-1:0] node1314;
	wire [15-1:0] node1315;
	wire [15-1:0] node1317;
	wire [15-1:0] node1320;
	wire [15-1:0] node1321;
	wire [15-1:0] node1324;
	wire [15-1:0] node1327;
	wire [15-1:0] node1328;
	wire [15-1:0] node1329;
	wire [15-1:0] node1330;
	wire [15-1:0] node1333;
	wire [15-1:0] node1336;
	wire [15-1:0] node1337;
	wire [15-1:0] node1340;
	wire [15-1:0] node1343;
	wire [15-1:0] node1344;
	wire [15-1:0] node1346;
	wire [15-1:0] node1349;
	wire [15-1:0] node1350;
	wire [15-1:0] node1353;
	wire [15-1:0] node1356;
	wire [15-1:0] node1357;
	wire [15-1:0] node1358;
	wire [15-1:0] node1359;
	wire [15-1:0] node1360;
	wire [15-1:0] node1361;
	wire [15-1:0] node1365;
	wire [15-1:0] node1367;
	wire [15-1:0] node1370;
	wire [15-1:0] node1371;
	wire [15-1:0] node1372;
	wire [15-1:0] node1375;
	wire [15-1:0] node1378;
	wire [15-1:0] node1379;
	wire [15-1:0] node1382;
	wire [15-1:0] node1385;
	wire [15-1:0] node1386;
	wire [15-1:0] node1387;
	wire [15-1:0] node1388;
	wire [15-1:0] node1391;
	wire [15-1:0] node1394;
	wire [15-1:0] node1395;
	wire [15-1:0] node1398;
	wire [15-1:0] node1401;
	wire [15-1:0] node1402;
	wire [15-1:0] node1403;
	wire [15-1:0] node1406;
	wire [15-1:0] node1409;
	wire [15-1:0] node1410;
	wire [15-1:0] node1413;
	wire [15-1:0] node1416;
	wire [15-1:0] node1417;
	wire [15-1:0] node1418;
	wire [15-1:0] node1419;
	wire [15-1:0] node1421;
	wire [15-1:0] node1425;
	wire [15-1:0] node1426;
	wire [15-1:0] node1427;
	wire [15-1:0] node1430;
	wire [15-1:0] node1433;
	wire [15-1:0] node1434;
	wire [15-1:0] node1437;
	wire [15-1:0] node1440;
	wire [15-1:0] node1441;
	wire [15-1:0] node1442;
	wire [15-1:0] node1443;
	wire [15-1:0] node1446;
	wire [15-1:0] node1449;
	wire [15-1:0] node1450;
	wire [15-1:0] node1453;
	wire [15-1:0] node1456;
	wire [15-1:0] node1457;
	wire [15-1:0] node1458;
	wire [15-1:0] node1461;
	wire [15-1:0] node1464;
	wire [15-1:0] node1466;
	wire [15-1:0] node1469;
	wire [15-1:0] node1470;
	wire [15-1:0] node1471;
	wire [15-1:0] node1472;
	wire [15-1:0] node1473;
	wire [15-1:0] node1474;
	wire [15-1:0] node1475;
	wire [15-1:0] node1476;
	wire [15-1:0] node1479;
	wire [15-1:0] node1482;
	wire [15-1:0] node1483;
	wire [15-1:0] node1486;
	wire [15-1:0] node1489;
	wire [15-1:0] node1490;
	wire [15-1:0] node1491;
	wire [15-1:0] node1494;
	wire [15-1:0] node1497;
	wire [15-1:0] node1498;
	wire [15-1:0] node1501;
	wire [15-1:0] node1504;
	wire [15-1:0] node1505;
	wire [15-1:0] node1506;
	wire [15-1:0] node1507;
	wire [15-1:0] node1510;
	wire [15-1:0] node1513;
	wire [15-1:0] node1514;
	wire [15-1:0] node1517;
	wire [15-1:0] node1520;
	wire [15-1:0] node1522;
	wire [15-1:0] node1523;
	wire [15-1:0] node1526;
	wire [15-1:0] node1529;
	wire [15-1:0] node1530;
	wire [15-1:0] node1531;
	wire [15-1:0] node1532;
	wire [15-1:0] node1533;
	wire [15-1:0] node1536;
	wire [15-1:0] node1539;
	wire [15-1:0] node1540;
	wire [15-1:0] node1543;
	wire [15-1:0] node1546;
	wire [15-1:0] node1547;
	wire [15-1:0] node1548;
	wire [15-1:0] node1551;
	wire [15-1:0] node1554;
	wire [15-1:0] node1555;
	wire [15-1:0] node1558;
	wire [15-1:0] node1561;
	wire [15-1:0] node1562;
	wire [15-1:0] node1563;
	wire [15-1:0] node1564;
	wire [15-1:0] node1568;
	wire [15-1:0] node1569;
	wire [15-1:0] node1572;
	wire [15-1:0] node1575;
	wire [15-1:0] node1576;
	wire [15-1:0] node1577;
	wire [15-1:0] node1581;
	wire [15-1:0] node1582;
	wire [15-1:0] node1585;
	wire [15-1:0] node1588;
	wire [15-1:0] node1589;
	wire [15-1:0] node1590;
	wire [15-1:0] node1591;
	wire [15-1:0] node1592;
	wire [15-1:0] node1593;
	wire [15-1:0] node1596;
	wire [15-1:0] node1599;
	wire [15-1:0] node1600;
	wire [15-1:0] node1603;
	wire [15-1:0] node1606;
	wire [15-1:0] node1607;
	wire [15-1:0] node1608;
	wire [15-1:0] node1611;
	wire [15-1:0] node1614;
	wire [15-1:0] node1615;
	wire [15-1:0] node1618;
	wire [15-1:0] node1621;
	wire [15-1:0] node1622;
	wire [15-1:0] node1623;
	wire [15-1:0] node1625;
	wire [15-1:0] node1628;
	wire [15-1:0] node1629;
	wire [15-1:0] node1632;
	wire [15-1:0] node1635;
	wire [15-1:0] node1636;
	wire [15-1:0] node1637;
	wire [15-1:0] node1640;
	wire [15-1:0] node1643;
	wire [15-1:0] node1645;
	wire [15-1:0] node1648;
	wire [15-1:0] node1649;
	wire [15-1:0] node1650;
	wire [15-1:0] node1651;
	wire [15-1:0] node1652;
	wire [15-1:0] node1655;
	wire [15-1:0] node1658;
	wire [15-1:0] node1659;
	wire [15-1:0] node1662;
	wire [15-1:0] node1665;
	wire [15-1:0] node1666;
	wire [15-1:0] node1668;
	wire [15-1:0] node1671;
	wire [15-1:0] node1672;
	wire [15-1:0] node1675;
	wire [15-1:0] node1678;
	wire [15-1:0] node1679;
	wire [15-1:0] node1680;
	wire [15-1:0] node1681;
	wire [15-1:0] node1684;
	wire [15-1:0] node1687;
	wire [15-1:0] node1688;
	wire [15-1:0] node1691;
	wire [15-1:0] node1694;
	wire [15-1:0] node1695;
	wire [15-1:0] node1697;
	wire [15-1:0] node1700;
	wire [15-1:0] node1702;
	wire [15-1:0] node1705;
	wire [15-1:0] node1706;
	wire [15-1:0] node1707;
	wire [15-1:0] node1708;
	wire [15-1:0] node1709;
	wire [15-1:0] node1710;
	wire [15-1:0] node1711;
	wire [15-1:0] node1714;
	wire [15-1:0] node1717;
	wire [15-1:0] node1718;
	wire [15-1:0] node1721;
	wire [15-1:0] node1724;
	wire [15-1:0] node1725;
	wire [15-1:0] node1726;
	wire [15-1:0] node1729;
	wire [15-1:0] node1732;
	wire [15-1:0] node1733;
	wire [15-1:0] node1736;
	wire [15-1:0] node1739;
	wire [15-1:0] node1740;
	wire [15-1:0] node1741;
	wire [15-1:0] node1742;
	wire [15-1:0] node1745;
	wire [15-1:0] node1748;
	wire [15-1:0] node1749;
	wire [15-1:0] node1752;
	wire [15-1:0] node1755;
	wire [15-1:0] node1756;
	wire [15-1:0] node1757;
	wire [15-1:0] node1760;
	wire [15-1:0] node1763;
	wire [15-1:0] node1764;
	wire [15-1:0] node1767;
	wire [15-1:0] node1770;
	wire [15-1:0] node1771;
	wire [15-1:0] node1772;
	wire [15-1:0] node1773;
	wire [15-1:0] node1774;
	wire [15-1:0] node1777;
	wire [15-1:0] node1780;
	wire [15-1:0] node1781;
	wire [15-1:0] node1784;
	wire [15-1:0] node1787;
	wire [15-1:0] node1788;
	wire [15-1:0] node1789;
	wire [15-1:0] node1792;
	wire [15-1:0] node1795;
	wire [15-1:0] node1796;
	wire [15-1:0] node1799;
	wire [15-1:0] node1802;
	wire [15-1:0] node1803;
	wire [15-1:0] node1804;
	wire [15-1:0] node1805;
	wire [15-1:0] node1808;
	wire [15-1:0] node1811;
	wire [15-1:0] node1812;
	wire [15-1:0] node1815;
	wire [15-1:0] node1818;
	wire [15-1:0] node1819;
	wire [15-1:0] node1820;
	wire [15-1:0] node1823;
	wire [15-1:0] node1826;
	wire [15-1:0] node1827;
	wire [15-1:0] node1830;
	wire [15-1:0] node1833;
	wire [15-1:0] node1834;
	wire [15-1:0] node1835;
	wire [15-1:0] node1836;
	wire [15-1:0] node1837;
	wire [15-1:0] node1838;
	wire [15-1:0] node1841;
	wire [15-1:0] node1844;
	wire [15-1:0] node1845;
	wire [15-1:0] node1848;
	wire [15-1:0] node1851;
	wire [15-1:0] node1852;
	wire [15-1:0] node1853;
	wire [15-1:0] node1856;
	wire [15-1:0] node1859;
	wire [15-1:0] node1860;
	wire [15-1:0] node1863;
	wire [15-1:0] node1866;
	wire [15-1:0] node1867;
	wire [15-1:0] node1868;
	wire [15-1:0] node1869;
	wire [15-1:0] node1872;
	wire [15-1:0] node1875;
	wire [15-1:0] node1877;
	wire [15-1:0] node1880;
	wire [15-1:0] node1881;
	wire [15-1:0] node1882;
	wire [15-1:0] node1885;
	wire [15-1:0] node1888;
	wire [15-1:0] node1889;
	wire [15-1:0] node1892;
	wire [15-1:0] node1895;
	wire [15-1:0] node1896;
	wire [15-1:0] node1897;
	wire [15-1:0] node1898;
	wire [15-1:0] node1899;
	wire [15-1:0] node1902;
	wire [15-1:0] node1905;
	wire [15-1:0] node1906;
	wire [15-1:0] node1909;
	wire [15-1:0] node1912;
	wire [15-1:0] node1913;
	wire [15-1:0] node1914;
	wire [15-1:0] node1918;
	wire [15-1:0] node1920;
	wire [15-1:0] node1923;
	wire [15-1:0] node1924;
	wire [15-1:0] node1925;
	wire [15-1:0] node1927;
	wire [15-1:0] node1930;
	wire [15-1:0] node1931;
	wire [15-1:0] node1934;
	wire [15-1:0] node1937;
	wire [15-1:0] node1938;
	wire [15-1:0] node1939;
	wire [15-1:0] node1942;
	wire [15-1:0] node1945;
	wire [15-1:0] node1946;
	wire [15-1:0] node1949;
	wire [15-1:0] node1952;
	wire [15-1:0] node1953;
	wire [15-1:0] node1954;
	wire [15-1:0] node1955;
	wire [15-1:0] node1956;
	wire [15-1:0] node1957;
	wire [15-1:0] node1958;
	wire [15-1:0] node1959;
	wire [15-1:0] node1960;
	wire [15-1:0] node1961;
	wire [15-1:0] node1964;
	wire [15-1:0] node1967;
	wire [15-1:0] node1968;
	wire [15-1:0] node1971;
	wire [15-1:0] node1974;
	wire [15-1:0] node1975;
	wire [15-1:0] node1976;
	wire [15-1:0] node1979;
	wire [15-1:0] node1982;
	wire [15-1:0] node1983;
	wire [15-1:0] node1986;
	wire [15-1:0] node1989;
	wire [15-1:0] node1990;
	wire [15-1:0] node1991;
	wire [15-1:0] node1992;
	wire [15-1:0] node1995;
	wire [15-1:0] node1998;
	wire [15-1:0] node1999;
	wire [15-1:0] node2002;
	wire [15-1:0] node2005;
	wire [15-1:0] node2006;
	wire [15-1:0] node2007;
	wire [15-1:0] node2010;
	wire [15-1:0] node2013;
	wire [15-1:0] node2014;
	wire [15-1:0] node2018;
	wire [15-1:0] node2019;
	wire [15-1:0] node2020;
	wire [15-1:0] node2021;
	wire [15-1:0] node2022;
	wire [15-1:0] node2025;
	wire [15-1:0] node2028;
	wire [15-1:0] node2029;
	wire [15-1:0] node2032;
	wire [15-1:0] node2035;
	wire [15-1:0] node2036;
	wire [15-1:0] node2037;
	wire [15-1:0] node2040;
	wire [15-1:0] node2043;
	wire [15-1:0] node2044;
	wire [15-1:0] node2047;
	wire [15-1:0] node2050;
	wire [15-1:0] node2051;
	wire [15-1:0] node2052;
	wire [15-1:0] node2053;
	wire [15-1:0] node2056;
	wire [15-1:0] node2059;
	wire [15-1:0] node2060;
	wire [15-1:0] node2063;
	wire [15-1:0] node2066;
	wire [15-1:0] node2067;
	wire [15-1:0] node2068;
	wire [15-1:0] node2071;
	wire [15-1:0] node2075;
	wire [15-1:0] node2076;
	wire [15-1:0] node2077;
	wire [15-1:0] node2078;
	wire [15-1:0] node2079;
	wire [15-1:0] node2080;
	wire [15-1:0] node2083;
	wire [15-1:0] node2086;
	wire [15-1:0] node2087;
	wire [15-1:0] node2090;
	wire [15-1:0] node2093;
	wire [15-1:0] node2094;
	wire [15-1:0] node2095;
	wire [15-1:0] node2098;
	wire [15-1:0] node2101;
	wire [15-1:0] node2102;
	wire [15-1:0] node2105;
	wire [15-1:0] node2108;
	wire [15-1:0] node2109;
	wire [15-1:0] node2110;
	wire [15-1:0] node2111;
	wire [15-1:0] node2114;
	wire [15-1:0] node2117;
	wire [15-1:0] node2118;
	wire [15-1:0] node2122;
	wire [15-1:0] node2123;
	wire [15-1:0] node2124;
	wire [15-1:0] node2127;
	wire [15-1:0] node2130;
	wire [15-1:0] node2131;
	wire [15-1:0] node2134;
	wire [15-1:0] node2137;
	wire [15-1:0] node2138;
	wire [15-1:0] node2139;
	wire [15-1:0] node2140;
	wire [15-1:0] node2141;
	wire [15-1:0] node2144;
	wire [15-1:0] node2147;
	wire [15-1:0] node2148;
	wire [15-1:0] node2151;
	wire [15-1:0] node2154;
	wire [15-1:0] node2155;
	wire [15-1:0] node2156;
	wire [15-1:0] node2160;
	wire [15-1:0] node2161;
	wire [15-1:0] node2164;
	wire [15-1:0] node2167;
	wire [15-1:0] node2168;
	wire [15-1:0] node2169;
	wire [15-1:0] node2170;
	wire [15-1:0] node2174;
	wire [15-1:0] node2175;
	wire [15-1:0] node2178;
	wire [15-1:0] node2181;
	wire [15-1:0] node2182;
	wire [15-1:0] node2183;
	wire [15-1:0] node2186;
	wire [15-1:0] node2189;
	wire [15-1:0] node2190;
	wire [15-1:0] node2193;
	wire [15-1:0] node2196;
	wire [15-1:0] node2197;
	wire [15-1:0] node2198;
	wire [15-1:0] node2199;
	wire [15-1:0] node2200;
	wire [15-1:0] node2201;
	wire [15-1:0] node2202;
	wire [15-1:0] node2205;
	wire [15-1:0] node2208;
	wire [15-1:0] node2209;
	wire [15-1:0] node2213;
	wire [15-1:0] node2214;
	wire [15-1:0] node2215;
	wire [15-1:0] node2218;
	wire [15-1:0] node2221;
	wire [15-1:0] node2222;
	wire [15-1:0] node2226;
	wire [15-1:0] node2227;
	wire [15-1:0] node2228;
	wire [15-1:0] node2229;
	wire [15-1:0] node2232;
	wire [15-1:0] node2235;
	wire [15-1:0] node2236;
	wire [15-1:0] node2239;
	wire [15-1:0] node2242;
	wire [15-1:0] node2243;
	wire [15-1:0] node2244;
	wire [15-1:0] node2247;
	wire [15-1:0] node2250;
	wire [15-1:0] node2251;
	wire [15-1:0] node2254;
	wire [15-1:0] node2257;
	wire [15-1:0] node2258;
	wire [15-1:0] node2259;
	wire [15-1:0] node2260;
	wire [15-1:0] node2261;
	wire [15-1:0] node2265;
	wire [15-1:0] node2266;
	wire [15-1:0] node2269;
	wire [15-1:0] node2272;
	wire [15-1:0] node2273;
	wire [15-1:0] node2274;
	wire [15-1:0] node2277;
	wire [15-1:0] node2280;
	wire [15-1:0] node2281;
	wire [15-1:0] node2284;
	wire [15-1:0] node2287;
	wire [15-1:0] node2288;
	wire [15-1:0] node2289;
	wire [15-1:0] node2290;
	wire [15-1:0] node2293;
	wire [15-1:0] node2296;
	wire [15-1:0] node2297;
	wire [15-1:0] node2300;
	wire [15-1:0] node2303;
	wire [15-1:0] node2304;
	wire [15-1:0] node2305;
	wire [15-1:0] node2308;
	wire [15-1:0] node2311;
	wire [15-1:0] node2312;
	wire [15-1:0] node2315;
	wire [15-1:0] node2318;
	wire [15-1:0] node2319;
	wire [15-1:0] node2320;
	wire [15-1:0] node2321;
	wire [15-1:0] node2322;
	wire [15-1:0] node2323;
	wire [15-1:0] node2326;
	wire [15-1:0] node2329;
	wire [15-1:0] node2330;
	wire [15-1:0] node2333;
	wire [15-1:0] node2336;
	wire [15-1:0] node2337;
	wire [15-1:0] node2338;
	wire [15-1:0] node2341;
	wire [15-1:0] node2344;
	wire [15-1:0] node2345;
	wire [15-1:0] node2348;
	wire [15-1:0] node2351;
	wire [15-1:0] node2352;
	wire [15-1:0] node2353;
	wire [15-1:0] node2354;
	wire [15-1:0] node2357;
	wire [15-1:0] node2360;
	wire [15-1:0] node2361;
	wire [15-1:0] node2364;
	wire [15-1:0] node2367;
	wire [15-1:0] node2368;
	wire [15-1:0] node2369;
	wire [15-1:0] node2372;
	wire [15-1:0] node2375;
	wire [15-1:0] node2376;
	wire [15-1:0] node2380;
	wire [15-1:0] node2381;
	wire [15-1:0] node2382;
	wire [15-1:0] node2383;
	wire [15-1:0] node2384;
	wire [15-1:0] node2387;
	wire [15-1:0] node2390;
	wire [15-1:0] node2391;
	wire [15-1:0] node2394;
	wire [15-1:0] node2397;
	wire [15-1:0] node2398;
	wire [15-1:0] node2399;
	wire [15-1:0] node2402;
	wire [15-1:0] node2405;
	wire [15-1:0] node2407;
	wire [15-1:0] node2410;
	wire [15-1:0] node2411;
	wire [15-1:0] node2412;
	wire [15-1:0] node2413;
	wire [15-1:0] node2416;
	wire [15-1:0] node2419;
	wire [15-1:0] node2420;
	wire [15-1:0] node2423;
	wire [15-1:0] node2426;
	wire [15-1:0] node2427;
	wire [15-1:0] node2428;
	wire [15-1:0] node2431;
	wire [15-1:0] node2434;
	wire [15-1:0] node2435;
	wire [15-1:0] node2438;
	wire [15-1:0] node2441;
	wire [15-1:0] node2442;
	wire [15-1:0] node2443;
	wire [15-1:0] node2444;
	wire [15-1:0] node2445;
	wire [15-1:0] node2446;
	wire [15-1:0] node2447;
	wire [15-1:0] node2448;
	wire [15-1:0] node2451;
	wire [15-1:0] node2454;
	wire [15-1:0] node2455;
	wire [15-1:0] node2458;
	wire [15-1:0] node2461;
	wire [15-1:0] node2462;
	wire [15-1:0] node2463;
	wire [15-1:0] node2466;
	wire [15-1:0] node2469;
	wire [15-1:0] node2470;
	wire [15-1:0] node2473;
	wire [15-1:0] node2476;
	wire [15-1:0] node2477;
	wire [15-1:0] node2478;
	wire [15-1:0] node2479;
	wire [15-1:0] node2482;
	wire [15-1:0] node2485;
	wire [15-1:0] node2486;
	wire [15-1:0] node2490;
	wire [15-1:0] node2491;
	wire [15-1:0] node2492;
	wire [15-1:0] node2495;
	wire [15-1:0] node2498;
	wire [15-1:0] node2501;
	wire [15-1:0] node2502;
	wire [15-1:0] node2503;
	wire [15-1:0] node2504;
	wire [15-1:0] node2505;
	wire [15-1:0] node2508;
	wire [15-1:0] node2511;
	wire [15-1:0] node2512;
	wire [15-1:0] node2515;
	wire [15-1:0] node2518;
	wire [15-1:0] node2519;
	wire [15-1:0] node2520;
	wire [15-1:0] node2524;
	wire [15-1:0] node2525;
	wire [15-1:0] node2528;
	wire [15-1:0] node2531;
	wire [15-1:0] node2532;
	wire [15-1:0] node2533;
	wire [15-1:0] node2534;
	wire [15-1:0] node2537;
	wire [15-1:0] node2540;
	wire [15-1:0] node2541;
	wire [15-1:0] node2545;
	wire [15-1:0] node2546;
	wire [15-1:0] node2547;
	wire [15-1:0] node2550;
	wire [15-1:0] node2553;
	wire [15-1:0] node2554;
	wire [15-1:0] node2557;
	wire [15-1:0] node2560;
	wire [15-1:0] node2561;
	wire [15-1:0] node2562;
	wire [15-1:0] node2563;
	wire [15-1:0] node2564;
	wire [15-1:0] node2565;
	wire [15-1:0] node2568;
	wire [15-1:0] node2571;
	wire [15-1:0] node2572;
	wire [15-1:0] node2576;
	wire [15-1:0] node2577;
	wire [15-1:0] node2578;
	wire [15-1:0] node2581;
	wire [15-1:0] node2584;
	wire [15-1:0] node2585;
	wire [15-1:0] node2588;
	wire [15-1:0] node2591;
	wire [15-1:0] node2592;
	wire [15-1:0] node2593;
	wire [15-1:0] node2594;
	wire [15-1:0] node2597;
	wire [15-1:0] node2600;
	wire [15-1:0] node2601;
	wire [15-1:0] node2604;
	wire [15-1:0] node2607;
	wire [15-1:0] node2608;
	wire [15-1:0] node2609;
	wire [15-1:0] node2612;
	wire [15-1:0] node2615;
	wire [15-1:0] node2616;
	wire [15-1:0] node2619;
	wire [15-1:0] node2622;
	wire [15-1:0] node2623;
	wire [15-1:0] node2624;
	wire [15-1:0] node2625;
	wire [15-1:0] node2626;
	wire [15-1:0] node2629;
	wire [15-1:0] node2632;
	wire [15-1:0] node2633;
	wire [15-1:0] node2636;
	wire [15-1:0] node2639;
	wire [15-1:0] node2640;
	wire [15-1:0] node2641;
	wire [15-1:0] node2644;
	wire [15-1:0] node2647;
	wire [15-1:0] node2648;
	wire [15-1:0] node2652;
	wire [15-1:0] node2653;
	wire [15-1:0] node2654;
	wire [15-1:0] node2655;
	wire [15-1:0] node2659;
	wire [15-1:0] node2660;
	wire [15-1:0] node2663;
	wire [15-1:0] node2666;
	wire [15-1:0] node2667;
	wire [15-1:0] node2668;
	wire [15-1:0] node2671;
	wire [15-1:0] node2674;
	wire [15-1:0] node2675;
	wire [15-1:0] node2678;
	wire [15-1:0] node2681;
	wire [15-1:0] node2682;
	wire [15-1:0] node2683;
	wire [15-1:0] node2684;
	wire [15-1:0] node2685;
	wire [15-1:0] node2686;
	wire [15-1:0] node2687;
	wire [15-1:0] node2690;
	wire [15-1:0] node2693;
	wire [15-1:0] node2694;
	wire [15-1:0] node2697;
	wire [15-1:0] node2700;
	wire [15-1:0] node2701;
	wire [15-1:0] node2702;
	wire [15-1:0] node2705;
	wire [15-1:0] node2708;
	wire [15-1:0] node2710;
	wire [15-1:0] node2713;
	wire [15-1:0] node2714;
	wire [15-1:0] node2715;
	wire [15-1:0] node2716;
	wire [15-1:0] node2719;
	wire [15-1:0] node2722;
	wire [15-1:0] node2723;
	wire [15-1:0] node2726;
	wire [15-1:0] node2729;
	wire [15-1:0] node2730;
	wire [15-1:0] node2732;
	wire [15-1:0] node2735;
	wire [15-1:0] node2736;
	wire [15-1:0] node2739;
	wire [15-1:0] node2742;
	wire [15-1:0] node2743;
	wire [15-1:0] node2744;
	wire [15-1:0] node2745;
	wire [15-1:0] node2746;
	wire [15-1:0] node2749;
	wire [15-1:0] node2752;
	wire [15-1:0] node2753;
	wire [15-1:0] node2756;
	wire [15-1:0] node2759;
	wire [15-1:0] node2760;
	wire [15-1:0] node2761;
	wire [15-1:0] node2764;
	wire [15-1:0] node2767;
	wire [15-1:0] node2768;
	wire [15-1:0] node2771;
	wire [15-1:0] node2774;
	wire [15-1:0] node2775;
	wire [15-1:0] node2776;
	wire [15-1:0] node2777;
	wire [15-1:0] node2780;
	wire [15-1:0] node2783;
	wire [15-1:0] node2784;
	wire [15-1:0] node2787;
	wire [15-1:0] node2790;
	wire [15-1:0] node2791;
	wire [15-1:0] node2792;
	wire [15-1:0] node2795;
	wire [15-1:0] node2798;
	wire [15-1:0] node2800;
	wire [15-1:0] node2803;
	wire [15-1:0] node2804;
	wire [15-1:0] node2805;
	wire [15-1:0] node2806;
	wire [15-1:0] node2807;
	wire [15-1:0] node2808;
	wire [15-1:0] node2812;
	wire [15-1:0] node2813;
	wire [15-1:0] node2816;
	wire [15-1:0] node2819;
	wire [15-1:0] node2820;
	wire [15-1:0] node2821;
	wire [15-1:0] node2824;
	wire [15-1:0] node2827;
	wire [15-1:0] node2828;
	wire [15-1:0] node2831;
	wire [15-1:0] node2834;
	wire [15-1:0] node2835;
	wire [15-1:0] node2836;
	wire [15-1:0] node2837;
	wire [15-1:0] node2841;
	wire [15-1:0] node2842;
	wire [15-1:0] node2846;
	wire [15-1:0] node2847;
	wire [15-1:0] node2848;
	wire [15-1:0] node2851;
	wire [15-1:0] node2854;
	wire [15-1:0] node2855;
	wire [15-1:0] node2858;
	wire [15-1:0] node2861;
	wire [15-1:0] node2862;
	wire [15-1:0] node2863;
	wire [15-1:0] node2864;
	wire [15-1:0] node2866;
	wire [15-1:0] node2869;
	wire [15-1:0] node2870;
	wire [15-1:0] node2873;
	wire [15-1:0] node2876;
	wire [15-1:0] node2877;
	wire [15-1:0] node2878;
	wire [15-1:0] node2881;
	wire [15-1:0] node2884;
	wire [15-1:0] node2885;
	wire [15-1:0] node2888;
	wire [15-1:0] node2891;
	wire [15-1:0] node2892;
	wire [15-1:0] node2893;
	wire [15-1:0] node2894;
	wire [15-1:0] node2897;
	wire [15-1:0] node2900;
	wire [15-1:0] node2901;
	wire [15-1:0] node2904;
	wire [15-1:0] node2907;
	wire [15-1:0] node2908;
	wire [15-1:0] node2909;
	wire [15-1:0] node2912;
	wire [15-1:0] node2915;
	wire [15-1:0] node2916;
	wire [15-1:0] node2919;
	wire [15-1:0] node2922;
	wire [15-1:0] node2923;
	wire [15-1:0] node2924;
	wire [15-1:0] node2925;
	wire [15-1:0] node2926;
	wire [15-1:0] node2927;
	wire [15-1:0] node2928;
	wire [15-1:0] node2929;
	wire [15-1:0] node2930;
	wire [15-1:0] node2933;
	wire [15-1:0] node2936;
	wire [15-1:0] node2937;
	wire [15-1:0] node2941;
	wire [15-1:0] node2942;
	wire [15-1:0] node2943;
	wire [15-1:0] node2946;
	wire [15-1:0] node2949;
	wire [15-1:0] node2950;
	wire [15-1:0] node2954;
	wire [15-1:0] node2955;
	wire [15-1:0] node2956;
	wire [15-1:0] node2958;
	wire [15-1:0] node2962;
	wire [15-1:0] node2963;
	wire [15-1:0] node2965;
	wire [15-1:0] node2968;
	wire [15-1:0] node2969;
	wire [15-1:0] node2972;
	wire [15-1:0] node2975;
	wire [15-1:0] node2976;
	wire [15-1:0] node2977;
	wire [15-1:0] node2978;
	wire [15-1:0] node2979;
	wire [15-1:0] node2982;
	wire [15-1:0] node2985;
	wire [15-1:0] node2986;
	wire [15-1:0] node2989;
	wire [15-1:0] node2992;
	wire [15-1:0] node2993;
	wire [15-1:0] node2994;
	wire [15-1:0] node2997;
	wire [15-1:0] node3000;
	wire [15-1:0] node3001;
	wire [15-1:0] node3004;
	wire [15-1:0] node3007;
	wire [15-1:0] node3008;
	wire [15-1:0] node3009;
	wire [15-1:0] node3010;
	wire [15-1:0] node3013;
	wire [15-1:0] node3016;
	wire [15-1:0] node3017;
	wire [15-1:0] node3020;
	wire [15-1:0] node3023;
	wire [15-1:0] node3024;
	wire [15-1:0] node3025;
	wire [15-1:0] node3028;
	wire [15-1:0] node3031;
	wire [15-1:0] node3033;
	wire [15-1:0] node3036;
	wire [15-1:0] node3037;
	wire [15-1:0] node3038;
	wire [15-1:0] node3039;
	wire [15-1:0] node3040;
	wire [15-1:0] node3041;
	wire [15-1:0] node3044;
	wire [15-1:0] node3047;
	wire [15-1:0] node3048;
	wire [15-1:0] node3051;
	wire [15-1:0] node3054;
	wire [15-1:0] node3055;
	wire [15-1:0] node3056;
	wire [15-1:0] node3059;
	wire [15-1:0] node3063;
	wire [15-1:0] node3064;
	wire [15-1:0] node3065;
	wire [15-1:0] node3066;
	wire [15-1:0] node3069;
	wire [15-1:0] node3072;
	wire [15-1:0] node3073;
	wire [15-1:0] node3077;
	wire [15-1:0] node3078;
	wire [15-1:0] node3080;
	wire [15-1:0] node3083;
	wire [15-1:0] node3084;
	wire [15-1:0] node3087;
	wire [15-1:0] node3090;
	wire [15-1:0] node3091;
	wire [15-1:0] node3092;
	wire [15-1:0] node3093;
	wire [15-1:0] node3094;
	wire [15-1:0] node3097;
	wire [15-1:0] node3100;
	wire [15-1:0] node3101;
	wire [15-1:0] node3105;
	wire [15-1:0] node3106;
	wire [15-1:0] node3107;
	wire [15-1:0] node3110;
	wire [15-1:0] node3113;
	wire [15-1:0] node3114;
	wire [15-1:0] node3118;
	wire [15-1:0] node3119;
	wire [15-1:0] node3120;
	wire [15-1:0] node3121;
	wire [15-1:0] node3124;
	wire [15-1:0] node3127;
	wire [15-1:0] node3128;
	wire [15-1:0] node3131;
	wire [15-1:0] node3134;
	wire [15-1:0] node3135;
	wire [15-1:0] node3137;
	wire [15-1:0] node3140;
	wire [15-1:0] node3142;
	wire [15-1:0] node3145;
	wire [15-1:0] node3146;
	wire [15-1:0] node3147;
	wire [15-1:0] node3148;
	wire [15-1:0] node3149;
	wire [15-1:0] node3150;
	wire [15-1:0] node3151;
	wire [15-1:0] node3154;
	wire [15-1:0] node3157;
	wire [15-1:0] node3158;
	wire [15-1:0] node3161;
	wire [15-1:0] node3164;
	wire [15-1:0] node3165;
	wire [15-1:0] node3166;
	wire [15-1:0] node3169;
	wire [15-1:0] node3172;
	wire [15-1:0] node3173;
	wire [15-1:0] node3176;
	wire [15-1:0] node3179;
	wire [15-1:0] node3180;
	wire [15-1:0] node3181;
	wire [15-1:0] node3182;
	wire [15-1:0] node3185;
	wire [15-1:0] node3188;
	wire [15-1:0] node3189;
	wire [15-1:0] node3192;
	wire [15-1:0] node3195;
	wire [15-1:0] node3196;
	wire [15-1:0] node3197;
	wire [15-1:0] node3200;
	wire [15-1:0] node3203;
	wire [15-1:0] node3204;
	wire [15-1:0] node3207;
	wire [15-1:0] node3210;
	wire [15-1:0] node3211;
	wire [15-1:0] node3212;
	wire [15-1:0] node3213;
	wire [15-1:0] node3214;
	wire [15-1:0] node3217;
	wire [15-1:0] node3220;
	wire [15-1:0] node3221;
	wire [15-1:0] node3224;
	wire [15-1:0] node3227;
	wire [15-1:0] node3228;
	wire [15-1:0] node3229;
	wire [15-1:0] node3232;
	wire [15-1:0] node3235;
	wire [15-1:0] node3236;
	wire [15-1:0] node3239;
	wire [15-1:0] node3242;
	wire [15-1:0] node3243;
	wire [15-1:0] node3244;
	wire [15-1:0] node3245;
	wire [15-1:0] node3248;
	wire [15-1:0] node3251;
	wire [15-1:0] node3252;
	wire [15-1:0] node3255;
	wire [15-1:0] node3258;
	wire [15-1:0] node3259;
	wire [15-1:0] node3260;
	wire [15-1:0] node3263;
	wire [15-1:0] node3266;
	wire [15-1:0] node3267;
	wire [15-1:0] node3270;
	wire [15-1:0] node3273;
	wire [15-1:0] node3274;
	wire [15-1:0] node3275;
	wire [15-1:0] node3276;
	wire [15-1:0] node3277;
	wire [15-1:0] node3278;
	wire [15-1:0] node3281;
	wire [15-1:0] node3284;
	wire [15-1:0] node3285;
	wire [15-1:0] node3288;
	wire [15-1:0] node3291;
	wire [15-1:0] node3292;
	wire [15-1:0] node3293;
	wire [15-1:0] node3296;
	wire [15-1:0] node3299;
	wire [15-1:0] node3300;
	wire [15-1:0] node3303;
	wire [15-1:0] node3306;
	wire [15-1:0] node3307;
	wire [15-1:0] node3308;
	wire [15-1:0] node3310;
	wire [15-1:0] node3313;
	wire [15-1:0] node3314;
	wire [15-1:0] node3317;
	wire [15-1:0] node3320;
	wire [15-1:0] node3321;
	wire [15-1:0] node3322;
	wire [15-1:0] node3325;
	wire [15-1:0] node3328;
	wire [15-1:0] node3329;
	wire [15-1:0] node3332;
	wire [15-1:0] node3335;
	wire [15-1:0] node3336;
	wire [15-1:0] node3337;
	wire [15-1:0] node3338;
	wire [15-1:0] node3339;
	wire [15-1:0] node3342;
	wire [15-1:0] node3345;
	wire [15-1:0] node3346;
	wire [15-1:0] node3349;
	wire [15-1:0] node3352;
	wire [15-1:0] node3353;
	wire [15-1:0] node3354;
	wire [15-1:0] node3357;
	wire [15-1:0] node3360;
	wire [15-1:0] node3361;
	wire [15-1:0] node3364;
	wire [15-1:0] node3367;
	wire [15-1:0] node3368;
	wire [15-1:0] node3369;
	wire [15-1:0] node3371;
	wire [15-1:0] node3374;
	wire [15-1:0] node3375;
	wire [15-1:0] node3378;
	wire [15-1:0] node3381;
	wire [15-1:0] node3382;
	wire [15-1:0] node3384;
	wire [15-1:0] node3387;
	wire [15-1:0] node3388;
	wire [15-1:0] node3391;
	wire [15-1:0] node3394;
	wire [15-1:0] node3395;
	wire [15-1:0] node3396;
	wire [15-1:0] node3397;
	wire [15-1:0] node3398;
	wire [15-1:0] node3399;
	wire [15-1:0] node3400;
	wire [15-1:0] node3401;
	wire [15-1:0] node3404;
	wire [15-1:0] node3407;
	wire [15-1:0] node3408;
	wire [15-1:0] node3411;
	wire [15-1:0] node3414;
	wire [15-1:0] node3415;
	wire [15-1:0] node3416;
	wire [15-1:0] node3419;
	wire [15-1:0] node3422;
	wire [15-1:0] node3423;
	wire [15-1:0] node3426;
	wire [15-1:0] node3429;
	wire [15-1:0] node3430;
	wire [15-1:0] node3431;
	wire [15-1:0] node3432;
	wire [15-1:0] node3435;
	wire [15-1:0] node3438;
	wire [15-1:0] node3439;
	wire [15-1:0] node3442;
	wire [15-1:0] node3445;
	wire [15-1:0] node3446;
	wire [15-1:0] node3447;
	wire [15-1:0] node3450;
	wire [15-1:0] node3453;
	wire [15-1:0] node3454;
	wire [15-1:0] node3457;
	wire [15-1:0] node3460;
	wire [15-1:0] node3461;
	wire [15-1:0] node3462;
	wire [15-1:0] node3463;
	wire [15-1:0] node3464;
	wire [15-1:0] node3467;
	wire [15-1:0] node3470;
	wire [15-1:0] node3471;
	wire [15-1:0] node3474;
	wire [15-1:0] node3477;
	wire [15-1:0] node3478;
	wire [15-1:0] node3479;
	wire [15-1:0] node3482;
	wire [15-1:0] node3485;
	wire [15-1:0] node3486;
	wire [15-1:0] node3489;
	wire [15-1:0] node3492;
	wire [15-1:0] node3493;
	wire [15-1:0] node3494;
	wire [15-1:0] node3495;
	wire [15-1:0] node3498;
	wire [15-1:0] node3501;
	wire [15-1:0] node3502;
	wire [15-1:0] node3505;
	wire [15-1:0] node3508;
	wire [15-1:0] node3509;
	wire [15-1:0] node3510;
	wire [15-1:0] node3513;
	wire [15-1:0] node3516;
	wire [15-1:0] node3517;
	wire [15-1:0] node3520;
	wire [15-1:0] node3523;
	wire [15-1:0] node3524;
	wire [15-1:0] node3525;
	wire [15-1:0] node3526;
	wire [15-1:0] node3527;
	wire [15-1:0] node3528;
	wire [15-1:0] node3531;
	wire [15-1:0] node3534;
	wire [15-1:0] node3535;
	wire [15-1:0] node3538;
	wire [15-1:0] node3541;
	wire [15-1:0] node3542;
	wire [15-1:0] node3544;
	wire [15-1:0] node3547;
	wire [15-1:0] node3548;
	wire [15-1:0] node3551;
	wire [15-1:0] node3554;
	wire [15-1:0] node3555;
	wire [15-1:0] node3556;
	wire [15-1:0] node3557;
	wire [15-1:0] node3560;
	wire [15-1:0] node3563;
	wire [15-1:0] node3564;
	wire [15-1:0] node3567;
	wire [15-1:0] node3570;
	wire [15-1:0] node3571;
	wire [15-1:0] node3572;
	wire [15-1:0] node3576;
	wire [15-1:0] node3577;
	wire [15-1:0] node3580;
	wire [15-1:0] node3583;
	wire [15-1:0] node3584;
	wire [15-1:0] node3585;
	wire [15-1:0] node3586;
	wire [15-1:0] node3587;
	wire [15-1:0] node3591;
	wire [15-1:0] node3592;
	wire [15-1:0] node3596;
	wire [15-1:0] node3597;
	wire [15-1:0] node3598;
	wire [15-1:0] node3601;
	wire [15-1:0] node3604;
	wire [15-1:0] node3605;
	wire [15-1:0] node3609;
	wire [15-1:0] node3610;
	wire [15-1:0] node3611;
	wire [15-1:0] node3612;
	wire [15-1:0] node3615;
	wire [15-1:0] node3618;
	wire [15-1:0] node3619;
	wire [15-1:0] node3622;
	wire [15-1:0] node3625;
	wire [15-1:0] node3626;
	wire [15-1:0] node3627;
	wire [15-1:0] node3630;
	wire [15-1:0] node3633;
	wire [15-1:0] node3634;
	wire [15-1:0] node3637;
	wire [15-1:0] node3640;
	wire [15-1:0] node3641;
	wire [15-1:0] node3642;
	wire [15-1:0] node3643;
	wire [15-1:0] node3644;
	wire [15-1:0] node3645;
	wire [15-1:0] node3646;
	wire [15-1:0] node3649;
	wire [15-1:0] node3652;
	wire [15-1:0] node3653;
	wire [15-1:0] node3656;
	wire [15-1:0] node3659;
	wire [15-1:0] node3660;
	wire [15-1:0] node3661;
	wire [15-1:0] node3664;
	wire [15-1:0] node3667;
	wire [15-1:0] node3668;
	wire [15-1:0] node3671;
	wire [15-1:0] node3674;
	wire [15-1:0] node3675;
	wire [15-1:0] node3676;
	wire [15-1:0] node3677;
	wire [15-1:0] node3680;
	wire [15-1:0] node3683;
	wire [15-1:0] node3684;
	wire [15-1:0] node3687;
	wire [15-1:0] node3690;
	wire [15-1:0] node3691;
	wire [15-1:0] node3692;
	wire [15-1:0] node3695;
	wire [15-1:0] node3698;
	wire [15-1:0] node3699;
	wire [15-1:0] node3702;
	wire [15-1:0] node3705;
	wire [15-1:0] node3706;
	wire [15-1:0] node3707;
	wire [15-1:0] node3708;
	wire [15-1:0] node3709;
	wire [15-1:0] node3712;
	wire [15-1:0] node3715;
	wire [15-1:0] node3716;
	wire [15-1:0] node3719;
	wire [15-1:0] node3722;
	wire [15-1:0] node3723;
	wire [15-1:0] node3724;
	wire [15-1:0] node3727;
	wire [15-1:0] node3730;
	wire [15-1:0] node3731;
	wire [15-1:0] node3734;
	wire [15-1:0] node3737;
	wire [15-1:0] node3738;
	wire [15-1:0] node3739;
	wire [15-1:0] node3741;
	wire [15-1:0] node3744;
	wire [15-1:0] node3745;
	wire [15-1:0] node3748;
	wire [15-1:0] node3751;
	wire [15-1:0] node3752;
	wire [15-1:0] node3753;
	wire [15-1:0] node3756;
	wire [15-1:0] node3759;
	wire [15-1:0] node3760;
	wire [15-1:0] node3764;
	wire [15-1:0] node3765;
	wire [15-1:0] node3766;
	wire [15-1:0] node3767;
	wire [15-1:0] node3768;
	wire [15-1:0] node3769;
	wire [15-1:0] node3772;
	wire [15-1:0] node3775;
	wire [15-1:0] node3776;
	wire [15-1:0] node3779;
	wire [15-1:0] node3782;
	wire [15-1:0] node3783;
	wire [15-1:0] node3784;
	wire [15-1:0] node3787;
	wire [15-1:0] node3790;
	wire [15-1:0] node3791;
	wire [15-1:0] node3795;
	wire [15-1:0] node3796;
	wire [15-1:0] node3797;
	wire [15-1:0] node3798;
	wire [15-1:0] node3801;
	wire [15-1:0] node3804;
	wire [15-1:0] node3805;
	wire [15-1:0] node3808;
	wire [15-1:0] node3811;
	wire [15-1:0] node3812;
	wire [15-1:0] node3814;
	wire [15-1:0] node3817;
	wire [15-1:0] node3818;
	wire [15-1:0] node3821;
	wire [15-1:0] node3824;
	wire [15-1:0] node3825;
	wire [15-1:0] node3826;
	wire [15-1:0] node3827;
	wire [15-1:0] node3828;
	wire [15-1:0] node3831;
	wire [15-1:0] node3834;
	wire [15-1:0] node3835;
	wire [15-1:0] node3838;
	wire [15-1:0] node3841;
	wire [15-1:0] node3842;
	wire [15-1:0] node3843;
	wire [15-1:0] node3846;
	wire [15-1:0] node3849;
	wire [15-1:0] node3850;
	wire [15-1:0] node3853;
	wire [15-1:0] node3856;
	wire [15-1:0] node3857;
	wire [15-1:0] node3858;
	wire [15-1:0] node3859;
	wire [15-1:0] node3862;
	wire [15-1:0] node3865;
	wire [15-1:0] node3866;
	wire [15-1:0] node3869;
	wire [15-1:0] node3872;
	wire [15-1:0] node3873;
	wire [15-1:0] node3874;
	wire [15-1:0] node3877;
	wire [15-1:0] node3880;
	wire [15-1:0] node3881;
	wire [15-1:0] node3884;
	wire [15-1:0] node3887;
	wire [15-1:0] node3888;
	wire [15-1:0] node3889;
	wire [15-1:0] node3890;
	wire [15-1:0] node3891;
	wire [15-1:0] node3892;
	wire [15-1:0] node3893;
	wire [15-1:0] node3894;
	wire [15-1:0] node3895;
	wire [15-1:0] node3896;
	wire [15-1:0] node3897;
	wire [15-1:0] node3900;
	wire [15-1:0] node3903;
	wire [15-1:0] node3904;
	wire [15-1:0] node3908;
	wire [15-1:0] node3909;
	wire [15-1:0] node3910;
	wire [15-1:0] node3913;
	wire [15-1:0] node3916;
	wire [15-1:0] node3917;
	wire [15-1:0] node3920;
	wire [15-1:0] node3923;
	wire [15-1:0] node3924;
	wire [15-1:0] node3925;
	wire [15-1:0] node3926;
	wire [15-1:0] node3929;
	wire [15-1:0] node3932;
	wire [15-1:0] node3933;
	wire [15-1:0] node3937;
	wire [15-1:0] node3938;
	wire [15-1:0] node3939;
	wire [15-1:0] node3942;
	wire [15-1:0] node3945;
	wire [15-1:0] node3946;
	wire [15-1:0] node3949;
	wire [15-1:0] node3952;
	wire [15-1:0] node3953;
	wire [15-1:0] node3954;
	wire [15-1:0] node3955;
	wire [15-1:0] node3956;
	wire [15-1:0] node3959;
	wire [15-1:0] node3962;
	wire [15-1:0] node3964;
	wire [15-1:0] node3967;
	wire [15-1:0] node3969;
	wire [15-1:0] node3970;
	wire [15-1:0] node3974;
	wire [15-1:0] node3975;
	wire [15-1:0] node3976;
	wire [15-1:0] node3977;
	wire [15-1:0] node3980;
	wire [15-1:0] node3983;
	wire [15-1:0] node3984;
	wire [15-1:0] node3987;
	wire [15-1:0] node3990;
	wire [15-1:0] node3991;
	wire [15-1:0] node3992;
	wire [15-1:0] node3995;
	wire [15-1:0] node3998;
	wire [15-1:0] node3999;
	wire [15-1:0] node4002;
	wire [15-1:0] node4005;
	wire [15-1:0] node4006;
	wire [15-1:0] node4007;
	wire [15-1:0] node4008;
	wire [15-1:0] node4009;
	wire [15-1:0] node4010;
	wire [15-1:0] node4013;
	wire [15-1:0] node4016;
	wire [15-1:0] node4017;
	wire [15-1:0] node4020;
	wire [15-1:0] node4023;
	wire [15-1:0] node4024;
	wire [15-1:0] node4025;
	wire [15-1:0] node4028;
	wire [15-1:0] node4031;
	wire [15-1:0] node4032;
	wire [15-1:0] node4035;
	wire [15-1:0] node4038;
	wire [15-1:0] node4039;
	wire [15-1:0] node4040;
	wire [15-1:0] node4041;
	wire [15-1:0] node4044;
	wire [15-1:0] node4047;
	wire [15-1:0] node4048;
	wire [15-1:0] node4051;
	wire [15-1:0] node4054;
	wire [15-1:0] node4055;
	wire [15-1:0] node4056;
	wire [15-1:0] node4059;
	wire [15-1:0] node4062;
	wire [15-1:0] node4063;
	wire [15-1:0] node4066;
	wire [15-1:0] node4069;
	wire [15-1:0] node4070;
	wire [15-1:0] node4071;
	wire [15-1:0] node4072;
	wire [15-1:0] node4073;
	wire [15-1:0] node4076;
	wire [15-1:0] node4079;
	wire [15-1:0] node4080;
	wire [15-1:0] node4083;
	wire [15-1:0] node4086;
	wire [15-1:0] node4087;
	wire [15-1:0] node4088;
	wire [15-1:0] node4091;
	wire [15-1:0] node4094;
	wire [15-1:0] node4095;
	wire [15-1:0] node4098;
	wire [15-1:0] node4101;
	wire [15-1:0] node4102;
	wire [15-1:0] node4103;
	wire [15-1:0] node4104;
	wire [15-1:0] node4107;
	wire [15-1:0] node4110;
	wire [15-1:0] node4111;
	wire [15-1:0] node4114;
	wire [15-1:0] node4117;
	wire [15-1:0] node4118;
	wire [15-1:0] node4119;
	wire [15-1:0] node4122;
	wire [15-1:0] node4125;
	wire [15-1:0] node4126;
	wire [15-1:0] node4129;
	wire [15-1:0] node4132;
	wire [15-1:0] node4133;
	wire [15-1:0] node4134;
	wire [15-1:0] node4135;
	wire [15-1:0] node4136;
	wire [15-1:0] node4137;
	wire [15-1:0] node4138;
	wire [15-1:0] node4141;
	wire [15-1:0] node4144;
	wire [15-1:0] node4145;
	wire [15-1:0] node4148;
	wire [15-1:0] node4151;
	wire [15-1:0] node4152;
	wire [15-1:0] node4154;
	wire [15-1:0] node4157;
	wire [15-1:0] node4160;
	wire [15-1:0] node4161;
	wire [15-1:0] node4162;
	wire [15-1:0] node4164;
	wire [15-1:0] node4167;
	wire [15-1:0] node4168;
	wire [15-1:0] node4171;
	wire [15-1:0] node4174;
	wire [15-1:0] node4175;
	wire [15-1:0] node4176;
	wire [15-1:0] node4179;
	wire [15-1:0] node4182;
	wire [15-1:0] node4183;
	wire [15-1:0] node4186;
	wire [15-1:0] node4189;
	wire [15-1:0] node4190;
	wire [15-1:0] node4191;
	wire [15-1:0] node4192;
	wire [15-1:0] node4193;
	wire [15-1:0] node4196;
	wire [15-1:0] node4199;
	wire [15-1:0] node4200;
	wire [15-1:0] node4203;
	wire [15-1:0] node4206;
	wire [15-1:0] node4207;
	wire [15-1:0] node4208;
	wire [15-1:0] node4212;
	wire [15-1:0] node4213;
	wire [15-1:0] node4217;
	wire [15-1:0] node4218;
	wire [15-1:0] node4219;
	wire [15-1:0] node4220;
	wire [15-1:0] node4223;
	wire [15-1:0] node4226;
	wire [15-1:0] node4227;
	wire [15-1:0] node4230;
	wire [15-1:0] node4233;
	wire [15-1:0] node4234;
	wire [15-1:0] node4235;
	wire [15-1:0] node4238;
	wire [15-1:0] node4241;
	wire [15-1:0] node4242;
	wire [15-1:0] node4245;
	wire [15-1:0] node4248;
	wire [15-1:0] node4249;
	wire [15-1:0] node4250;
	wire [15-1:0] node4251;
	wire [15-1:0] node4252;
	wire [15-1:0] node4254;
	wire [15-1:0] node4257;
	wire [15-1:0] node4258;
	wire [15-1:0] node4262;
	wire [15-1:0] node4263;
	wire [15-1:0] node4264;
	wire [15-1:0] node4267;
	wire [15-1:0] node4270;
	wire [15-1:0] node4271;
	wire [15-1:0] node4274;
	wire [15-1:0] node4277;
	wire [15-1:0] node4278;
	wire [15-1:0] node4279;
	wire [15-1:0] node4280;
	wire [15-1:0] node4283;
	wire [15-1:0] node4286;
	wire [15-1:0] node4287;
	wire [15-1:0] node4290;
	wire [15-1:0] node4293;
	wire [15-1:0] node4295;
	wire [15-1:0] node4296;
	wire [15-1:0] node4299;
	wire [15-1:0] node4302;
	wire [15-1:0] node4303;
	wire [15-1:0] node4304;
	wire [15-1:0] node4305;
	wire [15-1:0] node4306;
	wire [15-1:0] node4309;
	wire [15-1:0] node4312;
	wire [15-1:0] node4313;
	wire [15-1:0] node4316;
	wire [15-1:0] node4319;
	wire [15-1:0] node4320;
	wire [15-1:0] node4321;
	wire [15-1:0] node4324;
	wire [15-1:0] node4327;
	wire [15-1:0] node4328;
	wire [15-1:0] node4331;
	wire [15-1:0] node4334;
	wire [15-1:0] node4335;
	wire [15-1:0] node4336;
	wire [15-1:0] node4337;
	wire [15-1:0] node4341;
	wire [15-1:0] node4342;
	wire [15-1:0] node4345;
	wire [15-1:0] node4348;
	wire [15-1:0] node4349;
	wire [15-1:0] node4350;
	wire [15-1:0] node4353;
	wire [15-1:0] node4356;
	wire [15-1:0] node4357;
	wire [15-1:0] node4360;
	wire [15-1:0] node4363;
	wire [15-1:0] node4364;
	wire [15-1:0] node4365;
	wire [15-1:0] node4366;
	wire [15-1:0] node4367;
	wire [15-1:0] node4368;
	wire [15-1:0] node4369;
	wire [15-1:0] node4370;
	wire [15-1:0] node4373;
	wire [15-1:0] node4376;
	wire [15-1:0] node4377;
	wire [15-1:0] node4380;
	wire [15-1:0] node4383;
	wire [15-1:0] node4384;
	wire [15-1:0] node4385;
	wire [15-1:0] node4389;
	wire [15-1:0] node4390;
	wire [15-1:0] node4393;
	wire [15-1:0] node4396;
	wire [15-1:0] node4397;
	wire [15-1:0] node4398;
	wire [15-1:0] node4399;
	wire [15-1:0] node4402;
	wire [15-1:0] node4405;
	wire [15-1:0] node4406;
	wire [15-1:0] node4409;
	wire [15-1:0] node4412;
	wire [15-1:0] node4413;
	wire [15-1:0] node4414;
	wire [15-1:0] node4417;
	wire [15-1:0] node4420;
	wire [15-1:0] node4421;
	wire [15-1:0] node4424;
	wire [15-1:0] node4427;
	wire [15-1:0] node4428;
	wire [15-1:0] node4429;
	wire [15-1:0] node4430;
	wire [15-1:0] node4431;
	wire [15-1:0] node4434;
	wire [15-1:0] node4437;
	wire [15-1:0] node4438;
	wire [15-1:0] node4441;
	wire [15-1:0] node4444;
	wire [15-1:0] node4445;
	wire [15-1:0] node4446;
	wire [15-1:0] node4449;
	wire [15-1:0] node4452;
	wire [15-1:0] node4453;
	wire [15-1:0] node4456;
	wire [15-1:0] node4459;
	wire [15-1:0] node4460;
	wire [15-1:0] node4461;
	wire [15-1:0] node4462;
	wire [15-1:0] node4465;
	wire [15-1:0] node4468;
	wire [15-1:0] node4469;
	wire [15-1:0] node4472;
	wire [15-1:0] node4475;
	wire [15-1:0] node4476;
	wire [15-1:0] node4477;
	wire [15-1:0] node4480;
	wire [15-1:0] node4483;
	wire [15-1:0] node4484;
	wire [15-1:0] node4487;
	wire [15-1:0] node4490;
	wire [15-1:0] node4491;
	wire [15-1:0] node4492;
	wire [15-1:0] node4493;
	wire [15-1:0] node4494;
	wire [15-1:0] node4495;
	wire [15-1:0] node4498;
	wire [15-1:0] node4501;
	wire [15-1:0] node4502;
	wire [15-1:0] node4506;
	wire [15-1:0] node4507;
	wire [15-1:0] node4508;
	wire [15-1:0] node4511;
	wire [15-1:0] node4514;
	wire [15-1:0] node4515;
	wire [15-1:0] node4518;
	wire [15-1:0] node4521;
	wire [15-1:0] node4522;
	wire [15-1:0] node4523;
	wire [15-1:0] node4524;
	wire [15-1:0] node4527;
	wire [15-1:0] node4530;
	wire [15-1:0] node4531;
	wire [15-1:0] node4535;
	wire [15-1:0] node4536;
	wire [15-1:0] node4537;
	wire [15-1:0] node4540;
	wire [15-1:0] node4543;
	wire [15-1:0] node4544;
	wire [15-1:0] node4547;
	wire [15-1:0] node4550;
	wire [15-1:0] node4551;
	wire [15-1:0] node4552;
	wire [15-1:0] node4553;
	wire [15-1:0] node4554;
	wire [15-1:0] node4557;
	wire [15-1:0] node4560;
	wire [15-1:0] node4561;
	wire [15-1:0] node4565;
	wire [15-1:0] node4566;
	wire [15-1:0] node4567;
	wire [15-1:0] node4570;
	wire [15-1:0] node4573;
	wire [15-1:0] node4574;
	wire [15-1:0] node4577;
	wire [15-1:0] node4580;
	wire [15-1:0] node4581;
	wire [15-1:0] node4582;
	wire [15-1:0] node4583;
	wire [15-1:0] node4586;
	wire [15-1:0] node4589;
	wire [15-1:0] node4590;
	wire [15-1:0] node4593;
	wire [15-1:0] node4596;
	wire [15-1:0] node4597;
	wire [15-1:0] node4598;
	wire [15-1:0] node4602;
	wire [15-1:0] node4603;
	wire [15-1:0] node4606;
	wire [15-1:0] node4609;
	wire [15-1:0] node4610;
	wire [15-1:0] node4611;
	wire [15-1:0] node4612;
	wire [15-1:0] node4613;
	wire [15-1:0] node4614;
	wire [15-1:0] node4615;
	wire [15-1:0] node4618;
	wire [15-1:0] node4621;
	wire [15-1:0] node4622;
	wire [15-1:0] node4625;
	wire [15-1:0] node4628;
	wire [15-1:0] node4629;
	wire [15-1:0] node4630;
	wire [15-1:0] node4633;
	wire [15-1:0] node4636;
	wire [15-1:0] node4637;
	wire [15-1:0] node4641;
	wire [15-1:0] node4642;
	wire [15-1:0] node4643;
	wire [15-1:0] node4644;
	wire [15-1:0] node4647;
	wire [15-1:0] node4650;
	wire [15-1:0] node4651;
	wire [15-1:0] node4654;
	wire [15-1:0] node4657;
	wire [15-1:0] node4658;
	wire [15-1:0] node4659;
	wire [15-1:0] node4662;
	wire [15-1:0] node4665;
	wire [15-1:0] node4666;
	wire [15-1:0] node4670;
	wire [15-1:0] node4671;
	wire [15-1:0] node4672;
	wire [15-1:0] node4673;
	wire [15-1:0] node4674;
	wire [15-1:0] node4678;
	wire [15-1:0] node4679;
	wire [15-1:0] node4682;
	wire [15-1:0] node4685;
	wire [15-1:0] node4686;
	wire [15-1:0] node4687;
	wire [15-1:0] node4690;
	wire [15-1:0] node4693;
	wire [15-1:0] node4694;
	wire [15-1:0] node4697;
	wire [15-1:0] node4700;
	wire [15-1:0] node4701;
	wire [15-1:0] node4702;
	wire [15-1:0] node4703;
	wire [15-1:0] node4706;
	wire [15-1:0] node4709;
	wire [15-1:0] node4710;
	wire [15-1:0] node4713;
	wire [15-1:0] node4716;
	wire [15-1:0] node4717;
	wire [15-1:0] node4718;
	wire [15-1:0] node4721;
	wire [15-1:0] node4724;
	wire [15-1:0] node4725;
	wire [15-1:0] node4728;
	wire [15-1:0] node4731;
	wire [15-1:0] node4732;
	wire [15-1:0] node4733;
	wire [15-1:0] node4734;
	wire [15-1:0] node4735;
	wire [15-1:0] node4737;
	wire [15-1:0] node4740;
	wire [15-1:0] node4741;
	wire [15-1:0] node4744;
	wire [15-1:0] node4747;
	wire [15-1:0] node4748;
	wire [15-1:0] node4749;
	wire [15-1:0] node4752;
	wire [15-1:0] node4755;
	wire [15-1:0] node4756;
	wire [15-1:0] node4759;
	wire [15-1:0] node4762;
	wire [15-1:0] node4763;
	wire [15-1:0] node4764;
	wire [15-1:0] node4766;
	wire [15-1:0] node4769;
	wire [15-1:0] node4770;
	wire [15-1:0] node4773;
	wire [15-1:0] node4776;
	wire [15-1:0] node4777;
	wire [15-1:0] node4779;
	wire [15-1:0] node4782;
	wire [15-1:0] node4784;
	wire [15-1:0] node4787;
	wire [15-1:0] node4788;
	wire [15-1:0] node4789;
	wire [15-1:0] node4790;
	wire [15-1:0] node4791;
	wire [15-1:0] node4794;
	wire [15-1:0] node4797;
	wire [15-1:0] node4798;
	wire [15-1:0] node4801;
	wire [15-1:0] node4804;
	wire [15-1:0] node4805;
	wire [15-1:0] node4806;
	wire [15-1:0] node4809;
	wire [15-1:0] node4812;
	wire [15-1:0] node4813;
	wire [15-1:0] node4817;
	wire [15-1:0] node4818;
	wire [15-1:0] node4819;
	wire [15-1:0] node4820;
	wire [15-1:0] node4823;
	wire [15-1:0] node4826;
	wire [15-1:0] node4827;
	wire [15-1:0] node4830;
	wire [15-1:0] node4833;
	wire [15-1:0] node4834;
	wire [15-1:0] node4835;
	wire [15-1:0] node4838;
	wire [15-1:0] node4841;
	wire [15-1:0] node4842;
	wire [15-1:0] node4845;
	wire [15-1:0] node4848;
	wire [15-1:0] node4849;
	wire [15-1:0] node4850;
	wire [15-1:0] node4851;
	wire [15-1:0] node4852;
	wire [15-1:0] node4853;
	wire [15-1:0] node4854;
	wire [15-1:0] node4855;
	wire [15-1:0] node4856;
	wire [15-1:0] node4859;
	wire [15-1:0] node4862;
	wire [15-1:0] node4863;
	wire [15-1:0] node4866;
	wire [15-1:0] node4869;
	wire [15-1:0] node4871;
	wire [15-1:0] node4872;
	wire [15-1:0] node4875;
	wire [15-1:0] node4878;
	wire [15-1:0] node4879;
	wire [15-1:0] node4880;
	wire [15-1:0] node4881;
	wire [15-1:0] node4884;
	wire [15-1:0] node4887;
	wire [15-1:0] node4888;
	wire [15-1:0] node4891;
	wire [15-1:0] node4894;
	wire [15-1:0] node4895;
	wire [15-1:0] node4896;
	wire [15-1:0] node4899;
	wire [15-1:0] node4902;
	wire [15-1:0] node4903;
	wire [15-1:0] node4906;
	wire [15-1:0] node4909;
	wire [15-1:0] node4910;
	wire [15-1:0] node4911;
	wire [15-1:0] node4912;
	wire [15-1:0] node4913;
	wire [15-1:0] node4916;
	wire [15-1:0] node4919;
	wire [15-1:0] node4920;
	wire [15-1:0] node4923;
	wire [15-1:0] node4926;
	wire [15-1:0] node4927;
	wire [15-1:0] node4928;
	wire [15-1:0] node4931;
	wire [15-1:0] node4934;
	wire [15-1:0] node4935;
	wire [15-1:0] node4938;
	wire [15-1:0] node4941;
	wire [15-1:0] node4942;
	wire [15-1:0] node4943;
	wire [15-1:0] node4944;
	wire [15-1:0] node4948;
	wire [15-1:0] node4949;
	wire [15-1:0] node4952;
	wire [15-1:0] node4955;
	wire [15-1:0] node4956;
	wire [15-1:0] node4958;
	wire [15-1:0] node4961;
	wire [15-1:0] node4962;
	wire [15-1:0] node4965;
	wire [15-1:0] node4968;
	wire [15-1:0] node4969;
	wire [15-1:0] node4970;
	wire [15-1:0] node4971;
	wire [15-1:0] node4972;
	wire [15-1:0] node4973;
	wire [15-1:0] node4976;
	wire [15-1:0] node4979;
	wire [15-1:0] node4980;
	wire [15-1:0] node4983;
	wire [15-1:0] node4986;
	wire [15-1:0] node4987;
	wire [15-1:0] node4988;
	wire [15-1:0] node4992;
	wire [15-1:0] node4993;
	wire [15-1:0] node4996;
	wire [15-1:0] node4999;
	wire [15-1:0] node5000;
	wire [15-1:0] node5001;
	wire [15-1:0] node5002;
	wire [15-1:0] node5005;
	wire [15-1:0] node5008;
	wire [15-1:0] node5009;
	wire [15-1:0] node5012;
	wire [15-1:0] node5015;
	wire [15-1:0] node5016;
	wire [15-1:0] node5018;
	wire [15-1:0] node5021;
	wire [15-1:0] node5023;
	wire [15-1:0] node5026;
	wire [15-1:0] node5027;
	wire [15-1:0] node5028;
	wire [15-1:0] node5029;
	wire [15-1:0] node5030;
	wire [15-1:0] node5034;
	wire [15-1:0] node5035;
	wire [15-1:0] node5038;
	wire [15-1:0] node5041;
	wire [15-1:0] node5042;
	wire [15-1:0] node5043;
	wire [15-1:0] node5046;
	wire [15-1:0] node5049;
	wire [15-1:0] node5050;
	wire [15-1:0] node5053;
	wire [15-1:0] node5056;
	wire [15-1:0] node5057;
	wire [15-1:0] node5058;
	wire [15-1:0] node5059;
	wire [15-1:0] node5063;
	wire [15-1:0] node5064;
	wire [15-1:0] node5067;
	wire [15-1:0] node5070;
	wire [15-1:0] node5071;
	wire [15-1:0] node5072;
	wire [15-1:0] node5075;
	wire [15-1:0] node5078;
	wire [15-1:0] node5079;
	wire [15-1:0] node5083;
	wire [15-1:0] node5084;
	wire [15-1:0] node5085;
	wire [15-1:0] node5086;
	wire [15-1:0] node5087;
	wire [15-1:0] node5088;
	wire [15-1:0] node5090;
	wire [15-1:0] node5093;
	wire [15-1:0] node5094;
	wire [15-1:0] node5097;
	wire [15-1:0] node5100;
	wire [15-1:0] node5101;
	wire [15-1:0] node5102;
	wire [15-1:0] node5105;
	wire [15-1:0] node5108;
	wire [15-1:0] node5109;
	wire [15-1:0] node5112;
	wire [15-1:0] node5115;
	wire [15-1:0] node5116;
	wire [15-1:0] node5117;
	wire [15-1:0] node5118;
	wire [15-1:0] node5121;
	wire [15-1:0] node5124;
	wire [15-1:0] node5125;
	wire [15-1:0] node5128;
	wire [15-1:0] node5131;
	wire [15-1:0] node5132;
	wire [15-1:0] node5133;
	wire [15-1:0] node5136;
	wire [15-1:0] node5139;
	wire [15-1:0] node5140;
	wire [15-1:0] node5144;
	wire [15-1:0] node5145;
	wire [15-1:0] node5146;
	wire [15-1:0] node5147;
	wire [15-1:0] node5148;
	wire [15-1:0] node5151;
	wire [15-1:0] node5154;
	wire [15-1:0] node5155;
	wire [15-1:0] node5158;
	wire [15-1:0] node5161;
	wire [15-1:0] node5162;
	wire [15-1:0] node5163;
	wire [15-1:0] node5166;
	wire [15-1:0] node5169;
	wire [15-1:0] node5170;
	wire [15-1:0] node5173;
	wire [15-1:0] node5176;
	wire [15-1:0] node5177;
	wire [15-1:0] node5178;
	wire [15-1:0] node5179;
	wire [15-1:0] node5182;
	wire [15-1:0] node5185;
	wire [15-1:0] node5187;
	wire [15-1:0] node5190;
	wire [15-1:0] node5191;
	wire [15-1:0] node5192;
	wire [15-1:0] node5195;
	wire [15-1:0] node5198;
	wire [15-1:0] node5199;
	wire [15-1:0] node5202;
	wire [15-1:0] node5205;
	wire [15-1:0] node5206;
	wire [15-1:0] node5207;
	wire [15-1:0] node5208;
	wire [15-1:0] node5209;
	wire [15-1:0] node5210;
	wire [15-1:0] node5214;
	wire [15-1:0] node5215;
	wire [15-1:0] node5218;
	wire [15-1:0] node5221;
	wire [15-1:0] node5222;
	wire [15-1:0] node5223;
	wire [15-1:0] node5226;
	wire [15-1:0] node5229;
	wire [15-1:0] node5230;
	wire [15-1:0] node5233;
	wire [15-1:0] node5236;
	wire [15-1:0] node5237;
	wire [15-1:0] node5238;
	wire [15-1:0] node5239;
	wire [15-1:0] node5242;
	wire [15-1:0] node5245;
	wire [15-1:0] node5246;
	wire [15-1:0] node5249;
	wire [15-1:0] node5252;
	wire [15-1:0] node5253;
	wire [15-1:0] node5254;
	wire [15-1:0] node5257;
	wire [15-1:0] node5260;
	wire [15-1:0] node5261;
	wire [15-1:0] node5264;
	wire [15-1:0] node5267;
	wire [15-1:0] node5268;
	wire [15-1:0] node5269;
	wire [15-1:0] node5270;
	wire [15-1:0] node5271;
	wire [15-1:0] node5274;
	wire [15-1:0] node5277;
	wire [15-1:0] node5278;
	wire [15-1:0] node5281;
	wire [15-1:0] node5284;
	wire [15-1:0] node5285;
	wire [15-1:0] node5286;
	wire [15-1:0] node5289;
	wire [15-1:0] node5292;
	wire [15-1:0] node5293;
	wire [15-1:0] node5297;
	wire [15-1:0] node5298;
	wire [15-1:0] node5299;
	wire [15-1:0] node5300;
	wire [15-1:0] node5304;
	wire [15-1:0] node5305;
	wire [15-1:0] node5308;
	wire [15-1:0] node5311;
	wire [15-1:0] node5312;
	wire [15-1:0] node5313;
	wire [15-1:0] node5316;
	wire [15-1:0] node5319;
	wire [15-1:0] node5320;
	wire [15-1:0] node5323;
	wire [15-1:0] node5326;
	wire [15-1:0] node5327;
	wire [15-1:0] node5328;
	wire [15-1:0] node5329;
	wire [15-1:0] node5330;
	wire [15-1:0] node5331;
	wire [15-1:0] node5332;
	wire [15-1:0] node5333;
	wire [15-1:0] node5336;
	wire [15-1:0] node5339;
	wire [15-1:0] node5340;
	wire [15-1:0] node5343;
	wire [15-1:0] node5346;
	wire [15-1:0] node5347;
	wire [15-1:0] node5348;
	wire [15-1:0] node5351;
	wire [15-1:0] node5354;
	wire [15-1:0] node5356;
	wire [15-1:0] node5359;
	wire [15-1:0] node5360;
	wire [15-1:0] node5361;
	wire [15-1:0] node5362;
	wire [15-1:0] node5365;
	wire [15-1:0] node5368;
	wire [15-1:0] node5370;
	wire [15-1:0] node5373;
	wire [15-1:0] node5374;
	wire [15-1:0] node5375;
	wire [15-1:0] node5378;
	wire [15-1:0] node5381;
	wire [15-1:0] node5382;
	wire [15-1:0] node5385;
	wire [15-1:0] node5388;
	wire [15-1:0] node5389;
	wire [15-1:0] node5390;
	wire [15-1:0] node5391;
	wire [15-1:0] node5392;
	wire [15-1:0] node5395;
	wire [15-1:0] node5398;
	wire [15-1:0] node5399;
	wire [15-1:0] node5402;
	wire [15-1:0] node5405;
	wire [15-1:0] node5406;
	wire [15-1:0] node5407;
	wire [15-1:0] node5410;
	wire [15-1:0] node5413;
	wire [15-1:0] node5416;
	wire [15-1:0] node5417;
	wire [15-1:0] node5418;
	wire [15-1:0] node5419;
	wire [15-1:0] node5422;
	wire [15-1:0] node5425;
	wire [15-1:0] node5426;
	wire [15-1:0] node5429;
	wire [15-1:0] node5432;
	wire [15-1:0] node5433;
	wire [15-1:0] node5434;
	wire [15-1:0] node5437;
	wire [15-1:0] node5440;
	wire [15-1:0] node5441;
	wire [15-1:0] node5444;
	wire [15-1:0] node5447;
	wire [15-1:0] node5448;
	wire [15-1:0] node5449;
	wire [15-1:0] node5450;
	wire [15-1:0] node5451;
	wire [15-1:0] node5452;
	wire [15-1:0] node5455;
	wire [15-1:0] node5458;
	wire [15-1:0] node5459;
	wire [15-1:0] node5463;
	wire [15-1:0] node5464;
	wire [15-1:0] node5465;
	wire [15-1:0] node5468;
	wire [15-1:0] node5471;
	wire [15-1:0] node5472;
	wire [15-1:0] node5475;
	wire [15-1:0] node5478;
	wire [15-1:0] node5479;
	wire [15-1:0] node5480;
	wire [15-1:0] node5481;
	wire [15-1:0] node5484;
	wire [15-1:0] node5487;
	wire [15-1:0] node5488;
	wire [15-1:0] node5491;
	wire [15-1:0] node5494;
	wire [15-1:0] node5495;
	wire [15-1:0] node5496;
	wire [15-1:0] node5499;
	wire [15-1:0] node5502;
	wire [15-1:0] node5503;
	wire [15-1:0] node5506;
	wire [15-1:0] node5509;
	wire [15-1:0] node5510;
	wire [15-1:0] node5511;
	wire [15-1:0] node5512;
	wire [15-1:0] node5513;
	wire [15-1:0] node5516;
	wire [15-1:0] node5519;
	wire [15-1:0] node5520;
	wire [15-1:0] node5523;
	wire [15-1:0] node5526;
	wire [15-1:0] node5527;
	wire [15-1:0] node5528;
	wire [15-1:0] node5531;
	wire [15-1:0] node5534;
	wire [15-1:0] node5535;
	wire [15-1:0] node5538;
	wire [15-1:0] node5541;
	wire [15-1:0] node5542;
	wire [15-1:0] node5543;
	wire [15-1:0] node5544;
	wire [15-1:0] node5547;
	wire [15-1:0] node5550;
	wire [15-1:0] node5551;
	wire [15-1:0] node5554;
	wire [15-1:0] node5557;
	wire [15-1:0] node5558;
	wire [15-1:0] node5559;
	wire [15-1:0] node5562;
	wire [15-1:0] node5565;
	wire [15-1:0] node5566;
	wire [15-1:0] node5569;
	wire [15-1:0] node5572;
	wire [15-1:0] node5573;
	wire [15-1:0] node5574;
	wire [15-1:0] node5575;
	wire [15-1:0] node5576;
	wire [15-1:0] node5577;
	wire [15-1:0] node5578;
	wire [15-1:0] node5582;
	wire [15-1:0] node5585;
	wire [15-1:0] node5586;
	wire [15-1:0] node5587;
	wire [15-1:0] node5590;
	wire [15-1:0] node5593;
	wire [15-1:0] node5594;
	wire [15-1:0] node5597;
	wire [15-1:0] node5600;
	wire [15-1:0] node5601;
	wire [15-1:0] node5602;
	wire [15-1:0] node5603;
	wire [15-1:0] node5606;
	wire [15-1:0] node5609;
	wire [15-1:0] node5610;
	wire [15-1:0] node5613;
	wire [15-1:0] node5616;
	wire [15-1:0] node5617;
	wire [15-1:0] node5618;
	wire [15-1:0] node5621;
	wire [15-1:0] node5624;
	wire [15-1:0] node5625;
	wire [15-1:0] node5629;
	wire [15-1:0] node5630;
	wire [15-1:0] node5631;
	wire [15-1:0] node5632;
	wire [15-1:0] node5633;
	wire [15-1:0] node5636;
	wire [15-1:0] node5639;
	wire [15-1:0] node5640;
	wire [15-1:0] node5644;
	wire [15-1:0] node5645;
	wire [15-1:0] node5646;
	wire [15-1:0] node5649;
	wire [15-1:0] node5652;
	wire [15-1:0] node5653;
	wire [15-1:0] node5657;
	wire [15-1:0] node5658;
	wire [15-1:0] node5659;
	wire [15-1:0] node5660;
	wire [15-1:0] node5663;
	wire [15-1:0] node5666;
	wire [15-1:0] node5667;
	wire [15-1:0] node5670;
	wire [15-1:0] node5673;
	wire [15-1:0] node5674;
	wire [15-1:0] node5675;
	wire [15-1:0] node5678;
	wire [15-1:0] node5681;
	wire [15-1:0] node5683;
	wire [15-1:0] node5686;
	wire [15-1:0] node5687;
	wire [15-1:0] node5688;
	wire [15-1:0] node5689;
	wire [15-1:0] node5690;
	wire [15-1:0] node5692;
	wire [15-1:0] node5695;
	wire [15-1:0] node5696;
	wire [15-1:0] node5699;
	wire [15-1:0] node5702;
	wire [15-1:0] node5703;
	wire [15-1:0] node5704;
	wire [15-1:0] node5707;
	wire [15-1:0] node5710;
	wire [15-1:0] node5711;
	wire [15-1:0] node5714;
	wire [15-1:0] node5717;
	wire [15-1:0] node5718;
	wire [15-1:0] node5719;
	wire [15-1:0] node5720;
	wire [15-1:0] node5723;
	wire [15-1:0] node5726;
	wire [15-1:0] node5727;
	wire [15-1:0] node5730;
	wire [15-1:0] node5733;
	wire [15-1:0] node5734;
	wire [15-1:0] node5735;
	wire [15-1:0] node5738;
	wire [15-1:0] node5741;
	wire [15-1:0] node5743;
	wire [15-1:0] node5746;
	wire [15-1:0] node5747;
	wire [15-1:0] node5748;
	wire [15-1:0] node5749;
	wire [15-1:0] node5750;
	wire [15-1:0] node5753;
	wire [15-1:0] node5756;
	wire [15-1:0] node5757;
	wire [15-1:0] node5760;
	wire [15-1:0] node5763;
	wire [15-1:0] node5764;
	wire [15-1:0] node5765;
	wire [15-1:0] node5768;
	wire [15-1:0] node5771;
	wire [15-1:0] node5772;
	wire [15-1:0] node5775;
	wire [15-1:0] node5778;
	wire [15-1:0] node5779;
	wire [15-1:0] node5780;
	wire [15-1:0] node5781;
	wire [15-1:0] node5784;
	wire [15-1:0] node5787;
	wire [15-1:0] node5788;
	wire [15-1:0] node5791;
	wire [15-1:0] node5794;
	wire [15-1:0] node5795;
	wire [15-1:0] node5796;
	wire [15-1:0] node5799;
	wire [15-1:0] node5802;
	wire [15-1:0] node5803;
	wire [15-1:0] node5806;
	wire [15-1:0] node5809;
	wire [15-1:0] node5810;
	wire [15-1:0] node5811;
	wire [15-1:0] node5812;
	wire [15-1:0] node5813;
	wire [15-1:0] node5814;
	wire [15-1:0] node5815;
	wire [15-1:0] node5816;
	wire [15-1:0] node5817;
	wire [15-1:0] node5818;
	wire [15-1:0] node5821;
	wire [15-1:0] node5824;
	wire [15-1:0] node5825;
	wire [15-1:0] node5828;
	wire [15-1:0] node5831;
	wire [15-1:0] node5832;
	wire [15-1:0] node5833;
	wire [15-1:0] node5837;
	wire [15-1:0] node5838;
	wire [15-1:0] node5841;
	wire [15-1:0] node5844;
	wire [15-1:0] node5845;
	wire [15-1:0] node5846;
	wire [15-1:0] node5848;
	wire [15-1:0] node5851;
	wire [15-1:0] node5852;
	wire [15-1:0] node5855;
	wire [15-1:0] node5858;
	wire [15-1:0] node5859;
	wire [15-1:0] node5860;
	wire [15-1:0] node5863;
	wire [15-1:0] node5866;
	wire [15-1:0] node5867;
	wire [15-1:0] node5870;
	wire [15-1:0] node5873;
	wire [15-1:0] node5874;
	wire [15-1:0] node5875;
	wire [15-1:0] node5876;
	wire [15-1:0] node5877;
	wire [15-1:0] node5880;
	wire [15-1:0] node5883;
	wire [15-1:0] node5884;
	wire [15-1:0] node5887;
	wire [15-1:0] node5890;
	wire [15-1:0] node5891;
	wire [15-1:0] node5892;
	wire [15-1:0] node5895;
	wire [15-1:0] node5898;
	wire [15-1:0] node5899;
	wire [15-1:0] node5902;
	wire [15-1:0] node5905;
	wire [15-1:0] node5906;
	wire [15-1:0] node5907;
	wire [15-1:0] node5908;
	wire [15-1:0] node5911;
	wire [15-1:0] node5914;
	wire [15-1:0] node5915;
	wire [15-1:0] node5919;
	wire [15-1:0] node5920;
	wire [15-1:0] node5921;
	wire [15-1:0] node5924;
	wire [15-1:0] node5927;
	wire [15-1:0] node5928;
	wire [15-1:0] node5931;
	wire [15-1:0] node5934;
	wire [15-1:0] node5935;
	wire [15-1:0] node5936;
	wire [15-1:0] node5937;
	wire [15-1:0] node5938;
	wire [15-1:0] node5939;
	wire [15-1:0] node5942;
	wire [15-1:0] node5945;
	wire [15-1:0] node5946;
	wire [15-1:0] node5950;
	wire [15-1:0] node5951;
	wire [15-1:0] node5952;
	wire [15-1:0] node5955;
	wire [15-1:0] node5958;
	wire [15-1:0] node5959;
	wire [15-1:0] node5963;
	wire [15-1:0] node5964;
	wire [15-1:0] node5965;
	wire [15-1:0] node5966;
	wire [15-1:0] node5969;
	wire [15-1:0] node5972;
	wire [15-1:0] node5973;
	wire [15-1:0] node5977;
	wire [15-1:0] node5978;
	wire [15-1:0] node5979;
	wire [15-1:0] node5982;
	wire [15-1:0] node5985;
	wire [15-1:0] node5986;
	wire [15-1:0] node5989;
	wire [15-1:0] node5992;
	wire [15-1:0] node5993;
	wire [15-1:0] node5994;
	wire [15-1:0] node5995;
	wire [15-1:0] node5996;
	wire [15-1:0] node5999;
	wire [15-1:0] node6002;
	wire [15-1:0] node6003;
	wire [15-1:0] node6006;
	wire [15-1:0] node6009;
	wire [15-1:0] node6010;
	wire [15-1:0] node6011;
	wire [15-1:0] node6014;
	wire [15-1:0] node6017;
	wire [15-1:0] node6018;
	wire [15-1:0] node6021;
	wire [15-1:0] node6024;
	wire [15-1:0] node6025;
	wire [15-1:0] node6026;
	wire [15-1:0] node6027;
	wire [15-1:0] node6030;
	wire [15-1:0] node6033;
	wire [15-1:0] node6034;
	wire [15-1:0] node6037;
	wire [15-1:0] node6040;
	wire [15-1:0] node6041;
	wire [15-1:0] node6042;
	wire [15-1:0] node6045;
	wire [15-1:0] node6048;
	wire [15-1:0] node6049;
	wire [15-1:0] node6052;
	wire [15-1:0] node6055;
	wire [15-1:0] node6056;
	wire [15-1:0] node6057;
	wire [15-1:0] node6058;
	wire [15-1:0] node6059;
	wire [15-1:0] node6060;
	wire [15-1:0] node6061;
	wire [15-1:0] node6064;
	wire [15-1:0] node6067;
	wire [15-1:0] node6068;
	wire [15-1:0] node6072;
	wire [15-1:0] node6073;
	wire [15-1:0] node6074;
	wire [15-1:0] node6077;
	wire [15-1:0] node6080;
	wire [15-1:0] node6081;
	wire [15-1:0] node6084;
	wire [15-1:0] node6087;
	wire [15-1:0] node6088;
	wire [15-1:0] node6089;
	wire [15-1:0] node6090;
	wire [15-1:0] node6093;
	wire [15-1:0] node6096;
	wire [15-1:0] node6097;
	wire [15-1:0] node6100;
	wire [15-1:0] node6103;
	wire [15-1:0] node6104;
	wire [15-1:0] node6107;
	wire [15-1:0] node6109;
	wire [15-1:0] node6112;
	wire [15-1:0] node6113;
	wire [15-1:0] node6114;
	wire [15-1:0] node6115;
	wire [15-1:0] node6116;
	wire [15-1:0] node6120;
	wire [15-1:0] node6121;
	wire [15-1:0] node6124;
	wire [15-1:0] node6127;
	wire [15-1:0] node6128;
	wire [15-1:0] node6129;
	wire [15-1:0] node6132;
	wire [15-1:0] node6135;
	wire [15-1:0] node6136;
	wire [15-1:0] node6140;
	wire [15-1:0] node6141;
	wire [15-1:0] node6142;
	wire [15-1:0] node6143;
	wire [15-1:0] node6146;
	wire [15-1:0] node6149;
	wire [15-1:0] node6150;
	wire [15-1:0] node6153;
	wire [15-1:0] node6156;
	wire [15-1:0] node6157;
	wire [15-1:0] node6158;
	wire [15-1:0] node6161;
	wire [15-1:0] node6164;
	wire [15-1:0] node6165;
	wire [15-1:0] node6168;
	wire [15-1:0] node6171;
	wire [15-1:0] node6172;
	wire [15-1:0] node6173;
	wire [15-1:0] node6174;
	wire [15-1:0] node6175;
	wire [15-1:0] node6176;
	wire [15-1:0] node6179;
	wire [15-1:0] node6182;
	wire [15-1:0] node6185;
	wire [15-1:0] node6186;
	wire [15-1:0] node6188;
	wire [15-1:0] node6191;
	wire [15-1:0] node6192;
	wire [15-1:0] node6195;
	wire [15-1:0] node6198;
	wire [15-1:0] node6199;
	wire [15-1:0] node6200;
	wire [15-1:0] node6201;
	wire [15-1:0] node6204;
	wire [15-1:0] node6207;
	wire [15-1:0] node6208;
	wire [15-1:0] node6211;
	wire [15-1:0] node6214;
	wire [15-1:0] node6215;
	wire [15-1:0] node6216;
	wire [15-1:0] node6219;
	wire [15-1:0] node6222;
	wire [15-1:0] node6223;
	wire [15-1:0] node6226;
	wire [15-1:0] node6229;
	wire [15-1:0] node6230;
	wire [15-1:0] node6231;
	wire [15-1:0] node6232;
	wire [15-1:0] node6233;
	wire [15-1:0] node6236;
	wire [15-1:0] node6239;
	wire [15-1:0] node6240;
	wire [15-1:0] node6243;
	wire [15-1:0] node6246;
	wire [15-1:0] node6247;
	wire [15-1:0] node6248;
	wire [15-1:0] node6251;
	wire [15-1:0] node6254;
	wire [15-1:0] node6255;
	wire [15-1:0] node6258;
	wire [15-1:0] node6261;
	wire [15-1:0] node6262;
	wire [15-1:0] node6263;
	wire [15-1:0] node6266;
	wire [15-1:0] node6267;
	wire [15-1:0] node6270;
	wire [15-1:0] node6273;
	wire [15-1:0] node6274;
	wire [15-1:0] node6275;
	wire [15-1:0] node6278;
	wire [15-1:0] node6281;
	wire [15-1:0] node6283;
	wire [15-1:0] node6286;
	wire [15-1:0] node6287;
	wire [15-1:0] node6288;
	wire [15-1:0] node6289;
	wire [15-1:0] node6290;
	wire [15-1:0] node6291;
	wire [15-1:0] node6292;
	wire [15-1:0] node6293;
	wire [15-1:0] node6296;
	wire [15-1:0] node6299;
	wire [15-1:0] node6300;
	wire [15-1:0] node6303;
	wire [15-1:0] node6306;
	wire [15-1:0] node6307;
	wire [15-1:0] node6308;
	wire [15-1:0] node6311;
	wire [15-1:0] node6314;
	wire [15-1:0] node6315;
	wire [15-1:0] node6318;
	wire [15-1:0] node6321;
	wire [15-1:0] node6322;
	wire [15-1:0] node6323;
	wire [15-1:0] node6324;
	wire [15-1:0] node6327;
	wire [15-1:0] node6330;
	wire [15-1:0] node6331;
	wire [15-1:0] node6334;
	wire [15-1:0] node6337;
	wire [15-1:0] node6338;
	wire [15-1:0] node6339;
	wire [15-1:0] node6342;
	wire [15-1:0] node6345;
	wire [15-1:0] node6346;
	wire [15-1:0] node6350;
	wire [15-1:0] node6351;
	wire [15-1:0] node6352;
	wire [15-1:0] node6353;
	wire [15-1:0] node6354;
	wire [15-1:0] node6358;
	wire [15-1:0] node6359;
	wire [15-1:0] node6362;
	wire [15-1:0] node6365;
	wire [15-1:0] node6366;
	wire [15-1:0] node6367;
	wire [15-1:0] node6370;
	wire [15-1:0] node6373;
	wire [15-1:0] node6374;
	wire [15-1:0] node6377;
	wire [15-1:0] node6380;
	wire [15-1:0] node6381;
	wire [15-1:0] node6382;
	wire [15-1:0] node6383;
	wire [15-1:0] node6386;
	wire [15-1:0] node6389;
	wire [15-1:0] node6390;
	wire [15-1:0] node6393;
	wire [15-1:0] node6396;
	wire [15-1:0] node6397;
	wire [15-1:0] node6399;
	wire [15-1:0] node6402;
	wire [15-1:0] node6403;
	wire [15-1:0] node6406;
	wire [15-1:0] node6409;
	wire [15-1:0] node6410;
	wire [15-1:0] node6411;
	wire [15-1:0] node6412;
	wire [15-1:0] node6413;
	wire [15-1:0] node6414;
	wire [15-1:0] node6417;
	wire [15-1:0] node6420;
	wire [15-1:0] node6421;
	wire [15-1:0] node6424;
	wire [15-1:0] node6427;
	wire [15-1:0] node6428;
	wire [15-1:0] node6429;
	wire [15-1:0] node6432;
	wire [15-1:0] node6435;
	wire [15-1:0] node6436;
	wire [15-1:0] node6439;
	wire [15-1:0] node6442;
	wire [15-1:0] node6443;
	wire [15-1:0] node6444;
	wire [15-1:0] node6446;
	wire [15-1:0] node6449;
	wire [15-1:0] node6450;
	wire [15-1:0] node6453;
	wire [15-1:0] node6456;
	wire [15-1:0] node6457;
	wire [15-1:0] node6458;
	wire [15-1:0] node6461;
	wire [15-1:0] node6464;
	wire [15-1:0] node6465;
	wire [15-1:0] node6468;
	wire [15-1:0] node6471;
	wire [15-1:0] node6472;
	wire [15-1:0] node6473;
	wire [15-1:0] node6474;
	wire [15-1:0] node6475;
	wire [15-1:0] node6478;
	wire [15-1:0] node6481;
	wire [15-1:0] node6482;
	wire [15-1:0] node6485;
	wire [15-1:0] node6488;
	wire [15-1:0] node6489;
	wire [15-1:0] node6490;
	wire [15-1:0] node6493;
	wire [15-1:0] node6496;
	wire [15-1:0] node6497;
	wire [15-1:0] node6500;
	wire [15-1:0] node6503;
	wire [15-1:0] node6504;
	wire [15-1:0] node6505;
	wire [15-1:0] node6506;
	wire [15-1:0] node6509;
	wire [15-1:0] node6512;
	wire [15-1:0] node6513;
	wire [15-1:0] node6516;
	wire [15-1:0] node6519;
	wire [15-1:0] node6520;
	wire [15-1:0] node6521;
	wire [15-1:0] node6524;
	wire [15-1:0] node6527;
	wire [15-1:0] node6528;
	wire [15-1:0] node6531;
	wire [15-1:0] node6534;
	wire [15-1:0] node6535;
	wire [15-1:0] node6536;
	wire [15-1:0] node6537;
	wire [15-1:0] node6538;
	wire [15-1:0] node6539;
	wire [15-1:0] node6541;
	wire [15-1:0] node6544;
	wire [15-1:0] node6545;
	wire [15-1:0] node6548;
	wire [15-1:0] node6551;
	wire [15-1:0] node6552;
	wire [15-1:0] node6553;
	wire [15-1:0] node6556;
	wire [15-1:0] node6559;
	wire [15-1:0] node6560;
	wire [15-1:0] node6563;
	wire [15-1:0] node6566;
	wire [15-1:0] node6567;
	wire [15-1:0] node6568;
	wire [15-1:0] node6570;
	wire [15-1:0] node6573;
	wire [15-1:0] node6575;
	wire [15-1:0] node6578;
	wire [15-1:0] node6579;
	wire [15-1:0] node6581;
	wire [15-1:0] node6584;
	wire [15-1:0] node6585;
	wire [15-1:0] node6588;
	wire [15-1:0] node6591;
	wire [15-1:0] node6592;
	wire [15-1:0] node6593;
	wire [15-1:0] node6594;
	wire [15-1:0] node6595;
	wire [15-1:0] node6598;
	wire [15-1:0] node6601;
	wire [15-1:0] node6603;
	wire [15-1:0] node6606;
	wire [15-1:0] node6607;
	wire [15-1:0] node6608;
	wire [15-1:0] node6611;
	wire [15-1:0] node6614;
	wire [15-1:0] node6615;
	wire [15-1:0] node6618;
	wire [15-1:0] node6621;
	wire [15-1:0] node6622;
	wire [15-1:0] node6623;
	wire [15-1:0] node6625;
	wire [15-1:0] node6628;
	wire [15-1:0] node6629;
	wire [15-1:0] node6632;
	wire [15-1:0] node6635;
	wire [15-1:0] node6636;
	wire [15-1:0] node6638;
	wire [15-1:0] node6641;
	wire [15-1:0] node6642;
	wire [15-1:0] node6645;
	wire [15-1:0] node6648;
	wire [15-1:0] node6649;
	wire [15-1:0] node6650;
	wire [15-1:0] node6651;
	wire [15-1:0] node6652;
	wire [15-1:0] node6654;
	wire [15-1:0] node6657;
	wire [15-1:0] node6658;
	wire [15-1:0] node6662;
	wire [15-1:0] node6663;
	wire [15-1:0] node6664;
	wire [15-1:0] node6667;
	wire [15-1:0] node6670;
	wire [15-1:0] node6671;
	wire [15-1:0] node6674;
	wire [15-1:0] node6677;
	wire [15-1:0] node6678;
	wire [15-1:0] node6679;
	wire [15-1:0] node6680;
	wire [15-1:0] node6683;
	wire [15-1:0] node6686;
	wire [15-1:0] node6687;
	wire [15-1:0] node6690;
	wire [15-1:0] node6693;
	wire [15-1:0] node6694;
	wire [15-1:0] node6696;
	wire [15-1:0] node6699;
	wire [15-1:0] node6700;
	wire [15-1:0] node6704;
	wire [15-1:0] node6705;
	wire [15-1:0] node6706;
	wire [15-1:0] node6707;
	wire [15-1:0] node6708;
	wire [15-1:0] node6711;
	wire [15-1:0] node6714;
	wire [15-1:0] node6715;
	wire [15-1:0] node6718;
	wire [15-1:0] node6721;
	wire [15-1:0] node6722;
	wire [15-1:0] node6723;
	wire [15-1:0] node6726;
	wire [15-1:0] node6729;
	wire [15-1:0] node6730;
	wire [15-1:0] node6733;
	wire [15-1:0] node6736;
	wire [15-1:0] node6737;
	wire [15-1:0] node6738;
	wire [15-1:0] node6739;
	wire [15-1:0] node6742;
	wire [15-1:0] node6745;
	wire [15-1:0] node6746;
	wire [15-1:0] node6749;
	wire [15-1:0] node6752;
	wire [15-1:0] node6753;
	wire [15-1:0] node6754;
	wire [15-1:0] node6757;
	wire [15-1:0] node6760;
	wire [15-1:0] node6761;
	wire [15-1:0] node6764;
	wire [15-1:0] node6767;
	wire [15-1:0] node6768;
	wire [15-1:0] node6769;
	wire [15-1:0] node6770;
	wire [15-1:0] node6771;
	wire [15-1:0] node6772;
	wire [15-1:0] node6773;
	wire [15-1:0] node6774;
	wire [15-1:0] node6775;
	wire [15-1:0] node6778;
	wire [15-1:0] node6781;
	wire [15-1:0] node6782;
	wire [15-1:0] node6785;
	wire [15-1:0] node6788;
	wire [15-1:0] node6789;
	wire [15-1:0] node6790;
	wire [15-1:0] node6793;
	wire [15-1:0] node6796;
	wire [15-1:0] node6797;
	wire [15-1:0] node6800;
	wire [15-1:0] node6803;
	wire [15-1:0] node6804;
	wire [15-1:0] node6805;
	wire [15-1:0] node6806;
	wire [15-1:0] node6809;
	wire [15-1:0] node6812;
	wire [15-1:0] node6813;
	wire [15-1:0] node6817;
	wire [15-1:0] node6818;
	wire [15-1:0] node6819;
	wire [15-1:0] node6822;
	wire [15-1:0] node6825;
	wire [15-1:0] node6826;
	wire [15-1:0] node6829;
	wire [15-1:0] node6832;
	wire [15-1:0] node6833;
	wire [15-1:0] node6834;
	wire [15-1:0] node6835;
	wire [15-1:0] node6836;
	wire [15-1:0] node6839;
	wire [15-1:0] node6842;
	wire [15-1:0] node6843;
	wire [15-1:0] node6846;
	wire [15-1:0] node6849;
	wire [15-1:0] node6850;
	wire [15-1:0] node6851;
	wire [15-1:0] node6854;
	wire [15-1:0] node6857;
	wire [15-1:0] node6858;
	wire [15-1:0] node6861;
	wire [15-1:0] node6864;
	wire [15-1:0] node6865;
	wire [15-1:0] node6866;
	wire [15-1:0] node6868;
	wire [15-1:0] node6871;
	wire [15-1:0] node6872;
	wire [15-1:0] node6875;
	wire [15-1:0] node6878;
	wire [15-1:0] node6879;
	wire [15-1:0] node6880;
	wire [15-1:0] node6883;
	wire [15-1:0] node6886;
	wire [15-1:0] node6887;
	wire [15-1:0] node6890;
	wire [15-1:0] node6893;
	wire [15-1:0] node6894;
	wire [15-1:0] node6895;
	wire [15-1:0] node6896;
	wire [15-1:0] node6897;
	wire [15-1:0] node6898;
	wire [15-1:0] node6902;
	wire [15-1:0] node6903;
	wire [15-1:0] node6906;
	wire [15-1:0] node6909;
	wire [15-1:0] node6910;
	wire [15-1:0] node6911;
	wire [15-1:0] node6914;
	wire [15-1:0] node6917;
	wire [15-1:0] node6918;
	wire [15-1:0] node6921;
	wire [15-1:0] node6924;
	wire [15-1:0] node6925;
	wire [15-1:0] node6926;
	wire [15-1:0] node6927;
	wire [15-1:0] node6930;
	wire [15-1:0] node6933;
	wire [15-1:0] node6934;
	wire [15-1:0] node6937;
	wire [15-1:0] node6940;
	wire [15-1:0] node6941;
	wire [15-1:0] node6942;
	wire [15-1:0] node6945;
	wire [15-1:0] node6948;
	wire [15-1:0] node6949;
	wire [15-1:0] node6952;
	wire [15-1:0] node6955;
	wire [15-1:0] node6956;
	wire [15-1:0] node6957;
	wire [15-1:0] node6958;
	wire [15-1:0] node6959;
	wire [15-1:0] node6962;
	wire [15-1:0] node6965;
	wire [15-1:0] node6966;
	wire [15-1:0] node6969;
	wire [15-1:0] node6972;
	wire [15-1:0] node6973;
	wire [15-1:0] node6974;
	wire [15-1:0] node6977;
	wire [15-1:0] node6980;
	wire [15-1:0] node6981;
	wire [15-1:0] node6984;
	wire [15-1:0] node6987;
	wire [15-1:0] node6988;
	wire [15-1:0] node6989;
	wire [15-1:0] node6990;
	wire [15-1:0] node6993;
	wire [15-1:0] node6996;
	wire [15-1:0] node6997;
	wire [15-1:0] node7000;
	wire [15-1:0] node7003;
	wire [15-1:0] node7004;
	wire [15-1:0] node7005;
	wire [15-1:0] node7008;
	wire [15-1:0] node7011;
	wire [15-1:0] node7012;
	wire [15-1:0] node7015;
	wire [15-1:0] node7018;
	wire [15-1:0] node7019;
	wire [15-1:0] node7020;
	wire [15-1:0] node7021;
	wire [15-1:0] node7022;
	wire [15-1:0] node7023;
	wire [15-1:0] node7024;
	wire [15-1:0] node7027;
	wire [15-1:0] node7030;
	wire [15-1:0] node7031;
	wire [15-1:0] node7034;
	wire [15-1:0] node7037;
	wire [15-1:0] node7038;
	wire [15-1:0] node7039;
	wire [15-1:0] node7042;
	wire [15-1:0] node7045;
	wire [15-1:0] node7046;
	wire [15-1:0] node7049;
	wire [15-1:0] node7052;
	wire [15-1:0] node7053;
	wire [15-1:0] node7054;
	wire [15-1:0] node7055;
	wire [15-1:0] node7058;
	wire [15-1:0] node7061;
	wire [15-1:0] node7062;
	wire [15-1:0] node7065;
	wire [15-1:0] node7068;
	wire [15-1:0] node7069;
	wire [15-1:0] node7070;
	wire [15-1:0] node7073;
	wire [15-1:0] node7076;
	wire [15-1:0] node7077;
	wire [15-1:0] node7080;
	wire [15-1:0] node7083;
	wire [15-1:0] node7084;
	wire [15-1:0] node7085;
	wire [15-1:0] node7086;
	wire [15-1:0] node7087;
	wire [15-1:0] node7091;
	wire [15-1:0] node7092;
	wire [15-1:0] node7095;
	wire [15-1:0] node7098;
	wire [15-1:0] node7099;
	wire [15-1:0] node7100;
	wire [15-1:0] node7103;
	wire [15-1:0] node7106;
	wire [15-1:0] node7108;
	wire [15-1:0] node7111;
	wire [15-1:0] node7112;
	wire [15-1:0] node7113;
	wire [15-1:0] node7115;
	wire [15-1:0] node7118;
	wire [15-1:0] node7119;
	wire [15-1:0] node7122;
	wire [15-1:0] node7125;
	wire [15-1:0] node7126;
	wire [15-1:0] node7127;
	wire [15-1:0] node7130;
	wire [15-1:0] node7133;
	wire [15-1:0] node7134;
	wire [15-1:0] node7137;
	wire [15-1:0] node7140;
	wire [15-1:0] node7141;
	wire [15-1:0] node7142;
	wire [15-1:0] node7143;
	wire [15-1:0] node7144;
	wire [15-1:0] node7145;
	wire [15-1:0] node7149;
	wire [15-1:0] node7150;
	wire [15-1:0] node7153;
	wire [15-1:0] node7156;
	wire [15-1:0] node7157;
	wire [15-1:0] node7158;
	wire [15-1:0] node7161;
	wire [15-1:0] node7164;
	wire [15-1:0] node7165;
	wire [15-1:0] node7168;
	wire [15-1:0] node7171;
	wire [15-1:0] node7172;
	wire [15-1:0] node7173;
	wire [15-1:0] node7174;
	wire [15-1:0] node7177;
	wire [15-1:0] node7180;
	wire [15-1:0] node7181;
	wire [15-1:0] node7184;
	wire [15-1:0] node7187;
	wire [15-1:0] node7188;
	wire [15-1:0] node7189;
	wire [15-1:0] node7192;
	wire [15-1:0] node7195;
	wire [15-1:0] node7196;
	wire [15-1:0] node7199;
	wire [15-1:0] node7202;
	wire [15-1:0] node7203;
	wire [15-1:0] node7204;
	wire [15-1:0] node7205;
	wire [15-1:0] node7206;
	wire [15-1:0] node7209;
	wire [15-1:0] node7212;
	wire [15-1:0] node7213;
	wire [15-1:0] node7216;
	wire [15-1:0] node7219;
	wire [15-1:0] node7220;
	wire [15-1:0] node7221;
	wire [15-1:0] node7224;
	wire [15-1:0] node7227;
	wire [15-1:0] node7229;
	wire [15-1:0] node7232;
	wire [15-1:0] node7233;
	wire [15-1:0] node7234;
	wire [15-1:0] node7235;
	wire [15-1:0] node7238;
	wire [15-1:0] node7241;
	wire [15-1:0] node7242;
	wire [15-1:0] node7245;
	wire [15-1:0] node7248;
	wire [15-1:0] node7249;
	wire [15-1:0] node7251;
	wire [15-1:0] node7254;
	wire [15-1:0] node7255;
	wire [15-1:0] node7258;
	wire [15-1:0] node7261;
	wire [15-1:0] node7262;
	wire [15-1:0] node7263;
	wire [15-1:0] node7264;
	wire [15-1:0] node7265;
	wire [15-1:0] node7266;
	wire [15-1:0] node7267;
	wire [15-1:0] node7268;
	wire [15-1:0] node7271;
	wire [15-1:0] node7274;
	wire [15-1:0] node7275;
	wire [15-1:0] node7279;
	wire [15-1:0] node7280;
	wire [15-1:0] node7281;
	wire [15-1:0] node7284;
	wire [15-1:0] node7287;
	wire [15-1:0] node7288;
	wire [15-1:0] node7291;
	wire [15-1:0] node7294;
	wire [15-1:0] node7295;
	wire [15-1:0] node7296;
	wire [15-1:0] node7298;
	wire [15-1:0] node7301;
	wire [15-1:0] node7302;
	wire [15-1:0] node7305;
	wire [15-1:0] node7308;
	wire [15-1:0] node7309;
	wire [15-1:0] node7310;
	wire [15-1:0] node7313;
	wire [15-1:0] node7316;
	wire [15-1:0] node7318;
	wire [15-1:0] node7321;
	wire [15-1:0] node7322;
	wire [15-1:0] node7323;
	wire [15-1:0] node7324;
	wire [15-1:0] node7325;
	wire [15-1:0] node7328;
	wire [15-1:0] node7331;
	wire [15-1:0] node7332;
	wire [15-1:0] node7335;
	wire [15-1:0] node7338;
	wire [15-1:0] node7339;
	wire [15-1:0] node7340;
	wire [15-1:0] node7343;
	wire [15-1:0] node7346;
	wire [15-1:0] node7347;
	wire [15-1:0] node7350;
	wire [15-1:0] node7353;
	wire [15-1:0] node7354;
	wire [15-1:0] node7355;
	wire [15-1:0] node7356;
	wire [15-1:0] node7359;
	wire [15-1:0] node7362;
	wire [15-1:0] node7363;
	wire [15-1:0] node7367;
	wire [15-1:0] node7368;
	wire [15-1:0] node7369;
	wire [15-1:0] node7372;
	wire [15-1:0] node7375;
	wire [15-1:0] node7376;
	wire [15-1:0] node7379;
	wire [15-1:0] node7382;
	wire [15-1:0] node7383;
	wire [15-1:0] node7384;
	wire [15-1:0] node7385;
	wire [15-1:0] node7386;
	wire [15-1:0] node7387;
	wire [15-1:0] node7390;
	wire [15-1:0] node7393;
	wire [15-1:0] node7394;
	wire [15-1:0] node7397;
	wire [15-1:0] node7400;
	wire [15-1:0] node7401;
	wire [15-1:0] node7402;
	wire [15-1:0] node7405;
	wire [15-1:0] node7408;
	wire [15-1:0] node7409;
	wire [15-1:0] node7412;
	wire [15-1:0] node7415;
	wire [15-1:0] node7416;
	wire [15-1:0] node7417;
	wire [15-1:0] node7419;
	wire [15-1:0] node7422;
	wire [15-1:0] node7423;
	wire [15-1:0] node7426;
	wire [15-1:0] node7429;
	wire [15-1:0] node7430;
	wire [15-1:0] node7431;
	wire [15-1:0] node7434;
	wire [15-1:0] node7437;
	wire [15-1:0] node7438;
	wire [15-1:0] node7441;
	wire [15-1:0] node7444;
	wire [15-1:0] node7445;
	wire [15-1:0] node7446;
	wire [15-1:0] node7447;
	wire [15-1:0] node7448;
	wire [15-1:0] node7451;
	wire [15-1:0] node7454;
	wire [15-1:0] node7455;
	wire [15-1:0] node7458;
	wire [15-1:0] node7461;
	wire [15-1:0] node7462;
	wire [15-1:0] node7463;
	wire [15-1:0] node7466;
	wire [15-1:0] node7469;
	wire [15-1:0] node7470;
	wire [15-1:0] node7473;
	wire [15-1:0] node7476;
	wire [15-1:0] node7477;
	wire [15-1:0] node7478;
	wire [15-1:0] node7479;
	wire [15-1:0] node7483;
	wire [15-1:0] node7484;
	wire [15-1:0] node7487;
	wire [15-1:0] node7490;
	wire [15-1:0] node7491;
	wire [15-1:0] node7492;
	wire [15-1:0] node7495;
	wire [15-1:0] node7498;
	wire [15-1:0] node7499;
	wire [15-1:0] node7502;
	wire [15-1:0] node7505;
	wire [15-1:0] node7506;
	wire [15-1:0] node7507;
	wire [15-1:0] node7508;
	wire [15-1:0] node7509;
	wire [15-1:0] node7510;
	wire [15-1:0] node7511;
	wire [15-1:0] node7514;
	wire [15-1:0] node7517;
	wire [15-1:0] node7518;
	wire [15-1:0] node7521;
	wire [15-1:0] node7524;
	wire [15-1:0] node7525;
	wire [15-1:0] node7526;
	wire [15-1:0] node7530;
	wire [15-1:0] node7531;
	wire [15-1:0] node7534;
	wire [15-1:0] node7537;
	wire [15-1:0] node7538;
	wire [15-1:0] node7539;
	wire [15-1:0] node7540;
	wire [15-1:0] node7543;
	wire [15-1:0] node7546;
	wire [15-1:0] node7548;
	wire [15-1:0] node7551;
	wire [15-1:0] node7552;
	wire [15-1:0] node7553;
	wire [15-1:0] node7556;
	wire [15-1:0] node7559;
	wire [15-1:0] node7560;
	wire [15-1:0] node7563;
	wire [15-1:0] node7566;
	wire [15-1:0] node7567;
	wire [15-1:0] node7568;
	wire [15-1:0] node7569;
	wire [15-1:0] node7570;
	wire [15-1:0] node7573;
	wire [15-1:0] node7576;
	wire [15-1:0] node7577;
	wire [15-1:0] node7580;
	wire [15-1:0] node7583;
	wire [15-1:0] node7584;
	wire [15-1:0] node7585;
	wire [15-1:0] node7588;
	wire [15-1:0] node7591;
	wire [15-1:0] node7592;
	wire [15-1:0] node7595;
	wire [15-1:0] node7598;
	wire [15-1:0] node7599;
	wire [15-1:0] node7600;
	wire [15-1:0] node7601;
	wire [15-1:0] node7604;
	wire [15-1:0] node7607;
	wire [15-1:0] node7608;
	wire [15-1:0] node7611;
	wire [15-1:0] node7614;
	wire [15-1:0] node7615;
	wire [15-1:0] node7616;
	wire [15-1:0] node7619;
	wire [15-1:0] node7622;
	wire [15-1:0] node7623;
	wire [15-1:0] node7626;
	wire [15-1:0] node7629;
	wire [15-1:0] node7630;
	wire [15-1:0] node7631;
	wire [15-1:0] node7632;
	wire [15-1:0] node7633;
	wire [15-1:0] node7634;
	wire [15-1:0] node7637;
	wire [15-1:0] node7640;
	wire [15-1:0] node7641;
	wire [15-1:0] node7645;
	wire [15-1:0] node7646;
	wire [15-1:0] node7647;
	wire [15-1:0] node7650;
	wire [15-1:0] node7653;
	wire [15-1:0] node7654;
	wire [15-1:0] node7657;
	wire [15-1:0] node7660;
	wire [15-1:0] node7661;
	wire [15-1:0] node7662;
	wire [15-1:0] node7663;
	wire [15-1:0] node7666;
	wire [15-1:0] node7669;
	wire [15-1:0] node7670;
	wire [15-1:0] node7673;
	wire [15-1:0] node7676;
	wire [15-1:0] node7677;
	wire [15-1:0] node7678;
	wire [15-1:0] node7681;
	wire [15-1:0] node7684;
	wire [15-1:0] node7685;
	wire [15-1:0] node7688;
	wire [15-1:0] node7691;
	wire [15-1:0] node7692;
	wire [15-1:0] node7693;
	wire [15-1:0] node7694;
	wire [15-1:0] node7695;
	wire [15-1:0] node7698;
	wire [15-1:0] node7701;
	wire [15-1:0] node7702;
	wire [15-1:0] node7705;
	wire [15-1:0] node7708;
	wire [15-1:0] node7709;
	wire [15-1:0] node7710;
	wire [15-1:0] node7713;
	wire [15-1:0] node7716;
	wire [15-1:0] node7717;
	wire [15-1:0] node7720;
	wire [15-1:0] node7723;
	wire [15-1:0] node7724;
	wire [15-1:0] node7725;
	wire [15-1:0] node7726;
	wire [15-1:0] node7729;
	wire [15-1:0] node7732;
	wire [15-1:0] node7733;
	wire [15-1:0] node7736;
	wire [15-1:0] node7739;
	wire [15-1:0] node7740;
	wire [15-1:0] node7741;
	wire [15-1:0] node7744;
	wire [15-1:0] node7747;
	wire [15-1:0] node7748;
	wire [15-1:0] node7751;
	wire [15-1:0] node7754;
	wire [15-1:0] node7755;
	wire [15-1:0] node7756;
	wire [15-1:0] node7757;
	wire [15-1:0] node7758;
	wire [15-1:0] node7759;
	wire [15-1:0] node7760;
	wire [15-1:0] node7761;
	wire [15-1:0] node7762;
	wire [15-1:0] node7763;
	wire [15-1:0] node7764;
	wire [15-1:0] node7765;
	wire [15-1:0] node7768;
	wire [15-1:0] node7771;
	wire [15-1:0] node7772;
	wire [15-1:0] node7775;
	wire [15-1:0] node7778;
	wire [15-1:0] node7779;
	wire [15-1:0] node7781;
	wire [15-1:0] node7784;
	wire [15-1:0] node7785;
	wire [15-1:0] node7789;
	wire [15-1:0] node7790;
	wire [15-1:0] node7791;
	wire [15-1:0] node7792;
	wire [15-1:0] node7795;
	wire [15-1:0] node7798;
	wire [15-1:0] node7799;
	wire [15-1:0] node7802;
	wire [15-1:0] node7805;
	wire [15-1:0] node7806;
	wire [15-1:0] node7807;
	wire [15-1:0] node7811;
	wire [15-1:0] node7812;
	wire [15-1:0] node7815;
	wire [15-1:0] node7818;
	wire [15-1:0] node7819;
	wire [15-1:0] node7820;
	wire [15-1:0] node7821;
	wire [15-1:0] node7822;
	wire [15-1:0] node7825;
	wire [15-1:0] node7828;
	wire [15-1:0] node7829;
	wire [15-1:0] node7832;
	wire [15-1:0] node7835;
	wire [15-1:0] node7836;
	wire [15-1:0] node7837;
	wire [15-1:0] node7840;
	wire [15-1:0] node7843;
	wire [15-1:0] node7845;
	wire [15-1:0] node7848;
	wire [15-1:0] node7849;
	wire [15-1:0] node7850;
	wire [15-1:0] node7851;
	wire [15-1:0] node7854;
	wire [15-1:0] node7857;
	wire [15-1:0] node7858;
	wire [15-1:0] node7861;
	wire [15-1:0] node7864;
	wire [15-1:0] node7865;
	wire [15-1:0] node7866;
	wire [15-1:0] node7869;
	wire [15-1:0] node7872;
	wire [15-1:0] node7873;
	wire [15-1:0] node7876;
	wire [15-1:0] node7879;
	wire [15-1:0] node7880;
	wire [15-1:0] node7881;
	wire [15-1:0] node7882;
	wire [15-1:0] node7883;
	wire [15-1:0] node7884;
	wire [15-1:0] node7887;
	wire [15-1:0] node7890;
	wire [15-1:0] node7891;
	wire [15-1:0] node7894;
	wire [15-1:0] node7897;
	wire [15-1:0] node7898;
	wire [15-1:0] node7899;
	wire [15-1:0] node7902;
	wire [15-1:0] node7905;
	wire [15-1:0] node7906;
	wire [15-1:0] node7909;
	wire [15-1:0] node7912;
	wire [15-1:0] node7913;
	wire [15-1:0] node7914;
	wire [15-1:0] node7915;
	wire [15-1:0] node7918;
	wire [15-1:0] node7921;
	wire [15-1:0] node7922;
	wire [15-1:0] node7925;
	wire [15-1:0] node7928;
	wire [15-1:0] node7929;
	wire [15-1:0] node7930;
	wire [15-1:0] node7933;
	wire [15-1:0] node7936;
	wire [15-1:0] node7937;
	wire [15-1:0] node7940;
	wire [15-1:0] node7943;
	wire [15-1:0] node7944;
	wire [15-1:0] node7945;
	wire [15-1:0] node7946;
	wire [15-1:0] node7947;
	wire [15-1:0] node7950;
	wire [15-1:0] node7953;
	wire [15-1:0] node7954;
	wire [15-1:0] node7957;
	wire [15-1:0] node7960;
	wire [15-1:0] node7961;
	wire [15-1:0] node7962;
	wire [15-1:0] node7965;
	wire [15-1:0] node7968;
	wire [15-1:0] node7969;
	wire [15-1:0] node7972;
	wire [15-1:0] node7975;
	wire [15-1:0] node7976;
	wire [15-1:0] node7977;
	wire [15-1:0] node7978;
	wire [15-1:0] node7981;
	wire [15-1:0] node7984;
	wire [15-1:0] node7985;
	wire [15-1:0] node7988;
	wire [15-1:0] node7991;
	wire [15-1:0] node7992;
	wire [15-1:0] node7993;
	wire [15-1:0] node7996;
	wire [15-1:0] node7999;
	wire [15-1:0] node8000;
	wire [15-1:0] node8003;
	wire [15-1:0] node8006;
	wire [15-1:0] node8007;
	wire [15-1:0] node8008;
	wire [15-1:0] node8009;
	wire [15-1:0] node8010;
	wire [15-1:0] node8011;
	wire [15-1:0] node8012;
	wire [15-1:0] node8015;
	wire [15-1:0] node8018;
	wire [15-1:0] node8019;
	wire [15-1:0] node8022;
	wire [15-1:0] node8025;
	wire [15-1:0] node8026;
	wire [15-1:0] node8027;
	wire [15-1:0] node8030;
	wire [15-1:0] node8033;
	wire [15-1:0] node8034;
	wire [15-1:0] node8038;
	wire [15-1:0] node8039;
	wire [15-1:0] node8040;
	wire [15-1:0] node8041;
	wire [15-1:0] node8044;
	wire [15-1:0] node8047;
	wire [15-1:0] node8048;
	wire [15-1:0] node8051;
	wire [15-1:0] node8054;
	wire [15-1:0] node8055;
	wire [15-1:0] node8056;
	wire [15-1:0] node8059;
	wire [15-1:0] node8062;
	wire [15-1:0] node8063;
	wire [15-1:0] node8066;
	wire [15-1:0] node8069;
	wire [15-1:0] node8070;
	wire [15-1:0] node8071;
	wire [15-1:0] node8072;
	wire [15-1:0] node8073;
	wire [15-1:0] node8076;
	wire [15-1:0] node8079;
	wire [15-1:0] node8080;
	wire [15-1:0] node8083;
	wire [15-1:0] node8086;
	wire [15-1:0] node8087;
	wire [15-1:0] node8089;
	wire [15-1:0] node8092;
	wire [15-1:0] node8093;
	wire [15-1:0] node8096;
	wire [15-1:0] node8099;
	wire [15-1:0] node8100;
	wire [15-1:0] node8101;
	wire [15-1:0] node8102;
	wire [15-1:0] node8105;
	wire [15-1:0] node8108;
	wire [15-1:0] node8109;
	wire [15-1:0] node8112;
	wire [15-1:0] node8115;
	wire [15-1:0] node8116;
	wire [15-1:0] node8117;
	wire [15-1:0] node8120;
	wire [15-1:0] node8123;
	wire [15-1:0] node8124;
	wire [15-1:0] node8127;
	wire [15-1:0] node8130;
	wire [15-1:0] node8131;
	wire [15-1:0] node8132;
	wire [15-1:0] node8133;
	wire [15-1:0] node8134;
	wire [15-1:0] node8135;
	wire [15-1:0] node8138;
	wire [15-1:0] node8141;
	wire [15-1:0] node8142;
	wire [15-1:0] node8145;
	wire [15-1:0] node8148;
	wire [15-1:0] node8149;
	wire [15-1:0] node8150;
	wire [15-1:0] node8153;
	wire [15-1:0] node8156;
	wire [15-1:0] node8157;
	wire [15-1:0] node8160;
	wire [15-1:0] node8163;
	wire [15-1:0] node8164;
	wire [15-1:0] node8165;
	wire [15-1:0] node8166;
	wire [15-1:0] node8169;
	wire [15-1:0] node8172;
	wire [15-1:0] node8173;
	wire [15-1:0] node8176;
	wire [15-1:0] node8179;
	wire [15-1:0] node8180;
	wire [15-1:0] node8181;
	wire [15-1:0] node8184;
	wire [15-1:0] node8187;
	wire [15-1:0] node8188;
	wire [15-1:0] node8191;
	wire [15-1:0] node8194;
	wire [15-1:0] node8195;
	wire [15-1:0] node8196;
	wire [15-1:0] node8197;
	wire [15-1:0] node8198;
	wire [15-1:0] node8201;
	wire [15-1:0] node8204;
	wire [15-1:0] node8205;
	wire [15-1:0] node8208;
	wire [15-1:0] node8211;
	wire [15-1:0] node8212;
	wire [15-1:0] node8213;
	wire [15-1:0] node8216;
	wire [15-1:0] node8219;
	wire [15-1:0] node8220;
	wire [15-1:0] node8224;
	wire [15-1:0] node8225;
	wire [15-1:0] node8226;
	wire [15-1:0] node8227;
	wire [15-1:0] node8230;
	wire [15-1:0] node8233;
	wire [15-1:0] node8234;
	wire [15-1:0] node8237;
	wire [15-1:0] node8240;
	wire [15-1:0] node8241;
	wire [15-1:0] node8243;
	wire [15-1:0] node8246;
	wire [15-1:0] node8247;
	wire [15-1:0] node8250;
	wire [15-1:0] node8253;
	wire [15-1:0] node8254;
	wire [15-1:0] node8255;
	wire [15-1:0] node8256;
	wire [15-1:0] node8257;
	wire [15-1:0] node8258;
	wire [15-1:0] node8259;
	wire [15-1:0] node8260;
	wire [15-1:0] node8263;
	wire [15-1:0] node8266;
	wire [15-1:0] node8267;
	wire [15-1:0] node8270;
	wire [15-1:0] node8273;
	wire [15-1:0] node8274;
	wire [15-1:0] node8275;
	wire [15-1:0] node8278;
	wire [15-1:0] node8281;
	wire [15-1:0] node8282;
	wire [15-1:0] node8285;
	wire [15-1:0] node8288;
	wire [15-1:0] node8289;
	wire [15-1:0] node8290;
	wire [15-1:0] node8291;
	wire [15-1:0] node8294;
	wire [15-1:0] node8297;
	wire [15-1:0] node8298;
	wire [15-1:0] node8301;
	wire [15-1:0] node8304;
	wire [15-1:0] node8305;
	wire [15-1:0] node8306;
	wire [15-1:0] node8309;
	wire [15-1:0] node8312;
	wire [15-1:0] node8313;
	wire [15-1:0] node8316;
	wire [15-1:0] node8319;
	wire [15-1:0] node8320;
	wire [15-1:0] node8321;
	wire [15-1:0] node8322;
	wire [15-1:0] node8323;
	wire [15-1:0] node8326;
	wire [15-1:0] node8329;
	wire [15-1:0] node8330;
	wire [15-1:0] node8333;
	wire [15-1:0] node8336;
	wire [15-1:0] node8337;
	wire [15-1:0] node8338;
	wire [15-1:0] node8341;
	wire [15-1:0] node8344;
	wire [15-1:0] node8345;
	wire [15-1:0] node8348;
	wire [15-1:0] node8351;
	wire [15-1:0] node8352;
	wire [15-1:0] node8353;
	wire [15-1:0] node8354;
	wire [15-1:0] node8357;
	wire [15-1:0] node8360;
	wire [15-1:0] node8361;
	wire [15-1:0] node8364;
	wire [15-1:0] node8367;
	wire [15-1:0] node8368;
	wire [15-1:0] node8369;
	wire [15-1:0] node8372;
	wire [15-1:0] node8375;
	wire [15-1:0] node8376;
	wire [15-1:0] node8379;
	wire [15-1:0] node8382;
	wire [15-1:0] node8383;
	wire [15-1:0] node8384;
	wire [15-1:0] node8385;
	wire [15-1:0] node8386;
	wire [15-1:0] node8387;
	wire [15-1:0] node8390;
	wire [15-1:0] node8393;
	wire [15-1:0] node8394;
	wire [15-1:0] node8397;
	wire [15-1:0] node8400;
	wire [15-1:0] node8401;
	wire [15-1:0] node8402;
	wire [15-1:0] node8405;
	wire [15-1:0] node8408;
	wire [15-1:0] node8410;
	wire [15-1:0] node8413;
	wire [15-1:0] node8414;
	wire [15-1:0] node8415;
	wire [15-1:0] node8416;
	wire [15-1:0] node8419;
	wire [15-1:0] node8422;
	wire [15-1:0] node8423;
	wire [15-1:0] node8426;
	wire [15-1:0] node8429;
	wire [15-1:0] node8430;
	wire [15-1:0] node8431;
	wire [15-1:0] node8434;
	wire [15-1:0] node8437;
	wire [15-1:0] node8438;
	wire [15-1:0] node8441;
	wire [15-1:0] node8444;
	wire [15-1:0] node8445;
	wire [15-1:0] node8446;
	wire [15-1:0] node8447;
	wire [15-1:0] node8448;
	wire [15-1:0] node8451;
	wire [15-1:0] node8454;
	wire [15-1:0] node8455;
	wire [15-1:0] node8458;
	wire [15-1:0] node8461;
	wire [15-1:0] node8462;
	wire [15-1:0] node8463;
	wire [15-1:0] node8467;
	wire [15-1:0] node8469;
	wire [15-1:0] node8472;
	wire [15-1:0] node8473;
	wire [15-1:0] node8474;
	wire [15-1:0] node8475;
	wire [15-1:0] node8478;
	wire [15-1:0] node8481;
	wire [15-1:0] node8482;
	wire [15-1:0] node8485;
	wire [15-1:0] node8488;
	wire [15-1:0] node8489;
	wire [15-1:0] node8490;
	wire [15-1:0] node8493;
	wire [15-1:0] node8496;
	wire [15-1:0] node8497;
	wire [15-1:0] node8500;
	wire [15-1:0] node8503;
	wire [15-1:0] node8504;
	wire [15-1:0] node8505;
	wire [15-1:0] node8506;
	wire [15-1:0] node8507;
	wire [15-1:0] node8508;
	wire [15-1:0] node8509;
	wire [15-1:0] node8512;
	wire [15-1:0] node8515;
	wire [15-1:0] node8516;
	wire [15-1:0] node8520;
	wire [15-1:0] node8521;
	wire [15-1:0] node8522;
	wire [15-1:0] node8526;
	wire [15-1:0] node8527;
	wire [15-1:0] node8530;
	wire [15-1:0] node8533;
	wire [15-1:0] node8534;
	wire [15-1:0] node8535;
	wire [15-1:0] node8536;
	wire [15-1:0] node8539;
	wire [15-1:0] node8542;
	wire [15-1:0] node8543;
	wire [15-1:0] node8546;
	wire [15-1:0] node8549;
	wire [15-1:0] node8550;
	wire [15-1:0] node8551;
	wire [15-1:0] node8554;
	wire [15-1:0] node8557;
	wire [15-1:0] node8558;
	wire [15-1:0] node8561;
	wire [15-1:0] node8564;
	wire [15-1:0] node8565;
	wire [15-1:0] node8566;
	wire [15-1:0] node8567;
	wire [15-1:0] node8568;
	wire [15-1:0] node8571;
	wire [15-1:0] node8574;
	wire [15-1:0] node8575;
	wire [15-1:0] node8578;
	wire [15-1:0] node8581;
	wire [15-1:0] node8582;
	wire [15-1:0] node8583;
	wire [15-1:0] node8586;
	wire [15-1:0] node8589;
	wire [15-1:0] node8590;
	wire [15-1:0] node8593;
	wire [15-1:0] node8596;
	wire [15-1:0] node8597;
	wire [15-1:0] node8598;
	wire [15-1:0] node8599;
	wire [15-1:0] node8602;
	wire [15-1:0] node8605;
	wire [15-1:0] node8606;
	wire [15-1:0] node8609;
	wire [15-1:0] node8612;
	wire [15-1:0] node8613;
	wire [15-1:0] node8614;
	wire [15-1:0] node8617;
	wire [15-1:0] node8620;
	wire [15-1:0] node8621;
	wire [15-1:0] node8624;
	wire [15-1:0] node8627;
	wire [15-1:0] node8628;
	wire [15-1:0] node8629;
	wire [15-1:0] node8630;
	wire [15-1:0] node8631;
	wire [15-1:0] node8632;
	wire [15-1:0] node8635;
	wire [15-1:0] node8638;
	wire [15-1:0] node8639;
	wire [15-1:0] node8642;
	wire [15-1:0] node8645;
	wire [15-1:0] node8646;
	wire [15-1:0] node8647;
	wire [15-1:0] node8650;
	wire [15-1:0] node8653;
	wire [15-1:0] node8654;
	wire [15-1:0] node8657;
	wire [15-1:0] node8660;
	wire [15-1:0] node8661;
	wire [15-1:0] node8662;
	wire [15-1:0] node8664;
	wire [15-1:0] node8667;
	wire [15-1:0] node8668;
	wire [15-1:0] node8671;
	wire [15-1:0] node8674;
	wire [15-1:0] node8675;
	wire [15-1:0] node8676;
	wire [15-1:0] node8679;
	wire [15-1:0] node8682;
	wire [15-1:0] node8683;
	wire [15-1:0] node8686;
	wire [15-1:0] node8689;
	wire [15-1:0] node8690;
	wire [15-1:0] node8691;
	wire [15-1:0] node8692;
	wire [15-1:0] node8693;
	wire [15-1:0] node8696;
	wire [15-1:0] node8699;
	wire [15-1:0] node8700;
	wire [15-1:0] node8703;
	wire [15-1:0] node8706;
	wire [15-1:0] node8707;
	wire [15-1:0] node8708;
	wire [15-1:0] node8711;
	wire [15-1:0] node8714;
	wire [15-1:0] node8715;
	wire [15-1:0] node8718;
	wire [15-1:0] node8721;
	wire [15-1:0] node8722;
	wire [15-1:0] node8723;
	wire [15-1:0] node8724;
	wire [15-1:0] node8727;
	wire [15-1:0] node8730;
	wire [15-1:0] node8731;
	wire [15-1:0] node8734;
	wire [15-1:0] node8737;
	wire [15-1:0] node8738;
	wire [15-1:0] node8739;
	wire [15-1:0] node8742;
	wire [15-1:0] node8745;
	wire [15-1:0] node8746;
	wire [15-1:0] node8749;
	wire [15-1:0] node8752;
	wire [15-1:0] node8753;
	wire [15-1:0] node8754;
	wire [15-1:0] node8755;
	wire [15-1:0] node8756;
	wire [15-1:0] node8757;
	wire [15-1:0] node8758;
	wire [15-1:0] node8759;
	wire [15-1:0] node8760;
	wire [15-1:0] node8763;
	wire [15-1:0] node8766;
	wire [15-1:0] node8767;
	wire [15-1:0] node8771;
	wire [15-1:0] node8772;
	wire [15-1:0] node8773;
	wire [15-1:0] node8776;
	wire [15-1:0] node8779;
	wire [15-1:0] node8780;
	wire [15-1:0] node8783;
	wire [15-1:0] node8786;
	wire [15-1:0] node8787;
	wire [15-1:0] node8788;
	wire [15-1:0] node8789;
	wire [15-1:0] node8792;
	wire [15-1:0] node8795;
	wire [15-1:0] node8796;
	wire [15-1:0] node8800;
	wire [15-1:0] node8801;
	wire [15-1:0] node8802;
	wire [15-1:0] node8805;
	wire [15-1:0] node8808;
	wire [15-1:0] node8809;
	wire [15-1:0] node8812;
	wire [15-1:0] node8815;
	wire [15-1:0] node8816;
	wire [15-1:0] node8817;
	wire [15-1:0] node8818;
	wire [15-1:0] node8819;
	wire [15-1:0] node8822;
	wire [15-1:0] node8825;
	wire [15-1:0] node8826;
	wire [15-1:0] node8829;
	wire [15-1:0] node8832;
	wire [15-1:0] node8834;
	wire [15-1:0] node8835;
	wire [15-1:0] node8838;
	wire [15-1:0] node8841;
	wire [15-1:0] node8842;
	wire [15-1:0] node8843;
	wire [15-1:0] node8844;
	wire [15-1:0] node8847;
	wire [15-1:0] node8850;
	wire [15-1:0] node8851;
	wire [15-1:0] node8854;
	wire [15-1:0] node8857;
	wire [15-1:0] node8858;
	wire [15-1:0] node8859;
	wire [15-1:0] node8862;
	wire [15-1:0] node8865;
	wire [15-1:0] node8866;
	wire [15-1:0] node8869;
	wire [15-1:0] node8872;
	wire [15-1:0] node8873;
	wire [15-1:0] node8874;
	wire [15-1:0] node8875;
	wire [15-1:0] node8876;
	wire [15-1:0] node8877;
	wire [15-1:0] node8880;
	wire [15-1:0] node8883;
	wire [15-1:0] node8884;
	wire [15-1:0] node8887;
	wire [15-1:0] node8890;
	wire [15-1:0] node8891;
	wire [15-1:0] node8892;
	wire [15-1:0] node8895;
	wire [15-1:0] node8898;
	wire [15-1:0] node8899;
	wire [15-1:0] node8902;
	wire [15-1:0] node8905;
	wire [15-1:0] node8906;
	wire [15-1:0] node8907;
	wire [15-1:0] node8908;
	wire [15-1:0] node8911;
	wire [15-1:0] node8914;
	wire [15-1:0] node8915;
	wire [15-1:0] node8918;
	wire [15-1:0] node8921;
	wire [15-1:0] node8922;
	wire [15-1:0] node8923;
	wire [15-1:0] node8926;
	wire [15-1:0] node8929;
	wire [15-1:0] node8930;
	wire [15-1:0] node8933;
	wire [15-1:0] node8936;
	wire [15-1:0] node8937;
	wire [15-1:0] node8938;
	wire [15-1:0] node8939;
	wire [15-1:0] node8940;
	wire [15-1:0] node8943;
	wire [15-1:0] node8946;
	wire [15-1:0] node8947;
	wire [15-1:0] node8950;
	wire [15-1:0] node8953;
	wire [15-1:0] node8954;
	wire [15-1:0] node8955;
	wire [15-1:0] node8958;
	wire [15-1:0] node8961;
	wire [15-1:0] node8962;
	wire [15-1:0] node8965;
	wire [15-1:0] node8968;
	wire [15-1:0] node8969;
	wire [15-1:0] node8970;
	wire [15-1:0] node8971;
	wire [15-1:0] node8974;
	wire [15-1:0] node8977;
	wire [15-1:0] node8978;
	wire [15-1:0] node8981;
	wire [15-1:0] node8984;
	wire [15-1:0] node8985;
	wire [15-1:0] node8986;
	wire [15-1:0] node8989;
	wire [15-1:0] node8992;
	wire [15-1:0] node8993;
	wire [15-1:0] node8996;
	wire [15-1:0] node8999;
	wire [15-1:0] node9000;
	wire [15-1:0] node9001;
	wire [15-1:0] node9002;
	wire [15-1:0] node9003;
	wire [15-1:0] node9004;
	wire [15-1:0] node9005;
	wire [15-1:0] node9008;
	wire [15-1:0] node9011;
	wire [15-1:0] node9012;
	wire [15-1:0] node9015;
	wire [15-1:0] node9018;
	wire [15-1:0] node9019;
	wire [15-1:0] node9020;
	wire [15-1:0] node9023;
	wire [15-1:0] node9026;
	wire [15-1:0] node9027;
	wire [15-1:0] node9030;
	wire [15-1:0] node9033;
	wire [15-1:0] node9034;
	wire [15-1:0] node9035;
	wire [15-1:0] node9036;
	wire [15-1:0] node9039;
	wire [15-1:0] node9042;
	wire [15-1:0] node9043;
	wire [15-1:0] node9046;
	wire [15-1:0] node9049;
	wire [15-1:0] node9050;
	wire [15-1:0] node9051;
	wire [15-1:0] node9054;
	wire [15-1:0] node9057;
	wire [15-1:0] node9058;
	wire [15-1:0] node9061;
	wire [15-1:0] node9064;
	wire [15-1:0] node9065;
	wire [15-1:0] node9066;
	wire [15-1:0] node9067;
	wire [15-1:0] node9068;
	wire [15-1:0] node9072;
	wire [15-1:0] node9073;
	wire [15-1:0] node9076;
	wire [15-1:0] node9079;
	wire [15-1:0] node9080;
	wire [15-1:0] node9081;
	wire [15-1:0] node9084;
	wire [15-1:0] node9087;
	wire [15-1:0] node9088;
	wire [15-1:0] node9091;
	wire [15-1:0] node9094;
	wire [15-1:0] node9095;
	wire [15-1:0] node9096;
	wire [15-1:0] node9097;
	wire [15-1:0] node9100;
	wire [15-1:0] node9103;
	wire [15-1:0] node9105;
	wire [15-1:0] node9108;
	wire [15-1:0] node9109;
	wire [15-1:0] node9110;
	wire [15-1:0] node9113;
	wire [15-1:0] node9116;
	wire [15-1:0] node9117;
	wire [15-1:0] node9120;
	wire [15-1:0] node9123;
	wire [15-1:0] node9124;
	wire [15-1:0] node9125;
	wire [15-1:0] node9126;
	wire [15-1:0] node9128;
	wire [15-1:0] node9130;
	wire [15-1:0] node9133;
	wire [15-1:0] node9134;
	wire [15-1:0] node9135;
	wire [15-1:0] node9138;
	wire [15-1:0] node9141;
	wire [15-1:0] node9142;
	wire [15-1:0] node9145;
	wire [15-1:0] node9148;
	wire [15-1:0] node9149;
	wire [15-1:0] node9150;
	wire [15-1:0] node9151;
	wire [15-1:0] node9154;
	wire [15-1:0] node9157;
	wire [15-1:0] node9158;
	wire [15-1:0] node9161;
	wire [15-1:0] node9164;
	wire [15-1:0] node9165;
	wire [15-1:0] node9166;
	wire [15-1:0] node9169;
	wire [15-1:0] node9172;
	wire [15-1:0] node9174;
	wire [15-1:0] node9177;
	wire [15-1:0] node9178;
	wire [15-1:0] node9179;
	wire [15-1:0] node9180;
	wire [15-1:0] node9181;
	wire [15-1:0] node9184;
	wire [15-1:0] node9187;
	wire [15-1:0] node9188;
	wire [15-1:0] node9191;
	wire [15-1:0] node9194;
	wire [15-1:0] node9195;
	wire [15-1:0] node9196;
	wire [15-1:0] node9199;
	wire [15-1:0] node9202;
	wire [15-1:0] node9203;
	wire [15-1:0] node9206;
	wire [15-1:0] node9209;
	wire [15-1:0] node9210;
	wire [15-1:0] node9211;
	wire [15-1:0] node9212;
	wire [15-1:0] node9215;
	wire [15-1:0] node9218;
	wire [15-1:0] node9219;
	wire [15-1:0] node9222;
	wire [15-1:0] node9225;
	wire [15-1:0] node9226;
	wire [15-1:0] node9228;
	wire [15-1:0] node9231;
	wire [15-1:0] node9232;
	wire [15-1:0] node9235;
	wire [15-1:0] node9238;
	wire [15-1:0] node9239;
	wire [15-1:0] node9240;
	wire [15-1:0] node9241;
	wire [15-1:0] node9242;
	wire [15-1:0] node9243;
	wire [15-1:0] node9244;
	wire [15-1:0] node9245;
	wire [15-1:0] node9249;
	wire [15-1:0] node9250;
	wire [15-1:0] node9253;
	wire [15-1:0] node9256;
	wire [15-1:0] node9257;
	wire [15-1:0] node9258;
	wire [15-1:0] node9261;
	wire [15-1:0] node9264;
	wire [15-1:0] node9265;
	wire [15-1:0] node9269;
	wire [15-1:0] node9270;
	wire [15-1:0] node9271;
	wire [15-1:0] node9272;
	wire [15-1:0] node9275;
	wire [15-1:0] node9278;
	wire [15-1:0] node9279;
	wire [15-1:0] node9282;
	wire [15-1:0] node9285;
	wire [15-1:0] node9286;
	wire [15-1:0] node9287;
	wire [15-1:0] node9290;
	wire [15-1:0] node9293;
	wire [15-1:0] node9294;
	wire [15-1:0] node9297;
	wire [15-1:0] node9300;
	wire [15-1:0] node9301;
	wire [15-1:0] node9302;
	wire [15-1:0] node9303;
	wire [15-1:0] node9304;
	wire [15-1:0] node9308;
	wire [15-1:0] node9309;
	wire [15-1:0] node9312;
	wire [15-1:0] node9315;
	wire [15-1:0] node9316;
	wire [15-1:0] node9317;
	wire [15-1:0] node9320;
	wire [15-1:0] node9323;
	wire [15-1:0] node9325;
	wire [15-1:0] node9328;
	wire [15-1:0] node9329;
	wire [15-1:0] node9330;
	wire [15-1:0] node9331;
	wire [15-1:0] node9334;
	wire [15-1:0] node9337;
	wire [15-1:0] node9338;
	wire [15-1:0] node9341;
	wire [15-1:0] node9344;
	wire [15-1:0] node9345;
	wire [15-1:0] node9346;
	wire [15-1:0] node9349;
	wire [15-1:0] node9352;
	wire [15-1:0] node9353;
	wire [15-1:0] node9356;
	wire [15-1:0] node9359;
	wire [15-1:0] node9360;
	wire [15-1:0] node9361;
	wire [15-1:0] node9362;
	wire [15-1:0] node9363;
	wire [15-1:0] node9364;
	wire [15-1:0] node9367;
	wire [15-1:0] node9370;
	wire [15-1:0] node9372;
	wire [15-1:0] node9375;
	wire [15-1:0] node9376;
	wire [15-1:0] node9377;
	wire [15-1:0] node9380;
	wire [15-1:0] node9383;
	wire [15-1:0] node9384;
	wire [15-1:0] node9387;
	wire [15-1:0] node9390;
	wire [15-1:0] node9391;
	wire [15-1:0] node9392;
	wire [15-1:0] node9393;
	wire [15-1:0] node9396;
	wire [15-1:0] node9399;
	wire [15-1:0] node9400;
	wire [15-1:0] node9403;
	wire [15-1:0] node9406;
	wire [15-1:0] node9407;
	wire [15-1:0] node9408;
	wire [15-1:0] node9411;
	wire [15-1:0] node9414;
	wire [15-1:0] node9416;
	wire [15-1:0] node9419;
	wire [15-1:0] node9420;
	wire [15-1:0] node9421;
	wire [15-1:0] node9422;
	wire [15-1:0] node9423;
	wire [15-1:0] node9427;
	wire [15-1:0] node9429;
	wire [15-1:0] node9432;
	wire [15-1:0] node9433;
	wire [15-1:0] node9434;
	wire [15-1:0] node9437;
	wire [15-1:0] node9440;
	wire [15-1:0] node9441;
	wire [15-1:0] node9444;
	wire [15-1:0] node9447;
	wire [15-1:0] node9448;
	wire [15-1:0] node9449;
	wire [15-1:0] node9451;
	wire [15-1:0] node9454;
	wire [15-1:0] node9455;
	wire [15-1:0] node9458;
	wire [15-1:0] node9461;
	wire [15-1:0] node9462;
	wire [15-1:0] node9463;
	wire [15-1:0] node9466;
	wire [15-1:0] node9469;
	wire [15-1:0] node9470;
	wire [15-1:0] node9473;
	wire [15-1:0] node9476;
	wire [15-1:0] node9477;
	wire [15-1:0] node9478;
	wire [15-1:0] node9479;
	wire [15-1:0] node9480;
	wire [15-1:0] node9481;
	wire [15-1:0] node9482;
	wire [15-1:0] node9485;
	wire [15-1:0] node9488;
	wire [15-1:0] node9489;
	wire [15-1:0] node9492;
	wire [15-1:0] node9495;
	wire [15-1:0] node9496;
	wire [15-1:0] node9497;
	wire [15-1:0] node9500;
	wire [15-1:0] node9503;
	wire [15-1:0] node9504;
	wire [15-1:0] node9507;
	wire [15-1:0] node9510;
	wire [15-1:0] node9511;
	wire [15-1:0] node9512;
	wire [15-1:0] node9513;
	wire [15-1:0] node9516;
	wire [15-1:0] node9519;
	wire [15-1:0] node9520;
	wire [15-1:0] node9523;
	wire [15-1:0] node9526;
	wire [15-1:0] node9527;
	wire [15-1:0] node9528;
	wire [15-1:0] node9531;
	wire [15-1:0] node9534;
	wire [15-1:0] node9535;
	wire [15-1:0] node9538;
	wire [15-1:0] node9541;
	wire [15-1:0] node9542;
	wire [15-1:0] node9543;
	wire [15-1:0] node9544;
	wire [15-1:0] node9546;
	wire [15-1:0] node9549;
	wire [15-1:0] node9550;
	wire [15-1:0] node9553;
	wire [15-1:0] node9556;
	wire [15-1:0] node9557;
	wire [15-1:0] node9558;
	wire [15-1:0] node9561;
	wire [15-1:0] node9564;
	wire [15-1:0] node9565;
	wire [15-1:0] node9568;
	wire [15-1:0] node9571;
	wire [15-1:0] node9572;
	wire [15-1:0] node9573;
	wire [15-1:0] node9574;
	wire [15-1:0] node9577;
	wire [15-1:0] node9580;
	wire [15-1:0] node9581;
	wire [15-1:0] node9584;
	wire [15-1:0] node9587;
	wire [15-1:0] node9588;
	wire [15-1:0] node9589;
	wire [15-1:0] node9592;
	wire [15-1:0] node9595;
	wire [15-1:0] node9596;
	wire [15-1:0] node9599;
	wire [15-1:0] node9602;
	wire [15-1:0] node9603;
	wire [15-1:0] node9604;
	wire [15-1:0] node9605;
	wire [15-1:0] node9606;
	wire [15-1:0] node9607;
	wire [15-1:0] node9610;
	wire [15-1:0] node9613;
	wire [15-1:0] node9614;
	wire [15-1:0] node9617;
	wire [15-1:0] node9620;
	wire [15-1:0] node9621;
	wire [15-1:0] node9622;
	wire [15-1:0] node9625;
	wire [15-1:0] node9628;
	wire [15-1:0] node9629;
	wire [15-1:0] node9632;
	wire [15-1:0] node9635;
	wire [15-1:0] node9636;
	wire [15-1:0] node9637;
	wire [15-1:0] node9638;
	wire [15-1:0] node9641;
	wire [15-1:0] node9644;
	wire [15-1:0] node9645;
	wire [15-1:0] node9648;
	wire [15-1:0] node9651;
	wire [15-1:0] node9652;
	wire [15-1:0] node9653;
	wire [15-1:0] node9656;
	wire [15-1:0] node9659;
	wire [15-1:0] node9660;
	wire [15-1:0] node9663;
	wire [15-1:0] node9666;
	wire [15-1:0] node9667;
	wire [15-1:0] node9668;
	wire [15-1:0] node9669;
	wire [15-1:0] node9670;
	wire [15-1:0] node9673;
	wire [15-1:0] node9676;
	wire [15-1:0] node9677;
	wire [15-1:0] node9680;
	wire [15-1:0] node9683;
	wire [15-1:0] node9684;
	wire [15-1:0] node9685;
	wire [15-1:0] node9688;
	wire [15-1:0] node9691;
	wire [15-1:0] node9692;
	wire [15-1:0] node9695;
	wire [15-1:0] node9698;
	wire [15-1:0] node9699;
	wire [15-1:0] node9701;
	wire [15-1:0] node9702;
	wire [15-1:0] node9705;
	wire [15-1:0] node9708;
	wire [15-1:0] node9709;
	wire [15-1:0] node9710;
	wire [15-1:0] node9713;
	wire [15-1:0] node9716;
	wire [15-1:0] node9717;
	wire [15-1:0] node9720;
	wire [15-1:0] node9723;
	wire [15-1:0] node9724;
	wire [15-1:0] node9725;
	wire [15-1:0] node9726;
	wire [15-1:0] node9727;
	wire [15-1:0] node9728;
	wire [15-1:0] node9729;
	wire [15-1:0] node9730;
	wire [15-1:0] node9731;
	wire [15-1:0] node9732;
	wire [15-1:0] node9735;
	wire [15-1:0] node9738;
	wire [15-1:0] node9739;
	wire [15-1:0] node9743;
	wire [15-1:0] node9744;
	wire [15-1:0] node9745;
	wire [15-1:0] node9748;
	wire [15-1:0] node9751;
	wire [15-1:0] node9752;
	wire [15-1:0] node9756;
	wire [15-1:0] node9757;
	wire [15-1:0] node9758;
	wire [15-1:0] node9759;
	wire [15-1:0] node9762;
	wire [15-1:0] node9765;
	wire [15-1:0] node9766;
	wire [15-1:0] node9769;
	wire [15-1:0] node9772;
	wire [15-1:0] node9773;
	wire [15-1:0] node9774;
	wire [15-1:0] node9777;
	wire [15-1:0] node9780;
	wire [15-1:0] node9781;
	wire [15-1:0] node9784;
	wire [15-1:0] node9787;
	wire [15-1:0] node9788;
	wire [15-1:0] node9789;
	wire [15-1:0] node9790;
	wire [15-1:0] node9791;
	wire [15-1:0] node9794;
	wire [15-1:0] node9797;
	wire [15-1:0] node9798;
	wire [15-1:0] node9801;
	wire [15-1:0] node9804;
	wire [15-1:0] node9805;
	wire [15-1:0] node9807;
	wire [15-1:0] node9810;
	wire [15-1:0] node9811;
	wire [15-1:0] node9814;
	wire [15-1:0] node9817;
	wire [15-1:0] node9818;
	wire [15-1:0] node9819;
	wire [15-1:0] node9820;
	wire [15-1:0] node9823;
	wire [15-1:0] node9826;
	wire [15-1:0] node9827;
	wire [15-1:0] node9830;
	wire [15-1:0] node9833;
	wire [15-1:0] node9834;
	wire [15-1:0] node9835;
	wire [15-1:0] node9838;
	wire [15-1:0] node9841;
	wire [15-1:0] node9844;
	wire [15-1:0] node9845;
	wire [15-1:0] node9846;
	wire [15-1:0] node9847;
	wire [15-1:0] node9848;
	wire [15-1:0] node9850;
	wire [15-1:0] node9853;
	wire [15-1:0] node9854;
	wire [15-1:0] node9857;
	wire [15-1:0] node9860;
	wire [15-1:0] node9861;
	wire [15-1:0] node9862;
	wire [15-1:0] node9865;
	wire [15-1:0] node9868;
	wire [15-1:0] node9869;
	wire [15-1:0] node9872;
	wire [15-1:0] node9875;
	wire [15-1:0] node9876;
	wire [15-1:0] node9877;
	wire [15-1:0] node9878;
	wire [15-1:0] node9881;
	wire [15-1:0] node9884;
	wire [15-1:0] node9887;
	wire [15-1:0] node9888;
	wire [15-1:0] node9889;
	wire [15-1:0] node9892;
	wire [15-1:0] node9895;
	wire [15-1:0] node9896;
	wire [15-1:0] node9899;
	wire [15-1:0] node9902;
	wire [15-1:0] node9903;
	wire [15-1:0] node9904;
	wire [15-1:0] node9905;
	wire [15-1:0] node9907;
	wire [15-1:0] node9910;
	wire [15-1:0] node9911;
	wire [15-1:0] node9914;
	wire [15-1:0] node9917;
	wire [15-1:0] node9918;
	wire [15-1:0] node9919;
	wire [15-1:0] node9922;
	wire [15-1:0] node9925;
	wire [15-1:0] node9926;
	wire [15-1:0] node9929;
	wire [15-1:0] node9932;
	wire [15-1:0] node9933;
	wire [15-1:0] node9934;
	wire [15-1:0] node9935;
	wire [15-1:0] node9938;
	wire [15-1:0] node9941;
	wire [15-1:0] node9942;
	wire [15-1:0] node9946;
	wire [15-1:0] node9947;
	wire [15-1:0] node9948;
	wire [15-1:0] node9951;
	wire [15-1:0] node9954;
	wire [15-1:0] node9955;
	wire [15-1:0] node9958;
	wire [15-1:0] node9961;
	wire [15-1:0] node9962;
	wire [15-1:0] node9963;
	wire [15-1:0] node9964;
	wire [15-1:0] node9965;
	wire [15-1:0] node9966;
	wire [15-1:0] node9967;
	wire [15-1:0] node9970;
	wire [15-1:0] node9973;
	wire [15-1:0] node9974;
	wire [15-1:0] node9977;
	wire [15-1:0] node9980;
	wire [15-1:0] node9981;
	wire [15-1:0] node9982;
	wire [15-1:0] node9985;
	wire [15-1:0] node9988;
	wire [15-1:0] node9989;
	wire [15-1:0] node9992;
	wire [15-1:0] node9995;
	wire [15-1:0] node9996;
	wire [15-1:0] node9997;
	wire [15-1:0] node9999;
	wire [15-1:0] node10002;
	wire [15-1:0] node10003;
	wire [15-1:0] node10006;
	wire [15-1:0] node10009;
	wire [15-1:0] node10010;
	wire [15-1:0] node10011;
	wire [15-1:0] node10014;
	wire [15-1:0] node10017;
	wire [15-1:0] node10018;
	wire [15-1:0] node10021;
	wire [15-1:0] node10024;
	wire [15-1:0] node10025;
	wire [15-1:0] node10026;
	wire [15-1:0] node10027;
	wire [15-1:0] node10028;
	wire [15-1:0] node10031;
	wire [15-1:0] node10034;
	wire [15-1:0] node10035;
	wire [15-1:0] node10039;
	wire [15-1:0] node10040;
	wire [15-1:0] node10042;
	wire [15-1:0] node10045;
	wire [15-1:0] node10046;
	wire [15-1:0] node10049;
	wire [15-1:0] node10052;
	wire [15-1:0] node10053;
	wire [15-1:0] node10054;
	wire [15-1:0] node10055;
	wire [15-1:0] node10058;
	wire [15-1:0] node10061;
	wire [15-1:0] node10063;
	wire [15-1:0] node10066;
	wire [15-1:0] node10067;
	wire [15-1:0] node10068;
	wire [15-1:0] node10071;
	wire [15-1:0] node10074;
	wire [15-1:0] node10075;
	wire [15-1:0] node10078;
	wire [15-1:0] node10081;
	wire [15-1:0] node10082;
	wire [15-1:0] node10083;
	wire [15-1:0] node10084;
	wire [15-1:0] node10085;
	wire [15-1:0] node10086;
	wire [15-1:0] node10090;
	wire [15-1:0] node10091;
	wire [15-1:0] node10094;
	wire [15-1:0] node10097;
	wire [15-1:0] node10098;
	wire [15-1:0] node10099;
	wire [15-1:0] node10102;
	wire [15-1:0] node10105;
	wire [15-1:0] node10106;
	wire [15-1:0] node10109;
	wire [15-1:0] node10112;
	wire [15-1:0] node10113;
	wire [15-1:0] node10114;
	wire [15-1:0] node10115;
	wire [15-1:0] node10118;
	wire [15-1:0] node10121;
	wire [15-1:0] node10123;
	wire [15-1:0] node10126;
	wire [15-1:0] node10127;
	wire [15-1:0] node10128;
	wire [15-1:0] node10131;
	wire [15-1:0] node10134;
	wire [15-1:0] node10136;
	wire [15-1:0] node10139;
	wire [15-1:0] node10140;
	wire [15-1:0] node10141;
	wire [15-1:0] node10142;
	wire [15-1:0] node10143;
	wire [15-1:0] node10146;
	wire [15-1:0] node10149;
	wire [15-1:0] node10150;
	wire [15-1:0] node10153;
	wire [15-1:0] node10156;
	wire [15-1:0] node10157;
	wire [15-1:0] node10158;
	wire [15-1:0] node10161;
	wire [15-1:0] node10164;
	wire [15-1:0] node10165;
	wire [15-1:0] node10168;
	wire [15-1:0] node10171;
	wire [15-1:0] node10172;
	wire [15-1:0] node10173;
	wire [15-1:0] node10174;
	wire [15-1:0] node10177;
	wire [15-1:0] node10180;
	wire [15-1:0] node10181;
	wire [15-1:0] node10184;
	wire [15-1:0] node10187;
	wire [15-1:0] node10188;
	wire [15-1:0] node10189;
	wire [15-1:0] node10192;
	wire [15-1:0] node10195;
	wire [15-1:0] node10196;
	wire [15-1:0] node10200;
	wire [15-1:0] node10201;
	wire [15-1:0] node10202;
	wire [15-1:0] node10203;
	wire [15-1:0] node10204;
	wire [15-1:0] node10205;
	wire [15-1:0] node10206;
	wire [15-1:0] node10207;
	wire [15-1:0] node10211;
	wire [15-1:0] node10212;
	wire [15-1:0] node10215;
	wire [15-1:0] node10218;
	wire [15-1:0] node10219;
	wire [15-1:0] node10220;
	wire [15-1:0] node10224;
	wire [15-1:0] node10225;
	wire [15-1:0] node10228;
	wire [15-1:0] node10231;
	wire [15-1:0] node10232;
	wire [15-1:0] node10233;
	wire [15-1:0] node10234;
	wire [15-1:0] node10237;
	wire [15-1:0] node10240;
	wire [15-1:0] node10241;
	wire [15-1:0] node10244;
	wire [15-1:0] node10247;
	wire [15-1:0] node10248;
	wire [15-1:0] node10250;
	wire [15-1:0] node10253;
	wire [15-1:0] node10254;
	wire [15-1:0] node10257;
	wire [15-1:0] node10260;
	wire [15-1:0] node10261;
	wire [15-1:0] node10262;
	wire [15-1:0] node10263;
	wire [15-1:0] node10264;
	wire [15-1:0] node10267;
	wire [15-1:0] node10270;
	wire [15-1:0] node10271;
	wire [15-1:0] node10274;
	wire [15-1:0] node10277;
	wire [15-1:0] node10278;
	wire [15-1:0] node10279;
	wire [15-1:0] node10282;
	wire [15-1:0] node10285;
	wire [15-1:0] node10287;
	wire [15-1:0] node10290;
	wire [15-1:0] node10291;
	wire [15-1:0] node10292;
	wire [15-1:0] node10293;
	wire [15-1:0] node10296;
	wire [15-1:0] node10299;
	wire [15-1:0] node10300;
	wire [15-1:0] node10303;
	wire [15-1:0] node10306;
	wire [15-1:0] node10307;
	wire [15-1:0] node10308;
	wire [15-1:0] node10311;
	wire [15-1:0] node10314;
	wire [15-1:0] node10315;
	wire [15-1:0] node10318;
	wire [15-1:0] node10321;
	wire [15-1:0] node10322;
	wire [15-1:0] node10323;
	wire [15-1:0] node10324;
	wire [15-1:0] node10325;
	wire [15-1:0] node10326;
	wire [15-1:0] node10329;
	wire [15-1:0] node10332;
	wire [15-1:0] node10333;
	wire [15-1:0] node10337;
	wire [15-1:0] node10338;
	wire [15-1:0] node10339;
	wire [15-1:0] node10342;
	wire [15-1:0] node10345;
	wire [15-1:0] node10346;
	wire [15-1:0] node10350;
	wire [15-1:0] node10351;
	wire [15-1:0] node10352;
	wire [15-1:0] node10354;
	wire [15-1:0] node10357;
	wire [15-1:0] node10358;
	wire [15-1:0] node10361;
	wire [15-1:0] node10364;
	wire [15-1:0] node10365;
	wire [15-1:0] node10366;
	wire [15-1:0] node10369;
	wire [15-1:0] node10372;
	wire [15-1:0] node10373;
	wire [15-1:0] node10376;
	wire [15-1:0] node10379;
	wire [15-1:0] node10380;
	wire [15-1:0] node10381;
	wire [15-1:0] node10382;
	wire [15-1:0] node10383;
	wire [15-1:0] node10386;
	wire [15-1:0] node10389;
	wire [15-1:0] node10390;
	wire [15-1:0] node10393;
	wire [15-1:0] node10396;
	wire [15-1:0] node10397;
	wire [15-1:0] node10398;
	wire [15-1:0] node10401;
	wire [15-1:0] node10404;
	wire [15-1:0] node10405;
	wire [15-1:0] node10408;
	wire [15-1:0] node10411;
	wire [15-1:0] node10412;
	wire [15-1:0] node10413;
	wire [15-1:0] node10414;
	wire [15-1:0] node10417;
	wire [15-1:0] node10420;
	wire [15-1:0] node10421;
	wire [15-1:0] node10424;
	wire [15-1:0] node10427;
	wire [15-1:0] node10428;
	wire [15-1:0] node10429;
	wire [15-1:0] node10432;
	wire [15-1:0] node10435;
	wire [15-1:0] node10436;
	wire [15-1:0] node10440;
	wire [15-1:0] node10441;
	wire [15-1:0] node10442;
	wire [15-1:0] node10443;
	wire [15-1:0] node10444;
	wire [15-1:0] node10445;
	wire [15-1:0] node10446;
	wire [15-1:0] node10449;
	wire [15-1:0] node10452;
	wire [15-1:0] node10453;
	wire [15-1:0] node10456;
	wire [15-1:0] node10459;
	wire [15-1:0] node10460;
	wire [15-1:0] node10461;
	wire [15-1:0] node10464;
	wire [15-1:0] node10467;
	wire [15-1:0] node10468;
	wire [15-1:0] node10471;
	wire [15-1:0] node10474;
	wire [15-1:0] node10475;
	wire [15-1:0] node10476;
	wire [15-1:0] node10479;
	wire [15-1:0] node10480;
	wire [15-1:0] node10483;
	wire [15-1:0] node10486;
	wire [15-1:0] node10487;
	wire [15-1:0] node10488;
	wire [15-1:0] node10491;
	wire [15-1:0] node10494;
	wire [15-1:0] node10495;
	wire [15-1:0] node10498;
	wire [15-1:0] node10501;
	wire [15-1:0] node10502;
	wire [15-1:0] node10503;
	wire [15-1:0] node10504;
	wire [15-1:0] node10506;
	wire [15-1:0] node10509;
	wire [15-1:0] node10510;
	wire [15-1:0] node10514;
	wire [15-1:0] node10515;
	wire [15-1:0] node10517;
	wire [15-1:0] node10520;
	wire [15-1:0] node10522;
	wire [15-1:0] node10525;
	wire [15-1:0] node10526;
	wire [15-1:0] node10527;
	wire [15-1:0] node10528;
	wire [15-1:0] node10532;
	wire [15-1:0] node10533;
	wire [15-1:0] node10536;
	wire [15-1:0] node10539;
	wire [15-1:0] node10540;
	wire [15-1:0] node10541;
	wire [15-1:0] node10544;
	wire [15-1:0] node10547;
	wire [15-1:0] node10548;
	wire [15-1:0] node10551;
	wire [15-1:0] node10554;
	wire [15-1:0] node10555;
	wire [15-1:0] node10556;
	wire [15-1:0] node10557;
	wire [15-1:0] node10558;
	wire [15-1:0] node10560;
	wire [15-1:0] node10563;
	wire [15-1:0] node10564;
	wire [15-1:0] node10567;
	wire [15-1:0] node10570;
	wire [15-1:0] node10571;
	wire [15-1:0] node10572;
	wire [15-1:0] node10575;
	wire [15-1:0] node10578;
	wire [15-1:0] node10579;
	wire [15-1:0] node10582;
	wire [15-1:0] node10585;
	wire [15-1:0] node10586;
	wire [15-1:0] node10587;
	wire [15-1:0] node10588;
	wire [15-1:0] node10591;
	wire [15-1:0] node10594;
	wire [15-1:0] node10595;
	wire [15-1:0] node10598;
	wire [15-1:0] node10601;
	wire [15-1:0] node10602;
	wire [15-1:0] node10603;
	wire [15-1:0] node10606;
	wire [15-1:0] node10609;
	wire [15-1:0] node10610;
	wire [15-1:0] node10613;
	wire [15-1:0] node10616;
	wire [15-1:0] node10617;
	wire [15-1:0] node10618;
	wire [15-1:0] node10619;
	wire [15-1:0] node10620;
	wire [15-1:0] node10623;
	wire [15-1:0] node10626;
	wire [15-1:0] node10627;
	wire [15-1:0] node10630;
	wire [15-1:0] node10633;
	wire [15-1:0] node10634;
	wire [15-1:0] node10635;
	wire [15-1:0] node10638;
	wire [15-1:0] node10641;
	wire [15-1:0] node10642;
	wire [15-1:0] node10645;
	wire [15-1:0] node10648;
	wire [15-1:0] node10649;
	wire [15-1:0] node10650;
	wire [15-1:0] node10651;
	wire [15-1:0] node10654;
	wire [15-1:0] node10657;
	wire [15-1:0] node10658;
	wire [15-1:0] node10661;
	wire [15-1:0] node10664;
	wire [15-1:0] node10665;
	wire [15-1:0] node10666;
	wire [15-1:0] node10669;
	wire [15-1:0] node10672;
	wire [15-1:0] node10673;
	wire [15-1:0] node10676;
	wire [15-1:0] node10679;
	wire [15-1:0] node10680;
	wire [15-1:0] node10681;
	wire [15-1:0] node10682;
	wire [15-1:0] node10683;
	wire [15-1:0] node10684;
	wire [15-1:0] node10685;
	wire [15-1:0] node10686;
	wire [15-1:0] node10687;
	wire [15-1:0] node10690;
	wire [15-1:0] node10693;
	wire [15-1:0] node10695;
	wire [15-1:0] node10698;
	wire [15-1:0] node10699;
	wire [15-1:0] node10700;
	wire [15-1:0] node10703;
	wire [15-1:0] node10706;
	wire [15-1:0] node10707;
	wire [15-1:0] node10710;
	wire [15-1:0] node10713;
	wire [15-1:0] node10714;
	wire [15-1:0] node10715;
	wire [15-1:0] node10716;
	wire [15-1:0] node10719;
	wire [15-1:0] node10722;
	wire [15-1:0] node10723;
	wire [15-1:0] node10726;
	wire [15-1:0] node10729;
	wire [15-1:0] node10730;
	wire [15-1:0] node10731;
	wire [15-1:0] node10734;
	wire [15-1:0] node10737;
	wire [15-1:0] node10738;
	wire [15-1:0] node10741;
	wire [15-1:0] node10744;
	wire [15-1:0] node10745;
	wire [15-1:0] node10746;
	wire [15-1:0] node10747;
	wire [15-1:0] node10748;
	wire [15-1:0] node10751;
	wire [15-1:0] node10754;
	wire [15-1:0] node10755;
	wire [15-1:0] node10758;
	wire [15-1:0] node10761;
	wire [15-1:0] node10762;
	wire [15-1:0] node10763;
	wire [15-1:0] node10766;
	wire [15-1:0] node10769;
	wire [15-1:0] node10770;
	wire [15-1:0] node10773;
	wire [15-1:0] node10776;
	wire [15-1:0] node10777;
	wire [15-1:0] node10778;
	wire [15-1:0] node10779;
	wire [15-1:0] node10782;
	wire [15-1:0] node10785;
	wire [15-1:0] node10786;
	wire [15-1:0] node10790;
	wire [15-1:0] node10791;
	wire [15-1:0] node10792;
	wire [15-1:0] node10795;
	wire [15-1:0] node10798;
	wire [15-1:0] node10799;
	wire [15-1:0] node10802;
	wire [15-1:0] node10805;
	wire [15-1:0] node10806;
	wire [15-1:0] node10807;
	wire [15-1:0] node10808;
	wire [15-1:0] node10809;
	wire [15-1:0] node10810;
	wire [15-1:0] node10814;
	wire [15-1:0] node10816;
	wire [15-1:0] node10819;
	wire [15-1:0] node10820;
	wire [15-1:0] node10821;
	wire [15-1:0] node10825;
	wire [15-1:0] node10826;
	wire [15-1:0] node10829;
	wire [15-1:0] node10832;
	wire [15-1:0] node10833;
	wire [15-1:0] node10834;
	wire [15-1:0] node10835;
	wire [15-1:0] node10838;
	wire [15-1:0] node10841;
	wire [15-1:0] node10842;
	wire [15-1:0] node10845;
	wire [15-1:0] node10848;
	wire [15-1:0] node10849;
	wire [15-1:0] node10850;
	wire [15-1:0] node10853;
	wire [15-1:0] node10856;
	wire [15-1:0] node10857;
	wire [15-1:0] node10860;
	wire [15-1:0] node10863;
	wire [15-1:0] node10864;
	wire [15-1:0] node10865;
	wire [15-1:0] node10866;
	wire [15-1:0] node10868;
	wire [15-1:0] node10871;
	wire [15-1:0] node10872;
	wire [15-1:0] node10875;
	wire [15-1:0] node10878;
	wire [15-1:0] node10879;
	wire [15-1:0] node10880;
	wire [15-1:0] node10883;
	wire [15-1:0] node10886;
	wire [15-1:0] node10888;
	wire [15-1:0] node10891;
	wire [15-1:0] node10892;
	wire [15-1:0] node10893;
	wire [15-1:0] node10894;
	wire [15-1:0] node10897;
	wire [15-1:0] node10900;
	wire [15-1:0] node10901;
	wire [15-1:0] node10904;
	wire [15-1:0] node10907;
	wire [15-1:0] node10908;
	wire [15-1:0] node10909;
	wire [15-1:0] node10912;
	wire [15-1:0] node10915;
	wire [15-1:0] node10916;
	wire [15-1:0] node10920;
	wire [15-1:0] node10921;
	wire [15-1:0] node10922;
	wire [15-1:0] node10923;
	wire [15-1:0] node10924;
	wire [15-1:0] node10925;
	wire [15-1:0] node10926;
	wire [15-1:0] node10929;
	wire [15-1:0] node10933;
	wire [15-1:0] node10934;
	wire [15-1:0] node10935;
	wire [15-1:0] node10938;
	wire [15-1:0] node10941;
	wire [15-1:0] node10942;
	wire [15-1:0] node10945;
	wire [15-1:0] node10948;
	wire [15-1:0] node10949;
	wire [15-1:0] node10950;
	wire [15-1:0] node10951;
	wire [15-1:0] node10954;
	wire [15-1:0] node10957;
	wire [15-1:0] node10958;
	wire [15-1:0] node10961;
	wire [15-1:0] node10964;
	wire [15-1:0] node10965;
	wire [15-1:0] node10966;
	wire [15-1:0] node10969;
	wire [15-1:0] node10972;
	wire [15-1:0] node10974;
	wire [15-1:0] node10977;
	wire [15-1:0] node10978;
	wire [15-1:0] node10979;
	wire [15-1:0] node10980;
	wire [15-1:0] node10981;
	wire [15-1:0] node10985;
	wire [15-1:0] node10986;
	wire [15-1:0] node10990;
	wire [15-1:0] node10991;
	wire [15-1:0] node10992;
	wire [15-1:0] node10995;
	wire [15-1:0] node10998;
	wire [15-1:0] node10999;
	wire [15-1:0] node11002;
	wire [15-1:0] node11005;
	wire [15-1:0] node11006;
	wire [15-1:0] node11007;
	wire [15-1:0] node11008;
	wire [15-1:0] node11011;
	wire [15-1:0] node11014;
	wire [15-1:0] node11015;
	wire [15-1:0] node11018;
	wire [15-1:0] node11021;
	wire [15-1:0] node11022;
	wire [15-1:0] node11024;
	wire [15-1:0] node11027;
	wire [15-1:0] node11028;
	wire [15-1:0] node11031;
	wire [15-1:0] node11034;
	wire [15-1:0] node11035;
	wire [15-1:0] node11036;
	wire [15-1:0] node11037;
	wire [15-1:0] node11038;
	wire [15-1:0] node11039;
	wire [15-1:0] node11042;
	wire [15-1:0] node11045;
	wire [15-1:0] node11046;
	wire [15-1:0] node11049;
	wire [15-1:0] node11052;
	wire [15-1:0] node11053;
	wire [15-1:0] node11054;
	wire [15-1:0] node11057;
	wire [15-1:0] node11060;
	wire [15-1:0] node11061;
	wire [15-1:0] node11064;
	wire [15-1:0] node11067;
	wire [15-1:0] node11068;
	wire [15-1:0] node11069;
	wire [15-1:0] node11070;
	wire [15-1:0] node11073;
	wire [15-1:0] node11077;
	wire [15-1:0] node11078;
	wire [15-1:0] node11079;
	wire [15-1:0] node11082;
	wire [15-1:0] node11085;
	wire [15-1:0] node11086;
	wire [15-1:0] node11089;
	wire [15-1:0] node11092;
	wire [15-1:0] node11093;
	wire [15-1:0] node11094;
	wire [15-1:0] node11095;
	wire [15-1:0] node11096;
	wire [15-1:0] node11099;
	wire [15-1:0] node11102;
	wire [15-1:0] node11103;
	wire [15-1:0] node11106;
	wire [15-1:0] node11109;
	wire [15-1:0] node11110;
	wire [15-1:0] node11111;
	wire [15-1:0] node11114;
	wire [15-1:0] node11117;
	wire [15-1:0] node11118;
	wire [15-1:0] node11121;
	wire [15-1:0] node11124;
	wire [15-1:0] node11125;
	wire [15-1:0] node11126;
	wire [15-1:0] node11127;
	wire [15-1:0] node11130;
	wire [15-1:0] node11133;
	wire [15-1:0] node11134;
	wire [15-1:0] node11137;
	wire [15-1:0] node11140;
	wire [15-1:0] node11141;
	wire [15-1:0] node11142;
	wire [15-1:0] node11145;
	wire [15-1:0] node11148;
	wire [15-1:0] node11149;
	wire [15-1:0] node11152;
	wire [15-1:0] node11155;
	wire [15-1:0] node11156;
	wire [15-1:0] node11157;
	wire [15-1:0] node11158;
	wire [15-1:0] node11159;
	wire [15-1:0] node11160;
	wire [15-1:0] node11161;
	wire [15-1:0] node11162;
	wire [15-1:0] node11166;
	wire [15-1:0] node11167;
	wire [15-1:0] node11171;
	wire [15-1:0] node11172;
	wire [15-1:0] node11174;
	wire [15-1:0] node11177;
	wire [15-1:0] node11178;
	wire [15-1:0] node11181;
	wire [15-1:0] node11184;
	wire [15-1:0] node11185;
	wire [15-1:0] node11186;
	wire [15-1:0] node11187;
	wire [15-1:0] node11190;
	wire [15-1:0] node11193;
	wire [15-1:0] node11194;
	wire [15-1:0] node11197;
	wire [15-1:0] node11200;
	wire [15-1:0] node11201;
	wire [15-1:0] node11202;
	wire [15-1:0] node11205;
	wire [15-1:0] node11208;
	wire [15-1:0] node11209;
	wire [15-1:0] node11212;
	wire [15-1:0] node11215;
	wire [15-1:0] node11216;
	wire [15-1:0] node11217;
	wire [15-1:0] node11218;
	wire [15-1:0] node11219;
	wire [15-1:0] node11223;
	wire [15-1:0] node11224;
	wire [15-1:0] node11227;
	wire [15-1:0] node11230;
	wire [15-1:0] node11231;
	wire [15-1:0] node11232;
	wire [15-1:0] node11235;
	wire [15-1:0] node11238;
	wire [15-1:0] node11239;
	wire [15-1:0] node11242;
	wire [15-1:0] node11245;
	wire [15-1:0] node11246;
	wire [15-1:0] node11247;
	wire [15-1:0] node11249;
	wire [15-1:0] node11253;
	wire [15-1:0] node11254;
	wire [15-1:0] node11255;
	wire [15-1:0] node11258;
	wire [15-1:0] node11261;
	wire [15-1:0] node11262;
	wire [15-1:0] node11265;
	wire [15-1:0] node11268;
	wire [15-1:0] node11269;
	wire [15-1:0] node11270;
	wire [15-1:0] node11271;
	wire [15-1:0] node11272;
	wire [15-1:0] node11273;
	wire [15-1:0] node11276;
	wire [15-1:0] node11279;
	wire [15-1:0] node11280;
	wire [15-1:0] node11283;
	wire [15-1:0] node11286;
	wire [15-1:0] node11287;
	wire [15-1:0] node11288;
	wire [15-1:0] node11291;
	wire [15-1:0] node11294;
	wire [15-1:0] node11295;
	wire [15-1:0] node11298;
	wire [15-1:0] node11301;
	wire [15-1:0] node11302;
	wire [15-1:0] node11303;
	wire [15-1:0] node11304;
	wire [15-1:0] node11307;
	wire [15-1:0] node11310;
	wire [15-1:0] node11311;
	wire [15-1:0] node11314;
	wire [15-1:0] node11317;
	wire [15-1:0] node11318;
	wire [15-1:0] node11319;
	wire [15-1:0] node11322;
	wire [15-1:0] node11325;
	wire [15-1:0] node11326;
	wire [15-1:0] node11330;
	wire [15-1:0] node11331;
	wire [15-1:0] node11332;
	wire [15-1:0] node11333;
	wire [15-1:0] node11334;
	wire [15-1:0] node11337;
	wire [15-1:0] node11340;
	wire [15-1:0] node11342;
	wire [15-1:0] node11345;
	wire [15-1:0] node11346;
	wire [15-1:0] node11347;
	wire [15-1:0] node11350;
	wire [15-1:0] node11353;
	wire [15-1:0] node11355;
	wire [15-1:0] node11358;
	wire [15-1:0] node11359;
	wire [15-1:0] node11360;
	wire [15-1:0] node11361;
	wire [15-1:0] node11365;
	wire [15-1:0] node11366;
	wire [15-1:0] node11369;
	wire [15-1:0] node11372;
	wire [15-1:0] node11373;
	wire [15-1:0] node11374;
	wire [15-1:0] node11377;
	wire [15-1:0] node11380;
	wire [15-1:0] node11381;
	wire [15-1:0] node11384;
	wire [15-1:0] node11387;
	wire [15-1:0] node11388;
	wire [15-1:0] node11389;
	wire [15-1:0] node11390;
	wire [15-1:0] node11391;
	wire [15-1:0] node11392;
	wire [15-1:0] node11393;
	wire [15-1:0] node11396;
	wire [15-1:0] node11399;
	wire [15-1:0] node11401;
	wire [15-1:0] node11404;
	wire [15-1:0] node11405;
	wire [15-1:0] node11406;
	wire [15-1:0] node11409;
	wire [15-1:0] node11412;
	wire [15-1:0] node11413;
	wire [15-1:0] node11416;
	wire [15-1:0] node11419;
	wire [15-1:0] node11420;
	wire [15-1:0] node11421;
	wire [15-1:0] node11422;
	wire [15-1:0] node11425;
	wire [15-1:0] node11428;
	wire [15-1:0] node11429;
	wire [15-1:0] node11432;
	wire [15-1:0] node11435;
	wire [15-1:0] node11436;
	wire [15-1:0] node11437;
	wire [15-1:0] node11440;
	wire [15-1:0] node11443;
	wire [15-1:0] node11444;
	wire [15-1:0] node11447;
	wire [15-1:0] node11450;
	wire [15-1:0] node11451;
	wire [15-1:0] node11452;
	wire [15-1:0] node11453;
	wire [15-1:0] node11454;
	wire [15-1:0] node11457;
	wire [15-1:0] node11460;
	wire [15-1:0] node11461;
	wire [15-1:0] node11464;
	wire [15-1:0] node11467;
	wire [15-1:0] node11468;
	wire [15-1:0] node11469;
	wire [15-1:0] node11472;
	wire [15-1:0] node11475;
	wire [15-1:0] node11476;
	wire [15-1:0] node11479;
	wire [15-1:0] node11482;
	wire [15-1:0] node11483;
	wire [15-1:0] node11484;
	wire [15-1:0] node11485;
	wire [15-1:0] node11488;
	wire [15-1:0] node11491;
	wire [15-1:0] node11492;
	wire [15-1:0] node11495;
	wire [15-1:0] node11498;
	wire [15-1:0] node11499;
	wire [15-1:0] node11500;
	wire [15-1:0] node11503;
	wire [15-1:0] node11506;
	wire [15-1:0] node11507;
	wire [15-1:0] node11510;
	wire [15-1:0] node11513;
	wire [15-1:0] node11514;
	wire [15-1:0] node11515;
	wire [15-1:0] node11516;
	wire [15-1:0] node11517;
	wire [15-1:0] node11518;
	wire [15-1:0] node11521;
	wire [15-1:0] node11524;
	wire [15-1:0] node11525;
	wire [15-1:0] node11528;
	wire [15-1:0] node11531;
	wire [15-1:0] node11532;
	wire [15-1:0] node11533;
	wire [15-1:0] node11536;
	wire [15-1:0] node11539;
	wire [15-1:0] node11540;
	wire [15-1:0] node11543;
	wire [15-1:0] node11546;
	wire [15-1:0] node11547;
	wire [15-1:0] node11548;
	wire [15-1:0] node11549;
	wire [15-1:0] node11552;
	wire [15-1:0] node11555;
	wire [15-1:0] node11556;
	wire [15-1:0] node11559;
	wire [15-1:0] node11562;
	wire [15-1:0] node11563;
	wire [15-1:0] node11564;
	wire [15-1:0] node11567;
	wire [15-1:0] node11570;
	wire [15-1:0] node11571;
	wire [15-1:0] node11574;
	wire [15-1:0] node11577;
	wire [15-1:0] node11578;
	wire [15-1:0] node11579;
	wire [15-1:0] node11580;
	wire [15-1:0] node11581;
	wire [15-1:0] node11585;
	wire [15-1:0] node11586;
	wire [15-1:0] node11589;
	wire [15-1:0] node11592;
	wire [15-1:0] node11593;
	wire [15-1:0] node11594;
	wire [15-1:0] node11597;
	wire [15-1:0] node11600;
	wire [15-1:0] node11602;
	wire [15-1:0] node11605;
	wire [15-1:0] node11606;
	wire [15-1:0] node11607;
	wire [15-1:0] node11609;
	wire [15-1:0] node11612;
	wire [15-1:0] node11613;
	wire [15-1:0] node11616;
	wire [15-1:0] node11619;
	wire [15-1:0] node11620;
	wire [15-1:0] node11621;
	wire [15-1:0] node11624;
	wire [15-1:0] node11627;
	wire [15-1:0] node11628;
	wire [15-1:0] node11631;
	wire [15-1:0] node11634;
	wire [15-1:0] node11635;
	wire [15-1:0] node11636;
	wire [15-1:0] node11637;
	wire [15-1:0] node11638;
	wire [15-1:0] node11639;
	wire [15-1:0] node11640;
	wire [15-1:0] node11641;
	wire [15-1:0] node11642;
	wire [15-1:0] node11643;
	wire [15-1:0] node11644;
	wire [15-1:0] node11647;
	wire [15-1:0] node11650;
	wire [15-1:0] node11651;
	wire [15-1:0] node11654;
	wire [15-1:0] node11657;
	wire [15-1:0] node11658;
	wire [15-1:0] node11659;
	wire [15-1:0] node11662;
	wire [15-1:0] node11665;
	wire [15-1:0] node11666;
	wire [15-1:0] node11669;
	wire [15-1:0] node11672;
	wire [15-1:0] node11673;
	wire [15-1:0] node11674;
	wire [15-1:0] node11676;
	wire [15-1:0] node11679;
	wire [15-1:0] node11680;
	wire [15-1:0] node11683;
	wire [15-1:0] node11686;
	wire [15-1:0] node11687;
	wire [15-1:0] node11688;
	wire [15-1:0] node11691;
	wire [15-1:0] node11694;
	wire [15-1:0] node11695;
	wire [15-1:0] node11698;
	wire [15-1:0] node11701;
	wire [15-1:0] node11702;
	wire [15-1:0] node11703;
	wire [15-1:0] node11704;
	wire [15-1:0] node11705;
	wire [15-1:0] node11708;
	wire [15-1:0] node11711;
	wire [15-1:0] node11712;
	wire [15-1:0] node11715;
	wire [15-1:0] node11718;
	wire [15-1:0] node11719;
	wire [15-1:0] node11720;
	wire [15-1:0] node11723;
	wire [15-1:0] node11726;
	wire [15-1:0] node11727;
	wire [15-1:0] node11730;
	wire [15-1:0] node11733;
	wire [15-1:0] node11734;
	wire [15-1:0] node11735;
	wire [15-1:0] node11736;
	wire [15-1:0] node11739;
	wire [15-1:0] node11742;
	wire [15-1:0] node11743;
	wire [15-1:0] node11746;
	wire [15-1:0] node11749;
	wire [15-1:0] node11750;
	wire [15-1:0] node11751;
	wire [15-1:0] node11754;
	wire [15-1:0] node11757;
	wire [15-1:0] node11758;
	wire [15-1:0] node11761;
	wire [15-1:0] node11764;
	wire [15-1:0] node11765;
	wire [15-1:0] node11766;
	wire [15-1:0] node11767;
	wire [15-1:0] node11768;
	wire [15-1:0] node11769;
	wire [15-1:0] node11772;
	wire [15-1:0] node11775;
	wire [15-1:0] node11776;
	wire [15-1:0] node11779;
	wire [15-1:0] node11782;
	wire [15-1:0] node11783;
	wire [15-1:0] node11784;
	wire [15-1:0] node11787;
	wire [15-1:0] node11790;
	wire [15-1:0] node11791;
	wire [15-1:0] node11794;
	wire [15-1:0] node11797;
	wire [15-1:0] node11798;
	wire [15-1:0] node11799;
	wire [15-1:0] node11800;
	wire [15-1:0] node11803;
	wire [15-1:0] node11806;
	wire [15-1:0] node11807;
	wire [15-1:0] node11811;
	wire [15-1:0] node11812;
	wire [15-1:0] node11813;
	wire [15-1:0] node11816;
	wire [15-1:0] node11819;
	wire [15-1:0] node11821;
	wire [15-1:0] node11824;
	wire [15-1:0] node11825;
	wire [15-1:0] node11826;
	wire [15-1:0] node11827;
	wire [15-1:0] node11828;
	wire [15-1:0] node11831;
	wire [15-1:0] node11834;
	wire [15-1:0] node11835;
	wire [15-1:0] node11838;
	wire [15-1:0] node11841;
	wire [15-1:0] node11842;
	wire [15-1:0] node11843;
	wire [15-1:0] node11846;
	wire [15-1:0] node11849;
	wire [15-1:0] node11850;
	wire [15-1:0] node11853;
	wire [15-1:0] node11856;
	wire [15-1:0] node11857;
	wire [15-1:0] node11858;
	wire [15-1:0] node11859;
	wire [15-1:0] node11862;
	wire [15-1:0] node11865;
	wire [15-1:0] node11866;
	wire [15-1:0] node11869;
	wire [15-1:0] node11872;
	wire [15-1:0] node11873;
	wire [15-1:0] node11874;
	wire [15-1:0] node11877;
	wire [15-1:0] node11880;
	wire [15-1:0] node11882;
	wire [15-1:0] node11885;
	wire [15-1:0] node11886;
	wire [15-1:0] node11887;
	wire [15-1:0] node11888;
	wire [15-1:0] node11889;
	wire [15-1:0] node11890;
	wire [15-1:0] node11891;
	wire [15-1:0] node11894;
	wire [15-1:0] node11897;
	wire [15-1:0] node11898;
	wire [15-1:0] node11901;
	wire [15-1:0] node11904;
	wire [15-1:0] node11905;
	wire [15-1:0] node11906;
	wire [15-1:0] node11909;
	wire [15-1:0] node11912;
	wire [15-1:0] node11913;
	wire [15-1:0] node11916;
	wire [15-1:0] node11919;
	wire [15-1:0] node11920;
	wire [15-1:0] node11921;
	wire [15-1:0] node11922;
	wire [15-1:0] node11925;
	wire [15-1:0] node11928;
	wire [15-1:0] node11929;
	wire [15-1:0] node11932;
	wire [15-1:0] node11935;
	wire [15-1:0] node11936;
	wire [15-1:0] node11937;
	wire [15-1:0] node11940;
	wire [15-1:0] node11943;
	wire [15-1:0] node11944;
	wire [15-1:0] node11948;
	wire [15-1:0] node11949;
	wire [15-1:0] node11950;
	wire [15-1:0] node11951;
	wire [15-1:0] node11952;
	wire [15-1:0] node11955;
	wire [15-1:0] node11958;
	wire [15-1:0] node11959;
	wire [15-1:0] node11962;
	wire [15-1:0] node11965;
	wire [15-1:0] node11966;
	wire [15-1:0] node11967;
	wire [15-1:0] node11970;
	wire [15-1:0] node11973;
	wire [15-1:0] node11974;
	wire [15-1:0] node11978;
	wire [15-1:0] node11979;
	wire [15-1:0] node11980;
	wire [15-1:0] node11981;
	wire [15-1:0] node11984;
	wire [15-1:0] node11987;
	wire [15-1:0] node11988;
	wire [15-1:0] node11991;
	wire [15-1:0] node11994;
	wire [15-1:0] node11995;
	wire [15-1:0] node11997;
	wire [15-1:0] node12000;
	wire [15-1:0] node12001;
	wire [15-1:0] node12004;
	wire [15-1:0] node12007;
	wire [15-1:0] node12008;
	wire [15-1:0] node12009;
	wire [15-1:0] node12010;
	wire [15-1:0] node12011;
	wire [15-1:0] node12012;
	wire [15-1:0] node12015;
	wire [15-1:0] node12018;
	wire [15-1:0] node12019;
	wire [15-1:0] node12022;
	wire [15-1:0] node12025;
	wire [15-1:0] node12026;
	wire [15-1:0] node12027;
	wire [15-1:0] node12030;
	wire [15-1:0] node12033;
	wire [15-1:0] node12034;
	wire [15-1:0] node12037;
	wire [15-1:0] node12040;
	wire [15-1:0] node12041;
	wire [15-1:0] node12042;
	wire [15-1:0] node12043;
	wire [15-1:0] node12046;
	wire [15-1:0] node12049;
	wire [15-1:0] node12050;
	wire [15-1:0] node12053;
	wire [15-1:0] node12056;
	wire [15-1:0] node12057;
	wire [15-1:0] node12058;
	wire [15-1:0] node12062;
	wire [15-1:0] node12063;
	wire [15-1:0] node12066;
	wire [15-1:0] node12069;
	wire [15-1:0] node12070;
	wire [15-1:0] node12071;
	wire [15-1:0] node12072;
	wire [15-1:0] node12074;
	wire [15-1:0] node12077;
	wire [15-1:0] node12078;
	wire [15-1:0] node12081;
	wire [15-1:0] node12084;
	wire [15-1:0] node12085;
	wire [15-1:0] node12086;
	wire [15-1:0] node12089;
	wire [15-1:0] node12092;
	wire [15-1:0] node12093;
	wire [15-1:0] node12096;
	wire [15-1:0] node12099;
	wire [15-1:0] node12100;
	wire [15-1:0] node12101;
	wire [15-1:0] node12102;
	wire [15-1:0] node12105;
	wire [15-1:0] node12108;
	wire [15-1:0] node12109;
	wire [15-1:0] node12112;
	wire [15-1:0] node12115;
	wire [15-1:0] node12116;
	wire [15-1:0] node12117;
	wire [15-1:0] node12120;
	wire [15-1:0] node12123;
	wire [15-1:0] node12125;
	wire [15-1:0] node12128;
	wire [15-1:0] node12129;
	wire [15-1:0] node12130;
	wire [15-1:0] node12131;
	wire [15-1:0] node12132;
	wire [15-1:0] node12133;
	wire [15-1:0] node12134;
	wire [15-1:0] node12135;
	wire [15-1:0] node12139;
	wire [15-1:0] node12140;
	wire [15-1:0] node12143;
	wire [15-1:0] node12146;
	wire [15-1:0] node12147;
	wire [15-1:0] node12148;
	wire [15-1:0] node12151;
	wire [15-1:0] node12154;
	wire [15-1:0] node12155;
	wire [15-1:0] node12158;
	wire [15-1:0] node12161;
	wire [15-1:0] node12162;
	wire [15-1:0] node12163;
	wire [15-1:0] node12164;
	wire [15-1:0] node12167;
	wire [15-1:0] node12170;
	wire [15-1:0] node12171;
	wire [15-1:0] node12174;
	wire [15-1:0] node12177;
	wire [15-1:0] node12178;
	wire [15-1:0] node12179;
	wire [15-1:0] node12182;
	wire [15-1:0] node12185;
	wire [15-1:0] node12186;
	wire [15-1:0] node12190;
	wire [15-1:0] node12191;
	wire [15-1:0] node12192;
	wire [15-1:0] node12193;
	wire [15-1:0] node12194;
	wire [15-1:0] node12197;
	wire [15-1:0] node12200;
	wire [15-1:0] node12201;
	wire [15-1:0] node12204;
	wire [15-1:0] node12207;
	wire [15-1:0] node12208;
	wire [15-1:0] node12209;
	wire [15-1:0] node12212;
	wire [15-1:0] node12215;
	wire [15-1:0] node12216;
	wire [15-1:0] node12219;
	wire [15-1:0] node12222;
	wire [15-1:0] node12223;
	wire [15-1:0] node12224;
	wire [15-1:0] node12225;
	wire [15-1:0] node12228;
	wire [15-1:0] node12231;
	wire [15-1:0] node12232;
	wire [15-1:0] node12235;
	wire [15-1:0] node12238;
	wire [15-1:0] node12239;
	wire [15-1:0] node12241;
	wire [15-1:0] node12244;
	wire [15-1:0] node12245;
	wire [15-1:0] node12248;
	wire [15-1:0] node12251;
	wire [15-1:0] node12252;
	wire [15-1:0] node12253;
	wire [15-1:0] node12254;
	wire [15-1:0] node12255;
	wire [15-1:0] node12256;
	wire [15-1:0] node12259;
	wire [15-1:0] node12262;
	wire [15-1:0] node12263;
	wire [15-1:0] node12266;
	wire [15-1:0] node12269;
	wire [15-1:0] node12270;
	wire [15-1:0] node12271;
	wire [15-1:0] node12274;
	wire [15-1:0] node12277;
	wire [15-1:0] node12278;
	wire [15-1:0] node12281;
	wire [15-1:0] node12284;
	wire [15-1:0] node12285;
	wire [15-1:0] node12286;
	wire [15-1:0] node12287;
	wire [15-1:0] node12290;
	wire [15-1:0] node12293;
	wire [15-1:0] node12294;
	wire [15-1:0] node12297;
	wire [15-1:0] node12300;
	wire [15-1:0] node12301;
	wire [15-1:0] node12302;
	wire [15-1:0] node12305;
	wire [15-1:0] node12308;
	wire [15-1:0] node12309;
	wire [15-1:0] node12312;
	wire [15-1:0] node12315;
	wire [15-1:0] node12316;
	wire [15-1:0] node12317;
	wire [15-1:0] node12318;
	wire [15-1:0] node12320;
	wire [15-1:0] node12323;
	wire [15-1:0] node12324;
	wire [15-1:0] node12327;
	wire [15-1:0] node12330;
	wire [15-1:0] node12331;
	wire [15-1:0] node12332;
	wire [15-1:0] node12335;
	wire [15-1:0] node12338;
	wire [15-1:0] node12339;
	wire [15-1:0] node12342;
	wire [15-1:0] node12345;
	wire [15-1:0] node12346;
	wire [15-1:0] node12347;
	wire [15-1:0] node12348;
	wire [15-1:0] node12352;
	wire [15-1:0] node12353;
	wire [15-1:0] node12356;
	wire [15-1:0] node12359;
	wire [15-1:0] node12360;
	wire [15-1:0] node12361;
	wire [15-1:0] node12364;
	wire [15-1:0] node12367;
	wire [15-1:0] node12368;
	wire [15-1:0] node12371;
	wire [15-1:0] node12374;
	wire [15-1:0] node12375;
	wire [15-1:0] node12376;
	wire [15-1:0] node12377;
	wire [15-1:0] node12378;
	wire [15-1:0] node12379;
	wire [15-1:0] node12380;
	wire [15-1:0] node12384;
	wire [15-1:0] node12385;
	wire [15-1:0] node12388;
	wire [15-1:0] node12391;
	wire [15-1:0] node12392;
	wire [15-1:0] node12393;
	wire [15-1:0] node12396;
	wire [15-1:0] node12399;
	wire [15-1:0] node12400;
	wire [15-1:0] node12403;
	wire [15-1:0] node12406;
	wire [15-1:0] node12407;
	wire [15-1:0] node12408;
	wire [15-1:0] node12409;
	wire [15-1:0] node12412;
	wire [15-1:0] node12415;
	wire [15-1:0] node12416;
	wire [15-1:0] node12419;
	wire [15-1:0] node12422;
	wire [15-1:0] node12423;
	wire [15-1:0] node12424;
	wire [15-1:0] node12427;
	wire [15-1:0] node12430;
	wire [15-1:0] node12431;
	wire [15-1:0] node12434;
	wire [15-1:0] node12437;
	wire [15-1:0] node12438;
	wire [15-1:0] node12439;
	wire [15-1:0] node12440;
	wire [15-1:0] node12441;
	wire [15-1:0] node12444;
	wire [15-1:0] node12447;
	wire [15-1:0] node12448;
	wire [15-1:0] node12451;
	wire [15-1:0] node12454;
	wire [15-1:0] node12455;
	wire [15-1:0] node12457;
	wire [15-1:0] node12460;
	wire [15-1:0] node12463;
	wire [15-1:0] node12464;
	wire [15-1:0] node12465;
	wire [15-1:0] node12466;
	wire [15-1:0] node12469;
	wire [15-1:0] node12472;
	wire [15-1:0] node12473;
	wire [15-1:0] node12476;
	wire [15-1:0] node12479;
	wire [15-1:0] node12480;
	wire [15-1:0] node12481;
	wire [15-1:0] node12484;
	wire [15-1:0] node12487;
	wire [15-1:0] node12488;
	wire [15-1:0] node12491;
	wire [15-1:0] node12494;
	wire [15-1:0] node12495;
	wire [15-1:0] node12496;
	wire [15-1:0] node12497;
	wire [15-1:0] node12498;
	wire [15-1:0] node12499;
	wire [15-1:0] node12502;
	wire [15-1:0] node12505;
	wire [15-1:0] node12506;
	wire [15-1:0] node12509;
	wire [15-1:0] node12512;
	wire [15-1:0] node12513;
	wire [15-1:0] node12514;
	wire [15-1:0] node12517;
	wire [15-1:0] node12520;
	wire [15-1:0] node12521;
	wire [15-1:0] node12524;
	wire [15-1:0] node12527;
	wire [15-1:0] node12528;
	wire [15-1:0] node12529;
	wire [15-1:0] node12530;
	wire [15-1:0] node12533;
	wire [15-1:0] node12536;
	wire [15-1:0] node12537;
	wire [15-1:0] node12540;
	wire [15-1:0] node12543;
	wire [15-1:0] node12544;
	wire [15-1:0] node12545;
	wire [15-1:0] node12548;
	wire [15-1:0] node12551;
	wire [15-1:0] node12552;
	wire [15-1:0] node12555;
	wire [15-1:0] node12558;
	wire [15-1:0] node12559;
	wire [15-1:0] node12560;
	wire [15-1:0] node12561;
	wire [15-1:0] node12562;
	wire [15-1:0] node12565;
	wire [15-1:0] node12568;
	wire [15-1:0] node12569;
	wire [15-1:0] node12572;
	wire [15-1:0] node12575;
	wire [15-1:0] node12576;
	wire [15-1:0] node12577;
	wire [15-1:0] node12580;
	wire [15-1:0] node12583;
	wire [15-1:0] node12584;
	wire [15-1:0] node12587;
	wire [15-1:0] node12590;
	wire [15-1:0] node12591;
	wire [15-1:0] node12592;
	wire [15-1:0] node12593;
	wire [15-1:0] node12596;
	wire [15-1:0] node12599;
	wire [15-1:0] node12601;
	wire [15-1:0] node12604;
	wire [15-1:0] node12605;
	wire [15-1:0] node12606;
	wire [15-1:0] node12609;
	wire [15-1:0] node12612;
	wire [15-1:0] node12613;
	wire [15-1:0] node12616;
	wire [15-1:0] node12619;
	wire [15-1:0] node12620;
	wire [15-1:0] node12621;
	wire [15-1:0] node12622;
	wire [15-1:0] node12623;
	wire [15-1:0] node12624;
	wire [15-1:0] node12625;
	wire [15-1:0] node12626;
	wire [15-1:0] node12627;
	wire [15-1:0] node12631;
	wire [15-1:0] node12632;
	wire [15-1:0] node12635;
	wire [15-1:0] node12638;
	wire [15-1:0] node12639;
	wire [15-1:0] node12640;
	wire [15-1:0] node12643;
	wire [15-1:0] node12646;
	wire [15-1:0] node12647;
	wire [15-1:0] node12651;
	wire [15-1:0] node12652;
	wire [15-1:0] node12653;
	wire [15-1:0] node12654;
	wire [15-1:0] node12657;
	wire [15-1:0] node12660;
	wire [15-1:0] node12661;
	wire [15-1:0] node12664;
	wire [15-1:0] node12667;
	wire [15-1:0] node12668;
	wire [15-1:0] node12669;
	wire [15-1:0] node12672;
	wire [15-1:0] node12675;
	wire [15-1:0] node12676;
	wire [15-1:0] node12679;
	wire [15-1:0] node12682;
	wire [15-1:0] node12683;
	wire [15-1:0] node12684;
	wire [15-1:0] node12685;
	wire [15-1:0] node12686;
	wire [15-1:0] node12689;
	wire [15-1:0] node12692;
	wire [15-1:0] node12693;
	wire [15-1:0] node12697;
	wire [15-1:0] node12698;
	wire [15-1:0] node12699;
	wire [15-1:0] node12702;
	wire [15-1:0] node12705;
	wire [15-1:0] node12706;
	wire [15-1:0] node12709;
	wire [15-1:0] node12712;
	wire [15-1:0] node12713;
	wire [15-1:0] node12714;
	wire [15-1:0] node12715;
	wire [15-1:0] node12718;
	wire [15-1:0] node12721;
	wire [15-1:0] node12722;
	wire [15-1:0] node12725;
	wire [15-1:0] node12728;
	wire [15-1:0] node12729;
	wire [15-1:0] node12730;
	wire [15-1:0] node12733;
	wire [15-1:0] node12736;
	wire [15-1:0] node12737;
	wire [15-1:0] node12740;
	wire [15-1:0] node12743;
	wire [15-1:0] node12744;
	wire [15-1:0] node12745;
	wire [15-1:0] node12746;
	wire [15-1:0] node12747;
	wire [15-1:0] node12748;
	wire [15-1:0] node12751;
	wire [15-1:0] node12754;
	wire [15-1:0] node12755;
	wire [15-1:0] node12758;
	wire [15-1:0] node12761;
	wire [15-1:0] node12762;
	wire [15-1:0] node12763;
	wire [15-1:0] node12766;
	wire [15-1:0] node12769;
	wire [15-1:0] node12770;
	wire [15-1:0] node12773;
	wire [15-1:0] node12776;
	wire [15-1:0] node12777;
	wire [15-1:0] node12778;
	wire [15-1:0] node12779;
	wire [15-1:0] node12782;
	wire [15-1:0] node12785;
	wire [15-1:0] node12786;
	wire [15-1:0] node12789;
	wire [15-1:0] node12792;
	wire [15-1:0] node12793;
	wire [15-1:0] node12794;
	wire [15-1:0] node12797;
	wire [15-1:0] node12800;
	wire [15-1:0] node12802;
	wire [15-1:0] node12805;
	wire [15-1:0] node12806;
	wire [15-1:0] node12807;
	wire [15-1:0] node12808;
	wire [15-1:0] node12810;
	wire [15-1:0] node12813;
	wire [15-1:0] node12814;
	wire [15-1:0] node12818;
	wire [15-1:0] node12819;
	wire [15-1:0] node12821;
	wire [15-1:0] node12824;
	wire [15-1:0] node12825;
	wire [15-1:0] node12828;
	wire [15-1:0] node12831;
	wire [15-1:0] node12832;
	wire [15-1:0] node12833;
	wire [15-1:0] node12834;
	wire [15-1:0] node12837;
	wire [15-1:0] node12840;
	wire [15-1:0] node12841;
	wire [15-1:0] node12844;
	wire [15-1:0] node12847;
	wire [15-1:0] node12848;
	wire [15-1:0] node12849;
	wire [15-1:0] node12852;
	wire [15-1:0] node12855;
	wire [15-1:0] node12856;
	wire [15-1:0] node12860;
	wire [15-1:0] node12861;
	wire [15-1:0] node12862;
	wire [15-1:0] node12863;
	wire [15-1:0] node12864;
	wire [15-1:0] node12865;
	wire [15-1:0] node12866;
	wire [15-1:0] node12869;
	wire [15-1:0] node12872;
	wire [15-1:0] node12873;
	wire [15-1:0] node12876;
	wire [15-1:0] node12879;
	wire [15-1:0] node12880;
	wire [15-1:0] node12881;
	wire [15-1:0] node12884;
	wire [15-1:0] node12887;
	wire [15-1:0] node12888;
	wire [15-1:0] node12891;
	wire [15-1:0] node12894;
	wire [15-1:0] node12895;
	wire [15-1:0] node12896;
	wire [15-1:0] node12897;
	wire [15-1:0] node12900;
	wire [15-1:0] node12903;
	wire [15-1:0] node12904;
	wire [15-1:0] node12907;
	wire [15-1:0] node12910;
	wire [15-1:0] node12911;
	wire [15-1:0] node12912;
	wire [15-1:0] node12915;
	wire [15-1:0] node12918;
	wire [15-1:0] node12921;
	wire [15-1:0] node12922;
	wire [15-1:0] node12923;
	wire [15-1:0] node12924;
	wire [15-1:0] node12926;
	wire [15-1:0] node12929;
	wire [15-1:0] node12930;
	wire [15-1:0] node12933;
	wire [15-1:0] node12936;
	wire [15-1:0] node12937;
	wire [15-1:0] node12938;
	wire [15-1:0] node12941;
	wire [15-1:0] node12944;
	wire [15-1:0] node12945;
	wire [15-1:0] node12948;
	wire [15-1:0] node12951;
	wire [15-1:0] node12952;
	wire [15-1:0] node12953;
	wire [15-1:0] node12954;
	wire [15-1:0] node12957;
	wire [15-1:0] node12960;
	wire [15-1:0] node12961;
	wire [15-1:0] node12964;
	wire [15-1:0] node12967;
	wire [15-1:0] node12968;
	wire [15-1:0] node12969;
	wire [15-1:0] node12972;
	wire [15-1:0] node12975;
	wire [15-1:0] node12976;
	wire [15-1:0] node12979;
	wire [15-1:0] node12982;
	wire [15-1:0] node12983;
	wire [15-1:0] node12984;
	wire [15-1:0] node12985;
	wire [15-1:0] node12986;
	wire [15-1:0] node12987;
	wire [15-1:0] node12990;
	wire [15-1:0] node12993;
	wire [15-1:0] node12994;
	wire [15-1:0] node12997;
	wire [15-1:0] node13000;
	wire [15-1:0] node13001;
	wire [15-1:0] node13002;
	wire [15-1:0] node13005;
	wire [15-1:0] node13008;
	wire [15-1:0] node13009;
	wire [15-1:0] node13012;
	wire [15-1:0] node13015;
	wire [15-1:0] node13016;
	wire [15-1:0] node13017;
	wire [15-1:0] node13019;
	wire [15-1:0] node13022;
	wire [15-1:0] node13023;
	wire [15-1:0] node13026;
	wire [15-1:0] node13029;
	wire [15-1:0] node13030;
	wire [15-1:0] node13032;
	wire [15-1:0] node13035;
	wire [15-1:0] node13036;
	wire [15-1:0] node13039;
	wire [15-1:0] node13042;
	wire [15-1:0] node13043;
	wire [15-1:0] node13044;
	wire [15-1:0] node13045;
	wire [15-1:0] node13046;
	wire [15-1:0] node13050;
	wire [15-1:0] node13051;
	wire [15-1:0] node13054;
	wire [15-1:0] node13057;
	wire [15-1:0] node13058;
	wire [15-1:0] node13059;
	wire [15-1:0] node13062;
	wire [15-1:0] node13065;
	wire [15-1:0] node13066;
	wire [15-1:0] node13069;
	wire [15-1:0] node13072;
	wire [15-1:0] node13073;
	wire [15-1:0] node13074;
	wire [15-1:0] node13075;
	wire [15-1:0] node13078;
	wire [15-1:0] node13081;
	wire [15-1:0] node13083;
	wire [15-1:0] node13086;
	wire [15-1:0] node13087;
	wire [15-1:0] node13088;
	wire [15-1:0] node13091;
	wire [15-1:0] node13094;
	wire [15-1:0] node13095;
	wire [15-1:0] node13098;
	wire [15-1:0] node13101;
	wire [15-1:0] node13102;
	wire [15-1:0] node13103;
	wire [15-1:0] node13104;
	wire [15-1:0] node13105;
	wire [15-1:0] node13106;
	wire [15-1:0] node13107;
	wire [15-1:0] node13108;
	wire [15-1:0] node13112;
	wire [15-1:0] node13113;
	wire [15-1:0] node13116;
	wire [15-1:0] node13119;
	wire [15-1:0] node13120;
	wire [15-1:0] node13121;
	wire [15-1:0] node13124;
	wire [15-1:0] node13127;
	wire [15-1:0] node13128;
	wire [15-1:0] node13131;
	wire [15-1:0] node13134;
	wire [15-1:0] node13135;
	wire [15-1:0] node13136;
	wire [15-1:0] node13137;
	wire [15-1:0] node13140;
	wire [15-1:0] node13143;
	wire [15-1:0] node13144;
	wire [15-1:0] node13147;
	wire [15-1:0] node13150;
	wire [15-1:0] node13151;
	wire [15-1:0] node13152;
	wire [15-1:0] node13155;
	wire [15-1:0] node13158;
	wire [15-1:0] node13159;
	wire [15-1:0] node13162;
	wire [15-1:0] node13165;
	wire [15-1:0] node13166;
	wire [15-1:0] node13167;
	wire [15-1:0] node13168;
	wire [15-1:0] node13169;
	wire [15-1:0] node13172;
	wire [15-1:0] node13175;
	wire [15-1:0] node13176;
	wire [15-1:0] node13179;
	wire [15-1:0] node13182;
	wire [15-1:0] node13183;
	wire [15-1:0] node13184;
	wire [15-1:0] node13187;
	wire [15-1:0] node13190;
	wire [15-1:0] node13191;
	wire [15-1:0] node13194;
	wire [15-1:0] node13197;
	wire [15-1:0] node13198;
	wire [15-1:0] node13199;
	wire [15-1:0] node13200;
	wire [15-1:0] node13203;
	wire [15-1:0] node13206;
	wire [15-1:0] node13207;
	wire [15-1:0] node13210;
	wire [15-1:0] node13213;
	wire [15-1:0] node13214;
	wire [15-1:0] node13215;
	wire [15-1:0] node13218;
	wire [15-1:0] node13221;
	wire [15-1:0] node13222;
	wire [15-1:0] node13225;
	wire [15-1:0] node13228;
	wire [15-1:0] node13229;
	wire [15-1:0] node13230;
	wire [15-1:0] node13231;
	wire [15-1:0] node13232;
	wire [15-1:0] node13233;
	wire [15-1:0] node13236;
	wire [15-1:0] node13239;
	wire [15-1:0] node13240;
	wire [15-1:0] node13244;
	wire [15-1:0] node13245;
	wire [15-1:0] node13246;
	wire [15-1:0] node13249;
	wire [15-1:0] node13252;
	wire [15-1:0] node13253;
	wire [15-1:0] node13256;
	wire [15-1:0] node13259;
	wire [15-1:0] node13260;
	wire [15-1:0] node13261;
	wire [15-1:0] node13262;
	wire [15-1:0] node13265;
	wire [15-1:0] node13268;
	wire [15-1:0] node13269;
	wire [15-1:0] node13272;
	wire [15-1:0] node13275;
	wire [15-1:0] node13276;
	wire [15-1:0] node13277;
	wire [15-1:0] node13280;
	wire [15-1:0] node13283;
	wire [15-1:0] node13284;
	wire [15-1:0] node13287;
	wire [15-1:0] node13290;
	wire [15-1:0] node13291;
	wire [15-1:0] node13292;
	wire [15-1:0] node13293;
	wire [15-1:0] node13294;
	wire [15-1:0] node13297;
	wire [15-1:0] node13300;
	wire [15-1:0] node13301;
	wire [15-1:0] node13304;
	wire [15-1:0] node13307;
	wire [15-1:0] node13308;
	wire [15-1:0] node13309;
	wire [15-1:0] node13312;
	wire [15-1:0] node13315;
	wire [15-1:0] node13316;
	wire [15-1:0] node13319;
	wire [15-1:0] node13322;
	wire [15-1:0] node13323;
	wire [15-1:0] node13324;
	wire [15-1:0] node13325;
	wire [15-1:0] node13328;
	wire [15-1:0] node13331;
	wire [15-1:0] node13332;
	wire [15-1:0] node13335;
	wire [15-1:0] node13338;
	wire [15-1:0] node13339;
	wire [15-1:0] node13340;
	wire [15-1:0] node13343;
	wire [15-1:0] node13346;
	wire [15-1:0] node13347;
	wire [15-1:0] node13350;
	wire [15-1:0] node13353;
	wire [15-1:0] node13354;
	wire [15-1:0] node13355;
	wire [15-1:0] node13356;
	wire [15-1:0] node13357;
	wire [15-1:0] node13358;
	wire [15-1:0] node13359;
	wire [15-1:0] node13362;
	wire [15-1:0] node13365;
	wire [15-1:0] node13366;
	wire [15-1:0] node13369;
	wire [15-1:0] node13372;
	wire [15-1:0] node13373;
	wire [15-1:0] node13374;
	wire [15-1:0] node13377;
	wire [15-1:0] node13380;
	wire [15-1:0] node13381;
	wire [15-1:0] node13384;
	wire [15-1:0] node13387;
	wire [15-1:0] node13388;
	wire [15-1:0] node13389;
	wire [15-1:0] node13391;
	wire [15-1:0] node13394;
	wire [15-1:0] node13395;
	wire [15-1:0] node13398;
	wire [15-1:0] node13401;
	wire [15-1:0] node13402;
	wire [15-1:0] node13403;
	wire [15-1:0] node13406;
	wire [15-1:0] node13409;
	wire [15-1:0] node13410;
	wire [15-1:0] node13413;
	wire [15-1:0] node13416;
	wire [15-1:0] node13417;
	wire [15-1:0] node13418;
	wire [15-1:0] node13419;
	wire [15-1:0] node13420;
	wire [15-1:0] node13423;
	wire [15-1:0] node13426;
	wire [15-1:0] node13428;
	wire [15-1:0] node13431;
	wire [15-1:0] node13432;
	wire [15-1:0] node13433;
	wire [15-1:0] node13436;
	wire [15-1:0] node13439;
	wire [15-1:0] node13440;
	wire [15-1:0] node13443;
	wire [15-1:0] node13446;
	wire [15-1:0] node13447;
	wire [15-1:0] node13448;
	wire [15-1:0] node13449;
	wire [15-1:0] node13452;
	wire [15-1:0] node13455;
	wire [15-1:0] node13456;
	wire [15-1:0] node13459;
	wire [15-1:0] node13462;
	wire [15-1:0] node13463;
	wire [15-1:0] node13464;
	wire [15-1:0] node13467;
	wire [15-1:0] node13470;
	wire [15-1:0] node13471;
	wire [15-1:0] node13474;
	wire [15-1:0] node13477;
	wire [15-1:0] node13478;
	wire [15-1:0] node13479;
	wire [15-1:0] node13480;
	wire [15-1:0] node13481;
	wire [15-1:0] node13482;
	wire [15-1:0] node13485;
	wire [15-1:0] node13488;
	wire [15-1:0] node13489;
	wire [15-1:0] node13492;
	wire [15-1:0] node13495;
	wire [15-1:0] node13496;
	wire [15-1:0] node13497;
	wire [15-1:0] node13500;
	wire [15-1:0] node13503;
	wire [15-1:0] node13505;
	wire [15-1:0] node13508;
	wire [15-1:0] node13509;
	wire [15-1:0] node13510;
	wire [15-1:0] node13511;
	wire [15-1:0] node13514;
	wire [15-1:0] node13517;
	wire [15-1:0] node13518;
	wire [15-1:0] node13521;
	wire [15-1:0] node13524;
	wire [15-1:0] node13525;
	wire [15-1:0] node13526;
	wire [15-1:0] node13529;
	wire [15-1:0] node13532;
	wire [15-1:0] node13533;
	wire [15-1:0] node13536;
	wire [15-1:0] node13539;
	wire [15-1:0] node13540;
	wire [15-1:0] node13541;
	wire [15-1:0] node13542;
	wire [15-1:0] node13544;
	wire [15-1:0] node13547;
	wire [15-1:0] node13549;
	wire [15-1:0] node13552;
	wire [15-1:0] node13553;
	wire [15-1:0] node13554;
	wire [15-1:0] node13557;
	wire [15-1:0] node13560;
	wire [15-1:0] node13561;
	wire [15-1:0] node13564;
	wire [15-1:0] node13567;
	wire [15-1:0] node13568;
	wire [15-1:0] node13569;
	wire [15-1:0] node13570;
	wire [15-1:0] node13573;
	wire [15-1:0] node13576;
	wire [15-1:0] node13578;
	wire [15-1:0] node13581;
	wire [15-1:0] node13582;
	wire [15-1:0] node13583;
	wire [15-1:0] node13586;
	wire [15-1:0] node13589;
	wire [15-1:0] node13590;
	wire [15-1:0] node13593;
	wire [15-1:0] node13596;
	wire [15-1:0] node13597;
	wire [15-1:0] node13598;
	wire [15-1:0] node13599;
	wire [15-1:0] node13600;
	wire [15-1:0] node13601;
	wire [15-1:0] node13602;
	wire [15-1:0] node13603;
	wire [15-1:0] node13604;
	wire [15-1:0] node13605;
	wire [15-1:0] node13608;
	wire [15-1:0] node13611;
	wire [15-1:0] node13612;
	wire [15-1:0] node13615;
	wire [15-1:0] node13618;
	wire [15-1:0] node13619;
	wire [15-1:0] node13621;
	wire [15-1:0] node13624;
	wire [15-1:0] node13625;
	wire [15-1:0] node13628;
	wire [15-1:0] node13631;
	wire [15-1:0] node13632;
	wire [15-1:0] node13633;
	wire [15-1:0] node13634;
	wire [15-1:0] node13637;
	wire [15-1:0] node13640;
	wire [15-1:0] node13641;
	wire [15-1:0] node13644;
	wire [15-1:0] node13647;
	wire [15-1:0] node13648;
	wire [15-1:0] node13649;
	wire [15-1:0] node13652;
	wire [15-1:0] node13655;
	wire [15-1:0] node13656;
	wire [15-1:0] node13659;
	wire [15-1:0] node13662;
	wire [15-1:0] node13663;
	wire [15-1:0] node13664;
	wire [15-1:0] node13665;
	wire [15-1:0] node13666;
	wire [15-1:0] node13670;
	wire [15-1:0] node13671;
	wire [15-1:0] node13674;
	wire [15-1:0] node13677;
	wire [15-1:0] node13678;
	wire [15-1:0] node13679;
	wire [15-1:0] node13682;
	wire [15-1:0] node13685;
	wire [15-1:0] node13686;
	wire [15-1:0] node13689;
	wire [15-1:0] node13692;
	wire [15-1:0] node13693;
	wire [15-1:0] node13694;
	wire [15-1:0] node13695;
	wire [15-1:0] node13698;
	wire [15-1:0] node13701;
	wire [15-1:0] node13702;
	wire [15-1:0] node13705;
	wire [15-1:0] node13708;
	wire [15-1:0] node13709;
	wire [15-1:0] node13710;
	wire [15-1:0] node13713;
	wire [15-1:0] node13716;
	wire [15-1:0] node13717;
	wire [15-1:0] node13721;
	wire [15-1:0] node13722;
	wire [15-1:0] node13723;
	wire [15-1:0] node13724;
	wire [15-1:0] node13725;
	wire [15-1:0] node13726;
	wire [15-1:0] node13729;
	wire [15-1:0] node13732;
	wire [15-1:0] node13734;
	wire [15-1:0] node13737;
	wire [15-1:0] node13738;
	wire [15-1:0] node13739;
	wire [15-1:0] node13742;
	wire [15-1:0] node13745;
	wire [15-1:0] node13746;
	wire [15-1:0] node13749;
	wire [15-1:0] node13752;
	wire [15-1:0] node13753;
	wire [15-1:0] node13754;
	wire [15-1:0] node13756;
	wire [15-1:0] node13759;
	wire [15-1:0] node13760;
	wire [15-1:0] node13764;
	wire [15-1:0] node13765;
	wire [15-1:0] node13766;
	wire [15-1:0] node13769;
	wire [15-1:0] node13772;
	wire [15-1:0] node13773;
	wire [15-1:0] node13776;
	wire [15-1:0] node13779;
	wire [15-1:0] node13780;
	wire [15-1:0] node13781;
	wire [15-1:0] node13782;
	wire [15-1:0] node13783;
	wire [15-1:0] node13786;
	wire [15-1:0] node13789;
	wire [15-1:0] node13790;
	wire [15-1:0] node13794;
	wire [15-1:0] node13795;
	wire [15-1:0] node13796;
	wire [15-1:0] node13799;
	wire [15-1:0] node13802;
	wire [15-1:0] node13803;
	wire [15-1:0] node13806;
	wire [15-1:0] node13809;
	wire [15-1:0] node13810;
	wire [15-1:0] node13811;
	wire [15-1:0] node13812;
	wire [15-1:0] node13815;
	wire [15-1:0] node13818;
	wire [15-1:0] node13819;
	wire [15-1:0] node13822;
	wire [15-1:0] node13825;
	wire [15-1:0] node13826;
	wire [15-1:0] node13828;
	wire [15-1:0] node13831;
	wire [15-1:0] node13832;
	wire [15-1:0] node13835;
	wire [15-1:0] node13838;
	wire [15-1:0] node13839;
	wire [15-1:0] node13840;
	wire [15-1:0] node13841;
	wire [15-1:0] node13842;
	wire [15-1:0] node13843;
	wire [15-1:0] node13844;
	wire [15-1:0] node13847;
	wire [15-1:0] node13850;
	wire [15-1:0] node13851;
	wire [15-1:0] node13854;
	wire [15-1:0] node13857;
	wire [15-1:0] node13858;
	wire [15-1:0] node13859;
	wire [15-1:0] node13862;
	wire [15-1:0] node13865;
	wire [15-1:0] node13866;
	wire [15-1:0] node13869;
	wire [15-1:0] node13872;
	wire [15-1:0] node13873;
	wire [15-1:0] node13874;
	wire [15-1:0] node13875;
	wire [15-1:0] node13878;
	wire [15-1:0] node13881;
	wire [15-1:0] node13882;
	wire [15-1:0] node13885;
	wire [15-1:0] node13888;
	wire [15-1:0] node13889;
	wire [15-1:0] node13890;
	wire [15-1:0] node13893;
	wire [15-1:0] node13896;
	wire [15-1:0] node13897;
	wire [15-1:0] node13900;
	wire [15-1:0] node13903;
	wire [15-1:0] node13904;
	wire [15-1:0] node13905;
	wire [15-1:0] node13906;
	wire [15-1:0] node13908;
	wire [15-1:0] node13911;
	wire [15-1:0] node13912;
	wire [15-1:0] node13916;
	wire [15-1:0] node13917;
	wire [15-1:0] node13918;
	wire [15-1:0] node13921;
	wire [15-1:0] node13924;
	wire [15-1:0] node13925;
	wire [15-1:0] node13928;
	wire [15-1:0] node13931;
	wire [15-1:0] node13932;
	wire [15-1:0] node13933;
	wire [15-1:0] node13934;
	wire [15-1:0] node13937;
	wire [15-1:0] node13940;
	wire [15-1:0] node13941;
	wire [15-1:0] node13944;
	wire [15-1:0] node13947;
	wire [15-1:0] node13948;
	wire [15-1:0] node13949;
	wire [15-1:0] node13952;
	wire [15-1:0] node13955;
	wire [15-1:0] node13956;
	wire [15-1:0] node13959;
	wire [15-1:0] node13962;
	wire [15-1:0] node13963;
	wire [15-1:0] node13964;
	wire [15-1:0] node13965;
	wire [15-1:0] node13966;
	wire [15-1:0] node13967;
	wire [15-1:0] node13970;
	wire [15-1:0] node13973;
	wire [15-1:0] node13974;
	wire [15-1:0] node13977;
	wire [15-1:0] node13980;
	wire [15-1:0] node13981;
	wire [15-1:0] node13983;
	wire [15-1:0] node13986;
	wire [15-1:0] node13987;
	wire [15-1:0] node13990;
	wire [15-1:0] node13993;
	wire [15-1:0] node13994;
	wire [15-1:0] node13995;
	wire [15-1:0] node13996;
	wire [15-1:0] node13999;
	wire [15-1:0] node14002;
	wire [15-1:0] node14003;
	wire [15-1:0] node14006;
	wire [15-1:0] node14009;
	wire [15-1:0] node14010;
	wire [15-1:0] node14011;
	wire [15-1:0] node14014;
	wire [15-1:0] node14017;
	wire [15-1:0] node14018;
	wire [15-1:0] node14021;
	wire [15-1:0] node14024;
	wire [15-1:0] node14025;
	wire [15-1:0] node14026;
	wire [15-1:0] node14027;
	wire [15-1:0] node14028;
	wire [15-1:0] node14031;
	wire [15-1:0] node14034;
	wire [15-1:0] node14035;
	wire [15-1:0] node14039;
	wire [15-1:0] node14040;
	wire [15-1:0] node14041;
	wire [15-1:0] node14044;
	wire [15-1:0] node14047;
	wire [15-1:0] node14048;
	wire [15-1:0] node14051;
	wire [15-1:0] node14054;
	wire [15-1:0] node14055;
	wire [15-1:0] node14056;
	wire [15-1:0] node14057;
	wire [15-1:0] node14060;
	wire [15-1:0] node14063;
	wire [15-1:0] node14064;
	wire [15-1:0] node14067;
	wire [15-1:0] node14070;
	wire [15-1:0] node14071;
	wire [15-1:0] node14072;
	wire [15-1:0] node14075;
	wire [15-1:0] node14078;
	wire [15-1:0] node14079;
	wire [15-1:0] node14082;
	wire [15-1:0] node14085;
	wire [15-1:0] node14086;
	wire [15-1:0] node14087;
	wire [15-1:0] node14088;
	wire [15-1:0] node14089;
	wire [15-1:0] node14090;
	wire [15-1:0] node14091;
	wire [15-1:0] node14092;
	wire [15-1:0] node14095;
	wire [15-1:0] node14098;
	wire [15-1:0] node14099;
	wire [15-1:0] node14103;
	wire [15-1:0] node14104;
	wire [15-1:0] node14105;
	wire [15-1:0] node14108;
	wire [15-1:0] node14111;
	wire [15-1:0] node14112;
	wire [15-1:0] node14115;
	wire [15-1:0] node14118;
	wire [15-1:0] node14119;
	wire [15-1:0] node14120;
	wire [15-1:0] node14121;
	wire [15-1:0] node14124;
	wire [15-1:0] node14127;
	wire [15-1:0] node14128;
	wire [15-1:0] node14131;
	wire [15-1:0] node14134;
	wire [15-1:0] node14135;
	wire [15-1:0] node14137;
	wire [15-1:0] node14140;
	wire [15-1:0] node14141;
	wire [15-1:0] node14144;
	wire [15-1:0] node14147;
	wire [15-1:0] node14148;
	wire [15-1:0] node14149;
	wire [15-1:0] node14150;
	wire [15-1:0] node14151;
	wire [15-1:0] node14154;
	wire [15-1:0] node14157;
	wire [15-1:0] node14158;
	wire [15-1:0] node14161;
	wire [15-1:0] node14164;
	wire [15-1:0] node14165;
	wire [15-1:0] node14166;
	wire [15-1:0] node14169;
	wire [15-1:0] node14172;
	wire [15-1:0] node14173;
	wire [15-1:0] node14176;
	wire [15-1:0] node14179;
	wire [15-1:0] node14180;
	wire [15-1:0] node14181;
	wire [15-1:0] node14182;
	wire [15-1:0] node14185;
	wire [15-1:0] node14188;
	wire [15-1:0] node14189;
	wire [15-1:0] node14192;
	wire [15-1:0] node14195;
	wire [15-1:0] node14196;
	wire [15-1:0] node14197;
	wire [15-1:0] node14200;
	wire [15-1:0] node14203;
	wire [15-1:0] node14204;
	wire [15-1:0] node14207;
	wire [15-1:0] node14210;
	wire [15-1:0] node14211;
	wire [15-1:0] node14212;
	wire [15-1:0] node14213;
	wire [15-1:0] node14214;
	wire [15-1:0] node14215;
	wire [15-1:0] node14218;
	wire [15-1:0] node14221;
	wire [15-1:0] node14222;
	wire [15-1:0] node14225;
	wire [15-1:0] node14228;
	wire [15-1:0] node14229;
	wire [15-1:0] node14231;
	wire [15-1:0] node14234;
	wire [15-1:0] node14235;
	wire [15-1:0] node14239;
	wire [15-1:0] node14240;
	wire [15-1:0] node14241;
	wire [15-1:0] node14242;
	wire [15-1:0] node14245;
	wire [15-1:0] node14248;
	wire [15-1:0] node14249;
	wire [15-1:0] node14252;
	wire [15-1:0] node14255;
	wire [15-1:0] node14256;
	wire [15-1:0] node14257;
	wire [15-1:0] node14260;
	wire [15-1:0] node14263;
	wire [15-1:0] node14264;
	wire [15-1:0] node14267;
	wire [15-1:0] node14270;
	wire [15-1:0] node14271;
	wire [15-1:0] node14272;
	wire [15-1:0] node14273;
	wire [15-1:0] node14274;
	wire [15-1:0] node14277;
	wire [15-1:0] node14280;
	wire [15-1:0] node14281;
	wire [15-1:0] node14285;
	wire [15-1:0] node14286;
	wire [15-1:0] node14287;
	wire [15-1:0] node14290;
	wire [15-1:0] node14293;
	wire [15-1:0] node14294;
	wire [15-1:0] node14297;
	wire [15-1:0] node14300;
	wire [15-1:0] node14301;
	wire [15-1:0] node14302;
	wire [15-1:0] node14303;
	wire [15-1:0] node14306;
	wire [15-1:0] node14309;
	wire [15-1:0] node14310;
	wire [15-1:0] node14313;
	wire [15-1:0] node14316;
	wire [15-1:0] node14317;
	wire [15-1:0] node14318;
	wire [15-1:0] node14321;
	wire [15-1:0] node14324;
	wire [15-1:0] node14325;
	wire [15-1:0] node14328;
	wire [15-1:0] node14331;
	wire [15-1:0] node14332;
	wire [15-1:0] node14333;
	wire [15-1:0] node14334;
	wire [15-1:0] node14335;
	wire [15-1:0] node14336;
	wire [15-1:0] node14337;
	wire [15-1:0] node14340;
	wire [15-1:0] node14343;
	wire [15-1:0] node14344;
	wire [15-1:0] node14347;
	wire [15-1:0] node14350;
	wire [15-1:0] node14351;
	wire [15-1:0] node14352;
	wire [15-1:0] node14355;
	wire [15-1:0] node14358;
	wire [15-1:0] node14359;
	wire [15-1:0] node14362;
	wire [15-1:0] node14365;
	wire [15-1:0] node14366;
	wire [15-1:0] node14367;
	wire [15-1:0] node14368;
	wire [15-1:0] node14371;
	wire [15-1:0] node14374;
	wire [15-1:0] node14375;
	wire [15-1:0] node14379;
	wire [15-1:0] node14380;
	wire [15-1:0] node14381;
	wire [15-1:0] node14384;
	wire [15-1:0] node14387;
	wire [15-1:0] node14388;
	wire [15-1:0] node14391;
	wire [15-1:0] node14394;
	wire [15-1:0] node14395;
	wire [15-1:0] node14396;
	wire [15-1:0] node14397;
	wire [15-1:0] node14398;
	wire [15-1:0] node14401;
	wire [15-1:0] node14404;
	wire [15-1:0] node14405;
	wire [15-1:0] node14408;
	wire [15-1:0] node14411;
	wire [15-1:0] node14412;
	wire [15-1:0] node14414;
	wire [15-1:0] node14417;
	wire [15-1:0] node14418;
	wire [15-1:0] node14421;
	wire [15-1:0] node14424;
	wire [15-1:0] node14425;
	wire [15-1:0] node14426;
	wire [15-1:0] node14427;
	wire [15-1:0] node14430;
	wire [15-1:0] node14433;
	wire [15-1:0] node14434;
	wire [15-1:0] node14437;
	wire [15-1:0] node14440;
	wire [15-1:0] node14441;
	wire [15-1:0] node14444;
	wire [15-1:0] node14445;
	wire [15-1:0] node14448;
	wire [15-1:0] node14451;
	wire [15-1:0] node14452;
	wire [15-1:0] node14453;
	wire [15-1:0] node14454;
	wire [15-1:0] node14455;
	wire [15-1:0] node14457;
	wire [15-1:0] node14460;
	wire [15-1:0] node14461;
	wire [15-1:0] node14464;
	wire [15-1:0] node14467;
	wire [15-1:0] node14468;
	wire [15-1:0] node14469;
	wire [15-1:0] node14472;
	wire [15-1:0] node14475;
	wire [15-1:0] node14476;
	wire [15-1:0] node14479;
	wire [15-1:0] node14482;
	wire [15-1:0] node14483;
	wire [15-1:0] node14484;
	wire [15-1:0] node14485;
	wire [15-1:0] node14488;
	wire [15-1:0] node14491;
	wire [15-1:0] node14492;
	wire [15-1:0] node14495;
	wire [15-1:0] node14498;
	wire [15-1:0] node14499;
	wire [15-1:0] node14500;
	wire [15-1:0] node14503;
	wire [15-1:0] node14506;
	wire [15-1:0] node14507;
	wire [15-1:0] node14511;
	wire [15-1:0] node14512;
	wire [15-1:0] node14513;
	wire [15-1:0] node14514;
	wire [15-1:0] node14515;
	wire [15-1:0] node14518;
	wire [15-1:0] node14521;
	wire [15-1:0] node14522;
	wire [15-1:0] node14525;
	wire [15-1:0] node14528;
	wire [15-1:0] node14529;
	wire [15-1:0] node14530;
	wire [15-1:0] node14533;
	wire [15-1:0] node14536;
	wire [15-1:0] node14537;
	wire [15-1:0] node14540;
	wire [15-1:0] node14543;
	wire [15-1:0] node14544;
	wire [15-1:0] node14545;
	wire [15-1:0] node14546;
	wire [15-1:0] node14549;
	wire [15-1:0] node14552;
	wire [15-1:0] node14553;
	wire [15-1:0] node14556;
	wire [15-1:0] node14559;
	wire [15-1:0] node14560;
	wire [15-1:0] node14561;
	wire [15-1:0] node14564;
	wire [15-1:0] node14567;
	wire [15-1:0] node14568;
	wire [15-1:0] node14571;
	wire [15-1:0] node14574;
	wire [15-1:0] node14575;
	wire [15-1:0] node14576;
	wire [15-1:0] node14577;
	wire [15-1:0] node14578;
	wire [15-1:0] node14579;
	wire [15-1:0] node14580;
	wire [15-1:0] node14581;
	wire [15-1:0] node14582;
	wire [15-1:0] node14585;
	wire [15-1:0] node14588;
	wire [15-1:0] node14589;
	wire [15-1:0] node14592;
	wire [15-1:0] node14595;
	wire [15-1:0] node14596;
	wire [15-1:0] node14597;
	wire [15-1:0] node14600;
	wire [15-1:0] node14603;
	wire [15-1:0] node14604;
	wire [15-1:0] node14608;
	wire [15-1:0] node14609;
	wire [15-1:0] node14610;
	wire [15-1:0] node14611;
	wire [15-1:0] node14614;
	wire [15-1:0] node14617;
	wire [15-1:0] node14618;
	wire [15-1:0] node14621;
	wire [15-1:0] node14624;
	wire [15-1:0] node14625;
	wire [15-1:0] node14626;
	wire [15-1:0] node14629;
	wire [15-1:0] node14632;
	wire [15-1:0] node14633;
	wire [15-1:0] node14636;
	wire [15-1:0] node14639;
	wire [15-1:0] node14640;
	wire [15-1:0] node14641;
	wire [15-1:0] node14642;
	wire [15-1:0] node14643;
	wire [15-1:0] node14646;
	wire [15-1:0] node14649;
	wire [15-1:0] node14650;
	wire [15-1:0] node14653;
	wire [15-1:0] node14656;
	wire [15-1:0] node14657;
	wire [15-1:0] node14658;
	wire [15-1:0] node14661;
	wire [15-1:0] node14664;
	wire [15-1:0] node14665;
	wire [15-1:0] node14668;
	wire [15-1:0] node14671;
	wire [15-1:0] node14672;
	wire [15-1:0] node14673;
	wire [15-1:0] node14675;
	wire [15-1:0] node14678;
	wire [15-1:0] node14679;
	wire [15-1:0] node14682;
	wire [15-1:0] node14685;
	wire [15-1:0] node14686;
	wire [15-1:0] node14687;
	wire [15-1:0] node14690;
	wire [15-1:0] node14693;
	wire [15-1:0] node14694;
	wire [15-1:0] node14697;
	wire [15-1:0] node14700;
	wire [15-1:0] node14701;
	wire [15-1:0] node14702;
	wire [15-1:0] node14703;
	wire [15-1:0] node14704;
	wire [15-1:0] node14705;
	wire [15-1:0] node14708;
	wire [15-1:0] node14711;
	wire [15-1:0] node14712;
	wire [15-1:0] node14715;
	wire [15-1:0] node14718;
	wire [15-1:0] node14719;
	wire [15-1:0] node14720;
	wire [15-1:0] node14723;
	wire [15-1:0] node14726;
	wire [15-1:0] node14727;
	wire [15-1:0] node14730;
	wire [15-1:0] node14733;
	wire [15-1:0] node14734;
	wire [15-1:0] node14735;
	wire [15-1:0] node14736;
	wire [15-1:0] node14739;
	wire [15-1:0] node14742;
	wire [15-1:0] node14744;
	wire [15-1:0] node14747;
	wire [15-1:0] node14748;
	wire [15-1:0] node14749;
	wire [15-1:0] node14752;
	wire [15-1:0] node14755;
	wire [15-1:0] node14756;
	wire [15-1:0] node14759;
	wire [15-1:0] node14762;
	wire [15-1:0] node14763;
	wire [15-1:0] node14764;
	wire [15-1:0] node14765;
	wire [15-1:0] node14766;
	wire [15-1:0] node14769;
	wire [15-1:0] node14772;
	wire [15-1:0] node14773;
	wire [15-1:0] node14776;
	wire [15-1:0] node14779;
	wire [15-1:0] node14780;
	wire [15-1:0] node14781;
	wire [15-1:0] node14784;
	wire [15-1:0] node14787;
	wire [15-1:0] node14788;
	wire [15-1:0] node14791;
	wire [15-1:0] node14794;
	wire [15-1:0] node14795;
	wire [15-1:0] node14796;
	wire [15-1:0] node14797;
	wire [15-1:0] node14800;
	wire [15-1:0] node14803;
	wire [15-1:0] node14804;
	wire [15-1:0] node14807;
	wire [15-1:0] node14810;
	wire [15-1:0] node14811;
	wire [15-1:0] node14812;
	wire [15-1:0] node14815;
	wire [15-1:0] node14818;
	wire [15-1:0] node14819;
	wire [15-1:0] node14822;
	wire [15-1:0] node14825;
	wire [15-1:0] node14826;
	wire [15-1:0] node14827;
	wire [15-1:0] node14828;
	wire [15-1:0] node14829;
	wire [15-1:0] node14830;
	wire [15-1:0] node14831;
	wire [15-1:0] node14834;
	wire [15-1:0] node14837;
	wire [15-1:0] node14838;
	wire [15-1:0] node14841;
	wire [15-1:0] node14844;
	wire [15-1:0] node14845;
	wire [15-1:0] node14846;
	wire [15-1:0] node14849;
	wire [15-1:0] node14852;
	wire [15-1:0] node14853;
	wire [15-1:0] node14856;
	wire [15-1:0] node14859;
	wire [15-1:0] node14860;
	wire [15-1:0] node14861;
	wire [15-1:0] node14862;
	wire [15-1:0] node14865;
	wire [15-1:0] node14868;
	wire [15-1:0] node14870;
	wire [15-1:0] node14873;
	wire [15-1:0] node14874;
	wire [15-1:0] node14875;
	wire [15-1:0] node14878;
	wire [15-1:0] node14881;
	wire [15-1:0] node14882;
	wire [15-1:0] node14885;
	wire [15-1:0] node14888;
	wire [15-1:0] node14889;
	wire [15-1:0] node14890;
	wire [15-1:0] node14891;
	wire [15-1:0] node14892;
	wire [15-1:0] node14895;
	wire [15-1:0] node14898;
	wire [15-1:0] node14899;
	wire [15-1:0] node14902;
	wire [15-1:0] node14905;
	wire [15-1:0] node14906;
	wire [15-1:0] node14907;
	wire [15-1:0] node14910;
	wire [15-1:0] node14913;
	wire [15-1:0] node14914;
	wire [15-1:0] node14917;
	wire [15-1:0] node14920;
	wire [15-1:0] node14921;
	wire [15-1:0] node14922;
	wire [15-1:0] node14923;
	wire [15-1:0] node14926;
	wire [15-1:0] node14929;
	wire [15-1:0] node14930;
	wire [15-1:0] node14933;
	wire [15-1:0] node14936;
	wire [15-1:0] node14937;
	wire [15-1:0] node14938;
	wire [15-1:0] node14941;
	wire [15-1:0] node14944;
	wire [15-1:0] node14945;
	wire [15-1:0] node14948;
	wire [15-1:0] node14951;
	wire [15-1:0] node14952;
	wire [15-1:0] node14953;
	wire [15-1:0] node14954;
	wire [15-1:0] node14955;
	wire [15-1:0] node14956;
	wire [15-1:0] node14959;
	wire [15-1:0] node14962;
	wire [15-1:0] node14963;
	wire [15-1:0] node14966;
	wire [15-1:0] node14969;
	wire [15-1:0] node14970;
	wire [15-1:0] node14971;
	wire [15-1:0] node14975;
	wire [15-1:0] node14978;
	wire [15-1:0] node14979;
	wire [15-1:0] node14980;
	wire [15-1:0] node14981;
	wire [15-1:0] node14984;
	wire [15-1:0] node14987;
	wire [15-1:0] node14988;
	wire [15-1:0] node14991;
	wire [15-1:0] node14994;
	wire [15-1:0] node14995;
	wire [15-1:0] node14996;
	wire [15-1:0] node14999;
	wire [15-1:0] node15002;
	wire [15-1:0] node15003;
	wire [15-1:0] node15006;
	wire [15-1:0] node15009;
	wire [15-1:0] node15010;
	wire [15-1:0] node15011;
	wire [15-1:0] node15012;
	wire [15-1:0] node15013;
	wire [15-1:0] node15016;
	wire [15-1:0] node15019;
	wire [15-1:0] node15020;
	wire [15-1:0] node15023;
	wire [15-1:0] node15026;
	wire [15-1:0] node15027;
	wire [15-1:0] node15028;
	wire [15-1:0] node15031;
	wire [15-1:0] node15034;
	wire [15-1:0] node15035;
	wire [15-1:0] node15038;
	wire [15-1:0] node15041;
	wire [15-1:0] node15042;
	wire [15-1:0] node15043;
	wire [15-1:0] node15044;
	wire [15-1:0] node15047;
	wire [15-1:0] node15050;
	wire [15-1:0] node15051;
	wire [15-1:0] node15054;
	wire [15-1:0] node15057;
	wire [15-1:0] node15058;
	wire [15-1:0] node15059;
	wire [15-1:0] node15062;
	wire [15-1:0] node15065;
	wire [15-1:0] node15066;
	wire [15-1:0] node15069;
	wire [15-1:0] node15072;
	wire [15-1:0] node15073;
	wire [15-1:0] node15074;
	wire [15-1:0] node15075;
	wire [15-1:0] node15076;
	wire [15-1:0] node15077;
	wire [15-1:0] node15078;
	wire [15-1:0] node15079;
	wire [15-1:0] node15082;
	wire [15-1:0] node15085;
	wire [15-1:0] node15086;
	wire [15-1:0] node15089;
	wire [15-1:0] node15092;
	wire [15-1:0] node15093;
	wire [15-1:0] node15094;
	wire [15-1:0] node15097;
	wire [15-1:0] node15100;
	wire [15-1:0] node15101;
	wire [15-1:0] node15104;
	wire [15-1:0] node15107;
	wire [15-1:0] node15108;
	wire [15-1:0] node15109;
	wire [15-1:0] node15110;
	wire [15-1:0] node15113;
	wire [15-1:0] node15116;
	wire [15-1:0] node15117;
	wire [15-1:0] node15121;
	wire [15-1:0] node15122;
	wire [15-1:0] node15123;
	wire [15-1:0] node15126;
	wire [15-1:0] node15129;
	wire [15-1:0] node15130;
	wire [15-1:0] node15133;
	wire [15-1:0] node15136;
	wire [15-1:0] node15137;
	wire [15-1:0] node15138;
	wire [15-1:0] node15139;
	wire [15-1:0] node15140;
	wire [15-1:0] node15144;
	wire [15-1:0] node15145;
	wire [15-1:0] node15148;
	wire [15-1:0] node15151;
	wire [15-1:0] node15152;
	wire [15-1:0] node15153;
	wire [15-1:0] node15157;
	wire [15-1:0] node15158;
	wire [15-1:0] node15162;
	wire [15-1:0] node15163;
	wire [15-1:0] node15164;
	wire [15-1:0] node15165;
	wire [15-1:0] node15168;
	wire [15-1:0] node15171;
	wire [15-1:0] node15172;
	wire [15-1:0] node15175;
	wire [15-1:0] node15178;
	wire [15-1:0] node15179;
	wire [15-1:0] node15180;
	wire [15-1:0] node15183;
	wire [15-1:0] node15186;
	wire [15-1:0] node15187;
	wire [15-1:0] node15190;
	wire [15-1:0] node15193;
	wire [15-1:0] node15194;
	wire [15-1:0] node15195;
	wire [15-1:0] node15196;
	wire [15-1:0] node15197;
	wire [15-1:0] node15198;
	wire [15-1:0] node15202;
	wire [15-1:0] node15203;
	wire [15-1:0] node15207;
	wire [15-1:0] node15208;
	wire [15-1:0] node15209;
	wire [15-1:0] node15212;
	wire [15-1:0] node15215;
	wire [15-1:0] node15216;
	wire [15-1:0] node15219;
	wire [15-1:0] node15222;
	wire [15-1:0] node15223;
	wire [15-1:0] node15224;
	wire [15-1:0] node15225;
	wire [15-1:0] node15229;
	wire [15-1:0] node15230;
	wire [15-1:0] node15233;
	wire [15-1:0] node15236;
	wire [15-1:0] node15237;
	wire [15-1:0] node15238;
	wire [15-1:0] node15241;
	wire [15-1:0] node15244;
	wire [15-1:0] node15245;
	wire [15-1:0] node15248;
	wire [15-1:0] node15251;
	wire [15-1:0] node15252;
	wire [15-1:0] node15253;
	wire [15-1:0] node15254;
	wire [15-1:0] node15255;
	wire [15-1:0] node15258;
	wire [15-1:0] node15261;
	wire [15-1:0] node15262;
	wire [15-1:0] node15265;
	wire [15-1:0] node15268;
	wire [15-1:0] node15269;
	wire [15-1:0] node15271;
	wire [15-1:0] node15274;
	wire [15-1:0] node15275;
	wire [15-1:0] node15278;
	wire [15-1:0] node15281;
	wire [15-1:0] node15282;
	wire [15-1:0] node15283;
	wire [15-1:0] node15284;
	wire [15-1:0] node15287;
	wire [15-1:0] node15290;
	wire [15-1:0] node15291;
	wire [15-1:0] node15294;
	wire [15-1:0] node15297;
	wire [15-1:0] node15298;
	wire [15-1:0] node15301;
	wire [15-1:0] node15302;
	wire [15-1:0] node15305;
	wire [15-1:0] node15308;
	wire [15-1:0] node15309;
	wire [15-1:0] node15310;
	wire [15-1:0] node15311;
	wire [15-1:0] node15312;
	wire [15-1:0] node15313;
	wire [15-1:0] node15314;
	wire [15-1:0] node15317;
	wire [15-1:0] node15320;
	wire [15-1:0] node15321;
	wire [15-1:0] node15324;
	wire [15-1:0] node15327;
	wire [15-1:0] node15328;
	wire [15-1:0] node15329;
	wire [15-1:0] node15332;
	wire [15-1:0] node15335;
	wire [15-1:0] node15336;
	wire [15-1:0] node15339;
	wire [15-1:0] node15342;
	wire [15-1:0] node15343;
	wire [15-1:0] node15344;
	wire [15-1:0] node15345;
	wire [15-1:0] node15348;
	wire [15-1:0] node15351;
	wire [15-1:0] node15352;
	wire [15-1:0] node15355;
	wire [15-1:0] node15358;
	wire [15-1:0] node15359;
	wire [15-1:0] node15360;
	wire [15-1:0] node15363;
	wire [15-1:0] node15366;
	wire [15-1:0] node15367;
	wire [15-1:0] node15370;
	wire [15-1:0] node15373;
	wire [15-1:0] node15374;
	wire [15-1:0] node15375;
	wire [15-1:0] node15376;
	wire [15-1:0] node15378;
	wire [15-1:0] node15381;
	wire [15-1:0] node15382;
	wire [15-1:0] node15385;
	wire [15-1:0] node15388;
	wire [15-1:0] node15389;
	wire [15-1:0] node15391;
	wire [15-1:0] node15394;
	wire [15-1:0] node15395;
	wire [15-1:0] node15398;
	wire [15-1:0] node15401;
	wire [15-1:0] node15402;
	wire [15-1:0] node15403;
	wire [15-1:0] node15404;
	wire [15-1:0] node15407;
	wire [15-1:0] node15410;
	wire [15-1:0] node15411;
	wire [15-1:0] node15414;
	wire [15-1:0] node15417;
	wire [15-1:0] node15418;
	wire [15-1:0] node15419;
	wire [15-1:0] node15422;
	wire [15-1:0] node15425;
	wire [15-1:0] node15426;
	wire [15-1:0] node15429;
	wire [15-1:0] node15432;
	wire [15-1:0] node15433;
	wire [15-1:0] node15434;
	wire [15-1:0] node15435;
	wire [15-1:0] node15436;
	wire [15-1:0] node15437;
	wire [15-1:0] node15440;
	wire [15-1:0] node15443;
	wire [15-1:0] node15444;
	wire [15-1:0] node15447;
	wire [15-1:0] node15450;
	wire [15-1:0] node15451;
	wire [15-1:0] node15452;
	wire [15-1:0] node15455;
	wire [15-1:0] node15458;
	wire [15-1:0] node15459;
	wire [15-1:0] node15462;
	wire [15-1:0] node15465;
	wire [15-1:0] node15466;
	wire [15-1:0] node15467;
	wire [15-1:0] node15468;
	wire [15-1:0] node15471;
	wire [15-1:0] node15474;
	wire [15-1:0] node15475;
	wire [15-1:0] node15478;
	wire [15-1:0] node15481;
	wire [15-1:0] node15482;
	wire [15-1:0] node15483;
	wire [15-1:0] node15486;
	wire [15-1:0] node15489;
	wire [15-1:0] node15490;
	wire [15-1:0] node15493;
	wire [15-1:0] node15496;
	wire [15-1:0] node15497;
	wire [15-1:0] node15498;
	wire [15-1:0] node15499;
	wire [15-1:0] node15500;
	wire [15-1:0] node15503;
	wire [15-1:0] node15506;
	wire [15-1:0] node15507;
	wire [15-1:0] node15510;
	wire [15-1:0] node15513;
	wire [15-1:0] node15514;
	wire [15-1:0] node15515;
	wire [15-1:0] node15518;
	wire [15-1:0] node15521;
	wire [15-1:0] node15522;
	wire [15-1:0] node15525;
	wire [15-1:0] node15528;
	wire [15-1:0] node15529;
	wire [15-1:0] node15530;
	wire [15-1:0] node15532;
	wire [15-1:0] node15535;
	wire [15-1:0] node15536;
	wire [15-1:0] node15539;
	wire [15-1:0] node15542;
	wire [15-1:0] node15543;
	wire [15-1:0] node15544;
	wire [15-1:0] node15547;
	wire [15-1:0] node15550;
	wire [15-1:0] node15552;

	assign outp = (inp[6]) ? node7754 : node1;
		assign node1 = (inp[5]) ? node3887 : node2;
			assign node2 = (inp[9]) ? node1952 : node3;
				assign node3 = (inp[0]) ? node995 : node4;
					assign node4 = (inp[1]) ? node500 : node5;
						assign node5 = (inp[8]) ? node251 : node6;
							assign node6 = (inp[3]) ? node130 : node7;
								assign node7 = (inp[7]) ? node69 : node8;
									assign node8 = (inp[4]) ? node40 : node9;
										assign node9 = (inp[2]) ? node25 : node10;
											assign node10 = (inp[11]) ? node18 : node11;
												assign node11 = (inp[13]) ? node15 : node12;
													assign node12 = (inp[14]) ? 15'b001111111111111 : 15'b011111111111111;
													assign node15 = (inp[10]) ? 15'b000111111111111 : 15'b001111111111111;
												assign node18 = (inp[10]) ? node22 : node19;
													assign node19 = (inp[14]) ? 15'b000111111111111 : 15'b001111111111111;
													assign node22 = (inp[12]) ? 15'b000001111111111 : 15'b000111111111111;
											assign node25 = (inp[12]) ? node33 : node26;
												assign node26 = (inp[14]) ? node30 : node27;
													assign node27 = (inp[13]) ? 15'b000111111111111 : 15'b001111111111111;
													assign node30 = (inp[10]) ? 15'b000011111111111 : 15'b000111111111111;
												assign node33 = (inp[10]) ? node37 : node34;
													assign node34 = (inp[13]) ? 15'b000011111111111 : 15'b000111111111111;
													assign node37 = (inp[13]) ? 15'b000001111111111 : 15'b000011111111111;
										assign node40 = (inp[12]) ? node56 : node41;
											assign node41 = (inp[14]) ? node49 : node42;
												assign node42 = (inp[2]) ? node46 : node43;
													assign node43 = (inp[10]) ? 15'b000111111111111 : 15'b011111111111111;
													assign node46 = (inp[13]) ? 15'b000011111111111 : 15'b000111111111111;
												assign node49 = (inp[11]) ? node53 : node50;
													assign node50 = (inp[10]) ? 15'b000011111111111 : 15'b000111111111111;
													assign node53 = (inp[13]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node56 = (inp[10]) ? node64 : node57;
												assign node57 = (inp[11]) ? node61 : node58;
													assign node58 = (inp[2]) ? 15'b000011111111111 : 15'b000111111111111;
													assign node61 = (inp[13]) ? 15'b000000111111111 : 15'b000011111111111;
												assign node64 = (inp[2]) ? 15'b000001111111111 : node65;
													assign node65 = (inp[13]) ? 15'b000001111111111 : 15'b000011111111111;
									assign node69 = (inp[12]) ? node99 : node70;
										assign node70 = (inp[2]) ? node84 : node71;
											assign node71 = (inp[10]) ? node77 : node72;
												assign node72 = (inp[13]) ? node74 : 15'b001111111111111;
													assign node74 = (inp[11]) ? 15'b000011111111111 : 15'b000111111111111;
												assign node77 = (inp[11]) ? node81 : node78;
													assign node78 = (inp[4]) ? 15'b000011111111111 : 15'b000111111111111;
													assign node81 = (inp[14]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node84 = (inp[11]) ? node92 : node85;
												assign node85 = (inp[14]) ? node89 : node86;
													assign node86 = (inp[13]) ? 15'b000011111111111 : 15'b000111111111111;
													assign node89 = (inp[13]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node92 = (inp[4]) ? node96 : node93;
													assign node93 = (inp[10]) ? 15'b000001111111111 : 15'b000001111111111;
													assign node96 = (inp[10]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node99 = (inp[10]) ? node115 : node100;
											assign node100 = (inp[14]) ? node108 : node101;
												assign node101 = (inp[4]) ? node105 : node102;
													assign node102 = (inp[13]) ? 15'b000011111111111 : 15'b000111111111111;
													assign node105 = (inp[13]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node108 = (inp[13]) ? node112 : node109;
													assign node109 = (inp[2]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node112 = (inp[4]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node115 = (inp[11]) ? node123 : node116;
												assign node116 = (inp[14]) ? node120 : node117;
													assign node117 = (inp[13]) ? 15'b000001111111111 : 15'b000001111111111;
													assign node120 = (inp[4]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node123 = (inp[13]) ? node127 : node124;
													assign node124 = (inp[2]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node127 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
								assign node130 = (inp[2]) ? node192 : node131;
									assign node131 = (inp[14]) ? node163 : node132;
										assign node132 = (inp[10]) ? node148 : node133;
											assign node133 = (inp[12]) ? node141 : node134;
												assign node134 = (inp[7]) ? node138 : node135;
													assign node135 = (inp[13]) ? 15'b000111111111111 : 15'b001111111111111;
													assign node138 = (inp[4]) ? 15'b000011111111111 : 15'b000111111111111;
												assign node141 = (inp[11]) ? node145 : node142;
													assign node142 = (inp[13]) ? 15'b000011111111111 : 15'b000011111111111;
													assign node145 = (inp[7]) ? 15'b000001111111111 : 15'b000001111111111;
											assign node148 = (inp[7]) ? node156 : node149;
												assign node149 = (inp[11]) ? node153 : node150;
													assign node150 = (inp[4]) ? 15'b000011111111111 : 15'b000011111111111;
													assign node153 = (inp[12]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node156 = (inp[4]) ? node160 : node157;
													assign node157 = (inp[13]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node160 = (inp[13]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node163 = (inp[7]) ? node179 : node164;
											assign node164 = (inp[10]) ? node172 : node165;
												assign node165 = (inp[4]) ? node169 : node166;
													assign node166 = (inp[13]) ? 15'b000011111111111 : 15'b000111111111111;
													assign node169 = (inp[13]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node172 = (inp[12]) ? node176 : node173;
													assign node173 = (inp[13]) ? 15'b000000111111111 : 15'b000011111111111;
													assign node176 = (inp[4]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node179 = (inp[10]) ? node187 : node180;
												assign node180 = (inp[12]) ? node184 : node181;
													assign node181 = (inp[13]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node184 = (inp[11]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node187 = (inp[11]) ? 15'b000000011111111 : node188;
													assign node188 = (inp[12]) ? 15'b000000111111111 : 15'b000001111111111;
									assign node192 = (inp[14]) ? node224 : node193;
										assign node193 = (inp[13]) ? node209 : node194;
											assign node194 = (inp[7]) ? node202 : node195;
												assign node195 = (inp[12]) ? node199 : node196;
													assign node196 = (inp[4]) ? 15'b000011111111111 : 15'b000111111111111;
													assign node199 = (inp[10]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node202 = (inp[12]) ? node206 : node203;
													assign node203 = (inp[4]) ? 15'b000000111111111 : 15'b000011111111111;
													assign node206 = (inp[10]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node209 = (inp[10]) ? node217 : node210;
												assign node210 = (inp[12]) ? node214 : node211;
													assign node211 = (inp[11]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node214 = (inp[11]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node217 = (inp[4]) ? node221 : node218;
													assign node218 = (inp[7]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node221 = (inp[7]) ? 15'b000000011111111 : 15'b000000011111111;
										assign node224 = (inp[7]) ? node240 : node225;
											assign node225 = (inp[4]) ? node233 : node226;
												assign node226 = (inp[10]) ? node230 : node227;
													assign node227 = (inp[11]) ? 15'b000001111111111 : 15'b000001111111111;
													assign node230 = (inp[12]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node233 = (inp[12]) ? node237 : node234;
													assign node234 = (inp[11]) ? 15'b000000111111111 : 15'b000000111111111;
													assign node237 = (inp[10]) ? 15'b000000011111111 : 15'b000001111111111;
											assign node240 = (inp[4]) ? node246 : node241;
												assign node241 = (inp[10]) ? node243 : 15'b000000111111111;
													assign node243 = (inp[12]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node246 = (inp[10]) ? node248 : 15'b000000011111111;
													assign node248 = (inp[12]) ? 15'b000000000111111 : 15'b000000011111111;
							assign node251 = (inp[13]) ? node377 : node252;
								assign node252 = (inp[4]) ? node314 : node253;
									assign node253 = (inp[2]) ? node285 : node254;
										assign node254 = (inp[10]) ? node270 : node255;
											assign node255 = (inp[12]) ? node263 : node256;
												assign node256 = (inp[14]) ? node260 : node257;
													assign node257 = (inp[3]) ? 15'b000111111111111 : 15'b001111111111111;
													assign node260 = (inp[3]) ? 15'b000011111111111 : 15'b000111111111111;
												assign node263 = (inp[11]) ? node267 : node264;
													assign node264 = (inp[7]) ? 15'b000011111111111 : 15'b000111111111111;
													assign node267 = (inp[3]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node270 = (inp[12]) ? node278 : node271;
												assign node271 = (inp[11]) ? node275 : node272;
													assign node272 = (inp[3]) ? 15'b000011111111111 : 15'b000111111111111;
													assign node275 = (inp[14]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node278 = (inp[11]) ? node282 : node279;
													assign node279 = (inp[3]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node282 = (inp[3]) ? 15'b000000111111111 : 15'b000000111111111;
										assign node285 = (inp[10]) ? node299 : node286;
											assign node286 = (inp[14]) ? node294 : node287;
												assign node287 = (inp[3]) ? node291 : node288;
													assign node288 = (inp[12]) ? 15'b000011111111111 : 15'b000111111111111;
													assign node291 = (inp[12]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node294 = (inp[12]) ? 15'b000000011111111 : node295;
													assign node295 = (inp[7]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node299 = (inp[11]) ? node307 : node300;
												assign node300 = (inp[7]) ? node304 : node301;
													assign node301 = (inp[14]) ? 15'b000001111111111 : 15'b000001111111111;
													assign node304 = (inp[3]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node307 = (inp[14]) ? node311 : node308;
													assign node308 = (inp[7]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node311 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node314 = (inp[3]) ? node346 : node315;
										assign node315 = (inp[11]) ? node331 : node316;
											assign node316 = (inp[2]) ? node324 : node317;
												assign node317 = (inp[7]) ? node321 : node318;
													assign node318 = (inp[14]) ? 15'b000011111111111 : 15'b000111111111111;
													assign node321 = (inp[10]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node324 = (inp[14]) ? node328 : node325;
													assign node325 = (inp[10]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node328 = (inp[12]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node331 = (inp[12]) ? node339 : node332;
												assign node332 = (inp[7]) ? node336 : node333;
													assign node333 = (inp[2]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node336 = (inp[2]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node339 = (inp[2]) ? node343 : node340;
													assign node340 = (inp[7]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node343 = (inp[14]) ? 15'b000000111111111 : 15'b000000111111111;
										assign node346 = (inp[14]) ? node362 : node347;
											assign node347 = (inp[7]) ? node355 : node348;
												assign node348 = (inp[11]) ? node352 : node349;
													assign node349 = (inp[2]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node352 = (inp[10]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node355 = (inp[11]) ? node359 : node356;
													assign node356 = (inp[2]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node359 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node362 = (inp[10]) ? node370 : node363;
												assign node363 = (inp[7]) ? node367 : node364;
													assign node364 = (inp[11]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node367 = (inp[12]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node370 = (inp[11]) ? node374 : node371;
													assign node371 = (inp[7]) ? 15'b000000001111111 : 15'b000000111111111;
													assign node374 = (inp[12]) ? 15'b000000001111111 : 15'b000000001111111;
								assign node377 = (inp[7]) ? node441 : node378;
									assign node378 = (inp[3]) ? node410 : node379;
										assign node379 = (inp[4]) ? node395 : node380;
											assign node380 = (inp[10]) ? node388 : node381;
												assign node381 = (inp[2]) ? node385 : node382;
													assign node382 = (inp[11]) ? 15'b000011111111111 : 15'b000011111111111;
													assign node385 = (inp[14]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node388 = (inp[11]) ? node392 : node389;
													assign node389 = (inp[12]) ? 15'b000001111111111 : 15'b000111111111111;
													assign node392 = (inp[2]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node395 = (inp[11]) ? node403 : node396;
												assign node396 = (inp[14]) ? node400 : node397;
													assign node397 = (inp[12]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node400 = (inp[12]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node403 = (inp[10]) ? node407 : node404;
													assign node404 = (inp[12]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node407 = (inp[12]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node410 = (inp[2]) ? node426 : node411;
											assign node411 = (inp[10]) ? node419 : node412;
												assign node412 = (inp[14]) ? node416 : node413;
													assign node413 = (inp[4]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node416 = (inp[11]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node419 = (inp[12]) ? node423 : node420;
													assign node420 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node423 = (inp[4]) ? 15'b000000011111111 : 15'b000000011111111;
											assign node426 = (inp[11]) ? node434 : node427;
												assign node427 = (inp[4]) ? node431 : node428;
													assign node428 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node431 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node434 = (inp[10]) ? node438 : node435;
													assign node435 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node438 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node441 = (inp[2]) ? node471 : node442;
										assign node442 = (inp[4]) ? node456 : node443;
											assign node443 = (inp[14]) ? node449 : node444;
												assign node444 = (inp[12]) ? 15'b000001111111111 : node445;
													assign node445 = (inp[11]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node449 = (inp[10]) ? node453 : node450;
													assign node450 = (inp[3]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node453 = (inp[12]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node456 = (inp[11]) ? node464 : node457;
												assign node457 = (inp[12]) ? node461 : node458;
													assign node458 = (inp[3]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node461 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node464 = (inp[3]) ? node468 : node465;
													assign node465 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node468 = (inp[10]) ? 15'b000000000111111 : 15'b000000011111111;
										assign node471 = (inp[11]) ? node487 : node472;
											assign node472 = (inp[4]) ? node480 : node473;
												assign node473 = (inp[12]) ? node477 : node474;
													assign node474 = (inp[10]) ? 15'b000001111111111 : 15'b000000111111111;
													assign node477 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node480 = (inp[3]) ? node484 : node481;
													assign node481 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node484 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node487 = (inp[4]) ? node495 : node488;
												assign node488 = (inp[10]) ? node492 : node489;
													assign node489 = (inp[3]) ? 15'b000000011111111 : 15'b000000011111111;
													assign node492 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node495 = (inp[12]) ? node497 : 15'b000000011111111;
													assign node497 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
						assign node500 = (inp[4]) ? node742 : node501;
							assign node501 = (inp[2]) ? node621 : node502;
								assign node502 = (inp[10]) ? node560 : node503;
									assign node503 = (inp[13]) ? node535 : node504;
										assign node504 = (inp[14]) ? node520 : node505;
											assign node505 = (inp[3]) ? node513 : node506;
												assign node506 = (inp[7]) ? node510 : node507;
													assign node507 = (inp[8]) ? 15'b000111111111111 : 15'b001111111111111;
													assign node510 = (inp[8]) ? 15'b000011111111111 : 15'b000111111111111;
												assign node513 = (inp[12]) ? node517 : node514;
													assign node514 = (inp[7]) ? 15'b000011111111111 : 15'b000111111111111;
													assign node517 = (inp[8]) ? 15'b000011111111111 : 15'b000011111111111;
											assign node520 = (inp[3]) ? node528 : node521;
												assign node521 = (inp[11]) ? node525 : node522;
													assign node522 = (inp[12]) ? 15'b000011111111111 : 15'b000111111111111;
													assign node525 = (inp[12]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node528 = (inp[12]) ? node532 : node529;
													assign node529 = (inp[11]) ? 15'b000001111111111 : 15'b000111111111111;
													assign node532 = (inp[8]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node535 = (inp[11]) ? node551 : node536;
											assign node536 = (inp[8]) ? node544 : node537;
												assign node537 = (inp[3]) ? node541 : node538;
													assign node538 = (inp[14]) ? 15'b000111111111111 : 15'b000111111111111;
													assign node541 = (inp[12]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node544 = (inp[7]) ? node548 : node545;
													assign node545 = (inp[14]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node548 = (inp[14]) ? 15'b000000011111111 : 15'b000001111111111;
											assign node551 = (inp[8]) ? 15'b000000111111111 : node552;
												assign node552 = (inp[7]) ? node556 : node553;
													assign node553 = (inp[12]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node556 = (inp[3]) ? 15'b000000111111111 : 15'b000001111111111;
									assign node560 = (inp[11]) ? node592 : node561;
										assign node561 = (inp[3]) ? node577 : node562;
											assign node562 = (inp[12]) ? node570 : node563;
												assign node563 = (inp[7]) ? node567 : node564;
													assign node564 = (inp[8]) ? 15'b000011111111111 : 15'b000111111111111;
													assign node567 = (inp[8]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node570 = (inp[13]) ? node574 : node571;
													assign node571 = (inp[14]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node574 = (inp[8]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node577 = (inp[8]) ? node585 : node578;
												assign node578 = (inp[12]) ? node582 : node579;
													assign node579 = (inp[13]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node582 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node585 = (inp[13]) ? node589 : node586;
													assign node586 = (inp[12]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node589 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node592 = (inp[7]) ? node606 : node593;
											assign node593 = (inp[3]) ? node601 : node594;
												assign node594 = (inp[12]) ? node598 : node595;
													assign node595 = (inp[8]) ? 15'b000000111111111 : 15'b000011111111111;
													assign node598 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node601 = (inp[14]) ? 15'b000000111111111 : node602;
													assign node602 = (inp[12]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node606 = (inp[13]) ? node614 : node607;
												assign node607 = (inp[12]) ? node611 : node608;
													assign node608 = (inp[3]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node611 = (inp[14]) ? 15'b000000001111111 : 15'b000000111111111;
												assign node614 = (inp[3]) ? node618 : node615;
													assign node615 = (inp[8]) ? 15'b000000011111111 : 15'b000000011111111;
													assign node618 = (inp[8]) ? 15'b000000000111111 : 15'b000000011111111;
								assign node621 = (inp[7]) ? node683 : node622;
									assign node622 = (inp[12]) ? node652 : node623;
										assign node623 = (inp[10]) ? node639 : node624;
											assign node624 = (inp[11]) ? node632 : node625;
												assign node625 = (inp[14]) ? node629 : node626;
													assign node626 = (inp[3]) ? 15'b000011111111111 : 15'b000111111111111;
													assign node629 = (inp[3]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node632 = (inp[14]) ? node636 : node633;
													assign node633 = (inp[8]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node636 = (inp[3]) ? 15'b000000011111111 : 15'b000001111111111;
											assign node639 = (inp[13]) ? node645 : node640;
												assign node640 = (inp[11]) ? 15'b000000111111111 : node641;
													assign node641 = (inp[8]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node645 = (inp[8]) ? node649 : node646;
													assign node646 = (inp[3]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node649 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node652 = (inp[13]) ? node668 : node653;
											assign node653 = (inp[8]) ? node661 : node654;
												assign node654 = (inp[11]) ? node658 : node655;
													assign node655 = (inp[3]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node658 = (inp[10]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node661 = (inp[11]) ? node665 : node662;
													assign node662 = (inp[3]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node665 = (inp[10]) ? 15'b000000001111111 : 15'b000000111111111;
											assign node668 = (inp[14]) ? node676 : node669;
												assign node669 = (inp[8]) ? node673 : node670;
													assign node670 = (inp[3]) ? 15'b000000111111111 : 15'b000011111111111;
													assign node673 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node676 = (inp[3]) ? node680 : node677;
													assign node677 = (inp[11]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node680 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node683 = (inp[10]) ? node713 : node684;
										assign node684 = (inp[12]) ? node698 : node685;
											assign node685 = (inp[3]) ? node691 : node686;
												assign node686 = (inp[8]) ? 15'b000001111111111 : node687;
													assign node687 = (inp[11]) ? 15'b000000111111111 : 15'b000011111111111;
												assign node691 = (inp[11]) ? node695 : node692;
													assign node692 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node695 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node698 = (inp[8]) ? node706 : node699;
												assign node699 = (inp[13]) ? node703 : node700;
													assign node700 = (inp[11]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node703 = (inp[11]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node706 = (inp[14]) ? node710 : node707;
													assign node707 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node710 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node713 = (inp[12]) ? node729 : node714;
											assign node714 = (inp[3]) ? node722 : node715;
												assign node715 = (inp[13]) ? node719 : node716;
													assign node716 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node719 = (inp[11]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node722 = (inp[8]) ? node726 : node723;
													assign node723 = (inp[13]) ? 15'b000000011111111 : 15'b000000011111111;
													assign node726 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node729 = (inp[3]) ? node735 : node730;
												assign node730 = (inp[8]) ? node732 : 15'b000000011111111;
													assign node732 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node735 = (inp[13]) ? node739 : node736;
													assign node736 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node739 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
							assign node742 = (inp[11]) ? node868 : node743;
								assign node743 = (inp[14]) ? node805 : node744;
									assign node744 = (inp[13]) ? node776 : node745;
										assign node745 = (inp[2]) ? node761 : node746;
											assign node746 = (inp[8]) ? node754 : node747;
												assign node747 = (inp[7]) ? node751 : node748;
													assign node748 = (inp[10]) ? 15'b000011111111111 : 15'b000111111111111;
													assign node751 = (inp[10]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node754 = (inp[10]) ? node758 : node755;
													assign node755 = (inp[12]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node758 = (inp[7]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node761 = (inp[7]) ? node769 : node762;
												assign node762 = (inp[8]) ? node766 : node763;
													assign node763 = (inp[3]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node766 = (inp[10]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node769 = (inp[3]) ? node773 : node770;
													assign node770 = (inp[10]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node773 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node776 = (inp[10]) ? node792 : node777;
											assign node777 = (inp[12]) ? node785 : node778;
												assign node778 = (inp[3]) ? node782 : node779;
													assign node779 = (inp[7]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node782 = (inp[2]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node785 = (inp[8]) ? node789 : node786;
													assign node786 = (inp[7]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node789 = (inp[7]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node792 = (inp[3]) ? node798 : node793;
												assign node793 = (inp[7]) ? 15'b000000111111111 : node794;
													assign node794 = (inp[12]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node798 = (inp[7]) ? node802 : node799;
													assign node799 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node802 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node805 = (inp[7]) ? node837 : node806;
										assign node806 = (inp[10]) ? node822 : node807;
											assign node807 = (inp[13]) ? node815 : node808;
												assign node808 = (inp[12]) ? node812 : node809;
													assign node809 = (inp[8]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node812 = (inp[8]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node815 = (inp[2]) ? node819 : node816;
													assign node816 = (inp[12]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node819 = (inp[12]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node822 = (inp[8]) ? node830 : node823;
												assign node823 = (inp[12]) ? node827 : node824;
													assign node824 = (inp[2]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node827 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node830 = (inp[12]) ? node834 : node831;
													assign node831 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node834 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node837 = (inp[3]) ? node853 : node838;
											assign node838 = (inp[2]) ? node846 : node839;
												assign node839 = (inp[10]) ? node843 : node840;
													assign node840 = (inp[8]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node843 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node846 = (inp[8]) ? node850 : node847;
													assign node847 = (inp[13]) ? 15'b000000011111111 : 15'b000000011111111;
													assign node850 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node853 = (inp[8]) ? node861 : node854;
												assign node854 = (inp[13]) ? node858 : node855;
													assign node855 = (inp[12]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node858 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node861 = (inp[13]) ? node865 : node862;
													assign node862 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node865 = (inp[12]) ? 15'b000000000111111 : 15'b000000001111111;
								assign node868 = (inp[12]) ? node932 : node869;
									assign node869 = (inp[3]) ? node901 : node870;
										assign node870 = (inp[10]) ? node886 : node871;
											assign node871 = (inp[8]) ? node879 : node872;
												assign node872 = (inp[7]) ? node876 : node873;
													assign node873 = (inp[2]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node876 = (inp[13]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node879 = (inp[14]) ? node883 : node880;
													assign node880 = (inp[7]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node883 = (inp[7]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node886 = (inp[2]) ? node894 : node887;
												assign node887 = (inp[7]) ? node891 : node888;
													assign node888 = (inp[13]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node891 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node894 = (inp[14]) ? node898 : node895;
													assign node895 = (inp[13]) ? 15'b000000011111111 : 15'b000000011111111;
													assign node898 = (inp[7]) ? 15'b000000001111111 : 15'b000000001111111;
										assign node901 = (inp[8]) ? node917 : node902;
											assign node902 = (inp[14]) ? node910 : node903;
												assign node903 = (inp[13]) ? node907 : node904;
													assign node904 = (inp[10]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node907 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node910 = (inp[2]) ? node914 : node911;
													assign node911 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node914 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node917 = (inp[10]) ? node925 : node918;
												assign node918 = (inp[7]) ? node922 : node919;
													assign node919 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node922 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node925 = (inp[14]) ? node929 : node926;
													assign node926 = (inp[13]) ? 15'b000000001111111 : 15'b000000001111111;
													assign node929 = (inp[7]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node932 = (inp[13]) ? node964 : node933;
										assign node933 = (inp[2]) ? node949 : node934;
											assign node934 = (inp[14]) ? node942 : node935;
												assign node935 = (inp[10]) ? node939 : node936;
													assign node936 = (inp[7]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node939 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node942 = (inp[3]) ? node946 : node943;
													assign node943 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node946 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node949 = (inp[8]) ? node957 : node950;
												assign node950 = (inp[3]) ? node954 : node951;
													assign node951 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node954 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node957 = (inp[10]) ? node961 : node958;
													assign node958 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node961 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node964 = (inp[8]) ? node980 : node965;
											assign node965 = (inp[14]) ? node973 : node966;
												assign node966 = (inp[3]) ? node970 : node967;
													assign node967 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node970 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node973 = (inp[10]) ? node977 : node974;
													assign node974 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node977 = (inp[7]) ? 15'b000000000111111 : 15'b000000000111111;
											assign node980 = (inp[3]) ? node988 : node981;
												assign node981 = (inp[7]) ? node985 : node982;
													assign node982 = (inp[2]) ? 15'b000000000111111 : 15'b000000011111111;
													assign node985 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node988 = (inp[7]) ? node992 : node989;
													assign node989 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node992 = (inp[2]) ? 15'b000000000011111 : 15'b000000000111111;
					assign node995 = (inp[4]) ? node1469 : node996;
						assign node996 = (inp[3]) ? node1238 : node997;
							assign node997 = (inp[2]) ? node1119 : node998;
								assign node998 = (inp[13]) ? node1058 : node999;
									assign node999 = (inp[1]) ? node1029 : node1000;
										assign node1000 = (inp[14]) ? node1014 : node1001;
											assign node1001 = (inp[8]) ? node1009 : node1002;
												assign node1002 = (inp[7]) ? node1006 : node1003;
													assign node1003 = (inp[11]) ? 15'b000111111111111 : 15'b001111111111111;
													assign node1006 = (inp[10]) ? 15'b000011111111111 : 15'b000111111111111;
												assign node1009 = (inp[11]) ? 15'b000011111111111 : node1010;
													assign node1010 = (inp[10]) ? 15'b000011111111111 : 15'b000111111111111;
											assign node1014 = (inp[10]) ? node1022 : node1015;
												assign node1015 = (inp[7]) ? node1019 : node1016;
													assign node1016 = (inp[8]) ? 15'b000011111111111 : 15'b000111111111111;
													assign node1019 = (inp[12]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node1022 = (inp[12]) ? node1026 : node1023;
													assign node1023 = (inp[8]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node1026 = (inp[11]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node1029 = (inp[12]) ? node1043 : node1030;
											assign node1030 = (inp[11]) ? node1036 : node1031;
												assign node1031 = (inp[7]) ? node1033 : 15'b000111111111111;
													assign node1033 = (inp[10]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node1036 = (inp[10]) ? node1040 : node1037;
													assign node1037 = (inp[14]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node1040 = (inp[8]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node1043 = (inp[7]) ? node1051 : node1044;
												assign node1044 = (inp[14]) ? node1048 : node1045;
													assign node1045 = (inp[11]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node1048 = (inp[11]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node1051 = (inp[8]) ? node1055 : node1052;
													assign node1052 = (inp[10]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node1055 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node1058 = (inp[7]) ? node1090 : node1059;
										assign node1059 = (inp[11]) ? node1075 : node1060;
											assign node1060 = (inp[8]) ? node1068 : node1061;
												assign node1061 = (inp[10]) ? node1065 : node1062;
													assign node1062 = (inp[1]) ? 15'b000011111111111 : 15'b000111111111111;
													assign node1065 = (inp[1]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node1068 = (inp[10]) ? node1072 : node1069;
													assign node1069 = (inp[14]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node1072 = (inp[1]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node1075 = (inp[1]) ? node1083 : node1076;
												assign node1076 = (inp[14]) ? node1080 : node1077;
													assign node1077 = (inp[8]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node1080 = (inp[10]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node1083 = (inp[12]) ? node1087 : node1084;
													assign node1084 = (inp[10]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node1087 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node1090 = (inp[10]) ? node1106 : node1091;
											assign node1091 = (inp[14]) ? node1099 : node1092;
												assign node1092 = (inp[12]) ? node1096 : node1093;
													assign node1093 = (inp[8]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node1096 = (inp[1]) ? 15'b000000111111111 : 15'b000011111111111;
												assign node1099 = (inp[11]) ? node1103 : node1100;
													assign node1100 = (inp[8]) ? 15'b000000011111111 : 15'b000001111111111;
													assign node1103 = (inp[12]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node1106 = (inp[8]) ? node1114 : node1107;
												assign node1107 = (inp[1]) ? node1111 : node1108;
													assign node1108 = (inp[11]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node1111 = (inp[12]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node1114 = (inp[1]) ? 15'b000000011111111 : node1115;
													assign node1115 = (inp[11]) ? 15'b000000011111111 : 15'b000000111111111;
								assign node1119 = (inp[12]) ? node1183 : node1120;
									assign node1120 = (inp[7]) ? node1152 : node1121;
										assign node1121 = (inp[10]) ? node1137 : node1122;
											assign node1122 = (inp[11]) ? node1130 : node1123;
												assign node1123 = (inp[8]) ? node1127 : node1124;
													assign node1124 = (inp[13]) ? 15'b000011111111111 : 15'b000111111111111;
													assign node1127 = (inp[1]) ? 15'b000000111111111 : 15'b000011111111111;
												assign node1130 = (inp[13]) ? node1134 : node1131;
													assign node1131 = (inp[8]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node1134 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node1137 = (inp[13]) ? node1145 : node1138;
												assign node1138 = (inp[1]) ? node1142 : node1139;
													assign node1139 = (inp[8]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node1142 = (inp[11]) ? 15'b000000011111111 : 15'b000001111111111;
												assign node1145 = (inp[1]) ? node1149 : node1146;
													assign node1146 = (inp[8]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node1149 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node1152 = (inp[1]) ? node1168 : node1153;
											assign node1153 = (inp[13]) ? node1161 : node1154;
												assign node1154 = (inp[14]) ? node1158 : node1155;
													assign node1155 = (inp[11]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node1158 = (inp[8]) ? 15'b000000111111111 : 15'b000000111111111;
												assign node1161 = (inp[11]) ? node1165 : node1162;
													assign node1162 = (inp[10]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node1165 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node1168 = (inp[14]) ? node1176 : node1169;
												assign node1169 = (inp[13]) ? node1173 : node1170;
													assign node1170 = (inp[8]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node1173 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node1176 = (inp[10]) ? node1180 : node1177;
													assign node1177 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node1180 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node1183 = (inp[14]) ? node1209 : node1184;
										assign node1184 = (inp[11]) ? node1196 : node1185;
											assign node1185 = (inp[13]) ? node1189 : node1186;
												assign node1186 = (inp[10]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node1189 = (inp[1]) ? node1193 : node1190;
													assign node1190 = (inp[7]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node1193 = (inp[7]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node1196 = (inp[8]) ? node1202 : node1197;
												assign node1197 = (inp[1]) ? node1199 : 15'b000000111111111;
													assign node1199 = (inp[7]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node1202 = (inp[10]) ? node1206 : node1203;
													assign node1203 = (inp[7]) ? 15'b000000011111111 : 15'b000000011111111;
													assign node1206 = (inp[13]) ? 15'b000000001111111 : 15'b000000001111111;
										assign node1209 = (inp[10]) ? node1225 : node1210;
											assign node1210 = (inp[1]) ? node1218 : node1211;
												assign node1211 = (inp[13]) ? node1215 : node1212;
													assign node1212 = (inp[8]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node1215 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node1218 = (inp[8]) ? node1222 : node1219;
													assign node1219 = (inp[11]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node1222 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node1225 = (inp[11]) ? node1231 : node1226;
												assign node1226 = (inp[13]) ? node1228 : 15'b000000011111111;
													assign node1228 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node1231 = (inp[7]) ? node1235 : node1232;
													assign node1232 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node1235 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
							assign node1238 = (inp[8]) ? node1356 : node1239;
								assign node1239 = (inp[12]) ? node1299 : node1240;
									assign node1240 = (inp[14]) ? node1272 : node1241;
										assign node1241 = (inp[10]) ? node1257 : node1242;
											assign node1242 = (inp[2]) ? node1250 : node1243;
												assign node1243 = (inp[7]) ? node1247 : node1244;
													assign node1244 = (inp[11]) ? 15'b000011111111111 : 15'b000111111111111;
													assign node1247 = (inp[13]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node1250 = (inp[13]) ? node1254 : node1251;
													assign node1251 = (inp[7]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node1254 = (inp[1]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node1257 = (inp[1]) ? node1265 : node1258;
												assign node1258 = (inp[11]) ? node1262 : node1259;
													assign node1259 = (inp[2]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node1262 = (inp[7]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node1265 = (inp[13]) ? node1269 : node1266;
													assign node1266 = (inp[2]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node1269 = (inp[7]) ? 15'b000000001111111 : 15'b000000111111111;
										assign node1272 = (inp[13]) ? node1286 : node1273;
											assign node1273 = (inp[1]) ? node1279 : node1274;
												assign node1274 = (inp[11]) ? 15'b000001111111111 : node1275;
													assign node1275 = (inp[10]) ? 15'b000011111111111 : 15'b000001111111111;
												assign node1279 = (inp[7]) ? node1283 : node1280;
													assign node1280 = (inp[2]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node1283 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node1286 = (inp[7]) ? node1294 : node1287;
												assign node1287 = (inp[10]) ? node1291 : node1288;
													assign node1288 = (inp[1]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node1291 = (inp[1]) ? 15'b000000001111111 : 15'b000000111111111;
												assign node1294 = (inp[11]) ? 15'b000000011111111 : node1295;
													assign node1295 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node1299 = (inp[1]) ? node1327 : node1300;
										assign node1300 = (inp[10]) ? node1314 : node1301;
											assign node1301 = (inp[11]) ? node1309 : node1302;
												assign node1302 = (inp[13]) ? node1306 : node1303;
													assign node1303 = (inp[2]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node1306 = (inp[7]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node1309 = (inp[2]) ? 15'b000000011111111 : node1310;
													assign node1310 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node1314 = (inp[11]) ? node1320 : node1315;
												assign node1315 = (inp[13]) ? node1317 : 15'b000001111111111;
													assign node1317 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node1320 = (inp[14]) ? node1324 : node1321;
													assign node1321 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node1324 = (inp[7]) ? 15'b000000000111111 : 15'b000000011111111;
										assign node1327 = (inp[13]) ? node1343 : node1328;
											assign node1328 = (inp[11]) ? node1336 : node1329;
												assign node1329 = (inp[10]) ? node1333 : node1330;
													assign node1330 = (inp[7]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node1333 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node1336 = (inp[10]) ? node1340 : node1337;
													assign node1337 = (inp[7]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node1340 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node1343 = (inp[10]) ? node1349 : node1344;
												assign node1344 = (inp[11]) ? node1346 : 15'b000000011111111;
													assign node1346 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node1349 = (inp[11]) ? node1353 : node1350;
													assign node1350 = (inp[2]) ? 15'b000000001111111 : 15'b000000001111111;
													assign node1353 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
								assign node1356 = (inp[7]) ? node1416 : node1357;
									assign node1357 = (inp[13]) ? node1385 : node1358;
										assign node1358 = (inp[10]) ? node1370 : node1359;
											assign node1359 = (inp[2]) ? node1365 : node1360;
												assign node1360 = (inp[12]) ? 15'b000001111111111 : node1361;
													assign node1361 = (inp[1]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node1365 = (inp[11]) ? node1367 : 15'b000001111111111;
													assign node1367 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node1370 = (inp[14]) ? node1378 : node1371;
												assign node1371 = (inp[1]) ? node1375 : node1372;
													assign node1372 = (inp[2]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node1375 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node1378 = (inp[2]) ? node1382 : node1379;
													assign node1379 = (inp[12]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node1382 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node1385 = (inp[11]) ? node1401 : node1386;
											assign node1386 = (inp[2]) ? node1394 : node1387;
												assign node1387 = (inp[1]) ? node1391 : node1388;
													assign node1388 = (inp[12]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node1391 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node1394 = (inp[10]) ? node1398 : node1395;
													assign node1395 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node1398 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node1401 = (inp[1]) ? node1409 : node1402;
												assign node1402 = (inp[12]) ? node1406 : node1403;
													assign node1403 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node1406 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node1409 = (inp[2]) ? node1413 : node1410;
													assign node1410 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node1413 = (inp[14]) ? 15'b000000000111111 : 15'b000000000111111;
									assign node1416 = (inp[13]) ? node1440 : node1417;
										assign node1417 = (inp[10]) ? node1425 : node1418;
											assign node1418 = (inp[12]) ? 15'b000000011111111 : node1419;
												assign node1419 = (inp[11]) ? node1421 : 15'b000000111111111;
													assign node1421 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node1425 = (inp[11]) ? node1433 : node1426;
												assign node1426 = (inp[2]) ? node1430 : node1427;
													assign node1427 = (inp[12]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node1430 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node1433 = (inp[1]) ? node1437 : node1434;
													assign node1434 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node1437 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node1440 = (inp[1]) ? node1456 : node1441;
											assign node1441 = (inp[2]) ? node1449 : node1442;
												assign node1442 = (inp[11]) ? node1446 : node1443;
													assign node1443 = (inp[14]) ? 15'b000000011111111 : 15'b000000011111111;
													assign node1446 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node1449 = (inp[12]) ? node1453 : node1450;
													assign node1450 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node1453 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node1456 = (inp[11]) ? node1464 : node1457;
												assign node1457 = (inp[14]) ? node1461 : node1458;
													assign node1458 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node1461 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node1464 = (inp[14]) ? node1466 : 15'b000000000111111;
													assign node1466 = (inp[2]) ? 15'b000000000011111 : 15'b000000000111111;
						assign node1469 = (inp[13]) ? node1705 : node1470;
							assign node1470 = (inp[8]) ? node1588 : node1471;
								assign node1471 = (inp[2]) ? node1529 : node1472;
									assign node1472 = (inp[3]) ? node1504 : node1473;
										assign node1473 = (inp[14]) ? node1489 : node1474;
											assign node1474 = (inp[7]) ? node1482 : node1475;
												assign node1475 = (inp[10]) ? node1479 : node1476;
													assign node1476 = (inp[11]) ? 15'b000011111111111 : 15'b000111111111111;
													assign node1479 = (inp[12]) ? 15'b000000111111111 : 15'b000011111111111;
												assign node1482 = (inp[1]) ? node1486 : node1483;
													assign node1483 = (inp[11]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node1486 = (inp[10]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node1489 = (inp[12]) ? node1497 : node1490;
												assign node1490 = (inp[10]) ? node1494 : node1491;
													assign node1491 = (inp[11]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node1494 = (inp[1]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node1497 = (inp[11]) ? node1501 : node1498;
													assign node1498 = (inp[7]) ? 15'b000000011111111 : 15'b000001111111111;
													assign node1501 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node1504 = (inp[10]) ? node1520 : node1505;
											assign node1505 = (inp[1]) ? node1513 : node1506;
												assign node1506 = (inp[14]) ? node1510 : node1507;
													assign node1507 = (inp[7]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node1510 = (inp[7]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node1513 = (inp[7]) ? node1517 : node1514;
													assign node1514 = (inp[11]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node1517 = (inp[11]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node1520 = (inp[11]) ? node1522 : 15'b000000111111111;
												assign node1522 = (inp[14]) ? node1526 : node1523;
													assign node1523 = (inp[12]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node1526 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node1529 = (inp[12]) ? node1561 : node1530;
										assign node1530 = (inp[1]) ? node1546 : node1531;
											assign node1531 = (inp[10]) ? node1539 : node1532;
												assign node1532 = (inp[3]) ? node1536 : node1533;
													assign node1533 = (inp[7]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node1536 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node1539 = (inp[11]) ? node1543 : node1540;
													assign node1540 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node1543 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node1546 = (inp[3]) ? node1554 : node1547;
												assign node1547 = (inp[10]) ? node1551 : node1548;
													assign node1548 = (inp[7]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node1551 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node1554 = (inp[7]) ? node1558 : node1555;
													assign node1555 = (inp[11]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node1558 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node1561 = (inp[11]) ? node1575 : node1562;
											assign node1562 = (inp[7]) ? node1568 : node1563;
												assign node1563 = (inp[1]) ? 15'b000000111111111 : node1564;
													assign node1564 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node1568 = (inp[14]) ? node1572 : node1569;
													assign node1569 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node1572 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node1575 = (inp[10]) ? node1581 : node1576;
												assign node1576 = (inp[7]) ? 15'b000000011111111 : node1577;
													assign node1577 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node1581 = (inp[14]) ? node1585 : node1582;
													assign node1582 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node1585 = (inp[1]) ? 15'b000000000011111 : 15'b000000001111111;
								assign node1588 = (inp[14]) ? node1648 : node1589;
									assign node1589 = (inp[7]) ? node1621 : node1590;
										assign node1590 = (inp[12]) ? node1606 : node1591;
											assign node1591 = (inp[2]) ? node1599 : node1592;
												assign node1592 = (inp[3]) ? node1596 : node1593;
													assign node1593 = (inp[11]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node1596 = (inp[10]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node1599 = (inp[10]) ? node1603 : node1600;
													assign node1600 = (inp[3]) ? 15'b000000111111111 : 15'b000000111111111;
													assign node1603 = (inp[11]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node1606 = (inp[10]) ? node1614 : node1607;
												assign node1607 = (inp[1]) ? node1611 : node1608;
													assign node1608 = (inp[2]) ? 15'b000000111111111 : 15'b000000111111111;
													assign node1611 = (inp[11]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node1614 = (inp[2]) ? node1618 : node1615;
													assign node1615 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node1618 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node1621 = (inp[2]) ? node1635 : node1622;
											assign node1622 = (inp[1]) ? node1628 : node1623;
												assign node1623 = (inp[11]) ? node1625 : 15'b000001111111111;
													assign node1625 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node1628 = (inp[10]) ? node1632 : node1629;
													assign node1629 = (inp[11]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node1632 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node1635 = (inp[10]) ? node1643 : node1636;
												assign node1636 = (inp[11]) ? node1640 : node1637;
													assign node1637 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node1640 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node1643 = (inp[3]) ? node1645 : 15'b000000001111111;
													assign node1645 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node1648 = (inp[10]) ? node1678 : node1649;
										assign node1649 = (inp[1]) ? node1665 : node1650;
											assign node1650 = (inp[12]) ? node1658 : node1651;
												assign node1651 = (inp[2]) ? node1655 : node1652;
													assign node1652 = (inp[7]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node1655 = (inp[7]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node1658 = (inp[3]) ? node1662 : node1659;
													assign node1659 = (inp[2]) ? 15'b000000011111111 : 15'b000000011111111;
													assign node1662 = (inp[7]) ? 15'b000000000111111 : 15'b000000011111111;
											assign node1665 = (inp[3]) ? node1671 : node1666;
												assign node1666 = (inp[7]) ? node1668 : 15'b000000111111111;
													assign node1668 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node1671 = (inp[2]) ? node1675 : node1672;
													assign node1672 = (inp[11]) ? 15'b000000000111111 : 15'b000000011111111;
													assign node1675 = (inp[7]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node1678 = (inp[11]) ? node1694 : node1679;
											assign node1679 = (inp[2]) ? node1687 : node1680;
												assign node1680 = (inp[7]) ? node1684 : node1681;
													assign node1681 = (inp[12]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node1684 = (inp[3]) ? 15'b000000001111111 : 15'b000000001111111;
												assign node1687 = (inp[12]) ? node1691 : node1688;
													assign node1688 = (inp[7]) ? 15'b000000001111111 : 15'b000000001111111;
													assign node1691 = (inp[3]) ? 15'b000000000011111 : 15'b000000001111111;
											assign node1694 = (inp[12]) ? node1700 : node1695;
												assign node1695 = (inp[3]) ? node1697 : 15'b000000001111111;
													assign node1697 = (inp[2]) ? 15'b000000000111111 : 15'b000000000111111;
												assign node1700 = (inp[2]) ? node1702 : 15'b000000000111111;
													assign node1702 = (inp[1]) ? 15'b000000000011111 : 15'b000000000111111;
							assign node1705 = (inp[3]) ? node1833 : node1706;
								assign node1706 = (inp[2]) ? node1770 : node1707;
									assign node1707 = (inp[8]) ? node1739 : node1708;
										assign node1708 = (inp[11]) ? node1724 : node1709;
											assign node1709 = (inp[7]) ? node1717 : node1710;
												assign node1710 = (inp[10]) ? node1714 : node1711;
													assign node1711 = (inp[14]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node1714 = (inp[12]) ? 15'b000000011111111 : 15'b000001111111111;
												assign node1717 = (inp[12]) ? node1721 : node1718;
													assign node1718 = (inp[10]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node1721 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node1724 = (inp[1]) ? node1732 : node1725;
												assign node1725 = (inp[12]) ? node1729 : node1726;
													assign node1726 = (inp[7]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node1729 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node1732 = (inp[7]) ? node1736 : node1733;
													assign node1733 = (inp[10]) ? 15'b000000011111111 : 15'b000000011111111;
													assign node1736 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node1739 = (inp[14]) ? node1755 : node1740;
											assign node1740 = (inp[11]) ? node1748 : node1741;
												assign node1741 = (inp[10]) ? node1745 : node1742;
													assign node1742 = (inp[12]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node1745 = (inp[12]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node1748 = (inp[1]) ? node1752 : node1749;
													assign node1749 = (inp[10]) ? 15'b000000011111111 : 15'b000001111111111;
													assign node1752 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node1755 = (inp[1]) ? node1763 : node1756;
												assign node1756 = (inp[7]) ? node1760 : node1757;
													assign node1757 = (inp[10]) ? 15'b000000001111111 : 15'b000000111111111;
													assign node1760 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node1763 = (inp[11]) ? node1767 : node1764;
													assign node1764 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node1767 = (inp[7]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node1770 = (inp[1]) ? node1802 : node1771;
										assign node1771 = (inp[11]) ? node1787 : node1772;
											assign node1772 = (inp[7]) ? node1780 : node1773;
												assign node1773 = (inp[10]) ? node1777 : node1774;
													assign node1774 = (inp[12]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node1777 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node1780 = (inp[14]) ? node1784 : node1781;
													assign node1781 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node1784 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node1787 = (inp[7]) ? node1795 : node1788;
												assign node1788 = (inp[14]) ? node1792 : node1789;
													assign node1789 = (inp[12]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node1792 = (inp[12]) ? 15'b000000001111111 : 15'b000000001111111;
												assign node1795 = (inp[14]) ? node1799 : node1796;
													assign node1796 = (inp[10]) ? 15'b000000001111111 : 15'b000000001111111;
													assign node1799 = (inp[12]) ? 15'b000000000111111 : 15'b000000000111111;
										assign node1802 = (inp[8]) ? node1818 : node1803;
											assign node1803 = (inp[7]) ? node1811 : node1804;
												assign node1804 = (inp[14]) ? node1808 : node1805;
													assign node1805 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node1808 = (inp[10]) ? 15'b000000001111111 : 15'b000000001111111;
												assign node1811 = (inp[10]) ? node1815 : node1812;
													assign node1812 = (inp[12]) ? 15'b000000001111111 : 15'b000000111111111;
													assign node1815 = (inp[12]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node1818 = (inp[11]) ? node1826 : node1819;
												assign node1819 = (inp[10]) ? node1823 : node1820;
													assign node1820 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node1823 = (inp[12]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node1826 = (inp[10]) ? node1830 : node1827;
													assign node1827 = (inp[12]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node1830 = (inp[7]) ? 15'b000000000011111 : 15'b000000000011111;
								assign node1833 = (inp[10]) ? node1895 : node1834;
									assign node1834 = (inp[11]) ? node1866 : node1835;
										assign node1835 = (inp[1]) ? node1851 : node1836;
											assign node1836 = (inp[2]) ? node1844 : node1837;
												assign node1837 = (inp[8]) ? node1841 : node1838;
													assign node1838 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node1841 = (inp[12]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node1844 = (inp[14]) ? node1848 : node1845;
													assign node1845 = (inp[12]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node1848 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node1851 = (inp[12]) ? node1859 : node1852;
												assign node1852 = (inp[2]) ? node1856 : node1853;
													assign node1853 = (inp[7]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node1856 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node1859 = (inp[14]) ? node1863 : node1860;
													assign node1860 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node1863 = (inp[2]) ? 15'b000000000111111 : 15'b000000000111111;
										assign node1866 = (inp[8]) ? node1880 : node1867;
											assign node1867 = (inp[7]) ? node1875 : node1868;
												assign node1868 = (inp[2]) ? node1872 : node1869;
													assign node1869 = (inp[12]) ? 15'b000000011111111 : 15'b000001111111111;
													assign node1872 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node1875 = (inp[1]) ? node1877 : 15'b000000001111111;
													assign node1877 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node1880 = (inp[2]) ? node1888 : node1881;
												assign node1881 = (inp[12]) ? node1885 : node1882;
													assign node1882 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node1885 = (inp[7]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node1888 = (inp[1]) ? node1892 : node1889;
													assign node1889 = (inp[7]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node1892 = (inp[14]) ? 15'b000000000001111 : 15'b000000000111111;
									assign node1895 = (inp[7]) ? node1923 : node1896;
										assign node1896 = (inp[1]) ? node1912 : node1897;
											assign node1897 = (inp[11]) ? node1905 : node1898;
												assign node1898 = (inp[12]) ? node1902 : node1899;
													assign node1899 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node1902 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node1905 = (inp[8]) ? node1909 : node1906;
													assign node1906 = (inp[12]) ? 15'b000000001111111 : 15'b000000001111111;
													assign node1909 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node1912 = (inp[2]) ? node1918 : node1913;
												assign node1913 = (inp[12]) ? 15'b000000000111111 : node1914;
													assign node1914 = (inp[14]) ? 15'b000000000111111 : 15'b000000011111111;
												assign node1918 = (inp[14]) ? node1920 : 15'b000000000111111;
													assign node1920 = (inp[8]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node1923 = (inp[12]) ? node1937 : node1924;
											assign node1924 = (inp[1]) ? node1930 : node1925;
												assign node1925 = (inp[8]) ? node1927 : 15'b000000001111111;
													assign node1927 = (inp[11]) ? 15'b000000000011111 : 15'b000000001111111;
												assign node1930 = (inp[2]) ? node1934 : node1931;
													assign node1931 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node1934 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node1937 = (inp[14]) ? node1945 : node1938;
												assign node1938 = (inp[8]) ? node1942 : node1939;
													assign node1939 = (inp[1]) ? 15'b000000001111111 : 15'b000000001111111;
													assign node1942 = (inp[2]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node1945 = (inp[11]) ? node1949 : node1946;
													assign node1946 = (inp[8]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node1949 = (inp[8]) ? 15'b000000000001111 : 15'b000000000011111;
				assign node1952 = (inp[13]) ? node2922 : node1953;
					assign node1953 = (inp[11]) ? node2441 : node1954;
						assign node1954 = (inp[14]) ? node2196 : node1955;
							assign node1955 = (inp[7]) ? node2075 : node1956;
								assign node1956 = (inp[12]) ? node2018 : node1957;
									assign node1957 = (inp[3]) ? node1989 : node1958;
										assign node1958 = (inp[1]) ? node1974 : node1959;
											assign node1959 = (inp[4]) ? node1967 : node1960;
												assign node1960 = (inp[2]) ? node1964 : node1961;
													assign node1961 = (inp[10]) ? 15'b000111111111111 : 15'b001111111111111;
													assign node1964 = (inp[10]) ? 15'b000011111111111 : 15'b000111111111111;
												assign node1967 = (inp[0]) ? node1971 : node1968;
													assign node1968 = (inp[8]) ? 15'b000011111111111 : 15'b000111111111111;
													assign node1971 = (inp[8]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node1974 = (inp[0]) ? node1982 : node1975;
												assign node1975 = (inp[4]) ? node1979 : node1976;
													assign node1976 = (inp[10]) ? 15'b000001111111111 : 15'b000111111111111;
													assign node1979 = (inp[2]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node1982 = (inp[8]) ? node1986 : node1983;
													assign node1983 = (inp[10]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node1986 = (inp[2]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node1989 = (inp[10]) ? node2005 : node1990;
											assign node1990 = (inp[8]) ? node1998 : node1991;
												assign node1991 = (inp[2]) ? node1995 : node1992;
													assign node1992 = (inp[1]) ? 15'b000011111111111 : 15'b000111111111111;
													assign node1995 = (inp[1]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node1998 = (inp[0]) ? node2002 : node1999;
													assign node1999 = (inp[4]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node2002 = (inp[1]) ? 15'b000000011111111 : 15'b000001111111111;
											assign node2005 = (inp[1]) ? node2013 : node2006;
												assign node2006 = (inp[0]) ? node2010 : node2007;
													assign node2007 = (inp[2]) ? 15'b000001111111111 : 15'b000001111111111;
													assign node2010 = (inp[2]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node2013 = (inp[0]) ? 15'b000000111111111 : node2014;
													assign node2014 = (inp[8]) ? 15'b000000111111111 : 15'b000001111111111;
									assign node2018 = (inp[2]) ? node2050 : node2019;
										assign node2019 = (inp[8]) ? node2035 : node2020;
											assign node2020 = (inp[10]) ? node2028 : node2021;
												assign node2021 = (inp[3]) ? node2025 : node2022;
													assign node2022 = (inp[1]) ? 15'b000011111111111 : 15'b000111111111111;
													assign node2025 = (inp[4]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node2028 = (inp[0]) ? node2032 : node2029;
													assign node2029 = (inp[1]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node2032 = (inp[3]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node2035 = (inp[10]) ? node2043 : node2036;
												assign node2036 = (inp[3]) ? node2040 : node2037;
													assign node2037 = (inp[4]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node2040 = (inp[0]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node2043 = (inp[1]) ? node2047 : node2044;
													assign node2044 = (inp[0]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node2047 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node2050 = (inp[4]) ? node2066 : node2051;
											assign node2051 = (inp[1]) ? node2059 : node2052;
												assign node2052 = (inp[10]) ? node2056 : node2053;
													assign node2053 = (inp[0]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node2056 = (inp[0]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node2059 = (inp[10]) ? node2063 : node2060;
													assign node2060 = (inp[3]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node2063 = (inp[0]) ? 15'b000000011111111 : 15'b000000011111111;
											assign node2066 = (inp[1]) ? 15'b000000011111111 : node2067;
												assign node2067 = (inp[8]) ? node2071 : node2068;
													assign node2068 = (inp[0]) ? 15'b000000111111111 : 15'b000000111111111;
													assign node2071 = (inp[3]) ? 15'b000000001111111 : 15'b000000111111111;
								assign node2075 = (inp[10]) ? node2137 : node2076;
									assign node2076 = (inp[3]) ? node2108 : node2077;
										assign node2077 = (inp[0]) ? node2093 : node2078;
											assign node2078 = (inp[4]) ? node2086 : node2079;
												assign node2079 = (inp[8]) ? node2083 : node2080;
													assign node2080 = (inp[1]) ? 15'b000011111111111 : 15'b000111111111111;
													assign node2083 = (inp[12]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node2086 = (inp[2]) ? node2090 : node2087;
													assign node2087 = (inp[8]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node2090 = (inp[12]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node2093 = (inp[1]) ? node2101 : node2094;
												assign node2094 = (inp[12]) ? node2098 : node2095;
													assign node2095 = (inp[2]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node2098 = (inp[2]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node2101 = (inp[8]) ? node2105 : node2102;
													assign node2102 = (inp[4]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node2105 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node2108 = (inp[2]) ? node2122 : node2109;
											assign node2109 = (inp[1]) ? node2117 : node2110;
												assign node2110 = (inp[8]) ? node2114 : node2111;
													assign node2111 = (inp[4]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node2114 = (inp[0]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node2117 = (inp[12]) ? 15'b000000011111111 : node2118;
													assign node2118 = (inp[4]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node2122 = (inp[8]) ? node2130 : node2123;
												assign node2123 = (inp[0]) ? node2127 : node2124;
													assign node2124 = (inp[1]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node2127 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node2130 = (inp[4]) ? node2134 : node2131;
													assign node2131 = (inp[12]) ? 15'b000000011111111 : 15'b000001111111111;
													assign node2134 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node2137 = (inp[1]) ? node2167 : node2138;
										assign node2138 = (inp[2]) ? node2154 : node2139;
											assign node2139 = (inp[0]) ? node2147 : node2140;
												assign node2140 = (inp[8]) ? node2144 : node2141;
													assign node2141 = (inp[3]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node2144 = (inp[3]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node2147 = (inp[8]) ? node2151 : node2148;
													assign node2148 = (inp[4]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node2151 = (inp[12]) ? 15'b000000001111111 : 15'b000000111111111;
											assign node2154 = (inp[4]) ? node2160 : node2155;
												assign node2155 = (inp[0]) ? 15'b000000011111111 : node2156;
													assign node2156 = (inp[12]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node2160 = (inp[8]) ? node2164 : node2161;
													assign node2161 = (inp[12]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node2164 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node2167 = (inp[3]) ? node2181 : node2168;
											assign node2168 = (inp[12]) ? node2174 : node2169;
												assign node2169 = (inp[0]) ? 15'b000000111111111 : node2170;
													assign node2170 = (inp[2]) ? 15'b000000011111111 : 15'b000001111111111;
												assign node2174 = (inp[2]) ? node2178 : node2175;
													assign node2175 = (inp[8]) ? 15'b000000011111111 : 15'b000000011111111;
													assign node2178 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node2181 = (inp[12]) ? node2189 : node2182;
												assign node2182 = (inp[8]) ? node2186 : node2183;
													assign node2183 = (inp[2]) ? 15'b000000011111111 : 15'b000000011111111;
													assign node2186 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node2189 = (inp[0]) ? node2193 : node2190;
													assign node2190 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node2193 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
							assign node2196 = (inp[1]) ? node2318 : node2197;
								assign node2197 = (inp[12]) ? node2257 : node2198;
									assign node2198 = (inp[3]) ? node2226 : node2199;
										assign node2199 = (inp[7]) ? node2213 : node2200;
											assign node2200 = (inp[10]) ? node2208 : node2201;
												assign node2201 = (inp[4]) ? node2205 : node2202;
													assign node2202 = (inp[0]) ? 15'b000011111111111 : 15'b000111111111111;
													assign node2205 = (inp[2]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node2208 = (inp[0]) ? 15'b000001111111111 : node2209;
													assign node2209 = (inp[4]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node2213 = (inp[10]) ? node2221 : node2214;
												assign node2214 = (inp[0]) ? node2218 : node2215;
													assign node2215 = (inp[8]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node2218 = (inp[2]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node2221 = (inp[2]) ? 15'b000000111111111 : node2222;
													assign node2222 = (inp[8]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node2226 = (inp[2]) ? node2242 : node2227;
											assign node2227 = (inp[4]) ? node2235 : node2228;
												assign node2228 = (inp[7]) ? node2232 : node2229;
													assign node2229 = (inp[8]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node2232 = (inp[0]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node2235 = (inp[10]) ? node2239 : node2236;
													assign node2236 = (inp[7]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node2239 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node2242 = (inp[10]) ? node2250 : node2243;
												assign node2243 = (inp[4]) ? node2247 : node2244;
													assign node2244 = (inp[8]) ? 15'b000000111111111 : 15'b000000111111111;
													assign node2247 = (inp[7]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node2250 = (inp[7]) ? node2254 : node2251;
													assign node2251 = (inp[0]) ? 15'b000000011111111 : 15'b000001111111111;
													assign node2254 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node2257 = (inp[8]) ? node2287 : node2258;
										assign node2258 = (inp[4]) ? node2272 : node2259;
											assign node2259 = (inp[7]) ? node2265 : node2260;
												assign node2260 = (inp[2]) ? 15'b000001111111111 : node2261;
													assign node2261 = (inp[0]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node2265 = (inp[2]) ? node2269 : node2266;
													assign node2266 = (inp[0]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node2269 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node2272 = (inp[0]) ? node2280 : node2273;
												assign node2273 = (inp[2]) ? node2277 : node2274;
													assign node2274 = (inp[3]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node2277 = (inp[7]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node2280 = (inp[10]) ? node2284 : node2281;
													assign node2281 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node2284 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node2287 = (inp[4]) ? node2303 : node2288;
											assign node2288 = (inp[7]) ? node2296 : node2289;
												assign node2289 = (inp[2]) ? node2293 : node2290;
													assign node2290 = (inp[3]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node2293 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node2296 = (inp[10]) ? node2300 : node2297;
													assign node2297 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node2300 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node2303 = (inp[2]) ? node2311 : node2304;
												assign node2304 = (inp[3]) ? node2308 : node2305;
													assign node2305 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node2308 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node2311 = (inp[0]) ? node2315 : node2312;
													assign node2312 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node2315 = (inp[3]) ? 15'b000000000011111 : 15'b000000001111111;
								assign node2318 = (inp[0]) ? node2380 : node2319;
									assign node2319 = (inp[12]) ? node2351 : node2320;
										assign node2320 = (inp[8]) ? node2336 : node2321;
											assign node2321 = (inp[10]) ? node2329 : node2322;
												assign node2322 = (inp[7]) ? node2326 : node2323;
													assign node2323 = (inp[4]) ? 15'b000011111111111 : 15'b000011111111111;
													assign node2326 = (inp[3]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node2329 = (inp[3]) ? node2333 : node2330;
													assign node2330 = (inp[7]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node2333 = (inp[7]) ? 15'b000000111111111 : 15'b000000111111111;
											assign node2336 = (inp[2]) ? node2344 : node2337;
												assign node2337 = (inp[3]) ? node2341 : node2338;
													assign node2338 = (inp[10]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node2341 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node2344 = (inp[10]) ? node2348 : node2345;
													assign node2345 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node2348 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node2351 = (inp[3]) ? node2367 : node2352;
											assign node2352 = (inp[8]) ? node2360 : node2353;
												assign node2353 = (inp[2]) ? node2357 : node2354;
													assign node2354 = (inp[4]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node2357 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node2360 = (inp[4]) ? node2364 : node2361;
													assign node2361 = (inp[10]) ? 15'b000000011111111 : 15'b000000011111111;
													assign node2364 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node2367 = (inp[4]) ? node2375 : node2368;
												assign node2368 = (inp[8]) ? node2372 : node2369;
													assign node2369 = (inp[2]) ? 15'b000000011111111 : 15'b000000011111111;
													assign node2372 = (inp[2]) ? 15'b000000001111111 : 15'b000000001111111;
												assign node2375 = (inp[7]) ? 15'b000000000111111 : node2376;
													assign node2376 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node2380 = (inp[2]) ? node2410 : node2381;
										assign node2381 = (inp[10]) ? node2397 : node2382;
											assign node2382 = (inp[7]) ? node2390 : node2383;
												assign node2383 = (inp[3]) ? node2387 : node2384;
													assign node2384 = (inp[8]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node2387 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node2390 = (inp[8]) ? node2394 : node2391;
													assign node2391 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node2394 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node2397 = (inp[12]) ? node2405 : node2398;
												assign node2398 = (inp[4]) ? node2402 : node2399;
													assign node2399 = (inp[3]) ? 15'b000000011111111 : 15'b000000011111111;
													assign node2402 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node2405 = (inp[4]) ? node2407 : 15'b000000001111111;
													assign node2407 = (inp[3]) ? 15'b000000000111111 : 15'b000000000111111;
										assign node2410 = (inp[8]) ? node2426 : node2411;
											assign node2411 = (inp[3]) ? node2419 : node2412;
												assign node2412 = (inp[4]) ? node2416 : node2413;
													assign node2413 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node2416 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node2419 = (inp[7]) ? node2423 : node2420;
													assign node2420 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node2423 = (inp[12]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node2426 = (inp[12]) ? node2434 : node2427;
												assign node2427 = (inp[7]) ? node2431 : node2428;
													assign node2428 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node2431 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node2434 = (inp[10]) ? node2438 : node2435;
													assign node2435 = (inp[7]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node2438 = (inp[3]) ? 15'b000000000011111 : 15'b000000000111111;
						assign node2441 = (inp[3]) ? node2681 : node2442;
							assign node2442 = (inp[4]) ? node2560 : node2443;
								assign node2443 = (inp[8]) ? node2501 : node2444;
									assign node2444 = (inp[0]) ? node2476 : node2445;
										assign node2445 = (inp[7]) ? node2461 : node2446;
											assign node2446 = (inp[1]) ? node2454 : node2447;
												assign node2447 = (inp[2]) ? node2451 : node2448;
													assign node2448 = (inp[14]) ? 15'b000011111111111 : 15'b000111111111111;
													assign node2451 = (inp[12]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node2454 = (inp[10]) ? node2458 : node2455;
													assign node2455 = (inp[12]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node2458 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node2461 = (inp[10]) ? node2469 : node2462;
												assign node2462 = (inp[2]) ? node2466 : node2463;
													assign node2463 = (inp[14]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node2466 = (inp[12]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node2469 = (inp[2]) ? node2473 : node2470;
													assign node2470 = (inp[12]) ? 15'b000000011111111 : 15'b000001111111111;
													assign node2473 = (inp[14]) ? 15'b000000011111111 : 15'b000000011111111;
										assign node2476 = (inp[2]) ? node2490 : node2477;
											assign node2477 = (inp[7]) ? node2485 : node2478;
												assign node2478 = (inp[10]) ? node2482 : node2479;
													assign node2479 = (inp[12]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node2482 = (inp[12]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node2485 = (inp[12]) ? 15'b000000111111111 : node2486;
													assign node2486 = (inp[1]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node2490 = (inp[12]) ? node2498 : node2491;
												assign node2491 = (inp[1]) ? node2495 : node2492;
													assign node2492 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node2495 = (inp[14]) ? 15'b000000001111111 : 15'b000000111111111;
												assign node2498 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node2501 = (inp[0]) ? node2531 : node2502;
										assign node2502 = (inp[1]) ? node2518 : node2503;
											assign node2503 = (inp[7]) ? node2511 : node2504;
												assign node2504 = (inp[10]) ? node2508 : node2505;
													assign node2505 = (inp[2]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node2508 = (inp[12]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node2511 = (inp[14]) ? node2515 : node2512;
													assign node2512 = (inp[12]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node2515 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node2518 = (inp[10]) ? node2524 : node2519;
												assign node2519 = (inp[2]) ? 15'b000000011111111 : node2520;
													assign node2520 = (inp[12]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node2524 = (inp[7]) ? node2528 : node2525;
													assign node2525 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node2528 = (inp[12]) ? 15'b000000000111111 : 15'b000000011111111;
										assign node2531 = (inp[12]) ? node2545 : node2532;
											assign node2532 = (inp[14]) ? node2540 : node2533;
												assign node2533 = (inp[10]) ? node2537 : node2534;
													assign node2534 = (inp[7]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node2537 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node2540 = (inp[10]) ? 15'b000000001111111 : node2541;
													assign node2541 = (inp[1]) ? 15'b000000001111111 : 15'b000000111111111;
											assign node2545 = (inp[10]) ? node2553 : node2546;
												assign node2546 = (inp[14]) ? node2550 : node2547;
													assign node2547 = (inp[7]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node2550 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node2553 = (inp[1]) ? node2557 : node2554;
													assign node2554 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node2557 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
								assign node2560 = (inp[7]) ? node2622 : node2561;
									assign node2561 = (inp[0]) ? node2591 : node2562;
										assign node2562 = (inp[14]) ? node2576 : node2563;
											assign node2563 = (inp[8]) ? node2571 : node2564;
												assign node2564 = (inp[10]) ? node2568 : node2565;
													assign node2565 = (inp[12]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node2568 = (inp[12]) ? 15'b000000011111111 : 15'b000001111111111;
												assign node2571 = (inp[2]) ? 15'b000000111111111 : node2572;
													assign node2572 = (inp[1]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node2576 = (inp[12]) ? node2584 : node2577;
												assign node2577 = (inp[2]) ? node2581 : node2578;
													assign node2578 = (inp[10]) ? 15'b000001111111111 : 15'b000001111111111;
													assign node2581 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node2584 = (inp[10]) ? node2588 : node2585;
													assign node2585 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node2588 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node2591 = (inp[2]) ? node2607 : node2592;
											assign node2592 = (inp[10]) ? node2600 : node2593;
												assign node2593 = (inp[1]) ? node2597 : node2594;
													assign node2594 = (inp[12]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node2597 = (inp[12]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node2600 = (inp[14]) ? node2604 : node2601;
													assign node2601 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node2604 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node2607 = (inp[14]) ? node2615 : node2608;
												assign node2608 = (inp[10]) ? node2612 : node2609;
													assign node2609 = (inp[12]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node2612 = (inp[12]) ? 15'b000000001111111 : 15'b000000001111111;
												assign node2615 = (inp[8]) ? node2619 : node2616;
													assign node2616 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node2619 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node2622 = (inp[2]) ? node2652 : node2623;
										assign node2623 = (inp[12]) ? node2639 : node2624;
											assign node2624 = (inp[10]) ? node2632 : node2625;
												assign node2625 = (inp[8]) ? node2629 : node2626;
													assign node2626 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node2629 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node2632 = (inp[1]) ? node2636 : node2633;
													assign node2633 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node2636 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node2639 = (inp[0]) ? node2647 : node2640;
												assign node2640 = (inp[8]) ? node2644 : node2641;
													assign node2641 = (inp[1]) ? 15'b000000011111111 : 15'b000000011111111;
													assign node2644 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node2647 = (inp[14]) ? 15'b000000000111111 : node2648;
													assign node2648 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node2652 = (inp[14]) ? node2666 : node2653;
											assign node2653 = (inp[1]) ? node2659 : node2654;
												assign node2654 = (inp[0]) ? 15'b000000011111111 : node2655;
													assign node2655 = (inp[8]) ? 15'b000000011111111 : 15'b000000011111111;
												assign node2659 = (inp[0]) ? node2663 : node2660;
													assign node2660 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node2663 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node2666 = (inp[10]) ? node2674 : node2667;
												assign node2667 = (inp[12]) ? node2671 : node2668;
													assign node2668 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node2671 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node2674 = (inp[12]) ? node2678 : node2675;
													assign node2675 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node2678 = (inp[8]) ? 15'b000000000011111 : 15'b000000000111111;
							assign node2681 = (inp[8]) ? node2803 : node2682;
								assign node2682 = (inp[2]) ? node2742 : node2683;
									assign node2683 = (inp[4]) ? node2713 : node2684;
										assign node2684 = (inp[14]) ? node2700 : node2685;
											assign node2685 = (inp[12]) ? node2693 : node2686;
												assign node2686 = (inp[7]) ? node2690 : node2687;
													assign node2687 = (inp[1]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node2690 = (inp[10]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node2693 = (inp[1]) ? node2697 : node2694;
													assign node2694 = (inp[10]) ? 15'b000000111111111 : 15'b000011111111111;
													assign node2697 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node2700 = (inp[7]) ? node2708 : node2701;
												assign node2701 = (inp[10]) ? node2705 : node2702;
													assign node2702 = (inp[12]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node2705 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node2708 = (inp[1]) ? node2710 : 15'b000000111111111;
													assign node2710 = (inp[12]) ? 15'b000000000111111 : 15'b000000011111111;
										assign node2713 = (inp[12]) ? node2729 : node2714;
											assign node2714 = (inp[7]) ? node2722 : node2715;
												assign node2715 = (inp[1]) ? node2719 : node2716;
													assign node2716 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node2719 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node2722 = (inp[1]) ? node2726 : node2723;
													assign node2723 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node2726 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node2729 = (inp[1]) ? node2735 : node2730;
												assign node2730 = (inp[14]) ? node2732 : 15'b000000011111111;
													assign node2732 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node2735 = (inp[0]) ? node2739 : node2736;
													assign node2736 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node2739 = (inp[10]) ? 15'b000000001111111 : 15'b000000000111111;
									assign node2742 = (inp[14]) ? node2774 : node2743;
										assign node2743 = (inp[12]) ? node2759 : node2744;
											assign node2744 = (inp[0]) ? node2752 : node2745;
												assign node2745 = (inp[10]) ? node2749 : node2746;
													assign node2746 = (inp[1]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node2749 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node2752 = (inp[10]) ? node2756 : node2753;
													assign node2753 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node2756 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node2759 = (inp[10]) ? node2767 : node2760;
												assign node2760 = (inp[4]) ? node2764 : node2761;
													assign node2761 = (inp[7]) ? 15'b000000011111111 : 15'b000000011111111;
													assign node2764 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node2767 = (inp[4]) ? node2771 : node2768;
													assign node2768 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node2771 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node2774 = (inp[1]) ? node2790 : node2775;
											assign node2775 = (inp[7]) ? node2783 : node2776;
												assign node2776 = (inp[0]) ? node2780 : node2777;
													assign node2777 = (inp[12]) ? 15'b000000011111111 : 15'b000001111111111;
													assign node2780 = (inp[12]) ? 15'b000000000111111 : 15'b000000011111111;
												assign node2783 = (inp[10]) ? node2787 : node2784;
													assign node2784 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node2787 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node2790 = (inp[4]) ? node2798 : node2791;
												assign node2791 = (inp[12]) ? node2795 : node2792;
													assign node2792 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node2795 = (inp[7]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node2798 = (inp[7]) ? node2800 : 15'b000000000111111;
													assign node2800 = (inp[10]) ? 15'b000000000011111 : 15'b000000000011111;
								assign node2803 = (inp[10]) ? node2861 : node2804;
									assign node2804 = (inp[7]) ? node2834 : node2805;
										assign node2805 = (inp[0]) ? node2819 : node2806;
											assign node2806 = (inp[14]) ? node2812 : node2807;
												assign node2807 = (inp[4]) ? 15'b000000111111111 : node2808;
													assign node2808 = (inp[1]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node2812 = (inp[12]) ? node2816 : node2813;
													assign node2813 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node2816 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node2819 = (inp[12]) ? node2827 : node2820;
												assign node2820 = (inp[4]) ? node2824 : node2821;
													assign node2821 = (inp[14]) ? 15'b000000011111111 : 15'b000000011111111;
													assign node2824 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node2827 = (inp[14]) ? node2831 : node2828;
													assign node2828 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node2831 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node2834 = (inp[1]) ? node2846 : node2835;
											assign node2835 = (inp[0]) ? node2841 : node2836;
												assign node2836 = (inp[4]) ? 15'b000000011111111 : node2837;
													assign node2837 = (inp[12]) ? 15'b000000111111111 : 15'b000000111111111;
												assign node2841 = (inp[4]) ? 15'b000000000111111 : node2842;
													assign node2842 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node2846 = (inp[12]) ? node2854 : node2847;
												assign node2847 = (inp[0]) ? node2851 : node2848;
													assign node2848 = (inp[14]) ? 15'b000000001111111 : 15'b000000001111111;
													assign node2851 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node2854 = (inp[0]) ? node2858 : node2855;
													assign node2855 = (inp[14]) ? 15'b000000000111111 : 15'b000000000111111;
													assign node2858 = (inp[4]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node2861 = (inp[14]) ? node2891 : node2862;
										assign node2862 = (inp[4]) ? node2876 : node2863;
											assign node2863 = (inp[2]) ? node2869 : node2864;
												assign node2864 = (inp[12]) ? node2866 : 15'b000000111111111;
													assign node2866 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node2869 = (inp[12]) ? node2873 : node2870;
													assign node2870 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node2873 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node2876 = (inp[12]) ? node2884 : node2877;
												assign node2877 = (inp[1]) ? node2881 : node2878;
													assign node2878 = (inp[7]) ? 15'b000000001111111 : 15'b000000001111111;
													assign node2881 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node2884 = (inp[0]) ? node2888 : node2885;
													assign node2885 = (inp[7]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node2888 = (inp[7]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node2891 = (inp[12]) ? node2907 : node2892;
											assign node2892 = (inp[4]) ? node2900 : node2893;
												assign node2893 = (inp[1]) ? node2897 : node2894;
													assign node2894 = (inp[2]) ? 15'b000000001111111 : 15'b000000001111111;
													assign node2897 = (inp[7]) ? 15'b000000000011111 : 15'b000000001111111;
												assign node2900 = (inp[2]) ? node2904 : node2901;
													assign node2901 = (inp[7]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node2904 = (inp[1]) ? 15'b000000000011111 : 15'b000000000011111;
											assign node2907 = (inp[2]) ? node2915 : node2908;
												assign node2908 = (inp[0]) ? node2912 : node2909;
													assign node2909 = (inp[1]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node2912 = (inp[7]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node2915 = (inp[4]) ? node2919 : node2916;
													assign node2916 = (inp[0]) ? 15'b000000000011111 : 15'b000000000011111;
													assign node2919 = (inp[0]) ? 15'b000000000001111 : 15'b000000000001111;
					assign node2922 = (inp[8]) ? node3394 : node2923;
						assign node2923 = (inp[1]) ? node3145 : node2924;
							assign node2924 = (inp[12]) ? node3036 : node2925;
								assign node2925 = (inp[14]) ? node2975 : node2926;
									assign node2926 = (inp[10]) ? node2954 : node2927;
										assign node2927 = (inp[0]) ? node2941 : node2928;
											assign node2928 = (inp[2]) ? node2936 : node2929;
												assign node2929 = (inp[4]) ? node2933 : node2930;
													assign node2930 = (inp[11]) ? 15'b000011111111111 : 15'b000111111111111;
													assign node2933 = (inp[7]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node2936 = (inp[7]) ? 15'b000000111111111 : node2937;
													assign node2937 = (inp[3]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node2941 = (inp[2]) ? node2949 : node2942;
												assign node2942 = (inp[3]) ? node2946 : node2943;
													assign node2943 = (inp[11]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node2946 = (inp[7]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node2949 = (inp[11]) ? 15'b000000111111111 : node2950;
													assign node2950 = (inp[4]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node2954 = (inp[3]) ? node2962 : node2955;
											assign node2955 = (inp[4]) ? 15'b000000111111111 : node2956;
												assign node2956 = (inp[11]) ? node2958 : 15'b000001111111111;
													assign node2958 = (inp[2]) ? 15'b000000111111111 : 15'b000000111111111;
											assign node2962 = (inp[11]) ? node2968 : node2963;
												assign node2963 = (inp[4]) ? node2965 : 15'b000000111111111;
													assign node2965 = (inp[0]) ? 15'b000000011111111 : 15'b000001111111111;
												assign node2968 = (inp[2]) ? node2972 : node2969;
													assign node2969 = (inp[7]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node2972 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node2975 = (inp[11]) ? node3007 : node2976;
										assign node2976 = (inp[3]) ? node2992 : node2977;
											assign node2977 = (inp[4]) ? node2985 : node2978;
												assign node2978 = (inp[0]) ? node2982 : node2979;
													assign node2979 = (inp[2]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node2982 = (inp[2]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node2985 = (inp[2]) ? node2989 : node2986;
													assign node2986 = (inp[7]) ? 15'b000000111111111 : 15'b000000111111111;
													assign node2989 = (inp[10]) ? 15'b000000001111111 : 15'b000000111111111;
											assign node2992 = (inp[0]) ? node3000 : node2993;
												assign node2993 = (inp[7]) ? node2997 : node2994;
													assign node2994 = (inp[10]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node2997 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node3000 = (inp[4]) ? node3004 : node3001;
													assign node3001 = (inp[7]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node3004 = (inp[10]) ? 15'b000000000111111 : 15'b000000011111111;
										assign node3007 = (inp[10]) ? node3023 : node3008;
											assign node3008 = (inp[7]) ? node3016 : node3009;
												assign node3009 = (inp[2]) ? node3013 : node3010;
													assign node3010 = (inp[0]) ? 15'b000000111111111 : 15'b000000111111111;
													assign node3013 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node3016 = (inp[2]) ? node3020 : node3017;
													assign node3017 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node3020 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node3023 = (inp[3]) ? node3031 : node3024;
												assign node3024 = (inp[4]) ? node3028 : node3025;
													assign node3025 = (inp[2]) ? 15'b000000001111111 : 15'b000000111111111;
													assign node3028 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node3031 = (inp[4]) ? node3033 : 15'b000000001111111;
													assign node3033 = (inp[7]) ? 15'b000000000111111 : 15'b000000001111111;
								assign node3036 = (inp[4]) ? node3090 : node3037;
									assign node3037 = (inp[10]) ? node3063 : node3038;
										assign node3038 = (inp[14]) ? node3054 : node3039;
											assign node3039 = (inp[11]) ? node3047 : node3040;
												assign node3040 = (inp[3]) ? node3044 : node3041;
													assign node3041 = (inp[2]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node3044 = (inp[0]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node3047 = (inp[2]) ? node3051 : node3048;
													assign node3048 = (inp[3]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node3051 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node3054 = (inp[7]) ? 15'b000000011111111 : node3055;
												assign node3055 = (inp[3]) ? node3059 : node3056;
													assign node3056 = (inp[0]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node3059 = (inp[11]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node3063 = (inp[7]) ? node3077 : node3064;
											assign node3064 = (inp[2]) ? node3072 : node3065;
												assign node3065 = (inp[14]) ? node3069 : node3066;
													assign node3066 = (inp[3]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node3069 = (inp[11]) ? 15'b000000001111111 : 15'b000000111111111;
												assign node3072 = (inp[0]) ? 15'b000000011111111 : node3073;
													assign node3073 = (inp[11]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node3077 = (inp[11]) ? node3083 : node3078;
												assign node3078 = (inp[14]) ? node3080 : 15'b000000011111111;
													assign node3080 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node3083 = (inp[2]) ? node3087 : node3084;
													assign node3084 = (inp[3]) ? 15'b000000001111111 : 15'b000000111111111;
													assign node3087 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node3090 = (inp[7]) ? node3118 : node3091;
										assign node3091 = (inp[0]) ? node3105 : node3092;
											assign node3092 = (inp[14]) ? node3100 : node3093;
												assign node3093 = (inp[2]) ? node3097 : node3094;
													assign node3094 = (inp[11]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node3097 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node3100 = (inp[11]) ? 15'b000000011111111 : node3101;
													assign node3101 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node3105 = (inp[11]) ? node3113 : node3106;
												assign node3106 = (inp[14]) ? node3110 : node3107;
													assign node3107 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node3110 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node3113 = (inp[2]) ? 15'b000000000111111 : node3114;
													assign node3114 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node3118 = (inp[3]) ? node3134 : node3119;
											assign node3119 = (inp[11]) ? node3127 : node3120;
												assign node3120 = (inp[10]) ? node3124 : node3121;
													assign node3121 = (inp[2]) ? 15'b000000011111111 : 15'b000000011111111;
													assign node3124 = (inp[14]) ? 15'b000000000111111 : 15'b000000011111111;
												assign node3127 = (inp[0]) ? node3131 : node3128;
													assign node3128 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node3131 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node3134 = (inp[0]) ? node3140 : node3135;
												assign node3135 = (inp[14]) ? node3137 : 15'b000000011111111;
													assign node3137 = (inp[11]) ? 15'b000000000011111 : 15'b000000001111111;
												assign node3140 = (inp[2]) ? node3142 : 15'b000000000111111;
													assign node3142 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
							assign node3145 = (inp[3]) ? node3273 : node3146;
								assign node3146 = (inp[0]) ? node3210 : node3147;
									assign node3147 = (inp[11]) ? node3179 : node3148;
										assign node3148 = (inp[14]) ? node3164 : node3149;
											assign node3149 = (inp[4]) ? node3157 : node3150;
												assign node3150 = (inp[12]) ? node3154 : node3151;
													assign node3151 = (inp[10]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node3154 = (inp[2]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node3157 = (inp[2]) ? node3161 : node3158;
													assign node3158 = (inp[10]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node3161 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node3164 = (inp[10]) ? node3172 : node3165;
												assign node3165 = (inp[12]) ? node3169 : node3166;
													assign node3166 = (inp[2]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node3169 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node3172 = (inp[7]) ? node3176 : node3173;
													assign node3173 = (inp[12]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node3176 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node3179 = (inp[7]) ? node3195 : node3180;
											assign node3180 = (inp[14]) ? node3188 : node3181;
												assign node3181 = (inp[4]) ? node3185 : node3182;
													assign node3182 = (inp[2]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node3185 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node3188 = (inp[2]) ? node3192 : node3189;
													assign node3189 = (inp[12]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node3192 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node3195 = (inp[2]) ? node3203 : node3196;
												assign node3196 = (inp[4]) ? node3200 : node3197;
													assign node3197 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node3200 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node3203 = (inp[10]) ? node3207 : node3204;
													assign node3204 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node3207 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node3210 = (inp[4]) ? node3242 : node3211;
										assign node3211 = (inp[11]) ? node3227 : node3212;
											assign node3212 = (inp[7]) ? node3220 : node3213;
												assign node3213 = (inp[2]) ? node3217 : node3214;
													assign node3214 = (inp[14]) ? 15'b000000111111111 : 15'b000000111111111;
													assign node3217 = (inp[12]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node3220 = (inp[14]) ? node3224 : node3221;
													assign node3221 = (inp[2]) ? 15'b000000011111111 : 15'b000001111111111;
													assign node3224 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node3227 = (inp[10]) ? node3235 : node3228;
												assign node3228 = (inp[7]) ? node3232 : node3229;
													assign node3229 = (inp[12]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node3232 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node3235 = (inp[14]) ? node3239 : node3236;
													assign node3236 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node3239 = (inp[7]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node3242 = (inp[7]) ? node3258 : node3243;
											assign node3243 = (inp[11]) ? node3251 : node3244;
												assign node3244 = (inp[12]) ? node3248 : node3245;
													assign node3245 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node3248 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node3251 = (inp[12]) ? node3255 : node3252;
													assign node3252 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node3255 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node3258 = (inp[2]) ? node3266 : node3259;
												assign node3259 = (inp[14]) ? node3263 : node3260;
													assign node3260 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node3263 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node3266 = (inp[10]) ? node3270 : node3267;
													assign node3267 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node3270 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
								assign node3273 = (inp[0]) ? node3335 : node3274;
									assign node3274 = (inp[2]) ? node3306 : node3275;
										assign node3275 = (inp[7]) ? node3291 : node3276;
											assign node3276 = (inp[10]) ? node3284 : node3277;
												assign node3277 = (inp[4]) ? node3281 : node3278;
													assign node3278 = (inp[11]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node3281 = (inp[12]) ? 15'b000000011111111 : 15'b000000011111111;
												assign node3284 = (inp[12]) ? node3288 : node3285;
													assign node3285 = (inp[11]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node3288 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node3291 = (inp[14]) ? node3299 : node3292;
												assign node3292 = (inp[10]) ? node3296 : node3293;
													assign node3293 = (inp[11]) ? 15'b000000011111111 : 15'b000000011111111;
													assign node3296 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node3299 = (inp[11]) ? node3303 : node3300;
													assign node3300 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node3303 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node3306 = (inp[4]) ? node3320 : node3307;
											assign node3307 = (inp[12]) ? node3313 : node3308;
												assign node3308 = (inp[10]) ? node3310 : 15'b000000111111111;
													assign node3310 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node3313 = (inp[7]) ? node3317 : node3314;
													assign node3314 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node3317 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node3320 = (inp[11]) ? node3328 : node3321;
												assign node3321 = (inp[10]) ? node3325 : node3322;
													assign node3322 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node3325 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node3328 = (inp[7]) ? node3332 : node3329;
													assign node3329 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node3332 = (inp[12]) ? 15'b000000000011111 : 15'b000000000011111;
									assign node3335 = (inp[11]) ? node3367 : node3336;
										assign node3336 = (inp[2]) ? node3352 : node3337;
											assign node3337 = (inp[4]) ? node3345 : node3338;
												assign node3338 = (inp[12]) ? node3342 : node3339;
													assign node3339 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node3342 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node3345 = (inp[14]) ? node3349 : node3346;
													assign node3346 = (inp[7]) ? 15'b000000000111111 : 15'b000000011111111;
													assign node3349 = (inp[10]) ? 15'b000000000011111 : 15'b000000001111111;
											assign node3352 = (inp[10]) ? node3360 : node3353;
												assign node3353 = (inp[12]) ? node3357 : node3354;
													assign node3354 = (inp[7]) ? 15'b000000001111111 : 15'b000000001111111;
													assign node3357 = (inp[4]) ? 15'b000000000011111 : 15'b000000001111111;
												assign node3360 = (inp[4]) ? node3364 : node3361;
													assign node3361 = (inp[14]) ? 15'b000000000111111 : 15'b000000000111111;
													assign node3364 = (inp[12]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node3367 = (inp[12]) ? node3381 : node3368;
											assign node3368 = (inp[2]) ? node3374 : node3369;
												assign node3369 = (inp[4]) ? node3371 : 15'b000000011111111;
													assign node3371 = (inp[14]) ? 15'b000000001111111 : 15'b000000000111111;
												assign node3374 = (inp[7]) ? node3378 : node3375;
													assign node3375 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node3378 = (inp[4]) ? 15'b000000000001111 : 15'b000000000111111;
											assign node3381 = (inp[7]) ? node3387 : node3382;
												assign node3382 = (inp[14]) ? node3384 : 15'b000000000111111;
													assign node3384 = (inp[10]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node3387 = (inp[2]) ? node3391 : node3388;
													assign node3388 = (inp[10]) ? 15'b000000000011111 : 15'b000000000011111;
													assign node3391 = (inp[10]) ? 15'b000000000001111 : 15'b000000000011111;
						assign node3394 = (inp[14]) ? node3640 : node3395;
							assign node3395 = (inp[7]) ? node3523 : node3396;
								assign node3396 = (inp[11]) ? node3460 : node3397;
									assign node3397 = (inp[2]) ? node3429 : node3398;
										assign node3398 = (inp[10]) ? node3414 : node3399;
											assign node3399 = (inp[0]) ? node3407 : node3400;
												assign node3400 = (inp[12]) ? node3404 : node3401;
													assign node3401 = (inp[4]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node3404 = (inp[1]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node3407 = (inp[4]) ? node3411 : node3408;
													assign node3408 = (inp[3]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node3411 = (inp[12]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node3414 = (inp[12]) ? node3422 : node3415;
												assign node3415 = (inp[1]) ? node3419 : node3416;
													assign node3416 = (inp[0]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node3419 = (inp[3]) ? 15'b000000001111111 : 15'b000000111111111;
												assign node3422 = (inp[3]) ? node3426 : node3423;
													assign node3423 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node3426 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node3429 = (inp[12]) ? node3445 : node3430;
											assign node3430 = (inp[4]) ? node3438 : node3431;
												assign node3431 = (inp[10]) ? node3435 : node3432;
													assign node3432 = (inp[0]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node3435 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node3438 = (inp[1]) ? node3442 : node3439;
													assign node3439 = (inp[3]) ? 15'b000000011111111 : 15'b000001111111111;
													assign node3442 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node3445 = (inp[4]) ? node3453 : node3446;
												assign node3446 = (inp[0]) ? node3450 : node3447;
													assign node3447 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node3450 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node3453 = (inp[0]) ? node3457 : node3454;
													assign node3454 = (inp[3]) ? 15'b000000001111111 : 15'b000000001111111;
													assign node3457 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node3460 = (inp[4]) ? node3492 : node3461;
										assign node3461 = (inp[10]) ? node3477 : node3462;
											assign node3462 = (inp[12]) ? node3470 : node3463;
												assign node3463 = (inp[0]) ? node3467 : node3464;
													assign node3464 = (inp[1]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node3467 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node3470 = (inp[1]) ? node3474 : node3471;
													assign node3471 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node3474 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node3477 = (inp[0]) ? node3485 : node3478;
												assign node3478 = (inp[3]) ? node3482 : node3479;
													assign node3479 = (inp[12]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node3482 = (inp[1]) ? 15'b000000000111111 : 15'b000000011111111;
												assign node3485 = (inp[12]) ? node3489 : node3486;
													assign node3486 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node3489 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node3492 = (inp[2]) ? node3508 : node3493;
											assign node3493 = (inp[3]) ? node3501 : node3494;
												assign node3494 = (inp[10]) ? node3498 : node3495;
													assign node3495 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node3498 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node3501 = (inp[0]) ? node3505 : node3502;
													assign node3502 = (inp[12]) ? 15'b000000000111111 : 15'b000000011111111;
													assign node3505 = (inp[12]) ? 15'b000000000111111 : 15'b000000000111111;
											assign node3508 = (inp[3]) ? node3516 : node3509;
												assign node3509 = (inp[12]) ? node3513 : node3510;
													assign node3510 = (inp[0]) ? 15'b000000000111111 : 15'b000000011111111;
													assign node3513 = (inp[1]) ? 15'b000000000111111 : 15'b000000000111111;
												assign node3516 = (inp[10]) ? node3520 : node3517;
													assign node3517 = (inp[12]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node3520 = (inp[12]) ? 15'b000000000001111 : 15'b000000000011111;
								assign node3523 = (inp[12]) ? node3583 : node3524;
									assign node3524 = (inp[11]) ? node3554 : node3525;
										assign node3525 = (inp[0]) ? node3541 : node3526;
											assign node3526 = (inp[10]) ? node3534 : node3527;
												assign node3527 = (inp[1]) ? node3531 : node3528;
													assign node3528 = (inp[2]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node3531 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node3534 = (inp[1]) ? node3538 : node3535;
													assign node3535 = (inp[2]) ? 15'b000000011111111 : 15'b000000011111111;
													assign node3538 = (inp[4]) ? 15'b000000000111111 : 15'b000000011111111;
											assign node3541 = (inp[1]) ? node3547 : node3542;
												assign node3542 = (inp[3]) ? node3544 : 15'b000000111111111;
													assign node3544 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node3547 = (inp[3]) ? node3551 : node3548;
													assign node3548 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node3551 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node3554 = (inp[2]) ? node3570 : node3555;
											assign node3555 = (inp[10]) ? node3563 : node3556;
												assign node3556 = (inp[4]) ? node3560 : node3557;
													assign node3557 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node3560 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node3563 = (inp[4]) ? node3567 : node3564;
													assign node3564 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node3567 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node3570 = (inp[3]) ? node3576 : node3571;
												assign node3571 = (inp[0]) ? 15'b000000001111111 : node3572;
													assign node3572 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node3576 = (inp[0]) ? node3580 : node3577;
													assign node3577 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node3580 = (inp[10]) ? 15'b000000000001111 : 15'b000000000111111;
									assign node3583 = (inp[1]) ? node3609 : node3584;
										assign node3584 = (inp[0]) ? node3596 : node3585;
											assign node3585 = (inp[3]) ? node3591 : node3586;
												assign node3586 = (inp[10]) ? 15'b000000000111111 : node3587;
													assign node3587 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node3591 = (inp[11]) ? 15'b000000001111111 : node3592;
													assign node3592 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node3596 = (inp[11]) ? node3604 : node3597;
												assign node3597 = (inp[3]) ? node3601 : node3598;
													assign node3598 = (inp[2]) ? 15'b000000001111111 : 15'b000000001111111;
													assign node3601 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node3604 = (inp[4]) ? 15'b000000000011111 : node3605;
													assign node3605 = (inp[2]) ? 15'b000000000111111 : 15'b000000000111111;
										assign node3609 = (inp[4]) ? node3625 : node3610;
											assign node3610 = (inp[2]) ? node3618 : node3611;
												assign node3611 = (inp[10]) ? node3615 : node3612;
													assign node3612 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node3615 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node3618 = (inp[11]) ? node3622 : node3619;
													assign node3619 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node3622 = (inp[0]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node3625 = (inp[0]) ? node3633 : node3626;
												assign node3626 = (inp[2]) ? node3630 : node3627;
													assign node3627 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node3630 = (inp[10]) ? 15'b000000000011111 : 15'b000000000011111;
												assign node3633 = (inp[11]) ? node3637 : node3634;
													assign node3634 = (inp[10]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node3637 = (inp[10]) ? 15'b000000000001111 : 15'b000000000011111;
							assign node3640 = (inp[10]) ? node3764 : node3641;
								assign node3641 = (inp[3]) ? node3705 : node3642;
									assign node3642 = (inp[1]) ? node3674 : node3643;
										assign node3643 = (inp[7]) ? node3659 : node3644;
											assign node3644 = (inp[4]) ? node3652 : node3645;
												assign node3645 = (inp[11]) ? node3649 : node3646;
													assign node3646 = (inp[2]) ? 15'b000000011111111 : 15'b000001111111111;
													assign node3649 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node3652 = (inp[11]) ? node3656 : node3653;
													assign node3653 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node3656 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node3659 = (inp[11]) ? node3667 : node3660;
												assign node3660 = (inp[4]) ? node3664 : node3661;
													assign node3661 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node3664 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node3667 = (inp[0]) ? node3671 : node3668;
													assign node3668 = (inp[12]) ? 15'b000000000111111 : 15'b000000011111111;
													assign node3671 = (inp[2]) ? 15'b000000000011111 : 15'b000000001111111;
										assign node3674 = (inp[7]) ? node3690 : node3675;
											assign node3675 = (inp[0]) ? node3683 : node3676;
												assign node3676 = (inp[2]) ? node3680 : node3677;
													assign node3677 = (inp[11]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node3680 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node3683 = (inp[4]) ? node3687 : node3684;
													assign node3684 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node3687 = (inp[11]) ? 15'b000000000111111 : 15'b000000000111111;
											assign node3690 = (inp[12]) ? node3698 : node3691;
												assign node3691 = (inp[0]) ? node3695 : node3692;
													assign node3692 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node3695 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node3698 = (inp[4]) ? node3702 : node3699;
													assign node3699 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node3702 = (inp[11]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node3705 = (inp[7]) ? node3737 : node3706;
										assign node3706 = (inp[12]) ? node3722 : node3707;
											assign node3707 = (inp[1]) ? node3715 : node3708;
												assign node3708 = (inp[0]) ? node3712 : node3709;
													assign node3709 = (inp[11]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node3712 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node3715 = (inp[11]) ? node3719 : node3716;
													assign node3716 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node3719 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node3722 = (inp[11]) ? node3730 : node3723;
												assign node3723 = (inp[0]) ? node3727 : node3724;
													assign node3724 = (inp[4]) ? 15'b000000001111111 : 15'b000000001111111;
													assign node3727 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node3730 = (inp[1]) ? node3734 : node3731;
													assign node3731 = (inp[2]) ? 15'b000000000111111 : 15'b000000011111111;
													assign node3734 = (inp[4]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node3737 = (inp[4]) ? node3751 : node3738;
											assign node3738 = (inp[1]) ? node3744 : node3739;
												assign node3739 = (inp[0]) ? node3741 : 15'b000000001111111;
													assign node3741 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node3744 = (inp[2]) ? node3748 : node3745;
													assign node3745 = (inp[12]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node3748 = (inp[0]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node3751 = (inp[0]) ? node3759 : node3752;
												assign node3752 = (inp[11]) ? node3756 : node3753;
													assign node3753 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node3756 = (inp[2]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node3759 = (inp[1]) ? 15'b000000000001111 : node3760;
													assign node3760 = (inp[2]) ? 15'b000000000011111 : 15'b000000000111111;
								assign node3764 = (inp[4]) ? node3824 : node3765;
									assign node3765 = (inp[0]) ? node3795 : node3766;
										assign node3766 = (inp[3]) ? node3782 : node3767;
											assign node3767 = (inp[11]) ? node3775 : node3768;
												assign node3768 = (inp[7]) ? node3772 : node3769;
													assign node3769 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node3772 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node3775 = (inp[1]) ? node3779 : node3776;
													assign node3776 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node3779 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node3782 = (inp[1]) ? node3790 : node3783;
												assign node3783 = (inp[11]) ? node3787 : node3784;
													assign node3784 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node3787 = (inp[12]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node3790 = (inp[7]) ? 15'b000000000111111 : node3791;
													assign node3791 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node3795 = (inp[2]) ? node3811 : node3796;
											assign node3796 = (inp[1]) ? node3804 : node3797;
												assign node3797 = (inp[3]) ? node3801 : node3798;
													assign node3798 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node3801 = (inp[11]) ? 15'b000000000011111 : 15'b000000001111111;
												assign node3804 = (inp[3]) ? node3808 : node3805;
													assign node3805 = (inp[7]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node3808 = (inp[7]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node3811 = (inp[3]) ? node3817 : node3812;
												assign node3812 = (inp[11]) ? node3814 : 15'b000000000111111;
													assign node3814 = (inp[1]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node3817 = (inp[12]) ? node3821 : node3818;
													assign node3818 = (inp[11]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node3821 = (inp[11]) ? 15'b000000000001111 : 15'b000000000001111;
									assign node3824 = (inp[2]) ? node3856 : node3825;
										assign node3825 = (inp[1]) ? node3841 : node3826;
											assign node3826 = (inp[12]) ? node3834 : node3827;
												assign node3827 = (inp[0]) ? node3831 : node3828;
													assign node3828 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node3831 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node3834 = (inp[11]) ? node3838 : node3835;
													assign node3835 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node3838 = (inp[0]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node3841 = (inp[11]) ? node3849 : node3842;
												assign node3842 = (inp[3]) ? node3846 : node3843;
													assign node3843 = (inp[12]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node3846 = (inp[0]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node3849 = (inp[12]) ? node3853 : node3850;
													assign node3850 = (inp[0]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node3853 = (inp[0]) ? 15'b000000000000111 : 15'b000000000011111;
										assign node3856 = (inp[12]) ? node3872 : node3857;
											assign node3857 = (inp[1]) ? node3865 : node3858;
												assign node3858 = (inp[3]) ? node3862 : node3859;
													assign node3859 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node3862 = (inp[11]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node3865 = (inp[11]) ? node3869 : node3866;
													assign node3866 = (inp[3]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node3869 = (inp[7]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node3872 = (inp[7]) ? node3880 : node3873;
												assign node3873 = (inp[0]) ? node3877 : node3874;
													assign node3874 = (inp[3]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node3877 = (inp[11]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node3880 = (inp[3]) ? node3884 : node3881;
													assign node3881 = (inp[0]) ? 15'b000000000001111 : 15'b000000000011111;
													assign node3884 = (inp[0]) ? 15'b000000000000111 : 15'b000000000001111;
			assign node3887 = (inp[7]) ? node5809 : node3888;
				assign node3888 = (inp[12]) ? node4848 : node3889;
					assign node3889 = (inp[13]) ? node4363 : node3890;
						assign node3890 = (inp[11]) ? node4132 : node3891;
							assign node3891 = (inp[9]) ? node4005 : node3892;
								assign node3892 = (inp[3]) ? node3952 : node3893;
									assign node3893 = (inp[1]) ? node3923 : node3894;
										assign node3894 = (inp[4]) ? node3908 : node3895;
											assign node3895 = (inp[0]) ? node3903 : node3896;
												assign node3896 = (inp[2]) ? node3900 : node3897;
													assign node3897 = (inp[10]) ? 15'b000111111111111 : 15'b001111111111111;
													assign node3900 = (inp[8]) ? 15'b000011111111111 : 15'b000111111111111;
												assign node3903 = (inp[10]) ? 15'b000011111111111 : node3904;
													assign node3904 = (inp[14]) ? 15'b000011111111111 : 15'b000111111111111;
											assign node3908 = (inp[8]) ? node3916 : node3909;
												assign node3909 = (inp[2]) ? node3913 : node3910;
													assign node3910 = (inp[10]) ? 15'b000011111111111 : 15'b000111111111111;
													assign node3913 = (inp[0]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node3916 = (inp[14]) ? node3920 : node3917;
													assign node3917 = (inp[0]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node3920 = (inp[0]) ? 15'b000000011111111 : 15'b000001111111111;
										assign node3923 = (inp[10]) ? node3937 : node3924;
											assign node3924 = (inp[0]) ? node3932 : node3925;
												assign node3925 = (inp[2]) ? node3929 : node3926;
													assign node3926 = (inp[4]) ? 15'b000011111111111 : 15'b000111111111111;
													assign node3929 = (inp[8]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node3932 = (inp[8]) ? 15'b000001111111111 : node3933;
													assign node3933 = (inp[2]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node3937 = (inp[4]) ? node3945 : node3938;
												assign node3938 = (inp[2]) ? node3942 : node3939;
													assign node3939 = (inp[14]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node3942 = (inp[14]) ? 15'b000000011111111 : 15'b000001111111111;
												assign node3945 = (inp[0]) ? node3949 : node3946;
													assign node3946 = (inp[8]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node3949 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node3952 = (inp[2]) ? node3974 : node3953;
										assign node3953 = (inp[14]) ? node3967 : node3954;
											assign node3954 = (inp[1]) ? node3962 : node3955;
												assign node3955 = (inp[10]) ? node3959 : node3956;
													assign node3956 = (inp[0]) ? 15'b000011111111111 : 15'b000111111111111;
													assign node3959 = (inp[0]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node3962 = (inp[0]) ? node3964 : 15'b000001111111111;
													assign node3964 = (inp[10]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node3967 = (inp[4]) ? node3969 : 15'b000011111111111;
												assign node3969 = (inp[1]) ? 15'b000000111111111 : node3970;
													assign node3970 = (inp[10]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node3974 = (inp[8]) ? node3990 : node3975;
											assign node3975 = (inp[4]) ? node3983 : node3976;
												assign node3976 = (inp[0]) ? node3980 : node3977;
													assign node3977 = (inp[1]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node3980 = (inp[10]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node3983 = (inp[14]) ? node3987 : node3984;
													assign node3984 = (inp[10]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node3987 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node3990 = (inp[14]) ? node3998 : node3991;
												assign node3991 = (inp[0]) ? node3995 : node3992;
													assign node3992 = (inp[1]) ? 15'b000000111111111 : 15'b000000111111111;
													assign node3995 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node3998 = (inp[4]) ? node4002 : node3999;
													assign node3999 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node4002 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
								assign node4005 = (inp[3]) ? node4069 : node4006;
									assign node4006 = (inp[4]) ? node4038 : node4007;
										assign node4007 = (inp[14]) ? node4023 : node4008;
											assign node4008 = (inp[8]) ? node4016 : node4009;
												assign node4009 = (inp[0]) ? node4013 : node4010;
													assign node4010 = (inp[2]) ? 15'b000011111111111 : 15'b000111111111111;
													assign node4013 = (inp[1]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node4016 = (inp[2]) ? node4020 : node4017;
													assign node4017 = (inp[10]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node4020 = (inp[0]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node4023 = (inp[2]) ? node4031 : node4024;
												assign node4024 = (inp[8]) ? node4028 : node4025;
													assign node4025 = (inp[0]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node4028 = (inp[0]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node4031 = (inp[0]) ? node4035 : node4032;
													assign node4032 = (inp[1]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node4035 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node4038 = (inp[0]) ? node4054 : node4039;
											assign node4039 = (inp[1]) ? node4047 : node4040;
												assign node4040 = (inp[2]) ? node4044 : node4041;
													assign node4041 = (inp[14]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node4044 = (inp[10]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node4047 = (inp[2]) ? node4051 : node4048;
													assign node4048 = (inp[10]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node4051 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node4054 = (inp[10]) ? node4062 : node4055;
												assign node4055 = (inp[8]) ? node4059 : node4056;
													assign node4056 = (inp[1]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node4059 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node4062 = (inp[14]) ? node4066 : node4063;
													assign node4063 = (inp[8]) ? 15'b000000011111111 : 15'b000001111111111;
													assign node4066 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node4069 = (inp[8]) ? node4101 : node4070;
										assign node4070 = (inp[4]) ? node4086 : node4071;
											assign node4071 = (inp[0]) ? node4079 : node4072;
												assign node4072 = (inp[2]) ? node4076 : node4073;
													assign node4073 = (inp[14]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node4076 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node4079 = (inp[1]) ? node4083 : node4080;
													assign node4080 = (inp[2]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node4083 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node4086 = (inp[0]) ? node4094 : node4087;
												assign node4087 = (inp[10]) ? node4091 : node4088;
													assign node4088 = (inp[2]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node4091 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node4094 = (inp[14]) ? node4098 : node4095;
													assign node4095 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node4098 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node4101 = (inp[14]) ? node4117 : node4102;
											assign node4102 = (inp[10]) ? node4110 : node4103;
												assign node4103 = (inp[2]) ? node4107 : node4104;
													assign node4104 = (inp[4]) ? 15'b000000111111111 : 15'b000000111111111;
													assign node4107 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node4110 = (inp[2]) ? node4114 : node4111;
													assign node4111 = (inp[0]) ? 15'b000000011111111 : 15'b000000011111111;
													assign node4114 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node4117 = (inp[2]) ? node4125 : node4118;
												assign node4118 = (inp[4]) ? node4122 : node4119;
													assign node4119 = (inp[10]) ? 15'b000000111111111 : 15'b000000011111111;
													assign node4122 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node4125 = (inp[1]) ? node4129 : node4126;
													assign node4126 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node4129 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
							assign node4132 = (inp[2]) ? node4248 : node4133;
								assign node4133 = (inp[4]) ? node4189 : node4134;
									assign node4134 = (inp[14]) ? node4160 : node4135;
										assign node4135 = (inp[3]) ? node4151 : node4136;
											assign node4136 = (inp[1]) ? node4144 : node4137;
												assign node4137 = (inp[9]) ? node4141 : node4138;
													assign node4138 = (inp[0]) ? 15'b000001111111111 : 15'b000111111111111;
													assign node4141 = (inp[8]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node4144 = (inp[10]) ? node4148 : node4145;
													assign node4145 = (inp[9]) ? 15'b000001111111111 : 15'b000001111111111;
													assign node4148 = (inp[0]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node4151 = (inp[8]) ? node4157 : node4152;
												assign node4152 = (inp[1]) ? node4154 : 15'b000001111111111;
													assign node4154 = (inp[9]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node4157 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node4160 = (inp[8]) ? node4174 : node4161;
											assign node4161 = (inp[0]) ? node4167 : node4162;
												assign node4162 = (inp[1]) ? node4164 : 15'b000001111111111;
													assign node4164 = (inp[3]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node4167 = (inp[3]) ? node4171 : node4168;
													assign node4168 = (inp[1]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node4171 = (inp[9]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node4174 = (inp[10]) ? node4182 : node4175;
												assign node4175 = (inp[9]) ? node4179 : node4176;
													assign node4176 = (inp[1]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node4179 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node4182 = (inp[0]) ? node4186 : node4183;
													assign node4183 = (inp[9]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node4186 = (inp[9]) ? 15'b000000000111111 : 15'b000000011111111;
									assign node4189 = (inp[8]) ? node4217 : node4190;
										assign node4190 = (inp[1]) ? node4206 : node4191;
											assign node4191 = (inp[0]) ? node4199 : node4192;
												assign node4192 = (inp[3]) ? node4196 : node4193;
													assign node4193 = (inp[14]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node4196 = (inp[9]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node4199 = (inp[10]) ? node4203 : node4200;
													assign node4200 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node4203 = (inp[3]) ? 15'b000000001111111 : 15'b000000111111111;
											assign node4206 = (inp[14]) ? node4212 : node4207;
												assign node4207 = (inp[10]) ? 15'b000000111111111 : node4208;
													assign node4208 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node4212 = (inp[10]) ? 15'b000000001111111 : node4213;
													assign node4213 = (inp[3]) ? 15'b000000011111111 : 15'b000000011111111;
										assign node4217 = (inp[10]) ? node4233 : node4218;
											assign node4218 = (inp[0]) ? node4226 : node4219;
												assign node4219 = (inp[14]) ? node4223 : node4220;
													assign node4220 = (inp[1]) ? 15'b000000111111111 : 15'b000000111111111;
													assign node4223 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node4226 = (inp[9]) ? node4230 : node4227;
													assign node4227 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node4230 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node4233 = (inp[0]) ? node4241 : node4234;
												assign node4234 = (inp[14]) ? node4238 : node4235;
													assign node4235 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node4238 = (inp[9]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node4241 = (inp[1]) ? node4245 : node4242;
													assign node4242 = (inp[9]) ? 15'b000000001111111 : 15'b000000111111111;
													assign node4245 = (inp[9]) ? 15'b000000000111111 : 15'b000000001111111;
								assign node4248 = (inp[14]) ? node4302 : node4249;
									assign node4249 = (inp[10]) ? node4277 : node4250;
										assign node4250 = (inp[1]) ? node4262 : node4251;
											assign node4251 = (inp[0]) ? node4257 : node4252;
												assign node4252 = (inp[9]) ? node4254 : 15'b000011111111111;
													assign node4254 = (inp[8]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node4257 = (inp[3]) ? 15'b000000111111111 : node4258;
													assign node4258 = (inp[8]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node4262 = (inp[0]) ? node4270 : node4263;
												assign node4263 = (inp[8]) ? node4267 : node4264;
													assign node4264 = (inp[9]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node4267 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node4270 = (inp[4]) ? node4274 : node4271;
													assign node4271 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node4274 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node4277 = (inp[3]) ? node4293 : node4278;
											assign node4278 = (inp[8]) ? node4286 : node4279;
												assign node4279 = (inp[4]) ? node4283 : node4280;
													assign node4280 = (inp[1]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node4283 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node4286 = (inp[1]) ? node4290 : node4287;
													assign node4287 = (inp[9]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node4290 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node4293 = (inp[4]) ? node4295 : 15'b000000011111111;
												assign node4295 = (inp[0]) ? node4299 : node4296;
													assign node4296 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node4299 = (inp[9]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node4302 = (inp[4]) ? node4334 : node4303;
										assign node4303 = (inp[1]) ? node4319 : node4304;
											assign node4304 = (inp[10]) ? node4312 : node4305;
												assign node4305 = (inp[0]) ? node4309 : node4306;
													assign node4306 = (inp[8]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node4309 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node4312 = (inp[9]) ? node4316 : node4313;
													assign node4313 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node4316 = (inp[8]) ? 15'b000000000111111 : 15'b000000011111111;
											assign node4319 = (inp[9]) ? node4327 : node4320;
												assign node4320 = (inp[10]) ? node4324 : node4321;
													assign node4321 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node4324 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node4327 = (inp[8]) ? node4331 : node4328;
													assign node4328 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node4331 = (inp[10]) ? 15'b000000000011111 : 15'b000000001111111;
										assign node4334 = (inp[8]) ? node4348 : node4335;
											assign node4335 = (inp[3]) ? node4341 : node4336;
												assign node4336 = (inp[1]) ? 15'b000000011111111 : node4337;
													assign node4337 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node4341 = (inp[9]) ? node4345 : node4342;
													assign node4342 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node4345 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node4348 = (inp[0]) ? node4356 : node4349;
												assign node4349 = (inp[1]) ? node4353 : node4350;
													assign node4350 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node4353 = (inp[9]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node4356 = (inp[3]) ? node4360 : node4357;
													assign node4357 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node4360 = (inp[1]) ? 15'b000000000011111 : 15'b000000000111111;
						assign node4363 = (inp[9]) ? node4609 : node4364;
							assign node4364 = (inp[14]) ? node4490 : node4365;
								assign node4365 = (inp[4]) ? node4427 : node4366;
									assign node4366 = (inp[0]) ? node4396 : node4367;
										assign node4367 = (inp[2]) ? node4383 : node4368;
											assign node4368 = (inp[11]) ? node4376 : node4369;
												assign node4369 = (inp[10]) ? node4373 : node4370;
													assign node4370 = (inp[1]) ? 15'b000011111111111 : 15'b000111111111111;
													assign node4373 = (inp[8]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node4376 = (inp[10]) ? node4380 : node4377;
													assign node4377 = (inp[3]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node4380 = (inp[1]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node4383 = (inp[3]) ? node4389 : node4384;
												assign node4384 = (inp[1]) ? 15'b000001111111111 : node4385;
													assign node4385 = (inp[10]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node4389 = (inp[11]) ? node4393 : node4390;
													assign node4390 = (inp[10]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node4393 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node4396 = (inp[10]) ? node4412 : node4397;
											assign node4397 = (inp[8]) ? node4405 : node4398;
												assign node4398 = (inp[3]) ? node4402 : node4399;
													assign node4399 = (inp[11]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node4402 = (inp[11]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node4405 = (inp[1]) ? node4409 : node4406;
													assign node4406 = (inp[3]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node4409 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node4412 = (inp[3]) ? node4420 : node4413;
												assign node4413 = (inp[2]) ? node4417 : node4414;
													assign node4414 = (inp[1]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node4417 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node4420 = (inp[11]) ? node4424 : node4421;
													assign node4421 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node4424 = (inp[1]) ? 15'b000000001111111 : 15'b000000111111111;
									assign node4427 = (inp[1]) ? node4459 : node4428;
										assign node4428 = (inp[8]) ? node4444 : node4429;
											assign node4429 = (inp[2]) ? node4437 : node4430;
												assign node4430 = (inp[11]) ? node4434 : node4431;
													assign node4431 = (inp[3]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node4434 = (inp[3]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node4437 = (inp[3]) ? node4441 : node4438;
													assign node4438 = (inp[11]) ? 15'b000000111111111 : 15'b000000111111111;
													assign node4441 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node4444 = (inp[11]) ? node4452 : node4445;
												assign node4445 = (inp[0]) ? node4449 : node4446;
													assign node4446 = (inp[10]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node4449 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node4452 = (inp[3]) ? node4456 : node4453;
													assign node4453 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node4456 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node4459 = (inp[3]) ? node4475 : node4460;
											assign node4460 = (inp[2]) ? node4468 : node4461;
												assign node4461 = (inp[0]) ? node4465 : node4462;
													assign node4462 = (inp[8]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node4465 = (inp[11]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node4468 = (inp[0]) ? node4472 : node4469;
													assign node4469 = (inp[8]) ? 15'b000000011111111 : 15'b000000011111111;
													assign node4472 = (inp[8]) ? 15'b000000001111111 : 15'b000000001111111;
											assign node4475 = (inp[0]) ? node4483 : node4476;
												assign node4476 = (inp[10]) ? node4480 : node4477;
													assign node4477 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node4480 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node4483 = (inp[10]) ? node4487 : node4484;
													assign node4484 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node4487 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
								assign node4490 = (inp[2]) ? node4550 : node4491;
									assign node4491 = (inp[10]) ? node4521 : node4492;
										assign node4492 = (inp[8]) ? node4506 : node4493;
											assign node4493 = (inp[3]) ? node4501 : node4494;
												assign node4494 = (inp[0]) ? node4498 : node4495;
													assign node4495 = (inp[4]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node4498 = (inp[4]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node4501 = (inp[1]) ? 15'b000000111111111 : node4502;
													assign node4502 = (inp[0]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node4506 = (inp[1]) ? node4514 : node4507;
												assign node4507 = (inp[0]) ? node4511 : node4508;
													assign node4508 = (inp[3]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node4511 = (inp[11]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node4514 = (inp[4]) ? node4518 : node4515;
													assign node4515 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node4518 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node4521 = (inp[4]) ? node4535 : node4522;
											assign node4522 = (inp[0]) ? node4530 : node4523;
												assign node4523 = (inp[1]) ? node4527 : node4524;
													assign node4524 = (inp[11]) ? 15'b000000111111111 : 15'b000000111111111;
													assign node4527 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node4530 = (inp[8]) ? 15'b000000011111111 : node4531;
													assign node4531 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node4535 = (inp[1]) ? node4543 : node4536;
												assign node4536 = (inp[8]) ? node4540 : node4537;
													assign node4537 = (inp[11]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node4540 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node4543 = (inp[3]) ? node4547 : node4544;
													assign node4544 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node4547 = (inp[11]) ? 15'b000000000011111 : 15'b000000001111111;
									assign node4550 = (inp[10]) ? node4580 : node4551;
										assign node4551 = (inp[4]) ? node4565 : node4552;
											assign node4552 = (inp[3]) ? node4560 : node4553;
												assign node4553 = (inp[0]) ? node4557 : node4554;
													assign node4554 = (inp[8]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node4557 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node4560 = (inp[11]) ? 15'b000000011111111 : node4561;
													assign node4561 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node4565 = (inp[11]) ? node4573 : node4566;
												assign node4566 = (inp[1]) ? node4570 : node4567;
													assign node4567 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node4570 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node4573 = (inp[0]) ? node4577 : node4574;
													assign node4574 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node4577 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node4580 = (inp[8]) ? node4596 : node4581;
											assign node4581 = (inp[3]) ? node4589 : node4582;
												assign node4582 = (inp[1]) ? node4586 : node4583;
													assign node4583 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node4586 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node4589 = (inp[1]) ? node4593 : node4590;
													assign node4590 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node4593 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node4596 = (inp[11]) ? node4602 : node4597;
												assign node4597 = (inp[4]) ? 15'b000000000111111 : node4598;
													assign node4598 = (inp[3]) ? 15'b000000000111111 : 15'b000000011111111;
												assign node4602 = (inp[3]) ? node4606 : node4603;
													assign node4603 = (inp[0]) ? 15'b000000000011111 : 15'b000000001111111;
													assign node4606 = (inp[4]) ? 15'b000000000001111 : 15'b000000000011111;
							assign node4609 = (inp[1]) ? node4731 : node4610;
								assign node4610 = (inp[2]) ? node4670 : node4611;
									assign node4611 = (inp[14]) ? node4641 : node4612;
										assign node4612 = (inp[10]) ? node4628 : node4613;
											assign node4613 = (inp[4]) ? node4621 : node4614;
												assign node4614 = (inp[3]) ? node4618 : node4615;
													assign node4615 = (inp[11]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node4618 = (inp[0]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node4621 = (inp[11]) ? node4625 : node4622;
													assign node4622 = (inp[0]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node4625 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node4628 = (inp[3]) ? node4636 : node4629;
												assign node4629 = (inp[8]) ? node4633 : node4630;
													assign node4630 = (inp[4]) ? 15'b000000111111111 : 15'b000000111111111;
													assign node4633 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node4636 = (inp[8]) ? 15'b000000000111111 : node4637;
													assign node4637 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node4641 = (inp[3]) ? node4657 : node4642;
											assign node4642 = (inp[8]) ? node4650 : node4643;
												assign node4643 = (inp[0]) ? node4647 : node4644;
													assign node4644 = (inp[11]) ? 15'b000000111111111 : 15'b000011111111111;
													assign node4647 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node4650 = (inp[4]) ? node4654 : node4651;
													assign node4651 = (inp[10]) ? 15'b000000011111111 : 15'b000001111111111;
													assign node4654 = (inp[11]) ? 15'b000000000111111 : 15'b000000011111111;
											assign node4657 = (inp[4]) ? node4665 : node4658;
												assign node4658 = (inp[11]) ? node4662 : node4659;
													assign node4659 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node4662 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node4665 = (inp[0]) ? 15'b000000001111111 : node4666;
													assign node4666 = (inp[11]) ? 15'b000000000111111 : 15'b000000011111111;
									assign node4670 = (inp[0]) ? node4700 : node4671;
										assign node4671 = (inp[4]) ? node4685 : node4672;
											assign node4672 = (inp[3]) ? node4678 : node4673;
												assign node4673 = (inp[14]) ? 15'b000000111111111 : node4674;
													assign node4674 = (inp[8]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node4678 = (inp[10]) ? node4682 : node4679;
													assign node4679 = (inp[14]) ? 15'b000000001111111 : 15'b000000111111111;
													assign node4682 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node4685 = (inp[3]) ? node4693 : node4686;
												assign node4686 = (inp[14]) ? node4690 : node4687;
													assign node4687 = (inp[8]) ? 15'b000000011111111 : 15'b000000011111111;
													assign node4690 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node4693 = (inp[10]) ? node4697 : node4694;
													assign node4694 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node4697 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node4700 = (inp[10]) ? node4716 : node4701;
											assign node4701 = (inp[11]) ? node4709 : node4702;
												assign node4702 = (inp[14]) ? node4706 : node4703;
													assign node4703 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node4706 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node4709 = (inp[4]) ? node4713 : node4710;
													assign node4710 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node4713 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node4716 = (inp[8]) ? node4724 : node4717;
												assign node4717 = (inp[11]) ? node4721 : node4718;
													assign node4718 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node4721 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node4724 = (inp[11]) ? node4728 : node4725;
													assign node4725 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node4728 = (inp[14]) ? 15'b000000000011111 : 15'b000000000011111;
								assign node4731 = (inp[0]) ? node4787 : node4732;
									assign node4732 = (inp[11]) ? node4762 : node4733;
										assign node4733 = (inp[3]) ? node4747 : node4734;
											assign node4734 = (inp[8]) ? node4740 : node4735;
												assign node4735 = (inp[14]) ? node4737 : 15'b000000111111111;
													assign node4737 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node4740 = (inp[4]) ? node4744 : node4741;
													assign node4741 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node4744 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node4747 = (inp[14]) ? node4755 : node4748;
												assign node4748 = (inp[4]) ? node4752 : node4749;
													assign node4749 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node4752 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node4755 = (inp[4]) ? node4759 : node4756;
													assign node4756 = (inp[10]) ? 15'b000000001111111 : 15'b000000001111111;
													assign node4759 = (inp[8]) ? 15'b000000000111111 : 15'b000000011111111;
										assign node4762 = (inp[2]) ? node4776 : node4763;
											assign node4763 = (inp[4]) ? node4769 : node4764;
												assign node4764 = (inp[14]) ? node4766 : 15'b000000011111111;
													assign node4766 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node4769 = (inp[8]) ? node4773 : node4770;
													assign node4770 = (inp[14]) ? 15'b000000001111111 : 15'b000000001111111;
													assign node4773 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node4776 = (inp[14]) ? node4782 : node4777;
												assign node4777 = (inp[3]) ? node4779 : 15'b000000001111111;
													assign node4779 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node4782 = (inp[3]) ? node4784 : 15'b000000000111111;
													assign node4784 = (inp[8]) ? 15'b000000000011111 : 15'b000000000011111;
									assign node4787 = (inp[10]) ? node4817 : node4788;
										assign node4788 = (inp[14]) ? node4804 : node4789;
											assign node4789 = (inp[8]) ? node4797 : node4790;
												assign node4790 = (inp[4]) ? node4794 : node4791;
													assign node4791 = (inp[2]) ? 15'b000000011111111 : 15'b000000011111111;
													assign node4794 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node4797 = (inp[3]) ? node4801 : node4798;
													assign node4798 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node4801 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node4804 = (inp[11]) ? node4812 : node4805;
												assign node4805 = (inp[3]) ? node4809 : node4806;
													assign node4806 = (inp[8]) ? 15'b000000001111111 : 15'b000000001111111;
													assign node4809 = (inp[4]) ? 15'b000000000111111 : 15'b000000000111111;
												assign node4812 = (inp[3]) ? 15'b000000000111111 : node4813;
													assign node4813 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node4817 = (inp[4]) ? node4833 : node4818;
											assign node4818 = (inp[3]) ? node4826 : node4819;
												assign node4819 = (inp[8]) ? node4823 : node4820;
													assign node4820 = (inp[2]) ? 15'b000000001111111 : 15'b000000111111111;
													assign node4823 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node4826 = (inp[14]) ? node4830 : node4827;
													assign node4827 = (inp[2]) ? 15'b000000000111111 : 15'b000000000111111;
													assign node4830 = (inp[11]) ? 15'b000000000011111 : 15'b000000000011111;
											assign node4833 = (inp[3]) ? node4841 : node4834;
												assign node4834 = (inp[14]) ? node4838 : node4835;
													assign node4835 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node4838 = (inp[11]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node4841 = (inp[14]) ? node4845 : node4842;
													assign node4842 = (inp[2]) ? 15'b000000000011111 : 15'b000000000011111;
													assign node4845 = (inp[11]) ? 15'b000000000001111 : 15'b000000000001111;
					assign node4848 = (inp[11]) ? node5326 : node4849;
						assign node4849 = (inp[3]) ? node5083 : node4850;
							assign node4850 = (inp[2]) ? node4968 : node4851;
								assign node4851 = (inp[8]) ? node4909 : node4852;
									assign node4852 = (inp[4]) ? node4878 : node4853;
										assign node4853 = (inp[0]) ? node4869 : node4854;
											assign node4854 = (inp[9]) ? node4862 : node4855;
												assign node4855 = (inp[13]) ? node4859 : node4856;
													assign node4856 = (inp[1]) ? 15'b000011111111111 : 15'b000111111111111;
													assign node4859 = (inp[10]) ? 15'b000000111111111 : 15'b000011111111111;
												assign node4862 = (inp[1]) ? node4866 : node4863;
													assign node4863 = (inp[10]) ? 15'b000001111111111 : 15'b000001111111111;
													assign node4866 = (inp[10]) ? 15'b000001111111111 : 15'b000000111111111;
											assign node4869 = (inp[10]) ? node4871 : 15'b000001111111111;
												assign node4871 = (inp[1]) ? node4875 : node4872;
													assign node4872 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node4875 = (inp[9]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node4878 = (inp[13]) ? node4894 : node4879;
											assign node4879 = (inp[9]) ? node4887 : node4880;
												assign node4880 = (inp[0]) ? node4884 : node4881;
													assign node4881 = (inp[14]) ? 15'b000001111111111 : 15'b000001111111111;
													assign node4884 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node4887 = (inp[1]) ? node4891 : node4888;
													assign node4888 = (inp[10]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node4891 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node4894 = (inp[10]) ? node4902 : node4895;
												assign node4895 = (inp[1]) ? node4899 : node4896;
													assign node4896 = (inp[9]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node4899 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node4902 = (inp[14]) ? node4906 : node4903;
													assign node4903 = (inp[9]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node4906 = (inp[0]) ? 15'b000000001111111 : 15'b000000001111111;
									assign node4909 = (inp[13]) ? node4941 : node4910;
										assign node4910 = (inp[9]) ? node4926 : node4911;
											assign node4911 = (inp[0]) ? node4919 : node4912;
												assign node4912 = (inp[14]) ? node4916 : node4913;
													assign node4913 = (inp[4]) ? 15'b000001111111111 : 15'b000111111111111;
													assign node4916 = (inp[10]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node4919 = (inp[1]) ? node4923 : node4920;
													assign node4920 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node4923 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node4926 = (inp[14]) ? node4934 : node4927;
												assign node4927 = (inp[4]) ? node4931 : node4928;
													assign node4928 = (inp[10]) ? 15'b000000111111111 : 15'b000000111111111;
													assign node4931 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node4934 = (inp[1]) ? node4938 : node4935;
													assign node4935 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node4938 = (inp[0]) ? 15'b000000001111111 : 15'b000000001111111;
										assign node4941 = (inp[9]) ? node4955 : node4942;
											assign node4942 = (inp[14]) ? node4948 : node4943;
												assign node4943 = (inp[4]) ? 15'b000000111111111 : node4944;
													assign node4944 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node4948 = (inp[0]) ? node4952 : node4949;
													assign node4949 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node4952 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node4955 = (inp[1]) ? node4961 : node4956;
												assign node4956 = (inp[4]) ? node4958 : 15'b000000011111111;
													assign node4958 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node4961 = (inp[4]) ? node4965 : node4962;
													assign node4962 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node4965 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
								assign node4968 = (inp[0]) ? node5026 : node4969;
									assign node4969 = (inp[14]) ? node4999 : node4970;
										assign node4970 = (inp[4]) ? node4986 : node4971;
											assign node4971 = (inp[13]) ? node4979 : node4972;
												assign node4972 = (inp[10]) ? node4976 : node4973;
													assign node4973 = (inp[9]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node4976 = (inp[8]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node4979 = (inp[9]) ? node4983 : node4980;
													assign node4980 = (inp[1]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node4983 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node4986 = (inp[1]) ? node4992 : node4987;
												assign node4987 = (inp[8]) ? 15'b000000111111111 : node4988;
													assign node4988 = (inp[9]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node4992 = (inp[10]) ? node4996 : node4993;
													assign node4993 = (inp[9]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node4996 = (inp[13]) ? 15'b000000000111111 : 15'b000000011111111;
										assign node4999 = (inp[13]) ? node5015 : node5000;
											assign node5000 = (inp[1]) ? node5008 : node5001;
												assign node5001 = (inp[9]) ? node5005 : node5002;
													assign node5002 = (inp[4]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node5005 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node5008 = (inp[4]) ? node5012 : node5009;
													assign node5009 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node5012 = (inp[9]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node5015 = (inp[8]) ? node5021 : node5016;
												assign node5016 = (inp[1]) ? node5018 : 15'b000000111111111;
													assign node5018 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node5021 = (inp[10]) ? node5023 : 15'b000000001111111;
													assign node5023 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node5026 = (inp[4]) ? node5056 : node5027;
										assign node5027 = (inp[10]) ? node5041 : node5028;
											assign node5028 = (inp[13]) ? node5034 : node5029;
												assign node5029 = (inp[9]) ? 15'b000000111111111 : node5030;
													assign node5030 = (inp[1]) ? 15'b000000111111111 : 15'b000011111111111;
												assign node5034 = (inp[1]) ? node5038 : node5035;
													assign node5035 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node5038 = (inp[9]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node5041 = (inp[9]) ? node5049 : node5042;
												assign node5042 = (inp[1]) ? node5046 : node5043;
													assign node5043 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node5046 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node5049 = (inp[13]) ? node5053 : node5050;
													assign node5050 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node5053 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node5056 = (inp[10]) ? node5070 : node5057;
											assign node5057 = (inp[13]) ? node5063 : node5058;
												assign node5058 = (inp[1]) ? 15'b000000011111111 : node5059;
													assign node5059 = (inp[9]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node5063 = (inp[1]) ? node5067 : node5064;
													assign node5064 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node5067 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node5070 = (inp[1]) ? node5078 : node5071;
												assign node5071 = (inp[14]) ? node5075 : node5072;
													assign node5072 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node5075 = (inp[9]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node5078 = (inp[13]) ? 15'b000000000011111 : node5079;
													assign node5079 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
							assign node5083 = (inp[1]) ? node5205 : node5084;
								assign node5084 = (inp[9]) ? node5144 : node5085;
									assign node5085 = (inp[2]) ? node5115 : node5086;
										assign node5086 = (inp[14]) ? node5100 : node5087;
											assign node5087 = (inp[13]) ? node5093 : node5088;
												assign node5088 = (inp[0]) ? node5090 : 15'b000011111111111;
													assign node5090 = (inp[4]) ? 15'b000001111111111 : 15'b000001111111111;
												assign node5093 = (inp[0]) ? node5097 : node5094;
													assign node5094 = (inp[10]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node5097 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node5100 = (inp[10]) ? node5108 : node5101;
												assign node5101 = (inp[8]) ? node5105 : node5102;
													assign node5102 = (inp[13]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node5105 = (inp[4]) ? 15'b000000011111111 : 15'b000001111111111;
												assign node5108 = (inp[8]) ? node5112 : node5109;
													assign node5109 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node5112 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node5115 = (inp[0]) ? node5131 : node5116;
											assign node5116 = (inp[13]) ? node5124 : node5117;
												assign node5117 = (inp[10]) ? node5121 : node5118;
													assign node5118 = (inp[4]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node5121 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node5124 = (inp[4]) ? node5128 : node5125;
													assign node5125 = (inp[14]) ? 15'b000000011111111 : 15'b000001111111111;
													assign node5128 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node5131 = (inp[10]) ? node5139 : node5132;
												assign node5132 = (inp[4]) ? node5136 : node5133;
													assign node5133 = (inp[14]) ? 15'b000000011111111 : 15'b000000011111111;
													assign node5136 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node5139 = (inp[13]) ? 15'b000000001111111 : node5140;
													assign node5140 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node5144 = (inp[13]) ? node5176 : node5145;
										assign node5145 = (inp[14]) ? node5161 : node5146;
											assign node5146 = (inp[10]) ? node5154 : node5147;
												assign node5147 = (inp[8]) ? node5151 : node5148;
													assign node5148 = (inp[0]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node5151 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node5154 = (inp[0]) ? node5158 : node5155;
													assign node5155 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node5158 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node5161 = (inp[4]) ? node5169 : node5162;
												assign node5162 = (inp[8]) ? node5166 : node5163;
													assign node5163 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node5166 = (inp[0]) ? 15'b000000000111111 : 15'b000000011111111;
												assign node5169 = (inp[2]) ? node5173 : node5170;
													assign node5170 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node5173 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node5176 = (inp[8]) ? node5190 : node5177;
											assign node5177 = (inp[14]) ? node5185 : node5178;
												assign node5178 = (inp[10]) ? node5182 : node5179;
													assign node5179 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node5182 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node5185 = (inp[4]) ? node5187 : 15'b000000001111111;
													assign node5187 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node5190 = (inp[2]) ? node5198 : node5191;
												assign node5191 = (inp[0]) ? node5195 : node5192;
													assign node5192 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node5195 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node5198 = (inp[14]) ? node5202 : node5199;
													assign node5199 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node5202 = (inp[10]) ? 15'b000000000011111 : 15'b000000000111111;
								assign node5205 = (inp[9]) ? node5267 : node5206;
									assign node5206 = (inp[14]) ? node5236 : node5207;
										assign node5207 = (inp[8]) ? node5221 : node5208;
											assign node5208 = (inp[13]) ? node5214 : node5209;
												assign node5209 = (inp[2]) ? 15'b000000111111111 : node5210;
													assign node5210 = (inp[10]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node5214 = (inp[0]) ? node5218 : node5215;
													assign node5215 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node5218 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node5221 = (inp[13]) ? node5229 : node5222;
												assign node5222 = (inp[2]) ? node5226 : node5223;
													assign node5223 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node5226 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node5229 = (inp[4]) ? node5233 : node5230;
													assign node5230 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node5233 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node5236 = (inp[10]) ? node5252 : node5237;
											assign node5237 = (inp[4]) ? node5245 : node5238;
												assign node5238 = (inp[8]) ? node5242 : node5239;
													assign node5239 = (inp[0]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node5242 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node5245 = (inp[8]) ? node5249 : node5246;
													assign node5246 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node5249 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node5252 = (inp[0]) ? node5260 : node5253;
												assign node5253 = (inp[2]) ? node5257 : node5254;
													assign node5254 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node5257 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node5260 = (inp[8]) ? node5264 : node5261;
													assign node5261 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node5264 = (inp[4]) ? 15'b000000000011111 : 15'b000000000011111;
									assign node5267 = (inp[14]) ? node5297 : node5268;
										assign node5268 = (inp[0]) ? node5284 : node5269;
											assign node5269 = (inp[10]) ? node5277 : node5270;
												assign node5270 = (inp[2]) ? node5274 : node5271;
													assign node5271 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node5274 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node5277 = (inp[4]) ? node5281 : node5278;
													assign node5278 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node5281 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node5284 = (inp[8]) ? node5292 : node5285;
												assign node5285 = (inp[13]) ? node5289 : node5286;
													assign node5286 = (inp[4]) ? 15'b000000001111111 : 15'b000000001111111;
													assign node5289 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node5292 = (inp[2]) ? 15'b000000000011111 : node5293;
													assign node5293 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node5297 = (inp[4]) ? node5311 : node5298;
											assign node5298 = (inp[13]) ? node5304 : node5299;
												assign node5299 = (inp[10]) ? 15'b000000001111111 : node5300;
													assign node5300 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node5304 = (inp[8]) ? node5308 : node5305;
													assign node5305 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node5308 = (inp[2]) ? 15'b000000000001111 : 15'b000000000111111;
											assign node5311 = (inp[10]) ? node5319 : node5312;
												assign node5312 = (inp[8]) ? node5316 : node5313;
													assign node5313 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node5316 = (inp[0]) ? 15'b000000000011111 : 15'b000000000011111;
												assign node5319 = (inp[2]) ? node5323 : node5320;
													assign node5320 = (inp[8]) ? 15'b000000000011111 : 15'b000000000011111;
													assign node5323 = (inp[13]) ? 15'b000000000001111 : 15'b000000000011111;
						assign node5326 = (inp[0]) ? node5572 : node5327;
							assign node5327 = (inp[10]) ? node5447 : node5328;
								assign node5328 = (inp[1]) ? node5388 : node5329;
									assign node5329 = (inp[8]) ? node5359 : node5330;
										assign node5330 = (inp[14]) ? node5346 : node5331;
											assign node5331 = (inp[9]) ? node5339 : node5332;
												assign node5332 = (inp[3]) ? node5336 : node5333;
													assign node5333 = (inp[13]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node5336 = (inp[13]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node5339 = (inp[3]) ? node5343 : node5340;
													assign node5340 = (inp[4]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node5343 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node5346 = (inp[4]) ? node5354 : node5347;
												assign node5347 = (inp[13]) ? node5351 : node5348;
													assign node5348 = (inp[3]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node5351 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node5354 = (inp[2]) ? node5356 : 15'b000000011111111;
													assign node5356 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node5359 = (inp[13]) ? node5373 : node5360;
											assign node5360 = (inp[4]) ? node5368 : node5361;
												assign node5361 = (inp[9]) ? node5365 : node5362;
													assign node5362 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node5365 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node5368 = (inp[3]) ? node5370 : 15'b000000111111111;
													assign node5370 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node5373 = (inp[2]) ? node5381 : node5374;
												assign node5374 = (inp[3]) ? node5378 : node5375;
													assign node5375 = (inp[9]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node5378 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node5381 = (inp[9]) ? node5385 : node5382;
													assign node5382 = (inp[4]) ? 15'b000000001111111 : 15'b000000001111111;
													assign node5385 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node5388 = (inp[9]) ? node5416 : node5389;
										assign node5389 = (inp[14]) ? node5405 : node5390;
											assign node5390 = (inp[3]) ? node5398 : node5391;
												assign node5391 = (inp[13]) ? node5395 : node5392;
													assign node5392 = (inp[8]) ? 15'b000000111111111 : 15'b000000111111111;
													assign node5395 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node5398 = (inp[13]) ? node5402 : node5399;
													assign node5399 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node5402 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node5405 = (inp[4]) ? node5413 : node5406;
												assign node5406 = (inp[3]) ? node5410 : node5407;
													assign node5407 = (inp[2]) ? 15'b000000011111111 : 15'b000000011111111;
													assign node5410 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node5413 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node5416 = (inp[13]) ? node5432 : node5417;
											assign node5417 = (inp[3]) ? node5425 : node5418;
												assign node5418 = (inp[8]) ? node5422 : node5419;
													assign node5419 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node5422 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node5425 = (inp[4]) ? node5429 : node5426;
													assign node5426 = (inp[8]) ? 15'b000000001111111 : 15'b000000001111111;
													assign node5429 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node5432 = (inp[2]) ? node5440 : node5433;
												assign node5433 = (inp[8]) ? node5437 : node5434;
													assign node5434 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node5437 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node5440 = (inp[4]) ? node5444 : node5441;
													assign node5441 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node5444 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
								assign node5447 = (inp[4]) ? node5509 : node5448;
									assign node5448 = (inp[3]) ? node5478 : node5449;
										assign node5449 = (inp[8]) ? node5463 : node5450;
											assign node5450 = (inp[9]) ? node5458 : node5451;
												assign node5451 = (inp[1]) ? node5455 : node5452;
													assign node5452 = (inp[2]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node5455 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node5458 = (inp[13]) ? 15'b000000011111111 : node5459;
													assign node5459 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node5463 = (inp[2]) ? node5471 : node5464;
												assign node5464 = (inp[9]) ? node5468 : node5465;
													assign node5465 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node5468 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node5471 = (inp[1]) ? node5475 : node5472;
													assign node5472 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node5475 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node5478 = (inp[1]) ? node5494 : node5479;
											assign node5479 = (inp[14]) ? node5487 : node5480;
												assign node5480 = (inp[2]) ? node5484 : node5481;
													assign node5481 = (inp[9]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node5484 = (inp[9]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node5487 = (inp[13]) ? node5491 : node5488;
													assign node5488 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node5491 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node5494 = (inp[13]) ? node5502 : node5495;
												assign node5495 = (inp[14]) ? node5499 : node5496;
													assign node5496 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node5499 = (inp[2]) ? 15'b000000000111111 : 15'b000000000111111;
												assign node5502 = (inp[8]) ? node5506 : node5503;
													assign node5503 = (inp[14]) ? 15'b000000000111111 : 15'b000000000111111;
													assign node5506 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node5509 = (inp[9]) ? node5541 : node5510;
										assign node5510 = (inp[13]) ? node5526 : node5511;
											assign node5511 = (inp[2]) ? node5519 : node5512;
												assign node5512 = (inp[14]) ? node5516 : node5513;
													assign node5513 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node5516 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node5519 = (inp[14]) ? node5523 : node5520;
													assign node5520 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node5523 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node5526 = (inp[3]) ? node5534 : node5527;
												assign node5527 = (inp[8]) ? node5531 : node5528;
													assign node5528 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node5531 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node5534 = (inp[14]) ? node5538 : node5535;
													assign node5535 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node5538 = (inp[1]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node5541 = (inp[2]) ? node5557 : node5542;
											assign node5542 = (inp[3]) ? node5550 : node5543;
												assign node5543 = (inp[14]) ? node5547 : node5544;
													assign node5544 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node5547 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node5550 = (inp[8]) ? node5554 : node5551;
													assign node5551 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node5554 = (inp[1]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node5557 = (inp[14]) ? node5565 : node5558;
												assign node5558 = (inp[1]) ? node5562 : node5559;
													assign node5559 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node5562 = (inp[3]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node5565 = (inp[8]) ? node5569 : node5566;
													assign node5566 = (inp[13]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node5569 = (inp[1]) ? 15'b000000000001111 : 15'b000000000111111;
							assign node5572 = (inp[1]) ? node5686 : node5573;
								assign node5573 = (inp[3]) ? node5629 : node5574;
									assign node5574 = (inp[4]) ? node5600 : node5575;
										assign node5575 = (inp[10]) ? node5585 : node5576;
											assign node5576 = (inp[9]) ? node5582 : node5577;
												assign node5577 = (inp[13]) ? 15'b000000111111111 : node5578;
													assign node5578 = (inp[8]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node5582 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node5585 = (inp[14]) ? node5593 : node5586;
												assign node5586 = (inp[8]) ? node5590 : node5587;
													assign node5587 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node5590 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node5593 = (inp[13]) ? node5597 : node5594;
													assign node5594 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node5597 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node5600 = (inp[2]) ? node5616 : node5601;
											assign node5601 = (inp[14]) ? node5609 : node5602;
												assign node5602 = (inp[13]) ? node5606 : node5603;
													assign node5603 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node5606 = (inp[9]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node5609 = (inp[9]) ? node5613 : node5610;
													assign node5610 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node5613 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node5616 = (inp[8]) ? node5624 : node5617;
												assign node5617 = (inp[13]) ? node5621 : node5618;
													assign node5618 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node5621 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node5624 = (inp[14]) ? 15'b000000000011111 : node5625;
													assign node5625 = (inp[13]) ? 15'b000000000011111 : 15'b000000001111111;
									assign node5629 = (inp[13]) ? node5657 : node5630;
										assign node5630 = (inp[2]) ? node5644 : node5631;
											assign node5631 = (inp[4]) ? node5639 : node5632;
												assign node5632 = (inp[14]) ? node5636 : node5633;
													assign node5633 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node5636 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node5639 = (inp[9]) ? 15'b000000000111111 : node5640;
													assign node5640 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node5644 = (inp[14]) ? node5652 : node5645;
												assign node5645 = (inp[9]) ? node5649 : node5646;
													assign node5646 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node5649 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node5652 = (inp[9]) ? 15'b000000000011111 : node5653;
													assign node5653 = (inp[10]) ? 15'b000000000111111 : 15'b000000000111111;
										assign node5657 = (inp[4]) ? node5673 : node5658;
											assign node5658 = (inp[8]) ? node5666 : node5659;
												assign node5659 = (inp[2]) ? node5663 : node5660;
													assign node5660 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node5663 = (inp[10]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node5666 = (inp[10]) ? node5670 : node5667;
													assign node5667 = (inp[14]) ? 15'b000000000011111 : 15'b000000001111111;
													assign node5670 = (inp[9]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node5673 = (inp[14]) ? node5681 : node5674;
												assign node5674 = (inp[8]) ? node5678 : node5675;
													assign node5675 = (inp[9]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node5678 = (inp[2]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node5681 = (inp[2]) ? node5683 : 15'b000000000011111;
													assign node5683 = (inp[10]) ? 15'b000000000001111 : 15'b000000000011111;
								assign node5686 = (inp[9]) ? node5746 : node5687;
									assign node5687 = (inp[13]) ? node5717 : node5688;
										assign node5688 = (inp[3]) ? node5702 : node5689;
											assign node5689 = (inp[2]) ? node5695 : node5690;
												assign node5690 = (inp[4]) ? node5692 : 15'b000000011111111;
													assign node5692 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node5695 = (inp[10]) ? node5699 : node5696;
													assign node5696 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node5699 = (inp[14]) ? 15'b000000000111111 : 15'b000000000111111;
											assign node5702 = (inp[4]) ? node5710 : node5703;
												assign node5703 = (inp[2]) ? node5707 : node5704;
													assign node5704 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node5707 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node5710 = (inp[10]) ? node5714 : node5711;
													assign node5711 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node5714 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node5717 = (inp[10]) ? node5733 : node5718;
											assign node5718 = (inp[8]) ? node5726 : node5719;
												assign node5719 = (inp[2]) ? node5723 : node5720;
													assign node5720 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node5723 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node5726 = (inp[14]) ? node5730 : node5727;
													assign node5727 = (inp[2]) ? 15'b000000000011111 : 15'b000000001111111;
													assign node5730 = (inp[3]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node5733 = (inp[3]) ? node5741 : node5734;
												assign node5734 = (inp[8]) ? node5738 : node5735;
													assign node5735 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node5738 = (inp[2]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node5741 = (inp[14]) ? node5743 : 15'b000000000011111;
													assign node5743 = (inp[8]) ? 15'b000000000001111 : 15'b000000000011111;
									assign node5746 = (inp[8]) ? node5778 : node5747;
										assign node5747 = (inp[2]) ? node5763 : node5748;
											assign node5748 = (inp[14]) ? node5756 : node5749;
												assign node5749 = (inp[10]) ? node5753 : node5750;
													assign node5750 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node5753 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node5756 = (inp[4]) ? node5760 : node5757;
													assign node5757 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node5760 = (inp[3]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node5763 = (inp[10]) ? node5771 : node5764;
												assign node5764 = (inp[14]) ? node5768 : node5765;
													assign node5765 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node5768 = (inp[4]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node5771 = (inp[13]) ? node5775 : node5772;
													assign node5772 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node5775 = (inp[14]) ? 15'b000000000000111 : 15'b000000000001111;
										assign node5778 = (inp[4]) ? node5794 : node5779;
											assign node5779 = (inp[13]) ? node5787 : node5780;
												assign node5780 = (inp[14]) ? node5784 : node5781;
													assign node5781 = (inp[2]) ? 15'b000000000111111 : 15'b000000000111111;
													assign node5784 = (inp[10]) ? 15'b000000000001111 : 15'b000000000111111;
												assign node5787 = (inp[2]) ? node5791 : node5788;
													assign node5788 = (inp[3]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node5791 = (inp[14]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node5794 = (inp[3]) ? node5802 : node5795;
												assign node5795 = (inp[10]) ? node5799 : node5796;
													assign node5796 = (inp[14]) ? 15'b000000000011111 : 15'b000000000011111;
													assign node5799 = (inp[14]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node5802 = (inp[13]) ? node5806 : node5803;
													assign node5803 = (inp[10]) ? 15'b000000000001111 : 15'b000000000011111;
													assign node5806 = (inp[2]) ? 15'b000000000000111 : 15'b000000000001111;
				assign node5809 = (inp[13]) ? node6767 : node5810;
					assign node5810 = (inp[14]) ? node6286 : node5811;
						assign node5811 = (inp[9]) ? node6055 : node5812;
							assign node5812 = (inp[8]) ? node5934 : node5813;
								assign node5813 = (inp[3]) ? node5873 : node5814;
									assign node5814 = (inp[10]) ? node5844 : node5815;
										assign node5815 = (inp[11]) ? node5831 : node5816;
											assign node5816 = (inp[1]) ? node5824 : node5817;
												assign node5817 = (inp[4]) ? node5821 : node5818;
													assign node5818 = (inp[2]) ? 15'b000011111111111 : 15'b000111111111111;
													assign node5821 = (inp[12]) ? 15'b000001111111111 : 15'b000001111111111;
												assign node5824 = (inp[12]) ? node5828 : node5825;
													assign node5825 = (inp[2]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node5828 = (inp[4]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node5831 = (inp[0]) ? node5837 : node5832;
												assign node5832 = (inp[12]) ? 15'b000000111111111 : node5833;
													assign node5833 = (inp[1]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node5837 = (inp[4]) ? node5841 : node5838;
													assign node5838 = (inp[2]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node5841 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node5844 = (inp[1]) ? node5858 : node5845;
											assign node5845 = (inp[11]) ? node5851 : node5846;
												assign node5846 = (inp[0]) ? node5848 : 15'b000001111111111;
													assign node5848 = (inp[12]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node5851 = (inp[0]) ? node5855 : node5852;
													assign node5852 = (inp[12]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node5855 = (inp[12]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node5858 = (inp[11]) ? node5866 : node5859;
												assign node5859 = (inp[4]) ? node5863 : node5860;
													assign node5860 = (inp[2]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node5863 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node5866 = (inp[2]) ? node5870 : node5867;
													assign node5867 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node5870 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node5873 = (inp[2]) ? node5905 : node5874;
										assign node5874 = (inp[1]) ? node5890 : node5875;
											assign node5875 = (inp[12]) ? node5883 : node5876;
												assign node5876 = (inp[10]) ? node5880 : node5877;
													assign node5877 = (inp[4]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node5880 = (inp[0]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node5883 = (inp[11]) ? node5887 : node5884;
													assign node5884 = (inp[0]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node5887 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node5890 = (inp[4]) ? node5898 : node5891;
												assign node5891 = (inp[0]) ? node5895 : node5892;
													assign node5892 = (inp[11]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node5895 = (inp[11]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node5898 = (inp[11]) ? node5902 : node5899;
													assign node5899 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node5902 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node5905 = (inp[12]) ? node5919 : node5906;
											assign node5906 = (inp[1]) ? node5914 : node5907;
												assign node5907 = (inp[0]) ? node5911 : node5908;
													assign node5908 = (inp[11]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node5911 = (inp[10]) ? 15'b000000001111111 : 15'b000000111111111;
												assign node5914 = (inp[0]) ? 15'b000000011111111 : node5915;
													assign node5915 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node5919 = (inp[10]) ? node5927 : node5920;
												assign node5920 = (inp[11]) ? node5924 : node5921;
													assign node5921 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node5924 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node5927 = (inp[11]) ? node5931 : node5928;
													assign node5928 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node5931 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
								assign node5934 = (inp[0]) ? node5992 : node5935;
									assign node5935 = (inp[12]) ? node5963 : node5936;
										assign node5936 = (inp[11]) ? node5950 : node5937;
											assign node5937 = (inp[10]) ? node5945 : node5938;
												assign node5938 = (inp[3]) ? node5942 : node5939;
													assign node5939 = (inp[1]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node5942 = (inp[2]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node5945 = (inp[2]) ? 15'b000000111111111 : node5946;
													assign node5946 = (inp[4]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node5950 = (inp[2]) ? node5958 : node5951;
												assign node5951 = (inp[3]) ? node5955 : node5952;
													assign node5952 = (inp[1]) ? 15'b000000111111111 : 15'b000000111111111;
													assign node5955 = (inp[10]) ? 15'b000000111111111 : 15'b000000011111111;
												assign node5958 = (inp[3]) ? 15'b000000001111111 : node5959;
													assign node5959 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node5963 = (inp[4]) ? node5977 : node5964;
											assign node5964 = (inp[1]) ? node5972 : node5965;
												assign node5965 = (inp[3]) ? node5969 : node5966;
													assign node5966 = (inp[10]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node5969 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node5972 = (inp[2]) ? 15'b000000011111111 : node5973;
													assign node5973 = (inp[11]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node5977 = (inp[1]) ? node5985 : node5978;
												assign node5978 = (inp[3]) ? node5982 : node5979;
													assign node5979 = (inp[11]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node5982 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node5985 = (inp[2]) ? node5989 : node5986;
													assign node5986 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node5989 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node5992 = (inp[11]) ? node6024 : node5993;
										assign node5993 = (inp[2]) ? node6009 : node5994;
											assign node5994 = (inp[10]) ? node6002 : node5995;
												assign node5995 = (inp[4]) ? node5999 : node5996;
													assign node5996 = (inp[12]) ? 15'b000000111111111 : 15'b000000111111111;
													assign node5999 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node6002 = (inp[3]) ? node6006 : node6003;
													assign node6003 = (inp[12]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node6006 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node6009 = (inp[1]) ? node6017 : node6010;
												assign node6010 = (inp[12]) ? node6014 : node6011;
													assign node6011 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node6014 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node6017 = (inp[10]) ? node6021 : node6018;
													assign node6018 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node6021 = (inp[12]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node6024 = (inp[4]) ? node6040 : node6025;
											assign node6025 = (inp[1]) ? node6033 : node6026;
												assign node6026 = (inp[12]) ? node6030 : node6027;
													assign node6027 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node6030 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node6033 = (inp[10]) ? node6037 : node6034;
													assign node6034 = (inp[12]) ? 15'b000000000111111 : 15'b000000011111111;
													assign node6037 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node6040 = (inp[12]) ? node6048 : node6041;
												assign node6041 = (inp[1]) ? node6045 : node6042;
													assign node6042 = (inp[10]) ? 15'b000000001111111 : 15'b000000001111111;
													assign node6045 = (inp[2]) ? 15'b000000000011111 : 15'b000000001111111;
												assign node6048 = (inp[3]) ? node6052 : node6049;
													assign node6049 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node6052 = (inp[1]) ? 15'b000000000001111 : 15'b000000000111111;
							assign node6055 = (inp[11]) ? node6171 : node6056;
								assign node6056 = (inp[12]) ? node6112 : node6057;
									assign node6057 = (inp[3]) ? node6087 : node6058;
										assign node6058 = (inp[8]) ? node6072 : node6059;
											assign node6059 = (inp[1]) ? node6067 : node6060;
												assign node6060 = (inp[0]) ? node6064 : node6061;
													assign node6061 = (inp[10]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node6064 = (inp[2]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node6067 = (inp[4]) ? 15'b000000111111111 : node6068;
													assign node6068 = (inp[2]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node6072 = (inp[1]) ? node6080 : node6073;
												assign node6073 = (inp[10]) ? node6077 : node6074;
													assign node6074 = (inp[0]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node6077 = (inp[4]) ? 15'b000000011111111 : 15'b000000011111111;
												assign node6080 = (inp[2]) ? node6084 : node6081;
													assign node6081 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node6084 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node6087 = (inp[4]) ? node6103 : node6088;
											assign node6088 = (inp[0]) ? node6096 : node6089;
												assign node6089 = (inp[10]) ? node6093 : node6090;
													assign node6090 = (inp[2]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node6093 = (inp[2]) ? 15'b000000001111111 : 15'b000000111111111;
												assign node6096 = (inp[2]) ? node6100 : node6097;
													assign node6097 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node6100 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node6103 = (inp[2]) ? node6107 : node6104;
												assign node6104 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node6107 = (inp[1]) ? node6109 : 15'b000000001111111;
													assign node6109 = (inp[0]) ? 15'b000000000111111 : 15'b000000000111111;
									assign node6112 = (inp[0]) ? node6140 : node6113;
										assign node6113 = (inp[1]) ? node6127 : node6114;
											assign node6114 = (inp[10]) ? node6120 : node6115;
												assign node6115 = (inp[4]) ? 15'b000000111111111 : node6116;
													assign node6116 = (inp[8]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node6120 = (inp[8]) ? node6124 : node6121;
													assign node6121 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node6124 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node6127 = (inp[2]) ? node6135 : node6128;
												assign node6128 = (inp[10]) ? node6132 : node6129;
													assign node6129 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node6132 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node6135 = (inp[3]) ? 15'b000000001111111 : node6136;
													assign node6136 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node6140 = (inp[8]) ? node6156 : node6141;
											assign node6141 = (inp[1]) ? node6149 : node6142;
												assign node6142 = (inp[10]) ? node6146 : node6143;
													assign node6143 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node6146 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node6149 = (inp[4]) ? node6153 : node6150;
													assign node6150 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node6153 = (inp[2]) ? 15'b000000000011111 : 15'b000000001111111;
											assign node6156 = (inp[4]) ? node6164 : node6157;
												assign node6157 = (inp[10]) ? node6161 : node6158;
													assign node6158 = (inp[1]) ? 15'b000000001111111 : 15'b000000001111111;
													assign node6161 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node6164 = (inp[2]) ? node6168 : node6165;
													assign node6165 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node6168 = (inp[3]) ? 15'b000000000011111 : 15'b000000000111111;
								assign node6171 = (inp[10]) ? node6229 : node6172;
									assign node6172 = (inp[1]) ? node6198 : node6173;
										assign node6173 = (inp[0]) ? node6185 : node6174;
											assign node6174 = (inp[4]) ? node6182 : node6175;
												assign node6175 = (inp[8]) ? node6179 : node6176;
													assign node6176 = (inp[3]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node6179 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node6182 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node6185 = (inp[12]) ? node6191 : node6186;
												assign node6186 = (inp[3]) ? node6188 : 15'b000000111111111;
													assign node6188 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node6191 = (inp[3]) ? node6195 : node6192;
													assign node6192 = (inp[2]) ? 15'b000000001111111 : 15'b000000001111111;
													assign node6195 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node6198 = (inp[4]) ? node6214 : node6199;
											assign node6199 = (inp[2]) ? node6207 : node6200;
												assign node6200 = (inp[12]) ? node6204 : node6201;
													assign node6201 = (inp[3]) ? 15'b000000011111111 : 15'b000000011111111;
													assign node6204 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node6207 = (inp[8]) ? node6211 : node6208;
													assign node6208 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node6211 = (inp[12]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node6214 = (inp[3]) ? node6222 : node6215;
												assign node6215 = (inp[0]) ? node6219 : node6216;
													assign node6216 = (inp[2]) ? 15'b000000001111111 : 15'b000000001111111;
													assign node6219 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node6222 = (inp[0]) ? node6226 : node6223;
													assign node6223 = (inp[8]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node6226 = (inp[12]) ? 15'b000000000111111 : 15'b000000000111111;
									assign node6229 = (inp[12]) ? node6261 : node6230;
										assign node6230 = (inp[8]) ? node6246 : node6231;
											assign node6231 = (inp[3]) ? node6239 : node6232;
												assign node6232 = (inp[0]) ? node6236 : node6233;
													assign node6233 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node6236 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node6239 = (inp[2]) ? node6243 : node6240;
													assign node6240 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node6243 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node6246 = (inp[2]) ? node6254 : node6247;
												assign node6247 = (inp[1]) ? node6251 : node6248;
													assign node6248 = (inp[4]) ? 15'b000000001111111 : 15'b000000111111111;
													assign node6251 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node6254 = (inp[0]) ? node6258 : node6255;
													assign node6255 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node6258 = (inp[1]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node6261 = (inp[8]) ? node6273 : node6262;
											assign node6262 = (inp[1]) ? node6266 : node6263;
												assign node6263 = (inp[3]) ? 15'b000000011111111 : 15'b000000001111111;
												assign node6266 = (inp[3]) ? node6270 : node6267;
													assign node6267 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node6270 = (inp[2]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node6273 = (inp[1]) ? node6281 : node6274;
												assign node6274 = (inp[3]) ? node6278 : node6275;
													assign node6275 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node6278 = (inp[4]) ? 15'b000000000011111 : 15'b000000000011111;
												assign node6281 = (inp[2]) ? node6283 : 15'b000000000011111;
													assign node6283 = (inp[0]) ? 15'b000000000001111 : 15'b000000000011111;
						assign node6286 = (inp[12]) ? node6534 : node6287;
							assign node6287 = (inp[0]) ? node6409 : node6288;
								assign node6288 = (inp[9]) ? node6350 : node6289;
									assign node6289 = (inp[1]) ? node6321 : node6290;
										assign node6290 = (inp[4]) ? node6306 : node6291;
											assign node6291 = (inp[3]) ? node6299 : node6292;
												assign node6292 = (inp[8]) ? node6296 : node6293;
													assign node6293 = (inp[2]) ? 15'b000011111111111 : 15'b000011111111111;
													assign node6296 = (inp[10]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node6299 = (inp[8]) ? node6303 : node6300;
													assign node6300 = (inp[10]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node6303 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node6306 = (inp[11]) ? node6314 : node6307;
												assign node6307 = (inp[2]) ? node6311 : node6308;
													assign node6308 = (inp[8]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node6311 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node6314 = (inp[8]) ? node6318 : node6315;
													assign node6315 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node6318 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node6321 = (inp[3]) ? node6337 : node6322;
											assign node6322 = (inp[11]) ? node6330 : node6323;
												assign node6323 = (inp[2]) ? node6327 : node6324;
													assign node6324 = (inp[8]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node6327 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node6330 = (inp[10]) ? node6334 : node6331;
													assign node6331 = (inp[4]) ? 15'b000000011111111 : 15'b000000011111111;
													assign node6334 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node6337 = (inp[8]) ? node6345 : node6338;
												assign node6338 = (inp[11]) ? node6342 : node6339;
													assign node6339 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node6342 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node6345 = (inp[10]) ? 15'b000000001111111 : node6346;
													assign node6346 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node6350 = (inp[11]) ? node6380 : node6351;
										assign node6351 = (inp[4]) ? node6365 : node6352;
											assign node6352 = (inp[1]) ? node6358 : node6353;
												assign node6353 = (inp[8]) ? 15'b000000011111111 : node6354;
													assign node6354 = (inp[2]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node6358 = (inp[2]) ? node6362 : node6359;
													assign node6359 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node6362 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node6365 = (inp[3]) ? node6373 : node6366;
												assign node6366 = (inp[8]) ? node6370 : node6367;
													assign node6367 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node6370 = (inp[2]) ? 15'b000000001111111 : 15'b000000001111111;
												assign node6373 = (inp[1]) ? node6377 : node6374;
													assign node6374 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node6377 = (inp[8]) ? 15'b000000000111111 : 15'b000000000111111;
										assign node6380 = (inp[4]) ? node6396 : node6381;
											assign node6381 = (inp[3]) ? node6389 : node6382;
												assign node6382 = (inp[1]) ? node6386 : node6383;
													assign node6383 = (inp[8]) ? 15'b000000001111111 : 15'b000000111111111;
													assign node6386 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node6389 = (inp[2]) ? node6393 : node6390;
													assign node6390 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node6393 = (inp[8]) ? 15'b000000000111111 : 15'b000000000111111;
											assign node6396 = (inp[10]) ? node6402 : node6397;
												assign node6397 = (inp[2]) ? node6399 : 15'b000000011111111;
													assign node6399 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node6402 = (inp[2]) ? node6406 : node6403;
													assign node6403 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node6406 = (inp[1]) ? 15'b000000000001111 : 15'b000000000111111;
								assign node6409 = (inp[3]) ? node6471 : node6410;
									assign node6410 = (inp[10]) ? node6442 : node6411;
										assign node6411 = (inp[1]) ? node6427 : node6412;
											assign node6412 = (inp[8]) ? node6420 : node6413;
												assign node6413 = (inp[4]) ? node6417 : node6414;
													assign node6414 = (inp[2]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node6417 = (inp[9]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node6420 = (inp[11]) ? node6424 : node6421;
													assign node6421 = (inp[9]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node6424 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node6427 = (inp[11]) ? node6435 : node6428;
												assign node6428 = (inp[9]) ? node6432 : node6429;
													assign node6429 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node6432 = (inp[8]) ? 15'b000000001111111 : 15'b000000001111111;
												assign node6435 = (inp[4]) ? node6439 : node6436;
													assign node6436 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node6439 = (inp[9]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node6442 = (inp[9]) ? node6456 : node6443;
											assign node6443 = (inp[8]) ? node6449 : node6444;
												assign node6444 = (inp[2]) ? node6446 : 15'b000001111111111;
													assign node6446 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node6449 = (inp[1]) ? node6453 : node6450;
													assign node6450 = (inp[2]) ? 15'b000000001111111 : 15'b000000001111111;
													assign node6453 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node6456 = (inp[2]) ? node6464 : node6457;
												assign node6457 = (inp[4]) ? node6461 : node6458;
													assign node6458 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node6461 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node6464 = (inp[4]) ? node6468 : node6465;
													assign node6465 = (inp[11]) ? 15'b000000000011111 : 15'b000000001111111;
													assign node6468 = (inp[1]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node6471 = (inp[11]) ? node6503 : node6472;
										assign node6472 = (inp[2]) ? node6488 : node6473;
											assign node6473 = (inp[10]) ? node6481 : node6474;
												assign node6474 = (inp[9]) ? node6478 : node6475;
													assign node6475 = (inp[1]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node6478 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node6481 = (inp[1]) ? node6485 : node6482;
													assign node6482 = (inp[9]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node6485 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node6488 = (inp[4]) ? node6496 : node6489;
												assign node6489 = (inp[1]) ? node6493 : node6490;
													assign node6490 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node6493 = (inp[8]) ? 15'b000000000011111 : 15'b000000001111111;
												assign node6496 = (inp[9]) ? node6500 : node6497;
													assign node6497 = (inp[10]) ? 15'b000000000011111 : 15'b000000011111111;
													assign node6500 = (inp[10]) ? 15'b000000000011111 : 15'b000000000011111;
										assign node6503 = (inp[10]) ? node6519 : node6504;
											assign node6504 = (inp[1]) ? node6512 : node6505;
												assign node6505 = (inp[4]) ? node6509 : node6506;
													assign node6506 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node6509 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node6512 = (inp[4]) ? node6516 : node6513;
													assign node6513 = (inp[8]) ? 15'b000000000111111 : 15'b000000000111111;
													assign node6516 = (inp[2]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node6519 = (inp[4]) ? node6527 : node6520;
												assign node6520 = (inp[9]) ? node6524 : node6521;
													assign node6521 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node6524 = (inp[2]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node6527 = (inp[9]) ? node6531 : node6528;
													assign node6528 = (inp[8]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node6531 = (inp[8]) ? 15'b000000000001111 : 15'b000000000011111;
							assign node6534 = (inp[8]) ? node6648 : node6535;
								assign node6535 = (inp[2]) ? node6591 : node6536;
									assign node6536 = (inp[9]) ? node6566 : node6537;
										assign node6537 = (inp[1]) ? node6551 : node6538;
											assign node6538 = (inp[11]) ? node6544 : node6539;
												assign node6539 = (inp[10]) ? node6541 : 15'b000001111111111;
													assign node6541 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node6544 = (inp[10]) ? node6548 : node6545;
													assign node6545 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node6548 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node6551 = (inp[11]) ? node6559 : node6552;
												assign node6552 = (inp[10]) ? node6556 : node6553;
													assign node6553 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node6556 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node6559 = (inp[3]) ? node6563 : node6560;
													assign node6560 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node6563 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node6566 = (inp[1]) ? node6578 : node6567;
											assign node6567 = (inp[0]) ? node6573 : node6568;
												assign node6568 = (inp[11]) ? node6570 : 15'b000000111111111;
													assign node6570 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node6573 = (inp[4]) ? node6575 : 15'b000000001111111;
													assign node6575 = (inp[11]) ? 15'b000000000111111 : 15'b000000000111111;
											assign node6578 = (inp[3]) ? node6584 : node6579;
												assign node6579 = (inp[11]) ? node6581 : 15'b000000001111111;
													assign node6581 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node6584 = (inp[11]) ? node6588 : node6585;
													assign node6585 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node6588 = (inp[0]) ? 15'b000000000011111 : 15'b000000000011111;
									assign node6591 = (inp[9]) ? node6621 : node6592;
										assign node6592 = (inp[11]) ? node6606 : node6593;
											assign node6593 = (inp[1]) ? node6601 : node6594;
												assign node6594 = (inp[3]) ? node6598 : node6595;
													assign node6595 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node6598 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node6601 = (inp[3]) ? node6603 : 15'b000000001111111;
													assign node6603 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node6606 = (inp[3]) ? node6614 : node6607;
												assign node6607 = (inp[4]) ? node6611 : node6608;
													assign node6608 = (inp[0]) ? 15'b000000001111111 : 15'b000000001111111;
													assign node6611 = (inp[10]) ? 15'b000000000011111 : 15'b000000001111111;
												assign node6614 = (inp[10]) ? node6618 : node6615;
													assign node6615 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node6618 = (inp[0]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node6621 = (inp[0]) ? node6635 : node6622;
											assign node6622 = (inp[11]) ? node6628 : node6623;
												assign node6623 = (inp[1]) ? node6625 : 15'b000000011111111;
													assign node6625 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node6628 = (inp[3]) ? node6632 : node6629;
													assign node6629 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node6632 = (inp[10]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node6635 = (inp[10]) ? node6641 : node6636;
												assign node6636 = (inp[1]) ? node6638 : 15'b000000001111111;
													assign node6638 = (inp[4]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node6641 = (inp[1]) ? node6645 : node6642;
													assign node6642 = (inp[3]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node6645 = (inp[11]) ? 15'b000000000001111 : 15'b000000000001111;
								assign node6648 = (inp[4]) ? node6704 : node6649;
									assign node6649 = (inp[2]) ? node6677 : node6650;
										assign node6650 = (inp[3]) ? node6662 : node6651;
											assign node6651 = (inp[1]) ? node6657 : node6652;
												assign node6652 = (inp[11]) ? node6654 : 15'b000000111111111;
													assign node6654 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node6657 = (inp[0]) ? 15'b000000001111111 : node6658;
													assign node6658 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node6662 = (inp[11]) ? node6670 : node6663;
												assign node6663 = (inp[0]) ? node6667 : node6664;
													assign node6664 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node6667 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node6670 = (inp[1]) ? node6674 : node6671;
													assign node6671 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node6674 = (inp[9]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node6677 = (inp[3]) ? node6693 : node6678;
											assign node6678 = (inp[0]) ? node6686 : node6679;
												assign node6679 = (inp[10]) ? node6683 : node6680;
													assign node6680 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node6683 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node6686 = (inp[1]) ? node6690 : node6687;
													assign node6687 = (inp[10]) ? 15'b000000000011111 : 15'b000000001111111;
													assign node6690 = (inp[11]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node6693 = (inp[10]) ? node6699 : node6694;
												assign node6694 = (inp[11]) ? node6696 : 15'b000000000111111;
													assign node6696 = (inp[1]) ? 15'b000000000001111 : 15'b000000000111111;
												assign node6699 = (inp[0]) ? 15'b000000000011111 : node6700;
													assign node6700 = (inp[11]) ? 15'b000000000011111 : 15'b000000000011111;
									assign node6704 = (inp[1]) ? node6736 : node6705;
										assign node6705 = (inp[11]) ? node6721 : node6706;
											assign node6706 = (inp[3]) ? node6714 : node6707;
												assign node6707 = (inp[2]) ? node6711 : node6708;
													assign node6708 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node6711 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node6714 = (inp[10]) ? node6718 : node6715;
													assign node6715 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node6718 = (inp[0]) ? 15'b000000000011111 : 15'b000000000011111;
											assign node6721 = (inp[9]) ? node6729 : node6722;
												assign node6722 = (inp[10]) ? node6726 : node6723;
													assign node6723 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node6726 = (inp[0]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node6729 = (inp[0]) ? node6733 : node6730;
													assign node6730 = (inp[2]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node6733 = (inp[3]) ? 15'b000000000000111 : 15'b000000000011111;
										assign node6736 = (inp[9]) ? node6752 : node6737;
											assign node6737 = (inp[3]) ? node6745 : node6738;
												assign node6738 = (inp[10]) ? node6742 : node6739;
													assign node6739 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node6742 = (inp[11]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node6745 = (inp[0]) ? node6749 : node6746;
													assign node6746 = (inp[11]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node6749 = (inp[2]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node6752 = (inp[10]) ? node6760 : node6753;
												assign node6753 = (inp[3]) ? node6757 : node6754;
													assign node6754 = (inp[0]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node6757 = (inp[2]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node6760 = (inp[2]) ? node6764 : node6761;
													assign node6761 = (inp[3]) ? 15'b000000000001111 : 15'b000000000011111;
													assign node6764 = (inp[0]) ? 15'b000000000000111 : 15'b000000000001111;
					assign node6767 = (inp[2]) ? node7261 : node6768;
						assign node6768 = (inp[3]) ? node7018 : node6769;
							assign node6769 = (inp[8]) ? node6893 : node6770;
								assign node6770 = (inp[1]) ? node6832 : node6771;
									assign node6771 = (inp[12]) ? node6803 : node6772;
										assign node6772 = (inp[9]) ? node6788 : node6773;
											assign node6773 = (inp[10]) ? node6781 : node6774;
												assign node6774 = (inp[14]) ? node6778 : node6775;
													assign node6775 = (inp[0]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node6778 = (inp[11]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node6781 = (inp[4]) ? node6785 : node6782;
													assign node6782 = (inp[11]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node6785 = (inp[11]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node6788 = (inp[4]) ? node6796 : node6789;
												assign node6789 = (inp[14]) ? node6793 : node6790;
													assign node6790 = (inp[10]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node6793 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node6796 = (inp[11]) ? node6800 : node6797;
													assign node6797 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node6800 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node6803 = (inp[11]) ? node6817 : node6804;
											assign node6804 = (inp[0]) ? node6812 : node6805;
												assign node6805 = (inp[4]) ? node6809 : node6806;
													assign node6806 = (inp[10]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node6809 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node6812 = (inp[9]) ? 15'b000000011111111 : node6813;
													assign node6813 = (inp[4]) ? 15'b000000011111111 : 15'b000000011111111;
											assign node6817 = (inp[14]) ? node6825 : node6818;
												assign node6818 = (inp[0]) ? node6822 : node6819;
													assign node6819 = (inp[4]) ? 15'b000000011111111 : 15'b000001111111111;
													assign node6822 = (inp[9]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node6825 = (inp[10]) ? node6829 : node6826;
													assign node6826 = (inp[0]) ? 15'b000000001111111 : 15'b000000001111111;
													assign node6829 = (inp[4]) ? 15'b000000000011111 : 15'b000000001111111;
									assign node6832 = (inp[11]) ? node6864 : node6833;
										assign node6833 = (inp[9]) ? node6849 : node6834;
											assign node6834 = (inp[12]) ? node6842 : node6835;
												assign node6835 = (inp[14]) ? node6839 : node6836;
													assign node6836 = (inp[0]) ? 15'b000001111111111 : 15'b000001111111111;
													assign node6839 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node6842 = (inp[10]) ? node6846 : node6843;
													assign node6843 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node6846 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node6849 = (inp[10]) ? node6857 : node6850;
												assign node6850 = (inp[14]) ? node6854 : node6851;
													assign node6851 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node6854 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node6857 = (inp[12]) ? node6861 : node6858;
													assign node6858 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node6861 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node6864 = (inp[0]) ? node6878 : node6865;
											assign node6865 = (inp[14]) ? node6871 : node6866;
												assign node6866 = (inp[12]) ? node6868 : 15'b000000111111111;
													assign node6868 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node6871 = (inp[12]) ? node6875 : node6872;
													assign node6872 = (inp[9]) ? 15'b000000001111111 : 15'b000000001111111;
													assign node6875 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node6878 = (inp[10]) ? node6886 : node6879;
												assign node6879 = (inp[9]) ? node6883 : node6880;
													assign node6880 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node6883 = (inp[12]) ? 15'b000000000011111 : 15'b000000001111111;
												assign node6886 = (inp[4]) ? node6890 : node6887;
													assign node6887 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node6890 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
								assign node6893 = (inp[4]) ? node6955 : node6894;
									assign node6894 = (inp[14]) ? node6924 : node6895;
										assign node6895 = (inp[0]) ? node6909 : node6896;
											assign node6896 = (inp[11]) ? node6902 : node6897;
												assign node6897 = (inp[9]) ? 15'b000000111111111 : node6898;
													assign node6898 = (inp[1]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node6902 = (inp[10]) ? node6906 : node6903;
													assign node6903 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node6906 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node6909 = (inp[9]) ? node6917 : node6910;
												assign node6910 = (inp[10]) ? node6914 : node6911;
													assign node6911 = (inp[11]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node6914 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node6917 = (inp[10]) ? node6921 : node6918;
													assign node6918 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node6921 = (inp[1]) ? 15'b000000000011111 : 15'b000000001111111;
										assign node6924 = (inp[1]) ? node6940 : node6925;
											assign node6925 = (inp[11]) ? node6933 : node6926;
												assign node6926 = (inp[0]) ? node6930 : node6927;
													assign node6927 = (inp[12]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node6930 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node6933 = (inp[0]) ? node6937 : node6934;
													assign node6934 = (inp[12]) ? 15'b000000001111111 : 15'b000000001111111;
													assign node6937 = (inp[9]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node6940 = (inp[9]) ? node6948 : node6941;
												assign node6941 = (inp[0]) ? node6945 : node6942;
													assign node6942 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node6945 = (inp[12]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node6948 = (inp[12]) ? node6952 : node6949;
													assign node6949 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node6952 = (inp[11]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node6955 = (inp[12]) ? node6987 : node6956;
										assign node6956 = (inp[9]) ? node6972 : node6957;
											assign node6957 = (inp[1]) ? node6965 : node6958;
												assign node6958 = (inp[0]) ? node6962 : node6959;
													assign node6959 = (inp[14]) ? 15'b000000001111111 : 15'b000000111111111;
													assign node6962 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node6965 = (inp[0]) ? node6969 : node6966;
													assign node6966 = (inp[11]) ? 15'b000000001111111 : 15'b000000001111111;
													assign node6969 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node6972 = (inp[14]) ? node6980 : node6973;
												assign node6973 = (inp[0]) ? node6977 : node6974;
													assign node6974 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node6977 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node6980 = (inp[10]) ? node6984 : node6981;
													assign node6981 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node6984 = (inp[11]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node6987 = (inp[11]) ? node7003 : node6988;
											assign node6988 = (inp[0]) ? node6996 : node6989;
												assign node6989 = (inp[9]) ? node6993 : node6990;
													assign node6990 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node6993 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node6996 = (inp[10]) ? node7000 : node6997;
													assign node6997 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node7000 = (inp[1]) ? 15'b000000000001111 : 15'b000000000111111;
											assign node7003 = (inp[14]) ? node7011 : node7004;
												assign node7004 = (inp[9]) ? node7008 : node7005;
													assign node7005 = (inp[0]) ? 15'b000000000011111 : 15'b000000001111111;
													assign node7008 = (inp[1]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node7011 = (inp[1]) ? node7015 : node7012;
													assign node7012 = (inp[0]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node7015 = (inp[0]) ? 15'b000000000001111 : 15'b000000000011111;
							assign node7018 = (inp[11]) ? node7140 : node7019;
								assign node7019 = (inp[14]) ? node7083 : node7020;
									assign node7020 = (inp[0]) ? node7052 : node7021;
										assign node7021 = (inp[8]) ? node7037 : node7022;
											assign node7022 = (inp[4]) ? node7030 : node7023;
												assign node7023 = (inp[10]) ? node7027 : node7024;
													assign node7024 = (inp[12]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node7027 = (inp[12]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node7030 = (inp[9]) ? node7034 : node7031;
													assign node7031 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node7034 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node7037 = (inp[10]) ? node7045 : node7038;
												assign node7038 = (inp[9]) ? node7042 : node7039;
													assign node7039 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node7042 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node7045 = (inp[12]) ? node7049 : node7046;
													assign node7046 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node7049 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node7052 = (inp[9]) ? node7068 : node7053;
											assign node7053 = (inp[12]) ? node7061 : node7054;
												assign node7054 = (inp[4]) ? node7058 : node7055;
													assign node7055 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node7058 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node7061 = (inp[8]) ? node7065 : node7062;
													assign node7062 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node7065 = (inp[1]) ? 15'b000000000011111 : 15'b000000001111111;
											assign node7068 = (inp[8]) ? node7076 : node7069;
												assign node7069 = (inp[12]) ? node7073 : node7070;
													assign node7070 = (inp[10]) ? 15'b000000001111111 : 15'b000000001111111;
													assign node7073 = (inp[10]) ? 15'b000000000111111 : 15'b000000000111111;
												assign node7076 = (inp[10]) ? node7080 : node7077;
													assign node7077 = (inp[4]) ? 15'b000000000111111 : 15'b000000000111111;
													assign node7080 = (inp[4]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node7083 = (inp[9]) ? node7111 : node7084;
										assign node7084 = (inp[10]) ? node7098 : node7085;
											assign node7085 = (inp[0]) ? node7091 : node7086;
												assign node7086 = (inp[12]) ? 15'b000000011111111 : node7087;
													assign node7087 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node7091 = (inp[12]) ? node7095 : node7092;
													assign node7092 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node7095 = (inp[8]) ? 15'b000000000011111 : 15'b000000001111111;
											assign node7098 = (inp[1]) ? node7106 : node7099;
												assign node7099 = (inp[4]) ? node7103 : node7100;
													assign node7100 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node7103 = (inp[12]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node7106 = (inp[8]) ? node7108 : 15'b000000000111111;
													assign node7108 = (inp[4]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node7111 = (inp[12]) ? node7125 : node7112;
											assign node7112 = (inp[1]) ? node7118 : node7113;
												assign node7113 = (inp[4]) ? node7115 : 15'b000000001111111;
													assign node7115 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node7118 = (inp[8]) ? node7122 : node7119;
													assign node7119 = (inp[4]) ? 15'b000000000111111 : 15'b000000000111111;
													assign node7122 = (inp[4]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node7125 = (inp[4]) ? node7133 : node7126;
												assign node7126 = (inp[0]) ? node7130 : node7127;
													assign node7127 = (inp[8]) ? 15'b000000000011111 : 15'b000000001111111;
													assign node7130 = (inp[8]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node7133 = (inp[10]) ? node7137 : node7134;
													assign node7134 = (inp[8]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node7137 = (inp[1]) ? 15'b000000000001111 : 15'b000000000011111;
								assign node7140 = (inp[4]) ? node7202 : node7141;
									assign node7141 = (inp[10]) ? node7171 : node7142;
										assign node7142 = (inp[12]) ? node7156 : node7143;
											assign node7143 = (inp[8]) ? node7149 : node7144;
												assign node7144 = (inp[0]) ? 15'b000000011111111 : node7145;
													assign node7145 = (inp[1]) ? 15'b000000011111111 : 15'b000001111111111;
												assign node7149 = (inp[0]) ? node7153 : node7150;
													assign node7150 = (inp[9]) ? 15'b000000001111111 : 15'b000000111111111;
													assign node7153 = (inp[9]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node7156 = (inp[1]) ? node7164 : node7157;
												assign node7157 = (inp[8]) ? node7161 : node7158;
													assign node7158 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node7161 = (inp[0]) ? 15'b000000000111111 : 15'b000000000111111;
												assign node7164 = (inp[0]) ? node7168 : node7165;
													assign node7165 = (inp[9]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node7168 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node7171 = (inp[0]) ? node7187 : node7172;
											assign node7172 = (inp[8]) ? node7180 : node7173;
												assign node7173 = (inp[1]) ? node7177 : node7174;
													assign node7174 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node7177 = (inp[9]) ? 15'b000000000111111 : 15'b000000000111111;
												assign node7180 = (inp[9]) ? node7184 : node7181;
													assign node7181 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node7184 = (inp[1]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node7187 = (inp[12]) ? node7195 : node7188;
												assign node7188 = (inp[1]) ? node7192 : node7189;
													assign node7189 = (inp[14]) ? 15'b000000000111111 : 15'b000000011111111;
													assign node7192 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node7195 = (inp[9]) ? node7199 : node7196;
													assign node7196 = (inp[8]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node7199 = (inp[8]) ? 15'b000000000001111 : 15'b000000000011111;
									assign node7202 = (inp[9]) ? node7232 : node7203;
										assign node7203 = (inp[1]) ? node7219 : node7204;
											assign node7204 = (inp[12]) ? node7212 : node7205;
												assign node7205 = (inp[10]) ? node7209 : node7206;
													assign node7206 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node7209 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node7212 = (inp[14]) ? node7216 : node7213;
													assign node7213 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node7216 = (inp[10]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node7219 = (inp[0]) ? node7227 : node7220;
												assign node7220 = (inp[10]) ? node7224 : node7221;
													assign node7221 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node7224 = (inp[12]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node7227 = (inp[8]) ? node7229 : 15'b000000000011111;
													assign node7229 = (inp[14]) ? 15'b000000000000111 : 15'b000000000011111;
										assign node7232 = (inp[14]) ? node7248 : node7233;
											assign node7233 = (inp[8]) ? node7241 : node7234;
												assign node7234 = (inp[12]) ? node7238 : node7235;
													assign node7235 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node7238 = (inp[10]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node7241 = (inp[0]) ? node7245 : node7242;
													assign node7242 = (inp[10]) ? 15'b000000000011111 : 15'b000000000011111;
													assign node7245 = (inp[12]) ? 15'b000000000001111 : 15'b000000000001111;
											assign node7248 = (inp[10]) ? node7254 : node7249;
												assign node7249 = (inp[12]) ? node7251 : 15'b000000000011111;
													assign node7251 = (inp[1]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node7254 = (inp[1]) ? node7258 : node7255;
													assign node7255 = (inp[0]) ? 15'b000000000001111 : 15'b000000000001111;
													assign node7258 = (inp[8]) ? 15'b000000000000111 : 15'b000000000001111;
						assign node7261 = (inp[1]) ? node7505 : node7262;
							assign node7262 = (inp[9]) ? node7382 : node7263;
								assign node7263 = (inp[12]) ? node7321 : node7264;
									assign node7264 = (inp[4]) ? node7294 : node7265;
										assign node7265 = (inp[10]) ? node7279 : node7266;
											assign node7266 = (inp[11]) ? node7274 : node7267;
												assign node7267 = (inp[3]) ? node7271 : node7268;
													assign node7268 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node7271 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node7274 = (inp[3]) ? 15'b000000011111111 : node7275;
													assign node7275 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node7279 = (inp[8]) ? node7287 : node7280;
												assign node7280 = (inp[0]) ? node7284 : node7281;
													assign node7281 = (inp[3]) ? 15'b000000011111111 : 15'b000001111111111;
													assign node7284 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node7287 = (inp[0]) ? node7291 : node7288;
													assign node7288 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node7291 = (inp[14]) ? 15'b000000000011111 : 15'b000000001111111;
										assign node7294 = (inp[8]) ? node7308 : node7295;
											assign node7295 = (inp[3]) ? node7301 : node7296;
												assign node7296 = (inp[14]) ? node7298 : 15'b000000011111111;
													assign node7298 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node7301 = (inp[0]) ? node7305 : node7302;
													assign node7302 = (inp[14]) ? 15'b000000001111111 : 15'b000000111111111;
													assign node7305 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node7308 = (inp[0]) ? node7316 : node7309;
												assign node7309 = (inp[10]) ? node7313 : node7310;
													assign node7310 = (inp[11]) ? 15'b000000001111111 : 15'b000000001111111;
													assign node7313 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node7316 = (inp[11]) ? node7318 : 15'b000000000111111;
													assign node7318 = (inp[3]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node7321 = (inp[10]) ? node7353 : node7322;
										assign node7322 = (inp[14]) ? node7338 : node7323;
											assign node7323 = (inp[11]) ? node7331 : node7324;
												assign node7324 = (inp[8]) ? node7328 : node7325;
													assign node7325 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node7328 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node7331 = (inp[4]) ? node7335 : node7332;
													assign node7332 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node7335 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node7338 = (inp[0]) ? node7346 : node7339;
												assign node7339 = (inp[3]) ? node7343 : node7340;
													assign node7340 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node7343 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node7346 = (inp[8]) ? node7350 : node7347;
													assign node7347 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node7350 = (inp[3]) ? 15'b000000000001111 : 15'b000000000111111;
										assign node7353 = (inp[3]) ? node7367 : node7354;
											assign node7354 = (inp[0]) ? node7362 : node7355;
												assign node7355 = (inp[11]) ? node7359 : node7356;
													assign node7356 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node7359 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node7362 = (inp[4]) ? 15'b000000000011111 : node7363;
													assign node7363 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node7367 = (inp[4]) ? node7375 : node7368;
												assign node7368 = (inp[14]) ? node7372 : node7369;
													assign node7369 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node7372 = (inp[11]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node7375 = (inp[14]) ? node7379 : node7376;
													assign node7376 = (inp[0]) ? 15'b000000000011111 : 15'b000000000011111;
													assign node7379 = (inp[8]) ? 15'b000000000001111 : 15'b000000000011111;
								assign node7382 = (inp[8]) ? node7444 : node7383;
									assign node7383 = (inp[11]) ? node7415 : node7384;
										assign node7384 = (inp[0]) ? node7400 : node7385;
											assign node7385 = (inp[14]) ? node7393 : node7386;
												assign node7386 = (inp[4]) ? node7390 : node7387;
													assign node7387 = (inp[12]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node7390 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node7393 = (inp[4]) ? node7397 : node7394;
													assign node7394 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node7397 = (inp[10]) ? 15'b000000000011111 : 15'b000000001111111;
											assign node7400 = (inp[14]) ? node7408 : node7401;
												assign node7401 = (inp[10]) ? node7405 : node7402;
													assign node7402 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node7405 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node7408 = (inp[10]) ? node7412 : node7409;
													assign node7409 = (inp[12]) ? 15'b000000000111111 : 15'b000000000111111;
													assign node7412 = (inp[12]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node7415 = (inp[3]) ? node7429 : node7416;
											assign node7416 = (inp[10]) ? node7422 : node7417;
												assign node7417 = (inp[14]) ? node7419 : 15'b000000011111111;
													assign node7419 = (inp[12]) ? 15'b000000001111111 : 15'b000000001111111;
												assign node7422 = (inp[12]) ? node7426 : node7423;
													assign node7423 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node7426 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node7429 = (inp[10]) ? node7437 : node7430;
												assign node7430 = (inp[4]) ? node7434 : node7431;
													assign node7431 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node7434 = (inp[12]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node7437 = (inp[14]) ? node7441 : node7438;
													assign node7438 = (inp[12]) ? 15'b000000000011111 : 15'b000000000011111;
													assign node7441 = (inp[4]) ? 15'b000000000001111 : 15'b000000000011111;
									assign node7444 = (inp[0]) ? node7476 : node7445;
										assign node7445 = (inp[12]) ? node7461 : node7446;
											assign node7446 = (inp[14]) ? node7454 : node7447;
												assign node7447 = (inp[3]) ? node7451 : node7448;
													assign node7448 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node7451 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node7454 = (inp[4]) ? node7458 : node7455;
													assign node7455 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node7458 = (inp[11]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node7461 = (inp[11]) ? node7469 : node7462;
												assign node7462 = (inp[3]) ? node7466 : node7463;
													assign node7463 = (inp[14]) ? 15'b000000000111111 : 15'b000000000111111;
													assign node7466 = (inp[10]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node7469 = (inp[3]) ? node7473 : node7470;
													assign node7470 = (inp[10]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node7473 = (inp[4]) ? 15'b000000000001111 : 15'b000000000011111;
										assign node7476 = (inp[10]) ? node7490 : node7477;
											assign node7477 = (inp[12]) ? node7483 : node7478;
												assign node7478 = (inp[14]) ? 15'b000000000111111 : node7479;
													assign node7479 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node7483 = (inp[4]) ? node7487 : node7484;
													assign node7484 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node7487 = (inp[3]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node7490 = (inp[3]) ? node7498 : node7491;
												assign node7491 = (inp[4]) ? node7495 : node7492;
													assign node7492 = (inp[11]) ? 15'b000000000001111 : 15'b000000000111111;
													assign node7495 = (inp[12]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node7498 = (inp[4]) ? node7502 : node7499;
													assign node7499 = (inp[14]) ? 15'b000000000001111 : 15'b000000000001111;
													assign node7502 = (inp[14]) ? 15'b000000000000111 : 15'b000000000001111;
							assign node7505 = (inp[11]) ? node7629 : node7506;
								assign node7506 = (inp[8]) ? node7566 : node7507;
									assign node7507 = (inp[12]) ? node7537 : node7508;
										assign node7508 = (inp[3]) ? node7524 : node7509;
											assign node7509 = (inp[10]) ? node7517 : node7510;
												assign node7510 = (inp[9]) ? node7514 : node7511;
													assign node7511 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node7514 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node7517 = (inp[14]) ? node7521 : node7518;
													assign node7518 = (inp[9]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node7521 = (inp[9]) ? 15'b000000000011111 : 15'b000000001111111;
											assign node7524 = (inp[9]) ? node7530 : node7525;
												assign node7525 = (inp[14]) ? 15'b000000001111111 : node7526;
													assign node7526 = (inp[0]) ? 15'b000000001111111 : 15'b000000111111111;
												assign node7530 = (inp[10]) ? node7534 : node7531;
													assign node7531 = (inp[4]) ? 15'b000000000011111 : 15'b000000001111111;
													assign node7534 = (inp[0]) ? 15'b000000000111111 : 15'b000000000111111;
										assign node7537 = (inp[9]) ? node7551 : node7538;
											assign node7538 = (inp[3]) ? node7546 : node7539;
												assign node7539 = (inp[10]) ? node7543 : node7540;
													assign node7540 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node7543 = (inp[0]) ? 15'b000000000111111 : 15'b000000000111111;
												assign node7546 = (inp[10]) ? node7548 : 15'b000000000111111;
													assign node7548 = (inp[4]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node7551 = (inp[4]) ? node7559 : node7552;
												assign node7552 = (inp[10]) ? node7556 : node7553;
													assign node7553 = (inp[3]) ? 15'b000000000111111 : 15'b000000000111111;
													assign node7556 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node7559 = (inp[0]) ? node7563 : node7560;
													assign node7560 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node7563 = (inp[10]) ? 15'b000000000001111 : 15'b000000000011111;
									assign node7566 = (inp[4]) ? node7598 : node7567;
										assign node7567 = (inp[3]) ? node7583 : node7568;
											assign node7568 = (inp[9]) ? node7576 : node7569;
												assign node7569 = (inp[14]) ? node7573 : node7570;
													assign node7570 = (inp[0]) ? 15'b000000001111111 : 15'b000000001111111;
													assign node7573 = (inp[12]) ? 15'b000000000111111 : 15'b000000000111111;
												assign node7576 = (inp[10]) ? node7580 : node7577;
													assign node7577 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node7580 = (inp[0]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node7583 = (inp[14]) ? node7591 : node7584;
												assign node7584 = (inp[10]) ? node7588 : node7585;
													assign node7585 = (inp[12]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node7588 = (inp[9]) ? 15'b000000000011111 : 15'b000000000011111;
												assign node7591 = (inp[9]) ? node7595 : node7592;
													assign node7592 = (inp[0]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node7595 = (inp[0]) ? 15'b000000000001111 : 15'b000000000011111;
										assign node7598 = (inp[3]) ? node7614 : node7599;
											assign node7599 = (inp[14]) ? node7607 : node7600;
												assign node7600 = (inp[9]) ? node7604 : node7601;
													assign node7601 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node7604 = (inp[10]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node7607 = (inp[12]) ? node7611 : node7608;
													assign node7608 = (inp[9]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node7611 = (inp[10]) ? 15'b000000000001111 : 15'b000000000001111;
											assign node7614 = (inp[14]) ? node7622 : node7615;
												assign node7615 = (inp[9]) ? node7619 : node7616;
													assign node7616 = (inp[10]) ? 15'b000000000011111 : 15'b000000000011111;
													assign node7619 = (inp[0]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node7622 = (inp[10]) ? node7626 : node7623;
													assign node7623 = (inp[9]) ? 15'b000000000001111 : 15'b000000000011111;
													assign node7626 = (inp[12]) ? 15'b000000000000111 : 15'b000000000001111;
								assign node7629 = (inp[9]) ? node7691 : node7630;
									assign node7630 = (inp[10]) ? node7660 : node7631;
										assign node7631 = (inp[0]) ? node7645 : node7632;
											assign node7632 = (inp[12]) ? node7640 : node7633;
												assign node7633 = (inp[14]) ? node7637 : node7634;
													assign node7634 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node7637 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node7640 = (inp[8]) ? 15'b000000000111111 : node7641;
													assign node7641 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node7645 = (inp[14]) ? node7653 : node7646;
												assign node7646 = (inp[8]) ? node7650 : node7647;
													assign node7647 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node7650 = (inp[12]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node7653 = (inp[4]) ? node7657 : node7654;
													assign node7654 = (inp[8]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node7657 = (inp[3]) ? 15'b000000000001111 : 15'b000000000011111;
										assign node7660 = (inp[12]) ? node7676 : node7661;
											assign node7661 = (inp[4]) ? node7669 : node7662;
												assign node7662 = (inp[8]) ? node7666 : node7663;
													assign node7663 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node7666 = (inp[3]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node7669 = (inp[14]) ? node7673 : node7670;
													assign node7670 = (inp[0]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node7673 = (inp[0]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node7676 = (inp[14]) ? node7684 : node7677;
												assign node7677 = (inp[0]) ? node7681 : node7678;
													assign node7678 = (inp[4]) ? 15'b000000000011111 : 15'b000000000011111;
													assign node7681 = (inp[4]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node7684 = (inp[8]) ? node7688 : node7685;
													assign node7685 = (inp[0]) ? 15'b000000000001111 : 15'b000000000011111;
													assign node7688 = (inp[3]) ? 15'b000000000000111 : 15'b000000000001111;
									assign node7691 = (inp[8]) ? node7723 : node7692;
										assign node7692 = (inp[12]) ? node7708 : node7693;
											assign node7693 = (inp[3]) ? node7701 : node7694;
												assign node7694 = (inp[0]) ? node7698 : node7695;
													assign node7695 = (inp[14]) ? 15'b000000001111111 : 15'b000000001111111;
													assign node7698 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node7701 = (inp[14]) ? node7705 : node7702;
													assign node7702 = (inp[4]) ? 15'b000000000111111 : 15'b000000000011111;
													assign node7705 = (inp[0]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node7708 = (inp[10]) ? node7716 : node7709;
												assign node7709 = (inp[4]) ? node7713 : node7710;
													assign node7710 = (inp[0]) ? 15'b000000000011111 : 15'b000000000011111;
													assign node7713 = (inp[14]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node7716 = (inp[0]) ? node7720 : node7717;
													assign node7717 = (inp[14]) ? 15'b000000000001111 : 15'b000000000001111;
													assign node7720 = (inp[3]) ? 15'b000000000000111 : 15'b000000000001111;
										assign node7723 = (inp[12]) ? node7739 : node7724;
											assign node7724 = (inp[4]) ? node7732 : node7725;
												assign node7725 = (inp[0]) ? node7729 : node7726;
													assign node7726 = (inp[3]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node7729 = (inp[10]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node7732 = (inp[14]) ? node7736 : node7733;
													assign node7733 = (inp[10]) ? 15'b000000000001111 : 15'b000000000011111;
													assign node7736 = (inp[3]) ? 15'b000000000000111 : 15'b000000000001111;
											assign node7739 = (inp[4]) ? node7747 : node7740;
												assign node7740 = (inp[3]) ? node7744 : node7741;
													assign node7741 = (inp[0]) ? 15'b000000000001111 : 15'b000000000001111;
													assign node7744 = (inp[10]) ? 15'b000000000000111 : 15'b000000000001111;
												assign node7747 = (inp[14]) ? node7751 : node7748;
													assign node7748 = (inp[10]) ? 15'b000000000000111 : 15'b000000000001111;
													assign node7751 = (inp[3]) ? 15'b000000000000011 : 15'b000000000000111;
		assign node7754 = (inp[0]) ? node11634 : node7755;
			assign node7755 = (inp[13]) ? node9723 : node7756;
				assign node7756 = (inp[2]) ? node8752 : node7757;
					assign node7757 = (inp[5]) ? node8253 : node7758;
						assign node7758 = (inp[14]) ? node8006 : node7759;
							assign node7759 = (inp[9]) ? node7879 : node7760;
								assign node7760 = (inp[10]) ? node7818 : node7761;
									assign node7761 = (inp[12]) ? node7789 : node7762;
										assign node7762 = (inp[4]) ? node7778 : node7763;
											assign node7763 = (inp[11]) ? node7771 : node7764;
												assign node7764 = (inp[3]) ? node7768 : node7765;
													assign node7765 = (inp[8]) ? 15'b000111111111111 : 15'b001111111111111;
													assign node7768 = (inp[7]) ? 15'b000011111111111 : 15'b000111111111111;
												assign node7771 = (inp[8]) ? node7775 : node7772;
													assign node7772 = (inp[7]) ? 15'b000011111111111 : 15'b000111111111111;
													assign node7775 = (inp[1]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node7778 = (inp[11]) ? node7784 : node7779;
												assign node7779 = (inp[7]) ? node7781 : 15'b000011111111111;
													assign node7781 = (inp[1]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node7784 = (inp[1]) ? 15'b000001111111111 : node7785;
													assign node7785 = (inp[8]) ? 15'b000001111111111 : 15'b000011111111111;
										assign node7789 = (inp[4]) ? node7805 : node7790;
											assign node7790 = (inp[7]) ? node7798 : node7791;
												assign node7791 = (inp[1]) ? node7795 : node7792;
													assign node7792 = (inp[11]) ? 15'b000011111111111 : 15'b000011111111111;
													assign node7795 = (inp[8]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node7798 = (inp[11]) ? node7802 : node7799;
													assign node7799 = (inp[3]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node7802 = (inp[3]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node7805 = (inp[11]) ? node7811 : node7806;
												assign node7806 = (inp[1]) ? 15'b000000111111111 : node7807;
													assign node7807 = (inp[7]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node7811 = (inp[8]) ? node7815 : node7812;
													assign node7812 = (inp[3]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node7815 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node7818 = (inp[12]) ? node7848 : node7819;
										assign node7819 = (inp[11]) ? node7835 : node7820;
											assign node7820 = (inp[8]) ? node7828 : node7821;
												assign node7821 = (inp[4]) ? node7825 : node7822;
													assign node7822 = (inp[7]) ? 15'b000011111111111 : 15'b000111111111111;
													assign node7825 = (inp[3]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node7828 = (inp[4]) ? node7832 : node7829;
													assign node7829 = (inp[7]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node7832 = (inp[1]) ? 15'b000000011111111 : 15'b000001111111111;
											assign node7835 = (inp[3]) ? node7843 : node7836;
												assign node7836 = (inp[1]) ? node7840 : node7837;
													assign node7837 = (inp[4]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node7840 = (inp[7]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node7843 = (inp[1]) ? node7845 : 15'b000000111111111;
													assign node7845 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node7848 = (inp[4]) ? node7864 : node7849;
											assign node7849 = (inp[7]) ? node7857 : node7850;
												assign node7850 = (inp[11]) ? node7854 : node7851;
													assign node7851 = (inp[1]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node7854 = (inp[1]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node7857 = (inp[8]) ? node7861 : node7858;
													assign node7858 = (inp[1]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node7861 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node7864 = (inp[8]) ? node7872 : node7865;
												assign node7865 = (inp[1]) ? node7869 : node7866;
													assign node7866 = (inp[11]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node7869 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node7872 = (inp[1]) ? node7876 : node7873;
													assign node7873 = (inp[11]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node7876 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
								assign node7879 = (inp[7]) ? node7943 : node7880;
									assign node7880 = (inp[11]) ? node7912 : node7881;
										assign node7881 = (inp[3]) ? node7897 : node7882;
											assign node7882 = (inp[12]) ? node7890 : node7883;
												assign node7883 = (inp[1]) ? node7887 : node7884;
													assign node7884 = (inp[4]) ? 15'b000011111111111 : 15'b000111111111111;
													assign node7887 = (inp[10]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node7890 = (inp[4]) ? node7894 : node7891;
													assign node7891 = (inp[1]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node7894 = (inp[8]) ? 15'b000000111111111 : 15'b000011111111111;
											assign node7897 = (inp[4]) ? node7905 : node7898;
												assign node7898 = (inp[12]) ? node7902 : node7899;
													assign node7899 = (inp[8]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node7902 = (inp[1]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node7905 = (inp[1]) ? node7909 : node7906;
													assign node7906 = (inp[10]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node7909 = (inp[12]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node7912 = (inp[8]) ? node7928 : node7913;
											assign node7913 = (inp[4]) ? node7921 : node7914;
												assign node7914 = (inp[10]) ? node7918 : node7915;
													assign node7915 = (inp[1]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node7918 = (inp[12]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node7921 = (inp[1]) ? node7925 : node7922;
													assign node7922 = (inp[10]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node7925 = (inp[12]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node7928 = (inp[10]) ? node7936 : node7929;
												assign node7929 = (inp[12]) ? node7933 : node7930;
													assign node7930 = (inp[4]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node7933 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node7936 = (inp[4]) ? node7940 : node7937;
													assign node7937 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node7940 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node7943 = (inp[10]) ? node7975 : node7944;
										assign node7944 = (inp[4]) ? node7960 : node7945;
											assign node7945 = (inp[12]) ? node7953 : node7946;
												assign node7946 = (inp[8]) ? node7950 : node7947;
													assign node7947 = (inp[3]) ? 15'b000001111111111 : 15'b000001111111111;
													assign node7950 = (inp[11]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node7953 = (inp[3]) ? node7957 : node7954;
													assign node7954 = (inp[8]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node7957 = (inp[11]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node7960 = (inp[3]) ? node7968 : node7961;
												assign node7961 = (inp[8]) ? node7965 : node7962;
													assign node7962 = (inp[11]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node7965 = (inp[12]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node7968 = (inp[8]) ? node7972 : node7969;
													assign node7969 = (inp[11]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node7972 = (inp[12]) ? 15'b000000001111111 : 15'b000000001111111;
										assign node7975 = (inp[11]) ? node7991 : node7976;
											assign node7976 = (inp[12]) ? node7984 : node7977;
												assign node7977 = (inp[4]) ? node7981 : node7978;
													assign node7978 = (inp[8]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node7981 = (inp[1]) ? 15'b000000001111111 : 15'b000000111111111;
												assign node7984 = (inp[3]) ? node7988 : node7985;
													assign node7985 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node7988 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node7991 = (inp[1]) ? node7999 : node7992;
												assign node7992 = (inp[12]) ? node7996 : node7993;
													assign node7993 = (inp[4]) ? 15'b000000011111111 : 15'b000000011111111;
													assign node7996 = (inp[4]) ? 15'b000000000111111 : 15'b000000011111111;
												assign node7999 = (inp[12]) ? node8003 : node8000;
													assign node8000 = (inp[3]) ? 15'b000000001111111 : 15'b000000111111111;
													assign node8003 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
							assign node8006 = (inp[9]) ? node8130 : node8007;
								assign node8007 = (inp[12]) ? node8069 : node8008;
									assign node8008 = (inp[4]) ? node8038 : node8009;
										assign node8009 = (inp[10]) ? node8025 : node8010;
											assign node8010 = (inp[3]) ? node8018 : node8011;
												assign node8011 = (inp[8]) ? node8015 : node8012;
													assign node8012 = (inp[1]) ? 15'b000011111111111 : 15'b000111111111111;
													assign node8015 = (inp[11]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node8018 = (inp[1]) ? node8022 : node8019;
													assign node8019 = (inp[7]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node8022 = (inp[11]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node8025 = (inp[3]) ? node8033 : node8026;
												assign node8026 = (inp[8]) ? node8030 : node8027;
													assign node8027 = (inp[7]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node8030 = (inp[1]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node8033 = (inp[11]) ? 15'b000000111111111 : node8034;
													assign node8034 = (inp[1]) ? 15'b000000111111111 : 15'b000000111111111;
										assign node8038 = (inp[8]) ? node8054 : node8039;
											assign node8039 = (inp[1]) ? node8047 : node8040;
												assign node8040 = (inp[7]) ? node8044 : node8041;
													assign node8041 = (inp[11]) ? 15'b000001111111111 : 15'b000001111111111;
													assign node8044 = (inp[3]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node8047 = (inp[10]) ? node8051 : node8048;
													assign node8048 = (inp[3]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node8051 = (inp[11]) ? 15'b000000001111111 : 15'b000000111111111;
											assign node8054 = (inp[3]) ? node8062 : node8055;
												assign node8055 = (inp[7]) ? node8059 : node8056;
													assign node8056 = (inp[11]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node8059 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node8062 = (inp[11]) ? node8066 : node8063;
													assign node8063 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node8066 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node8069 = (inp[1]) ? node8099 : node8070;
										assign node8070 = (inp[11]) ? node8086 : node8071;
											assign node8071 = (inp[4]) ? node8079 : node8072;
												assign node8072 = (inp[10]) ? node8076 : node8073;
													assign node8073 = (inp[3]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node8076 = (inp[7]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node8079 = (inp[8]) ? node8083 : node8080;
													assign node8080 = (inp[3]) ? 15'b000000111111111 : 15'b000000111111111;
													assign node8083 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node8086 = (inp[10]) ? node8092 : node8087;
												assign node8087 = (inp[8]) ? node8089 : 15'b000000111111111;
													assign node8089 = (inp[7]) ? 15'b000000011111111 : 15'b000001111111111;
												assign node8092 = (inp[3]) ? node8096 : node8093;
													assign node8093 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node8096 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node8099 = (inp[8]) ? node8115 : node8100;
											assign node8100 = (inp[7]) ? node8108 : node8101;
												assign node8101 = (inp[10]) ? node8105 : node8102;
													assign node8102 = (inp[11]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node8105 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node8108 = (inp[10]) ? node8112 : node8109;
													assign node8109 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node8112 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node8115 = (inp[3]) ? node8123 : node8116;
												assign node8116 = (inp[4]) ? node8120 : node8117;
													assign node8117 = (inp[7]) ? 15'b000000011111111 : 15'b000001111111111;
													assign node8120 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node8123 = (inp[10]) ? node8127 : node8124;
													assign node8124 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node8127 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
								assign node8130 = (inp[10]) ? node8194 : node8131;
									assign node8131 = (inp[8]) ? node8163 : node8132;
										assign node8132 = (inp[1]) ? node8148 : node8133;
											assign node8133 = (inp[11]) ? node8141 : node8134;
												assign node8134 = (inp[3]) ? node8138 : node8135;
													assign node8135 = (inp[12]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node8138 = (inp[4]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node8141 = (inp[3]) ? node8145 : node8142;
													assign node8142 = (inp[4]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node8145 = (inp[4]) ? 15'b000000001111111 : 15'b000000111111111;
											assign node8148 = (inp[4]) ? node8156 : node8149;
												assign node8149 = (inp[3]) ? node8153 : node8150;
													assign node8150 = (inp[12]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node8153 = (inp[11]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node8156 = (inp[3]) ? node8160 : node8157;
													assign node8157 = (inp[11]) ? 15'b000000011111111 : 15'b000000011111111;
													assign node8160 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node8163 = (inp[12]) ? node8179 : node8164;
											assign node8164 = (inp[4]) ? node8172 : node8165;
												assign node8165 = (inp[7]) ? node8169 : node8166;
													assign node8166 = (inp[1]) ? 15'b000000111111111 : 15'b000000111111111;
													assign node8169 = (inp[3]) ? 15'b000000001111111 : 15'b000000111111111;
												assign node8172 = (inp[3]) ? node8176 : node8173;
													assign node8173 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node8176 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node8179 = (inp[3]) ? node8187 : node8180;
												assign node8180 = (inp[11]) ? node8184 : node8181;
													assign node8181 = (inp[7]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node8184 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node8187 = (inp[7]) ? node8191 : node8188;
													assign node8188 = (inp[1]) ? 15'b000000000111111 : 15'b000000011111111;
													assign node8191 = (inp[11]) ? 15'b000000000111111 : 15'b000000000111111;
									assign node8194 = (inp[11]) ? node8224 : node8195;
										assign node8195 = (inp[4]) ? node8211 : node8196;
											assign node8196 = (inp[7]) ? node8204 : node8197;
												assign node8197 = (inp[12]) ? node8201 : node8198;
													assign node8198 = (inp[8]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node8201 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node8204 = (inp[1]) ? node8208 : node8205;
													assign node8205 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node8208 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node8211 = (inp[8]) ? node8219 : node8212;
												assign node8212 = (inp[3]) ? node8216 : node8213;
													assign node8213 = (inp[1]) ? 15'b000000011111111 : 15'b000000011111111;
													assign node8216 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node8219 = (inp[1]) ? 15'b000000000111111 : node8220;
													assign node8220 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node8224 = (inp[4]) ? node8240 : node8225;
											assign node8225 = (inp[1]) ? node8233 : node8226;
												assign node8226 = (inp[8]) ? node8230 : node8227;
													assign node8227 = (inp[7]) ? 15'b000000011111111 : 15'b000000011111111;
													assign node8230 = (inp[7]) ? 15'b000000000111111 : 15'b000000011111111;
												assign node8233 = (inp[3]) ? node8237 : node8234;
													assign node8234 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node8237 = (inp[7]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node8240 = (inp[7]) ? node8246 : node8241;
												assign node8241 = (inp[8]) ? node8243 : 15'b000000001111111;
													assign node8243 = (inp[12]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node8246 = (inp[3]) ? node8250 : node8247;
													assign node8247 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node8250 = (inp[1]) ? 15'b000000000011111 : 15'b000000000111111;
						assign node8253 = (inp[11]) ? node8503 : node8254;
							assign node8254 = (inp[10]) ? node8382 : node8255;
								assign node8255 = (inp[1]) ? node8319 : node8256;
									assign node8256 = (inp[8]) ? node8288 : node8257;
										assign node8257 = (inp[3]) ? node8273 : node8258;
											assign node8258 = (inp[14]) ? node8266 : node8259;
												assign node8259 = (inp[9]) ? node8263 : node8260;
													assign node8260 = (inp[4]) ? 15'b000011111111111 : 15'b000111111111111;
													assign node8263 = (inp[12]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node8266 = (inp[7]) ? node8270 : node8267;
													assign node8267 = (inp[4]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node8270 = (inp[9]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node8273 = (inp[4]) ? node8281 : node8274;
												assign node8274 = (inp[9]) ? node8278 : node8275;
													assign node8275 = (inp[12]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node8278 = (inp[7]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node8281 = (inp[14]) ? node8285 : node8282;
													assign node8282 = (inp[12]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node8285 = (inp[7]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node8288 = (inp[12]) ? node8304 : node8289;
											assign node8289 = (inp[4]) ? node8297 : node8290;
												assign node8290 = (inp[14]) ? node8294 : node8291;
													assign node8291 = (inp[7]) ? 15'b000001111111111 : 15'b000001111111111;
													assign node8294 = (inp[9]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node8297 = (inp[9]) ? node8301 : node8298;
													assign node8298 = (inp[3]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node8301 = (inp[7]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node8304 = (inp[9]) ? node8312 : node8305;
												assign node8305 = (inp[7]) ? node8309 : node8306;
													assign node8306 = (inp[14]) ? 15'b000000111111111 : 15'b000000111111111;
													assign node8309 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node8312 = (inp[3]) ? node8316 : node8313;
													assign node8313 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node8316 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node8319 = (inp[14]) ? node8351 : node8320;
										assign node8320 = (inp[4]) ? node8336 : node8321;
											assign node8321 = (inp[9]) ? node8329 : node8322;
												assign node8322 = (inp[7]) ? node8326 : node8323;
													assign node8323 = (inp[12]) ? 15'b000001111111111 : 15'b000001111111111;
													assign node8326 = (inp[3]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node8329 = (inp[12]) ? node8333 : node8330;
													assign node8330 = (inp[3]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node8333 = (inp[8]) ? 15'b000000001111111 : 15'b000000111111111;
											assign node8336 = (inp[3]) ? node8344 : node8337;
												assign node8337 = (inp[9]) ? node8341 : node8338;
													assign node8338 = (inp[7]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node8341 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node8344 = (inp[8]) ? node8348 : node8345;
													assign node8345 = (inp[12]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node8348 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node8351 = (inp[7]) ? node8367 : node8352;
											assign node8352 = (inp[4]) ? node8360 : node8353;
												assign node8353 = (inp[12]) ? node8357 : node8354;
													assign node8354 = (inp[9]) ? 15'b000000011111111 : 15'b000001111111111;
													assign node8357 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node8360 = (inp[12]) ? node8364 : node8361;
													assign node8361 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node8364 = (inp[3]) ? 15'b000000000111111 : 15'b000000011111111;
											assign node8367 = (inp[8]) ? node8375 : node8368;
												assign node8368 = (inp[9]) ? node8372 : node8369;
													assign node8369 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node8372 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node8375 = (inp[4]) ? node8379 : node8376;
													assign node8376 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node8379 = (inp[3]) ? 15'b000000000011111 : 15'b000000001111111;
								assign node8382 = (inp[3]) ? node8444 : node8383;
									assign node8383 = (inp[9]) ? node8413 : node8384;
										assign node8384 = (inp[12]) ? node8400 : node8385;
											assign node8385 = (inp[4]) ? node8393 : node8386;
												assign node8386 = (inp[1]) ? node8390 : node8387;
													assign node8387 = (inp[14]) ? 15'b000011111111111 : 15'b000011111111111;
													assign node8390 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node8393 = (inp[7]) ? node8397 : node8394;
													assign node8394 = (inp[8]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node8397 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node8400 = (inp[4]) ? node8408 : node8401;
												assign node8401 = (inp[14]) ? node8405 : node8402;
													assign node8402 = (inp[7]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node8405 = (inp[8]) ? 15'b000000111111111 : 15'b000000011111111;
												assign node8408 = (inp[1]) ? node8410 : 15'b000000011111111;
													assign node8410 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node8413 = (inp[8]) ? node8429 : node8414;
											assign node8414 = (inp[14]) ? node8422 : node8415;
												assign node8415 = (inp[1]) ? node8419 : node8416;
													assign node8416 = (inp[4]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node8419 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node8422 = (inp[7]) ? node8426 : node8423;
													assign node8423 = (inp[12]) ? 15'b000000011111111 : 15'b000001111111111;
													assign node8426 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node8429 = (inp[1]) ? node8437 : node8430;
												assign node8430 = (inp[14]) ? node8434 : node8431;
													assign node8431 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node8434 = (inp[7]) ? 15'b000000001111111 : 15'b000000111111111;
												assign node8437 = (inp[14]) ? node8441 : node8438;
													assign node8438 = (inp[4]) ? 15'b000000001111111 : 15'b000000001111111;
													assign node8441 = (inp[12]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node8444 = (inp[8]) ? node8472 : node8445;
										assign node8445 = (inp[14]) ? node8461 : node8446;
											assign node8446 = (inp[1]) ? node8454 : node8447;
												assign node8447 = (inp[9]) ? node8451 : node8448;
													assign node8448 = (inp[12]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node8451 = (inp[7]) ? 15'b000000011111111 : 15'b000000011111111;
												assign node8454 = (inp[7]) ? node8458 : node8455;
													assign node8455 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node8458 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node8461 = (inp[7]) ? node8467 : node8462;
												assign node8462 = (inp[9]) ? 15'b000000011111111 : node8463;
													assign node8463 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node8467 = (inp[12]) ? node8469 : 15'b000000001111111;
													assign node8469 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node8472 = (inp[1]) ? node8488 : node8473;
											assign node8473 = (inp[12]) ? node8481 : node8474;
												assign node8474 = (inp[4]) ? node8478 : node8475;
													assign node8475 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node8478 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node8481 = (inp[9]) ? node8485 : node8482;
													assign node8482 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node8485 = (inp[4]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node8488 = (inp[14]) ? node8496 : node8489;
												assign node8489 = (inp[12]) ? node8493 : node8490;
													assign node8490 = (inp[9]) ? 15'b000000000111111 : 15'b000000011111111;
													assign node8493 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node8496 = (inp[9]) ? node8500 : node8497;
													assign node8497 = (inp[12]) ? 15'b000000000111111 : 15'b000000000111111;
													assign node8500 = (inp[4]) ? 15'b000000000011111 : 15'b000000000011111;
							assign node8503 = (inp[12]) ? node8627 : node8504;
								assign node8504 = (inp[7]) ? node8564 : node8505;
									assign node8505 = (inp[4]) ? node8533 : node8506;
										assign node8506 = (inp[3]) ? node8520 : node8507;
											assign node8507 = (inp[14]) ? node8515 : node8508;
												assign node8508 = (inp[1]) ? node8512 : node8509;
													assign node8509 = (inp[9]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node8512 = (inp[8]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node8515 = (inp[8]) ? 15'b000000111111111 : node8516;
													assign node8516 = (inp[1]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node8520 = (inp[10]) ? node8526 : node8521;
												assign node8521 = (inp[1]) ? 15'b000000111111111 : node8522;
													assign node8522 = (inp[8]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node8526 = (inp[14]) ? node8530 : node8527;
													assign node8527 = (inp[9]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node8530 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node8533 = (inp[9]) ? node8549 : node8534;
											assign node8534 = (inp[14]) ? node8542 : node8535;
												assign node8535 = (inp[1]) ? node8539 : node8536;
													assign node8536 = (inp[10]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node8539 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node8542 = (inp[1]) ? node8546 : node8543;
													assign node8543 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node8546 = (inp[8]) ? 15'b000000000111111 : 15'b000000011111111;
											assign node8549 = (inp[10]) ? node8557 : node8550;
												assign node8550 = (inp[1]) ? node8554 : node8551;
													assign node8551 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node8554 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node8557 = (inp[8]) ? node8561 : node8558;
													assign node8558 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node8561 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node8564 = (inp[8]) ? node8596 : node8565;
										assign node8565 = (inp[14]) ? node8581 : node8566;
											assign node8566 = (inp[9]) ? node8574 : node8567;
												assign node8567 = (inp[4]) ? node8571 : node8568;
													assign node8568 = (inp[10]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node8571 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node8574 = (inp[10]) ? node8578 : node8575;
													assign node8575 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node8578 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node8581 = (inp[4]) ? node8589 : node8582;
												assign node8582 = (inp[10]) ? node8586 : node8583;
													assign node8583 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node8586 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node8589 = (inp[9]) ? node8593 : node8590;
													assign node8590 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node8593 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node8596 = (inp[9]) ? node8612 : node8597;
											assign node8597 = (inp[3]) ? node8605 : node8598;
												assign node8598 = (inp[4]) ? node8602 : node8599;
													assign node8599 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node8602 = (inp[14]) ? 15'b000000001111111 : 15'b000000001111111;
												assign node8605 = (inp[10]) ? node8609 : node8606;
													assign node8606 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node8609 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node8612 = (inp[4]) ? node8620 : node8613;
												assign node8613 = (inp[1]) ? node8617 : node8614;
													assign node8614 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node8617 = (inp[10]) ? 15'b000000000111111 : 15'b000000000111111;
												assign node8620 = (inp[14]) ? node8624 : node8621;
													assign node8621 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node8624 = (inp[1]) ? 15'b000000000011111 : 15'b000000000111111;
								assign node8627 = (inp[1]) ? node8689 : node8628;
									assign node8628 = (inp[4]) ? node8660 : node8629;
										assign node8629 = (inp[3]) ? node8645 : node8630;
											assign node8630 = (inp[9]) ? node8638 : node8631;
												assign node8631 = (inp[8]) ? node8635 : node8632;
													assign node8632 = (inp[7]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node8635 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node8638 = (inp[10]) ? node8642 : node8639;
													assign node8639 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node8642 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node8645 = (inp[10]) ? node8653 : node8646;
												assign node8646 = (inp[14]) ? node8650 : node8647;
													assign node8647 = (inp[8]) ? 15'b000000011111111 : 15'b000000011111111;
													assign node8650 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node8653 = (inp[14]) ? node8657 : node8654;
													assign node8654 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node8657 = (inp[9]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node8660 = (inp[14]) ? node8674 : node8661;
											assign node8661 = (inp[3]) ? node8667 : node8662;
												assign node8662 = (inp[10]) ? node8664 : 15'b000000111111111;
													assign node8664 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node8667 = (inp[7]) ? node8671 : node8668;
													assign node8668 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node8671 = (inp[9]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node8674 = (inp[3]) ? node8682 : node8675;
												assign node8675 = (inp[7]) ? node8679 : node8676;
													assign node8676 = (inp[9]) ? 15'b000000001111111 : 15'b000000001111111;
													assign node8679 = (inp[9]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node8682 = (inp[8]) ? node8686 : node8683;
													assign node8683 = (inp[10]) ? 15'b000000000011111 : 15'b000000001111111;
													assign node8686 = (inp[9]) ? 15'b000000000011111 : 15'b000000000011111;
									assign node8689 = (inp[8]) ? node8721 : node8690;
										assign node8690 = (inp[10]) ? node8706 : node8691;
											assign node8691 = (inp[4]) ? node8699 : node8692;
												assign node8692 = (inp[9]) ? node8696 : node8693;
													assign node8693 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node8696 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node8699 = (inp[7]) ? node8703 : node8700;
													assign node8700 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node8703 = (inp[9]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node8706 = (inp[9]) ? node8714 : node8707;
												assign node8707 = (inp[14]) ? node8711 : node8708;
													assign node8708 = (inp[7]) ? 15'b000000001111111 : 15'b000000111111111;
													assign node8711 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node8714 = (inp[7]) ? node8718 : node8715;
													assign node8715 = (inp[4]) ? 15'b000000000111111 : 15'b000000011111111;
													assign node8718 = (inp[4]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node8721 = (inp[10]) ? node8737 : node8722;
											assign node8722 = (inp[3]) ? node8730 : node8723;
												assign node8723 = (inp[4]) ? node8727 : node8724;
													assign node8724 = (inp[9]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node8727 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node8730 = (inp[7]) ? node8734 : node8731;
													assign node8731 = (inp[9]) ? 15'b000000000111111 : 15'b000000000111111;
													assign node8734 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node8737 = (inp[7]) ? node8745 : node8738;
												assign node8738 = (inp[9]) ? node8742 : node8739;
													assign node8739 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node8742 = (inp[3]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node8745 = (inp[9]) ? node8749 : node8746;
													assign node8746 = (inp[4]) ? 15'b000000000001111 : 15'b000000000111111;
													assign node8749 = (inp[14]) ? 15'b000000000001111 : 15'b000000000011111;
					assign node8752 = (inp[3]) ? node9238 : node8753;
						assign node8753 = (inp[9]) ? node8999 : node8754;
							assign node8754 = (inp[7]) ? node8872 : node8755;
								assign node8755 = (inp[12]) ? node8815 : node8756;
									assign node8756 = (inp[14]) ? node8786 : node8757;
										assign node8757 = (inp[10]) ? node8771 : node8758;
											assign node8758 = (inp[11]) ? node8766 : node8759;
												assign node8759 = (inp[5]) ? node8763 : node8760;
													assign node8760 = (inp[8]) ? 15'b000111111111111 : 15'b000111111111111;
													assign node8763 = (inp[8]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node8766 = (inp[1]) ? 15'b000000111111111 : node8767;
													assign node8767 = (inp[4]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node8771 = (inp[8]) ? node8779 : node8772;
												assign node8772 = (inp[5]) ? node8776 : node8773;
													assign node8773 = (inp[11]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node8776 = (inp[4]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node8779 = (inp[5]) ? node8783 : node8780;
													assign node8780 = (inp[4]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node8783 = (inp[1]) ? 15'b000000111111111 : 15'b000000111111111;
										assign node8786 = (inp[11]) ? node8800 : node8787;
											assign node8787 = (inp[5]) ? node8795 : node8788;
												assign node8788 = (inp[8]) ? node8792 : node8789;
													assign node8789 = (inp[4]) ? 15'b000001111111111 : 15'b000001111111111;
													assign node8792 = (inp[10]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node8795 = (inp[1]) ? 15'b000000011111111 : node8796;
													assign node8796 = (inp[4]) ? 15'b000000111111111 : 15'b000000111111111;
											assign node8800 = (inp[1]) ? node8808 : node8801;
												assign node8801 = (inp[8]) ? node8805 : node8802;
													assign node8802 = (inp[5]) ? 15'b000000111111111 : 15'b000000111111111;
													assign node8805 = (inp[5]) ? 15'b000000111111111 : 15'b000000111111111;
												assign node8808 = (inp[4]) ? node8812 : node8809;
													assign node8809 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node8812 = (inp[8]) ? 15'b000000001111111 : 15'b000000001111111;
									assign node8815 = (inp[10]) ? node8841 : node8816;
										assign node8816 = (inp[5]) ? node8832 : node8817;
											assign node8817 = (inp[4]) ? node8825 : node8818;
												assign node8818 = (inp[1]) ? node8822 : node8819;
													assign node8819 = (inp[14]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node8822 = (inp[8]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node8825 = (inp[8]) ? node8829 : node8826;
													assign node8826 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node8829 = (inp[14]) ? 15'b000000001111111 : 15'b000000111111111;
											assign node8832 = (inp[11]) ? node8834 : 15'b000000111111111;
												assign node8834 = (inp[14]) ? node8838 : node8835;
													assign node8835 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node8838 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node8841 = (inp[1]) ? node8857 : node8842;
											assign node8842 = (inp[11]) ? node8850 : node8843;
												assign node8843 = (inp[4]) ? node8847 : node8844;
													assign node8844 = (inp[8]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node8847 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node8850 = (inp[5]) ? node8854 : node8851;
													assign node8851 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node8854 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node8857 = (inp[4]) ? node8865 : node8858;
												assign node8858 = (inp[8]) ? node8862 : node8859;
													assign node8859 = (inp[11]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node8862 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node8865 = (inp[11]) ? node8869 : node8866;
													assign node8866 = (inp[8]) ? 15'b000000000111111 : 15'b000000011111111;
													assign node8869 = (inp[8]) ? 15'b000000000111111 : 15'b000000000111111;
								assign node8872 = (inp[4]) ? node8936 : node8873;
									assign node8873 = (inp[5]) ? node8905 : node8874;
										assign node8874 = (inp[1]) ? node8890 : node8875;
											assign node8875 = (inp[12]) ? node8883 : node8876;
												assign node8876 = (inp[10]) ? node8880 : node8877;
													assign node8877 = (inp[11]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node8880 = (inp[8]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node8883 = (inp[10]) ? node8887 : node8884;
													assign node8884 = (inp[11]) ? 15'b000000111111111 : 15'b000011111111111;
													assign node8887 = (inp[11]) ? 15'b000000001111111 : 15'b000000111111111;
											assign node8890 = (inp[12]) ? node8898 : node8891;
												assign node8891 = (inp[10]) ? node8895 : node8892;
													assign node8892 = (inp[11]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node8895 = (inp[8]) ? 15'b000000001111111 : 15'b000000111111111;
												assign node8898 = (inp[14]) ? node8902 : node8899;
													assign node8899 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node8902 = (inp[8]) ? 15'b000000001111111 : 15'b000000001111111;
										assign node8905 = (inp[1]) ? node8921 : node8906;
											assign node8906 = (inp[11]) ? node8914 : node8907;
												assign node8907 = (inp[12]) ? node8911 : node8908;
													assign node8908 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node8911 = (inp[14]) ? 15'b000000011111111 : 15'b000000011111111;
												assign node8914 = (inp[8]) ? node8918 : node8915;
													assign node8915 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node8918 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node8921 = (inp[14]) ? node8929 : node8922;
												assign node8922 = (inp[12]) ? node8926 : node8923;
													assign node8923 = (inp[11]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node8926 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node8929 = (inp[11]) ? node8933 : node8930;
													assign node8930 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node8933 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node8936 = (inp[5]) ? node8968 : node8937;
										assign node8937 = (inp[14]) ? node8953 : node8938;
											assign node8938 = (inp[8]) ? node8946 : node8939;
												assign node8939 = (inp[10]) ? node8943 : node8940;
													assign node8940 = (inp[1]) ? 15'b000000111111111 : 15'b000011111111111;
													assign node8943 = (inp[12]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node8946 = (inp[11]) ? node8950 : node8947;
													assign node8947 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node8950 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node8953 = (inp[12]) ? node8961 : node8954;
												assign node8954 = (inp[1]) ? node8958 : node8955;
													assign node8955 = (inp[8]) ? 15'b000000011111111 : 15'b000000011111111;
													assign node8958 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node8961 = (inp[10]) ? node8965 : node8962;
													assign node8962 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node8965 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node8968 = (inp[1]) ? node8984 : node8969;
											assign node8969 = (inp[11]) ? node8977 : node8970;
												assign node8970 = (inp[12]) ? node8974 : node8971;
													assign node8971 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node8974 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node8977 = (inp[12]) ? node8981 : node8978;
													assign node8978 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node8981 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node8984 = (inp[8]) ? node8992 : node8985;
												assign node8985 = (inp[12]) ? node8989 : node8986;
													assign node8986 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node8989 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node8992 = (inp[11]) ? node8996 : node8993;
													assign node8993 = (inp[12]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node8996 = (inp[10]) ? 15'b000000000011111 : 15'b000000000111111;
							assign node8999 = (inp[12]) ? node9123 : node9000;
								assign node9000 = (inp[1]) ? node9064 : node9001;
									assign node9001 = (inp[8]) ? node9033 : node9002;
										assign node9002 = (inp[10]) ? node9018 : node9003;
											assign node9003 = (inp[5]) ? node9011 : node9004;
												assign node9004 = (inp[7]) ? node9008 : node9005;
													assign node9005 = (inp[4]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node9008 = (inp[4]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node9011 = (inp[11]) ? node9015 : node9012;
													assign node9012 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node9015 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node9018 = (inp[4]) ? node9026 : node9019;
												assign node9019 = (inp[14]) ? node9023 : node9020;
													assign node9020 = (inp[7]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node9023 = (inp[11]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node9026 = (inp[7]) ? node9030 : node9027;
													assign node9027 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node9030 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node9033 = (inp[4]) ? node9049 : node9034;
											assign node9034 = (inp[11]) ? node9042 : node9035;
												assign node9035 = (inp[5]) ? node9039 : node9036;
													assign node9036 = (inp[10]) ? 15'b000000111111111 : 15'b000011111111111;
													assign node9039 = (inp[7]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node9042 = (inp[10]) ? node9046 : node9043;
													assign node9043 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node9046 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node9049 = (inp[10]) ? node9057 : node9050;
												assign node9050 = (inp[5]) ? node9054 : node9051;
													assign node9051 = (inp[7]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node9054 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node9057 = (inp[5]) ? node9061 : node9058;
													assign node9058 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node9061 = (inp[7]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node9064 = (inp[5]) ? node9094 : node9065;
										assign node9065 = (inp[7]) ? node9079 : node9066;
											assign node9066 = (inp[8]) ? node9072 : node9067;
												assign node9067 = (inp[14]) ? 15'b000000111111111 : node9068;
													assign node9068 = (inp[11]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node9072 = (inp[10]) ? node9076 : node9073;
													assign node9073 = (inp[11]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node9076 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node9079 = (inp[4]) ? node9087 : node9080;
												assign node9080 = (inp[10]) ? node9084 : node9081;
													assign node9081 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node9084 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node9087 = (inp[8]) ? node9091 : node9088;
													assign node9088 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node9091 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node9094 = (inp[14]) ? node9108 : node9095;
											assign node9095 = (inp[10]) ? node9103 : node9096;
												assign node9096 = (inp[8]) ? node9100 : node9097;
													assign node9097 = (inp[4]) ? 15'b000000011111111 : 15'b000001111111111;
													assign node9100 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node9103 = (inp[4]) ? node9105 : 15'b000000001111111;
													assign node9105 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node9108 = (inp[11]) ? node9116 : node9109;
												assign node9109 = (inp[4]) ? node9113 : node9110;
													assign node9110 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node9113 = (inp[7]) ? 15'b000000000011111 : 15'b000000001111111;
												assign node9116 = (inp[8]) ? node9120 : node9117;
													assign node9117 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node9120 = (inp[10]) ? 15'b000000000011111 : 15'b000000000111111;
								assign node9123 = (inp[8]) ? node9177 : node9124;
									assign node9124 = (inp[5]) ? node9148 : node9125;
										assign node9125 = (inp[7]) ? node9133 : node9126;
											assign node9126 = (inp[1]) ? node9128 : 15'b000000111111111;
												assign node9128 = (inp[14]) ? node9130 : 15'b000000111111111;
													assign node9130 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node9133 = (inp[10]) ? node9141 : node9134;
												assign node9134 = (inp[14]) ? node9138 : node9135;
													assign node9135 = (inp[1]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node9138 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node9141 = (inp[1]) ? node9145 : node9142;
													assign node9142 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node9145 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node9148 = (inp[10]) ? node9164 : node9149;
											assign node9149 = (inp[4]) ? node9157 : node9150;
												assign node9150 = (inp[1]) ? node9154 : node9151;
													assign node9151 = (inp[14]) ? 15'b000000011111111 : 15'b000000011111111;
													assign node9154 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node9157 = (inp[14]) ? node9161 : node9158;
													assign node9158 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node9161 = (inp[1]) ? 15'b000000000111111 : 15'b000000000111111;
											assign node9164 = (inp[14]) ? node9172 : node9165;
												assign node9165 = (inp[11]) ? node9169 : node9166;
													assign node9166 = (inp[7]) ? 15'b000000001111111 : 15'b000000001111111;
													assign node9169 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node9172 = (inp[4]) ? node9174 : 15'b000000001111111;
													assign node9174 = (inp[1]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node9177 = (inp[7]) ? node9209 : node9178;
										assign node9178 = (inp[1]) ? node9194 : node9179;
											assign node9179 = (inp[11]) ? node9187 : node9180;
												assign node9180 = (inp[10]) ? node9184 : node9181;
													assign node9181 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node9184 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node9187 = (inp[5]) ? node9191 : node9188;
													assign node9188 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node9191 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node9194 = (inp[5]) ? node9202 : node9195;
												assign node9195 = (inp[14]) ? node9199 : node9196;
													assign node9196 = (inp[11]) ? 15'b000000001111111 : 15'b000000001111111;
													assign node9199 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node9202 = (inp[10]) ? node9206 : node9203;
													assign node9203 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node9206 = (inp[4]) ? 15'b000000000011111 : 15'b000000000011111;
										assign node9209 = (inp[10]) ? node9225 : node9210;
											assign node9210 = (inp[14]) ? node9218 : node9211;
												assign node9211 = (inp[4]) ? node9215 : node9212;
													assign node9212 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node9215 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node9218 = (inp[4]) ? node9222 : node9219;
													assign node9219 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node9222 = (inp[11]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node9225 = (inp[5]) ? node9231 : node9226;
												assign node9226 = (inp[4]) ? node9228 : 15'b000000000111111;
													assign node9228 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node9231 = (inp[1]) ? node9235 : node9232;
													assign node9232 = (inp[11]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node9235 = (inp[4]) ? 15'b000000000000111 : 15'b000000000011111;
						assign node9238 = (inp[10]) ? node9476 : node9239;
							assign node9239 = (inp[5]) ? node9359 : node9240;
								assign node9240 = (inp[11]) ? node9300 : node9241;
									assign node9241 = (inp[9]) ? node9269 : node9242;
										assign node9242 = (inp[4]) ? node9256 : node9243;
											assign node9243 = (inp[1]) ? node9249 : node9244;
												assign node9244 = (inp[14]) ? 15'b000001111111111 : node9245;
													assign node9245 = (inp[7]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node9249 = (inp[8]) ? node9253 : node9250;
													assign node9250 = (inp[12]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node9253 = (inp[12]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node9256 = (inp[12]) ? node9264 : node9257;
												assign node9257 = (inp[1]) ? node9261 : node9258;
													assign node9258 = (inp[7]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node9261 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node9264 = (inp[8]) ? 15'b000000001111111 : node9265;
													assign node9265 = (inp[7]) ? 15'b000000001111111 : 15'b000000111111111;
										assign node9269 = (inp[8]) ? node9285 : node9270;
											assign node9270 = (inp[7]) ? node9278 : node9271;
												assign node9271 = (inp[12]) ? node9275 : node9272;
													assign node9272 = (inp[1]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node9275 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node9278 = (inp[4]) ? node9282 : node9279;
													assign node9279 = (inp[1]) ? 15'b000000001111111 : 15'b000000111111111;
													assign node9282 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node9285 = (inp[12]) ? node9293 : node9286;
												assign node9286 = (inp[1]) ? node9290 : node9287;
													assign node9287 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node9290 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node9293 = (inp[1]) ? node9297 : node9294;
													assign node9294 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node9297 = (inp[7]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node9300 = (inp[4]) ? node9328 : node9301;
										assign node9301 = (inp[9]) ? node9315 : node9302;
											assign node9302 = (inp[1]) ? node9308 : node9303;
												assign node9303 = (inp[8]) ? 15'b000000111111111 : node9304;
													assign node9304 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node9308 = (inp[14]) ? node9312 : node9309;
													assign node9309 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node9312 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node9315 = (inp[1]) ? node9323 : node9316;
												assign node9316 = (inp[14]) ? node9320 : node9317;
													assign node9317 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node9320 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node9323 = (inp[14]) ? node9325 : 15'b000000001111111;
													assign node9325 = (inp[12]) ? 15'b000000000011111 : 15'b000000001111111;
										assign node9328 = (inp[12]) ? node9344 : node9329;
											assign node9329 = (inp[8]) ? node9337 : node9330;
												assign node9330 = (inp[14]) ? node9334 : node9331;
													assign node9331 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node9334 = (inp[1]) ? 15'b000000001111111 : 15'b000000001111111;
												assign node9337 = (inp[9]) ? node9341 : node9338;
													assign node9338 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node9341 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node9344 = (inp[7]) ? node9352 : node9345;
												assign node9345 = (inp[14]) ? node9349 : node9346;
													assign node9346 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node9349 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node9352 = (inp[9]) ? node9356 : node9353;
													assign node9353 = (inp[14]) ? 15'b000000000111111 : 15'b000000000111111;
													assign node9356 = (inp[1]) ? 15'b000000000011111 : 15'b000000000111111;
								assign node9359 = (inp[1]) ? node9419 : node9360;
									assign node9360 = (inp[11]) ? node9390 : node9361;
										assign node9361 = (inp[8]) ? node9375 : node9362;
											assign node9362 = (inp[12]) ? node9370 : node9363;
												assign node9363 = (inp[7]) ? node9367 : node9364;
													assign node9364 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node9367 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node9370 = (inp[14]) ? node9372 : 15'b000000111111111;
													assign node9372 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node9375 = (inp[7]) ? node9383 : node9376;
												assign node9376 = (inp[14]) ? node9380 : node9377;
													assign node9377 = (inp[9]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node9380 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node9383 = (inp[9]) ? node9387 : node9384;
													assign node9384 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node9387 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node9390 = (inp[4]) ? node9406 : node9391;
											assign node9391 = (inp[7]) ? node9399 : node9392;
												assign node9392 = (inp[12]) ? node9396 : node9393;
													assign node9393 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node9396 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node9399 = (inp[14]) ? node9403 : node9400;
													assign node9400 = (inp[9]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node9403 = (inp[9]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node9406 = (inp[9]) ? node9414 : node9407;
												assign node9407 = (inp[14]) ? node9411 : node9408;
													assign node9408 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node9411 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node9414 = (inp[7]) ? node9416 : 15'b000000000111111;
													assign node9416 = (inp[12]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node9419 = (inp[4]) ? node9447 : node9420;
										assign node9420 = (inp[9]) ? node9432 : node9421;
											assign node9421 = (inp[14]) ? node9427 : node9422;
												assign node9422 = (inp[7]) ? 15'b000000011111111 : node9423;
													assign node9423 = (inp[12]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node9427 = (inp[12]) ? node9429 : 15'b000000011111111;
													assign node9429 = (inp[7]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node9432 = (inp[11]) ? node9440 : node9433;
												assign node9433 = (inp[12]) ? node9437 : node9434;
													assign node9434 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node9437 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node9440 = (inp[14]) ? node9444 : node9441;
													assign node9441 = (inp[12]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node9444 = (inp[7]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node9447 = (inp[8]) ? node9461 : node9448;
											assign node9448 = (inp[9]) ? node9454 : node9449;
												assign node9449 = (inp[7]) ? node9451 : 15'b000000011111111;
													assign node9451 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node9454 = (inp[12]) ? node9458 : node9455;
													assign node9455 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node9458 = (inp[11]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node9461 = (inp[14]) ? node9469 : node9462;
												assign node9462 = (inp[9]) ? node9466 : node9463;
													assign node9463 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node9466 = (inp[7]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node9469 = (inp[12]) ? node9473 : node9470;
													assign node9470 = (inp[9]) ? 15'b000000000011111 : 15'b000000000011111;
													assign node9473 = (inp[11]) ? 15'b000000000001111 : 15'b000000000011111;
							assign node9476 = (inp[4]) ? node9602 : node9477;
								assign node9477 = (inp[1]) ? node9541 : node9478;
									assign node9478 = (inp[8]) ? node9510 : node9479;
										assign node9479 = (inp[14]) ? node9495 : node9480;
											assign node9480 = (inp[12]) ? node9488 : node9481;
												assign node9481 = (inp[11]) ? node9485 : node9482;
													assign node9482 = (inp[7]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node9485 = (inp[9]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node9488 = (inp[5]) ? node9492 : node9489;
													assign node9489 = (inp[7]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node9492 = (inp[9]) ? 15'b000000000111111 : 15'b000000011111111;
											assign node9495 = (inp[9]) ? node9503 : node9496;
												assign node9496 = (inp[12]) ? node9500 : node9497;
													assign node9497 = (inp[11]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node9500 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node9503 = (inp[5]) ? node9507 : node9504;
													assign node9504 = (inp[7]) ? 15'b000000001111111 : 15'b000000111111111;
													assign node9507 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node9510 = (inp[5]) ? node9526 : node9511;
											assign node9511 = (inp[9]) ? node9519 : node9512;
												assign node9512 = (inp[11]) ? node9516 : node9513;
													assign node9513 = (inp[14]) ? 15'b000000001111111 : 15'b000000111111111;
													assign node9516 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node9519 = (inp[7]) ? node9523 : node9520;
													assign node9520 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node9523 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node9526 = (inp[9]) ? node9534 : node9527;
												assign node9527 = (inp[12]) ? node9531 : node9528;
													assign node9528 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node9531 = (inp[7]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node9534 = (inp[11]) ? node9538 : node9535;
													assign node9535 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node9538 = (inp[12]) ? 15'b000000000001111 : 15'b000000000111111;
									assign node9541 = (inp[12]) ? node9571 : node9542;
										assign node9542 = (inp[5]) ? node9556 : node9543;
											assign node9543 = (inp[7]) ? node9549 : node9544;
												assign node9544 = (inp[8]) ? node9546 : 15'b000000011111111;
													assign node9546 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node9549 = (inp[8]) ? node9553 : node9550;
													assign node9550 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node9553 = (inp[14]) ? 15'b000000000011111 : 15'b000000001111111;
											assign node9556 = (inp[11]) ? node9564 : node9557;
												assign node9557 = (inp[7]) ? node9561 : node9558;
													assign node9558 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node9561 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node9564 = (inp[9]) ? node9568 : node9565;
													assign node9565 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node9568 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node9571 = (inp[14]) ? node9587 : node9572;
											assign node9572 = (inp[11]) ? node9580 : node9573;
												assign node9573 = (inp[5]) ? node9577 : node9574;
													assign node9574 = (inp[7]) ? 15'b000000001111111 : 15'b000000001111111;
													assign node9577 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node9580 = (inp[9]) ? node9584 : node9581;
													assign node9581 = (inp[7]) ? 15'b000000000111111 : 15'b000000000111111;
													assign node9584 = (inp[5]) ? 15'b000000000001111 : 15'b000000000111111;
											assign node9587 = (inp[11]) ? node9595 : node9588;
												assign node9588 = (inp[9]) ? node9592 : node9589;
													assign node9589 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node9592 = (inp[8]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node9595 = (inp[5]) ? node9599 : node9596;
													assign node9596 = (inp[8]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node9599 = (inp[8]) ? 15'b000000000001111 : 15'b000000000011111;
								assign node9602 = (inp[7]) ? node9666 : node9603;
									assign node9603 = (inp[14]) ? node9635 : node9604;
										assign node9604 = (inp[11]) ? node9620 : node9605;
											assign node9605 = (inp[12]) ? node9613 : node9606;
												assign node9606 = (inp[5]) ? node9610 : node9607;
													assign node9607 = (inp[1]) ? 15'b000000011111111 : 15'b000000011111111;
													assign node9610 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node9613 = (inp[9]) ? node9617 : node9614;
													assign node9614 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node9617 = (inp[5]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node9620 = (inp[9]) ? node9628 : node9621;
												assign node9621 = (inp[1]) ? node9625 : node9622;
													assign node9622 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node9625 = (inp[5]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node9628 = (inp[8]) ? node9632 : node9629;
													assign node9629 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node9632 = (inp[1]) ? 15'b000000000001111 : 15'b000000000111111;
										assign node9635 = (inp[8]) ? node9651 : node9636;
											assign node9636 = (inp[5]) ? node9644 : node9637;
												assign node9637 = (inp[12]) ? node9641 : node9638;
													assign node9638 = (inp[9]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node9641 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node9644 = (inp[11]) ? node9648 : node9645;
													assign node9645 = (inp[1]) ? 15'b000000000111111 : 15'b000000000111111;
													assign node9648 = (inp[1]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node9651 = (inp[11]) ? node9659 : node9652;
												assign node9652 = (inp[12]) ? node9656 : node9653;
													assign node9653 = (inp[5]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node9656 = (inp[5]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node9659 = (inp[1]) ? node9663 : node9660;
													assign node9660 = (inp[5]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node9663 = (inp[5]) ? 15'b000000000001111 : 15'b000000000011111;
									assign node9666 = (inp[1]) ? node9698 : node9667;
										assign node9667 = (inp[11]) ? node9683 : node9668;
											assign node9668 = (inp[9]) ? node9676 : node9669;
												assign node9669 = (inp[5]) ? node9673 : node9670;
													assign node9670 = (inp[12]) ? 15'b000000001111111 : 15'b000000001111111;
													assign node9673 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node9676 = (inp[8]) ? node9680 : node9677;
													assign node9677 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node9680 = (inp[5]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node9683 = (inp[9]) ? node9691 : node9684;
												assign node9684 = (inp[12]) ? node9688 : node9685;
													assign node9685 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node9688 = (inp[5]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node9691 = (inp[12]) ? node9695 : node9692;
													assign node9692 = (inp[14]) ? 15'b000000000011111 : 15'b000000000011111;
													assign node9695 = (inp[5]) ? 15'b000000000001111 : 15'b000000000011111;
										assign node9698 = (inp[8]) ? node9708 : node9699;
											assign node9699 = (inp[9]) ? node9701 : 15'b000000000111111;
												assign node9701 = (inp[14]) ? node9705 : node9702;
													assign node9702 = (inp[5]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node9705 = (inp[11]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node9708 = (inp[5]) ? node9716 : node9709;
												assign node9709 = (inp[14]) ? node9713 : node9710;
													assign node9710 = (inp[9]) ? 15'b000000000011111 : 15'b000000001111111;
													assign node9713 = (inp[9]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node9716 = (inp[12]) ? node9720 : node9717;
													assign node9717 = (inp[9]) ? 15'b000000000001111 : 15'b000000000001111;
													assign node9720 = (inp[14]) ? 15'b000000000000111 : 15'b000000000001111;
				assign node9723 = (inp[10]) ? node10679 : node9724;
					assign node9724 = (inp[1]) ? node10200 : node9725;
						assign node9725 = (inp[8]) ? node9961 : node9726;
							assign node9726 = (inp[12]) ? node9844 : node9727;
								assign node9727 = (inp[3]) ? node9787 : node9728;
									assign node9728 = (inp[2]) ? node9756 : node9729;
										assign node9729 = (inp[5]) ? node9743 : node9730;
											assign node9730 = (inp[4]) ? node9738 : node9731;
												assign node9731 = (inp[11]) ? node9735 : node9732;
													assign node9732 = (inp[7]) ? 15'b000011111111111 : 15'b000111111111111;
													assign node9735 = (inp[14]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node9738 = (inp[14]) ? 15'b000001111111111 : node9739;
													assign node9739 = (inp[9]) ? 15'b000001111111111 : 15'b000001111111111;
											assign node9743 = (inp[14]) ? node9751 : node9744;
												assign node9744 = (inp[4]) ? node9748 : node9745;
													assign node9745 = (inp[11]) ? 15'b000001111111111 : 15'b000001111111111;
													assign node9748 = (inp[11]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node9751 = (inp[7]) ? 15'b000000111111111 : node9752;
													assign node9752 = (inp[4]) ? 15'b000000111111111 : 15'b000011111111111;
										assign node9756 = (inp[14]) ? node9772 : node9757;
											assign node9757 = (inp[11]) ? node9765 : node9758;
												assign node9758 = (inp[4]) ? node9762 : node9759;
													assign node9759 = (inp[7]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node9762 = (inp[9]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node9765 = (inp[4]) ? node9769 : node9766;
													assign node9766 = (inp[7]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node9769 = (inp[9]) ? 15'b000000001111111 : 15'b000000111111111;
											assign node9772 = (inp[5]) ? node9780 : node9773;
												assign node9773 = (inp[9]) ? node9777 : node9774;
													assign node9774 = (inp[7]) ? 15'b000000111111111 : 15'b000000111111111;
													assign node9777 = (inp[11]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node9780 = (inp[11]) ? node9784 : node9781;
													assign node9781 = (inp[7]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node9784 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node9787 = (inp[14]) ? node9817 : node9788;
										assign node9788 = (inp[9]) ? node9804 : node9789;
											assign node9789 = (inp[2]) ? node9797 : node9790;
												assign node9790 = (inp[7]) ? node9794 : node9791;
													assign node9791 = (inp[5]) ? 15'b000000111111111 : 15'b000011111111111;
													assign node9794 = (inp[11]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node9797 = (inp[11]) ? node9801 : node9798;
													assign node9798 = (inp[4]) ? 15'b000000011111111 : 15'b000001111111111;
													assign node9801 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node9804 = (inp[4]) ? node9810 : node9805;
												assign node9805 = (inp[11]) ? node9807 : 15'b000000111111111;
													assign node9807 = (inp[7]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node9810 = (inp[2]) ? node9814 : node9811;
													assign node9811 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node9814 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node9817 = (inp[7]) ? node9833 : node9818;
											assign node9818 = (inp[4]) ? node9826 : node9819;
												assign node9819 = (inp[11]) ? node9823 : node9820;
													assign node9820 = (inp[5]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node9823 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node9826 = (inp[2]) ? node9830 : node9827;
													assign node9827 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node9830 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node9833 = (inp[9]) ? node9841 : node9834;
												assign node9834 = (inp[2]) ? node9838 : node9835;
													assign node9835 = (inp[5]) ? 15'b000000001111111 : 15'b000000111111111;
													assign node9838 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node9841 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
								assign node9844 = (inp[11]) ? node9902 : node9845;
									assign node9845 = (inp[3]) ? node9875 : node9846;
										assign node9846 = (inp[14]) ? node9860 : node9847;
											assign node9847 = (inp[4]) ? node9853 : node9848;
												assign node9848 = (inp[7]) ? node9850 : 15'b000011111111111;
													assign node9850 = (inp[9]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node9853 = (inp[2]) ? node9857 : node9854;
													assign node9854 = (inp[5]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node9857 = (inp[7]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node9860 = (inp[5]) ? node9868 : node9861;
												assign node9861 = (inp[2]) ? node9865 : node9862;
													assign node9862 = (inp[7]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node9865 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node9868 = (inp[7]) ? node9872 : node9869;
													assign node9869 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node9872 = (inp[9]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node9875 = (inp[7]) ? node9887 : node9876;
											assign node9876 = (inp[9]) ? node9884 : node9877;
												assign node9877 = (inp[4]) ? node9881 : node9878;
													assign node9878 = (inp[2]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node9881 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node9884 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node9887 = (inp[2]) ? node9895 : node9888;
												assign node9888 = (inp[14]) ? node9892 : node9889;
													assign node9889 = (inp[9]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node9892 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node9895 = (inp[4]) ? node9899 : node9896;
													assign node9896 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node9899 = (inp[14]) ? 15'b000000000111111 : 15'b000000000111111;
									assign node9902 = (inp[5]) ? node9932 : node9903;
										assign node9903 = (inp[7]) ? node9917 : node9904;
											assign node9904 = (inp[14]) ? node9910 : node9905;
												assign node9905 = (inp[9]) ? node9907 : 15'b000001111111111;
													assign node9907 = (inp[4]) ? 15'b000000111111111 : 15'b000000111111111;
												assign node9910 = (inp[9]) ? node9914 : node9911;
													assign node9911 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node9914 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node9917 = (inp[3]) ? node9925 : node9918;
												assign node9918 = (inp[4]) ? node9922 : node9919;
													assign node9919 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node9922 = (inp[9]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node9925 = (inp[2]) ? node9929 : node9926;
													assign node9926 = (inp[9]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node9929 = (inp[9]) ? 15'b000000000111111 : 15'b000000000111111;
										assign node9932 = (inp[2]) ? node9946 : node9933;
											assign node9933 = (inp[9]) ? node9941 : node9934;
												assign node9934 = (inp[4]) ? node9938 : node9935;
													assign node9935 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node9938 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node9941 = (inp[14]) ? 15'b000000000111111 : node9942;
													assign node9942 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node9946 = (inp[7]) ? node9954 : node9947;
												assign node9947 = (inp[14]) ? node9951 : node9948;
													assign node9948 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node9951 = (inp[9]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node9954 = (inp[3]) ? node9958 : node9955;
													assign node9955 = (inp[9]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node9958 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
							assign node9961 = (inp[11]) ? node10081 : node9962;
								assign node9962 = (inp[2]) ? node10024 : node9963;
									assign node9963 = (inp[4]) ? node9995 : node9964;
										assign node9964 = (inp[14]) ? node9980 : node9965;
											assign node9965 = (inp[12]) ? node9973 : node9966;
												assign node9966 = (inp[9]) ? node9970 : node9967;
													assign node9967 = (inp[5]) ? 15'b000000111111111 : 15'b000011111111111;
													assign node9970 = (inp[3]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node9973 = (inp[7]) ? node9977 : node9974;
													assign node9974 = (inp[5]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node9977 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node9980 = (inp[5]) ? node9988 : node9981;
												assign node9981 = (inp[3]) ? node9985 : node9982;
													assign node9982 = (inp[7]) ? 15'b000000111111111 : 15'b000011111111111;
													assign node9985 = (inp[7]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node9988 = (inp[12]) ? node9992 : node9989;
													assign node9989 = (inp[9]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node9992 = (inp[9]) ? 15'b000000000111111 : 15'b000000011111111;
										assign node9995 = (inp[14]) ? node10009 : node9996;
											assign node9996 = (inp[12]) ? node10002 : node9997;
												assign node9997 = (inp[5]) ? node9999 : 15'b000001111111111;
													assign node9999 = (inp[9]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node10002 = (inp[5]) ? node10006 : node10003;
													assign node10003 = (inp[7]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node10006 = (inp[9]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node10009 = (inp[3]) ? node10017 : node10010;
												assign node10010 = (inp[5]) ? node10014 : node10011;
													assign node10011 = (inp[12]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node10014 = (inp[7]) ? 15'b000000001111111 : 15'b000000001111111;
												assign node10017 = (inp[9]) ? node10021 : node10018;
													assign node10018 = (inp[5]) ? 15'b000000001111111 : 15'b000000001111111;
													assign node10021 = (inp[5]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node10024 = (inp[12]) ? node10052 : node10025;
										assign node10025 = (inp[9]) ? node10039 : node10026;
											assign node10026 = (inp[7]) ? node10034 : node10027;
												assign node10027 = (inp[14]) ? node10031 : node10028;
													assign node10028 = (inp[5]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node10031 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node10034 = (inp[4]) ? 15'b000000001111111 : node10035;
													assign node10035 = (inp[14]) ? 15'b000000001111111 : 15'b000000111111111;
											assign node10039 = (inp[7]) ? node10045 : node10040;
												assign node10040 = (inp[3]) ? node10042 : 15'b000000011111111;
													assign node10042 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node10045 = (inp[5]) ? node10049 : node10046;
													assign node10046 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node10049 = (inp[14]) ? 15'b000000000011111 : 15'b000000001111111;
										assign node10052 = (inp[5]) ? node10066 : node10053;
											assign node10053 = (inp[3]) ? node10061 : node10054;
												assign node10054 = (inp[14]) ? node10058 : node10055;
													assign node10055 = (inp[7]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node10058 = (inp[9]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node10061 = (inp[9]) ? node10063 : 15'b000000001111111;
													assign node10063 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node10066 = (inp[9]) ? node10074 : node10067;
												assign node10067 = (inp[14]) ? node10071 : node10068;
													assign node10068 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node10071 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node10074 = (inp[3]) ? node10078 : node10075;
													assign node10075 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node10078 = (inp[4]) ? 15'b000000000011111 : 15'b000000000111111;
								assign node10081 = (inp[9]) ? node10139 : node10082;
									assign node10082 = (inp[5]) ? node10112 : node10083;
										assign node10083 = (inp[14]) ? node10097 : node10084;
											assign node10084 = (inp[12]) ? node10090 : node10085;
												assign node10085 = (inp[3]) ? 15'b000000111111111 : node10086;
													assign node10086 = (inp[2]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node10090 = (inp[7]) ? node10094 : node10091;
													assign node10091 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node10094 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node10097 = (inp[4]) ? node10105 : node10098;
												assign node10098 = (inp[3]) ? node10102 : node10099;
													assign node10099 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node10102 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node10105 = (inp[7]) ? node10109 : node10106;
													assign node10106 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node10109 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node10112 = (inp[7]) ? node10126 : node10113;
											assign node10113 = (inp[4]) ? node10121 : node10114;
												assign node10114 = (inp[3]) ? node10118 : node10115;
													assign node10115 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node10118 = (inp[2]) ? 15'b000000001111111 : 15'b000000001111111;
												assign node10121 = (inp[12]) ? node10123 : 15'b000000001111111;
													assign node10123 = (inp[2]) ? 15'b000000001111111 : 15'b000000001111111;
											assign node10126 = (inp[2]) ? node10134 : node10127;
												assign node10127 = (inp[3]) ? node10131 : node10128;
													assign node10128 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node10131 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node10134 = (inp[12]) ? node10136 : 15'b000000000111111;
													assign node10136 = (inp[4]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node10139 = (inp[14]) ? node10171 : node10140;
										assign node10140 = (inp[4]) ? node10156 : node10141;
											assign node10141 = (inp[5]) ? node10149 : node10142;
												assign node10142 = (inp[3]) ? node10146 : node10143;
													assign node10143 = (inp[7]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node10146 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node10149 = (inp[2]) ? node10153 : node10150;
													assign node10150 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node10153 = (inp[3]) ? 15'b000000000111111 : 15'b000000000111111;
											assign node10156 = (inp[3]) ? node10164 : node10157;
												assign node10157 = (inp[5]) ? node10161 : node10158;
													assign node10158 = (inp[12]) ? 15'b000000011111111 : 15'b000000001111111;
													assign node10161 = (inp[7]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node10164 = (inp[2]) ? node10168 : node10165;
													assign node10165 = (inp[12]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node10168 = (inp[5]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node10171 = (inp[3]) ? node10187 : node10172;
											assign node10172 = (inp[12]) ? node10180 : node10173;
												assign node10173 = (inp[2]) ? node10177 : node10174;
													assign node10174 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node10177 = (inp[5]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node10180 = (inp[7]) ? node10184 : node10181;
													assign node10181 = (inp[5]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node10184 = (inp[2]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node10187 = (inp[12]) ? node10195 : node10188;
												assign node10188 = (inp[5]) ? node10192 : node10189;
													assign node10189 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node10192 = (inp[2]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node10195 = (inp[5]) ? 15'b000000000011111 : node10196;
													assign node10196 = (inp[7]) ? 15'b000000000011111 : 15'b000000000111111;
						assign node10200 = (inp[12]) ? node10440 : node10201;
							assign node10201 = (inp[5]) ? node10321 : node10202;
								assign node10202 = (inp[4]) ? node10260 : node10203;
									assign node10203 = (inp[14]) ? node10231 : node10204;
										assign node10204 = (inp[9]) ? node10218 : node10205;
											assign node10205 = (inp[2]) ? node10211 : node10206;
												assign node10206 = (inp[3]) ? 15'b000001111111111 : node10207;
													assign node10207 = (inp[11]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node10211 = (inp[8]) ? node10215 : node10212;
													assign node10212 = (inp[11]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node10215 = (inp[7]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node10218 = (inp[3]) ? node10224 : node10219;
												assign node10219 = (inp[11]) ? 15'b000000111111111 : node10220;
													assign node10220 = (inp[7]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node10224 = (inp[7]) ? node10228 : node10225;
													assign node10225 = (inp[11]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node10228 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node10231 = (inp[2]) ? node10247 : node10232;
											assign node10232 = (inp[3]) ? node10240 : node10233;
												assign node10233 = (inp[8]) ? node10237 : node10234;
													assign node10234 = (inp[9]) ? 15'b000000111111111 : 15'b000000111111111;
													assign node10237 = (inp[9]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node10240 = (inp[7]) ? node10244 : node10241;
													assign node10241 = (inp[11]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node10244 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node10247 = (inp[7]) ? node10253 : node10248;
												assign node10248 = (inp[3]) ? node10250 : 15'b000000111111111;
													assign node10250 = (inp[9]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node10253 = (inp[8]) ? node10257 : node10254;
													assign node10254 = (inp[9]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node10257 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node10260 = (inp[7]) ? node10290 : node10261;
										assign node10261 = (inp[2]) ? node10277 : node10262;
											assign node10262 = (inp[3]) ? node10270 : node10263;
												assign node10263 = (inp[8]) ? node10267 : node10264;
													assign node10264 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node10267 = (inp[11]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node10270 = (inp[9]) ? node10274 : node10271;
													assign node10271 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node10274 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node10277 = (inp[8]) ? node10285 : node10278;
												assign node10278 = (inp[11]) ? node10282 : node10279;
													assign node10279 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node10282 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node10285 = (inp[11]) ? node10287 : 15'b000000001111111;
													assign node10287 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node10290 = (inp[3]) ? node10306 : node10291;
											assign node10291 = (inp[14]) ? node10299 : node10292;
												assign node10292 = (inp[8]) ? node10296 : node10293;
													assign node10293 = (inp[11]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node10296 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node10299 = (inp[8]) ? node10303 : node10300;
													assign node10300 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node10303 = (inp[9]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node10306 = (inp[2]) ? node10314 : node10307;
												assign node10307 = (inp[9]) ? node10311 : node10308;
													assign node10308 = (inp[14]) ? 15'b000000001111111 : 15'b000000001111111;
													assign node10311 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node10314 = (inp[14]) ? node10318 : node10315;
													assign node10315 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node10318 = (inp[11]) ? 15'b000000000011111 : 15'b000000000111111;
								assign node10321 = (inp[2]) ? node10379 : node10322;
									assign node10322 = (inp[3]) ? node10350 : node10323;
										assign node10323 = (inp[7]) ? node10337 : node10324;
											assign node10324 = (inp[8]) ? node10332 : node10325;
												assign node10325 = (inp[11]) ? node10329 : node10326;
													assign node10326 = (inp[9]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node10329 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node10332 = (inp[4]) ? 15'b000000011111111 : node10333;
													assign node10333 = (inp[11]) ? 15'b000000011111111 : 15'b000000011111111;
											assign node10337 = (inp[14]) ? node10345 : node10338;
												assign node10338 = (inp[11]) ? node10342 : node10339;
													assign node10339 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node10342 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node10345 = (inp[4]) ? 15'b000000001111111 : node10346;
													assign node10346 = (inp[9]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node10350 = (inp[14]) ? node10364 : node10351;
											assign node10351 = (inp[4]) ? node10357 : node10352;
												assign node10352 = (inp[11]) ? node10354 : 15'b000000011111111;
													assign node10354 = (inp[9]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node10357 = (inp[8]) ? node10361 : node10358;
													assign node10358 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node10361 = (inp[7]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node10364 = (inp[8]) ? node10372 : node10365;
												assign node10365 = (inp[4]) ? node10369 : node10366;
													assign node10366 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node10369 = (inp[7]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node10372 = (inp[7]) ? node10376 : node10373;
													assign node10373 = (inp[11]) ? 15'b000000000111111 : 15'b000000000111111;
													assign node10376 = (inp[9]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node10379 = (inp[9]) ? node10411 : node10380;
										assign node10380 = (inp[7]) ? node10396 : node10381;
											assign node10381 = (inp[14]) ? node10389 : node10382;
												assign node10382 = (inp[3]) ? node10386 : node10383;
													assign node10383 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node10386 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node10389 = (inp[4]) ? node10393 : node10390;
													assign node10390 = (inp[11]) ? 15'b000000001111111 : 15'b000000001111111;
													assign node10393 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node10396 = (inp[8]) ? node10404 : node10397;
												assign node10397 = (inp[3]) ? node10401 : node10398;
													assign node10398 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node10401 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node10404 = (inp[4]) ? node10408 : node10405;
													assign node10405 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node10408 = (inp[11]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node10411 = (inp[3]) ? node10427 : node10412;
											assign node10412 = (inp[14]) ? node10420 : node10413;
												assign node10413 = (inp[4]) ? node10417 : node10414;
													assign node10414 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node10417 = (inp[7]) ? 15'b000000000011111 : 15'b000000001111111;
												assign node10420 = (inp[8]) ? node10424 : node10421;
													assign node10421 = (inp[7]) ? 15'b000000000111111 : 15'b000000000111111;
													assign node10424 = (inp[4]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node10427 = (inp[11]) ? node10435 : node10428;
												assign node10428 = (inp[7]) ? node10432 : node10429;
													assign node10429 = (inp[8]) ? 15'b000000000111111 : 15'b000000000111111;
													assign node10432 = (inp[8]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node10435 = (inp[14]) ? 15'b000000000001111 : node10436;
													assign node10436 = (inp[4]) ? 15'b000000000011111 : 15'b000000000011111;
							assign node10440 = (inp[4]) ? node10554 : node10441;
								assign node10441 = (inp[8]) ? node10501 : node10442;
									assign node10442 = (inp[14]) ? node10474 : node10443;
										assign node10443 = (inp[11]) ? node10459 : node10444;
											assign node10444 = (inp[2]) ? node10452 : node10445;
												assign node10445 = (inp[9]) ? node10449 : node10446;
													assign node10446 = (inp[7]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node10449 = (inp[7]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node10452 = (inp[3]) ? node10456 : node10453;
													assign node10453 = (inp[7]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node10456 = (inp[9]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node10459 = (inp[5]) ? node10467 : node10460;
												assign node10460 = (inp[2]) ? node10464 : node10461;
													assign node10461 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node10464 = (inp[3]) ? 15'b000000001111111 : 15'b000000001111111;
												assign node10467 = (inp[9]) ? node10471 : node10468;
													assign node10468 = (inp[2]) ? 15'b000000001111111 : 15'b000000001111111;
													assign node10471 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node10474 = (inp[9]) ? node10486 : node10475;
											assign node10475 = (inp[5]) ? node10479 : node10476;
												assign node10476 = (inp[2]) ? 15'b000000111111111 : 15'b000000011111111;
												assign node10479 = (inp[11]) ? node10483 : node10480;
													assign node10480 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node10483 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node10486 = (inp[3]) ? node10494 : node10487;
												assign node10487 = (inp[7]) ? node10491 : node10488;
													assign node10488 = (inp[11]) ? 15'b000000001111111 : 15'b000000001111111;
													assign node10491 = (inp[5]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node10494 = (inp[2]) ? node10498 : node10495;
													assign node10495 = (inp[7]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node10498 = (inp[7]) ? 15'b000000000001111 : 15'b000000000111111;
									assign node10501 = (inp[5]) ? node10525 : node10502;
										assign node10502 = (inp[3]) ? node10514 : node10503;
											assign node10503 = (inp[14]) ? node10509 : node10504;
												assign node10504 = (inp[9]) ? node10506 : 15'b000000111111111;
													assign node10506 = (inp[7]) ? 15'b000000011111111 : 15'b000000011111111;
												assign node10509 = (inp[11]) ? 15'b000000001111111 : node10510;
													assign node10510 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node10514 = (inp[11]) ? node10520 : node10515;
												assign node10515 = (inp[7]) ? node10517 : 15'b000000011111111;
													assign node10517 = (inp[14]) ? 15'b000000000011111 : 15'b000000001111111;
												assign node10520 = (inp[14]) ? node10522 : 15'b000000000111111;
													assign node10522 = (inp[2]) ? 15'b000000000111111 : 15'b000000000111111;
										assign node10525 = (inp[3]) ? node10539 : node10526;
											assign node10526 = (inp[14]) ? node10532 : node10527;
												assign node10527 = (inp[2]) ? 15'b000000001111111 : node10528;
													assign node10528 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node10532 = (inp[9]) ? node10536 : node10533;
													assign node10533 = (inp[7]) ? 15'b000000000011111 : 15'b000000001111111;
													assign node10536 = (inp[2]) ? 15'b000000000011111 : 15'b000000000011111;
											assign node10539 = (inp[11]) ? node10547 : node10540;
												assign node10540 = (inp[2]) ? node10544 : node10541;
													assign node10541 = (inp[7]) ? 15'b000000000111111 : 15'b000000000111111;
													assign node10544 = (inp[9]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node10547 = (inp[9]) ? node10551 : node10548;
													assign node10548 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node10551 = (inp[14]) ? 15'b000000000001111 : 15'b000000000011111;
								assign node10554 = (inp[5]) ? node10616 : node10555;
									assign node10555 = (inp[14]) ? node10585 : node10556;
										assign node10556 = (inp[9]) ? node10570 : node10557;
											assign node10557 = (inp[8]) ? node10563 : node10558;
												assign node10558 = (inp[3]) ? node10560 : 15'b000000011111111;
													assign node10560 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node10563 = (inp[7]) ? node10567 : node10564;
													assign node10564 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node10567 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node10570 = (inp[7]) ? node10578 : node10571;
												assign node10571 = (inp[8]) ? node10575 : node10572;
													assign node10572 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node10575 = (inp[2]) ? 15'b000000000111111 : 15'b000000000111111;
												assign node10578 = (inp[11]) ? node10582 : node10579;
													assign node10579 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node10582 = (inp[8]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node10585 = (inp[11]) ? node10601 : node10586;
											assign node10586 = (inp[3]) ? node10594 : node10587;
												assign node10587 = (inp[7]) ? node10591 : node10588;
													assign node10588 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node10591 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node10594 = (inp[9]) ? node10598 : node10595;
													assign node10595 = (inp[2]) ? 15'b000000000111111 : 15'b000000000111111;
													assign node10598 = (inp[7]) ? 15'b000000000001111 : 15'b000000000111111;
											assign node10601 = (inp[8]) ? node10609 : node10602;
												assign node10602 = (inp[3]) ? node10606 : node10603;
													assign node10603 = (inp[9]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node10606 = (inp[2]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node10609 = (inp[2]) ? node10613 : node10610;
													assign node10610 = (inp[7]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node10613 = (inp[9]) ? 15'b000000000001111 : 15'b000000000011111;
									assign node10616 = (inp[14]) ? node10648 : node10617;
										assign node10617 = (inp[9]) ? node10633 : node10618;
											assign node10618 = (inp[11]) ? node10626 : node10619;
												assign node10619 = (inp[7]) ? node10623 : node10620;
													assign node10620 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node10623 = (inp[8]) ? 15'b000000000111111 : 15'b000000000111111;
												assign node10626 = (inp[8]) ? node10630 : node10627;
													assign node10627 = (inp[7]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node10630 = (inp[3]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node10633 = (inp[2]) ? node10641 : node10634;
												assign node10634 = (inp[7]) ? node10638 : node10635;
													assign node10635 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node10638 = (inp[8]) ? 15'b000000000001111 : 15'b000000000111111;
												assign node10641 = (inp[11]) ? node10645 : node10642;
													assign node10642 = (inp[8]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node10645 = (inp[7]) ? 15'b000000000000111 : 15'b000000000001111;
										assign node10648 = (inp[2]) ? node10664 : node10649;
											assign node10649 = (inp[9]) ? node10657 : node10650;
												assign node10650 = (inp[8]) ? node10654 : node10651;
													assign node10651 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node10654 = (inp[7]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node10657 = (inp[11]) ? node10661 : node10658;
													assign node10658 = (inp[7]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node10661 = (inp[3]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node10664 = (inp[8]) ? node10672 : node10665;
												assign node10665 = (inp[7]) ? node10669 : node10666;
													assign node10666 = (inp[11]) ? 15'b000000000011111 : 15'b000000000011111;
													assign node10669 = (inp[9]) ? 15'b000000000000111 : 15'b000000000011111;
												assign node10672 = (inp[9]) ? node10676 : node10673;
													assign node10673 = (inp[11]) ? 15'b000000000001111 : 15'b000000000011111;
													assign node10676 = (inp[11]) ? 15'b000000000000111 : 15'b000000000000111;
					assign node10679 = (inp[7]) ? node11155 : node10680;
						assign node10680 = (inp[12]) ? node10920 : node10681;
							assign node10681 = (inp[11]) ? node10805 : node10682;
								assign node10682 = (inp[9]) ? node10744 : node10683;
									assign node10683 = (inp[5]) ? node10713 : node10684;
										assign node10684 = (inp[14]) ? node10698 : node10685;
											assign node10685 = (inp[4]) ? node10693 : node10686;
												assign node10686 = (inp[8]) ? node10690 : node10687;
													assign node10687 = (inp[2]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node10690 = (inp[1]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node10693 = (inp[8]) ? node10695 : 15'b000001111111111;
													assign node10695 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node10698 = (inp[8]) ? node10706 : node10699;
												assign node10699 = (inp[4]) ? node10703 : node10700;
													assign node10700 = (inp[1]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node10703 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node10706 = (inp[1]) ? node10710 : node10707;
													assign node10707 = (inp[4]) ? 15'b000000011111111 : 15'b000000011111111;
													assign node10710 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node10713 = (inp[4]) ? node10729 : node10714;
											assign node10714 = (inp[3]) ? node10722 : node10715;
												assign node10715 = (inp[8]) ? node10719 : node10716;
													assign node10716 = (inp[2]) ? 15'b000000111111111 : 15'b000011111111111;
													assign node10719 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node10722 = (inp[8]) ? node10726 : node10723;
													assign node10723 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node10726 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node10729 = (inp[14]) ? node10737 : node10730;
												assign node10730 = (inp[8]) ? node10734 : node10731;
													assign node10731 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node10734 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node10737 = (inp[2]) ? node10741 : node10738;
													assign node10738 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node10741 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node10744 = (inp[8]) ? node10776 : node10745;
										assign node10745 = (inp[1]) ? node10761 : node10746;
											assign node10746 = (inp[14]) ? node10754 : node10747;
												assign node10747 = (inp[3]) ? node10751 : node10748;
													assign node10748 = (inp[5]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node10751 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node10754 = (inp[2]) ? node10758 : node10755;
													assign node10755 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node10758 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node10761 = (inp[3]) ? node10769 : node10762;
												assign node10762 = (inp[2]) ? node10766 : node10763;
													assign node10763 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node10766 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node10769 = (inp[5]) ? node10773 : node10770;
													assign node10770 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node10773 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node10776 = (inp[3]) ? node10790 : node10777;
											assign node10777 = (inp[2]) ? node10785 : node10778;
												assign node10778 = (inp[1]) ? node10782 : node10779;
													assign node10779 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node10782 = (inp[14]) ? 15'b000000000111111 : 15'b000000011111111;
												assign node10785 = (inp[4]) ? 15'b000000000111111 : node10786;
													assign node10786 = (inp[5]) ? 15'b000000001111111 : 15'b000000001111111;
											assign node10790 = (inp[5]) ? node10798 : node10791;
												assign node10791 = (inp[2]) ? node10795 : node10792;
													assign node10792 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node10795 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node10798 = (inp[1]) ? node10802 : node10799;
													assign node10799 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node10802 = (inp[2]) ? 15'b000000000011111 : 15'b000000000111111;
								assign node10805 = (inp[8]) ? node10863 : node10806;
									assign node10806 = (inp[9]) ? node10832 : node10807;
										assign node10807 = (inp[4]) ? node10819 : node10808;
											assign node10808 = (inp[14]) ? node10814 : node10809;
												assign node10809 = (inp[1]) ? 15'b000000111111111 : node10810;
													assign node10810 = (inp[5]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node10814 = (inp[3]) ? node10816 : 15'b000000111111111;
													assign node10816 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node10819 = (inp[2]) ? node10825 : node10820;
												assign node10820 = (inp[1]) ? 15'b000000011111111 : node10821;
													assign node10821 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node10825 = (inp[14]) ? node10829 : node10826;
													assign node10826 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node10829 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node10832 = (inp[3]) ? node10848 : node10833;
											assign node10833 = (inp[14]) ? node10841 : node10834;
												assign node10834 = (inp[1]) ? node10838 : node10835;
													assign node10835 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node10838 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node10841 = (inp[4]) ? node10845 : node10842;
													assign node10842 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node10845 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node10848 = (inp[14]) ? node10856 : node10849;
												assign node10849 = (inp[5]) ? node10853 : node10850;
													assign node10850 = (inp[1]) ? 15'b000000001111111 : 15'b000000001111111;
													assign node10853 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node10856 = (inp[1]) ? node10860 : node10857;
													assign node10857 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node10860 = (inp[4]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node10863 = (inp[9]) ? node10891 : node10864;
										assign node10864 = (inp[1]) ? node10878 : node10865;
											assign node10865 = (inp[3]) ? node10871 : node10866;
												assign node10866 = (inp[14]) ? node10868 : 15'b000000011111111;
													assign node10868 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node10871 = (inp[2]) ? node10875 : node10872;
													assign node10872 = (inp[14]) ? 15'b000000001111111 : 15'b000000001111111;
													assign node10875 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node10878 = (inp[14]) ? node10886 : node10879;
												assign node10879 = (inp[5]) ? node10883 : node10880;
													assign node10880 = (inp[4]) ? 15'b000000001111111 : 15'b000000001111111;
													assign node10883 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node10886 = (inp[3]) ? node10888 : 15'b000000000111111;
													assign node10888 = (inp[5]) ? 15'b000000000011111 : 15'b000000000011111;
										assign node10891 = (inp[4]) ? node10907 : node10892;
											assign node10892 = (inp[14]) ? node10900 : node10893;
												assign node10893 = (inp[5]) ? node10897 : node10894;
													assign node10894 = (inp[2]) ? 15'b000000001111111 : 15'b000000111111111;
													assign node10897 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node10900 = (inp[3]) ? node10904 : node10901;
													assign node10901 = (inp[5]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node10904 = (inp[2]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node10907 = (inp[2]) ? node10915 : node10908;
												assign node10908 = (inp[5]) ? node10912 : node10909;
													assign node10909 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node10912 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node10915 = (inp[5]) ? 15'b000000000011111 : node10916;
													assign node10916 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
							assign node10920 = (inp[8]) ? node11034 : node10921;
								assign node10921 = (inp[11]) ? node10977 : node10922;
									assign node10922 = (inp[5]) ? node10948 : node10923;
										assign node10923 = (inp[1]) ? node10933 : node10924;
											assign node10924 = (inp[2]) ? 15'b000000111111111 : node10925;
												assign node10925 = (inp[4]) ? node10929 : node10926;
													assign node10926 = (inp[3]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node10929 = (inp[9]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node10933 = (inp[4]) ? node10941 : node10934;
												assign node10934 = (inp[3]) ? node10938 : node10935;
													assign node10935 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node10938 = (inp[9]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node10941 = (inp[2]) ? node10945 : node10942;
													assign node10942 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node10945 = (inp[3]) ? 15'b000000000111111 : 15'b000000000111111;
										assign node10948 = (inp[9]) ? node10964 : node10949;
											assign node10949 = (inp[2]) ? node10957 : node10950;
												assign node10950 = (inp[14]) ? node10954 : node10951;
													assign node10951 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node10954 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node10957 = (inp[3]) ? node10961 : node10958;
													assign node10958 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node10961 = (inp[14]) ? 15'b000000000111111 : 15'b000000000111111;
											assign node10964 = (inp[3]) ? node10972 : node10965;
												assign node10965 = (inp[1]) ? node10969 : node10966;
													assign node10966 = (inp[2]) ? 15'b000000000111111 : 15'b000000011111111;
													assign node10969 = (inp[14]) ? 15'b000000000011111 : 15'b000000001111111;
												assign node10972 = (inp[1]) ? node10974 : 15'b000000000111111;
													assign node10974 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node10977 = (inp[1]) ? node11005 : node10978;
										assign node10978 = (inp[2]) ? node10990 : node10979;
											assign node10979 = (inp[9]) ? node10985 : node10980;
												assign node10980 = (inp[3]) ? 15'b000000011111111 : node10981;
													assign node10981 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node10985 = (inp[3]) ? 15'b000000000111111 : node10986;
													assign node10986 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node10990 = (inp[14]) ? node10998 : node10991;
												assign node10991 = (inp[5]) ? node10995 : node10992;
													assign node10992 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node10995 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node10998 = (inp[3]) ? node11002 : node10999;
													assign node10999 = (inp[5]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node11002 = (inp[4]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node11005 = (inp[3]) ? node11021 : node11006;
											assign node11006 = (inp[2]) ? node11014 : node11007;
												assign node11007 = (inp[5]) ? node11011 : node11008;
													assign node11008 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node11011 = (inp[9]) ? 15'b000000000011111 : 15'b000000001111111;
												assign node11014 = (inp[4]) ? node11018 : node11015;
													assign node11015 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node11018 = (inp[9]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node11021 = (inp[4]) ? node11027 : node11022;
												assign node11022 = (inp[9]) ? node11024 : 15'b000000000111111;
													assign node11024 = (inp[5]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node11027 = (inp[2]) ? node11031 : node11028;
													assign node11028 = (inp[5]) ? 15'b000000000011111 : 15'b000000000011111;
													assign node11031 = (inp[5]) ? 15'b000000000000111 : 15'b000000000001111;
								assign node11034 = (inp[1]) ? node11092 : node11035;
									assign node11035 = (inp[11]) ? node11067 : node11036;
										assign node11036 = (inp[4]) ? node11052 : node11037;
											assign node11037 = (inp[9]) ? node11045 : node11038;
												assign node11038 = (inp[3]) ? node11042 : node11039;
													assign node11039 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node11042 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node11045 = (inp[2]) ? node11049 : node11046;
													assign node11046 = (inp[14]) ? 15'b000000000111111 : 15'b000000011111111;
													assign node11049 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node11052 = (inp[2]) ? node11060 : node11053;
												assign node11053 = (inp[3]) ? node11057 : node11054;
													assign node11054 = (inp[5]) ? 15'b000000001111111 : 15'b000000111111111;
													assign node11057 = (inp[9]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node11060 = (inp[9]) ? node11064 : node11061;
													assign node11061 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node11064 = (inp[5]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node11067 = (inp[5]) ? node11077 : node11068;
											assign node11068 = (inp[3]) ? 15'b000000000111111 : node11069;
												assign node11069 = (inp[4]) ? node11073 : node11070;
													assign node11070 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node11073 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node11077 = (inp[14]) ? node11085 : node11078;
												assign node11078 = (inp[9]) ? node11082 : node11079;
													assign node11079 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node11082 = (inp[4]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node11085 = (inp[2]) ? node11089 : node11086;
													assign node11086 = (inp[4]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node11089 = (inp[9]) ? 15'b000000000001111 : 15'b000000000011111;
									assign node11092 = (inp[2]) ? node11124 : node11093;
										assign node11093 = (inp[3]) ? node11109 : node11094;
											assign node11094 = (inp[14]) ? node11102 : node11095;
												assign node11095 = (inp[5]) ? node11099 : node11096;
													assign node11096 = (inp[9]) ? 15'b000000001111111 : 15'b000000111111111;
													assign node11099 = (inp[9]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node11102 = (inp[9]) ? node11106 : node11103;
													assign node11103 = (inp[11]) ? 15'b000000000111111 : 15'b000000011111111;
													assign node11106 = (inp[11]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node11109 = (inp[14]) ? node11117 : node11110;
												assign node11110 = (inp[4]) ? node11114 : node11111;
													assign node11111 = (inp[9]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node11114 = (inp[11]) ? 15'b000000000001111 : 15'b000000000111111;
												assign node11117 = (inp[9]) ? node11121 : node11118;
													assign node11118 = (inp[11]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node11121 = (inp[5]) ? 15'b000000000001111 : 15'b000000000011111;
										assign node11124 = (inp[11]) ? node11140 : node11125;
											assign node11125 = (inp[9]) ? node11133 : node11126;
												assign node11126 = (inp[5]) ? node11130 : node11127;
													assign node11127 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node11130 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node11133 = (inp[4]) ? node11137 : node11134;
													assign node11134 = (inp[14]) ? 15'b000000000001111 : 15'b000000000111111;
													assign node11137 = (inp[14]) ? 15'b000000000001111 : 15'b000000000001111;
											assign node11140 = (inp[14]) ? node11148 : node11141;
												assign node11141 = (inp[3]) ? node11145 : node11142;
													assign node11142 = (inp[9]) ? 15'b000000000111111 : 15'b000000000011111;
													assign node11145 = (inp[4]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node11148 = (inp[5]) ? node11152 : node11149;
													assign node11149 = (inp[9]) ? 15'b000000000001111 : 15'b000000000011111;
													assign node11152 = (inp[9]) ? 15'b000000000000111 : 15'b000000000001111;
						assign node11155 = (inp[9]) ? node11387 : node11156;
							assign node11156 = (inp[14]) ? node11268 : node11157;
								assign node11157 = (inp[12]) ? node11215 : node11158;
									assign node11158 = (inp[8]) ? node11184 : node11159;
										assign node11159 = (inp[1]) ? node11171 : node11160;
											assign node11160 = (inp[3]) ? node11166 : node11161;
												assign node11161 = (inp[2]) ? 15'b000000011111111 : node11162;
													assign node11162 = (inp[11]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node11166 = (inp[5]) ? 15'b000000011111111 : node11167;
													assign node11167 = (inp[11]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node11171 = (inp[2]) ? node11177 : node11172;
												assign node11172 = (inp[3]) ? node11174 : 15'b000000111111111;
													assign node11174 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node11177 = (inp[5]) ? node11181 : node11178;
													assign node11178 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node11181 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node11184 = (inp[5]) ? node11200 : node11185;
											assign node11185 = (inp[4]) ? node11193 : node11186;
												assign node11186 = (inp[3]) ? node11190 : node11187;
													assign node11187 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node11190 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node11193 = (inp[1]) ? node11197 : node11194;
													assign node11194 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node11197 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node11200 = (inp[4]) ? node11208 : node11201;
												assign node11201 = (inp[11]) ? node11205 : node11202;
													assign node11202 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node11205 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node11208 = (inp[11]) ? node11212 : node11209;
													assign node11209 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node11212 = (inp[3]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node11215 = (inp[8]) ? node11245 : node11216;
										assign node11216 = (inp[1]) ? node11230 : node11217;
											assign node11217 = (inp[4]) ? node11223 : node11218;
												assign node11218 = (inp[5]) ? 15'b000000011111111 : node11219;
													assign node11219 = (inp[11]) ? 15'b000000011111111 : 15'b000001111111111;
												assign node11223 = (inp[5]) ? node11227 : node11224;
													assign node11224 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node11227 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node11230 = (inp[3]) ? node11238 : node11231;
												assign node11231 = (inp[4]) ? node11235 : node11232;
													assign node11232 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node11235 = (inp[5]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node11238 = (inp[5]) ? node11242 : node11239;
													assign node11239 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node11242 = (inp[2]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node11245 = (inp[2]) ? node11253 : node11246;
											assign node11246 = (inp[4]) ? 15'b000000000111111 : node11247;
												assign node11247 = (inp[3]) ? node11249 : 15'b000000001111111;
													assign node11249 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node11253 = (inp[3]) ? node11261 : node11254;
												assign node11254 = (inp[1]) ? node11258 : node11255;
													assign node11255 = (inp[5]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node11258 = (inp[4]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node11261 = (inp[11]) ? node11265 : node11262;
													assign node11262 = (inp[4]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node11265 = (inp[5]) ? 15'b000000000001111 : 15'b000000000011111;
								assign node11268 = (inp[5]) ? node11330 : node11269;
									assign node11269 = (inp[8]) ? node11301 : node11270;
										assign node11270 = (inp[4]) ? node11286 : node11271;
											assign node11271 = (inp[1]) ? node11279 : node11272;
												assign node11272 = (inp[3]) ? node11276 : node11273;
													assign node11273 = (inp[12]) ? 15'b000000011111111 : 15'b000000011111111;
													assign node11276 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node11279 = (inp[2]) ? node11283 : node11280;
													assign node11280 = (inp[11]) ? 15'b000000001111111 : 15'b000000001111111;
													assign node11283 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node11286 = (inp[12]) ? node11294 : node11287;
												assign node11287 = (inp[11]) ? node11291 : node11288;
													assign node11288 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node11291 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node11294 = (inp[1]) ? node11298 : node11295;
													assign node11295 = (inp[3]) ? 15'b000000000111111 : 15'b000000000111111;
													assign node11298 = (inp[11]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node11301 = (inp[1]) ? node11317 : node11302;
											assign node11302 = (inp[2]) ? node11310 : node11303;
												assign node11303 = (inp[11]) ? node11307 : node11304;
													assign node11304 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node11307 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node11310 = (inp[11]) ? node11314 : node11311;
													assign node11311 = (inp[12]) ? 15'b000000000111111 : 15'b000000000111111;
													assign node11314 = (inp[3]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node11317 = (inp[3]) ? node11325 : node11318;
												assign node11318 = (inp[12]) ? node11322 : node11319;
													assign node11319 = (inp[2]) ? 15'b000000000111111 : 15'b000000000111111;
													assign node11322 = (inp[2]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node11325 = (inp[2]) ? 15'b000000000001111 : node11326;
													assign node11326 = (inp[12]) ? 15'b000000000011111 : 15'b000000000011111;
									assign node11330 = (inp[11]) ? node11358 : node11331;
										assign node11331 = (inp[2]) ? node11345 : node11332;
											assign node11332 = (inp[1]) ? node11340 : node11333;
												assign node11333 = (inp[8]) ? node11337 : node11334;
													assign node11334 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node11337 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node11340 = (inp[3]) ? node11342 : 15'b000000000111111;
													assign node11342 = (inp[12]) ? 15'b000000000111111 : 15'b000000000011111;
											assign node11345 = (inp[4]) ? node11353 : node11346;
												assign node11346 = (inp[8]) ? node11350 : node11347;
													assign node11347 = (inp[3]) ? 15'b000000000111111 : 15'b000000000111111;
													assign node11350 = (inp[12]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node11353 = (inp[3]) ? node11355 : 15'b000000001111111;
													assign node11355 = (inp[8]) ? 15'b000000000000111 : 15'b000000000001111;
										assign node11358 = (inp[4]) ? node11372 : node11359;
											assign node11359 = (inp[12]) ? node11365 : node11360;
												assign node11360 = (inp[2]) ? 15'b000000001111111 : node11361;
													assign node11361 = (inp[8]) ? 15'b000000000111111 : 15'b000000000111111;
												assign node11365 = (inp[1]) ? node11369 : node11366;
													assign node11366 = (inp[3]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node11369 = (inp[8]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node11372 = (inp[2]) ? node11380 : node11373;
												assign node11373 = (inp[12]) ? node11377 : node11374;
													assign node11374 = (inp[8]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node11377 = (inp[3]) ? 15'b000000000000111 : 15'b000000000011111;
												assign node11380 = (inp[8]) ? node11384 : node11381;
													assign node11381 = (inp[1]) ? 15'b000000000001111 : 15'b000000000001111;
													assign node11384 = (inp[3]) ? 15'b000000000000111 : 15'b000000000001111;
							assign node11387 = (inp[8]) ? node11513 : node11388;
								assign node11388 = (inp[3]) ? node11450 : node11389;
									assign node11389 = (inp[12]) ? node11419 : node11390;
										assign node11390 = (inp[5]) ? node11404 : node11391;
											assign node11391 = (inp[11]) ? node11399 : node11392;
												assign node11392 = (inp[2]) ? node11396 : node11393;
													assign node11393 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node11396 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node11399 = (inp[4]) ? node11401 : 15'b000000011111111;
													assign node11401 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node11404 = (inp[4]) ? node11412 : node11405;
												assign node11405 = (inp[14]) ? node11409 : node11406;
													assign node11406 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node11409 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node11412 = (inp[2]) ? node11416 : node11413;
													assign node11413 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node11416 = (inp[11]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node11419 = (inp[11]) ? node11435 : node11420;
											assign node11420 = (inp[5]) ? node11428 : node11421;
												assign node11421 = (inp[1]) ? node11425 : node11422;
													assign node11422 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node11425 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node11428 = (inp[4]) ? node11432 : node11429;
													assign node11429 = (inp[14]) ? 15'b000000000111111 : 15'b000000000111111;
													assign node11432 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node11435 = (inp[4]) ? node11443 : node11436;
												assign node11436 = (inp[2]) ? node11440 : node11437;
													assign node11437 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node11440 = (inp[1]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node11443 = (inp[5]) ? node11447 : node11444;
													assign node11444 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node11447 = (inp[14]) ? 15'b000000000001111 : 15'b000000000011111;
									assign node11450 = (inp[4]) ? node11482 : node11451;
										assign node11451 = (inp[14]) ? node11467 : node11452;
											assign node11452 = (inp[11]) ? node11460 : node11453;
												assign node11453 = (inp[12]) ? node11457 : node11454;
													assign node11454 = (inp[5]) ? 15'b000000001111111 : 15'b000000111111111;
													assign node11457 = (inp[5]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node11460 = (inp[12]) ? node11464 : node11461;
													assign node11461 = (inp[5]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node11464 = (inp[2]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node11467 = (inp[12]) ? node11475 : node11468;
												assign node11468 = (inp[2]) ? node11472 : node11469;
													assign node11469 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node11472 = (inp[1]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node11475 = (inp[2]) ? node11479 : node11476;
													assign node11476 = (inp[11]) ? 15'b000000000001111 : 15'b000000000111111;
													assign node11479 = (inp[5]) ? 15'b000000000001111 : 15'b000000000011111;
										assign node11482 = (inp[5]) ? node11498 : node11483;
											assign node11483 = (inp[2]) ? node11491 : node11484;
												assign node11484 = (inp[11]) ? node11488 : node11485;
													assign node11485 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node11488 = (inp[1]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node11491 = (inp[14]) ? node11495 : node11492;
													assign node11492 = (inp[12]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node11495 = (inp[11]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node11498 = (inp[12]) ? node11506 : node11499;
												assign node11499 = (inp[11]) ? node11503 : node11500;
													assign node11500 = (inp[2]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node11503 = (inp[2]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node11506 = (inp[1]) ? node11510 : node11507;
													assign node11507 = (inp[11]) ? 15'b000000000001111 : 15'b000000000011111;
													assign node11510 = (inp[11]) ? 15'b000000000000111 : 15'b000000000001111;
								assign node11513 = (inp[2]) ? node11577 : node11514;
									assign node11514 = (inp[3]) ? node11546 : node11515;
										assign node11515 = (inp[11]) ? node11531 : node11516;
											assign node11516 = (inp[5]) ? node11524 : node11517;
												assign node11517 = (inp[4]) ? node11521 : node11518;
													assign node11518 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node11521 = (inp[12]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node11524 = (inp[14]) ? node11528 : node11525;
													assign node11525 = (inp[12]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node11528 = (inp[4]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node11531 = (inp[5]) ? node11539 : node11532;
												assign node11532 = (inp[1]) ? node11536 : node11533;
													assign node11533 = (inp[12]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node11536 = (inp[4]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node11539 = (inp[1]) ? node11543 : node11540;
													assign node11540 = (inp[4]) ? 15'b000000000011111 : 15'b000000000011111;
													assign node11543 = (inp[4]) ? 15'b000000000000111 : 15'b000000000011111;
										assign node11546 = (inp[12]) ? node11562 : node11547;
											assign node11547 = (inp[1]) ? node11555 : node11548;
												assign node11548 = (inp[14]) ? node11552 : node11549;
													assign node11549 = (inp[5]) ? 15'b000000000111111 : 15'b000000000111111;
													assign node11552 = (inp[5]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node11555 = (inp[14]) ? node11559 : node11556;
													assign node11556 = (inp[4]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node11559 = (inp[5]) ? 15'b000000000001111 : 15'b000000000001111;
											assign node11562 = (inp[14]) ? node11570 : node11563;
												assign node11563 = (inp[4]) ? node11567 : node11564;
													assign node11564 = (inp[1]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node11567 = (inp[11]) ? 15'b000000000000111 : 15'b000000000011111;
												assign node11570 = (inp[11]) ? node11574 : node11571;
													assign node11571 = (inp[4]) ? 15'b000000000001111 : 15'b000000000001111;
													assign node11574 = (inp[5]) ? 15'b000000000000111 : 15'b000000000001111;
									assign node11577 = (inp[4]) ? node11605 : node11578;
										assign node11578 = (inp[3]) ? node11592 : node11579;
											assign node11579 = (inp[1]) ? node11585 : node11580;
												assign node11580 = (inp[5]) ? 15'b000000000111111 : node11581;
													assign node11581 = (inp[12]) ? 15'b000000001111111 : 15'b000000001111111;
												assign node11585 = (inp[11]) ? node11589 : node11586;
													assign node11586 = (inp[5]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node11589 = (inp[12]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node11592 = (inp[12]) ? node11600 : node11593;
												assign node11593 = (inp[14]) ? node11597 : node11594;
													assign node11594 = (inp[5]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node11597 = (inp[11]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node11600 = (inp[11]) ? node11602 : 15'b000000000001111;
													assign node11602 = (inp[1]) ? 15'b000000000000111 : 15'b000000000001111;
										assign node11605 = (inp[12]) ? node11619 : node11606;
											assign node11606 = (inp[11]) ? node11612 : node11607;
												assign node11607 = (inp[14]) ? node11609 : 15'b000000000011111;
													assign node11609 = (inp[3]) ? 15'b000000000000111 : 15'b000000000011111;
												assign node11612 = (inp[3]) ? node11616 : node11613;
													assign node11613 = (inp[5]) ? 15'b000000000001111 : 15'b000000000011111;
													assign node11616 = (inp[1]) ? 15'b000000000000111 : 15'b000000000001111;
											assign node11619 = (inp[5]) ? node11627 : node11620;
												assign node11620 = (inp[11]) ? node11624 : node11621;
													assign node11621 = (inp[1]) ? 15'b000000000000111 : 15'b000000000011111;
													assign node11624 = (inp[14]) ? 15'b000000000000111 : 15'b000000000001111;
												assign node11627 = (inp[14]) ? node11631 : node11628;
													assign node11628 = (inp[1]) ? 15'b000000000000111 : 15'b000000000001111;
													assign node11631 = (inp[3]) ? 15'b000000000000011 : 15'b000000000000111;
			assign node11634 = (inp[3]) ? node13596 : node11635;
				assign node11635 = (inp[12]) ? node12619 : node11636;
					assign node11636 = (inp[9]) ? node12128 : node11637;
						assign node11637 = (inp[14]) ? node11885 : node11638;
							assign node11638 = (inp[4]) ? node11764 : node11639;
								assign node11639 = (inp[7]) ? node11701 : node11640;
									assign node11640 = (inp[10]) ? node11672 : node11641;
										assign node11641 = (inp[5]) ? node11657 : node11642;
											assign node11642 = (inp[2]) ? node11650 : node11643;
												assign node11643 = (inp[13]) ? node11647 : node11644;
													assign node11644 = (inp[11]) ? 15'b000011111111111 : 15'b000111111111111;
													assign node11647 = (inp[8]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node11650 = (inp[1]) ? node11654 : node11651;
													assign node11651 = (inp[8]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node11654 = (inp[8]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node11657 = (inp[1]) ? node11665 : node11658;
												assign node11658 = (inp[11]) ? node11662 : node11659;
													assign node11659 = (inp[8]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node11662 = (inp[8]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node11665 = (inp[13]) ? node11669 : node11666;
													assign node11666 = (inp[2]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node11669 = (inp[11]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node11672 = (inp[8]) ? node11686 : node11673;
											assign node11673 = (inp[2]) ? node11679 : node11674;
												assign node11674 = (inp[1]) ? node11676 : 15'b000011111111111;
													assign node11676 = (inp[5]) ? 15'b000000011111111 : 15'b000001111111111;
												assign node11679 = (inp[13]) ? node11683 : node11680;
													assign node11680 = (inp[5]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node11683 = (inp[11]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node11686 = (inp[1]) ? node11694 : node11687;
												assign node11687 = (inp[13]) ? node11691 : node11688;
													assign node11688 = (inp[11]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node11691 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node11694 = (inp[5]) ? node11698 : node11695;
													assign node11695 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node11698 = (inp[2]) ? 15'b000000000111111 : 15'b000000011111111;
									assign node11701 = (inp[5]) ? node11733 : node11702;
										assign node11702 = (inp[8]) ? node11718 : node11703;
											assign node11703 = (inp[11]) ? node11711 : node11704;
												assign node11704 = (inp[10]) ? node11708 : node11705;
													assign node11705 = (inp[13]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node11708 = (inp[1]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node11711 = (inp[1]) ? node11715 : node11712;
													assign node11712 = (inp[10]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node11715 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node11718 = (inp[2]) ? node11726 : node11719;
												assign node11719 = (inp[10]) ? node11723 : node11720;
													assign node11720 = (inp[11]) ? 15'b000000111111111 : 15'b000000111111111;
													assign node11723 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node11726 = (inp[10]) ? node11730 : node11727;
													assign node11727 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node11730 = (inp[1]) ? 15'b000000000111111 : 15'b000000011111111;
										assign node11733 = (inp[8]) ? node11749 : node11734;
											assign node11734 = (inp[11]) ? node11742 : node11735;
												assign node11735 = (inp[2]) ? node11739 : node11736;
													assign node11736 = (inp[13]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node11739 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node11742 = (inp[1]) ? node11746 : node11743;
													assign node11743 = (inp[2]) ? 15'b000000011111111 : 15'b000000011111111;
													assign node11746 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node11749 = (inp[10]) ? node11757 : node11750;
												assign node11750 = (inp[2]) ? node11754 : node11751;
													assign node11751 = (inp[11]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node11754 = (inp[13]) ? 15'b000000000111111 : 15'b000000011111111;
												assign node11757 = (inp[1]) ? node11761 : node11758;
													assign node11758 = (inp[2]) ? 15'b000000001111111 : 15'b000000001111111;
													assign node11761 = (inp[11]) ? 15'b000000000011111 : 15'b000000001111111;
								assign node11764 = (inp[1]) ? node11824 : node11765;
									assign node11765 = (inp[13]) ? node11797 : node11766;
										assign node11766 = (inp[10]) ? node11782 : node11767;
											assign node11767 = (inp[7]) ? node11775 : node11768;
												assign node11768 = (inp[5]) ? node11772 : node11769;
													assign node11769 = (inp[2]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node11772 = (inp[11]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node11775 = (inp[5]) ? node11779 : node11776;
													assign node11776 = (inp[2]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node11779 = (inp[8]) ? 15'b000000011111111 : 15'b000001111111111;
											assign node11782 = (inp[8]) ? node11790 : node11783;
												assign node11783 = (inp[5]) ? node11787 : node11784;
													assign node11784 = (inp[11]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node11787 = (inp[7]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node11790 = (inp[2]) ? node11794 : node11791;
													assign node11791 = (inp[11]) ? 15'b000000011111111 : 15'b000001111111111;
													assign node11794 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node11797 = (inp[2]) ? node11811 : node11798;
											assign node11798 = (inp[7]) ? node11806 : node11799;
												assign node11799 = (inp[11]) ? node11803 : node11800;
													assign node11800 = (inp[10]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node11803 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node11806 = (inp[10]) ? 15'b000000001111111 : node11807;
													assign node11807 = (inp[11]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node11811 = (inp[7]) ? node11819 : node11812;
												assign node11812 = (inp[10]) ? node11816 : node11813;
													assign node11813 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node11816 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node11819 = (inp[5]) ? node11821 : 15'b000000011111111;
													assign node11821 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node11824 = (inp[2]) ? node11856 : node11825;
										assign node11825 = (inp[11]) ? node11841 : node11826;
											assign node11826 = (inp[8]) ? node11834 : node11827;
												assign node11827 = (inp[7]) ? node11831 : node11828;
													assign node11828 = (inp[10]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node11831 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node11834 = (inp[13]) ? node11838 : node11835;
													assign node11835 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node11838 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node11841 = (inp[13]) ? node11849 : node11842;
												assign node11842 = (inp[5]) ? node11846 : node11843;
													assign node11843 = (inp[7]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node11846 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node11849 = (inp[10]) ? node11853 : node11850;
													assign node11850 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node11853 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node11856 = (inp[5]) ? node11872 : node11857;
											assign node11857 = (inp[13]) ? node11865 : node11858;
												assign node11858 = (inp[11]) ? node11862 : node11859;
													assign node11859 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node11862 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node11865 = (inp[11]) ? node11869 : node11866;
													assign node11866 = (inp[10]) ? 15'b000000001111111 : 15'b000000001111111;
													assign node11869 = (inp[7]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node11872 = (inp[10]) ? node11880 : node11873;
												assign node11873 = (inp[7]) ? node11877 : node11874;
													assign node11874 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node11877 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node11880 = (inp[8]) ? node11882 : 15'b000000000111111;
													assign node11882 = (inp[13]) ? 15'b000000000011111 : 15'b000000000111111;
							assign node11885 = (inp[8]) ? node12007 : node11886;
								assign node11886 = (inp[7]) ? node11948 : node11887;
									assign node11887 = (inp[1]) ? node11919 : node11888;
										assign node11888 = (inp[4]) ? node11904 : node11889;
											assign node11889 = (inp[13]) ? node11897 : node11890;
												assign node11890 = (inp[2]) ? node11894 : node11891;
													assign node11891 = (inp[5]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node11894 = (inp[5]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node11897 = (inp[5]) ? node11901 : node11898;
													assign node11898 = (inp[11]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node11901 = (inp[10]) ? 15'b000000011111111 : 15'b000000011111111;
											assign node11904 = (inp[11]) ? node11912 : node11905;
												assign node11905 = (inp[2]) ? node11909 : node11906;
													assign node11906 = (inp[10]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node11909 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node11912 = (inp[10]) ? node11916 : node11913;
													assign node11913 = (inp[13]) ? 15'b000000011111111 : 15'b000000011111111;
													assign node11916 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node11919 = (inp[11]) ? node11935 : node11920;
											assign node11920 = (inp[13]) ? node11928 : node11921;
												assign node11921 = (inp[10]) ? node11925 : node11922;
													assign node11922 = (inp[5]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node11925 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node11928 = (inp[2]) ? node11932 : node11929;
													assign node11929 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node11932 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node11935 = (inp[13]) ? node11943 : node11936;
												assign node11936 = (inp[4]) ? node11940 : node11937;
													assign node11937 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node11940 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node11943 = (inp[4]) ? 15'b000000000111111 : node11944;
													assign node11944 = (inp[5]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node11948 = (inp[13]) ? node11978 : node11949;
										assign node11949 = (inp[11]) ? node11965 : node11950;
											assign node11950 = (inp[1]) ? node11958 : node11951;
												assign node11951 = (inp[2]) ? node11955 : node11952;
													assign node11952 = (inp[4]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node11955 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node11958 = (inp[5]) ? node11962 : node11959;
													assign node11959 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node11962 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node11965 = (inp[2]) ? node11973 : node11966;
												assign node11966 = (inp[1]) ? node11970 : node11967;
													assign node11967 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node11970 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node11973 = (inp[1]) ? 15'b000000000111111 : node11974;
													assign node11974 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node11978 = (inp[10]) ? node11994 : node11979;
											assign node11979 = (inp[5]) ? node11987 : node11980;
												assign node11980 = (inp[4]) ? node11984 : node11981;
													assign node11981 = (inp[2]) ? 15'b000000011111111 : 15'b000000011111111;
													assign node11984 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node11987 = (inp[11]) ? node11991 : node11988;
													assign node11988 = (inp[4]) ? 15'b000000001111111 : 15'b000000111111111;
													assign node11991 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node11994 = (inp[2]) ? node12000 : node11995;
												assign node11995 = (inp[4]) ? node11997 : 15'b000000001111111;
													assign node11997 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node12000 = (inp[11]) ? node12004 : node12001;
													assign node12001 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node12004 = (inp[5]) ? 15'b000000000011111 : 15'b000000000011111;
								assign node12007 = (inp[10]) ? node12069 : node12008;
									assign node12008 = (inp[4]) ? node12040 : node12009;
										assign node12009 = (inp[1]) ? node12025 : node12010;
											assign node12010 = (inp[13]) ? node12018 : node12011;
												assign node12011 = (inp[5]) ? node12015 : node12012;
													assign node12012 = (inp[11]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node12015 = (inp[7]) ? 15'b000000111111111 : 15'b000000111111111;
												assign node12018 = (inp[5]) ? node12022 : node12019;
													assign node12019 = (inp[11]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node12022 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node12025 = (inp[13]) ? node12033 : node12026;
												assign node12026 = (inp[5]) ? node12030 : node12027;
													assign node12027 = (inp[7]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node12030 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node12033 = (inp[11]) ? node12037 : node12034;
													assign node12034 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node12037 = (inp[7]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node12040 = (inp[1]) ? node12056 : node12041;
											assign node12041 = (inp[13]) ? node12049 : node12042;
												assign node12042 = (inp[5]) ? node12046 : node12043;
													assign node12043 = (inp[11]) ? 15'b000000011111111 : 15'b000000011111111;
													assign node12046 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node12049 = (inp[7]) ? node12053 : node12050;
													assign node12050 = (inp[2]) ? 15'b000000000111111 : 15'b000000011111111;
													assign node12053 = (inp[2]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node12056 = (inp[11]) ? node12062 : node12057;
												assign node12057 = (inp[5]) ? 15'b000000000111111 : node12058;
													assign node12058 = (inp[13]) ? 15'b000000001111111 : 15'b000000001111111;
												assign node12062 = (inp[2]) ? node12066 : node12063;
													assign node12063 = (inp[13]) ? 15'b000000000111111 : 15'b000000000111111;
													assign node12066 = (inp[5]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node12069 = (inp[2]) ? node12099 : node12070;
										assign node12070 = (inp[11]) ? node12084 : node12071;
											assign node12071 = (inp[1]) ? node12077 : node12072;
												assign node12072 = (inp[7]) ? node12074 : 15'b000000011111111;
													assign node12074 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node12077 = (inp[4]) ? node12081 : node12078;
													assign node12078 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node12081 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node12084 = (inp[7]) ? node12092 : node12085;
												assign node12085 = (inp[13]) ? node12089 : node12086;
													assign node12086 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node12089 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node12092 = (inp[4]) ? node12096 : node12093;
													assign node12093 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node12096 = (inp[5]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node12099 = (inp[7]) ? node12115 : node12100;
											assign node12100 = (inp[11]) ? node12108 : node12101;
												assign node12101 = (inp[4]) ? node12105 : node12102;
													assign node12102 = (inp[13]) ? 15'b000000011111111 : 15'b000000001111111;
													assign node12105 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node12108 = (inp[1]) ? node12112 : node12109;
													assign node12109 = (inp[5]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node12112 = (inp[5]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node12115 = (inp[13]) ? node12123 : node12116;
												assign node12116 = (inp[4]) ? node12120 : node12117;
													assign node12117 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node12120 = (inp[11]) ? 15'b000000000011111 : 15'b000000000011111;
												assign node12123 = (inp[4]) ? node12125 : 15'b000000000011111;
													assign node12125 = (inp[5]) ? 15'b000000000001111 : 15'b000000000011111;
						assign node12128 = (inp[11]) ? node12374 : node12129;
							assign node12129 = (inp[13]) ? node12251 : node12130;
								assign node12130 = (inp[10]) ? node12190 : node12131;
									assign node12131 = (inp[7]) ? node12161 : node12132;
										assign node12132 = (inp[5]) ? node12146 : node12133;
											assign node12133 = (inp[14]) ? node12139 : node12134;
												assign node12134 = (inp[4]) ? 15'b000001111111111 : node12135;
													assign node12135 = (inp[8]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node12139 = (inp[8]) ? node12143 : node12140;
													assign node12140 = (inp[2]) ? 15'b000000011111111 : 15'b000001111111111;
													assign node12143 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node12146 = (inp[2]) ? node12154 : node12147;
												assign node12147 = (inp[8]) ? node12151 : node12148;
													assign node12148 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node12151 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node12154 = (inp[8]) ? node12158 : node12155;
													assign node12155 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node12158 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node12161 = (inp[14]) ? node12177 : node12162;
											assign node12162 = (inp[1]) ? node12170 : node12163;
												assign node12163 = (inp[4]) ? node12167 : node12164;
													assign node12164 = (inp[2]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node12167 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node12170 = (inp[5]) ? node12174 : node12171;
													assign node12171 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node12174 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node12177 = (inp[5]) ? node12185 : node12178;
												assign node12178 = (inp[2]) ? node12182 : node12179;
													assign node12179 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node12182 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node12185 = (inp[1]) ? 15'b000000001111111 : node12186;
													assign node12186 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node12190 = (inp[2]) ? node12222 : node12191;
										assign node12191 = (inp[4]) ? node12207 : node12192;
											assign node12192 = (inp[7]) ? node12200 : node12193;
												assign node12193 = (inp[1]) ? node12197 : node12194;
													assign node12194 = (inp[8]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node12197 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node12200 = (inp[14]) ? node12204 : node12201;
													assign node12201 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node12204 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node12207 = (inp[14]) ? node12215 : node12208;
												assign node12208 = (inp[8]) ? node12212 : node12209;
													assign node12209 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node12212 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node12215 = (inp[7]) ? node12219 : node12216;
													assign node12216 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node12219 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node12222 = (inp[1]) ? node12238 : node12223;
											assign node12223 = (inp[5]) ? node12231 : node12224;
												assign node12224 = (inp[8]) ? node12228 : node12225;
													assign node12225 = (inp[7]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node12228 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node12231 = (inp[7]) ? node12235 : node12232;
													assign node12232 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node12235 = (inp[4]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node12238 = (inp[8]) ? node12244 : node12239;
												assign node12239 = (inp[7]) ? node12241 : 15'b000000001111111;
													assign node12241 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node12244 = (inp[5]) ? node12248 : node12245;
													assign node12245 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node12248 = (inp[4]) ? 15'b000000000011111 : 15'b000000000111111;
								assign node12251 = (inp[5]) ? node12315 : node12252;
									assign node12252 = (inp[10]) ? node12284 : node12253;
										assign node12253 = (inp[4]) ? node12269 : node12254;
											assign node12254 = (inp[1]) ? node12262 : node12255;
												assign node12255 = (inp[8]) ? node12259 : node12256;
													assign node12256 = (inp[7]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node12259 = (inp[7]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node12262 = (inp[2]) ? node12266 : node12263;
													assign node12263 = (inp[7]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node12266 = (inp[14]) ? 15'b000000001111111 : 15'b000000111111111;
											assign node12269 = (inp[8]) ? node12277 : node12270;
												assign node12270 = (inp[14]) ? node12274 : node12271;
													assign node12271 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node12274 = (inp[1]) ? 15'b000000001111111 : 15'b000000001111111;
												assign node12277 = (inp[2]) ? node12281 : node12278;
													assign node12278 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node12281 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node12284 = (inp[4]) ? node12300 : node12285;
											assign node12285 = (inp[7]) ? node12293 : node12286;
												assign node12286 = (inp[1]) ? node12290 : node12287;
													assign node12287 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node12290 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node12293 = (inp[2]) ? node12297 : node12294;
													assign node12294 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node12297 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node12300 = (inp[2]) ? node12308 : node12301;
												assign node12301 = (inp[8]) ? node12305 : node12302;
													assign node12302 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node12305 = (inp[7]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node12308 = (inp[7]) ? node12312 : node12309;
													assign node12309 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node12312 = (inp[8]) ? 15'b000000000001111 : 15'b000000000111111;
									assign node12315 = (inp[7]) ? node12345 : node12316;
										assign node12316 = (inp[4]) ? node12330 : node12317;
											assign node12317 = (inp[10]) ? node12323 : node12318;
												assign node12318 = (inp[8]) ? node12320 : 15'b000000011111111;
													assign node12320 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node12323 = (inp[14]) ? node12327 : node12324;
													assign node12324 = (inp[2]) ? 15'b000000001111111 : 15'b000000111111111;
													assign node12327 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node12330 = (inp[8]) ? node12338 : node12331;
												assign node12331 = (inp[10]) ? node12335 : node12332;
													assign node12332 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node12335 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node12338 = (inp[10]) ? node12342 : node12339;
													assign node12339 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node12342 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node12345 = (inp[2]) ? node12359 : node12346;
											assign node12346 = (inp[14]) ? node12352 : node12347;
												assign node12347 = (inp[8]) ? 15'b000000001111111 : node12348;
													assign node12348 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node12352 = (inp[10]) ? node12356 : node12353;
													assign node12353 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node12356 = (inp[1]) ? 15'b000000000011111 : 15'b000000000011111;
											assign node12359 = (inp[4]) ? node12367 : node12360;
												assign node12360 = (inp[10]) ? node12364 : node12361;
													assign node12361 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node12364 = (inp[1]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node12367 = (inp[8]) ? node12371 : node12368;
													assign node12368 = (inp[14]) ? 15'b000000000001111 : 15'b000000000111111;
													assign node12371 = (inp[1]) ? 15'b000000000001111 : 15'b000000000011111;
							assign node12374 = (inp[8]) ? node12494 : node12375;
								assign node12375 = (inp[1]) ? node12437 : node12376;
									assign node12376 = (inp[2]) ? node12406 : node12377;
										assign node12377 = (inp[4]) ? node12391 : node12378;
											assign node12378 = (inp[7]) ? node12384 : node12379;
												assign node12379 = (inp[13]) ? 15'b000000111111111 : node12380;
													assign node12380 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node12384 = (inp[5]) ? node12388 : node12385;
													assign node12385 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node12388 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node12391 = (inp[14]) ? node12399 : node12392;
												assign node12392 = (inp[13]) ? node12396 : node12393;
													assign node12393 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node12396 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node12399 = (inp[5]) ? node12403 : node12400;
													assign node12400 = (inp[13]) ? 15'b000000011111111 : 15'b000000001111111;
													assign node12403 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node12406 = (inp[7]) ? node12422 : node12407;
											assign node12407 = (inp[10]) ? node12415 : node12408;
												assign node12408 = (inp[5]) ? node12412 : node12409;
													assign node12409 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node12412 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node12415 = (inp[13]) ? node12419 : node12416;
													assign node12416 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node12419 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node12422 = (inp[10]) ? node12430 : node12423;
												assign node12423 = (inp[4]) ? node12427 : node12424;
													assign node12424 = (inp[14]) ? 15'b000000000111111 : 15'b000000011111111;
													assign node12427 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node12430 = (inp[13]) ? node12434 : node12431;
													assign node12431 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node12434 = (inp[4]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node12437 = (inp[13]) ? node12463 : node12438;
										assign node12438 = (inp[5]) ? node12454 : node12439;
											assign node12439 = (inp[14]) ? node12447 : node12440;
												assign node12440 = (inp[2]) ? node12444 : node12441;
													assign node12441 = (inp[10]) ? 15'b000000011111111 : 15'b000001111111111;
													assign node12444 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node12447 = (inp[2]) ? node12451 : node12448;
													assign node12448 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node12451 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node12454 = (inp[14]) ? node12460 : node12455;
												assign node12455 = (inp[4]) ? node12457 : 15'b000000001111111;
													assign node12457 = (inp[2]) ? 15'b000000000011111 : 15'b000000001111111;
												assign node12460 = (inp[7]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node12463 = (inp[7]) ? node12479 : node12464;
											assign node12464 = (inp[14]) ? node12472 : node12465;
												assign node12465 = (inp[5]) ? node12469 : node12466;
													assign node12466 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node12469 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node12472 = (inp[10]) ? node12476 : node12473;
													assign node12473 = (inp[5]) ? 15'b000000000111111 : 15'b000000000111111;
													assign node12476 = (inp[4]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node12479 = (inp[5]) ? node12487 : node12480;
												assign node12480 = (inp[2]) ? node12484 : node12481;
													assign node12481 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node12484 = (inp[4]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node12487 = (inp[14]) ? node12491 : node12488;
													assign node12488 = (inp[4]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node12491 = (inp[2]) ? 15'b000000000001111 : 15'b000000000011111;
								assign node12494 = (inp[7]) ? node12558 : node12495;
									assign node12495 = (inp[2]) ? node12527 : node12496;
										assign node12496 = (inp[10]) ? node12512 : node12497;
											assign node12497 = (inp[13]) ? node12505 : node12498;
												assign node12498 = (inp[1]) ? node12502 : node12499;
													assign node12499 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node12502 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node12505 = (inp[14]) ? node12509 : node12506;
													assign node12506 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node12509 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node12512 = (inp[5]) ? node12520 : node12513;
												assign node12513 = (inp[1]) ? node12517 : node12514;
													assign node12514 = (inp[13]) ? 15'b000000000111111 : 15'b000000011111111;
													assign node12517 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node12520 = (inp[14]) ? node12524 : node12521;
													assign node12521 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node12524 = (inp[13]) ? 15'b000000000001111 : 15'b000000000111111;
										assign node12527 = (inp[13]) ? node12543 : node12528;
											assign node12528 = (inp[10]) ? node12536 : node12529;
												assign node12529 = (inp[14]) ? node12533 : node12530;
													assign node12530 = (inp[1]) ? 15'b000000001111111 : 15'b000000111111111;
													assign node12533 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node12536 = (inp[14]) ? node12540 : node12537;
													assign node12537 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node12540 = (inp[1]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node12543 = (inp[10]) ? node12551 : node12544;
												assign node12544 = (inp[4]) ? node12548 : node12545;
													assign node12545 = (inp[5]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node12548 = (inp[5]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node12551 = (inp[1]) ? node12555 : node12552;
													assign node12552 = (inp[14]) ? 15'b000000000011111 : 15'b000000000011111;
													assign node12555 = (inp[14]) ? 15'b000000000001111 : 15'b000000000011111;
									assign node12558 = (inp[5]) ? node12590 : node12559;
										assign node12559 = (inp[4]) ? node12575 : node12560;
											assign node12560 = (inp[13]) ? node12568 : node12561;
												assign node12561 = (inp[10]) ? node12565 : node12562;
													assign node12562 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node12565 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node12568 = (inp[10]) ? node12572 : node12569;
													assign node12569 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node12572 = (inp[14]) ? 15'b000000000011111 : 15'b000000000011111;
											assign node12575 = (inp[2]) ? node12583 : node12576;
												assign node12576 = (inp[1]) ? node12580 : node12577;
													assign node12577 = (inp[14]) ? 15'b000000000111111 : 15'b000000000111111;
													assign node12580 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node12583 = (inp[14]) ? node12587 : node12584;
													assign node12584 = (inp[10]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node12587 = (inp[10]) ? 15'b000000000001111 : 15'b000000000011111;
										assign node12590 = (inp[10]) ? node12604 : node12591;
											assign node12591 = (inp[14]) ? node12599 : node12592;
												assign node12592 = (inp[13]) ? node12596 : node12593;
													assign node12593 = (inp[2]) ? 15'b000000000111111 : 15'b000000000111111;
													assign node12596 = (inp[4]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node12599 = (inp[2]) ? node12601 : 15'b000000000011111;
													assign node12601 = (inp[4]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node12604 = (inp[13]) ? node12612 : node12605;
												assign node12605 = (inp[2]) ? node12609 : node12606;
													assign node12606 = (inp[4]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node12609 = (inp[4]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node12612 = (inp[4]) ? node12616 : node12613;
													assign node12613 = (inp[1]) ? 15'b000000000001111 : 15'b000000000011111;
													assign node12616 = (inp[2]) ? 15'b000000000000111 : 15'b000000000001111;
					assign node12619 = (inp[7]) ? node13101 : node12620;
						assign node12620 = (inp[5]) ? node12860 : node12621;
							assign node12621 = (inp[1]) ? node12743 : node12622;
								assign node12622 = (inp[4]) ? node12682 : node12623;
									assign node12623 = (inp[8]) ? node12651 : node12624;
										assign node12624 = (inp[14]) ? node12638 : node12625;
											assign node12625 = (inp[13]) ? node12631 : node12626;
												assign node12626 = (inp[2]) ? 15'b000001111111111 : node12627;
													assign node12627 = (inp[9]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node12631 = (inp[2]) ? node12635 : node12632;
													assign node12632 = (inp[10]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node12635 = (inp[9]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node12638 = (inp[13]) ? node12646 : node12639;
												assign node12639 = (inp[11]) ? node12643 : node12640;
													assign node12640 = (inp[10]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node12643 = (inp[9]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node12646 = (inp[11]) ? 15'b000000011111111 : node12647;
													assign node12647 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node12651 = (inp[2]) ? node12667 : node12652;
											assign node12652 = (inp[9]) ? node12660 : node12653;
												assign node12653 = (inp[11]) ? node12657 : node12654;
													assign node12654 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node12657 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node12660 = (inp[11]) ? node12664 : node12661;
													assign node12661 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node12664 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node12667 = (inp[13]) ? node12675 : node12668;
												assign node12668 = (inp[11]) ? node12672 : node12669;
													assign node12669 = (inp[9]) ? 15'b000000011111111 : 15'b000001111111111;
													assign node12672 = (inp[9]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node12675 = (inp[9]) ? node12679 : node12676;
													assign node12676 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node12679 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node12682 = (inp[10]) ? node12712 : node12683;
										assign node12683 = (inp[9]) ? node12697 : node12684;
											assign node12684 = (inp[11]) ? node12692 : node12685;
												assign node12685 = (inp[14]) ? node12689 : node12686;
													assign node12686 = (inp[2]) ? 15'b000000111111111 : 15'b000011111111111;
													assign node12689 = (inp[2]) ? 15'b000000001111111 : 15'b000000111111111;
												assign node12692 = (inp[14]) ? 15'b000000011111111 : node12693;
													assign node12693 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node12697 = (inp[13]) ? node12705 : node12698;
												assign node12698 = (inp[11]) ? node12702 : node12699;
													assign node12699 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node12702 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node12705 = (inp[8]) ? node12709 : node12706;
													assign node12706 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node12709 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node12712 = (inp[2]) ? node12728 : node12713;
											assign node12713 = (inp[9]) ? node12721 : node12714;
												assign node12714 = (inp[13]) ? node12718 : node12715;
													assign node12715 = (inp[11]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node12718 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node12721 = (inp[13]) ? node12725 : node12722;
													assign node12722 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node12725 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node12728 = (inp[11]) ? node12736 : node12729;
												assign node12729 = (inp[9]) ? node12733 : node12730;
													assign node12730 = (inp[13]) ? 15'b000000001111111 : 15'b000000001111111;
													assign node12733 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node12736 = (inp[14]) ? node12740 : node12737;
													assign node12737 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node12740 = (inp[13]) ? 15'b000000000011111 : 15'b000000000111111;
								assign node12743 = (inp[9]) ? node12805 : node12744;
									assign node12744 = (inp[11]) ? node12776 : node12745;
										assign node12745 = (inp[14]) ? node12761 : node12746;
											assign node12746 = (inp[13]) ? node12754 : node12747;
												assign node12747 = (inp[10]) ? node12751 : node12748;
													assign node12748 = (inp[2]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node12751 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node12754 = (inp[4]) ? node12758 : node12755;
													assign node12755 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node12758 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node12761 = (inp[10]) ? node12769 : node12762;
												assign node12762 = (inp[13]) ? node12766 : node12763;
													assign node12763 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node12766 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node12769 = (inp[4]) ? node12773 : node12770;
													assign node12770 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node12773 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node12776 = (inp[14]) ? node12792 : node12777;
											assign node12777 = (inp[10]) ? node12785 : node12778;
												assign node12778 = (inp[4]) ? node12782 : node12779;
													assign node12779 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node12782 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node12785 = (inp[2]) ? node12789 : node12786;
													assign node12786 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node12789 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node12792 = (inp[4]) ? node12800 : node12793;
												assign node12793 = (inp[2]) ? node12797 : node12794;
													assign node12794 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node12797 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node12800 = (inp[10]) ? node12802 : 15'b000000000111111;
													assign node12802 = (inp[2]) ? 15'b000000000001111 : 15'b000000000011111;
									assign node12805 = (inp[14]) ? node12831 : node12806;
										assign node12806 = (inp[13]) ? node12818 : node12807;
											assign node12807 = (inp[8]) ? node12813 : node12808;
												assign node12808 = (inp[10]) ? node12810 : 15'b000000011111111;
													assign node12810 = (inp[4]) ? 15'b000000001111111 : 15'b000000111111111;
												assign node12813 = (inp[4]) ? 15'b000000001111111 : node12814;
													assign node12814 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node12818 = (inp[8]) ? node12824 : node12819;
												assign node12819 = (inp[10]) ? node12821 : 15'b000000001111111;
													assign node12821 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node12824 = (inp[11]) ? node12828 : node12825;
													assign node12825 = (inp[4]) ? 15'b000000000111111 : 15'b000000011111111;
													assign node12828 = (inp[2]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node12831 = (inp[13]) ? node12847 : node12832;
											assign node12832 = (inp[2]) ? node12840 : node12833;
												assign node12833 = (inp[4]) ? node12837 : node12834;
													assign node12834 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node12837 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node12840 = (inp[4]) ? node12844 : node12841;
													assign node12841 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node12844 = (inp[10]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node12847 = (inp[2]) ? node12855 : node12848;
												assign node12848 = (inp[10]) ? node12852 : node12849;
													assign node12849 = (inp[8]) ? 15'b000000000111111 : 15'b000000000111111;
													assign node12852 = (inp[4]) ? 15'b000000000001111 : 15'b000000000111111;
												assign node12855 = (inp[4]) ? 15'b000000000011111 : node12856;
													assign node12856 = (inp[8]) ? 15'b000000000011111 : 15'b000000000111111;
							assign node12860 = (inp[2]) ? node12982 : node12861;
								assign node12861 = (inp[4]) ? node12921 : node12862;
									assign node12862 = (inp[8]) ? node12894 : node12863;
										assign node12863 = (inp[1]) ? node12879 : node12864;
											assign node12864 = (inp[9]) ? node12872 : node12865;
												assign node12865 = (inp[10]) ? node12869 : node12866;
													assign node12866 = (inp[13]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node12869 = (inp[11]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node12872 = (inp[11]) ? node12876 : node12873;
													assign node12873 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node12876 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node12879 = (inp[11]) ? node12887 : node12880;
												assign node12880 = (inp[14]) ? node12884 : node12881;
													assign node12881 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node12884 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node12887 = (inp[10]) ? node12891 : node12888;
													assign node12888 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node12891 = (inp[9]) ? 15'b000000000111111 : 15'b000000000111111;
										assign node12894 = (inp[13]) ? node12910 : node12895;
											assign node12895 = (inp[9]) ? node12903 : node12896;
												assign node12896 = (inp[11]) ? node12900 : node12897;
													assign node12897 = (inp[14]) ? 15'b000000011111111 : 15'b000000011111111;
													assign node12900 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node12903 = (inp[11]) ? node12907 : node12904;
													assign node12904 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node12907 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node12910 = (inp[11]) ? node12918 : node12911;
												assign node12911 = (inp[10]) ? node12915 : node12912;
													assign node12912 = (inp[9]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node12915 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node12918 = (inp[9]) ? 15'b000000000001111 : 15'b000000000111111;
									assign node12921 = (inp[1]) ? node12951 : node12922;
										assign node12922 = (inp[14]) ? node12936 : node12923;
											assign node12923 = (inp[9]) ? node12929 : node12924;
												assign node12924 = (inp[10]) ? node12926 : 15'b000000011111111;
													assign node12926 = (inp[11]) ? 15'b000000011111111 : 15'b000000011111111;
												assign node12929 = (inp[11]) ? node12933 : node12930;
													assign node12930 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node12933 = (inp[8]) ? 15'b000000000011111 : 15'b000000001111111;
											assign node12936 = (inp[13]) ? node12944 : node12937;
												assign node12937 = (inp[9]) ? node12941 : node12938;
													assign node12938 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node12941 = (inp[10]) ? 15'b000000000111111 : 15'b000000000111111;
												assign node12944 = (inp[11]) ? node12948 : node12945;
													assign node12945 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node12948 = (inp[8]) ? 15'b000000000001111 : 15'b000000000111111;
										assign node12951 = (inp[13]) ? node12967 : node12952;
											assign node12952 = (inp[8]) ? node12960 : node12953;
												assign node12953 = (inp[11]) ? node12957 : node12954;
													assign node12954 = (inp[10]) ? 15'b000000001111111 : 15'b000000001111111;
													assign node12957 = (inp[9]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node12960 = (inp[10]) ? node12964 : node12961;
													assign node12961 = (inp[11]) ? 15'b000000000111111 : 15'b000000000111111;
													assign node12964 = (inp[11]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node12967 = (inp[11]) ? node12975 : node12968;
												assign node12968 = (inp[10]) ? node12972 : node12969;
													assign node12969 = (inp[9]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node12972 = (inp[8]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node12975 = (inp[8]) ? node12979 : node12976;
													assign node12976 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node12979 = (inp[14]) ? 15'b000000000001111 : 15'b000000000011111;
								assign node12982 = (inp[9]) ? node13042 : node12983;
									assign node12983 = (inp[8]) ? node13015 : node12984;
										assign node12984 = (inp[14]) ? node13000 : node12985;
											assign node12985 = (inp[4]) ? node12993 : node12986;
												assign node12986 = (inp[13]) ? node12990 : node12987;
													assign node12987 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node12990 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node12993 = (inp[11]) ? node12997 : node12994;
													assign node12994 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node12997 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node13000 = (inp[11]) ? node13008 : node13001;
												assign node13001 = (inp[1]) ? node13005 : node13002;
													assign node13002 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node13005 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node13008 = (inp[1]) ? node13012 : node13009;
													assign node13009 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node13012 = (inp[10]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node13015 = (inp[10]) ? node13029 : node13016;
											assign node13016 = (inp[1]) ? node13022 : node13017;
												assign node13017 = (inp[4]) ? node13019 : 15'b000000001111111;
													assign node13019 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node13022 = (inp[11]) ? node13026 : node13023;
													assign node13023 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node13026 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node13029 = (inp[13]) ? node13035 : node13030;
												assign node13030 = (inp[14]) ? node13032 : 15'b000000001111111;
													assign node13032 = (inp[1]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node13035 = (inp[14]) ? node13039 : node13036;
													assign node13036 = (inp[11]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node13039 = (inp[4]) ? 15'b000000000001111 : 15'b000000000011111;
									assign node13042 = (inp[13]) ? node13072 : node13043;
										assign node13043 = (inp[8]) ? node13057 : node13044;
											assign node13044 = (inp[14]) ? node13050 : node13045;
												assign node13045 = (inp[11]) ? 15'b000000000111111 : node13046;
													assign node13046 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node13050 = (inp[1]) ? node13054 : node13051;
													assign node13051 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node13054 = (inp[10]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node13057 = (inp[14]) ? node13065 : node13058;
												assign node13058 = (inp[1]) ? node13062 : node13059;
													assign node13059 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node13062 = (inp[4]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node13065 = (inp[10]) ? node13069 : node13066;
													assign node13066 = (inp[4]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node13069 = (inp[4]) ? 15'b000000000001111 : 15'b000000000011111;
										assign node13072 = (inp[8]) ? node13086 : node13073;
											assign node13073 = (inp[1]) ? node13081 : node13074;
												assign node13074 = (inp[14]) ? node13078 : node13075;
													assign node13075 = (inp[11]) ? 15'b000000000111111 : 15'b000000000111111;
													assign node13078 = (inp[10]) ? 15'b000000000011111 : 15'b000000000011111;
												assign node13081 = (inp[14]) ? node13083 : 15'b000000000011111;
													assign node13083 = (inp[4]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node13086 = (inp[14]) ? node13094 : node13087;
												assign node13087 = (inp[4]) ? node13091 : node13088;
													assign node13088 = (inp[11]) ? 15'b000000000001111 : 15'b000000000111111;
													assign node13091 = (inp[1]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node13094 = (inp[10]) ? node13098 : node13095;
													assign node13095 = (inp[11]) ? 15'b000000000001111 : 15'b000000000011111;
													assign node13098 = (inp[11]) ? 15'b000000000000111 : 15'b000000000001111;
						assign node13101 = (inp[4]) ? node13353 : node13102;
							assign node13102 = (inp[14]) ? node13228 : node13103;
								assign node13103 = (inp[1]) ? node13165 : node13104;
									assign node13104 = (inp[9]) ? node13134 : node13105;
										assign node13105 = (inp[13]) ? node13119 : node13106;
											assign node13106 = (inp[2]) ? node13112 : node13107;
												assign node13107 = (inp[5]) ? 15'b000000111111111 : node13108;
													assign node13108 = (inp[11]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node13112 = (inp[8]) ? node13116 : node13113;
													assign node13113 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node13116 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node13119 = (inp[8]) ? node13127 : node13120;
												assign node13120 = (inp[5]) ? node13124 : node13121;
													assign node13121 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node13124 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node13127 = (inp[2]) ? node13131 : node13128;
													assign node13128 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node13131 = (inp[5]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node13134 = (inp[11]) ? node13150 : node13135;
											assign node13135 = (inp[8]) ? node13143 : node13136;
												assign node13136 = (inp[13]) ? node13140 : node13137;
													assign node13137 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node13140 = (inp[5]) ? 15'b000000000111111 : 15'b000000011111111;
												assign node13143 = (inp[5]) ? node13147 : node13144;
													assign node13144 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node13147 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node13150 = (inp[2]) ? node13158 : node13151;
												assign node13151 = (inp[8]) ? node13155 : node13152;
													assign node13152 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node13155 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node13158 = (inp[5]) ? node13162 : node13159;
													assign node13159 = (inp[10]) ? 15'b000000000011111 : 15'b000000001111111;
													assign node13162 = (inp[8]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node13165 = (inp[10]) ? node13197 : node13166;
										assign node13166 = (inp[2]) ? node13182 : node13167;
											assign node13167 = (inp[9]) ? node13175 : node13168;
												assign node13168 = (inp[13]) ? node13172 : node13169;
													assign node13169 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node13172 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node13175 = (inp[13]) ? node13179 : node13176;
													assign node13176 = (inp[5]) ? 15'b000000001111111 : 15'b000000001111111;
													assign node13179 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node13182 = (inp[13]) ? node13190 : node13183;
												assign node13183 = (inp[11]) ? node13187 : node13184;
													assign node13184 = (inp[9]) ? 15'b000000001111111 : 15'b000000111111111;
													assign node13187 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node13190 = (inp[5]) ? node13194 : node13191;
													assign node13191 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node13194 = (inp[8]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node13197 = (inp[8]) ? node13213 : node13198;
											assign node13198 = (inp[9]) ? node13206 : node13199;
												assign node13199 = (inp[13]) ? node13203 : node13200;
													assign node13200 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node13203 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node13206 = (inp[2]) ? node13210 : node13207;
													assign node13207 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node13210 = (inp[11]) ? 15'b000000000001111 : 15'b000000000111111;
											assign node13213 = (inp[5]) ? node13221 : node13214;
												assign node13214 = (inp[13]) ? node13218 : node13215;
													assign node13215 = (inp[2]) ? 15'b000000000011111 : 15'b000000001111111;
													assign node13218 = (inp[11]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node13221 = (inp[2]) ? node13225 : node13222;
													assign node13222 = (inp[9]) ? 15'b000000000011111 : 15'b000000000011111;
													assign node13225 = (inp[11]) ? 15'b000000000001111 : 15'b000000000011111;
								assign node13228 = (inp[11]) ? node13290 : node13229;
									assign node13229 = (inp[10]) ? node13259 : node13230;
										assign node13230 = (inp[8]) ? node13244 : node13231;
											assign node13231 = (inp[5]) ? node13239 : node13232;
												assign node13232 = (inp[2]) ? node13236 : node13233;
													assign node13233 = (inp[13]) ? 15'b000000111111111 : 15'b000000111111111;
													assign node13236 = (inp[9]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node13239 = (inp[2]) ? 15'b000000000111111 : node13240;
													assign node13240 = (inp[9]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node13244 = (inp[5]) ? node13252 : node13245;
												assign node13245 = (inp[1]) ? node13249 : node13246;
													assign node13246 = (inp[13]) ? 15'b000000001111111 : 15'b000000111111111;
													assign node13249 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node13252 = (inp[13]) ? node13256 : node13253;
													assign node13253 = (inp[9]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node13256 = (inp[1]) ? 15'b000000000111111 : 15'b000000000111111;
										assign node13259 = (inp[9]) ? node13275 : node13260;
											assign node13260 = (inp[1]) ? node13268 : node13261;
												assign node13261 = (inp[13]) ? node13265 : node13262;
													assign node13262 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node13265 = (inp[5]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node13268 = (inp[5]) ? node13272 : node13269;
													assign node13269 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node13272 = (inp[13]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node13275 = (inp[5]) ? node13283 : node13276;
												assign node13276 = (inp[13]) ? node13280 : node13277;
													assign node13277 = (inp[1]) ? 15'b000000000111111 : 15'b000000000111111;
													assign node13280 = (inp[2]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node13283 = (inp[2]) ? node13287 : node13284;
													assign node13284 = (inp[8]) ? 15'b000000000001111 : 15'b000000000111111;
													assign node13287 = (inp[13]) ? 15'b000000000001111 : 15'b000000000001111;
									assign node13290 = (inp[1]) ? node13322 : node13291;
										assign node13291 = (inp[10]) ? node13307 : node13292;
											assign node13292 = (inp[9]) ? node13300 : node13293;
												assign node13293 = (inp[2]) ? node13297 : node13294;
													assign node13294 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node13297 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node13300 = (inp[5]) ? node13304 : node13301;
													assign node13301 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node13304 = (inp[2]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node13307 = (inp[5]) ? node13315 : node13308;
												assign node13308 = (inp[9]) ? node13312 : node13309;
													assign node13309 = (inp[8]) ? 15'b000000000111111 : 15'b000000000111111;
													assign node13312 = (inp[8]) ? 15'b000000000011111 : 15'b000000000011111;
												assign node13315 = (inp[13]) ? node13319 : node13316;
													assign node13316 = (inp[8]) ? 15'b000000000011111 : 15'b000000000011111;
													assign node13319 = (inp[8]) ? 15'b000000000001111 : 15'b000000000001111;
										assign node13322 = (inp[13]) ? node13338 : node13323;
											assign node13323 = (inp[9]) ? node13331 : node13324;
												assign node13324 = (inp[10]) ? node13328 : node13325;
													assign node13325 = (inp[8]) ? 15'b000000000111111 : 15'b000000011111111;
													assign node13328 = (inp[8]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node13331 = (inp[8]) ? node13335 : node13332;
													assign node13332 = (inp[10]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node13335 = (inp[10]) ? 15'b000000000000111 : 15'b000000000011111;
											assign node13338 = (inp[5]) ? node13346 : node13339;
												assign node13339 = (inp[2]) ? node13343 : node13340;
													assign node13340 = (inp[9]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node13343 = (inp[8]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node13346 = (inp[9]) ? node13350 : node13347;
													assign node13347 = (inp[10]) ? 15'b000000000001111 : 15'b000000000011111;
													assign node13350 = (inp[2]) ? 15'b000000000000111 : 15'b000000000001111;
							assign node13353 = (inp[10]) ? node13477 : node13354;
								assign node13354 = (inp[9]) ? node13416 : node13355;
									assign node13355 = (inp[14]) ? node13387 : node13356;
										assign node13356 = (inp[8]) ? node13372 : node13357;
											assign node13357 = (inp[11]) ? node13365 : node13358;
												assign node13358 = (inp[2]) ? node13362 : node13359;
													assign node13359 = (inp[5]) ? 15'b000000011111111 : 15'b000000011111111;
													assign node13362 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node13365 = (inp[1]) ? node13369 : node13366;
													assign node13366 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node13369 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node13372 = (inp[2]) ? node13380 : node13373;
												assign node13373 = (inp[11]) ? node13377 : node13374;
													assign node13374 = (inp[1]) ? 15'b000000001111111 : 15'b000000001111111;
													assign node13377 = (inp[1]) ? 15'b000000000111111 : 15'b000000000111111;
												assign node13380 = (inp[13]) ? node13384 : node13381;
													assign node13381 = (inp[1]) ? 15'b000000000111111 : 15'b000000011111111;
													assign node13384 = (inp[5]) ? 15'b000000000011111 : 15'b000000000011111;
										assign node13387 = (inp[5]) ? node13401 : node13388;
											assign node13388 = (inp[13]) ? node13394 : node13389;
												assign node13389 = (inp[8]) ? node13391 : 15'b000000001111111;
													assign node13391 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node13394 = (inp[1]) ? node13398 : node13395;
													assign node13395 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node13398 = (inp[8]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node13401 = (inp[11]) ? node13409 : node13402;
												assign node13402 = (inp[2]) ? node13406 : node13403;
													assign node13403 = (inp[13]) ? 15'b000000000111111 : 15'b000000000111111;
													assign node13406 = (inp[13]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node13409 = (inp[8]) ? node13413 : node13410;
													assign node13410 = (inp[13]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node13413 = (inp[1]) ? 15'b000000000001111 : 15'b000000000011111;
									assign node13416 = (inp[1]) ? node13446 : node13417;
										assign node13417 = (inp[8]) ? node13431 : node13418;
											assign node13418 = (inp[5]) ? node13426 : node13419;
												assign node13419 = (inp[14]) ? node13423 : node13420;
													assign node13420 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node13423 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node13426 = (inp[14]) ? node13428 : 15'b000000000111111;
													assign node13428 = (inp[2]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node13431 = (inp[2]) ? node13439 : node13432;
												assign node13432 = (inp[13]) ? node13436 : node13433;
													assign node13433 = (inp[14]) ? 15'b000000000111111 : 15'b000000000111111;
													assign node13436 = (inp[11]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node13439 = (inp[11]) ? node13443 : node13440;
													assign node13440 = (inp[13]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node13443 = (inp[14]) ? 15'b000000000001111 : 15'b000000000011111;
										assign node13446 = (inp[8]) ? node13462 : node13447;
											assign node13447 = (inp[2]) ? node13455 : node13448;
												assign node13448 = (inp[14]) ? node13452 : node13449;
													assign node13449 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node13452 = (inp[5]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node13455 = (inp[11]) ? node13459 : node13456;
													assign node13456 = (inp[5]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node13459 = (inp[13]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node13462 = (inp[11]) ? node13470 : node13463;
												assign node13463 = (inp[5]) ? node13467 : node13464;
													assign node13464 = (inp[2]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node13467 = (inp[2]) ? 15'b000000000001111 : 15'b000000000001111;
												assign node13470 = (inp[13]) ? node13474 : node13471;
													assign node13471 = (inp[14]) ? 15'b000000000001111 : 15'b000000000011111;
													assign node13474 = (inp[2]) ? 15'b000000000000111 : 15'b000000000001111;
								assign node13477 = (inp[9]) ? node13539 : node13478;
									assign node13478 = (inp[13]) ? node13508 : node13479;
										assign node13479 = (inp[2]) ? node13495 : node13480;
											assign node13480 = (inp[14]) ? node13488 : node13481;
												assign node13481 = (inp[5]) ? node13485 : node13482;
													assign node13482 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node13485 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node13488 = (inp[11]) ? node13492 : node13489;
													assign node13489 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node13492 = (inp[5]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node13495 = (inp[11]) ? node13503 : node13496;
												assign node13496 = (inp[8]) ? node13500 : node13497;
													assign node13497 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node13500 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node13503 = (inp[5]) ? node13505 : 15'b000000000011111;
													assign node13505 = (inp[8]) ? 15'b000000000000111 : 15'b000000000001111;
										assign node13508 = (inp[1]) ? node13524 : node13509;
											assign node13509 = (inp[11]) ? node13517 : node13510;
												assign node13510 = (inp[8]) ? node13514 : node13511;
													assign node13511 = (inp[5]) ? 15'b000000000111111 : 15'b000000000111111;
													assign node13514 = (inp[2]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node13517 = (inp[14]) ? node13521 : node13518;
													assign node13518 = (inp[8]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node13521 = (inp[8]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node13524 = (inp[2]) ? node13532 : node13525;
												assign node13525 = (inp[11]) ? node13529 : node13526;
													assign node13526 = (inp[5]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node13529 = (inp[8]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node13532 = (inp[5]) ? node13536 : node13533;
													assign node13533 = (inp[8]) ? 15'b000000000001111 : 15'b000000000011111;
													assign node13536 = (inp[8]) ? 15'b000000000000111 : 15'b000000000001111;
									assign node13539 = (inp[5]) ? node13567 : node13540;
										assign node13540 = (inp[11]) ? node13552 : node13541;
											assign node13541 = (inp[1]) ? node13547 : node13542;
												assign node13542 = (inp[2]) ? node13544 : 15'b000000001111111;
													assign node13544 = (inp[8]) ? 15'b000000000011111 : 15'b000000000011111;
												assign node13547 = (inp[8]) ? node13549 : 15'b000000000011111;
													assign node13549 = (inp[2]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node13552 = (inp[13]) ? node13560 : node13553;
												assign node13553 = (inp[14]) ? node13557 : node13554;
													assign node13554 = (inp[8]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node13557 = (inp[1]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node13560 = (inp[1]) ? node13564 : node13561;
													assign node13561 = (inp[2]) ? 15'b000000000001111 : 15'b000000000001111;
													assign node13564 = (inp[8]) ? 15'b000000000000011 : 15'b000000000001111;
										assign node13567 = (inp[14]) ? node13581 : node13568;
											assign node13568 = (inp[11]) ? node13576 : node13569;
												assign node13569 = (inp[1]) ? node13573 : node13570;
													assign node13570 = (inp[2]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node13573 = (inp[13]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node13576 = (inp[8]) ? node13578 : 15'b000000000011111;
													assign node13578 = (inp[2]) ? 15'b000000000000111 : 15'b000000000001111;
											assign node13581 = (inp[2]) ? node13589 : node13582;
												assign node13582 = (inp[1]) ? node13586 : node13583;
													assign node13583 = (inp[11]) ? 15'b000000000000111 : 15'b000000000011111;
													assign node13586 = (inp[13]) ? 15'b000000000000111 : 15'b000000000001111;
												assign node13589 = (inp[8]) ? node13593 : node13590;
													assign node13590 = (inp[1]) ? 15'b000000000000111 : 15'b000000000001111;
													assign node13593 = (inp[13]) ? 15'b000000000000001 : 15'b000000000000111;
				assign node13596 = (inp[11]) ? node14574 : node13597;
					assign node13597 = (inp[8]) ? node14085 : node13598;
						assign node13598 = (inp[7]) ? node13838 : node13599;
							assign node13599 = (inp[9]) ? node13721 : node13600;
								assign node13600 = (inp[10]) ? node13662 : node13601;
									assign node13601 = (inp[13]) ? node13631 : node13602;
										assign node13602 = (inp[12]) ? node13618 : node13603;
											assign node13603 = (inp[1]) ? node13611 : node13604;
												assign node13604 = (inp[2]) ? node13608 : node13605;
													assign node13605 = (inp[4]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node13608 = (inp[4]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node13611 = (inp[14]) ? node13615 : node13612;
													assign node13612 = (inp[2]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node13615 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node13618 = (inp[1]) ? node13624 : node13619;
												assign node13619 = (inp[14]) ? node13621 : 15'b000001111111111;
													assign node13621 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node13624 = (inp[2]) ? node13628 : node13625;
													assign node13625 = (inp[4]) ? 15'b000000011111111 : 15'b000000011111111;
													assign node13628 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node13631 = (inp[4]) ? node13647 : node13632;
											assign node13632 = (inp[2]) ? node13640 : node13633;
												assign node13633 = (inp[5]) ? node13637 : node13634;
													assign node13634 = (inp[12]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node13637 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node13640 = (inp[12]) ? node13644 : node13641;
													assign node13641 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node13644 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node13647 = (inp[1]) ? node13655 : node13648;
												assign node13648 = (inp[2]) ? node13652 : node13649;
													assign node13649 = (inp[12]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node13652 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node13655 = (inp[12]) ? node13659 : node13656;
													assign node13656 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node13659 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node13662 = (inp[2]) ? node13692 : node13663;
										assign node13663 = (inp[13]) ? node13677 : node13664;
											assign node13664 = (inp[5]) ? node13670 : node13665;
												assign node13665 = (inp[14]) ? 15'b000000111111111 : node13666;
													assign node13666 = (inp[1]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node13670 = (inp[1]) ? node13674 : node13671;
													assign node13671 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node13674 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node13677 = (inp[1]) ? node13685 : node13678;
												assign node13678 = (inp[14]) ? node13682 : node13679;
													assign node13679 = (inp[12]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node13682 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node13685 = (inp[4]) ? node13689 : node13686;
													assign node13686 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node13689 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node13692 = (inp[14]) ? node13708 : node13693;
											assign node13693 = (inp[5]) ? node13701 : node13694;
												assign node13694 = (inp[13]) ? node13698 : node13695;
													assign node13695 = (inp[12]) ? 15'b000000001111111 : 15'b000000111111111;
													assign node13698 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node13701 = (inp[13]) ? node13705 : node13702;
													assign node13702 = (inp[4]) ? 15'b000000001111111 : 15'b000000001111111;
													assign node13705 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node13708 = (inp[1]) ? node13716 : node13709;
												assign node13709 = (inp[12]) ? node13713 : node13710;
													assign node13710 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node13713 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node13716 = (inp[5]) ? 15'b000000000011111 : node13717;
													assign node13717 = (inp[13]) ? 15'b000000000111111 : 15'b000000000111111;
								assign node13721 = (inp[14]) ? node13779 : node13722;
									assign node13722 = (inp[5]) ? node13752 : node13723;
										assign node13723 = (inp[1]) ? node13737 : node13724;
											assign node13724 = (inp[4]) ? node13732 : node13725;
												assign node13725 = (inp[13]) ? node13729 : node13726;
													assign node13726 = (inp[10]) ? 15'b000001111111111 : 15'b000001111111111;
													assign node13729 = (inp[12]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node13732 = (inp[10]) ? node13734 : 15'b000000011111111;
													assign node13734 = (inp[13]) ? 15'b000000001111111 : 15'b000000001111111;
											assign node13737 = (inp[13]) ? node13745 : node13738;
												assign node13738 = (inp[2]) ? node13742 : node13739;
													assign node13739 = (inp[12]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node13742 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node13745 = (inp[12]) ? node13749 : node13746;
													assign node13746 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node13749 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node13752 = (inp[13]) ? node13764 : node13753;
											assign node13753 = (inp[1]) ? node13759 : node13754;
												assign node13754 = (inp[10]) ? node13756 : 15'b000000111111111;
													assign node13756 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node13759 = (inp[4]) ? 15'b000000000111111 : node13760;
													assign node13760 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node13764 = (inp[10]) ? node13772 : node13765;
												assign node13765 = (inp[2]) ? node13769 : node13766;
													assign node13766 = (inp[1]) ? 15'b000000001111111 : 15'b000000111111111;
													assign node13769 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node13772 = (inp[12]) ? node13776 : node13773;
													assign node13773 = (inp[4]) ? 15'b000000000111111 : 15'b000000000111111;
													assign node13776 = (inp[1]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node13779 = (inp[13]) ? node13809 : node13780;
										assign node13780 = (inp[2]) ? node13794 : node13781;
											assign node13781 = (inp[10]) ? node13789 : node13782;
												assign node13782 = (inp[12]) ? node13786 : node13783;
													assign node13783 = (inp[5]) ? 15'b000000011111111 : 15'b000000011111111;
													assign node13786 = (inp[5]) ? 15'b000000000111111 : 15'b000000011111111;
												assign node13789 = (inp[1]) ? 15'b000000001111111 : node13790;
													assign node13790 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node13794 = (inp[4]) ? node13802 : node13795;
												assign node13795 = (inp[1]) ? node13799 : node13796;
													assign node13796 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node13799 = (inp[5]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node13802 = (inp[10]) ? node13806 : node13803;
													assign node13803 = (inp[5]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node13806 = (inp[5]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node13809 = (inp[12]) ? node13825 : node13810;
											assign node13810 = (inp[4]) ? node13818 : node13811;
												assign node13811 = (inp[1]) ? node13815 : node13812;
													assign node13812 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node13815 = (inp[5]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node13818 = (inp[1]) ? node13822 : node13819;
													assign node13819 = (inp[10]) ? 15'b000000000011111 : 15'b000000001111111;
													assign node13822 = (inp[5]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node13825 = (inp[2]) ? node13831 : node13826;
												assign node13826 = (inp[10]) ? node13828 : 15'b000000000111111;
													assign node13828 = (inp[1]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node13831 = (inp[4]) ? node13835 : node13832;
													assign node13832 = (inp[10]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node13835 = (inp[1]) ? 15'b000000000001111 : 15'b000000000001111;
							assign node13838 = (inp[4]) ? node13962 : node13839;
								assign node13839 = (inp[10]) ? node13903 : node13840;
									assign node13840 = (inp[14]) ? node13872 : node13841;
										assign node13841 = (inp[2]) ? node13857 : node13842;
											assign node13842 = (inp[5]) ? node13850 : node13843;
												assign node13843 = (inp[13]) ? node13847 : node13844;
													assign node13844 = (inp[9]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node13847 = (inp[9]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node13850 = (inp[12]) ? node13854 : node13851;
													assign node13851 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node13854 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node13857 = (inp[13]) ? node13865 : node13858;
												assign node13858 = (inp[5]) ? node13862 : node13859;
													assign node13859 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node13862 = (inp[9]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node13865 = (inp[1]) ? node13869 : node13866;
													assign node13866 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node13869 = (inp[9]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node13872 = (inp[13]) ? node13888 : node13873;
											assign node13873 = (inp[2]) ? node13881 : node13874;
												assign node13874 = (inp[1]) ? node13878 : node13875;
													assign node13875 = (inp[5]) ? 15'b000000001111111 : 15'b000000111111111;
													assign node13878 = (inp[9]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node13881 = (inp[9]) ? node13885 : node13882;
													assign node13882 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node13885 = (inp[5]) ? 15'b000000000011111 : 15'b000000001111111;
											assign node13888 = (inp[2]) ? node13896 : node13889;
												assign node13889 = (inp[12]) ? node13893 : node13890;
													assign node13890 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node13893 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node13896 = (inp[9]) ? node13900 : node13897;
													assign node13897 = (inp[5]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node13900 = (inp[12]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node13903 = (inp[2]) ? node13931 : node13904;
										assign node13904 = (inp[5]) ? node13916 : node13905;
											assign node13905 = (inp[1]) ? node13911 : node13906;
												assign node13906 = (inp[13]) ? node13908 : 15'b000000011111111;
													assign node13908 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node13911 = (inp[12]) ? 15'b000000001111111 : node13912;
													assign node13912 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node13916 = (inp[1]) ? node13924 : node13917;
												assign node13917 = (inp[12]) ? node13921 : node13918;
													assign node13918 = (inp[9]) ? 15'b000000001111111 : 15'b000000001111111;
													assign node13921 = (inp[9]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node13924 = (inp[14]) ? node13928 : node13925;
													assign node13925 = (inp[9]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node13928 = (inp[13]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node13931 = (inp[9]) ? node13947 : node13932;
											assign node13932 = (inp[13]) ? node13940 : node13933;
												assign node13933 = (inp[1]) ? node13937 : node13934;
													assign node13934 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node13937 = (inp[12]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node13940 = (inp[14]) ? node13944 : node13941;
													assign node13941 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node13944 = (inp[5]) ? 15'b000000000011111 : 15'b000000000011111;
											assign node13947 = (inp[1]) ? node13955 : node13948;
												assign node13948 = (inp[14]) ? node13952 : node13949;
													assign node13949 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node13952 = (inp[5]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node13955 = (inp[5]) ? node13959 : node13956;
													assign node13956 = (inp[13]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node13959 = (inp[12]) ? 15'b000000000001111 : 15'b000000000011111;
								assign node13962 = (inp[1]) ? node14024 : node13963;
									assign node13963 = (inp[13]) ? node13993 : node13964;
										assign node13964 = (inp[5]) ? node13980 : node13965;
											assign node13965 = (inp[2]) ? node13973 : node13966;
												assign node13966 = (inp[10]) ? node13970 : node13967;
													assign node13967 = (inp[9]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node13970 = (inp[9]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node13973 = (inp[12]) ? node13977 : node13974;
													assign node13974 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node13977 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node13980 = (inp[12]) ? node13986 : node13981;
												assign node13981 = (inp[10]) ? node13983 : 15'b000000011111111;
													assign node13983 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node13986 = (inp[9]) ? node13990 : node13987;
													assign node13987 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node13990 = (inp[10]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node13993 = (inp[2]) ? node14009 : node13994;
											assign node13994 = (inp[5]) ? node14002 : node13995;
												assign node13995 = (inp[10]) ? node13999 : node13996;
													assign node13996 = (inp[9]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node13999 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node14002 = (inp[9]) ? node14006 : node14003;
													assign node14003 = (inp[12]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node14006 = (inp[10]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node14009 = (inp[12]) ? node14017 : node14010;
												assign node14010 = (inp[5]) ? node14014 : node14011;
													assign node14011 = (inp[9]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node14014 = (inp[9]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node14017 = (inp[10]) ? node14021 : node14018;
													assign node14018 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node14021 = (inp[9]) ? 15'b000000000000111 : 15'b000000000001111;
									assign node14024 = (inp[9]) ? node14054 : node14025;
										assign node14025 = (inp[2]) ? node14039 : node14026;
											assign node14026 = (inp[5]) ? node14034 : node14027;
												assign node14027 = (inp[13]) ? node14031 : node14028;
													assign node14028 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node14031 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node14034 = (inp[12]) ? 15'b000000000011111 : node14035;
													assign node14035 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node14039 = (inp[12]) ? node14047 : node14040;
												assign node14040 = (inp[10]) ? node14044 : node14041;
													assign node14041 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node14044 = (inp[5]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node14047 = (inp[13]) ? node14051 : node14048;
													assign node14048 = (inp[5]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node14051 = (inp[5]) ? 15'b000000000001111 : 15'b000000000011111;
										assign node14054 = (inp[14]) ? node14070 : node14055;
											assign node14055 = (inp[10]) ? node14063 : node14056;
												assign node14056 = (inp[5]) ? node14060 : node14057;
													assign node14057 = (inp[12]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node14060 = (inp[2]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node14063 = (inp[12]) ? node14067 : node14064;
													assign node14064 = (inp[2]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node14067 = (inp[2]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node14070 = (inp[13]) ? node14078 : node14071;
												assign node14071 = (inp[10]) ? node14075 : node14072;
													assign node14072 = (inp[12]) ? 15'b000000000001111 : 15'b000000000111111;
													assign node14075 = (inp[5]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node14078 = (inp[5]) ? node14082 : node14079;
													assign node14079 = (inp[2]) ? 15'b000000000001111 : 15'b000000000001111;
													assign node14082 = (inp[12]) ? 15'b000000000000111 : 15'b000000000001111;
						assign node14085 = (inp[1]) ? node14331 : node14086;
							assign node14086 = (inp[4]) ? node14210 : node14087;
								assign node14087 = (inp[12]) ? node14147 : node14088;
									assign node14088 = (inp[10]) ? node14118 : node14089;
										assign node14089 = (inp[7]) ? node14103 : node14090;
											assign node14090 = (inp[5]) ? node14098 : node14091;
												assign node14091 = (inp[14]) ? node14095 : node14092;
													assign node14092 = (inp[9]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node14095 = (inp[9]) ? 15'b000000111111111 : 15'b000000011111111;
												assign node14098 = (inp[14]) ? 15'b000000011111111 : node14099;
													assign node14099 = (inp[9]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node14103 = (inp[14]) ? node14111 : node14104;
												assign node14104 = (inp[5]) ? node14108 : node14105;
													assign node14105 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node14108 = (inp[9]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node14111 = (inp[5]) ? node14115 : node14112;
													assign node14112 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node14115 = (inp[9]) ? 15'b000000000111111 : 15'b000000011111111;
										assign node14118 = (inp[9]) ? node14134 : node14119;
											assign node14119 = (inp[7]) ? node14127 : node14120;
												assign node14120 = (inp[5]) ? node14124 : node14121;
													assign node14121 = (inp[13]) ? 15'b000000001111111 : 15'b000000111111111;
													assign node14124 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node14127 = (inp[14]) ? node14131 : node14128;
													assign node14128 = (inp[5]) ? 15'b000000000111111 : 15'b000000011111111;
													assign node14131 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node14134 = (inp[7]) ? node14140 : node14135;
												assign node14135 = (inp[5]) ? node14137 : 15'b000000001111111;
													assign node14137 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node14140 = (inp[5]) ? node14144 : node14141;
													assign node14141 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node14144 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node14147 = (inp[2]) ? node14179 : node14148;
										assign node14148 = (inp[13]) ? node14164 : node14149;
											assign node14149 = (inp[5]) ? node14157 : node14150;
												assign node14150 = (inp[14]) ? node14154 : node14151;
													assign node14151 = (inp[9]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node14154 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node14157 = (inp[10]) ? node14161 : node14158;
													assign node14158 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node14161 = (inp[9]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node14164 = (inp[10]) ? node14172 : node14165;
												assign node14165 = (inp[9]) ? node14169 : node14166;
													assign node14166 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node14169 = (inp[7]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node14172 = (inp[7]) ? node14176 : node14173;
													assign node14173 = (inp[9]) ? 15'b000000000011111 : 15'b000000001111111;
													assign node14176 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node14179 = (inp[7]) ? node14195 : node14180;
											assign node14180 = (inp[5]) ? node14188 : node14181;
												assign node14181 = (inp[13]) ? node14185 : node14182;
													assign node14182 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node14185 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node14188 = (inp[14]) ? node14192 : node14189;
													assign node14189 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node14192 = (inp[9]) ? 15'b000000000011111 : 15'b000000000011111;
											assign node14195 = (inp[10]) ? node14203 : node14196;
												assign node14196 = (inp[13]) ? node14200 : node14197;
													assign node14197 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node14200 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node14203 = (inp[9]) ? node14207 : node14204;
													assign node14204 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node14207 = (inp[14]) ? 15'b000000000001111 : 15'b000000000001111;
								assign node14210 = (inp[9]) ? node14270 : node14211;
									assign node14211 = (inp[13]) ? node14239 : node14212;
										assign node14212 = (inp[14]) ? node14228 : node14213;
											assign node14213 = (inp[10]) ? node14221 : node14214;
												assign node14214 = (inp[12]) ? node14218 : node14215;
													assign node14215 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node14218 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node14221 = (inp[7]) ? node14225 : node14222;
													assign node14222 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node14225 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node14228 = (inp[5]) ? node14234 : node14229;
												assign node14229 = (inp[12]) ? node14231 : 15'b000000111111111;
													assign node14231 = (inp[7]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node14234 = (inp[7]) ? 15'b000000000011111 : node14235;
													assign node14235 = (inp[12]) ? 15'b000000000111111 : 15'b000000000111111;
										assign node14239 = (inp[5]) ? node14255 : node14240;
											assign node14240 = (inp[12]) ? node14248 : node14241;
												assign node14241 = (inp[14]) ? node14245 : node14242;
													assign node14242 = (inp[2]) ? 15'b000000011111111 : 15'b000000011111111;
													assign node14245 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node14248 = (inp[14]) ? node14252 : node14249;
													assign node14249 = (inp[7]) ? 15'b000000000111111 : 15'b000000000111111;
													assign node14252 = (inp[7]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node14255 = (inp[7]) ? node14263 : node14256;
												assign node14256 = (inp[12]) ? node14260 : node14257;
													assign node14257 = (inp[10]) ? 15'b000000000111111 : 15'b000000000111111;
													assign node14260 = (inp[2]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node14263 = (inp[14]) ? node14267 : node14264;
													assign node14264 = (inp[2]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node14267 = (inp[12]) ? 15'b000000000001111 : 15'b000000000011111;
									assign node14270 = (inp[2]) ? node14300 : node14271;
										assign node14271 = (inp[13]) ? node14285 : node14272;
											assign node14272 = (inp[5]) ? node14280 : node14273;
												assign node14273 = (inp[10]) ? node14277 : node14274;
													assign node14274 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node14277 = (inp[12]) ? 15'b000000000011111 : 15'b000000001111111;
												assign node14280 = (inp[14]) ? 15'b000000000111111 : node14281;
													assign node14281 = (inp[7]) ? 15'b000000000111111 : 15'b000000000111111;
											assign node14285 = (inp[12]) ? node14293 : node14286;
												assign node14286 = (inp[7]) ? node14290 : node14287;
													assign node14287 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node14290 = (inp[5]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node14293 = (inp[14]) ? node14297 : node14294;
													assign node14294 = (inp[7]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node14297 = (inp[10]) ? 15'b000000000001111 : 15'b000000000011111;
										assign node14300 = (inp[14]) ? node14316 : node14301;
											assign node14301 = (inp[10]) ? node14309 : node14302;
												assign node14302 = (inp[13]) ? node14306 : node14303;
													assign node14303 = (inp[12]) ? 15'b000000000111111 : 15'b000000000111111;
													assign node14306 = (inp[5]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node14309 = (inp[13]) ? node14313 : node14310;
													assign node14310 = (inp[7]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node14313 = (inp[7]) ? 15'b000000000001111 : 15'b000000000001111;
											assign node14316 = (inp[10]) ? node14324 : node14317;
												assign node14317 = (inp[13]) ? node14321 : node14318;
													assign node14318 = (inp[5]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node14321 = (inp[5]) ? 15'b000000000000111 : 15'b000000000001111;
												assign node14324 = (inp[12]) ? node14328 : node14325;
													assign node14325 = (inp[5]) ? 15'b000000000001111 : 15'b000000000011111;
													assign node14328 = (inp[13]) ? 15'b000000000000111 : 15'b000000000000111;
							assign node14331 = (inp[13]) ? node14451 : node14332;
								assign node14332 = (inp[10]) ? node14394 : node14333;
									assign node14333 = (inp[5]) ? node14365 : node14334;
										assign node14334 = (inp[14]) ? node14350 : node14335;
											assign node14335 = (inp[9]) ? node14343 : node14336;
												assign node14336 = (inp[7]) ? node14340 : node14337;
													assign node14337 = (inp[12]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node14340 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node14343 = (inp[7]) ? node14347 : node14344;
													assign node14344 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node14347 = (inp[12]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node14350 = (inp[9]) ? node14358 : node14351;
												assign node14351 = (inp[4]) ? node14355 : node14352;
													assign node14352 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node14355 = (inp[7]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node14358 = (inp[4]) ? node14362 : node14359;
													assign node14359 = (inp[7]) ? 15'b000000000011111 : 15'b000000001111111;
													assign node14362 = (inp[2]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node14365 = (inp[7]) ? node14379 : node14366;
											assign node14366 = (inp[4]) ? node14374 : node14367;
												assign node14367 = (inp[9]) ? node14371 : node14368;
													assign node14368 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node14371 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node14374 = (inp[2]) ? 15'b000000000011111 : node14375;
													assign node14375 = (inp[9]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node14379 = (inp[2]) ? node14387 : node14380;
												assign node14380 = (inp[9]) ? node14384 : node14381;
													assign node14381 = (inp[12]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node14384 = (inp[4]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node14387 = (inp[14]) ? node14391 : node14388;
													assign node14388 = (inp[12]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node14391 = (inp[9]) ? 15'b000000000000111 : 15'b000000000011111;
									assign node14394 = (inp[2]) ? node14424 : node14395;
										assign node14395 = (inp[4]) ? node14411 : node14396;
											assign node14396 = (inp[12]) ? node14404 : node14397;
												assign node14397 = (inp[5]) ? node14401 : node14398;
													assign node14398 = (inp[9]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node14401 = (inp[7]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node14404 = (inp[14]) ? node14408 : node14405;
													assign node14405 = (inp[9]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node14408 = (inp[5]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node14411 = (inp[7]) ? node14417 : node14412;
												assign node14412 = (inp[12]) ? node14414 : 15'b000000000111111;
													assign node14414 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node14417 = (inp[14]) ? node14421 : node14418;
													assign node14418 = (inp[5]) ? 15'b000000000011111 : 15'b000000000011111;
													assign node14421 = (inp[12]) ? 15'b000000000000111 : 15'b000000000011111;
										assign node14424 = (inp[9]) ? node14440 : node14425;
											assign node14425 = (inp[12]) ? node14433 : node14426;
												assign node14426 = (inp[14]) ? node14430 : node14427;
													assign node14427 = (inp[7]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node14430 = (inp[7]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node14433 = (inp[4]) ? node14437 : node14434;
													assign node14434 = (inp[5]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node14437 = (inp[5]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node14440 = (inp[7]) ? node14444 : node14441;
												assign node14441 = (inp[12]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node14444 = (inp[14]) ? node14448 : node14445;
													assign node14445 = (inp[4]) ? 15'b000000000001111 : 15'b000000000011111;
													assign node14448 = (inp[12]) ? 15'b000000000000111 : 15'b000000000000111;
								assign node14451 = (inp[14]) ? node14511 : node14452;
									assign node14452 = (inp[2]) ? node14482 : node14453;
										assign node14453 = (inp[9]) ? node14467 : node14454;
											assign node14454 = (inp[12]) ? node14460 : node14455;
												assign node14455 = (inp[10]) ? node14457 : 15'b000000001111111;
													assign node14457 = (inp[5]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node14460 = (inp[10]) ? node14464 : node14461;
													assign node14461 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node14464 = (inp[4]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node14467 = (inp[12]) ? node14475 : node14468;
												assign node14468 = (inp[10]) ? node14472 : node14469;
													assign node14469 = (inp[5]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node14472 = (inp[5]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node14475 = (inp[10]) ? node14479 : node14476;
													assign node14476 = (inp[5]) ? 15'b000000000011111 : 15'b000000000011111;
													assign node14479 = (inp[5]) ? 15'b000000000000111 : 15'b000000000011111;
										assign node14482 = (inp[4]) ? node14498 : node14483;
											assign node14483 = (inp[7]) ? node14491 : node14484;
												assign node14484 = (inp[12]) ? node14488 : node14485;
													assign node14485 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node14488 = (inp[10]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node14491 = (inp[5]) ? node14495 : node14492;
													assign node14492 = (inp[10]) ? 15'b000000000001111 : 15'b000000000111111;
													assign node14495 = (inp[12]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node14498 = (inp[12]) ? node14506 : node14499;
												assign node14499 = (inp[9]) ? node14503 : node14500;
													assign node14500 = (inp[5]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node14503 = (inp[7]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node14506 = (inp[9]) ? 15'b000000000001111 : node14507;
													assign node14507 = (inp[7]) ? 15'b000000000001111 : 15'b000000000011111;
									assign node14511 = (inp[9]) ? node14543 : node14512;
										assign node14512 = (inp[4]) ? node14528 : node14513;
											assign node14513 = (inp[7]) ? node14521 : node14514;
												assign node14514 = (inp[5]) ? node14518 : node14515;
													assign node14515 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node14518 = (inp[10]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node14521 = (inp[2]) ? node14525 : node14522;
													assign node14522 = (inp[10]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node14525 = (inp[12]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node14528 = (inp[5]) ? node14536 : node14529;
												assign node14529 = (inp[10]) ? node14533 : node14530;
													assign node14530 = (inp[2]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node14533 = (inp[12]) ? 15'b000000000000111 : 15'b000000000011111;
												assign node14536 = (inp[7]) ? node14540 : node14537;
													assign node14537 = (inp[2]) ? 15'b000000000001111 : 15'b000000000011111;
													assign node14540 = (inp[12]) ? 15'b000000000000111 : 15'b000000000001111;
										assign node14543 = (inp[2]) ? node14559 : node14544;
											assign node14544 = (inp[12]) ? node14552 : node14545;
												assign node14545 = (inp[7]) ? node14549 : node14546;
													assign node14546 = (inp[5]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node14549 = (inp[4]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node14552 = (inp[10]) ? node14556 : node14553;
													assign node14553 = (inp[4]) ? 15'b000000000001111 : 15'b000000000011111;
													assign node14556 = (inp[4]) ? 15'b000000000000111 : 15'b000000000001111;
											assign node14559 = (inp[7]) ? node14567 : node14560;
												assign node14560 = (inp[5]) ? node14564 : node14561;
													assign node14561 = (inp[10]) ? 15'b000000000000111 : 15'b000000000011111;
													assign node14564 = (inp[4]) ? 15'b000000000000111 : 15'b000000000000111;
												assign node14567 = (inp[10]) ? node14571 : node14568;
													assign node14568 = (inp[5]) ? 15'b000000000000111 : 15'b000000000001111;
													assign node14571 = (inp[4]) ? 15'b000000000000011 : 15'b000000000000111;
					assign node14574 = (inp[1]) ? node15072 : node14575;
						assign node14575 = (inp[2]) ? node14825 : node14576;
							assign node14576 = (inp[9]) ? node14700 : node14577;
								assign node14577 = (inp[14]) ? node14639 : node14578;
									assign node14578 = (inp[8]) ? node14608 : node14579;
										assign node14579 = (inp[13]) ? node14595 : node14580;
											assign node14580 = (inp[5]) ? node14588 : node14581;
												assign node14581 = (inp[7]) ? node14585 : node14582;
													assign node14582 = (inp[4]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node14585 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node14588 = (inp[12]) ? node14592 : node14589;
													assign node14589 = (inp[7]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node14592 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node14595 = (inp[12]) ? node14603 : node14596;
												assign node14596 = (inp[5]) ? node14600 : node14597;
													assign node14597 = (inp[7]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node14600 = (inp[7]) ? 15'b000000000111111 : 15'b000000011111111;
												assign node14603 = (inp[7]) ? 15'b000000001111111 : node14604;
													assign node14604 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node14608 = (inp[13]) ? node14624 : node14609;
											assign node14609 = (inp[5]) ? node14617 : node14610;
												assign node14610 = (inp[12]) ? node14614 : node14611;
													assign node14611 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node14614 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node14617 = (inp[12]) ? node14621 : node14618;
													assign node14618 = (inp[7]) ? 15'b000000001111111 : 15'b000000001111111;
													assign node14621 = (inp[7]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node14624 = (inp[4]) ? node14632 : node14625;
												assign node14625 = (inp[5]) ? node14629 : node14626;
													assign node14626 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node14629 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node14632 = (inp[12]) ? node14636 : node14633;
													assign node14633 = (inp[7]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node14636 = (inp[5]) ? 15'b000000000001111 : 15'b000000000011111;
									assign node14639 = (inp[8]) ? node14671 : node14640;
										assign node14640 = (inp[5]) ? node14656 : node14641;
											assign node14641 = (inp[10]) ? node14649 : node14642;
												assign node14642 = (inp[4]) ? node14646 : node14643;
													assign node14643 = (inp[7]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node14646 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node14649 = (inp[13]) ? node14653 : node14650;
													assign node14650 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node14653 = (inp[12]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node14656 = (inp[4]) ? node14664 : node14657;
												assign node14657 = (inp[7]) ? node14661 : node14658;
													assign node14658 = (inp[12]) ? 15'b000000001111111 : 15'b000000111111111;
													assign node14661 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node14664 = (inp[12]) ? node14668 : node14665;
													assign node14665 = (inp[7]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node14668 = (inp[7]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node14671 = (inp[7]) ? node14685 : node14672;
											assign node14672 = (inp[13]) ? node14678 : node14673;
												assign node14673 = (inp[12]) ? node14675 : 15'b000000001111111;
													assign node14675 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node14678 = (inp[10]) ? node14682 : node14679;
													assign node14679 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node14682 = (inp[12]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node14685 = (inp[13]) ? node14693 : node14686;
												assign node14686 = (inp[5]) ? node14690 : node14687;
													assign node14687 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node14690 = (inp[12]) ? 15'b000000000001111 : 15'b000000000111111;
												assign node14693 = (inp[12]) ? node14697 : node14694;
													assign node14694 = (inp[4]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node14697 = (inp[10]) ? 15'b000000000000111 : 15'b000000000011111;
								assign node14700 = (inp[4]) ? node14762 : node14701;
									assign node14701 = (inp[13]) ? node14733 : node14702;
										assign node14702 = (inp[10]) ? node14718 : node14703;
											assign node14703 = (inp[5]) ? node14711 : node14704;
												assign node14704 = (inp[7]) ? node14708 : node14705;
													assign node14705 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node14708 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node14711 = (inp[8]) ? node14715 : node14712;
													assign node14712 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node14715 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node14718 = (inp[5]) ? node14726 : node14719;
												assign node14719 = (inp[12]) ? node14723 : node14720;
													assign node14720 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node14723 = (inp[7]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node14726 = (inp[7]) ? node14730 : node14727;
													assign node14727 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node14730 = (inp[12]) ? 15'b000000000011111 : 15'b000000000011111;
										assign node14733 = (inp[8]) ? node14747 : node14734;
											assign node14734 = (inp[7]) ? node14742 : node14735;
												assign node14735 = (inp[10]) ? node14739 : node14736;
													assign node14736 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node14739 = (inp[5]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node14742 = (inp[10]) ? node14744 : 15'b000000001111111;
													assign node14744 = (inp[5]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node14747 = (inp[10]) ? node14755 : node14748;
												assign node14748 = (inp[5]) ? node14752 : node14749;
													assign node14749 = (inp[12]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node14752 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node14755 = (inp[14]) ? node14759 : node14756;
													assign node14756 = (inp[12]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node14759 = (inp[12]) ? 15'b000000000001111 : 15'b000000000001111;
									assign node14762 = (inp[14]) ? node14794 : node14763;
										assign node14763 = (inp[8]) ? node14779 : node14764;
											assign node14764 = (inp[10]) ? node14772 : node14765;
												assign node14765 = (inp[7]) ? node14769 : node14766;
													assign node14766 = (inp[5]) ? 15'b000000001111111 : 15'b000000001111111;
													assign node14769 = (inp[12]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node14772 = (inp[5]) ? node14776 : node14773;
													assign node14773 = (inp[7]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node14776 = (inp[12]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node14779 = (inp[12]) ? node14787 : node14780;
												assign node14780 = (inp[5]) ? node14784 : node14781;
													assign node14781 = (inp[13]) ? 15'b000000000111111 : 15'b000000000111111;
													assign node14784 = (inp[7]) ? 15'b000000000011111 : 15'b000000000011111;
												assign node14787 = (inp[5]) ? node14791 : node14788;
													assign node14788 = (inp[13]) ? 15'b000000000011111 : 15'b000000000011111;
													assign node14791 = (inp[10]) ? 15'b000000000001111 : 15'b000000000011111;
										assign node14794 = (inp[12]) ? node14810 : node14795;
											assign node14795 = (inp[10]) ? node14803 : node14796;
												assign node14796 = (inp[13]) ? node14800 : node14797;
													assign node14797 = (inp[7]) ? 15'b000000000011111 : 15'b000000001111111;
													assign node14800 = (inp[5]) ? 15'b000000000011111 : 15'b000000000011111;
												assign node14803 = (inp[8]) ? node14807 : node14804;
													assign node14804 = (inp[7]) ? 15'b000000000011111 : 15'b000000000011111;
													assign node14807 = (inp[7]) ? 15'b000000000001111 : 15'b000000000001111;
											assign node14810 = (inp[8]) ? node14818 : node14811;
												assign node14811 = (inp[5]) ? node14815 : node14812;
													assign node14812 = (inp[7]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node14815 = (inp[10]) ? 15'b000000000000111 : 15'b000000000011111;
												assign node14818 = (inp[7]) ? node14822 : node14819;
													assign node14819 = (inp[13]) ? 15'b000000000000111 : 15'b000000000001111;
													assign node14822 = (inp[13]) ? 15'b000000000000011 : 15'b000000000000111;
							assign node14825 = (inp[7]) ? node14951 : node14826;
								assign node14826 = (inp[13]) ? node14888 : node14827;
									assign node14827 = (inp[14]) ? node14859 : node14828;
										assign node14828 = (inp[8]) ? node14844 : node14829;
											assign node14829 = (inp[4]) ? node14837 : node14830;
												assign node14830 = (inp[5]) ? node14834 : node14831;
													assign node14831 = (inp[10]) ? 15'b000000011111111 : 15'b000001111111111;
													assign node14834 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node14837 = (inp[9]) ? node14841 : node14838;
													assign node14838 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node14841 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node14844 = (inp[10]) ? node14852 : node14845;
												assign node14845 = (inp[5]) ? node14849 : node14846;
													assign node14846 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node14849 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node14852 = (inp[4]) ? node14856 : node14853;
													assign node14853 = (inp[9]) ? 15'b000000000111111 : 15'b000000000111111;
													assign node14856 = (inp[12]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node14859 = (inp[8]) ? node14873 : node14860;
											assign node14860 = (inp[5]) ? node14868 : node14861;
												assign node14861 = (inp[9]) ? node14865 : node14862;
													assign node14862 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node14865 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node14868 = (inp[4]) ? node14870 : 15'b000000000111111;
													assign node14870 = (inp[9]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node14873 = (inp[5]) ? node14881 : node14874;
												assign node14874 = (inp[9]) ? node14878 : node14875;
													assign node14875 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node14878 = (inp[12]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node14881 = (inp[9]) ? node14885 : node14882;
													assign node14882 = (inp[12]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node14885 = (inp[12]) ? 15'b000000000000111 : 15'b000000000001111;
									assign node14888 = (inp[12]) ? node14920 : node14889;
										assign node14889 = (inp[14]) ? node14905 : node14890;
											assign node14890 = (inp[10]) ? node14898 : node14891;
												assign node14891 = (inp[9]) ? node14895 : node14892;
													assign node14892 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node14895 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node14898 = (inp[8]) ? node14902 : node14899;
													assign node14899 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node14902 = (inp[9]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node14905 = (inp[10]) ? node14913 : node14906;
												assign node14906 = (inp[4]) ? node14910 : node14907;
													assign node14907 = (inp[9]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node14910 = (inp[8]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node14913 = (inp[9]) ? node14917 : node14914;
													assign node14914 = (inp[4]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node14917 = (inp[5]) ? 15'b000000000001111 : 15'b000000000011111;
										assign node14920 = (inp[4]) ? node14936 : node14921;
											assign node14921 = (inp[8]) ? node14929 : node14922;
												assign node14922 = (inp[5]) ? node14926 : node14923;
													assign node14923 = (inp[14]) ? 15'b000000000111111 : 15'b000000000111111;
													assign node14926 = (inp[10]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node14929 = (inp[14]) ? node14933 : node14930;
													assign node14930 = (inp[9]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node14933 = (inp[10]) ? 15'b000000000000111 : 15'b000000000011111;
											assign node14936 = (inp[5]) ? node14944 : node14937;
												assign node14937 = (inp[10]) ? node14941 : node14938;
													assign node14938 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node14941 = (inp[14]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node14944 = (inp[9]) ? node14948 : node14945;
													assign node14945 = (inp[8]) ? 15'b000000000001111 : 15'b000000000001111;
													assign node14948 = (inp[8]) ? 15'b000000000000011 : 15'b000000000001111;
								assign node14951 = (inp[8]) ? node15009 : node14952;
									assign node14952 = (inp[12]) ? node14978 : node14953;
										assign node14953 = (inp[13]) ? node14969 : node14954;
											assign node14954 = (inp[5]) ? node14962 : node14955;
												assign node14955 = (inp[4]) ? node14959 : node14956;
													assign node14956 = (inp[10]) ? 15'b000000001111111 : 15'b000000001111111;
													assign node14959 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node14962 = (inp[10]) ? node14966 : node14963;
													assign node14963 = (inp[9]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node14966 = (inp[9]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node14969 = (inp[4]) ? node14975 : node14970;
												assign node14970 = (inp[9]) ? 15'b000000000111111 : node14971;
													assign node14971 = (inp[5]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node14975 = (inp[9]) ? 15'b000000000001111 : 15'b000000000011111;
										assign node14978 = (inp[5]) ? node14994 : node14979;
											assign node14979 = (inp[9]) ? node14987 : node14980;
												assign node14980 = (inp[4]) ? node14984 : node14981;
													assign node14981 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node14984 = (inp[10]) ? 15'b000000000011111 : 15'b000000000011111;
												assign node14987 = (inp[4]) ? node14991 : node14988;
													assign node14988 = (inp[13]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node14991 = (inp[10]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node14994 = (inp[14]) ? node15002 : node14995;
												assign node14995 = (inp[9]) ? node14999 : node14996;
													assign node14996 = (inp[13]) ? 15'b000000000001111 : 15'b000000000111111;
													assign node14999 = (inp[10]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node15002 = (inp[10]) ? node15006 : node15003;
													assign node15003 = (inp[9]) ? 15'b000000000001111 : 15'b000000000001111;
													assign node15006 = (inp[9]) ? 15'b000000000000011 : 15'b000000000001111;
									assign node15009 = (inp[4]) ? node15041 : node15010;
										assign node15010 = (inp[5]) ? node15026 : node15011;
											assign node15011 = (inp[10]) ? node15019 : node15012;
												assign node15012 = (inp[12]) ? node15016 : node15013;
													assign node15013 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node15016 = (inp[13]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node15019 = (inp[9]) ? node15023 : node15020;
													assign node15020 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node15023 = (inp[14]) ? 15'b000000000000111 : 15'b000000000011111;
											assign node15026 = (inp[12]) ? node15034 : node15027;
												assign node15027 = (inp[10]) ? node15031 : node15028;
													assign node15028 = (inp[13]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node15031 = (inp[13]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node15034 = (inp[13]) ? node15038 : node15035;
													assign node15035 = (inp[9]) ? 15'b000000000001111 : 15'b000000000011111;
													assign node15038 = (inp[14]) ? 15'b000000000000111 : 15'b000000000001111;
										assign node15041 = (inp[14]) ? node15057 : node15042;
											assign node15042 = (inp[10]) ? node15050 : node15043;
												assign node15043 = (inp[13]) ? node15047 : node15044;
													assign node15044 = (inp[9]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node15047 = (inp[9]) ? 15'b000000000001111 : 15'b000000000001111;
												assign node15050 = (inp[9]) ? node15054 : node15051;
													assign node15051 = (inp[12]) ? 15'b000000000001111 : 15'b000000000011111;
													assign node15054 = (inp[13]) ? 15'b000000000000111 : 15'b000000000001111;
											assign node15057 = (inp[12]) ? node15065 : node15058;
												assign node15058 = (inp[5]) ? node15062 : node15059;
													assign node15059 = (inp[10]) ? 15'b000000000001111 : 15'b000000000011111;
													assign node15062 = (inp[13]) ? 15'b000000000000111 : 15'b000000000001111;
												assign node15065 = (inp[9]) ? node15069 : node15066;
													assign node15066 = (inp[10]) ? 15'b000000000000111 : 15'b000000000001111;
													assign node15069 = (inp[5]) ? 15'b000000000000001 : 15'b000000000000111;
						assign node15072 = (inp[12]) ? node15308 : node15073;
							assign node15073 = (inp[4]) ? node15193 : node15074;
								assign node15074 = (inp[13]) ? node15136 : node15075;
									assign node15075 = (inp[14]) ? node15107 : node15076;
										assign node15076 = (inp[2]) ? node15092 : node15077;
											assign node15077 = (inp[7]) ? node15085 : node15078;
												assign node15078 = (inp[9]) ? node15082 : node15079;
													assign node15079 = (inp[8]) ? 15'b000000011111111 : 15'b000001111111111;
													assign node15082 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node15085 = (inp[5]) ? node15089 : node15086;
													assign node15086 = (inp[9]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node15089 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node15092 = (inp[10]) ? node15100 : node15093;
												assign node15093 = (inp[9]) ? node15097 : node15094;
													assign node15094 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node15097 = (inp[7]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node15100 = (inp[8]) ? node15104 : node15101;
													assign node15101 = (inp[9]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node15104 = (inp[5]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node15107 = (inp[10]) ? node15121 : node15108;
											assign node15108 = (inp[9]) ? node15116 : node15109;
												assign node15109 = (inp[2]) ? node15113 : node15110;
													assign node15110 = (inp[5]) ? 15'b000000001111111 : 15'b000000111111111;
													assign node15113 = (inp[7]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node15116 = (inp[7]) ? 15'b000000000011111 : node15117;
													assign node15117 = (inp[5]) ? 15'b000000000111111 : 15'b000000000111111;
											assign node15121 = (inp[5]) ? node15129 : node15122;
												assign node15122 = (inp[2]) ? node15126 : node15123;
													assign node15123 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node15126 = (inp[8]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node15129 = (inp[7]) ? node15133 : node15130;
													assign node15130 = (inp[2]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node15133 = (inp[8]) ? 15'b000000000001111 : 15'b000000000111111;
									assign node15136 = (inp[8]) ? node15162 : node15137;
										assign node15137 = (inp[5]) ? node15151 : node15138;
											assign node15138 = (inp[14]) ? node15144 : node15139;
												assign node15139 = (inp[7]) ? 15'b000000001111111 : node15140;
													assign node15140 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node15144 = (inp[7]) ? node15148 : node15145;
													assign node15145 = (inp[9]) ? 15'b000000000111111 : 15'b000000011111111;
													assign node15148 = (inp[9]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node15151 = (inp[7]) ? node15157 : node15152;
												assign node15152 = (inp[10]) ? 15'b000000000011111 : node15153;
													assign node15153 = (inp[9]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node15157 = (inp[2]) ? 15'b000000000011111 : node15158;
													assign node15158 = (inp[9]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node15162 = (inp[5]) ? node15178 : node15163;
											assign node15163 = (inp[14]) ? node15171 : node15164;
												assign node15164 = (inp[7]) ? node15168 : node15165;
													assign node15165 = (inp[10]) ? 15'b000000000111111 : 15'b000000000111111;
													assign node15168 = (inp[9]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node15171 = (inp[10]) ? node15175 : node15172;
													assign node15172 = (inp[7]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node15175 = (inp[7]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node15178 = (inp[10]) ? node15186 : node15179;
												assign node15179 = (inp[9]) ? node15183 : node15180;
													assign node15180 = (inp[2]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node15183 = (inp[14]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node15186 = (inp[7]) ? node15190 : node15187;
													assign node15187 = (inp[2]) ? 15'b000000000001111 : 15'b000000000011111;
													assign node15190 = (inp[2]) ? 15'b000000000000111 : 15'b000000000001111;
								assign node15193 = (inp[10]) ? node15251 : node15194;
									assign node15194 = (inp[5]) ? node15222 : node15195;
										assign node15195 = (inp[13]) ? node15207 : node15196;
											assign node15196 = (inp[2]) ? node15202 : node15197;
												assign node15197 = (inp[7]) ? 15'b000000001111111 : node15198;
													assign node15198 = (inp[14]) ? 15'b000000001111111 : 15'b000000111111111;
												assign node15202 = (inp[8]) ? 15'b000000000111111 : node15203;
													assign node15203 = (inp[7]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node15207 = (inp[8]) ? node15215 : node15208;
												assign node15208 = (inp[14]) ? node15212 : node15209;
													assign node15209 = (inp[7]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node15212 = (inp[2]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node15215 = (inp[2]) ? node15219 : node15216;
													assign node15216 = (inp[7]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node15219 = (inp[9]) ? 15'b000000000001111 : 15'b000000000011111;
										assign node15222 = (inp[2]) ? node15236 : node15223;
											assign node15223 = (inp[7]) ? node15229 : node15224;
												assign node15224 = (inp[8]) ? 15'b000000000011111 : node15225;
													assign node15225 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node15229 = (inp[9]) ? node15233 : node15230;
													assign node15230 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node15233 = (inp[8]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node15236 = (inp[7]) ? node15244 : node15237;
												assign node15237 = (inp[8]) ? node15241 : node15238;
													assign node15238 = (inp[9]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node15241 = (inp[9]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node15244 = (inp[13]) ? node15248 : node15245;
													assign node15245 = (inp[8]) ? 15'b000000000001111 : 15'b000000000011111;
													assign node15248 = (inp[9]) ? 15'b000000000000111 : 15'b000000000001111;
									assign node15251 = (inp[9]) ? node15281 : node15252;
										assign node15252 = (inp[13]) ? node15268 : node15253;
											assign node15253 = (inp[14]) ? node15261 : node15254;
												assign node15254 = (inp[8]) ? node15258 : node15255;
													assign node15255 = (inp[5]) ? 15'b000000001111111 : 15'b000000000111111;
													assign node15258 = (inp[7]) ? 15'b000000000011111 : 15'b000000000011111;
												assign node15261 = (inp[7]) ? node15265 : node15262;
													assign node15262 = (inp[5]) ? 15'b000000000001111 : 15'b000000000111111;
													assign node15265 = (inp[2]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node15268 = (inp[2]) ? node15274 : node15269;
												assign node15269 = (inp[8]) ? node15271 : 15'b000000000011111;
													assign node15271 = (inp[14]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node15274 = (inp[14]) ? node15278 : node15275;
													assign node15275 = (inp[5]) ? 15'b000000000011111 : 15'b000000000001111;
													assign node15278 = (inp[5]) ? 15'b000000000000011 : 15'b000000000000111;
										assign node15281 = (inp[2]) ? node15297 : node15282;
											assign node15282 = (inp[8]) ? node15290 : node15283;
												assign node15283 = (inp[13]) ? node15287 : node15284;
													assign node15284 = (inp[5]) ? 15'b000000000011111 : 15'b000000000011111;
													assign node15287 = (inp[14]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node15290 = (inp[13]) ? node15294 : node15291;
													assign node15291 = (inp[5]) ? 15'b000000000001111 : 15'b000000000011111;
													assign node15294 = (inp[5]) ? 15'b000000000000111 : 15'b000000000001111;
											assign node15297 = (inp[5]) ? node15301 : node15298;
												assign node15298 = (inp[7]) ? 15'b000000000000011 : 15'b000000000001111;
												assign node15301 = (inp[8]) ? node15305 : node15302;
													assign node15302 = (inp[13]) ? 15'b000000000000111 : 15'b000000000000111;
													assign node15305 = (inp[14]) ? 15'b000000000000001 : 15'b000000000000111;
							assign node15308 = (inp[7]) ? node15432 : node15309;
								assign node15309 = (inp[14]) ? node15373 : node15310;
									assign node15310 = (inp[10]) ? node15342 : node15311;
										assign node15311 = (inp[2]) ? node15327 : node15312;
											assign node15312 = (inp[13]) ? node15320 : node15313;
												assign node15313 = (inp[4]) ? node15317 : node15314;
													assign node15314 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node15317 = (inp[9]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node15320 = (inp[4]) ? node15324 : node15321;
													assign node15321 = (inp[5]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node15324 = (inp[8]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node15327 = (inp[9]) ? node15335 : node15328;
												assign node15328 = (inp[5]) ? node15332 : node15329;
													assign node15329 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node15332 = (inp[8]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node15335 = (inp[13]) ? node15339 : node15336;
													assign node15336 = (inp[8]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node15339 = (inp[4]) ? 15'b000000000001111 : 15'b000000000001111;
										assign node15342 = (inp[9]) ? node15358 : node15343;
											assign node15343 = (inp[4]) ? node15351 : node15344;
												assign node15344 = (inp[13]) ? node15348 : node15345;
													assign node15345 = (inp[8]) ? 15'b000000000111111 : 15'b000000000111111;
													assign node15348 = (inp[5]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node15351 = (inp[2]) ? node15355 : node15352;
													assign node15352 = (inp[5]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node15355 = (inp[13]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node15358 = (inp[2]) ? node15366 : node15359;
												assign node15359 = (inp[4]) ? node15363 : node15360;
													assign node15360 = (inp[5]) ? 15'b000000000011111 : 15'b000000000011111;
													assign node15363 = (inp[13]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node15366 = (inp[8]) ? node15370 : node15367;
													assign node15367 = (inp[4]) ? 15'b000000000001111 : 15'b000000000011111;
													assign node15370 = (inp[5]) ? 15'b000000000000111 : 15'b000000000001111;
									assign node15373 = (inp[5]) ? node15401 : node15374;
										assign node15374 = (inp[2]) ? node15388 : node15375;
											assign node15375 = (inp[4]) ? node15381 : node15376;
												assign node15376 = (inp[13]) ? node15378 : 15'b000000000111111;
													assign node15378 = (inp[10]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node15381 = (inp[9]) ? node15385 : node15382;
													assign node15382 = (inp[8]) ? 15'b000000000011111 : 15'b000000000011111;
													assign node15385 = (inp[10]) ? 15'b000000000000111 : 15'b000000000011111;
											assign node15388 = (inp[13]) ? node15394 : node15389;
												assign node15389 = (inp[8]) ? node15391 : 15'b000000000111111;
													assign node15391 = (inp[10]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node15394 = (inp[8]) ? node15398 : node15395;
													assign node15395 = (inp[4]) ? 15'b000000000001111 : 15'b000000000011111;
													assign node15398 = (inp[4]) ? 15'b000000000000111 : 15'b000000000001111;
										assign node15401 = (inp[2]) ? node15417 : node15402;
											assign node15402 = (inp[10]) ? node15410 : node15403;
												assign node15403 = (inp[9]) ? node15407 : node15404;
													assign node15404 = (inp[13]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node15407 = (inp[4]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node15410 = (inp[13]) ? node15414 : node15411;
													assign node15411 = (inp[8]) ? 15'b000000000001111 : 15'b000000000011111;
													assign node15414 = (inp[9]) ? 15'b000000000000111 : 15'b000000000001111;
											assign node15417 = (inp[4]) ? node15425 : node15418;
												assign node15418 = (inp[9]) ? node15422 : node15419;
													assign node15419 = (inp[8]) ? 15'b000000000001111 : 15'b000000000011111;
													assign node15422 = (inp[13]) ? 15'b000000000000111 : 15'b000000000001111;
												assign node15425 = (inp[10]) ? node15429 : node15426;
													assign node15426 = (inp[9]) ? 15'b000000000000111 : 15'b000000000001111;
													assign node15429 = (inp[13]) ? 15'b000000000000011 : 15'b000000000000111;
								assign node15432 = (inp[13]) ? node15496 : node15433;
									assign node15433 = (inp[14]) ? node15465 : node15434;
										assign node15434 = (inp[8]) ? node15450 : node15435;
											assign node15435 = (inp[4]) ? node15443 : node15436;
												assign node15436 = (inp[10]) ? node15440 : node15437;
													assign node15437 = (inp[5]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node15440 = (inp[5]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node15443 = (inp[5]) ? node15447 : node15444;
													assign node15444 = (inp[9]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node15447 = (inp[10]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node15450 = (inp[9]) ? node15458 : node15451;
												assign node15451 = (inp[5]) ? node15455 : node15452;
													assign node15452 = (inp[4]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node15455 = (inp[4]) ? 15'b000000000000111 : 15'b000000000011111;
												assign node15458 = (inp[2]) ? node15462 : node15459;
													assign node15459 = (inp[4]) ? 15'b000000000001111 : 15'b000000000011111;
													assign node15462 = (inp[10]) ? 15'b000000000000111 : 15'b000000000001111;
										assign node15465 = (inp[4]) ? node15481 : node15466;
											assign node15466 = (inp[2]) ? node15474 : node15467;
												assign node15467 = (inp[5]) ? node15471 : node15468;
													assign node15468 = (inp[10]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node15471 = (inp[8]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node15474 = (inp[9]) ? node15478 : node15475;
													assign node15475 = (inp[8]) ? 15'b000000000001111 : 15'b000000000011111;
													assign node15478 = (inp[5]) ? 15'b000000000000111 : 15'b000000000001111;
											assign node15481 = (inp[5]) ? node15489 : node15482;
												assign node15482 = (inp[9]) ? node15486 : node15483;
													assign node15483 = (inp[8]) ? 15'b000000000001111 : 15'b000000000011111;
													assign node15486 = (inp[10]) ? 15'b000000000000111 : 15'b000000000001111;
												assign node15489 = (inp[2]) ? node15493 : node15490;
													assign node15490 = (inp[8]) ? 15'b000000000000111 : 15'b000000000001111;
													assign node15493 = (inp[9]) ? 15'b000000000000011 : 15'b000000000000111;
									assign node15496 = (inp[5]) ? node15528 : node15497;
										assign node15497 = (inp[2]) ? node15513 : node15498;
											assign node15498 = (inp[9]) ? node15506 : node15499;
												assign node15499 = (inp[10]) ? node15503 : node15500;
													assign node15500 = (inp[4]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node15503 = (inp[8]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node15506 = (inp[4]) ? node15510 : node15507;
													assign node15507 = (inp[14]) ? 15'b000000000000111 : 15'b000000000011111;
													assign node15510 = (inp[8]) ? 15'b000000000000111 : 15'b000000000000111;
											assign node15513 = (inp[10]) ? node15521 : node15514;
												assign node15514 = (inp[14]) ? node15518 : node15515;
													assign node15515 = (inp[9]) ? 15'b000000000001111 : 15'b000000000001111;
													assign node15518 = (inp[9]) ? 15'b000000000000111 : 15'b000000000001111;
												assign node15521 = (inp[4]) ? node15525 : node15522;
													assign node15522 = (inp[8]) ? 15'b000000000000111 : 15'b000000000001111;
													assign node15525 = (inp[14]) ? 15'b000000000000011 : 15'b000000000000111;
										assign node15528 = (inp[8]) ? node15542 : node15529;
											assign node15529 = (inp[2]) ? node15535 : node15530;
												assign node15530 = (inp[10]) ? node15532 : 15'b000000000001111;
													assign node15532 = (inp[4]) ? 15'b000000000000111 : 15'b000000000001111;
												assign node15535 = (inp[4]) ? node15539 : node15536;
													assign node15536 = (inp[10]) ? 15'b000000000000111 : 15'b000000000001111;
													assign node15539 = (inp[9]) ? 15'b000000000000001 : 15'b000000000000111;
											assign node15542 = (inp[14]) ? node15550 : node15543;
												assign node15543 = (inp[9]) ? node15547 : node15544;
													assign node15544 = (inp[4]) ? 15'b000000000000111 : 15'b000000000001111;
													assign node15547 = (inp[10]) ? 15'b000000000000011 : 15'b000000000000011;
												assign node15550 = (inp[10]) ? node15552 : 15'b000000000000011;
													assign node15552 = (inp[4]) ? 15'b000000000000001 : 15'b000000000000011;

endmodule