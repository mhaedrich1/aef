module dtc_split75_bm56 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node7;
	wire [3-1:0] node8;
	wire [3-1:0] node9;
	wire [3-1:0] node12;
	wire [3-1:0] node15;
	wire [3-1:0] node16;
	wire [3-1:0] node17;
	wire [3-1:0] node19;
	wire [3-1:0] node23;
	wire [3-1:0] node25;
	wire [3-1:0] node28;
	wire [3-1:0] node29;
	wire [3-1:0] node30;
	wire [3-1:0] node32;
	wire [3-1:0] node33;
	wire [3-1:0] node36;
	wire [3-1:0] node39;
	wire [3-1:0] node40;
	wire [3-1:0] node41;
	wire [3-1:0] node44;
	wire [3-1:0] node47;
	wire [3-1:0] node48;
	wire [3-1:0] node52;
	wire [3-1:0] node53;
	wire [3-1:0] node54;
	wire [3-1:0] node55;
	wire [3-1:0] node59;
	wire [3-1:0] node60;
	wire [3-1:0] node64;
	wire [3-1:0] node65;
	wire [3-1:0] node67;
	wire [3-1:0] node71;
	wire [3-1:0] node72;
	wire [3-1:0] node73;
	wire [3-1:0] node74;
	wire [3-1:0] node75;
	wire [3-1:0] node78;
	wire [3-1:0] node81;
	wire [3-1:0] node82;
	wire [3-1:0] node85;
	wire [3-1:0] node88;
	wire [3-1:0] node89;
	wire [3-1:0] node90;
	wire [3-1:0] node93;
	wire [3-1:0] node96;
	wire [3-1:0] node98;
	wire [3-1:0] node99;
	wire [3-1:0] node102;
	wire [3-1:0] node105;
	wire [3-1:0] node106;
	wire [3-1:0] node107;
	wire [3-1:0] node108;
	wire [3-1:0] node112;
	wire [3-1:0] node113;
	wire [3-1:0] node117;
	wire [3-1:0] node118;
	wire [3-1:0] node120;
	wire [3-1:0] node122;
	wire [3-1:0] node125;
	wire [3-1:0] node126;
	wire [3-1:0] node127;
	wire [3-1:0] node130;
	wire [3-1:0] node133;
	wire [3-1:0] node134;
	wire [3-1:0] node138;
	wire [3-1:0] node139;
	wire [3-1:0] node140;
	wire [3-1:0] node141;
	wire [3-1:0] node142;
	wire [3-1:0] node143;
	wire [3-1:0] node144;
	wire [3-1:0] node147;
	wire [3-1:0] node151;
	wire [3-1:0] node152;
	wire [3-1:0] node153;
	wire [3-1:0] node156;
	wire [3-1:0] node159;
	wire [3-1:0] node160;
	wire [3-1:0] node163;
	wire [3-1:0] node166;
	wire [3-1:0] node167;
	wire [3-1:0] node168;
	wire [3-1:0] node170;
	wire [3-1:0] node174;
	wire [3-1:0] node175;
	wire [3-1:0] node176;
	wire [3-1:0] node181;
	wire [3-1:0] node182;
	wire [3-1:0] node184;
	wire [3-1:0] node186;
	wire [3-1:0] node188;
	wire [3-1:0] node191;
	wire [3-1:0] node192;
	wire [3-1:0] node193;
	wire [3-1:0] node195;
	wire [3-1:0] node199;
	wire [3-1:0] node200;
	wire [3-1:0] node203;
	wire [3-1:0] node206;
	wire [3-1:0] node207;
	wire [3-1:0] node208;
	wire [3-1:0] node209;
	wire [3-1:0] node210;
	wire [3-1:0] node212;
	wire [3-1:0] node215;
	wire [3-1:0] node216;
	wire [3-1:0] node219;
	wire [3-1:0] node222;
	wire [3-1:0] node224;
	wire [3-1:0] node225;
	wire [3-1:0] node229;
	wire [3-1:0] node230;
	wire [3-1:0] node231;
	wire [3-1:0] node232;
	wire [3-1:0] node237;
	wire [3-1:0] node238;
	wire [3-1:0] node242;
	wire [3-1:0] node243;
	wire [3-1:0] node244;
	wire [3-1:0] node245;
	wire [3-1:0] node247;
	wire [3-1:0] node250;
	wire [3-1:0] node251;
	wire [3-1:0] node255;
	wire [3-1:0] node256;
	wire [3-1:0] node259;
	wire [3-1:0] node262;
	wire [3-1:0] node263;
	wire [3-1:0] node265;
	wire [3-1:0] node267;
	wire [3-1:0] node270;
	wire [3-1:0] node272;
	wire [3-1:0] node275;
	wire [3-1:0] node276;
	wire [3-1:0] node277;
	wire [3-1:0] node278;
	wire [3-1:0] node279;
	wire [3-1:0] node280;
	wire [3-1:0] node281;
	wire [3-1:0] node285;
	wire [3-1:0] node287;
	wire [3-1:0] node288;
	wire [3-1:0] node291;
	wire [3-1:0] node294;
	wire [3-1:0] node295;
	wire [3-1:0] node296;
	wire [3-1:0] node300;
	wire [3-1:0] node301;
	wire [3-1:0] node304;
	wire [3-1:0] node307;
	wire [3-1:0] node308;
	wire [3-1:0] node309;
	wire [3-1:0] node310;
	wire [3-1:0] node313;
	wire [3-1:0] node316;
	wire [3-1:0] node317;
	wire [3-1:0] node319;
	wire [3-1:0] node323;
	wire [3-1:0] node324;
	wire [3-1:0] node325;
	wire [3-1:0] node329;
	wire [3-1:0] node331;
	wire [3-1:0] node332;
	wire [3-1:0] node335;
	wire [3-1:0] node338;
	wire [3-1:0] node339;
	wire [3-1:0] node340;
	wire [3-1:0] node341;
	wire [3-1:0] node342;
	wire [3-1:0] node345;
	wire [3-1:0] node348;
	wire [3-1:0] node349;
	wire [3-1:0] node350;
	wire [3-1:0] node353;
	wire [3-1:0] node356;
	wire [3-1:0] node357;
	wire [3-1:0] node360;
	wire [3-1:0] node363;
	wire [3-1:0] node364;
	wire [3-1:0] node365;
	wire [3-1:0] node368;
	wire [3-1:0] node371;
	wire [3-1:0] node372;
	wire [3-1:0] node374;
	wire [3-1:0] node377;
	wire [3-1:0] node380;
	wire [3-1:0] node381;
	wire [3-1:0] node382;
	wire [3-1:0] node384;
	wire [3-1:0] node385;
	wire [3-1:0] node388;
	wire [3-1:0] node391;
	wire [3-1:0] node392;
	wire [3-1:0] node394;
	wire [3-1:0] node397;
	wire [3-1:0] node400;
	wire [3-1:0] node401;
	wire [3-1:0] node403;
	wire [3-1:0] node404;
	wire [3-1:0] node407;
	wire [3-1:0] node410;
	wire [3-1:0] node411;
	wire [3-1:0] node412;
	wire [3-1:0] node415;
	wire [3-1:0] node418;
	wire [3-1:0] node419;
	wire [3-1:0] node422;
	wire [3-1:0] node425;
	wire [3-1:0] node426;
	wire [3-1:0] node427;
	wire [3-1:0] node428;
	wire [3-1:0] node429;
	wire [3-1:0] node431;
	wire [3-1:0] node434;
	wire [3-1:0] node436;
	wire [3-1:0] node439;
	wire [3-1:0] node440;
	wire [3-1:0] node442;
	wire [3-1:0] node445;
	wire [3-1:0] node446;
	wire [3-1:0] node449;
	wire [3-1:0] node452;
	wire [3-1:0] node453;
	wire [3-1:0] node454;
	wire [3-1:0] node455;
	wire [3-1:0] node457;
	wire [3-1:0] node460;
	wire [3-1:0] node462;
	wire [3-1:0] node465;
	wire [3-1:0] node466;
	wire [3-1:0] node469;
	wire [3-1:0] node471;
	wire [3-1:0] node474;
	wire [3-1:0] node475;
	wire [3-1:0] node477;
	wire [3-1:0] node478;
	wire [3-1:0] node482;
	wire [3-1:0] node483;
	wire [3-1:0] node486;
	wire [3-1:0] node489;
	wire [3-1:0] node490;
	wire [3-1:0] node491;
	wire [3-1:0] node492;
	wire [3-1:0] node494;
	wire [3-1:0] node497;
	wire [3-1:0] node499;
	wire [3-1:0] node501;
	wire [3-1:0] node504;
	wire [3-1:0] node505;
	wire [3-1:0] node506;
	wire [3-1:0] node510;
	wire [3-1:0] node511;
	wire [3-1:0] node515;
	wire [3-1:0] node516;
	wire [3-1:0] node517;
	wire [3-1:0] node518;
	wire [3-1:0] node521;
	wire [3-1:0] node522;
	wire [3-1:0] node526;
	wire [3-1:0] node527;
	wire [3-1:0] node530;
	wire [3-1:0] node533;
	wire [3-1:0] node534;
	wire [3-1:0] node536;
	wire [3-1:0] node537;
	wire [3-1:0] node540;
	wire [3-1:0] node543;
	wire [3-1:0] node544;
	wire [3-1:0] node546;
	wire [3-1:0] node549;
	wire [3-1:0] node551;
	wire [3-1:0] node554;
	wire [3-1:0] node555;
	wire [3-1:0] node556;
	wire [3-1:0] node557;
	wire [3-1:0] node558;
	wire [3-1:0] node559;
	wire [3-1:0] node562;
	wire [3-1:0] node564;
	wire [3-1:0] node567;
	wire [3-1:0] node568;
	wire [3-1:0] node569;
	wire [3-1:0] node572;
	wire [3-1:0] node575;
	wire [3-1:0] node576;
	wire [3-1:0] node579;
	wire [3-1:0] node582;
	wire [3-1:0] node583;
	wire [3-1:0] node584;
	wire [3-1:0] node587;
	wire [3-1:0] node589;
	wire [3-1:0] node592;
	wire [3-1:0] node593;
	wire [3-1:0] node594;
	wire [3-1:0] node597;
	wire [3-1:0] node600;
	wire [3-1:0] node601;
	wire [3-1:0] node604;
	wire [3-1:0] node607;
	wire [3-1:0] node608;
	wire [3-1:0] node609;
	wire [3-1:0] node610;
	wire [3-1:0] node611;
	wire [3-1:0] node614;
	wire [3-1:0] node617;
	wire [3-1:0] node618;
	wire [3-1:0] node621;
	wire [3-1:0] node624;
	wire [3-1:0] node625;
	wire [3-1:0] node626;
	wire [3-1:0] node629;
	wire [3-1:0] node632;
	wire [3-1:0] node633;
	wire [3-1:0] node636;
	wire [3-1:0] node639;
	wire [3-1:0] node640;
	wire [3-1:0] node641;
	wire [3-1:0] node644;
	wire [3-1:0] node646;
	wire [3-1:0] node649;
	wire [3-1:0] node650;
	wire [3-1:0] node651;
	wire [3-1:0] node654;
	wire [3-1:0] node657;
	wire [3-1:0] node658;
	wire [3-1:0] node661;
	wire [3-1:0] node664;
	wire [3-1:0] node665;
	wire [3-1:0] node666;
	wire [3-1:0] node667;
	wire [3-1:0] node668;
	wire [3-1:0] node669;
	wire [3-1:0] node670;
	wire [3-1:0] node673;
	wire [3-1:0] node675;
	wire [3-1:0] node678;
	wire [3-1:0] node679;
	wire [3-1:0] node681;
	wire [3-1:0] node684;
	wire [3-1:0] node685;
	wire [3-1:0] node689;
	wire [3-1:0] node690;
	wire [3-1:0] node691;
	wire [3-1:0] node694;
	wire [3-1:0] node697;
	wire [3-1:0] node699;
	wire [3-1:0] node702;
	wire [3-1:0] node703;
	wire [3-1:0] node704;
	wire [3-1:0] node708;
	wire [3-1:0] node709;
	wire [3-1:0] node710;
	wire [3-1:0] node713;
	wire [3-1:0] node716;
	wire [3-1:0] node717;
	wire [3-1:0] node720;
	wire [3-1:0] node723;
	wire [3-1:0] node724;
	wire [3-1:0] node725;
	wire [3-1:0] node726;
	wire [3-1:0] node727;
	wire [3-1:0] node730;
	wire [3-1:0] node733;
	wire [3-1:0] node734;
	wire [3-1:0] node738;
	wire [3-1:0] node739;
	wire [3-1:0] node740;
	wire [3-1:0] node743;
	wire [3-1:0] node746;
	wire [3-1:0] node748;
	wire [3-1:0] node751;
	wire [3-1:0] node752;
	wire [3-1:0] node753;
	wire [3-1:0] node756;
	wire [3-1:0] node758;
	wire [3-1:0] node761;
	wire [3-1:0] node762;
	wire [3-1:0] node763;
	wire [3-1:0] node766;
	wire [3-1:0] node769;
	wire [3-1:0] node770;
	wire [3-1:0] node773;
	wire [3-1:0] node776;
	wire [3-1:0] node777;
	wire [3-1:0] node778;
	wire [3-1:0] node779;
	wire [3-1:0] node780;
	wire [3-1:0] node781;
	wire [3-1:0] node785;
	wire [3-1:0] node786;
	wire [3-1:0] node787;
	wire [3-1:0] node790;
	wire [3-1:0] node793;
	wire [3-1:0] node794;
	wire [3-1:0] node797;
	wire [3-1:0] node800;
	wire [3-1:0] node801;
	wire [3-1:0] node802;
	wire [3-1:0] node803;
	wire [3-1:0] node806;
	wire [3-1:0] node809;
	wire [3-1:0] node810;
	wire [3-1:0] node813;
	wire [3-1:0] node816;
	wire [3-1:0] node817;
	wire [3-1:0] node818;
	wire [3-1:0] node821;
	wire [3-1:0] node824;
	wire [3-1:0] node825;
	wire [3-1:0] node828;
	wire [3-1:0] node831;
	wire [3-1:0] node832;
	wire [3-1:0] node833;
	wire [3-1:0] node834;
	wire [3-1:0] node837;
	wire [3-1:0] node840;
	wire [3-1:0] node841;
	wire [3-1:0] node842;
	wire [3-1:0] node846;
	wire [3-1:0] node847;
	wire [3-1:0] node850;
	wire [3-1:0] node853;
	wire [3-1:0] node854;
	wire [3-1:0] node855;
	wire [3-1:0] node858;
	wire [3-1:0] node861;
	wire [3-1:0] node862;
	wire [3-1:0] node863;
	wire [3-1:0] node867;
	wire [3-1:0] node868;
	wire [3-1:0] node872;
	wire [3-1:0] node873;
	wire [3-1:0] node874;
	wire [3-1:0] node875;
	wire [3-1:0] node877;
	wire [3-1:0] node878;
	wire [3-1:0] node883;
	wire [3-1:0] node884;
	wire [3-1:0] node885;
	wire [3-1:0] node886;
	wire [3-1:0] node891;
	wire [3-1:0] node892;
	wire [3-1:0] node893;
	wire [3-1:0] node897;
	wire [3-1:0] node898;
	wire [3-1:0] node902;
	wire [3-1:0] node903;
	wire [3-1:0] node904;
	wire [3-1:0] node905;
	wire [3-1:0] node908;
	wire [3-1:0] node909;
	wire [3-1:0] node913;
	wire [3-1:0] node915;
	wire [3-1:0] node918;
	wire [3-1:0] node919;
	wire [3-1:0] node921;
	wire [3-1:0] node922;
	wire [3-1:0] node926;
	wire [3-1:0] node927;
	wire [3-1:0] node930;
	wire [3-1:0] node933;
	wire [3-1:0] node934;
	wire [3-1:0] node935;
	wire [3-1:0] node936;
	wire [3-1:0] node937;
	wire [3-1:0] node938;
	wire [3-1:0] node939;
	wire [3-1:0] node940;
	wire [3-1:0] node941;
	wire [3-1:0] node944;
	wire [3-1:0] node947;
	wire [3-1:0] node948;
	wire [3-1:0] node950;
	wire [3-1:0] node954;
	wire [3-1:0] node955;
	wire [3-1:0] node958;
	wire [3-1:0] node959;
	wire [3-1:0] node961;
	wire [3-1:0] node964;
	wire [3-1:0] node967;
	wire [3-1:0] node968;
	wire [3-1:0] node969;
	wire [3-1:0] node970;
	wire [3-1:0] node972;
	wire [3-1:0] node975;
	wire [3-1:0] node977;
	wire [3-1:0] node980;
	wire [3-1:0] node981;
	wire [3-1:0] node983;
	wire [3-1:0] node986;
	wire [3-1:0] node988;
	wire [3-1:0] node991;
	wire [3-1:0] node992;
	wire [3-1:0] node994;
	wire [3-1:0] node995;
	wire [3-1:0] node998;
	wire [3-1:0] node1001;
	wire [3-1:0] node1002;
	wire [3-1:0] node1005;
	wire [3-1:0] node1007;
	wire [3-1:0] node1010;
	wire [3-1:0] node1011;
	wire [3-1:0] node1012;
	wire [3-1:0] node1013;
	wire [3-1:0] node1014;
	wire [3-1:0] node1017;
	wire [3-1:0] node1020;
	wire [3-1:0] node1022;
	wire [3-1:0] node1023;
	wire [3-1:0] node1026;
	wire [3-1:0] node1029;
	wire [3-1:0] node1030;
	wire [3-1:0] node1031;
	wire [3-1:0] node1033;
	wire [3-1:0] node1037;
	wire [3-1:0] node1038;
	wire [3-1:0] node1040;
	wire [3-1:0] node1043;
	wire [3-1:0] node1045;
	wire [3-1:0] node1048;
	wire [3-1:0] node1049;
	wire [3-1:0] node1050;
	wire [3-1:0] node1051;
	wire [3-1:0] node1053;
	wire [3-1:0] node1056;
	wire [3-1:0] node1058;
	wire [3-1:0] node1061;
	wire [3-1:0] node1062;
	wire [3-1:0] node1065;
	wire [3-1:0] node1067;
	wire [3-1:0] node1070;
	wire [3-1:0] node1071;
	wire [3-1:0] node1072;
	wire [3-1:0] node1073;
	wire [3-1:0] node1076;
	wire [3-1:0] node1079;
	wire [3-1:0] node1081;
	wire [3-1:0] node1084;
	wire [3-1:0] node1086;
	wire [3-1:0] node1088;
	wire [3-1:0] node1091;
	wire [3-1:0] node1092;
	wire [3-1:0] node1093;
	wire [3-1:0] node1094;
	wire [3-1:0] node1095;
	wire [3-1:0] node1097;
	wire [3-1:0] node1100;
	wire [3-1:0] node1102;
	wire [3-1:0] node1105;
	wire [3-1:0] node1106;
	wire [3-1:0] node1108;
	wire [3-1:0] node1110;
	wire [3-1:0] node1113;
	wire [3-1:0] node1115;
	wire [3-1:0] node1118;
	wire [3-1:0] node1119;
	wire [3-1:0] node1120;
	wire [3-1:0] node1121;
	wire [3-1:0] node1125;
	wire [3-1:0] node1126;
	wire [3-1:0] node1128;
	wire [3-1:0] node1131;
	wire [3-1:0] node1133;
	wire [3-1:0] node1136;
	wire [3-1:0] node1137;
	wire [3-1:0] node1138;
	wire [3-1:0] node1141;
	wire [3-1:0] node1144;
	wire [3-1:0] node1145;
	wire [3-1:0] node1146;
	wire [3-1:0] node1149;
	wire [3-1:0] node1152;
	wire [3-1:0] node1153;
	wire [3-1:0] node1156;
	wire [3-1:0] node1159;
	wire [3-1:0] node1160;
	wire [3-1:0] node1161;
	wire [3-1:0] node1162;
	wire [3-1:0] node1164;
	wire [3-1:0] node1167;
	wire [3-1:0] node1169;
	wire [3-1:0] node1172;
	wire [3-1:0] node1174;
	wire [3-1:0] node1175;
	wire [3-1:0] node1178;
	wire [3-1:0] node1181;
	wire [3-1:0] node1182;
	wire [3-1:0] node1183;
	wire [3-1:0] node1184;
	wire [3-1:0] node1188;
	wire [3-1:0] node1189;
	wire [3-1:0] node1192;
	wire [3-1:0] node1193;
	wire [3-1:0] node1196;
	wire [3-1:0] node1199;
	wire [3-1:0] node1200;
	wire [3-1:0] node1202;
	wire [3-1:0] node1204;
	wire [3-1:0] node1207;
	wire [3-1:0] node1208;
	wire [3-1:0] node1209;
	wire [3-1:0] node1214;
	wire [3-1:0] node1215;
	wire [3-1:0] node1216;
	wire [3-1:0] node1217;
	wire [3-1:0] node1218;
	wire [3-1:0] node1219;
	wire [3-1:0] node1220;
	wire [3-1:0] node1224;
	wire [3-1:0] node1225;
	wire [3-1:0] node1226;
	wire [3-1:0] node1231;
	wire [3-1:0] node1232;
	wire [3-1:0] node1233;
	wire [3-1:0] node1234;
	wire [3-1:0] node1238;
	wire [3-1:0] node1239;
	wire [3-1:0] node1244;
	wire [3-1:0] node1245;
	wire [3-1:0] node1246;
	wire [3-1:0] node1248;
	wire [3-1:0] node1251;
	wire [3-1:0] node1252;
	wire [3-1:0] node1253;
	wire [3-1:0] node1258;
	wire [3-1:0] node1259;
	wire [3-1:0] node1260;
	wire [3-1:0] node1261;
	wire [3-1:0] node1265;
	wire [3-1:0] node1266;
	wire [3-1:0] node1270;
	wire [3-1:0] node1271;
	wire [3-1:0] node1272;
	wire [3-1:0] node1277;
	wire [3-1:0] node1278;
	wire [3-1:0] node1279;
	wire [3-1:0] node1280;
	wire [3-1:0] node1281;
	wire [3-1:0] node1285;
	wire [3-1:0] node1286;
	wire [3-1:0] node1287;
	wire [3-1:0] node1292;
	wire [3-1:0] node1293;
	wire [3-1:0] node1295;
	wire [3-1:0] node1298;
	wire [3-1:0] node1300;
	wire [3-1:0] node1303;
	wire [3-1:0] node1304;
	wire [3-1:0] node1305;
	wire [3-1:0] node1307;
	wire [3-1:0] node1310;
	wire [3-1:0] node1311;
	wire [3-1:0] node1315;
	wire [3-1:0] node1316;
	wire [3-1:0] node1317;
	wire [3-1:0] node1321;
	wire [3-1:0] node1324;
	wire [3-1:0] node1325;
	wire [3-1:0] node1326;
	wire [3-1:0] node1327;
	wire [3-1:0] node1328;
	wire [3-1:0] node1329;
	wire [3-1:0] node1331;
	wire [3-1:0] node1334;
	wire [3-1:0] node1336;
	wire [3-1:0] node1339;
	wire [3-1:0] node1341;
	wire [3-1:0] node1343;
	wire [3-1:0] node1346;
	wire [3-1:0] node1347;
	wire [3-1:0] node1349;
	wire [3-1:0] node1352;
	wire [3-1:0] node1354;
	wire [3-1:0] node1357;
	wire [3-1:0] node1358;
	wire [3-1:0] node1359;
	wire [3-1:0] node1360;
	wire [3-1:0] node1362;
	wire [3-1:0] node1366;
	wire [3-1:0] node1368;
	wire [3-1:0] node1371;
	wire [3-1:0] node1372;
	wire [3-1:0] node1373;
	wire [3-1:0] node1377;
	wire [3-1:0] node1378;
	wire [3-1:0] node1382;
	wire [3-1:0] node1383;
	wire [3-1:0] node1384;
	wire [3-1:0] node1385;
	wire [3-1:0] node1387;
	wire [3-1:0] node1390;
	wire [3-1:0] node1391;
	wire [3-1:0] node1392;
	wire [3-1:0] node1395;
	wire [3-1:0] node1399;
	wire [3-1:0] node1400;
	wire [3-1:0] node1401;
	wire [3-1:0] node1405;
	wire [3-1:0] node1408;
	wire [3-1:0] node1409;
	wire [3-1:0] node1410;
	wire [3-1:0] node1411;
	wire [3-1:0] node1414;
	wire [3-1:0] node1415;
	wire [3-1:0] node1419;
	wire [3-1:0] node1421;
	wire [3-1:0] node1422;
	wire [3-1:0] node1426;
	wire [3-1:0] node1427;
	wire [3-1:0] node1428;
	wire [3-1:0] node1432;
	wire [3-1:0] node1433;
	wire [3-1:0] node1437;
	wire [3-1:0] node1438;
	wire [3-1:0] node1439;
	wire [3-1:0] node1440;
	wire [3-1:0] node1441;
	wire [3-1:0] node1442;
	wire [3-1:0] node1443;
	wire [3-1:0] node1444;
	wire [3-1:0] node1445;
	wire [3-1:0] node1449;
	wire [3-1:0] node1450;
	wire [3-1:0] node1455;
	wire [3-1:0] node1456;
	wire [3-1:0] node1459;
	wire [3-1:0] node1461;
	wire [3-1:0] node1462;
	wire [3-1:0] node1466;
	wire [3-1:0] node1467;
	wire [3-1:0] node1468;
	wire [3-1:0] node1469;
	wire [3-1:0] node1473;
	wire [3-1:0] node1474;
	wire [3-1:0] node1478;
	wire [3-1:0] node1479;
	wire [3-1:0] node1480;
	wire [3-1:0] node1484;
	wire [3-1:0] node1485;
	wire [3-1:0] node1489;
	wire [3-1:0] node1490;
	wire [3-1:0] node1491;
	wire [3-1:0] node1493;
	wire [3-1:0] node1494;
	wire [3-1:0] node1498;
	wire [3-1:0] node1499;
	wire [3-1:0] node1500;
	wire [3-1:0] node1504;
	wire [3-1:0] node1505;
	wire [3-1:0] node1509;
	wire [3-1:0] node1510;
	wire [3-1:0] node1511;
	wire [3-1:0] node1512;
	wire [3-1:0] node1514;
	wire [3-1:0] node1517;
	wire [3-1:0] node1520;
	wire [3-1:0] node1522;
	wire [3-1:0] node1525;
	wire [3-1:0] node1526;
	wire [3-1:0] node1529;
	wire [3-1:0] node1532;
	wire [3-1:0] node1533;
	wire [3-1:0] node1534;
	wire [3-1:0] node1535;
	wire [3-1:0] node1536;
	wire [3-1:0] node1537;
	wire [3-1:0] node1541;
	wire [3-1:0] node1542;
	wire [3-1:0] node1546;
	wire [3-1:0] node1547;
	wire [3-1:0] node1548;
	wire [3-1:0] node1552;
	wire [3-1:0] node1553;
	wire [3-1:0] node1557;
	wire [3-1:0] node1558;
	wire [3-1:0] node1559;
	wire [3-1:0] node1560;
	wire [3-1:0] node1564;
	wire [3-1:0] node1565;
	wire [3-1:0] node1569;
	wire [3-1:0] node1570;
	wire [3-1:0] node1573;
	wire [3-1:0] node1575;
	wire [3-1:0] node1578;
	wire [3-1:0] node1579;
	wire [3-1:0] node1580;
	wire [3-1:0] node1581;
	wire [3-1:0] node1582;
	wire [3-1:0] node1586;
	wire [3-1:0] node1589;
	wire [3-1:0] node1590;
	wire [3-1:0] node1591;
	wire [3-1:0] node1595;
	wire [3-1:0] node1596;
	wire [3-1:0] node1600;
	wire [3-1:0] node1601;
	wire [3-1:0] node1602;
	wire [3-1:0] node1603;
	wire [3-1:0] node1607;
	wire [3-1:0] node1608;
	wire [3-1:0] node1612;
	wire [3-1:0] node1613;
	wire [3-1:0] node1614;
	wire [3-1:0] node1618;
	wire [3-1:0] node1619;
	wire [3-1:0] node1623;
	wire [3-1:0] node1624;
	wire [3-1:0] node1625;
	wire [3-1:0] node1626;
	wire [3-1:0] node1627;
	wire [3-1:0] node1628;
	wire [3-1:0] node1629;
	wire [3-1:0] node1631;
	wire [3-1:0] node1634;
	wire [3-1:0] node1636;
	wire [3-1:0] node1639;
	wire [3-1:0] node1640;
	wire [3-1:0] node1641;
	wire [3-1:0] node1645;
	wire [3-1:0] node1646;
	wire [3-1:0] node1649;
	wire [3-1:0] node1652;
	wire [3-1:0] node1653;
	wire [3-1:0] node1654;
	wire [3-1:0] node1655;
	wire [3-1:0] node1659;
	wire [3-1:0] node1660;
	wire [3-1:0] node1664;
	wire [3-1:0] node1665;
	wire [3-1:0] node1668;
	wire [3-1:0] node1669;
	wire [3-1:0] node1673;
	wire [3-1:0] node1674;
	wire [3-1:0] node1675;
	wire [3-1:0] node1676;
	wire [3-1:0] node1680;
	wire [3-1:0] node1683;
	wire [3-1:0] node1684;
	wire [3-1:0] node1685;
	wire [3-1:0] node1689;
	wire [3-1:0] node1690;
	wire [3-1:0] node1694;
	wire [3-1:0] node1695;
	wire [3-1:0] node1696;
	wire [3-1:0] node1697;
	wire [3-1:0] node1698;
	wire [3-1:0] node1702;
	wire [3-1:0] node1703;
	wire [3-1:0] node1707;
	wire [3-1:0] node1708;
	wire [3-1:0] node1709;
	wire [3-1:0] node1713;
	wire [3-1:0] node1716;
	wire [3-1:0] node1717;
	wire [3-1:0] node1718;
	wire [3-1:0] node1719;
	wire [3-1:0] node1724;
	wire [3-1:0] node1725;
	wire [3-1:0] node1726;
	wire [3-1:0] node1730;
	wire [3-1:0] node1731;
	wire [3-1:0] node1735;
	wire [3-1:0] node1736;
	wire [3-1:0] node1737;
	wire [3-1:0] node1738;
	wire [3-1:0] node1739;
	wire [3-1:0] node1740;
	wire [3-1:0] node1743;
	wire [3-1:0] node1746;
	wire [3-1:0] node1747;
	wire [3-1:0] node1750;
	wire [3-1:0] node1753;
	wire [3-1:0] node1754;
	wire [3-1:0] node1757;
	wire [3-1:0] node1760;
	wire [3-1:0] node1761;
	wire [3-1:0] node1762;
	wire [3-1:0] node1763;
	wire [3-1:0] node1764;
	wire [3-1:0] node1769;
	wire [3-1:0] node1770;
	wire [3-1:0] node1774;
	wire [3-1:0] node1775;
	wire [3-1:0] node1776;
	wire [3-1:0] node1780;
	wire [3-1:0] node1781;
	wire [3-1:0] node1785;
	wire [3-1:0] node1786;
	wire [3-1:0] node1787;
	wire [3-1:0] node1788;
	wire [3-1:0] node1789;
	wire [3-1:0] node1793;
	wire [3-1:0] node1794;
	wire [3-1:0] node1798;
	wire [3-1:0] node1799;
	wire [3-1:0] node1800;
	wire [3-1:0] node1804;
	wire [3-1:0] node1805;
	wire [3-1:0] node1809;
	wire [3-1:0] node1810;
	wire [3-1:0] node1811;
	wire [3-1:0] node1812;
	wire [3-1:0] node1815;
	wire [3-1:0] node1818;
	wire [3-1:0] node1819;
	wire [3-1:0] node1822;
	wire [3-1:0] node1825;
	wire [3-1:0] node1826;
	wire [3-1:0] node1829;
	wire [3-1:0] node1832;
	wire [3-1:0] node1833;
	wire [3-1:0] node1834;
	wire [3-1:0] node1835;
	wire [3-1:0] node1836;
	wire [3-1:0] node1837;
	wire [3-1:0] node1838;
	wire [3-1:0] node1839;
	wire [3-1:0] node1840;
	wire [3-1:0] node1843;
	wire [3-1:0] node1846;
	wire [3-1:0] node1847;
	wire [3-1:0] node1848;
	wire [3-1:0] node1849;
	wire [3-1:0] node1852;
	wire [3-1:0] node1855;
	wire [3-1:0] node1856;
	wire [3-1:0] node1859;
	wire [3-1:0] node1862;
	wire [3-1:0] node1863;
	wire [3-1:0] node1867;
	wire [3-1:0] node1868;
	wire [3-1:0] node1869;
	wire [3-1:0] node1870;
	wire [3-1:0] node1873;
	wire [3-1:0] node1876;
	wire [3-1:0] node1877;
	wire [3-1:0] node1880;
	wire [3-1:0] node1883;
	wire [3-1:0] node1884;
	wire [3-1:0] node1886;
	wire [3-1:0] node1887;
	wire [3-1:0] node1890;
	wire [3-1:0] node1893;
	wire [3-1:0] node1894;
	wire [3-1:0] node1895;
	wire [3-1:0] node1898;
	wire [3-1:0] node1901;
	wire [3-1:0] node1903;
	wire [3-1:0] node1906;
	wire [3-1:0] node1907;
	wire [3-1:0] node1908;
	wire [3-1:0] node1909;
	wire [3-1:0] node1911;
	wire [3-1:0] node1914;
	wire [3-1:0] node1916;
	wire [3-1:0] node1919;
	wire [3-1:0] node1920;
	wire [3-1:0] node1922;
	wire [3-1:0] node1925;
	wire [3-1:0] node1927;
	wire [3-1:0] node1930;
	wire [3-1:0] node1931;
	wire [3-1:0] node1932;
	wire [3-1:0] node1933;
	wire [3-1:0] node1937;
	wire [3-1:0] node1940;
	wire [3-1:0] node1941;
	wire [3-1:0] node1942;
	wire [3-1:0] node1946;
	wire [3-1:0] node1947;
	wire [3-1:0] node1951;
	wire [3-1:0] node1952;
	wire [3-1:0] node1953;
	wire [3-1:0] node1954;
	wire [3-1:0] node1955;
	wire [3-1:0] node1956;
	wire [3-1:0] node1958;
	wire [3-1:0] node1961;
	wire [3-1:0] node1962;
	wire [3-1:0] node1966;
	wire [3-1:0] node1967;
	wire [3-1:0] node1968;
	wire [3-1:0] node1971;
	wire [3-1:0] node1975;
	wire [3-1:0] node1976;
	wire [3-1:0] node1977;
	wire [3-1:0] node1979;
	wire [3-1:0] node1983;
	wire [3-1:0] node1984;
	wire [3-1:0] node1986;
	wire [3-1:0] node1989;
	wire [3-1:0] node1990;
	wire [3-1:0] node1993;
	wire [3-1:0] node1996;
	wire [3-1:0] node1997;
	wire [3-1:0] node1998;
	wire [3-1:0] node1999;
	wire [3-1:0] node2000;
	wire [3-1:0] node2003;
	wire [3-1:0] node2008;
	wire [3-1:0] node2009;
	wire [3-1:0] node2010;
	wire [3-1:0] node2011;
	wire [3-1:0] node2014;
	wire [3-1:0] node2018;
	wire [3-1:0] node2019;
	wire [3-1:0] node2020;
	wire [3-1:0] node2023;
	wire [3-1:0] node2027;
	wire [3-1:0] node2028;
	wire [3-1:0] node2029;
	wire [3-1:0] node2030;
	wire [3-1:0] node2032;
	wire [3-1:0] node2033;
	wire [3-1:0] node2036;
	wire [3-1:0] node2039;
	wire [3-1:0] node2040;
	wire [3-1:0] node2043;
	wire [3-1:0] node2045;
	wire [3-1:0] node2048;
	wire [3-1:0] node2049;
	wire [3-1:0] node2050;
	wire [3-1:0] node2051;
	wire [3-1:0] node2055;
	wire [3-1:0] node2058;
	wire [3-1:0] node2059;
	wire [3-1:0] node2060;
	wire [3-1:0] node2063;
	wire [3-1:0] node2066;
	wire [3-1:0] node2068;
	wire [3-1:0] node2071;
	wire [3-1:0] node2072;
	wire [3-1:0] node2073;
	wire [3-1:0] node2074;
	wire [3-1:0] node2075;
	wire [3-1:0] node2079;
	wire [3-1:0] node2080;
	wire [3-1:0] node2083;
	wire [3-1:0] node2086;
	wire [3-1:0] node2087;
	wire [3-1:0] node2090;
	wire [3-1:0] node2093;
	wire [3-1:0] node2094;
	wire [3-1:0] node2095;
	wire [3-1:0] node2098;
	wire [3-1:0] node2101;
	wire [3-1:0] node2102;
	wire [3-1:0] node2103;
	wire [3-1:0] node2106;
	wire [3-1:0] node2109;
	wire [3-1:0] node2110;
	wire [3-1:0] node2113;
	wire [3-1:0] node2116;
	wire [3-1:0] node2117;
	wire [3-1:0] node2118;
	wire [3-1:0] node2119;
	wire [3-1:0] node2120;
	wire [3-1:0] node2121;
	wire [3-1:0] node2122;
	wire [3-1:0] node2123;
	wire [3-1:0] node2126;
	wire [3-1:0] node2129;
	wire [3-1:0] node2130;
	wire [3-1:0] node2134;
	wire [3-1:0] node2136;
	wire [3-1:0] node2139;
	wire [3-1:0] node2140;
	wire [3-1:0] node2141;
	wire [3-1:0] node2142;
	wire [3-1:0] node2146;
	wire [3-1:0] node2149;
	wire [3-1:0] node2150;
	wire [3-1:0] node2153;
	wire [3-1:0] node2154;
	wire [3-1:0] node2158;
	wire [3-1:0] node2159;
	wire [3-1:0] node2160;
	wire [3-1:0] node2161;
	wire [3-1:0] node2164;
	wire [3-1:0] node2167;
	wire [3-1:0] node2168;
	wire [3-1:0] node2171;
	wire [3-1:0] node2172;
	wire [3-1:0] node2176;
	wire [3-1:0] node2177;
	wire [3-1:0] node2180;
	wire [3-1:0] node2181;
	wire [3-1:0] node2185;
	wire [3-1:0] node2186;
	wire [3-1:0] node2187;
	wire [3-1:0] node2188;
	wire [3-1:0] node2189;
	wire [3-1:0] node2190;
	wire [3-1:0] node2194;
	wire [3-1:0] node2195;
	wire [3-1:0] node2199;
	wire [3-1:0] node2200;
	wire [3-1:0] node2204;
	wire [3-1:0] node2205;
	wire [3-1:0] node2206;
	wire [3-1:0] node2209;
	wire [3-1:0] node2210;
	wire [3-1:0] node2214;
	wire [3-1:0] node2215;
	wire [3-1:0] node2216;
	wire [3-1:0] node2221;
	wire [3-1:0] node2222;
	wire [3-1:0] node2223;
	wire [3-1:0] node2224;
	wire [3-1:0] node2228;
	wire [3-1:0] node2231;
	wire [3-1:0] node2232;
	wire [3-1:0] node2234;
	wire [3-1:0] node2237;
	wire [3-1:0] node2238;
	wire [3-1:0] node2239;
	wire [3-1:0] node2243;
	wire [3-1:0] node2246;
	wire [3-1:0] node2247;
	wire [3-1:0] node2248;
	wire [3-1:0] node2249;
	wire [3-1:0] node2250;
	wire [3-1:0] node2251;
	wire [3-1:0] node2252;
	wire [3-1:0] node2256;
	wire [3-1:0] node2257;
	wire [3-1:0] node2261;
	wire [3-1:0] node2262;
	wire [3-1:0] node2263;
	wire [3-1:0] node2267;
	wire [3-1:0] node2268;
	wire [3-1:0] node2272;
	wire [3-1:0] node2273;
	wire [3-1:0] node2274;
	wire [3-1:0] node2275;
	wire [3-1:0] node2279;
	wire [3-1:0] node2280;
	wire [3-1:0] node2285;
	wire [3-1:0] node2286;
	wire [3-1:0] node2287;
	wire [3-1:0] node2289;
	wire [3-1:0] node2290;
	wire [3-1:0] node2294;
	wire [3-1:0] node2296;
	wire [3-1:0] node2299;
	wire [3-1:0] node2300;
	wire [3-1:0] node2301;
	wire [3-1:0] node2302;
	wire [3-1:0] node2307;
	wire [3-1:0] node2308;
	wire [3-1:0] node2311;
	wire [3-1:0] node2314;
	wire [3-1:0] node2315;
	wire [3-1:0] node2316;
	wire [3-1:0] node2317;
	wire [3-1:0] node2318;
	wire [3-1:0] node2319;
	wire [3-1:0] node2323;
	wire [3-1:0] node2325;
	wire [3-1:0] node2328;
	wire [3-1:0] node2330;
	wire [3-1:0] node2333;
	wire [3-1:0] node2334;
	wire [3-1:0] node2335;
	wire [3-1:0] node2336;
	wire [3-1:0] node2340;
	wire [3-1:0] node2343;
	wire [3-1:0] node2345;
	wire [3-1:0] node2346;
	wire [3-1:0] node2350;
	wire [3-1:0] node2351;
	wire [3-1:0] node2352;
	wire [3-1:0] node2353;
	wire [3-1:0] node2356;
	wire [3-1:0] node2357;
	wire [3-1:0] node2361;
	wire [3-1:0] node2362;
	wire [3-1:0] node2363;
	wire [3-1:0] node2367;
	wire [3-1:0] node2368;
	wire [3-1:0] node2372;
	wire [3-1:0] node2373;
	wire [3-1:0] node2374;
	wire [3-1:0] node2378;
	wire [3-1:0] node2379;
	wire [3-1:0] node2383;
	wire [3-1:0] node2384;
	wire [3-1:0] node2385;
	wire [3-1:0] node2386;
	wire [3-1:0] node2387;
	wire [3-1:0] node2388;
	wire [3-1:0] node2389;
	wire [3-1:0] node2392;
	wire [3-1:0] node2394;
	wire [3-1:0] node2397;
	wire [3-1:0] node2398;
	wire [3-1:0] node2399;
	wire [3-1:0] node2403;
	wire [3-1:0] node2405;
	wire [3-1:0] node2406;
	wire [3-1:0] node2409;
	wire [3-1:0] node2412;
	wire [3-1:0] node2413;
	wire [3-1:0] node2414;
	wire [3-1:0] node2415;
	wire [3-1:0] node2418;
	wire [3-1:0] node2421;
	wire [3-1:0] node2422;
	wire [3-1:0] node2425;
	wire [3-1:0] node2428;
	wire [3-1:0] node2429;
	wire [3-1:0] node2430;
	wire [3-1:0] node2433;
	wire [3-1:0] node2436;
	wire [3-1:0] node2437;
	wire [3-1:0] node2440;
	wire [3-1:0] node2443;
	wire [3-1:0] node2444;
	wire [3-1:0] node2445;
	wire [3-1:0] node2446;
	wire [3-1:0] node2449;
	wire [3-1:0] node2451;
	wire [3-1:0] node2454;
	wire [3-1:0] node2455;
	wire [3-1:0] node2456;
	wire [3-1:0] node2460;
	wire [3-1:0] node2461;
	wire [3-1:0] node2464;
	wire [3-1:0] node2467;
	wire [3-1:0] node2468;
	wire [3-1:0] node2469;
	wire [3-1:0] node2470;
	wire [3-1:0] node2473;
	wire [3-1:0] node2476;
	wire [3-1:0] node2478;
	wire [3-1:0] node2481;
	wire [3-1:0] node2482;
	wire [3-1:0] node2483;
	wire [3-1:0] node2484;
	wire [3-1:0] node2489;
	wire [3-1:0] node2490;
	wire [3-1:0] node2494;
	wire [3-1:0] node2495;
	wire [3-1:0] node2496;
	wire [3-1:0] node2497;
	wire [3-1:0] node2498;
	wire [3-1:0] node2501;
	wire [3-1:0] node2504;
	wire [3-1:0] node2505;
	wire [3-1:0] node2508;
	wire [3-1:0] node2510;
	wire [3-1:0] node2513;
	wire [3-1:0] node2514;
	wire [3-1:0] node2515;
	wire [3-1:0] node2516;
	wire [3-1:0] node2517;
	wire [3-1:0] node2521;
	wire [3-1:0] node2522;
	wire [3-1:0] node2526;
	wire [3-1:0] node2527;
	wire [3-1:0] node2528;
	wire [3-1:0] node2532;
	wire [3-1:0] node2533;
	wire [3-1:0] node2537;
	wire [3-1:0] node2538;
	wire [3-1:0] node2540;
	wire [3-1:0] node2541;
	wire [3-1:0] node2545;
	wire [3-1:0] node2546;
	wire [3-1:0] node2547;
	wire [3-1:0] node2551;
	wire [3-1:0] node2552;
	wire [3-1:0] node2556;
	wire [3-1:0] node2557;
	wire [3-1:0] node2558;
	wire [3-1:0] node2559;
	wire [3-1:0] node2560;
	wire [3-1:0] node2561;
	wire [3-1:0] node2564;
	wire [3-1:0] node2567;
	wire [3-1:0] node2568;
	wire [3-1:0] node2572;
	wire [3-1:0] node2574;
	wire [3-1:0] node2577;
	wire [3-1:0] node2578;
	wire [3-1:0] node2579;
	wire [3-1:0] node2580;
	wire [3-1:0] node2583;
	wire [3-1:0] node2587;
	wire [3-1:0] node2588;
	wire [3-1:0] node2589;
	wire [3-1:0] node2593;
	wire [3-1:0] node2596;
	wire [3-1:0] node2597;
	wire [3-1:0] node2598;
	wire [3-1:0] node2599;
	wire [3-1:0] node2601;
	wire [3-1:0] node2604;
	wire [3-1:0] node2605;
	wire [3-1:0] node2609;
	wire [3-1:0] node2610;
	wire [3-1:0] node2611;
	wire [3-1:0] node2614;
	wire [3-1:0] node2617;
	wire [3-1:0] node2618;
	wire [3-1:0] node2622;
	wire [3-1:0] node2623;
	wire [3-1:0] node2626;
	wire [3-1:0] node2629;
	wire [3-1:0] node2630;
	wire [3-1:0] node2631;
	wire [3-1:0] node2632;
	wire [3-1:0] node2633;
	wire [3-1:0] node2634;
	wire [3-1:0] node2637;
	wire [3-1:0] node2640;
	wire [3-1:0] node2641;
	wire [3-1:0] node2642;
	wire [3-1:0] node2645;
	wire [3-1:0] node2648;
	wire [3-1:0] node2649;
	wire [3-1:0] node2653;
	wire [3-1:0] node2654;
	wire [3-1:0] node2655;
	wire [3-1:0] node2656;
	wire [3-1:0] node2661;
	wire [3-1:0] node2662;
	wire [3-1:0] node2663;
	wire [3-1:0] node2666;
	wire [3-1:0] node2669;
	wire [3-1:0] node2670;
	wire [3-1:0] node2671;
	wire [3-1:0] node2676;
	wire [3-1:0] node2677;
	wire [3-1:0] node2678;
	wire [3-1:0] node2680;
	wire [3-1:0] node2681;
	wire [3-1:0] node2684;
	wire [3-1:0] node2687;
	wire [3-1:0] node2688;
	wire [3-1:0] node2689;
	wire [3-1:0] node2690;
	wire [3-1:0] node2693;
	wire [3-1:0] node2697;
	wire [3-1:0] node2699;
	wire [3-1:0] node2702;
	wire [3-1:0] node2703;
	wire [3-1:0] node2704;
	wire [3-1:0] node2705;
	wire [3-1:0] node2708;
	wire [3-1:0] node2712;
	wire [3-1:0] node2713;
	wire [3-1:0] node2714;
	wire [3-1:0] node2717;
	wire [3-1:0] node2720;
	wire [3-1:0] node2721;
	wire [3-1:0] node2722;
	wire [3-1:0] node2726;
	wire [3-1:0] node2727;
	wire [3-1:0] node2730;
	wire [3-1:0] node2733;
	wire [3-1:0] node2734;
	wire [3-1:0] node2735;
	wire [3-1:0] node2736;
	wire [3-1:0] node2737;
	wire [3-1:0] node2740;
	wire [3-1:0] node2741;
	wire [3-1:0] node2742;
	wire [3-1:0] node2745;
	wire [3-1:0] node2748;
	wire [3-1:0] node2749;
	wire [3-1:0] node2752;
	wire [3-1:0] node2755;
	wire [3-1:0] node2756;
	wire [3-1:0] node2757;
	wire [3-1:0] node2758;
	wire [3-1:0] node2762;
	wire [3-1:0] node2763;
	wire [3-1:0] node2766;
	wire [3-1:0] node2769;
	wire [3-1:0] node2770;
	wire [3-1:0] node2771;
	wire [3-1:0] node2774;
	wire [3-1:0] node2777;
	wire [3-1:0] node2778;
	wire [3-1:0] node2782;
	wire [3-1:0] node2783;
	wire [3-1:0] node2784;
	wire [3-1:0] node2785;
	wire [3-1:0] node2786;
	wire [3-1:0] node2789;
	wire [3-1:0] node2792;
	wire [3-1:0] node2793;
	wire [3-1:0] node2797;
	wire [3-1:0] node2798;
	wire [3-1:0] node2802;
	wire [3-1:0] node2803;
	wire [3-1:0] node2804;
	wire [3-1:0] node2807;
	wire [3-1:0] node2810;
	wire [3-1:0] node2811;
	wire [3-1:0] node2814;
	wire [3-1:0] node2815;
	wire [3-1:0] node2819;
	wire [3-1:0] node2820;
	wire [3-1:0] node2821;
	wire [3-1:0] node2822;
	wire [3-1:0] node2823;
	wire [3-1:0] node2827;
	wire [3-1:0] node2830;
	wire [3-1:0] node2831;
	wire [3-1:0] node2832;
	wire [3-1:0] node2835;
	wire [3-1:0] node2839;
	wire [3-1:0] node2840;
	wire [3-1:0] node2841;
	wire [3-1:0] node2842;
	wire [3-1:0] node2846;
	wire [3-1:0] node2849;
	wire [3-1:0] node2850;
	wire [3-1:0] node2852;
	wire [3-1:0] node2855;
	wire [3-1:0] node2858;
	wire [3-1:0] node2859;
	wire [3-1:0] node2860;
	wire [3-1:0] node2861;
	wire [3-1:0] node2862;
	wire [3-1:0] node2863;
	wire [3-1:0] node2864;
	wire [3-1:0] node2865;
	wire [3-1:0] node2866;
	wire [3-1:0] node2869;
	wire [3-1:0] node2872;
	wire [3-1:0] node2873;
	wire [3-1:0] node2876;
	wire [3-1:0] node2879;
	wire [3-1:0] node2880;
	wire [3-1:0] node2882;
	wire [3-1:0] node2885;
	wire [3-1:0] node2886;
	wire [3-1:0] node2887;
	wire [3-1:0] node2890;
	wire [3-1:0] node2893;
	wire [3-1:0] node2894;
	wire [3-1:0] node2898;
	wire [3-1:0] node2899;
	wire [3-1:0] node2900;
	wire [3-1:0] node2901;
	wire [3-1:0] node2904;
	wire [3-1:0] node2907;
	wire [3-1:0] node2908;
	wire [3-1:0] node2909;
	wire [3-1:0] node2912;
	wire [3-1:0] node2916;
	wire [3-1:0] node2917;
	wire [3-1:0] node2918;
	wire [3-1:0] node2921;
	wire [3-1:0] node2924;
	wire [3-1:0] node2925;
	wire [3-1:0] node2929;
	wire [3-1:0] node2930;
	wire [3-1:0] node2931;
	wire [3-1:0] node2932;
	wire [3-1:0] node2933;
	wire [3-1:0] node2937;
	wire [3-1:0] node2939;
	wire [3-1:0] node2940;
	wire [3-1:0] node2944;
	wire [3-1:0] node2945;
	wire [3-1:0] node2946;
	wire [3-1:0] node2947;
	wire [3-1:0] node2950;
	wire [3-1:0] node2953;
	wire [3-1:0] node2954;
	wire [3-1:0] node2957;
	wire [3-1:0] node2960;
	wire [3-1:0] node2961;
	wire [3-1:0] node2965;
	wire [3-1:0] node2966;
	wire [3-1:0] node2967;
	wire [3-1:0] node2968;
	wire [3-1:0] node2969;
	wire [3-1:0] node2973;
	wire [3-1:0] node2974;
	wire [3-1:0] node2977;
	wire [3-1:0] node2980;
	wire [3-1:0] node2981;
	wire [3-1:0] node2985;
	wire [3-1:0] node2987;
	wire [3-1:0] node2988;
	wire [3-1:0] node2991;
	wire [3-1:0] node2994;
	wire [3-1:0] node2995;
	wire [3-1:0] node2996;
	wire [3-1:0] node2997;
	wire [3-1:0] node2998;
	wire [3-1:0] node2999;
	wire [3-1:0] node3000;
	wire [3-1:0] node3004;
	wire [3-1:0] node3005;
	wire [3-1:0] node3008;
	wire [3-1:0] node3011;
	wire [3-1:0] node3013;
	wire [3-1:0] node3015;
	wire [3-1:0] node3018;
	wire [3-1:0] node3019;
	wire [3-1:0] node3020;
	wire [3-1:0] node3024;
	wire [3-1:0] node3025;
	wire [3-1:0] node3026;
	wire [3-1:0] node3029;
	wire [3-1:0] node3032;
	wire [3-1:0] node3033;
	wire [3-1:0] node3036;
	wire [3-1:0] node3039;
	wire [3-1:0] node3040;
	wire [3-1:0] node3041;
	wire [3-1:0] node3042;
	wire [3-1:0] node3044;
	wire [3-1:0] node3048;
	wire [3-1:0] node3049;
	wire [3-1:0] node3052;
	wire [3-1:0] node3055;
	wire [3-1:0] node3056;
	wire [3-1:0] node3059;
	wire [3-1:0] node3062;
	wire [3-1:0] node3063;
	wire [3-1:0] node3064;
	wire [3-1:0] node3065;
	wire [3-1:0] node3066;
	wire [3-1:0] node3067;
	wire [3-1:0] node3070;
	wire [3-1:0] node3073;
	wire [3-1:0] node3075;
	wire [3-1:0] node3078;
	wire [3-1:0] node3079;
	wire [3-1:0] node3082;
	wire [3-1:0] node3085;
	wire [3-1:0] node3086;
	wire [3-1:0] node3087;
	wire [3-1:0] node3090;
	wire [3-1:0] node3093;
	wire [3-1:0] node3095;
	wire [3-1:0] node3098;
	wire [3-1:0] node3099;
	wire [3-1:0] node3100;
	wire [3-1:0] node3101;
	wire [3-1:0] node3102;
	wire [3-1:0] node3105;
	wire [3-1:0] node3109;
	wire [3-1:0] node3111;
	wire [3-1:0] node3114;
	wire [3-1:0] node3115;
	wire [3-1:0] node3118;
	wire [3-1:0] node3121;
	wire [3-1:0] node3122;
	wire [3-1:0] node3123;
	wire [3-1:0] node3124;
	wire [3-1:0] node3125;
	wire [3-1:0] node3126;
	wire [3-1:0] node3127;
	wire [3-1:0] node3129;
	wire [3-1:0] node3133;
	wire [3-1:0] node3134;
	wire [3-1:0] node3138;
	wire [3-1:0] node3139;
	wire [3-1:0] node3140;
	wire [3-1:0] node3142;
	wire [3-1:0] node3145;
	wire [3-1:0] node3146;
	wire [3-1:0] node3149;
	wire [3-1:0] node3153;
	wire [3-1:0] node3154;
	wire [3-1:0] node3155;
	wire [3-1:0] node3156;
	wire [3-1:0] node3158;
	wire [3-1:0] node3161;
	wire [3-1:0] node3164;
	wire [3-1:0] node3165;
	wire [3-1:0] node3167;
	wire [3-1:0] node3170;
	wire [3-1:0] node3173;
	wire [3-1:0] node3174;
	wire [3-1:0] node3177;
	wire [3-1:0] node3179;
	wire [3-1:0] node3180;
	wire [3-1:0] node3184;
	wire [3-1:0] node3185;
	wire [3-1:0] node3186;
	wire [3-1:0] node3187;
	wire [3-1:0] node3188;
	wire [3-1:0] node3189;
	wire [3-1:0] node3192;
	wire [3-1:0] node3195;
	wire [3-1:0] node3197;
	wire [3-1:0] node3200;
	wire [3-1:0] node3201;
	wire [3-1:0] node3204;
	wire [3-1:0] node3207;
	wire [3-1:0] node3208;
	wire [3-1:0] node3210;
	wire [3-1:0] node3213;
	wire [3-1:0] node3214;
	wire [3-1:0] node3215;
	wire [3-1:0] node3219;
	wire [3-1:0] node3220;
	wire [3-1:0] node3224;
	wire [3-1:0] node3225;
	wire [3-1:0] node3226;
	wire [3-1:0] node3227;
	wire [3-1:0] node3228;
	wire [3-1:0] node3231;
	wire [3-1:0] node3234;
	wire [3-1:0] node3235;
	wire [3-1:0] node3238;
	wire [3-1:0] node3241;
	wire [3-1:0] node3243;
	wire [3-1:0] node3246;
	wire [3-1:0] node3247;
	wire [3-1:0] node3248;
	wire [3-1:0] node3249;
	wire [3-1:0] node3253;
	wire [3-1:0] node3254;
	wire [3-1:0] node3258;
	wire [3-1:0] node3259;
	wire [3-1:0] node3262;
	wire [3-1:0] node3265;
	wire [3-1:0] node3266;
	wire [3-1:0] node3267;
	wire [3-1:0] node3268;
	wire [3-1:0] node3269;
	wire [3-1:0] node3270;
	wire [3-1:0] node3271;
	wire [3-1:0] node3275;
	wire [3-1:0] node3277;
	wire [3-1:0] node3280;
	wire [3-1:0] node3281;
	wire [3-1:0] node3282;
	wire [3-1:0] node3286;
	wire [3-1:0] node3287;
	wire [3-1:0] node3291;
	wire [3-1:0] node3292;
	wire [3-1:0] node3293;
	wire [3-1:0] node3294;
	wire [3-1:0] node3298;
	wire [3-1:0] node3300;
	wire [3-1:0] node3303;
	wire [3-1:0] node3304;
	wire [3-1:0] node3307;
	wire [3-1:0] node3310;
	wire [3-1:0] node3311;
	wire [3-1:0] node3312;
	wire [3-1:0] node3314;
	wire [3-1:0] node3315;
	wire [3-1:0] node3318;
	wire [3-1:0] node3321;
	wire [3-1:0] node3323;
	wire [3-1:0] node3326;
	wire [3-1:0] node3327;
	wire [3-1:0] node3330;
	wire [3-1:0] node3333;
	wire [3-1:0] node3334;
	wire [3-1:0] node3335;
	wire [3-1:0] node3336;
	wire [3-1:0] node3338;
	wire [3-1:0] node3339;
	wire [3-1:0] node3343;
	wire [3-1:0] node3344;
	wire [3-1:0] node3348;
	wire [3-1:0] node3349;
	wire [3-1:0] node3350;
	wire [3-1:0] node3351;
	wire [3-1:0] node3354;
	wire [3-1:0] node3357;
	wire [3-1:0] node3358;
	wire [3-1:0] node3362;
	wire [3-1:0] node3363;
	wire [3-1:0] node3366;
	wire [3-1:0] node3369;
	wire [3-1:0] node3370;
	wire [3-1:0] node3371;
	wire [3-1:0] node3373;
	wire [3-1:0] node3376;
	wire [3-1:0] node3378;
	wire [3-1:0] node3381;
	wire [3-1:0] node3382;
	wire [3-1:0] node3385;
	wire [3-1:0] node3388;
	wire [3-1:0] node3389;
	wire [3-1:0] node3390;
	wire [3-1:0] node3391;
	wire [3-1:0] node3392;
	wire [3-1:0] node3393;
	wire [3-1:0] node3394;
	wire [3-1:0] node3395;
	wire [3-1:0] node3398;
	wire [3-1:0] node3402;
	wire [3-1:0] node3403;
	wire [3-1:0] node3404;
	wire [3-1:0] node3405;
	wire [3-1:0] node3408;
	wire [3-1:0] node3411;
	wire [3-1:0] node3413;
	wire [3-1:0] node3416;
	wire [3-1:0] node3417;
	wire [3-1:0] node3421;
	wire [3-1:0] node3422;
	wire [3-1:0] node3423;
	wire [3-1:0] node3424;
	wire [3-1:0] node3428;
	wire [3-1:0] node3431;
	wire [3-1:0] node3432;
	wire [3-1:0] node3433;
	wire [3-1:0] node3437;
	wire [3-1:0] node3438;
	wire [3-1:0] node3442;
	wire [3-1:0] node3443;
	wire [3-1:0] node3444;
	wire [3-1:0] node3445;
	wire [3-1:0] node3447;
	wire [3-1:0] node3448;
	wire [3-1:0] node3452;
	wire [3-1:0] node3453;
	wire [3-1:0] node3456;
	wire [3-1:0] node3459;
	wire [3-1:0] node3460;
	wire [3-1:0] node3463;
	wire [3-1:0] node3466;
	wire [3-1:0] node3467;
	wire [3-1:0] node3469;
	wire [3-1:0] node3470;
	wire [3-1:0] node3474;
	wire [3-1:0] node3475;
	wire [3-1:0] node3477;
	wire [3-1:0] node3480;
	wire [3-1:0] node3481;
	wire [3-1:0] node3485;
	wire [3-1:0] node3486;
	wire [3-1:0] node3487;
	wire [3-1:0] node3488;
	wire [3-1:0] node3489;
	wire [3-1:0] node3491;
	wire [3-1:0] node3494;
	wire [3-1:0] node3495;
	wire [3-1:0] node3497;
	wire [3-1:0] node3500;
	wire [3-1:0] node3501;
	wire [3-1:0] node3504;
	wire [3-1:0] node3507;
	wire [3-1:0] node3508;
	wire [3-1:0] node3509;
	wire [3-1:0] node3510;
	wire [3-1:0] node3513;
	wire [3-1:0] node3516;
	wire [3-1:0] node3517;
	wire [3-1:0] node3521;
	wire [3-1:0] node3522;
	wire [3-1:0] node3525;
	wire [3-1:0] node3528;
	wire [3-1:0] node3529;
	wire [3-1:0] node3530;
	wire [3-1:0] node3531;
	wire [3-1:0] node3535;
	wire [3-1:0] node3536;
	wire [3-1:0] node3540;
	wire [3-1:0] node3541;
	wire [3-1:0] node3542;
	wire [3-1:0] node3546;
	wire [3-1:0] node3547;
	wire [3-1:0] node3551;
	wire [3-1:0] node3552;
	wire [3-1:0] node3553;
	wire [3-1:0] node3554;
	wire [3-1:0] node3555;
	wire [3-1:0] node3559;
	wire [3-1:0] node3560;
	wire [3-1:0] node3564;
	wire [3-1:0] node3565;
	wire [3-1:0] node3566;
	wire [3-1:0] node3570;
	wire [3-1:0] node3571;
	wire [3-1:0] node3575;
	wire [3-1:0] node3576;
	wire [3-1:0] node3577;
	wire [3-1:0] node3578;
	wire [3-1:0] node3582;
	wire [3-1:0] node3585;
	wire [3-1:0] node3586;
	wire [3-1:0] node3587;
	wire [3-1:0] node3591;
	wire [3-1:0] node3594;
	wire [3-1:0] node3595;
	wire [3-1:0] node3596;
	wire [3-1:0] node3597;
	wire [3-1:0] node3598;
	wire [3-1:0] node3599;
	wire [3-1:0] node3600;
	wire [3-1:0] node3604;
	wire [3-1:0] node3606;
	wire [3-1:0] node3609;
	wire [3-1:0] node3610;
	wire [3-1:0] node3611;
	wire [3-1:0] node3614;
	wire [3-1:0] node3617;
	wire [3-1:0] node3618;
	wire [3-1:0] node3620;
	wire [3-1:0] node3624;
	wire [3-1:0] node3625;
	wire [3-1:0] node3626;
	wire [3-1:0] node3627;
	wire [3-1:0] node3628;
	wire [3-1:0] node3633;
	wire [3-1:0] node3635;
	wire [3-1:0] node3638;
	wire [3-1:0] node3639;
	wire [3-1:0] node3641;
	wire [3-1:0] node3642;
	wire [3-1:0] node3645;
	wire [3-1:0] node3648;
	wire [3-1:0] node3650;
	wire [3-1:0] node3653;
	wire [3-1:0] node3654;
	wire [3-1:0] node3655;
	wire [3-1:0] node3656;
	wire [3-1:0] node3657;
	wire [3-1:0] node3658;
	wire [3-1:0] node3662;
	wire [3-1:0] node3664;
	wire [3-1:0] node3667;
	wire [3-1:0] node3668;
	wire [3-1:0] node3669;
	wire [3-1:0] node3672;
	wire [3-1:0] node3675;
	wire [3-1:0] node3677;
	wire [3-1:0] node3680;
	wire [3-1:0] node3681;
	wire [3-1:0] node3684;
	wire [3-1:0] node3685;
	wire [3-1:0] node3686;
	wire [3-1:0] node3689;
	wire [3-1:0] node3692;
	wire [3-1:0] node3695;
	wire [3-1:0] node3696;
	wire [3-1:0] node3697;
	wire [3-1:0] node3698;
	wire [3-1:0] node3701;
	wire [3-1:0] node3704;
	wire [3-1:0] node3705;
	wire [3-1:0] node3706;
	wire [3-1:0] node3709;
	wire [3-1:0] node3712;
	wire [3-1:0] node3713;
	wire [3-1:0] node3716;
	wire [3-1:0] node3719;
	wire [3-1:0] node3720;
	wire [3-1:0] node3721;
	wire [3-1:0] node3724;
	wire [3-1:0] node3727;
	wire [3-1:0] node3728;
	wire [3-1:0] node3729;
	wire [3-1:0] node3732;
	wire [3-1:0] node3735;
	wire [3-1:0] node3736;
	wire [3-1:0] node3739;
	wire [3-1:0] node3742;
	wire [3-1:0] node3743;
	wire [3-1:0] node3744;
	wire [3-1:0] node3745;
	wire [3-1:0] node3746;
	wire [3-1:0] node3749;
	wire [3-1:0] node3752;
	wire [3-1:0] node3753;
	wire [3-1:0] node3756;
	wire [3-1:0] node3759;
	wire [3-1:0] node3760;
	wire [3-1:0] node3761;
	wire [3-1:0] node3764;
	wire [3-1:0] node3767;
	wire [3-1:0] node3768;
	wire [3-1:0] node3771;
	wire [3-1:0] node3774;
	wire [3-1:0] node3775;
	wire [3-1:0] node3776;
	wire [3-1:0] node3777;
	wire [3-1:0] node3778;
	wire [3-1:0] node3781;
	wire [3-1:0] node3783;
	wire [3-1:0] node3786;
	wire [3-1:0] node3787;
	wire [3-1:0] node3791;
	wire [3-1:0] node3792;
	wire [3-1:0] node3793;
	wire [3-1:0] node3796;
	wire [3-1:0] node3799;
	wire [3-1:0] node3800;
	wire [3-1:0] node3803;
	wire [3-1:0] node3806;
	wire [3-1:0] node3807;
	wire [3-1:0] node3808;
	wire [3-1:0] node3811;
	wire [3-1:0] node3814;
	wire [3-1:0] node3815;
	wire [3-1:0] node3817;
	wire [3-1:0] node3820;
	wire [3-1:0] node3821;
	wire [3-1:0] node3824;

	assign outp = (inp[10]) ? node1832 : node1;
		assign node1 = (inp[6]) ? node933 : node2;
			assign node2 = (inp[11]) ? node554 : node3;
				assign node3 = (inp[1]) ? node275 : node4;
					assign node4 = (inp[0]) ? node138 : node5;
						assign node5 = (inp[8]) ? node71 : node6;
							assign node6 = (inp[4]) ? node28 : node7;
								assign node7 = (inp[5]) ? node15 : node8;
									assign node8 = (inp[9]) ? node12 : node9;
										assign node9 = (inp[7]) ? 3'b110 : 3'b111;
										assign node12 = (inp[7]) ? 3'b111 : 3'b110;
									assign node15 = (inp[3]) ? node23 : node16;
										assign node16 = (inp[2]) ? 3'b111 : node17;
											assign node17 = (inp[7]) ? node19 : 3'b110;
												assign node19 = (inp[9]) ? 3'b111 : 3'b110;
										assign node23 = (inp[9]) ? node25 : 3'b100;
											assign node25 = (inp[7]) ? 3'b101 : 3'b100;
								assign node28 = (inp[5]) ? node52 : node29;
									assign node29 = (inp[2]) ? node39 : node30;
										assign node30 = (inp[3]) ? node32 : 3'b100;
											assign node32 = (inp[7]) ? node36 : node33;
												assign node33 = (inp[9]) ? 3'b100 : 3'b101;
												assign node36 = (inp[9]) ? 3'b101 : 3'b100;
										assign node39 = (inp[3]) ? node47 : node40;
											assign node40 = (inp[9]) ? node44 : node41;
												assign node41 = (inp[7]) ? 3'b100 : 3'b101;
												assign node44 = (inp[7]) ? 3'b101 : 3'b100;
											assign node47 = (inp[9]) ? 3'b101 : node48;
												assign node48 = (inp[7]) ? 3'b100 : 3'b101;
									assign node52 = (inp[3]) ? node64 : node53;
										assign node53 = (inp[2]) ? node59 : node54;
											assign node54 = (inp[7]) ? 3'b101 : node55;
												assign node55 = (inp[9]) ? 3'b100 : 3'b101;
											assign node59 = (inp[9]) ? 3'b101 : node60;
												assign node60 = (inp[7]) ? 3'b100 : 3'b101;
										assign node64 = (inp[7]) ? 3'b110 : node65;
											assign node65 = (inp[9]) ? node67 : 3'b111;
												assign node67 = (inp[2]) ? 3'b111 : 3'b110;
							assign node71 = (inp[4]) ? node105 : node72;
								assign node72 = (inp[5]) ? node88 : node73;
									assign node73 = (inp[3]) ? node81 : node74;
										assign node74 = (inp[9]) ? node78 : node75;
											assign node75 = (inp[7]) ? 3'b100 : 3'b101;
											assign node78 = (inp[7]) ? 3'b101 : 3'b100;
										assign node81 = (inp[7]) ? node85 : node82;
											assign node82 = (inp[9]) ? 3'b100 : 3'b101;
											assign node85 = (inp[9]) ? 3'b101 : 3'b100;
									assign node88 = (inp[3]) ? node96 : node89;
										assign node89 = (inp[9]) ? node93 : node90;
											assign node90 = (inp[7]) ? 3'b100 : 3'b101;
											assign node93 = (inp[7]) ? 3'b101 : 3'b100;
										assign node96 = (inp[2]) ? node98 : 3'b111;
											assign node98 = (inp[7]) ? node102 : node99;
												assign node99 = (inp[9]) ? 3'b111 : 3'b110;
												assign node102 = (inp[9]) ? 3'b110 : 3'b111;
								assign node105 = (inp[5]) ? node117 : node106;
									assign node106 = (inp[2]) ? node112 : node107;
										assign node107 = (inp[7]) ? 3'b111 : node108;
											assign node108 = (inp[9]) ? 3'b110 : 3'b111;
										assign node112 = (inp[7]) ? 3'b110 : node113;
											assign node113 = (inp[9]) ? 3'b111 : 3'b110;
									assign node117 = (inp[3]) ? node125 : node118;
										assign node118 = (inp[9]) ? node120 : 3'b111;
											assign node120 = (inp[7]) ? node122 : 3'b111;
												assign node122 = (inp[2]) ? 3'b110 : 3'b111;
										assign node125 = (inp[7]) ? node133 : node126;
											assign node126 = (inp[2]) ? node130 : node127;
												assign node127 = (inp[9]) ? 3'b100 : 3'b101;
												assign node130 = (inp[9]) ? 3'b101 : 3'b100;
											assign node133 = (inp[9]) ? 3'b101 : node134;
												assign node134 = (inp[2]) ? 3'b101 : 3'b100;
						assign node138 = (inp[4]) ? node206 : node139;
							assign node139 = (inp[8]) ? node181 : node140;
								assign node140 = (inp[3]) ? node166 : node141;
									assign node141 = (inp[5]) ? node151 : node142;
										assign node142 = (inp[2]) ? 3'b111 : node143;
											assign node143 = (inp[9]) ? node147 : node144;
												assign node144 = (inp[7]) ? 3'b110 : 3'b111;
												assign node147 = (inp[7]) ? 3'b111 : 3'b110;
										assign node151 = (inp[9]) ? node159 : node152;
											assign node152 = (inp[7]) ? node156 : node153;
												assign node153 = (inp[2]) ? 3'b110 : 3'b111;
												assign node156 = (inp[2]) ? 3'b111 : 3'b110;
											assign node159 = (inp[7]) ? node163 : node160;
												assign node160 = (inp[2]) ? 3'b111 : 3'b110;
												assign node163 = (inp[2]) ? 3'b110 : 3'b111;
									assign node166 = (inp[5]) ? node174 : node167;
										assign node167 = (inp[2]) ? 3'b110 : node168;
											assign node168 = (inp[7]) ? node170 : 3'b111;
												assign node170 = (inp[9]) ? 3'b111 : 3'b110;
										assign node174 = (inp[9]) ? 3'b100 : node175;
											assign node175 = (inp[7]) ? 3'b101 : node176;
												assign node176 = (inp[2]) ? 3'b100 : 3'b101;
								assign node181 = (inp[5]) ? node191 : node182;
									assign node182 = (inp[3]) ? node184 : 3'b100;
										assign node184 = (inp[7]) ? node186 : 3'b100;
											assign node186 = (inp[2]) ? node188 : 3'b100;
												assign node188 = (inp[9]) ? 3'b100 : 3'b101;
									assign node191 = (inp[3]) ? node199 : node192;
										assign node192 = (inp[2]) ? 3'b101 : node193;
											assign node193 = (inp[9]) ? node195 : 3'b100;
												assign node195 = (inp[7]) ? 3'b101 : 3'b100;
										assign node199 = (inp[7]) ? node203 : node200;
											assign node200 = (inp[9]) ? 3'b111 : 3'b110;
											assign node203 = (inp[9]) ? 3'b110 : 3'b111;
							assign node206 = (inp[8]) ? node242 : node207;
								assign node207 = (inp[3]) ? node229 : node208;
									assign node208 = (inp[5]) ? node222 : node209;
										assign node209 = (inp[7]) ? node215 : node210;
											assign node210 = (inp[9]) ? node212 : 3'b101;
												assign node212 = (inp[2]) ? 3'b101 : 3'b100;
											assign node215 = (inp[9]) ? node219 : node216;
												assign node216 = (inp[2]) ? 3'b101 : 3'b100;
												assign node219 = (inp[2]) ? 3'b100 : 3'b101;
										assign node222 = (inp[7]) ? node224 : 3'b100;
											assign node224 = (inp[2]) ? 3'b101 : node225;
												assign node225 = (inp[9]) ? 3'b101 : 3'b100;
									assign node229 = (inp[5]) ? node237 : node230;
										assign node230 = (inp[2]) ? 3'b101 : node231;
											assign node231 = (inp[9]) ? 3'b101 : node232;
												assign node232 = (inp[7]) ? 3'b100 : 3'b101;
										assign node237 = (inp[9]) ? 3'b111 : node238;
											assign node238 = (inp[7]) ? 3'b111 : 3'b110;
								assign node242 = (inp[3]) ? node262 : node243;
									assign node243 = (inp[2]) ? node255 : node244;
										assign node244 = (inp[5]) ? node250 : node245;
											assign node245 = (inp[7]) ? node247 : 3'b111;
												assign node247 = (inp[9]) ? 3'b110 : 3'b111;
											assign node250 = (inp[9]) ? 3'b111 : node251;
												assign node251 = (inp[7]) ? 3'b111 : 3'b110;
										assign node255 = (inp[9]) ? node259 : node256;
											assign node256 = (inp[7]) ? 3'b111 : 3'b110;
											assign node259 = (inp[7]) ? 3'b110 : 3'b111;
									assign node262 = (inp[5]) ? node270 : node263;
										assign node263 = (inp[2]) ? node265 : 3'b110;
											assign node265 = (inp[7]) ? node267 : 3'b111;
												assign node267 = (inp[9]) ? 3'b110 : 3'b111;
										assign node270 = (inp[9]) ? node272 : 3'b100;
											assign node272 = (inp[7]) ? 3'b100 : 3'b101;
					assign node275 = (inp[7]) ? node425 : node276;
						assign node276 = (inp[9]) ? node338 : node277;
							assign node277 = (inp[0]) ? node307 : node278;
								assign node278 = (inp[2]) ? node294 : node279;
									assign node279 = (inp[4]) ? node285 : node280;
										assign node280 = (inp[8]) ? 3'b001 : node281;
											assign node281 = (inp[5]) ? 3'b001 : 3'b011;
										assign node285 = (inp[3]) ? node287 : 3'b011;
											assign node287 = (inp[8]) ? node291 : node288;
												assign node288 = (inp[5]) ? 3'b011 : 3'b001;
												assign node291 = (inp[5]) ? 3'b001 : 3'b011;
									assign node294 = (inp[8]) ? node300 : node295;
										assign node295 = (inp[4]) ? 3'b001 : node296;
											assign node296 = (inp[5]) ? 3'b001 : 3'b011;
										assign node300 = (inp[4]) ? node304 : node301;
											assign node301 = (inp[5]) ? 3'b010 : 3'b001;
											assign node304 = (inp[3]) ? 3'b000 : 3'b010;
								assign node307 = (inp[2]) ? node323 : node308;
									assign node308 = (inp[3]) ? node316 : node309;
										assign node309 = (inp[4]) ? node313 : node310;
											assign node310 = (inp[8]) ? 3'b001 : 3'b011;
											assign node313 = (inp[8]) ? 3'b010 : 3'b001;
										assign node316 = (inp[5]) ? 3'b010 : node317;
											assign node317 = (inp[4]) ? node319 : 3'b001;
												assign node319 = (inp[8]) ? 3'b010 : 3'b001;
									assign node323 = (inp[3]) ? node329 : node324;
										assign node324 = (inp[8]) ? 3'b010 : node325;
											assign node325 = (inp[4]) ? 3'b000 : 3'b010;
										assign node329 = (inp[4]) ? node331 : 3'b000;
											assign node331 = (inp[5]) ? node335 : node332;
												assign node332 = (inp[8]) ? 3'b010 : 3'b000;
												assign node335 = (inp[8]) ? 3'b000 : 3'b010;
							assign node338 = (inp[2]) ? node380 : node339;
								assign node339 = (inp[0]) ? node363 : node340;
									assign node340 = (inp[3]) ? node348 : node341;
										assign node341 = (inp[8]) ? node345 : node342;
											assign node342 = (inp[4]) ? 3'b000 : 3'b010;
											assign node345 = (inp[5]) ? 3'b000 : 3'b010;
										assign node348 = (inp[8]) ? node356 : node349;
											assign node349 = (inp[5]) ? node353 : node350;
												assign node350 = (inp[4]) ? 3'b000 : 3'b010;
												assign node353 = (inp[4]) ? 3'b010 : 3'b000;
											assign node356 = (inp[4]) ? node360 : node357;
												assign node357 = (inp[5]) ? 3'b010 : 3'b000;
												assign node360 = (inp[5]) ? 3'b000 : 3'b010;
									assign node363 = (inp[8]) ? node371 : node364;
										assign node364 = (inp[3]) ? node368 : node365;
											assign node365 = (inp[4]) ? 3'b000 : 3'b010;
											assign node368 = (inp[4]) ? 3'b011 : 3'b000;
										assign node371 = (inp[4]) ? node377 : node372;
											assign node372 = (inp[5]) ? node374 : 3'b000;
												assign node374 = (inp[3]) ? 3'b011 : 3'b000;
											assign node377 = (inp[3]) ? 3'b001 : 3'b011;
								assign node380 = (inp[0]) ? node400 : node381;
									assign node381 = (inp[4]) ? node391 : node382;
										assign node382 = (inp[5]) ? node384 : 3'b000;
											assign node384 = (inp[8]) ? node388 : node385;
												assign node385 = (inp[3]) ? 3'b000 : 3'b010;
												assign node388 = (inp[3]) ? 3'b011 : 3'b000;
										assign node391 = (inp[8]) ? node397 : node392;
											assign node392 = (inp[3]) ? node394 : 3'b000;
												assign node394 = (inp[5]) ? 3'b011 : 3'b000;
											assign node397 = (inp[3]) ? 3'b001 : 3'b011;
									assign node400 = (inp[5]) ? node410 : node401;
										assign node401 = (inp[3]) ? node403 : 3'b001;
											assign node403 = (inp[4]) ? node407 : node404;
												assign node404 = (inp[8]) ? 3'b001 : 3'b011;
												assign node407 = (inp[8]) ? 3'b011 : 3'b001;
										assign node410 = (inp[3]) ? node418 : node411;
											assign node411 = (inp[8]) ? node415 : node412;
												assign node412 = (inp[4]) ? 3'b001 : 3'b011;
												assign node415 = (inp[4]) ? 3'b011 : 3'b001;
											assign node418 = (inp[4]) ? node422 : node419;
												assign node419 = (inp[8]) ? 3'b011 : 3'b001;
												assign node422 = (inp[8]) ? 3'b001 : 3'b011;
						assign node425 = (inp[9]) ? node489 : node426;
							assign node426 = (inp[0]) ? node452 : node427;
								assign node427 = (inp[4]) ? node439 : node428;
									assign node428 = (inp[8]) ? node434 : node429;
										assign node429 = (inp[5]) ? node431 : 3'b010;
											assign node431 = (inp[3]) ? 3'b000 : 3'b010;
										assign node434 = (inp[3]) ? node436 : 3'b000;
											assign node436 = (inp[5]) ? 3'b010 : 3'b000;
									assign node439 = (inp[2]) ? node445 : node440;
										assign node440 = (inp[8]) ? node442 : 3'b000;
											assign node442 = (inp[3]) ? 3'b000 : 3'b010;
										assign node445 = (inp[8]) ? node449 : node446;
											assign node446 = (inp[5]) ? 3'b011 : 3'b000;
											assign node449 = (inp[3]) ? 3'b001 : 3'b011;
								assign node452 = (inp[2]) ? node474 : node453;
									assign node453 = (inp[4]) ? node465 : node454;
										assign node454 = (inp[8]) ? node460 : node455;
											assign node455 = (inp[5]) ? node457 : 3'b010;
												assign node457 = (inp[3]) ? 3'b000 : 3'b010;
											assign node460 = (inp[5]) ? node462 : 3'b000;
												assign node462 = (inp[3]) ? 3'b011 : 3'b000;
										assign node465 = (inp[8]) ? node469 : node466;
											assign node466 = (inp[5]) ? 3'b011 : 3'b000;
											assign node469 = (inp[3]) ? node471 : 3'b011;
												assign node471 = (inp[5]) ? 3'b001 : 3'b011;
									assign node474 = (inp[8]) ? node482 : node475;
										assign node475 = (inp[3]) ? node477 : 3'b011;
											assign node477 = (inp[4]) ? 3'b011 : node478;
												assign node478 = (inp[5]) ? 3'b001 : 3'b011;
										assign node482 = (inp[5]) ? node486 : node483;
											assign node483 = (inp[4]) ? 3'b011 : 3'b001;
											assign node486 = (inp[4]) ? 3'b001 : 3'b011;
							assign node489 = (inp[2]) ? node515 : node490;
								assign node490 = (inp[8]) ? node504 : node491;
									assign node491 = (inp[4]) ? node497 : node492;
										assign node492 = (inp[5]) ? node494 : 3'b011;
											assign node494 = (inp[3]) ? 3'b001 : 3'b011;
										assign node497 = (inp[3]) ? node499 : 3'b001;
											assign node499 = (inp[5]) ? node501 : 3'b001;
												assign node501 = (inp[0]) ? 3'b010 : 3'b011;
									assign node504 = (inp[0]) ? node510 : node505;
										assign node505 = (inp[4]) ? 3'b011 : node506;
											assign node506 = (inp[5]) ? 3'b011 : 3'b001;
										assign node510 = (inp[3]) ? 3'b010 : node511;
											assign node511 = (inp[4]) ? 3'b010 : 3'b001;
								assign node515 = (inp[0]) ? node533 : node516;
									assign node516 = (inp[8]) ? node526 : node517;
										assign node517 = (inp[3]) ? node521 : node518;
											assign node518 = (inp[4]) ? 3'b001 : 3'b011;
											assign node521 = (inp[4]) ? 3'b010 : node522;
												assign node522 = (inp[5]) ? 3'b001 : 3'b011;
										assign node526 = (inp[5]) ? node530 : node527;
											assign node527 = (inp[4]) ? 3'b010 : 3'b001;
											assign node530 = (inp[4]) ? 3'b000 : 3'b010;
									assign node533 = (inp[8]) ? node543 : node534;
										assign node534 = (inp[3]) ? node536 : 3'b000;
											assign node536 = (inp[4]) ? node540 : node537;
												assign node537 = (inp[5]) ? 3'b000 : 3'b010;
												assign node540 = (inp[5]) ? 3'b010 : 3'b000;
										assign node543 = (inp[4]) ? node549 : node544;
											assign node544 = (inp[5]) ? node546 : 3'b000;
												assign node546 = (inp[3]) ? 3'b010 : 3'b000;
											assign node549 = (inp[5]) ? node551 : 3'b010;
												assign node551 = (inp[3]) ? 3'b000 : 3'b010;
				assign node554 = (inp[3]) ? node664 : node555;
					assign node555 = (inp[7]) ? node607 : node556;
						assign node556 = (inp[9]) ? node582 : node557;
							assign node557 = (inp[0]) ? node567 : node558;
								assign node558 = (inp[8]) ? node562 : node559;
									assign node559 = (inp[4]) ? 3'b001 : 3'b011;
									assign node562 = (inp[4]) ? node564 : 3'b001;
										assign node564 = (inp[2]) ? 3'b010 : 3'b011;
								assign node567 = (inp[2]) ? node575 : node568;
									assign node568 = (inp[8]) ? node572 : node569;
										assign node569 = (inp[4]) ? 3'b001 : 3'b011;
										assign node572 = (inp[4]) ? 3'b010 : 3'b001;
									assign node575 = (inp[8]) ? node579 : node576;
										assign node576 = (inp[4]) ? 3'b000 : 3'b010;
										assign node579 = (inp[4]) ? 3'b010 : 3'b000;
							assign node582 = (inp[0]) ? node592 : node583;
								assign node583 = (inp[4]) ? node587 : node584;
									assign node584 = (inp[8]) ? 3'b000 : 3'b010;
									assign node587 = (inp[8]) ? node589 : 3'b000;
										assign node589 = (inp[2]) ? 3'b011 : 3'b010;
								assign node592 = (inp[2]) ? node600 : node593;
									assign node593 = (inp[4]) ? node597 : node594;
										assign node594 = (inp[8]) ? 3'b000 : 3'b010;
										assign node597 = (inp[8]) ? 3'b011 : 3'b000;
									assign node600 = (inp[8]) ? node604 : node601;
										assign node601 = (inp[4]) ? 3'b001 : 3'b011;
										assign node604 = (inp[4]) ? 3'b011 : 3'b001;
						assign node607 = (inp[9]) ? node639 : node608;
							assign node608 = (inp[0]) ? node624 : node609;
								assign node609 = (inp[2]) ? node617 : node610;
									assign node610 = (inp[8]) ? node614 : node611;
										assign node611 = (inp[4]) ? 3'b000 : 3'b010;
										assign node614 = (inp[4]) ? 3'b010 : 3'b000;
									assign node617 = (inp[4]) ? node621 : node618;
										assign node618 = (inp[8]) ? 3'b000 : 3'b010;
										assign node621 = (inp[8]) ? 3'b011 : 3'b000;
								assign node624 = (inp[2]) ? node632 : node625;
									assign node625 = (inp[8]) ? node629 : node626;
										assign node626 = (inp[4]) ? 3'b000 : 3'b010;
										assign node629 = (inp[4]) ? 3'b011 : 3'b000;
									assign node632 = (inp[8]) ? node636 : node633;
										assign node633 = (inp[4]) ? 3'b001 : 3'b011;
										assign node636 = (inp[4]) ? 3'b011 : 3'b001;
							assign node639 = (inp[0]) ? node649 : node640;
								assign node640 = (inp[8]) ? node644 : node641;
									assign node641 = (inp[4]) ? 3'b001 : 3'b011;
									assign node644 = (inp[4]) ? node646 : 3'b001;
										assign node646 = (inp[2]) ? 3'b010 : 3'b011;
								assign node649 = (inp[2]) ? node657 : node650;
									assign node650 = (inp[4]) ? node654 : node651;
										assign node651 = (inp[8]) ? 3'b001 : 3'b011;
										assign node654 = (inp[8]) ? 3'b010 : 3'b001;
									assign node657 = (inp[8]) ? node661 : node658;
										assign node658 = (inp[4]) ? 3'b000 : 3'b010;
										assign node661 = (inp[4]) ? 3'b010 : 3'b000;
					assign node664 = (inp[8]) ? node776 : node665;
						assign node665 = (inp[7]) ? node723 : node666;
							assign node666 = (inp[9]) ? node702 : node667;
								assign node667 = (inp[0]) ? node689 : node668;
									assign node668 = (inp[1]) ? node678 : node669;
										assign node669 = (inp[5]) ? node673 : node670;
											assign node670 = (inp[4]) ? 3'b001 : 3'b011;
											assign node673 = (inp[4]) ? node675 : 3'b001;
												assign node675 = (inp[2]) ? 3'b010 : 3'b011;
										assign node678 = (inp[2]) ? node684 : node679;
											assign node679 = (inp[4]) ? node681 : 3'b001;
												assign node681 = (inp[5]) ? 3'b011 : 3'b001;
											assign node684 = (inp[4]) ? 3'b001 : node685;
												assign node685 = (inp[5]) ? 3'b001 : 3'b011;
									assign node689 = (inp[2]) ? node697 : node690;
										assign node690 = (inp[4]) ? node694 : node691;
											assign node691 = (inp[5]) ? 3'b001 : 3'b011;
											assign node694 = (inp[5]) ? 3'b010 : 3'b001;
										assign node697 = (inp[4]) ? node699 : 3'b000;
											assign node699 = (inp[5]) ? 3'b010 : 3'b000;
								assign node702 = (inp[2]) ? node708 : node703;
									assign node703 = (inp[5]) ? 3'b000 : node704;
										assign node704 = (inp[4]) ? 3'b000 : 3'b010;
									assign node708 = (inp[0]) ? node716 : node709;
										assign node709 = (inp[5]) ? node713 : node710;
											assign node710 = (inp[4]) ? 3'b000 : 3'b010;
											assign node713 = (inp[4]) ? 3'b011 : 3'b000;
										assign node716 = (inp[4]) ? node720 : node717;
											assign node717 = (inp[5]) ? 3'b001 : 3'b011;
											assign node720 = (inp[5]) ? 3'b011 : 3'b001;
							assign node723 = (inp[9]) ? node751 : node724;
								assign node724 = (inp[0]) ? node738 : node725;
									assign node725 = (inp[2]) ? node733 : node726;
										assign node726 = (inp[5]) ? node730 : node727;
											assign node727 = (inp[4]) ? 3'b000 : 3'b010;
											assign node730 = (inp[4]) ? 3'b010 : 3'b000;
										assign node733 = (inp[4]) ? 3'b011 : node734;
											assign node734 = (inp[5]) ? 3'b000 : 3'b010;
									assign node738 = (inp[2]) ? node746 : node739;
										assign node739 = (inp[4]) ? node743 : node740;
											assign node740 = (inp[5]) ? 3'b000 : 3'b010;
											assign node743 = (inp[5]) ? 3'b011 : 3'b000;
										assign node746 = (inp[4]) ? node748 : 3'b011;
											assign node748 = (inp[5]) ? 3'b011 : 3'b001;
								assign node751 = (inp[0]) ? node761 : node752;
									assign node752 = (inp[5]) ? node756 : node753;
										assign node753 = (inp[4]) ? 3'b001 : 3'b011;
										assign node756 = (inp[4]) ? node758 : 3'b001;
											assign node758 = (inp[2]) ? 3'b010 : 3'b011;
									assign node761 = (inp[2]) ? node769 : node762;
										assign node762 = (inp[5]) ? node766 : node763;
											assign node763 = (inp[4]) ? 3'b001 : 3'b011;
											assign node766 = (inp[4]) ? 3'b010 : 3'b001;
										assign node769 = (inp[4]) ? node773 : node770;
											assign node770 = (inp[5]) ? 3'b000 : 3'b010;
											assign node773 = (inp[5]) ? 3'b010 : 3'b000;
						assign node776 = (inp[1]) ? node872 : node777;
							assign node777 = (inp[0]) ? node831 : node778;
								assign node778 = (inp[7]) ? node800 : node779;
									assign node779 = (inp[5]) ? node785 : node780;
										assign node780 = (inp[4]) ? 3'b011 : node781;
											assign node781 = (inp[9]) ? 3'b000 : 3'b001;
										assign node785 = (inp[4]) ? node793 : node786;
											assign node786 = (inp[2]) ? node790 : node787;
												assign node787 = (inp[9]) ? 3'b010 : 3'b011;
												assign node790 = (inp[9]) ? 3'b011 : 3'b010;
											assign node793 = (inp[2]) ? node797 : node794;
												assign node794 = (inp[9]) ? 3'b000 : 3'b001;
												assign node797 = (inp[9]) ? 3'b001 : 3'b000;
									assign node800 = (inp[9]) ? node816 : node801;
										assign node801 = (inp[2]) ? node809 : node802;
											assign node802 = (inp[5]) ? node806 : node803;
												assign node803 = (inp[4]) ? 3'b010 : 3'b000;
												assign node806 = (inp[4]) ? 3'b000 : 3'b010;
											assign node809 = (inp[4]) ? node813 : node810;
												assign node810 = (inp[5]) ? 3'b011 : 3'b000;
												assign node813 = (inp[5]) ? 3'b001 : 3'b011;
										assign node816 = (inp[2]) ? node824 : node817;
											assign node817 = (inp[4]) ? node821 : node818;
												assign node818 = (inp[5]) ? 3'b011 : 3'b001;
												assign node821 = (inp[5]) ? 3'b001 : 3'b011;
											assign node824 = (inp[5]) ? node828 : node825;
												assign node825 = (inp[4]) ? 3'b010 : 3'b001;
												assign node828 = (inp[4]) ? 3'b000 : 3'b010;
								assign node831 = (inp[4]) ? node853 : node832;
									assign node832 = (inp[5]) ? node840 : node833;
										assign node833 = (inp[2]) ? node837 : node834;
											assign node834 = (inp[7]) ? 3'b001 : 3'b000;
											assign node837 = (inp[7]) ? 3'b000 : 3'b001;
										assign node840 = (inp[2]) ? node846 : node841;
											assign node841 = (inp[7]) ? 3'b010 : node842;
												assign node842 = (inp[9]) ? 3'b011 : 3'b010;
											assign node846 = (inp[7]) ? node850 : node847;
												assign node847 = (inp[9]) ? 3'b011 : 3'b010;
												assign node850 = (inp[9]) ? 3'b010 : 3'b011;
									assign node853 = (inp[5]) ? node861 : node854;
										assign node854 = (inp[9]) ? node858 : node855;
											assign node855 = (inp[7]) ? 3'b011 : 3'b010;
											assign node858 = (inp[7]) ? 3'b010 : 3'b011;
										assign node861 = (inp[2]) ? node867 : node862;
											assign node862 = (inp[9]) ? 3'b000 : node863;
												assign node863 = (inp[7]) ? 3'b001 : 3'b000;
											assign node867 = (inp[7]) ? 3'b001 : node868;
												assign node868 = (inp[9]) ? 3'b001 : 3'b000;
							assign node872 = (inp[5]) ? node902 : node873;
								assign node873 = (inp[4]) ? node883 : node874;
									assign node874 = (inp[9]) ? 3'b001 : node875;
										assign node875 = (inp[0]) ? node877 : 3'b000;
											assign node877 = (inp[2]) ? 3'b001 : node878;
												assign node878 = (inp[7]) ? 3'b000 : 3'b001;
									assign node883 = (inp[7]) ? node891 : node884;
										assign node884 = (inp[9]) ? 3'b011 : node885;
											assign node885 = (inp[2]) ? 3'b010 : node886;
												assign node886 = (inp[0]) ? 3'b010 : 3'b011;
										assign node891 = (inp[9]) ? node897 : node892;
											assign node892 = (inp[0]) ? 3'b011 : node893;
												assign node893 = (inp[2]) ? 3'b011 : 3'b010;
											assign node897 = (inp[0]) ? 3'b010 : node898;
												assign node898 = (inp[2]) ? 3'b010 : 3'b011;
								assign node902 = (inp[4]) ? node918 : node903;
									assign node903 = (inp[7]) ? node913 : node904;
										assign node904 = (inp[9]) ? node908 : node905;
											assign node905 = (inp[2]) ? 3'b010 : 3'b011;
											assign node908 = (inp[0]) ? 3'b011 : node909;
												assign node909 = (inp[2]) ? 3'b011 : 3'b010;
										assign node913 = (inp[9]) ? node915 : 3'b011;
											assign node915 = (inp[0]) ? 3'b010 : 3'b011;
									assign node918 = (inp[0]) ? node926 : node919;
										assign node919 = (inp[9]) ? node921 : 3'b001;
											assign node921 = (inp[7]) ? 3'b000 : node922;
												assign node922 = (inp[2]) ? 3'b001 : 3'b000;
										assign node926 = (inp[9]) ? node930 : node927;
											assign node927 = (inp[7]) ? 3'b001 : 3'b000;
											assign node930 = (inp[7]) ? 3'b000 : 3'b001;
			assign node933 = (inp[1]) ? node1437 : node934;
				assign node934 = (inp[11]) ? node1214 : node935;
					assign node935 = (inp[9]) ? node1091 : node936;
						assign node936 = (inp[7]) ? node1010 : node937;
							assign node937 = (inp[2]) ? node967 : node938;
								assign node938 = (inp[0]) ? node954 : node939;
									assign node939 = (inp[5]) ? node947 : node940;
										assign node940 = (inp[8]) ? node944 : node941;
											assign node941 = (inp[4]) ? 3'b001 : 3'b011;
											assign node944 = (inp[4]) ? 3'b011 : 3'b001;
										assign node947 = (inp[3]) ? 3'b001 : node948;
											assign node948 = (inp[8]) ? node950 : 3'b001;
												assign node950 = (inp[4]) ? 3'b011 : 3'b001;
									assign node954 = (inp[4]) ? node958 : node955;
										assign node955 = (inp[8]) ? 3'b001 : 3'b011;
										assign node958 = (inp[8]) ? node964 : node959;
											assign node959 = (inp[3]) ? node961 : 3'b001;
												assign node961 = (inp[5]) ? 3'b010 : 3'b001;
											assign node964 = (inp[3]) ? 3'b000 : 3'b010;
								assign node967 = (inp[0]) ? node991 : node968;
									assign node968 = (inp[8]) ? node980 : node969;
										assign node969 = (inp[4]) ? node975 : node970;
											assign node970 = (inp[5]) ? node972 : 3'b011;
												assign node972 = (inp[3]) ? 3'b001 : 3'b011;
											assign node975 = (inp[3]) ? node977 : 3'b001;
												assign node977 = (inp[5]) ? 3'b010 : 3'b001;
										assign node980 = (inp[4]) ? node986 : node981;
											assign node981 = (inp[3]) ? node983 : 3'b001;
												assign node983 = (inp[5]) ? 3'b010 : 3'b001;
											assign node986 = (inp[5]) ? node988 : 3'b010;
												assign node988 = (inp[3]) ? 3'b000 : 3'b010;
									assign node991 = (inp[8]) ? node1001 : node992;
										assign node992 = (inp[3]) ? node994 : 3'b000;
											assign node994 = (inp[5]) ? node998 : node995;
												assign node995 = (inp[4]) ? 3'b000 : 3'b010;
												assign node998 = (inp[4]) ? 3'b010 : 3'b000;
										assign node1001 = (inp[4]) ? node1005 : node1002;
											assign node1002 = (inp[5]) ? 3'b010 : 3'b000;
											assign node1005 = (inp[5]) ? node1007 : 3'b010;
												assign node1007 = (inp[3]) ? 3'b000 : 3'b010;
							assign node1010 = (inp[2]) ? node1048 : node1011;
								assign node1011 = (inp[0]) ? node1029 : node1012;
									assign node1012 = (inp[5]) ? node1020 : node1013;
										assign node1013 = (inp[4]) ? node1017 : node1014;
											assign node1014 = (inp[8]) ? 3'b000 : 3'b010;
											assign node1017 = (inp[8]) ? 3'b010 : 3'b000;
										assign node1020 = (inp[8]) ? node1022 : 3'b010;
											assign node1022 = (inp[3]) ? node1026 : node1023;
												assign node1023 = (inp[4]) ? 3'b010 : 3'b000;
												assign node1026 = (inp[4]) ? 3'b000 : 3'b010;
									assign node1029 = (inp[8]) ? node1037 : node1030;
										assign node1030 = (inp[4]) ? 3'b000 : node1031;
											assign node1031 = (inp[5]) ? node1033 : 3'b010;
												assign node1033 = (inp[3]) ? 3'b000 : 3'b010;
										assign node1037 = (inp[4]) ? node1043 : node1038;
											assign node1038 = (inp[3]) ? node1040 : 3'b000;
												assign node1040 = (inp[5]) ? 3'b011 : 3'b000;
											assign node1043 = (inp[5]) ? node1045 : 3'b011;
												assign node1045 = (inp[3]) ? 3'b001 : 3'b011;
								assign node1048 = (inp[0]) ? node1070 : node1049;
									assign node1049 = (inp[4]) ? node1061 : node1050;
										assign node1050 = (inp[8]) ? node1056 : node1051;
											assign node1051 = (inp[3]) ? node1053 : 3'b010;
												assign node1053 = (inp[5]) ? 3'b000 : 3'b010;
											assign node1056 = (inp[5]) ? node1058 : 3'b000;
												assign node1058 = (inp[3]) ? 3'b011 : 3'b000;
										assign node1061 = (inp[8]) ? node1065 : node1062;
											assign node1062 = (inp[5]) ? 3'b011 : 3'b000;
											assign node1065 = (inp[3]) ? node1067 : 3'b011;
												assign node1067 = (inp[5]) ? 3'b001 : 3'b011;
									assign node1070 = (inp[5]) ? node1084 : node1071;
										assign node1071 = (inp[3]) ? node1079 : node1072;
											assign node1072 = (inp[8]) ? node1076 : node1073;
												assign node1073 = (inp[4]) ? 3'b001 : 3'b011;
												assign node1076 = (inp[4]) ? 3'b011 : 3'b001;
											assign node1079 = (inp[4]) ? node1081 : 3'b001;
												assign node1081 = (inp[8]) ? 3'b011 : 3'b001;
										assign node1084 = (inp[3]) ? node1086 : 3'b001;
											assign node1086 = (inp[8]) ? node1088 : 3'b001;
												assign node1088 = (inp[4]) ? 3'b001 : 3'b011;
						assign node1091 = (inp[7]) ? node1159 : node1092;
							assign node1092 = (inp[2]) ? node1118 : node1093;
								assign node1093 = (inp[8]) ? node1105 : node1094;
									assign node1094 = (inp[4]) ? node1100 : node1095;
										assign node1095 = (inp[5]) ? node1097 : 3'b010;
											assign node1097 = (inp[0]) ? 3'b010 : 3'b000;
										assign node1100 = (inp[5]) ? node1102 : 3'b000;
											assign node1102 = (inp[3]) ? 3'b010 : 3'b000;
									assign node1105 = (inp[4]) ? node1113 : node1106;
										assign node1106 = (inp[3]) ? node1108 : 3'b000;
											assign node1108 = (inp[5]) ? node1110 : 3'b000;
												assign node1110 = (inp[0]) ? 3'b011 : 3'b010;
										assign node1113 = (inp[0]) ? node1115 : 3'b010;
											assign node1115 = (inp[5]) ? 3'b001 : 3'b011;
								assign node1118 = (inp[0]) ? node1136 : node1119;
									assign node1119 = (inp[8]) ? node1125 : node1120;
										assign node1120 = (inp[4]) ? 3'b000 : node1121;
											assign node1121 = (inp[5]) ? 3'b000 : 3'b010;
										assign node1125 = (inp[4]) ? node1131 : node1126;
											assign node1126 = (inp[5]) ? node1128 : 3'b000;
												assign node1128 = (inp[3]) ? 3'b011 : 3'b000;
											assign node1131 = (inp[5]) ? node1133 : 3'b011;
												assign node1133 = (inp[3]) ? 3'b001 : 3'b011;
									assign node1136 = (inp[3]) ? node1144 : node1137;
										assign node1137 = (inp[8]) ? node1141 : node1138;
											assign node1138 = (inp[5]) ? 3'b011 : 3'b001;
											assign node1141 = (inp[4]) ? 3'b011 : 3'b001;
										assign node1144 = (inp[5]) ? node1152 : node1145;
											assign node1145 = (inp[8]) ? node1149 : node1146;
												assign node1146 = (inp[4]) ? 3'b001 : 3'b011;
												assign node1149 = (inp[4]) ? 3'b011 : 3'b001;
											assign node1152 = (inp[4]) ? node1156 : node1153;
												assign node1153 = (inp[8]) ? 3'b011 : 3'b001;
												assign node1156 = (inp[8]) ? 3'b001 : 3'b011;
							assign node1159 = (inp[2]) ? node1181 : node1160;
								assign node1160 = (inp[4]) ? node1172 : node1161;
									assign node1161 = (inp[8]) ? node1167 : node1162;
										assign node1162 = (inp[5]) ? node1164 : 3'b011;
											assign node1164 = (inp[3]) ? 3'b001 : 3'b011;
										assign node1167 = (inp[5]) ? node1169 : 3'b001;
											assign node1169 = (inp[3]) ? 3'b011 : 3'b001;
									assign node1172 = (inp[8]) ? node1174 : 3'b001;
										assign node1174 = (inp[0]) ? node1178 : node1175;
											assign node1175 = (inp[3]) ? 3'b001 : 3'b011;
											assign node1178 = (inp[3]) ? 3'b000 : 3'b010;
								assign node1181 = (inp[0]) ? node1199 : node1182;
									assign node1182 = (inp[5]) ? node1188 : node1183;
										assign node1183 = (inp[4]) ? 3'b001 : node1184;
											assign node1184 = (inp[8]) ? 3'b001 : 3'b011;
										assign node1188 = (inp[4]) ? node1192 : node1189;
											assign node1189 = (inp[8]) ? 3'b001 : 3'b011;
											assign node1192 = (inp[8]) ? node1196 : node1193;
												assign node1193 = (inp[3]) ? 3'b010 : 3'b001;
												assign node1196 = (inp[3]) ? 3'b000 : 3'b010;
									assign node1199 = (inp[3]) ? node1207 : node1200;
										assign node1200 = (inp[5]) ? node1202 : 3'b010;
											assign node1202 = (inp[4]) ? node1204 : 3'b000;
												assign node1204 = (inp[8]) ? 3'b010 : 3'b000;
										assign node1207 = (inp[4]) ? 3'b000 : node1208;
											assign node1208 = (inp[8]) ? 3'b000 : node1209;
												assign node1209 = (inp[5]) ? 3'b000 : 3'b010;
					assign node1214 = (inp[9]) ? node1324 : node1215;
						assign node1215 = (inp[7]) ? node1277 : node1216;
							assign node1216 = (inp[0]) ? node1244 : node1217;
								assign node1217 = (inp[2]) ? node1231 : node1218;
									assign node1218 = (inp[8]) ? node1224 : node1219;
										assign node1219 = (inp[4]) ? 3'b111 : node1220;
											assign node1220 = (inp[5]) ? 3'b101 : 3'b111;
										assign node1224 = (inp[4]) ? 3'b101 : node1225;
											assign node1225 = (inp[3]) ? 3'b111 : node1226;
												assign node1226 = (inp[5]) ? 3'b111 : 3'b101;
									assign node1231 = (inp[4]) ? 3'b110 : node1232;
										assign node1232 = (inp[8]) ? node1238 : node1233;
											assign node1233 = (inp[5]) ? 3'b101 : node1234;
												assign node1234 = (inp[3]) ? 3'b101 : 3'b111;
											assign node1238 = (inp[5]) ? 3'b110 : node1239;
												assign node1239 = (inp[3]) ? 3'b110 : 3'b101;
								assign node1244 = (inp[2]) ? node1258 : node1245;
									assign node1245 = (inp[4]) ? node1251 : node1246;
										assign node1246 = (inp[8]) ? node1248 : 3'b101;
											assign node1248 = (inp[3]) ? 3'b110 : 3'b101;
										assign node1251 = (inp[8]) ? 3'b100 : node1252;
											assign node1252 = (inp[3]) ? 3'b110 : node1253;
												assign node1253 = (inp[5]) ? 3'b110 : 3'b101;
									assign node1258 = (inp[4]) ? node1270 : node1259;
										assign node1259 = (inp[8]) ? node1265 : node1260;
											assign node1260 = (inp[3]) ? 3'b100 : node1261;
												assign node1261 = (inp[5]) ? 3'b100 : 3'b110;
											assign node1265 = (inp[5]) ? 3'b110 : node1266;
												assign node1266 = (inp[3]) ? 3'b110 : 3'b100;
										assign node1270 = (inp[8]) ? 3'b100 : node1271;
											assign node1271 = (inp[5]) ? 3'b110 : node1272;
												assign node1272 = (inp[3]) ? 3'b110 : 3'b100;
							assign node1277 = (inp[0]) ? node1303 : node1278;
								assign node1278 = (inp[4]) ? node1292 : node1279;
									assign node1279 = (inp[2]) ? node1285 : node1280;
										assign node1280 = (inp[8]) ? 3'b110 : node1281;
											assign node1281 = (inp[3]) ? 3'b100 : 3'b110;
										assign node1285 = (inp[3]) ? 3'b100 : node1286;
											assign node1286 = (inp[8]) ? 3'b100 : node1287;
												assign node1287 = (inp[5]) ? 3'b100 : 3'b110;
									assign node1292 = (inp[2]) ? node1298 : node1293;
										assign node1293 = (inp[3]) ? node1295 : 3'b110;
											assign node1295 = (inp[8]) ? 3'b100 : 3'b110;
										assign node1298 = (inp[8]) ? node1300 : 3'b111;
											assign node1300 = (inp[5]) ? 3'b101 : 3'b111;
								assign node1303 = (inp[8]) ? node1315 : node1304;
									assign node1304 = (inp[4]) ? node1310 : node1305;
										assign node1305 = (inp[2]) ? node1307 : 3'b100;
											assign node1307 = (inp[3]) ? 3'b101 : 3'b111;
										assign node1310 = (inp[3]) ? 3'b111 : node1311;
											assign node1311 = (inp[5]) ? 3'b111 : 3'b101;
									assign node1315 = (inp[4]) ? node1321 : node1316;
										assign node1316 = (inp[3]) ? 3'b111 : node1317;
											assign node1317 = (inp[5]) ? 3'b111 : 3'b101;
										assign node1321 = (inp[3]) ? 3'b101 : 3'b111;
						assign node1324 = (inp[4]) ? node1382 : node1325;
							assign node1325 = (inp[8]) ? node1357 : node1326;
								assign node1326 = (inp[3]) ? node1346 : node1327;
									assign node1327 = (inp[5]) ? node1339 : node1328;
										assign node1328 = (inp[7]) ? node1334 : node1329;
											assign node1329 = (inp[2]) ? node1331 : 3'b110;
												assign node1331 = (inp[0]) ? 3'b111 : 3'b110;
											assign node1334 = (inp[0]) ? node1336 : 3'b111;
												assign node1336 = (inp[2]) ? 3'b110 : 3'b111;
										assign node1339 = (inp[7]) ? node1341 : 3'b100;
											assign node1341 = (inp[0]) ? node1343 : 3'b101;
												assign node1343 = (inp[2]) ? 3'b100 : 3'b101;
									assign node1346 = (inp[7]) ? node1352 : node1347;
										assign node1347 = (inp[2]) ? node1349 : 3'b100;
											assign node1349 = (inp[0]) ? 3'b101 : 3'b100;
										assign node1352 = (inp[0]) ? node1354 : 3'b101;
											assign node1354 = (inp[2]) ? 3'b100 : 3'b101;
								assign node1357 = (inp[3]) ? node1371 : node1358;
									assign node1358 = (inp[5]) ? node1366 : node1359;
										assign node1359 = (inp[7]) ? 3'b101 : node1360;
											assign node1360 = (inp[0]) ? node1362 : 3'b100;
												assign node1362 = (inp[2]) ? 3'b101 : 3'b100;
										assign node1366 = (inp[7]) ? node1368 : 3'b111;
											assign node1368 = (inp[0]) ? 3'b110 : 3'b111;
									assign node1371 = (inp[7]) ? node1377 : node1372;
										assign node1372 = (inp[0]) ? 3'b111 : node1373;
											assign node1373 = (inp[2]) ? 3'b111 : 3'b110;
										assign node1377 = (inp[2]) ? 3'b110 : node1378;
											assign node1378 = (inp[0]) ? 3'b110 : 3'b111;
							assign node1382 = (inp[8]) ? node1408 : node1383;
								assign node1383 = (inp[5]) ? node1399 : node1384;
									assign node1384 = (inp[3]) ? node1390 : node1385;
										assign node1385 = (inp[7]) ? node1387 : 3'b100;
											assign node1387 = (inp[2]) ? 3'b100 : 3'b101;
										assign node1390 = (inp[0]) ? 3'b110 : node1391;
											assign node1391 = (inp[7]) ? node1395 : node1392;
												assign node1392 = (inp[2]) ? 3'b111 : 3'b110;
												assign node1395 = (inp[2]) ? 3'b110 : 3'b111;
									assign node1399 = (inp[7]) ? node1405 : node1400;
										assign node1400 = (inp[2]) ? 3'b111 : node1401;
											assign node1401 = (inp[0]) ? 3'b111 : 3'b110;
										assign node1405 = (inp[2]) ? 3'b110 : 3'b111;
								assign node1408 = (inp[3]) ? node1426 : node1409;
									assign node1409 = (inp[5]) ? node1419 : node1410;
										assign node1410 = (inp[7]) ? node1414 : node1411;
											assign node1411 = (inp[0]) ? 3'b111 : 3'b110;
											assign node1414 = (inp[0]) ? 3'b110 : node1415;
												assign node1415 = (inp[2]) ? 3'b110 : 3'b111;
										assign node1419 = (inp[7]) ? node1421 : 3'b101;
											assign node1421 = (inp[0]) ? 3'b100 : node1422;
												assign node1422 = (inp[2]) ? 3'b100 : 3'b101;
									assign node1426 = (inp[7]) ? node1432 : node1427;
										assign node1427 = (inp[2]) ? 3'b101 : node1428;
											assign node1428 = (inp[0]) ? 3'b101 : 3'b100;
										assign node1432 = (inp[2]) ? 3'b100 : node1433;
											assign node1433 = (inp[0]) ? 3'b100 : 3'b101;
				assign node1437 = (inp[9]) ? node1623 : node1438;
					assign node1438 = (inp[7]) ? node1532 : node1439;
						assign node1439 = (inp[2]) ? node1489 : node1440;
							assign node1440 = (inp[0]) ? node1466 : node1441;
								assign node1441 = (inp[11]) ? node1455 : node1442;
									assign node1442 = (inp[8]) ? 3'b111 : node1443;
										assign node1443 = (inp[4]) ? node1449 : node1444;
											assign node1444 = (inp[5]) ? 3'b101 : node1445;
												assign node1445 = (inp[3]) ? 3'b101 : 3'b111;
											assign node1449 = (inp[3]) ? 3'b111 : node1450;
												assign node1450 = (inp[5]) ? 3'b111 : 3'b101;
									assign node1455 = (inp[4]) ? node1459 : node1456;
										assign node1456 = (inp[8]) ? 3'b111 : 3'b101;
										assign node1459 = (inp[8]) ? node1461 : 3'b111;
											assign node1461 = (inp[5]) ? 3'b101 : node1462;
												assign node1462 = (inp[3]) ? 3'b101 : 3'b111;
								assign node1466 = (inp[4]) ? node1478 : node1467;
									assign node1467 = (inp[8]) ? node1473 : node1468;
										assign node1468 = (inp[3]) ? 3'b101 : node1469;
											assign node1469 = (inp[5]) ? 3'b101 : 3'b111;
										assign node1473 = (inp[3]) ? 3'b110 : node1474;
											assign node1474 = (inp[5]) ? 3'b110 : 3'b101;
									assign node1478 = (inp[8]) ? node1484 : node1479;
										assign node1479 = (inp[3]) ? 3'b110 : node1480;
											assign node1480 = (inp[5]) ? 3'b110 : 3'b101;
										assign node1484 = (inp[3]) ? 3'b100 : node1485;
											assign node1485 = (inp[5]) ? 3'b100 : 3'b110;
							assign node1489 = (inp[0]) ? node1509 : node1490;
								assign node1490 = (inp[4]) ? node1498 : node1491;
									assign node1491 = (inp[8]) ? node1493 : 3'b101;
										assign node1493 = (inp[3]) ? 3'b110 : node1494;
											assign node1494 = (inp[11]) ? 3'b110 : 3'b101;
									assign node1498 = (inp[8]) ? node1504 : node1499;
										assign node1499 = (inp[3]) ? 3'b110 : node1500;
											assign node1500 = (inp[5]) ? 3'b110 : 3'b101;
										assign node1504 = (inp[5]) ? 3'b100 : node1505;
											assign node1505 = (inp[3]) ? 3'b100 : 3'b110;
								assign node1509 = (inp[3]) ? node1525 : node1510;
									assign node1510 = (inp[8]) ? node1520 : node1511;
										assign node1511 = (inp[11]) ? node1517 : node1512;
											assign node1512 = (inp[5]) ? node1514 : 3'b100;
												assign node1514 = (inp[4]) ? 3'b110 : 3'b100;
											assign node1517 = (inp[4]) ? 3'b100 : 3'b110;
										assign node1520 = (inp[4]) ? node1522 : 3'b100;
											assign node1522 = (inp[5]) ? 3'b100 : 3'b110;
									assign node1525 = (inp[4]) ? node1529 : node1526;
										assign node1526 = (inp[8]) ? 3'b110 : 3'b100;
										assign node1529 = (inp[8]) ? 3'b100 : 3'b110;
						assign node1532 = (inp[2]) ? node1578 : node1533;
							assign node1533 = (inp[0]) ? node1557 : node1534;
								assign node1534 = (inp[4]) ? node1546 : node1535;
									assign node1535 = (inp[8]) ? node1541 : node1536;
										assign node1536 = (inp[3]) ? 3'b100 : node1537;
											assign node1537 = (inp[5]) ? 3'b100 : 3'b110;
										assign node1541 = (inp[3]) ? 3'b110 : node1542;
											assign node1542 = (inp[5]) ? 3'b110 : 3'b100;
									assign node1546 = (inp[8]) ? node1552 : node1547;
										assign node1547 = (inp[5]) ? 3'b110 : node1548;
											assign node1548 = (inp[3]) ? 3'b110 : 3'b100;
										assign node1552 = (inp[5]) ? 3'b100 : node1553;
											assign node1553 = (inp[3]) ? 3'b100 : 3'b110;
								assign node1557 = (inp[4]) ? node1569 : node1558;
									assign node1558 = (inp[8]) ? node1564 : node1559;
										assign node1559 = (inp[3]) ? 3'b100 : node1560;
											assign node1560 = (inp[5]) ? 3'b100 : 3'b110;
										assign node1564 = (inp[5]) ? 3'b111 : node1565;
											assign node1565 = (inp[3]) ? 3'b111 : 3'b100;
									assign node1569 = (inp[11]) ? node1573 : node1570;
										assign node1570 = (inp[8]) ? 3'b101 : 3'b100;
										assign node1573 = (inp[8]) ? node1575 : 3'b111;
											assign node1575 = (inp[5]) ? 3'b101 : 3'b111;
							assign node1578 = (inp[0]) ? node1600 : node1579;
								assign node1579 = (inp[4]) ? node1589 : node1580;
									assign node1580 = (inp[8]) ? node1586 : node1581;
										assign node1581 = (inp[3]) ? 3'b100 : node1582;
											assign node1582 = (inp[5]) ? 3'b100 : 3'b110;
										assign node1586 = (inp[5]) ? 3'b111 : 3'b100;
									assign node1589 = (inp[8]) ? node1595 : node1590;
										assign node1590 = (inp[3]) ? 3'b111 : node1591;
											assign node1591 = (inp[5]) ? 3'b111 : 3'b100;
										assign node1595 = (inp[5]) ? 3'b101 : node1596;
											assign node1596 = (inp[3]) ? 3'b101 : 3'b111;
								assign node1600 = (inp[8]) ? node1612 : node1601;
									assign node1601 = (inp[4]) ? node1607 : node1602;
										assign node1602 = (inp[5]) ? 3'b101 : node1603;
											assign node1603 = (inp[3]) ? 3'b101 : 3'b111;
										assign node1607 = (inp[3]) ? 3'b111 : node1608;
											assign node1608 = (inp[11]) ? 3'b101 : 3'b111;
									assign node1612 = (inp[4]) ? node1618 : node1613;
										assign node1613 = (inp[3]) ? 3'b111 : node1614;
											assign node1614 = (inp[5]) ? 3'b111 : 3'b101;
										assign node1618 = (inp[3]) ? 3'b101 : node1619;
											assign node1619 = (inp[5]) ? 3'b101 : 3'b111;
					assign node1623 = (inp[7]) ? node1735 : node1624;
						assign node1624 = (inp[0]) ? node1694 : node1625;
							assign node1625 = (inp[2]) ? node1673 : node1626;
								assign node1626 = (inp[11]) ? node1652 : node1627;
									assign node1627 = (inp[5]) ? node1639 : node1628;
										assign node1628 = (inp[3]) ? node1634 : node1629;
											assign node1629 = (inp[8]) ? node1631 : 3'b100;
												assign node1631 = (inp[4]) ? 3'b110 : 3'b100;
											assign node1634 = (inp[8]) ? node1636 : 3'b110;
												assign node1636 = (inp[4]) ? 3'b100 : 3'b110;
										assign node1639 = (inp[3]) ? node1645 : node1640;
											assign node1640 = (inp[4]) ? 3'b110 : node1641;
												assign node1641 = (inp[8]) ? 3'b110 : 3'b100;
											assign node1645 = (inp[4]) ? node1649 : node1646;
												assign node1646 = (inp[8]) ? 3'b110 : 3'b100;
												assign node1649 = (inp[8]) ? 3'b100 : 3'b110;
									assign node1652 = (inp[4]) ? node1664 : node1653;
										assign node1653 = (inp[8]) ? node1659 : node1654;
											assign node1654 = (inp[5]) ? 3'b100 : node1655;
												assign node1655 = (inp[3]) ? 3'b100 : 3'b110;
											assign node1659 = (inp[3]) ? 3'b110 : node1660;
												assign node1660 = (inp[5]) ? 3'b110 : 3'b100;
										assign node1664 = (inp[8]) ? node1668 : node1665;
											assign node1665 = (inp[3]) ? 3'b110 : 3'b100;
											assign node1668 = (inp[5]) ? 3'b100 : node1669;
												assign node1669 = (inp[3]) ? 3'b100 : 3'b110;
								assign node1673 = (inp[4]) ? node1683 : node1674;
									assign node1674 = (inp[8]) ? node1680 : node1675;
										assign node1675 = (inp[3]) ? 3'b100 : node1676;
											assign node1676 = (inp[5]) ? 3'b100 : 3'b110;
										assign node1680 = (inp[5]) ? 3'b111 : 3'b100;
									assign node1683 = (inp[8]) ? node1689 : node1684;
										assign node1684 = (inp[3]) ? 3'b111 : node1685;
											assign node1685 = (inp[5]) ? 3'b111 : 3'b100;
										assign node1689 = (inp[3]) ? 3'b101 : node1690;
											assign node1690 = (inp[5]) ? 3'b101 : 3'b111;
							assign node1694 = (inp[2]) ? node1716 : node1695;
								assign node1695 = (inp[8]) ? node1707 : node1696;
									assign node1696 = (inp[4]) ? node1702 : node1697;
										assign node1697 = (inp[3]) ? 3'b100 : node1698;
											assign node1698 = (inp[5]) ? 3'b100 : 3'b110;
										assign node1702 = (inp[3]) ? 3'b111 : node1703;
											assign node1703 = (inp[5]) ? 3'b111 : 3'b100;
									assign node1707 = (inp[4]) ? node1713 : node1708;
										assign node1708 = (inp[5]) ? 3'b111 : node1709;
											assign node1709 = (inp[3]) ? 3'b111 : 3'b100;
										assign node1713 = (inp[3]) ? 3'b101 : 3'b111;
								assign node1716 = (inp[8]) ? node1724 : node1717;
									assign node1717 = (inp[4]) ? 3'b111 : node1718;
										assign node1718 = (inp[3]) ? 3'b101 : node1719;
											assign node1719 = (inp[5]) ? 3'b101 : 3'b111;
									assign node1724 = (inp[4]) ? node1730 : node1725;
										assign node1725 = (inp[3]) ? 3'b111 : node1726;
											assign node1726 = (inp[5]) ? 3'b111 : 3'b101;
										assign node1730 = (inp[3]) ? 3'b101 : node1731;
											assign node1731 = (inp[5]) ? 3'b101 : 3'b111;
						assign node1735 = (inp[2]) ? node1785 : node1736;
							assign node1736 = (inp[0]) ? node1760 : node1737;
								assign node1737 = (inp[3]) ? node1753 : node1738;
									assign node1738 = (inp[8]) ? node1746 : node1739;
										assign node1739 = (inp[4]) ? node1743 : node1740;
											assign node1740 = (inp[5]) ? 3'b101 : 3'b111;
											assign node1743 = (inp[5]) ? 3'b111 : 3'b101;
										assign node1746 = (inp[4]) ? node1750 : node1747;
											assign node1747 = (inp[5]) ? 3'b111 : 3'b101;
											assign node1750 = (inp[5]) ? 3'b101 : 3'b111;
									assign node1753 = (inp[8]) ? node1757 : node1754;
										assign node1754 = (inp[4]) ? 3'b111 : 3'b101;
										assign node1757 = (inp[4]) ? 3'b101 : 3'b111;
								assign node1760 = (inp[4]) ? node1774 : node1761;
									assign node1761 = (inp[8]) ? node1769 : node1762;
										assign node1762 = (inp[11]) ? 3'b101 : node1763;
											assign node1763 = (inp[5]) ? 3'b101 : node1764;
												assign node1764 = (inp[3]) ? 3'b101 : 3'b111;
										assign node1769 = (inp[5]) ? 3'b110 : node1770;
											assign node1770 = (inp[3]) ? 3'b110 : 3'b101;
									assign node1774 = (inp[8]) ? node1780 : node1775;
										assign node1775 = (inp[3]) ? 3'b110 : node1776;
											assign node1776 = (inp[5]) ? 3'b110 : 3'b101;
										assign node1780 = (inp[5]) ? 3'b100 : node1781;
											assign node1781 = (inp[3]) ? 3'b100 : 3'b110;
							assign node1785 = (inp[0]) ? node1809 : node1786;
								assign node1786 = (inp[8]) ? node1798 : node1787;
									assign node1787 = (inp[4]) ? node1793 : node1788;
										assign node1788 = (inp[3]) ? 3'b101 : node1789;
											assign node1789 = (inp[5]) ? 3'b101 : 3'b111;
										assign node1793 = (inp[5]) ? 3'b110 : node1794;
											assign node1794 = (inp[3]) ? 3'b110 : 3'b101;
									assign node1798 = (inp[4]) ? node1804 : node1799;
										assign node1799 = (inp[5]) ? 3'b110 : node1800;
											assign node1800 = (inp[3]) ? 3'b110 : 3'b101;
										assign node1804 = (inp[5]) ? 3'b100 : node1805;
											assign node1805 = (inp[3]) ? 3'b100 : 3'b110;
								assign node1809 = (inp[5]) ? node1825 : node1810;
									assign node1810 = (inp[4]) ? node1818 : node1811;
										assign node1811 = (inp[3]) ? node1815 : node1812;
											assign node1812 = (inp[8]) ? 3'b100 : 3'b110;
											assign node1815 = (inp[8]) ? 3'b110 : 3'b100;
										assign node1818 = (inp[3]) ? node1822 : node1819;
											assign node1819 = (inp[8]) ? 3'b110 : 3'b100;
											assign node1822 = (inp[8]) ? 3'b100 : 3'b110;
									assign node1825 = (inp[8]) ? node1829 : node1826;
										assign node1826 = (inp[4]) ? 3'b110 : 3'b100;
										assign node1829 = (inp[4]) ? 3'b100 : 3'b110;
		assign node1832 = (inp[6]) ? node2858 : node1833;
			assign node1833 = (inp[11]) ? node2383 : node1834;
				assign node1834 = (inp[1]) ? node2116 : node1835;
					assign node1835 = (inp[3]) ? node1951 : node1836;
						assign node1836 = (inp[8]) ? node1906 : node1837;
							assign node1837 = (inp[4]) ? node1867 : node1838;
								assign node1838 = (inp[0]) ? node1846 : node1839;
									assign node1839 = (inp[9]) ? node1843 : node1840;
										assign node1840 = (inp[7]) ? 3'b010 : 3'b011;
										assign node1843 = (inp[7]) ? 3'b011 : 3'b010;
									assign node1846 = (inp[5]) ? node1862 : node1847;
										assign node1847 = (inp[9]) ? node1855 : node1848;
											assign node1848 = (inp[2]) ? node1852 : node1849;
												assign node1849 = (inp[7]) ? 3'b010 : 3'b011;
												assign node1852 = (inp[7]) ? 3'b011 : 3'b010;
											assign node1855 = (inp[2]) ? node1859 : node1856;
												assign node1856 = (inp[7]) ? 3'b011 : 3'b010;
												assign node1859 = (inp[7]) ? 3'b010 : 3'b011;
										assign node1862 = (inp[7]) ? 3'b011 : node1863;
											assign node1863 = (inp[2]) ? 3'b010 : 3'b011;
								assign node1867 = (inp[2]) ? node1883 : node1868;
									assign node1868 = (inp[5]) ? node1876 : node1869;
										assign node1869 = (inp[9]) ? node1873 : node1870;
											assign node1870 = (inp[7]) ? 3'b000 : 3'b001;
											assign node1873 = (inp[7]) ? 3'b001 : 3'b000;
										assign node1876 = (inp[9]) ? node1880 : node1877;
											assign node1877 = (inp[7]) ? 3'b000 : 3'b001;
											assign node1880 = (inp[7]) ? 3'b001 : 3'b000;
									assign node1883 = (inp[5]) ? node1893 : node1884;
										assign node1884 = (inp[7]) ? node1886 : 3'b000;
											assign node1886 = (inp[9]) ? node1890 : node1887;
												assign node1887 = (inp[0]) ? 3'b001 : 3'b000;
												assign node1890 = (inp[0]) ? 3'b000 : 3'b001;
										assign node1893 = (inp[9]) ? node1901 : node1894;
											assign node1894 = (inp[7]) ? node1898 : node1895;
												assign node1895 = (inp[0]) ? 3'b000 : 3'b001;
												assign node1898 = (inp[0]) ? 3'b001 : 3'b000;
											assign node1901 = (inp[7]) ? node1903 : 3'b001;
												assign node1903 = (inp[0]) ? 3'b000 : 3'b001;
							assign node1906 = (inp[4]) ? node1930 : node1907;
								assign node1907 = (inp[7]) ? node1919 : node1908;
									assign node1908 = (inp[9]) ? node1914 : node1909;
										assign node1909 = (inp[2]) ? node1911 : 3'b001;
											assign node1911 = (inp[0]) ? 3'b000 : 3'b001;
										assign node1914 = (inp[0]) ? node1916 : 3'b000;
											assign node1916 = (inp[2]) ? 3'b001 : 3'b000;
									assign node1919 = (inp[9]) ? node1925 : node1920;
										assign node1920 = (inp[0]) ? node1922 : 3'b000;
											assign node1922 = (inp[2]) ? 3'b001 : 3'b000;
										assign node1925 = (inp[0]) ? node1927 : 3'b001;
											assign node1927 = (inp[2]) ? 3'b000 : 3'b001;
								assign node1930 = (inp[7]) ? node1940 : node1931;
									assign node1931 = (inp[9]) ? node1937 : node1932;
										assign node1932 = (inp[0]) ? 3'b010 : node1933;
											assign node1933 = (inp[2]) ? 3'b010 : 3'b011;
										assign node1937 = (inp[0]) ? 3'b011 : 3'b010;
									assign node1940 = (inp[9]) ? node1946 : node1941;
										assign node1941 = (inp[2]) ? 3'b011 : node1942;
											assign node1942 = (inp[0]) ? 3'b011 : 3'b010;
										assign node1946 = (inp[2]) ? 3'b010 : node1947;
											assign node1947 = (inp[0]) ? 3'b010 : 3'b011;
						assign node1951 = (inp[0]) ? node2027 : node1952;
							assign node1952 = (inp[9]) ? node1996 : node1953;
								assign node1953 = (inp[7]) ? node1975 : node1954;
									assign node1954 = (inp[2]) ? node1966 : node1955;
										assign node1955 = (inp[5]) ? node1961 : node1956;
											assign node1956 = (inp[4]) ? node1958 : 3'b011;
												assign node1958 = (inp[8]) ? 3'b011 : 3'b001;
											assign node1961 = (inp[4]) ? 3'b001 : node1962;
												assign node1962 = (inp[8]) ? 3'b011 : 3'b001;
										assign node1966 = (inp[4]) ? 3'b010 : node1967;
											assign node1967 = (inp[8]) ? node1971 : node1968;
												assign node1968 = (inp[5]) ? 3'b001 : 3'b011;
												assign node1971 = (inp[5]) ? 3'b010 : 3'b001;
									assign node1975 = (inp[2]) ? node1983 : node1976;
										assign node1976 = (inp[4]) ? 3'b010 : node1977;
											assign node1977 = (inp[5]) ? node1979 : 3'b000;
												assign node1979 = (inp[8]) ? 3'b010 : 3'b000;
										assign node1983 = (inp[8]) ? node1989 : node1984;
											assign node1984 = (inp[5]) ? node1986 : 3'b000;
												assign node1986 = (inp[4]) ? 3'b011 : 3'b000;
											assign node1989 = (inp[5]) ? node1993 : node1990;
												assign node1990 = (inp[4]) ? 3'b011 : 3'b000;
												assign node1993 = (inp[4]) ? 3'b001 : 3'b011;
								assign node1996 = (inp[7]) ? node2008 : node1997;
									assign node1997 = (inp[2]) ? 3'b011 : node1998;
										assign node1998 = (inp[8]) ? 3'b010 : node1999;
											assign node1999 = (inp[4]) ? node2003 : node2000;
												assign node2000 = (inp[5]) ? 3'b000 : 3'b010;
												assign node2003 = (inp[5]) ? 3'b010 : 3'b000;
									assign node2008 = (inp[2]) ? node2018 : node2009;
										assign node2009 = (inp[8]) ? 3'b011 : node2010;
											assign node2010 = (inp[4]) ? node2014 : node2011;
												assign node2011 = (inp[5]) ? 3'b001 : 3'b011;
												assign node2014 = (inp[5]) ? 3'b011 : 3'b001;
										assign node2018 = (inp[4]) ? 3'b010 : node2019;
											assign node2019 = (inp[8]) ? node2023 : node2020;
												assign node2020 = (inp[5]) ? 3'b001 : 3'b011;
												assign node2023 = (inp[5]) ? 3'b010 : 3'b001;
							assign node2027 = (inp[8]) ? node2071 : node2028;
								assign node2028 = (inp[7]) ? node2048 : node2029;
									assign node2029 = (inp[9]) ? node2039 : node2030;
										assign node2030 = (inp[2]) ? node2032 : 3'b001;
											assign node2032 = (inp[5]) ? node2036 : node2033;
												assign node2033 = (inp[4]) ? 3'b000 : 3'b010;
												assign node2036 = (inp[4]) ? 3'b010 : 3'b000;
										assign node2039 = (inp[2]) ? node2043 : node2040;
											assign node2040 = (inp[5]) ? 3'b000 : 3'b010;
											assign node2043 = (inp[5]) ? node2045 : 3'b001;
												assign node2045 = (inp[4]) ? 3'b011 : 3'b001;
									assign node2048 = (inp[9]) ? node2058 : node2049;
										assign node2049 = (inp[5]) ? node2055 : node2050;
											assign node2050 = (inp[2]) ? 3'b001 : node2051;
												assign node2051 = (inp[4]) ? 3'b000 : 3'b010;
											assign node2055 = (inp[4]) ? 3'b011 : 3'b001;
										assign node2058 = (inp[2]) ? node2066 : node2059;
											assign node2059 = (inp[4]) ? node2063 : node2060;
												assign node2060 = (inp[5]) ? 3'b001 : 3'b011;
												assign node2063 = (inp[5]) ? 3'b010 : 3'b001;
											assign node2066 = (inp[5]) ? node2068 : 3'b000;
												assign node2068 = (inp[4]) ? 3'b010 : 3'b000;
								assign node2071 = (inp[5]) ? node2093 : node2072;
									assign node2072 = (inp[4]) ? node2086 : node2073;
										assign node2073 = (inp[2]) ? node2079 : node2074;
											assign node2074 = (inp[9]) ? 3'b001 : node2075;
												assign node2075 = (inp[7]) ? 3'b000 : 3'b001;
											assign node2079 = (inp[7]) ? node2083 : node2080;
												assign node2080 = (inp[9]) ? 3'b001 : 3'b000;
												assign node2083 = (inp[9]) ? 3'b000 : 3'b001;
										assign node2086 = (inp[7]) ? node2090 : node2087;
											assign node2087 = (inp[9]) ? 3'b011 : 3'b010;
											assign node2090 = (inp[9]) ? 3'b010 : 3'b011;
									assign node2093 = (inp[4]) ? node2101 : node2094;
										assign node2094 = (inp[7]) ? node2098 : node2095;
											assign node2095 = (inp[9]) ? 3'b011 : 3'b010;
											assign node2098 = (inp[9]) ? 3'b010 : 3'b011;
										assign node2101 = (inp[2]) ? node2109 : node2102;
											assign node2102 = (inp[7]) ? node2106 : node2103;
												assign node2103 = (inp[9]) ? 3'b001 : 3'b000;
												assign node2106 = (inp[9]) ? 3'b000 : 3'b001;
											assign node2109 = (inp[9]) ? node2113 : node2110;
												assign node2110 = (inp[7]) ? 3'b001 : 3'b000;
												assign node2113 = (inp[7]) ? 3'b000 : 3'b001;
					assign node2116 = (inp[7]) ? node2246 : node2117;
						assign node2117 = (inp[9]) ? node2185 : node2118;
							assign node2118 = (inp[2]) ? node2158 : node2119;
								assign node2119 = (inp[0]) ? node2139 : node2120;
									assign node2120 = (inp[3]) ? node2134 : node2121;
										assign node2121 = (inp[8]) ? node2129 : node2122;
											assign node2122 = (inp[4]) ? node2126 : node2123;
												assign node2123 = (inp[5]) ? 3'b101 : 3'b111;
												assign node2126 = (inp[5]) ? 3'b111 : 3'b101;
											assign node2129 = (inp[4]) ? 3'b101 : node2130;
												assign node2130 = (inp[5]) ? 3'b111 : 3'b101;
										assign node2134 = (inp[8]) ? node2136 : 3'b111;
											assign node2136 = (inp[4]) ? 3'b101 : 3'b111;
									assign node2139 = (inp[8]) ? node2149 : node2140;
										assign node2140 = (inp[3]) ? node2146 : node2141;
											assign node2141 = (inp[4]) ? 3'b101 : node2142;
												assign node2142 = (inp[5]) ? 3'b101 : 3'b111;
											assign node2146 = (inp[4]) ? 3'b110 : 3'b101;
										assign node2149 = (inp[4]) ? node2153 : node2150;
											assign node2150 = (inp[5]) ? 3'b110 : 3'b101;
											assign node2153 = (inp[5]) ? 3'b100 : node2154;
												assign node2154 = (inp[3]) ? 3'b100 : 3'b110;
								assign node2158 = (inp[8]) ? node2176 : node2159;
									assign node2159 = (inp[0]) ? node2167 : node2160;
										assign node2160 = (inp[4]) ? node2164 : node2161;
											assign node2161 = (inp[3]) ? 3'b101 : 3'b111;
											assign node2164 = (inp[3]) ? 3'b110 : 3'b101;
										assign node2167 = (inp[4]) ? node2171 : node2168;
											assign node2168 = (inp[3]) ? 3'b100 : 3'b110;
											assign node2171 = (inp[3]) ? 3'b110 : node2172;
												assign node2172 = (inp[5]) ? 3'b110 : 3'b100;
									assign node2176 = (inp[4]) ? node2180 : node2177;
										assign node2177 = (inp[5]) ? 3'b110 : 3'b100;
										assign node2180 = (inp[5]) ? 3'b100 : node2181;
											assign node2181 = (inp[3]) ? 3'b100 : 3'b110;
							assign node2185 = (inp[0]) ? node2221 : node2186;
								assign node2186 = (inp[2]) ? node2204 : node2187;
									assign node2187 = (inp[4]) ? node2199 : node2188;
										assign node2188 = (inp[8]) ? node2194 : node2189;
											assign node2189 = (inp[3]) ? 3'b100 : node2190;
												assign node2190 = (inp[5]) ? 3'b100 : 3'b110;
											assign node2194 = (inp[3]) ? 3'b110 : node2195;
												assign node2195 = (inp[5]) ? 3'b110 : 3'b100;
										assign node2199 = (inp[8]) ? 3'b100 : node2200;
											assign node2200 = (inp[3]) ? 3'b110 : 3'b100;
									assign node2204 = (inp[4]) ? node2214 : node2205;
										assign node2205 = (inp[8]) ? node2209 : node2206;
											assign node2206 = (inp[5]) ? 3'b100 : 3'b110;
											assign node2209 = (inp[3]) ? 3'b111 : node2210;
												assign node2210 = (inp[5]) ? 3'b111 : 3'b100;
										assign node2214 = (inp[8]) ? 3'b101 : node2215;
											assign node2215 = (inp[3]) ? 3'b111 : node2216;
												assign node2216 = (inp[5]) ? 3'b111 : 3'b100;
								assign node2221 = (inp[2]) ? node2231 : node2222;
									assign node2222 = (inp[8]) ? node2228 : node2223;
										assign node2223 = (inp[4]) ? 3'b111 : node2224;
											assign node2224 = (inp[3]) ? 3'b100 : 3'b110;
										assign node2228 = (inp[4]) ? 3'b101 : 3'b111;
									assign node2231 = (inp[8]) ? node2237 : node2232;
										assign node2232 = (inp[4]) ? node2234 : 3'b101;
											assign node2234 = (inp[5]) ? 3'b111 : 3'b101;
										assign node2237 = (inp[4]) ? node2243 : node2238;
											assign node2238 = (inp[5]) ? 3'b111 : node2239;
												assign node2239 = (inp[3]) ? 3'b111 : 3'b101;
											assign node2243 = (inp[3]) ? 3'b101 : 3'b111;
						assign node2246 = (inp[9]) ? node2314 : node2247;
							assign node2247 = (inp[2]) ? node2285 : node2248;
								assign node2248 = (inp[0]) ? node2272 : node2249;
									assign node2249 = (inp[8]) ? node2261 : node2250;
										assign node2250 = (inp[4]) ? node2256 : node2251;
											assign node2251 = (inp[5]) ? 3'b100 : node2252;
												assign node2252 = (inp[3]) ? 3'b100 : 3'b110;
											assign node2256 = (inp[3]) ? 3'b110 : node2257;
												assign node2257 = (inp[5]) ? 3'b110 : 3'b100;
										assign node2261 = (inp[4]) ? node2267 : node2262;
											assign node2262 = (inp[5]) ? 3'b110 : node2263;
												assign node2263 = (inp[3]) ? 3'b110 : 3'b100;
											assign node2267 = (inp[5]) ? 3'b100 : node2268;
												assign node2268 = (inp[3]) ? 3'b100 : 3'b110;
									assign node2272 = (inp[4]) ? 3'b111 : node2273;
										assign node2273 = (inp[8]) ? node2279 : node2274;
											assign node2274 = (inp[5]) ? 3'b100 : node2275;
												assign node2275 = (inp[3]) ? 3'b100 : 3'b110;
											assign node2279 = (inp[3]) ? 3'b111 : node2280;
												assign node2280 = (inp[5]) ? 3'b111 : 3'b100;
								assign node2285 = (inp[0]) ? node2299 : node2286;
									assign node2286 = (inp[8]) ? node2294 : node2287;
										assign node2287 = (inp[4]) ? node2289 : 3'b100;
											assign node2289 = (inp[5]) ? 3'b111 : node2290;
												assign node2290 = (inp[3]) ? 3'b111 : 3'b100;
										assign node2294 = (inp[4]) ? node2296 : 3'b111;
											assign node2296 = (inp[5]) ? 3'b101 : 3'b111;
									assign node2299 = (inp[8]) ? node2307 : node2300;
										assign node2300 = (inp[4]) ? 3'b111 : node2301;
											assign node2301 = (inp[3]) ? 3'b101 : node2302;
												assign node2302 = (inp[5]) ? 3'b101 : 3'b111;
										assign node2307 = (inp[4]) ? node2311 : node2308;
											assign node2308 = (inp[3]) ? 3'b111 : 3'b101;
											assign node2311 = (inp[5]) ? 3'b101 : 3'b111;
							assign node2314 = (inp[0]) ? node2350 : node2315;
								assign node2315 = (inp[2]) ? node2333 : node2316;
									assign node2316 = (inp[5]) ? node2328 : node2317;
										assign node2317 = (inp[8]) ? node2323 : node2318;
											assign node2318 = (inp[3]) ? 3'b111 : node2319;
												assign node2319 = (inp[4]) ? 3'b101 : 3'b111;
											assign node2323 = (inp[4]) ? node2325 : 3'b101;
												assign node2325 = (inp[3]) ? 3'b101 : 3'b111;
										assign node2328 = (inp[8]) ? node2330 : 3'b101;
											assign node2330 = (inp[4]) ? 3'b101 : 3'b111;
									assign node2333 = (inp[4]) ? node2343 : node2334;
										assign node2334 = (inp[8]) ? node2340 : node2335;
											assign node2335 = (inp[3]) ? 3'b101 : node2336;
												assign node2336 = (inp[5]) ? 3'b101 : 3'b111;
											assign node2340 = (inp[5]) ? 3'b110 : 3'b101;
										assign node2343 = (inp[8]) ? node2345 : 3'b110;
											assign node2345 = (inp[3]) ? 3'b100 : node2346;
												assign node2346 = (inp[5]) ? 3'b100 : 3'b110;
								assign node2350 = (inp[2]) ? node2372 : node2351;
									assign node2351 = (inp[4]) ? node2361 : node2352;
										assign node2352 = (inp[8]) ? node2356 : node2353;
											assign node2353 = (inp[3]) ? 3'b101 : 3'b111;
											assign node2356 = (inp[5]) ? 3'b110 : node2357;
												assign node2357 = (inp[3]) ? 3'b110 : 3'b101;
										assign node2361 = (inp[8]) ? node2367 : node2362;
											assign node2362 = (inp[5]) ? 3'b110 : node2363;
												assign node2363 = (inp[3]) ? 3'b110 : 3'b101;
											assign node2367 = (inp[3]) ? 3'b100 : node2368;
												assign node2368 = (inp[5]) ? 3'b100 : 3'b110;
									assign node2372 = (inp[8]) ? node2378 : node2373;
										assign node2373 = (inp[4]) ? 3'b110 : node2374;
											assign node2374 = (inp[3]) ? 3'b100 : 3'b110;
										assign node2378 = (inp[4]) ? 3'b100 : node2379;
											assign node2379 = (inp[3]) ? 3'b110 : 3'b100;
				assign node2383 = (inp[5]) ? node2629 : node2384;
					assign node2384 = (inp[4]) ? node2494 : node2385;
						assign node2385 = (inp[9]) ? node2443 : node2386;
							assign node2386 = (inp[7]) ? node2412 : node2387;
								assign node2387 = (inp[2]) ? node2397 : node2388;
									assign node2388 = (inp[8]) ? node2392 : node2389;
										assign node2389 = (inp[3]) ? 3'b101 : 3'b111;
										assign node2392 = (inp[3]) ? node2394 : 3'b101;
											assign node2394 = (inp[0]) ? 3'b110 : 3'b111;
									assign node2397 = (inp[0]) ? node2403 : node2398;
										assign node2398 = (inp[3]) ? 3'b110 : node2399;
											assign node2399 = (inp[8]) ? 3'b101 : 3'b111;
										assign node2403 = (inp[1]) ? node2405 : 3'b110;
											assign node2405 = (inp[3]) ? node2409 : node2406;
												assign node2406 = (inp[8]) ? 3'b100 : 3'b110;
												assign node2409 = (inp[8]) ? 3'b110 : 3'b100;
								assign node2412 = (inp[2]) ? node2428 : node2413;
									assign node2413 = (inp[0]) ? node2421 : node2414;
										assign node2414 = (inp[3]) ? node2418 : node2415;
											assign node2415 = (inp[8]) ? 3'b100 : 3'b110;
											assign node2418 = (inp[8]) ? 3'b110 : 3'b100;
										assign node2421 = (inp[3]) ? node2425 : node2422;
											assign node2422 = (inp[8]) ? 3'b100 : 3'b110;
											assign node2425 = (inp[8]) ? 3'b111 : 3'b100;
									assign node2428 = (inp[0]) ? node2436 : node2429;
										assign node2429 = (inp[3]) ? node2433 : node2430;
											assign node2430 = (inp[8]) ? 3'b100 : 3'b110;
											assign node2433 = (inp[8]) ? 3'b111 : 3'b100;
										assign node2436 = (inp[8]) ? node2440 : node2437;
											assign node2437 = (inp[3]) ? 3'b101 : 3'b111;
											assign node2440 = (inp[3]) ? 3'b111 : 3'b101;
							assign node2443 = (inp[7]) ? node2467 : node2444;
								assign node2444 = (inp[0]) ? node2454 : node2445;
									assign node2445 = (inp[8]) ? node2449 : node2446;
										assign node2446 = (inp[3]) ? 3'b100 : 3'b110;
										assign node2449 = (inp[3]) ? node2451 : 3'b100;
											assign node2451 = (inp[2]) ? 3'b111 : 3'b110;
									assign node2454 = (inp[2]) ? node2460 : node2455;
										assign node2455 = (inp[3]) ? 3'b111 : node2456;
											assign node2456 = (inp[8]) ? 3'b100 : 3'b110;
										assign node2460 = (inp[8]) ? node2464 : node2461;
											assign node2461 = (inp[3]) ? 3'b101 : 3'b111;
											assign node2464 = (inp[3]) ? 3'b111 : 3'b101;
								assign node2467 = (inp[0]) ? node2481 : node2468;
									assign node2468 = (inp[1]) ? node2476 : node2469;
										assign node2469 = (inp[8]) ? node2473 : node2470;
											assign node2470 = (inp[3]) ? 3'b101 : 3'b111;
											assign node2473 = (inp[3]) ? 3'b111 : 3'b101;
										assign node2476 = (inp[3]) ? node2478 : 3'b101;
											assign node2478 = (inp[8]) ? 3'b111 : 3'b101;
									assign node2481 = (inp[2]) ? node2489 : node2482;
										assign node2482 = (inp[1]) ? 3'b101 : node2483;
											assign node2483 = (inp[3]) ? 3'b110 : node2484;
												assign node2484 = (inp[8]) ? 3'b101 : 3'b111;
										assign node2489 = (inp[3]) ? 3'b100 : node2490;
											assign node2490 = (inp[8]) ? 3'b100 : 3'b110;
						assign node2494 = (inp[3]) ? node2556 : node2495;
							assign node2495 = (inp[8]) ? node2513 : node2496;
								assign node2496 = (inp[9]) ? node2504 : node2497;
									assign node2497 = (inp[7]) ? node2501 : node2498;
										assign node2498 = (inp[0]) ? 3'b100 : 3'b101;
										assign node2501 = (inp[0]) ? 3'b101 : 3'b100;
									assign node2504 = (inp[7]) ? node2508 : node2505;
										assign node2505 = (inp[0]) ? 3'b101 : 3'b100;
										assign node2508 = (inp[0]) ? node2510 : 3'b101;
											assign node2510 = (inp[2]) ? 3'b100 : 3'b101;
								assign node2513 = (inp[1]) ? node2537 : node2514;
									assign node2514 = (inp[9]) ? node2526 : node2515;
										assign node2515 = (inp[7]) ? node2521 : node2516;
											assign node2516 = (inp[0]) ? 3'b110 : node2517;
												assign node2517 = (inp[2]) ? 3'b110 : 3'b111;
											assign node2521 = (inp[2]) ? 3'b111 : node2522;
												assign node2522 = (inp[0]) ? 3'b111 : 3'b110;
										assign node2526 = (inp[7]) ? node2532 : node2527;
											assign node2527 = (inp[2]) ? 3'b111 : node2528;
												assign node2528 = (inp[0]) ? 3'b111 : 3'b110;
											assign node2532 = (inp[2]) ? 3'b110 : node2533;
												assign node2533 = (inp[0]) ? 3'b110 : 3'b111;
									assign node2537 = (inp[9]) ? node2545 : node2538;
										assign node2538 = (inp[7]) ? node2540 : 3'b110;
											assign node2540 = (inp[2]) ? 3'b111 : node2541;
												assign node2541 = (inp[0]) ? 3'b111 : 3'b110;
										assign node2545 = (inp[7]) ? node2551 : node2546;
											assign node2546 = (inp[2]) ? 3'b111 : node2547;
												assign node2547 = (inp[0]) ? 3'b111 : 3'b110;
											assign node2551 = (inp[0]) ? 3'b110 : node2552;
												assign node2552 = (inp[2]) ? 3'b110 : 3'b111;
							assign node2556 = (inp[8]) ? node2596 : node2557;
								assign node2557 = (inp[1]) ? node2577 : node2558;
									assign node2558 = (inp[2]) ? node2572 : node2559;
										assign node2559 = (inp[0]) ? node2567 : node2560;
											assign node2560 = (inp[7]) ? node2564 : node2561;
												assign node2561 = (inp[9]) ? 3'b110 : 3'b111;
												assign node2564 = (inp[9]) ? 3'b111 : 3'b110;
											assign node2567 = (inp[9]) ? 3'b111 : node2568;
												assign node2568 = (inp[7]) ? 3'b111 : 3'b110;
										assign node2572 = (inp[9]) ? node2574 : 3'b110;
											assign node2574 = (inp[7]) ? 3'b110 : 3'b111;
									assign node2577 = (inp[7]) ? node2587 : node2578;
										assign node2578 = (inp[0]) ? 3'b111 : node2579;
											assign node2579 = (inp[9]) ? node2583 : node2580;
												assign node2580 = (inp[2]) ? 3'b110 : 3'b111;
												assign node2583 = (inp[2]) ? 3'b111 : 3'b110;
										assign node2587 = (inp[2]) ? node2593 : node2588;
											assign node2588 = (inp[0]) ? 3'b110 : node2589;
												assign node2589 = (inp[9]) ? 3'b111 : 3'b110;
											assign node2593 = (inp[9]) ? 3'b110 : 3'b111;
								assign node2596 = (inp[2]) ? node2622 : node2597;
									assign node2597 = (inp[0]) ? node2609 : node2598;
										assign node2598 = (inp[1]) ? node2604 : node2599;
											assign node2599 = (inp[9]) ? node2601 : 3'b100;
												assign node2601 = (inp[7]) ? 3'b101 : 3'b100;
											assign node2604 = (inp[7]) ? 3'b100 : node2605;
												assign node2605 = (inp[9]) ? 3'b100 : 3'b101;
										assign node2609 = (inp[1]) ? node2617 : node2610;
											assign node2610 = (inp[9]) ? node2614 : node2611;
												assign node2611 = (inp[7]) ? 3'b101 : 3'b100;
												assign node2614 = (inp[7]) ? 3'b100 : 3'b101;
											assign node2617 = (inp[7]) ? 3'b101 : node2618;
												assign node2618 = (inp[9]) ? 3'b101 : 3'b100;
									assign node2622 = (inp[9]) ? node2626 : node2623;
										assign node2623 = (inp[7]) ? 3'b101 : 3'b100;
										assign node2626 = (inp[7]) ? 3'b100 : 3'b101;
					assign node2629 = (inp[2]) ? node2733 : node2630;
						assign node2630 = (inp[8]) ? node2676 : node2631;
							assign node2631 = (inp[4]) ? node2653 : node2632;
								assign node2632 = (inp[3]) ? node2640 : node2633;
									assign node2633 = (inp[9]) ? node2637 : node2634;
										assign node2634 = (inp[7]) ? 3'b100 : 3'b101;
										assign node2637 = (inp[7]) ? 3'b101 : 3'b100;
									assign node2640 = (inp[0]) ? node2648 : node2641;
										assign node2641 = (inp[9]) ? node2645 : node2642;
											assign node2642 = (inp[7]) ? 3'b100 : 3'b101;
											assign node2645 = (inp[7]) ? 3'b101 : 3'b100;
										assign node2648 = (inp[7]) ? 3'b101 : node2649;
											assign node2649 = (inp[9]) ? 3'b100 : 3'b101;
								assign node2653 = (inp[1]) ? node2661 : node2654;
									assign node2654 = (inp[3]) ? 3'b110 : node2655;
										assign node2655 = (inp[7]) ? 3'b110 : node2656;
											assign node2656 = (inp[9]) ? 3'b110 : 3'b111;
									assign node2661 = (inp[7]) ? node2669 : node2662;
										assign node2662 = (inp[0]) ? node2666 : node2663;
											assign node2663 = (inp[9]) ? 3'b110 : 3'b111;
											assign node2666 = (inp[9]) ? 3'b111 : 3'b110;
										assign node2669 = (inp[3]) ? 3'b111 : node2670;
											assign node2670 = (inp[0]) ? 3'b110 : node2671;
												assign node2671 = (inp[9]) ? 3'b111 : 3'b110;
							assign node2676 = (inp[4]) ? node2702 : node2677;
								assign node2677 = (inp[0]) ? node2687 : node2678;
									assign node2678 = (inp[3]) ? node2680 : 3'b111;
										assign node2680 = (inp[9]) ? node2684 : node2681;
											assign node2681 = (inp[7]) ? 3'b110 : 3'b111;
											assign node2684 = (inp[7]) ? 3'b111 : 3'b110;
									assign node2687 = (inp[1]) ? node2697 : node2688;
										assign node2688 = (inp[3]) ? 3'b110 : node2689;
											assign node2689 = (inp[9]) ? node2693 : node2690;
												assign node2690 = (inp[7]) ? 3'b111 : 3'b110;
												assign node2693 = (inp[7]) ? 3'b110 : 3'b111;
										assign node2697 = (inp[7]) ? node2699 : 3'b110;
											assign node2699 = (inp[9]) ? 3'b110 : 3'b111;
								assign node2702 = (inp[7]) ? node2712 : node2703;
									assign node2703 = (inp[3]) ? 3'b101 : node2704;
										assign node2704 = (inp[0]) ? node2708 : node2705;
											assign node2705 = (inp[9]) ? 3'b100 : 3'b101;
											assign node2708 = (inp[9]) ? 3'b101 : 3'b100;
									assign node2712 = (inp[3]) ? node2720 : node2713;
										assign node2713 = (inp[9]) ? node2717 : node2714;
											assign node2714 = (inp[0]) ? 3'b101 : 3'b100;
											assign node2717 = (inp[0]) ? 3'b100 : 3'b101;
										assign node2720 = (inp[1]) ? node2726 : node2721;
											assign node2721 = (inp[9]) ? 3'b100 : node2722;
												assign node2722 = (inp[0]) ? 3'b101 : 3'b100;
											assign node2726 = (inp[9]) ? node2730 : node2727;
												assign node2727 = (inp[0]) ? 3'b101 : 3'b100;
												assign node2730 = (inp[0]) ? 3'b100 : 3'b101;
						assign node2733 = (inp[1]) ? node2819 : node2734;
							assign node2734 = (inp[3]) ? node2782 : node2735;
								assign node2735 = (inp[8]) ? node2755 : node2736;
									assign node2736 = (inp[4]) ? node2740 : node2737;
										assign node2737 = (inp[9]) ? 3'b101 : 3'b100;
										assign node2740 = (inp[0]) ? node2748 : node2741;
											assign node2741 = (inp[7]) ? node2745 : node2742;
												assign node2742 = (inp[9]) ? 3'b111 : 3'b110;
												assign node2745 = (inp[9]) ? 3'b110 : 3'b111;
											assign node2748 = (inp[9]) ? node2752 : node2749;
												assign node2749 = (inp[7]) ? 3'b111 : 3'b110;
												assign node2752 = (inp[7]) ? 3'b110 : 3'b111;
									assign node2755 = (inp[4]) ? node2769 : node2756;
										assign node2756 = (inp[0]) ? node2762 : node2757;
											assign node2757 = (inp[9]) ? 3'b110 : node2758;
												assign node2758 = (inp[7]) ? 3'b111 : 3'b110;
											assign node2762 = (inp[9]) ? node2766 : node2763;
												assign node2763 = (inp[7]) ? 3'b111 : 3'b110;
												assign node2766 = (inp[7]) ? 3'b110 : 3'b111;
										assign node2769 = (inp[0]) ? node2777 : node2770;
											assign node2770 = (inp[9]) ? node2774 : node2771;
												assign node2771 = (inp[7]) ? 3'b101 : 3'b100;
												assign node2774 = (inp[7]) ? 3'b100 : 3'b101;
											assign node2777 = (inp[9]) ? 3'b100 : node2778;
												assign node2778 = (inp[7]) ? 3'b101 : 3'b100;
								assign node2782 = (inp[8]) ? node2802 : node2783;
									assign node2783 = (inp[4]) ? node2797 : node2784;
										assign node2784 = (inp[7]) ? node2792 : node2785;
											assign node2785 = (inp[9]) ? node2789 : node2786;
												assign node2786 = (inp[0]) ? 3'b100 : 3'b101;
												assign node2789 = (inp[0]) ? 3'b101 : 3'b100;
											assign node2792 = (inp[9]) ? 3'b101 : node2793;
												assign node2793 = (inp[0]) ? 3'b101 : 3'b100;
										assign node2797 = (inp[9]) ? 3'b111 : node2798;
											assign node2798 = (inp[7]) ? 3'b111 : 3'b110;
									assign node2802 = (inp[4]) ? node2810 : node2803;
										assign node2803 = (inp[9]) ? node2807 : node2804;
											assign node2804 = (inp[7]) ? 3'b111 : 3'b110;
											assign node2807 = (inp[7]) ? 3'b110 : 3'b111;
										assign node2810 = (inp[0]) ? node2814 : node2811;
											assign node2811 = (inp[7]) ? 3'b100 : 3'b101;
											assign node2814 = (inp[7]) ? 3'b101 : node2815;
												assign node2815 = (inp[9]) ? 3'b101 : 3'b100;
							assign node2819 = (inp[7]) ? node2839 : node2820;
								assign node2820 = (inp[9]) ? node2830 : node2821;
									assign node2821 = (inp[8]) ? node2827 : node2822;
										assign node2822 = (inp[4]) ? 3'b110 : node2823;
											assign node2823 = (inp[0]) ? 3'b100 : 3'b101;
										assign node2827 = (inp[4]) ? 3'b100 : 3'b110;
									assign node2830 = (inp[0]) ? 3'b101 : node2831;
										assign node2831 = (inp[4]) ? node2835 : node2832;
											assign node2832 = (inp[8]) ? 3'b111 : 3'b100;
											assign node2835 = (inp[8]) ? 3'b101 : 3'b111;
								assign node2839 = (inp[9]) ? node2849 : node2840;
									assign node2840 = (inp[4]) ? node2846 : node2841;
										assign node2841 = (inp[8]) ? 3'b111 : node2842;
											assign node2842 = (inp[0]) ? 3'b101 : 3'b100;
										assign node2846 = (inp[8]) ? 3'b101 : 3'b111;
									assign node2849 = (inp[8]) ? node2855 : node2850;
										assign node2850 = (inp[0]) ? node2852 : 3'b101;
											assign node2852 = (inp[4]) ? 3'b110 : 3'b100;
										assign node2855 = (inp[4]) ? 3'b100 : 3'b110;
			assign node2858 = (inp[1]) ? node3388 : node2859;
				assign node2859 = (inp[11]) ? node3121 : node2860;
					assign node2860 = (inp[0]) ? node2994 : node2861;
						assign node2861 = (inp[8]) ? node2929 : node2862;
							assign node2862 = (inp[4]) ? node2898 : node2863;
								assign node2863 = (inp[5]) ? node2879 : node2864;
									assign node2864 = (inp[3]) ? node2872 : node2865;
										assign node2865 = (inp[9]) ? node2869 : node2866;
											assign node2866 = (inp[7]) ? 3'b110 : 3'b111;
											assign node2869 = (inp[7]) ? 3'b111 : 3'b110;
										assign node2872 = (inp[7]) ? node2876 : node2873;
											assign node2873 = (inp[9]) ? 3'b100 : 3'b101;
											assign node2876 = (inp[9]) ? 3'b101 : 3'b100;
									assign node2879 = (inp[2]) ? node2885 : node2880;
										assign node2880 = (inp[7]) ? node2882 : 3'b101;
											assign node2882 = (inp[9]) ? 3'b101 : 3'b100;
										assign node2885 = (inp[3]) ? node2893 : node2886;
											assign node2886 = (inp[7]) ? node2890 : node2887;
												assign node2887 = (inp[9]) ? 3'b100 : 3'b101;
												assign node2890 = (inp[9]) ? 3'b101 : 3'b100;
											assign node2893 = (inp[9]) ? 3'b100 : node2894;
												assign node2894 = (inp[7]) ? 3'b100 : 3'b101;
								assign node2898 = (inp[3]) ? node2916 : node2899;
									assign node2899 = (inp[5]) ? node2907 : node2900;
										assign node2900 = (inp[9]) ? node2904 : node2901;
											assign node2901 = (inp[7]) ? 3'b100 : 3'b101;
											assign node2904 = (inp[7]) ? 3'b101 : 3'b100;
										assign node2907 = (inp[7]) ? 3'b110 : node2908;
											assign node2908 = (inp[2]) ? node2912 : node2909;
												assign node2909 = (inp[9]) ? 3'b110 : 3'b111;
												assign node2912 = (inp[9]) ? 3'b111 : 3'b110;
									assign node2916 = (inp[9]) ? node2924 : node2917;
										assign node2917 = (inp[7]) ? node2921 : node2918;
											assign node2918 = (inp[2]) ? 3'b110 : 3'b111;
											assign node2921 = (inp[2]) ? 3'b111 : 3'b110;
										assign node2924 = (inp[2]) ? 3'b110 : node2925;
											assign node2925 = (inp[7]) ? 3'b111 : 3'b110;
							assign node2929 = (inp[4]) ? node2965 : node2930;
								assign node2930 = (inp[5]) ? node2944 : node2931;
									assign node2931 = (inp[3]) ? node2937 : node2932;
										assign node2932 = (inp[9]) ? 3'b100 : node2933;
											assign node2933 = (inp[7]) ? 3'b100 : 3'b101;
										assign node2937 = (inp[9]) ? node2939 : 3'b111;
											assign node2939 = (inp[2]) ? 3'b111 : node2940;
												assign node2940 = (inp[7]) ? 3'b111 : 3'b110;
									assign node2944 = (inp[9]) ? node2960 : node2945;
										assign node2945 = (inp[3]) ? node2953 : node2946;
											assign node2946 = (inp[2]) ? node2950 : node2947;
												assign node2947 = (inp[7]) ? 3'b110 : 3'b111;
												assign node2950 = (inp[7]) ? 3'b111 : 3'b110;
											assign node2953 = (inp[2]) ? node2957 : node2954;
												assign node2954 = (inp[7]) ? 3'b110 : 3'b111;
												assign node2957 = (inp[7]) ? 3'b111 : 3'b110;
										assign node2960 = (inp[7]) ? 3'b111 : node2961;
											assign node2961 = (inp[2]) ? 3'b111 : 3'b110;
								assign node2965 = (inp[3]) ? node2985 : node2966;
									assign node2966 = (inp[5]) ? node2980 : node2967;
										assign node2967 = (inp[2]) ? node2973 : node2968;
											assign node2968 = (inp[9]) ? 3'b110 : node2969;
												assign node2969 = (inp[7]) ? 3'b110 : 3'b111;
											assign node2973 = (inp[9]) ? node2977 : node2974;
												assign node2974 = (inp[7]) ? 3'b111 : 3'b110;
												assign node2977 = (inp[7]) ? 3'b110 : 3'b111;
										assign node2980 = (inp[2]) ? 3'b101 : node2981;
											assign node2981 = (inp[9]) ? 3'b101 : 3'b100;
									assign node2985 = (inp[2]) ? node2987 : 3'b101;
										assign node2987 = (inp[7]) ? node2991 : node2988;
											assign node2988 = (inp[9]) ? 3'b101 : 3'b100;
											assign node2991 = (inp[9]) ? 3'b100 : 3'b101;
						assign node2994 = (inp[4]) ? node3062 : node2995;
							assign node2995 = (inp[8]) ? node3039 : node2996;
								assign node2996 = (inp[5]) ? node3018 : node2997;
									assign node2997 = (inp[3]) ? node3011 : node2998;
										assign node2998 = (inp[2]) ? node3004 : node2999;
											assign node2999 = (inp[9]) ? 3'b111 : node3000;
												assign node3000 = (inp[7]) ? 3'b110 : 3'b111;
											assign node3004 = (inp[9]) ? node3008 : node3005;
												assign node3005 = (inp[7]) ? 3'b111 : 3'b110;
												assign node3008 = (inp[7]) ? 3'b110 : 3'b111;
										assign node3011 = (inp[9]) ? node3013 : 3'b100;
											assign node3013 = (inp[2]) ? node3015 : 3'b100;
												assign node3015 = (inp[7]) ? 3'b100 : 3'b101;
									assign node3018 = (inp[7]) ? node3024 : node3019;
										assign node3019 = (inp[9]) ? 3'b100 : node3020;
											assign node3020 = (inp[2]) ? 3'b100 : 3'b101;
										assign node3024 = (inp[3]) ? node3032 : node3025;
											assign node3025 = (inp[2]) ? node3029 : node3026;
												assign node3026 = (inp[9]) ? 3'b101 : 3'b100;
												assign node3029 = (inp[9]) ? 3'b100 : 3'b101;
											assign node3032 = (inp[9]) ? node3036 : node3033;
												assign node3033 = (inp[2]) ? 3'b101 : 3'b100;
												assign node3036 = (inp[2]) ? 3'b100 : 3'b101;
								assign node3039 = (inp[5]) ? node3055 : node3040;
									assign node3040 = (inp[3]) ? node3048 : node3041;
										assign node3041 = (inp[7]) ? 3'b100 : node3042;
											assign node3042 = (inp[2]) ? node3044 : 3'b100;
												assign node3044 = (inp[9]) ? 3'b101 : 3'b100;
										assign node3048 = (inp[7]) ? node3052 : node3049;
											assign node3049 = (inp[9]) ? 3'b111 : 3'b110;
											assign node3052 = (inp[9]) ? 3'b110 : 3'b111;
									assign node3055 = (inp[9]) ? node3059 : node3056;
										assign node3056 = (inp[7]) ? 3'b111 : 3'b110;
										assign node3059 = (inp[7]) ? 3'b110 : 3'b111;
							assign node3062 = (inp[8]) ? node3098 : node3063;
								assign node3063 = (inp[5]) ? node3085 : node3064;
									assign node3064 = (inp[3]) ? node3078 : node3065;
										assign node3065 = (inp[7]) ? node3073 : node3066;
											assign node3066 = (inp[9]) ? node3070 : node3067;
												assign node3067 = (inp[2]) ? 3'b100 : 3'b101;
												assign node3070 = (inp[2]) ? 3'b101 : 3'b100;
											assign node3073 = (inp[9]) ? node3075 : 3'b100;
												assign node3075 = (inp[2]) ? 3'b100 : 3'b101;
										assign node3078 = (inp[7]) ? node3082 : node3079;
											assign node3079 = (inp[9]) ? 3'b111 : 3'b110;
											assign node3082 = (inp[9]) ? 3'b110 : 3'b111;
									assign node3085 = (inp[2]) ? node3093 : node3086;
										assign node3086 = (inp[7]) ? node3090 : node3087;
											assign node3087 = (inp[9]) ? 3'b111 : 3'b110;
											assign node3090 = (inp[9]) ? 3'b110 : 3'b111;
										assign node3093 = (inp[7]) ? node3095 : 3'b111;
											assign node3095 = (inp[9]) ? 3'b110 : 3'b111;
								assign node3098 = (inp[5]) ? node3114 : node3099;
									assign node3099 = (inp[3]) ? node3109 : node3100;
										assign node3100 = (inp[2]) ? 3'b111 : node3101;
											assign node3101 = (inp[7]) ? node3105 : node3102;
												assign node3102 = (inp[9]) ? 3'b111 : 3'b110;
												assign node3105 = (inp[9]) ? 3'b110 : 3'b111;
										assign node3109 = (inp[7]) ? node3111 : 3'b101;
											assign node3111 = (inp[9]) ? 3'b100 : 3'b101;
									assign node3114 = (inp[7]) ? node3118 : node3115;
										assign node3115 = (inp[9]) ? 3'b101 : 3'b100;
										assign node3118 = (inp[9]) ? 3'b100 : 3'b101;
					assign node3121 = (inp[2]) ? node3265 : node3122;
						assign node3122 = (inp[5]) ? node3184 : node3123;
							assign node3123 = (inp[0]) ? node3153 : node3124;
								assign node3124 = (inp[9]) ? node3138 : node3125;
									assign node3125 = (inp[7]) ? node3133 : node3126;
										assign node3126 = (inp[4]) ? 3'b001 : node3127;
											assign node3127 = (inp[8]) ? node3129 : 3'b011;
												assign node3129 = (inp[3]) ? 3'b011 : 3'b001;
										assign node3133 = (inp[8]) ? 3'b000 : node3134;
											assign node3134 = (inp[3]) ? 3'b010 : 3'b000;
									assign node3138 = (inp[7]) ? 3'b011 : node3139;
										assign node3139 = (inp[3]) ? node3145 : node3140;
											assign node3140 = (inp[4]) ? node3142 : 3'b010;
												assign node3142 = (inp[8]) ? 3'b010 : 3'b000;
											assign node3145 = (inp[8]) ? node3149 : node3146;
												assign node3146 = (inp[4]) ? 3'b010 : 3'b000;
												assign node3149 = (inp[4]) ? 3'b000 : 3'b010;
								assign node3153 = (inp[3]) ? node3173 : node3154;
									assign node3154 = (inp[7]) ? node3164 : node3155;
										assign node3155 = (inp[4]) ? node3161 : node3156;
											assign node3156 = (inp[8]) ? node3158 : 3'b010;
												assign node3158 = (inp[9]) ? 3'b000 : 3'b001;
											assign node3161 = (inp[9]) ? 3'b011 : 3'b010;
										assign node3164 = (inp[8]) ? node3170 : node3165;
											assign node3165 = (inp[9]) ? node3167 : 3'b010;
												assign node3167 = (inp[4]) ? 3'b001 : 3'b011;
											assign node3170 = (inp[9]) ? 3'b010 : 3'b011;
									assign node3173 = (inp[9]) ? node3177 : node3174;
										assign node3174 = (inp[7]) ? 3'b011 : 3'b010;
										assign node3177 = (inp[7]) ? node3179 : 3'b011;
											assign node3179 = (inp[8]) ? 3'b010 : node3180;
												assign node3180 = (inp[4]) ? 3'b010 : 3'b001;
							assign node3184 = (inp[0]) ? node3224 : node3185;
								assign node3185 = (inp[4]) ? node3207 : node3186;
									assign node3186 = (inp[8]) ? node3200 : node3187;
										assign node3187 = (inp[3]) ? node3195 : node3188;
											assign node3188 = (inp[9]) ? node3192 : node3189;
												assign node3189 = (inp[7]) ? 3'b000 : 3'b001;
												assign node3192 = (inp[7]) ? 3'b001 : 3'b000;
											assign node3195 = (inp[7]) ? node3197 : 3'b000;
												assign node3197 = (inp[9]) ? 3'b001 : 3'b000;
										assign node3200 = (inp[9]) ? node3204 : node3201;
											assign node3201 = (inp[7]) ? 3'b010 : 3'b011;
											assign node3204 = (inp[7]) ? 3'b011 : 3'b010;
									assign node3207 = (inp[8]) ? node3213 : node3208;
										assign node3208 = (inp[9]) ? node3210 : 3'b011;
											assign node3210 = (inp[7]) ? 3'b011 : 3'b010;
										assign node3213 = (inp[3]) ? node3219 : node3214;
											assign node3214 = (inp[9]) ? 3'b000 : node3215;
												assign node3215 = (inp[7]) ? 3'b000 : 3'b001;
											assign node3219 = (inp[9]) ? 3'b001 : node3220;
												assign node3220 = (inp[7]) ? 3'b000 : 3'b001;
								assign node3224 = (inp[4]) ? node3246 : node3225;
									assign node3225 = (inp[8]) ? node3241 : node3226;
										assign node3226 = (inp[3]) ? node3234 : node3227;
											assign node3227 = (inp[9]) ? node3231 : node3228;
												assign node3228 = (inp[7]) ? 3'b000 : 3'b001;
												assign node3231 = (inp[7]) ? 3'b001 : 3'b000;
											assign node3234 = (inp[7]) ? node3238 : node3235;
												assign node3235 = (inp[9]) ? 3'b000 : 3'b001;
												assign node3238 = (inp[9]) ? 3'b001 : 3'b000;
										assign node3241 = (inp[7]) ? node3243 : 3'b010;
											assign node3243 = (inp[9]) ? 3'b010 : 3'b011;
									assign node3246 = (inp[8]) ? node3258 : node3247;
										assign node3247 = (inp[3]) ? node3253 : node3248;
											assign node3248 = (inp[7]) ? 3'b010 : node3249;
												assign node3249 = (inp[9]) ? 3'b011 : 3'b010;
											assign node3253 = (inp[9]) ? 3'b010 : node3254;
												assign node3254 = (inp[7]) ? 3'b011 : 3'b010;
										assign node3258 = (inp[7]) ? node3262 : node3259;
											assign node3259 = (inp[3]) ? 3'b000 : 3'b001;
											assign node3262 = (inp[9]) ? 3'b000 : 3'b001;
						assign node3265 = (inp[4]) ? node3333 : node3266;
							assign node3266 = (inp[8]) ? node3310 : node3267;
								assign node3267 = (inp[5]) ? node3291 : node3268;
									assign node3268 = (inp[3]) ? node3280 : node3269;
										assign node3269 = (inp[0]) ? node3275 : node3270;
											assign node3270 = (inp[7]) ? 3'b011 : node3271;
												assign node3271 = (inp[9]) ? 3'b010 : 3'b011;
											assign node3275 = (inp[9]) ? node3277 : 3'b010;
												assign node3277 = (inp[7]) ? 3'b010 : 3'b011;
										assign node3280 = (inp[7]) ? node3286 : node3281;
											assign node3281 = (inp[0]) ? 3'b000 : node3282;
												assign node3282 = (inp[9]) ? 3'b000 : 3'b001;
											assign node3286 = (inp[0]) ? 3'b001 : node3287;
												assign node3287 = (inp[9]) ? 3'b001 : 3'b000;
									assign node3291 = (inp[7]) ? node3303 : node3292;
										assign node3292 = (inp[3]) ? node3298 : node3293;
											assign node3293 = (inp[0]) ? 3'b001 : node3294;
												assign node3294 = (inp[9]) ? 3'b000 : 3'b001;
											assign node3298 = (inp[0]) ? node3300 : 3'b001;
												assign node3300 = (inp[9]) ? 3'b001 : 3'b000;
										assign node3303 = (inp[9]) ? node3307 : node3304;
											assign node3304 = (inp[0]) ? 3'b001 : 3'b000;
											assign node3307 = (inp[0]) ? 3'b000 : 3'b001;
								assign node3310 = (inp[5]) ? node3326 : node3311;
									assign node3311 = (inp[3]) ? node3321 : node3312;
										assign node3312 = (inp[9]) ? node3314 : 3'b001;
											assign node3314 = (inp[0]) ? node3318 : node3315;
												assign node3315 = (inp[7]) ? 3'b001 : 3'b000;
												assign node3318 = (inp[7]) ? 3'b000 : 3'b001;
										assign node3321 = (inp[9]) ? node3323 : 3'b011;
											assign node3323 = (inp[7]) ? 3'b010 : 3'b011;
									assign node3326 = (inp[7]) ? node3330 : node3327;
										assign node3327 = (inp[9]) ? 3'b011 : 3'b010;
										assign node3330 = (inp[9]) ? 3'b010 : 3'b011;
							assign node3333 = (inp[8]) ? node3369 : node3334;
								assign node3334 = (inp[3]) ? node3348 : node3335;
									assign node3335 = (inp[5]) ? node3343 : node3336;
										assign node3336 = (inp[0]) ? node3338 : 3'b000;
											assign node3338 = (inp[9]) ? 3'b001 : node3339;
												assign node3339 = (inp[7]) ? 3'b001 : 3'b000;
										assign node3343 = (inp[7]) ? 3'b010 : node3344;
											assign node3344 = (inp[9]) ? 3'b011 : 3'b010;
									assign node3348 = (inp[0]) ? node3362 : node3349;
										assign node3349 = (inp[5]) ? node3357 : node3350;
											assign node3350 = (inp[7]) ? node3354 : node3351;
												assign node3351 = (inp[9]) ? 3'b011 : 3'b010;
												assign node3354 = (inp[9]) ? 3'b010 : 3'b011;
											assign node3357 = (inp[9]) ? 3'b011 : node3358;
												assign node3358 = (inp[7]) ? 3'b011 : 3'b010;
										assign node3362 = (inp[7]) ? node3366 : node3363;
											assign node3363 = (inp[9]) ? 3'b011 : 3'b010;
											assign node3366 = (inp[9]) ? 3'b010 : 3'b011;
								assign node3369 = (inp[3]) ? node3381 : node3370;
									assign node3370 = (inp[5]) ? node3376 : node3371;
										assign node3371 = (inp[7]) ? node3373 : 3'b011;
											assign node3373 = (inp[9]) ? 3'b010 : 3'b011;
										assign node3376 = (inp[9]) ? node3378 : 3'b000;
											assign node3378 = (inp[7]) ? 3'b000 : 3'b001;
									assign node3381 = (inp[9]) ? node3385 : node3382;
										assign node3382 = (inp[7]) ? 3'b001 : 3'b000;
										assign node3385 = (inp[7]) ? 3'b000 : 3'b001;
				assign node3388 = (inp[0]) ? node3594 : node3389;
					assign node3389 = (inp[9]) ? node3485 : node3390;
						assign node3390 = (inp[7]) ? node3442 : node3391;
							assign node3391 = (inp[2]) ? node3421 : node3392;
								assign node3392 = (inp[3]) ? node3402 : node3393;
									assign node3393 = (inp[8]) ? 3'b001 : node3394;
										assign node3394 = (inp[5]) ? node3398 : node3395;
											assign node3395 = (inp[4]) ? 3'b001 : 3'b011;
											assign node3398 = (inp[4]) ? 3'b011 : 3'b001;
									assign node3402 = (inp[5]) ? node3416 : node3403;
										assign node3403 = (inp[11]) ? node3411 : node3404;
											assign node3404 = (inp[4]) ? node3408 : node3405;
												assign node3405 = (inp[8]) ? 3'b011 : 3'b001;
												assign node3408 = (inp[8]) ? 3'b001 : 3'b011;
											assign node3411 = (inp[4]) ? node3413 : 3'b001;
												assign node3413 = (inp[8]) ? 3'b001 : 3'b011;
										assign node3416 = (inp[4]) ? 3'b011 : node3417;
											assign node3417 = (inp[8]) ? 3'b011 : 3'b001;
								assign node3421 = (inp[4]) ? node3431 : node3422;
									assign node3422 = (inp[8]) ? node3428 : node3423;
										assign node3423 = (inp[5]) ? 3'b001 : node3424;
											assign node3424 = (inp[3]) ? 3'b001 : 3'b011;
										assign node3428 = (inp[5]) ? 3'b010 : 3'b001;
									assign node3431 = (inp[8]) ? node3437 : node3432;
										assign node3432 = (inp[5]) ? 3'b010 : node3433;
											assign node3433 = (inp[3]) ? 3'b010 : 3'b001;
										assign node3437 = (inp[5]) ? 3'b000 : node3438;
											assign node3438 = (inp[3]) ? 3'b000 : 3'b010;
							assign node3442 = (inp[2]) ? node3466 : node3443;
								assign node3443 = (inp[3]) ? node3459 : node3444;
									assign node3444 = (inp[8]) ? node3452 : node3445;
										assign node3445 = (inp[11]) ? node3447 : 3'b000;
											assign node3447 = (inp[5]) ? 3'b000 : node3448;
												assign node3448 = (inp[4]) ? 3'b000 : 3'b010;
										assign node3452 = (inp[5]) ? node3456 : node3453;
											assign node3453 = (inp[11]) ? 3'b000 : 3'b010;
											assign node3456 = (inp[4]) ? 3'b000 : 3'b010;
									assign node3459 = (inp[4]) ? node3463 : node3460;
										assign node3460 = (inp[8]) ? 3'b010 : 3'b000;
										assign node3463 = (inp[8]) ? 3'b000 : 3'b010;
								assign node3466 = (inp[4]) ? node3474 : node3467;
									assign node3467 = (inp[8]) ? node3469 : 3'b000;
										assign node3469 = (inp[5]) ? 3'b011 : node3470;
											assign node3470 = (inp[3]) ? 3'b011 : 3'b000;
									assign node3474 = (inp[8]) ? node3480 : node3475;
										assign node3475 = (inp[11]) ? node3477 : 3'b011;
											assign node3477 = (inp[3]) ? 3'b011 : 3'b000;
										assign node3480 = (inp[3]) ? 3'b001 : node3481;
											assign node3481 = (inp[5]) ? 3'b001 : 3'b011;
						assign node3485 = (inp[7]) ? node3551 : node3486;
							assign node3486 = (inp[2]) ? node3528 : node3487;
								assign node3487 = (inp[3]) ? node3507 : node3488;
									assign node3488 = (inp[4]) ? node3494 : node3489;
										assign node3489 = (inp[8]) ? node3491 : 3'b010;
											assign node3491 = (inp[5]) ? 3'b010 : 3'b000;
										assign node3494 = (inp[11]) ? node3500 : node3495;
											assign node3495 = (inp[8]) ? node3497 : 3'b000;
												assign node3497 = (inp[5]) ? 3'b000 : 3'b010;
											assign node3500 = (inp[5]) ? node3504 : node3501;
												assign node3501 = (inp[8]) ? 3'b010 : 3'b000;
												assign node3504 = (inp[8]) ? 3'b000 : 3'b010;
									assign node3507 = (inp[5]) ? node3521 : node3508;
										assign node3508 = (inp[11]) ? node3516 : node3509;
											assign node3509 = (inp[8]) ? node3513 : node3510;
												assign node3510 = (inp[4]) ? 3'b010 : 3'b000;
												assign node3513 = (inp[4]) ? 3'b000 : 3'b010;
											assign node3516 = (inp[8]) ? 3'b000 : node3517;
												assign node3517 = (inp[4]) ? 3'b010 : 3'b000;
										assign node3521 = (inp[8]) ? node3525 : node3522;
											assign node3522 = (inp[4]) ? 3'b010 : 3'b000;
											assign node3525 = (inp[4]) ? 3'b000 : 3'b010;
								assign node3528 = (inp[8]) ? node3540 : node3529;
									assign node3529 = (inp[4]) ? node3535 : node3530;
										assign node3530 = (inp[3]) ? 3'b000 : node3531;
											assign node3531 = (inp[5]) ? 3'b000 : 3'b010;
										assign node3535 = (inp[5]) ? 3'b011 : node3536;
											assign node3536 = (inp[3]) ? 3'b011 : 3'b000;
									assign node3540 = (inp[4]) ? node3546 : node3541;
										assign node3541 = (inp[3]) ? 3'b011 : node3542;
											assign node3542 = (inp[5]) ? 3'b011 : 3'b000;
										assign node3546 = (inp[5]) ? 3'b001 : node3547;
											assign node3547 = (inp[3]) ? 3'b001 : 3'b011;
							assign node3551 = (inp[2]) ? node3575 : node3552;
								assign node3552 = (inp[8]) ? node3564 : node3553;
									assign node3553 = (inp[4]) ? node3559 : node3554;
										assign node3554 = (inp[3]) ? 3'b001 : node3555;
											assign node3555 = (inp[5]) ? 3'b001 : 3'b011;
										assign node3559 = (inp[3]) ? 3'b011 : node3560;
											assign node3560 = (inp[5]) ? 3'b011 : 3'b001;
									assign node3564 = (inp[4]) ? node3570 : node3565;
										assign node3565 = (inp[5]) ? 3'b011 : node3566;
											assign node3566 = (inp[3]) ? 3'b011 : 3'b001;
										assign node3570 = (inp[3]) ? 3'b001 : node3571;
											assign node3571 = (inp[5]) ? 3'b001 : 3'b011;
								assign node3575 = (inp[8]) ? node3585 : node3576;
									assign node3576 = (inp[5]) ? node3582 : node3577;
										assign node3577 = (inp[4]) ? 3'b001 : node3578;
											assign node3578 = (inp[3]) ? 3'b001 : 3'b011;
										assign node3582 = (inp[4]) ? 3'b010 : 3'b001;
									assign node3585 = (inp[4]) ? node3591 : node3586;
										assign node3586 = (inp[3]) ? 3'b010 : node3587;
											assign node3587 = (inp[5]) ? 3'b010 : 3'b001;
										assign node3591 = (inp[3]) ? 3'b000 : 3'b010;
					assign node3594 = (inp[5]) ? node3742 : node3595;
						assign node3595 = (inp[2]) ? node3653 : node3596;
							assign node3596 = (inp[9]) ? node3624 : node3597;
								assign node3597 = (inp[7]) ? node3609 : node3598;
									assign node3598 = (inp[4]) ? node3604 : node3599;
										assign node3599 = (inp[3]) ? 3'b010 : node3600;
											assign node3600 = (inp[8]) ? 3'b001 : 3'b011;
										assign node3604 = (inp[8]) ? node3606 : 3'b010;
											assign node3606 = (inp[3]) ? 3'b000 : 3'b010;
									assign node3609 = (inp[3]) ? node3617 : node3610;
										assign node3610 = (inp[4]) ? node3614 : node3611;
											assign node3611 = (inp[8]) ? 3'b000 : 3'b010;
											assign node3614 = (inp[8]) ? 3'b011 : 3'b000;
										assign node3617 = (inp[11]) ? 3'b011 : node3618;
											assign node3618 = (inp[8]) ? node3620 : 3'b011;
												assign node3620 = (inp[4]) ? 3'b001 : 3'b011;
								assign node3624 = (inp[8]) ? node3638 : node3625;
									assign node3625 = (inp[7]) ? node3633 : node3626;
										assign node3626 = (inp[11]) ? 3'b000 : node3627;
											assign node3627 = (inp[3]) ? 3'b011 : node3628;
												assign node3628 = (inp[4]) ? 3'b000 : 3'b010;
										assign node3633 = (inp[3]) ? node3635 : 3'b001;
											assign node3635 = (inp[4]) ? 3'b010 : 3'b001;
									assign node3638 = (inp[7]) ? node3648 : node3639;
										assign node3639 = (inp[11]) ? node3641 : 3'b011;
											assign node3641 = (inp[4]) ? node3645 : node3642;
												assign node3642 = (inp[3]) ? 3'b011 : 3'b000;
												assign node3645 = (inp[3]) ? 3'b001 : 3'b011;
										assign node3648 = (inp[3]) ? node3650 : 3'b010;
											assign node3650 = (inp[4]) ? 3'b000 : 3'b010;
							assign node3653 = (inp[8]) ? node3695 : node3654;
								assign node3654 = (inp[11]) ? node3680 : node3655;
									assign node3655 = (inp[9]) ? node3667 : node3656;
										assign node3656 = (inp[7]) ? node3662 : node3657;
											assign node3657 = (inp[4]) ? 3'b000 : node3658;
												assign node3658 = (inp[3]) ? 3'b000 : 3'b010;
											assign node3662 = (inp[3]) ? node3664 : 3'b001;
												assign node3664 = (inp[4]) ? 3'b011 : 3'b001;
										assign node3667 = (inp[7]) ? node3675 : node3668;
											assign node3668 = (inp[3]) ? node3672 : node3669;
												assign node3669 = (inp[4]) ? 3'b001 : 3'b011;
												assign node3672 = (inp[4]) ? 3'b011 : 3'b001;
											assign node3675 = (inp[3]) ? node3677 : 3'b010;
												assign node3677 = (inp[4]) ? 3'b010 : 3'b000;
									assign node3680 = (inp[7]) ? node3684 : node3681;
										assign node3681 = (inp[9]) ? 3'b011 : 3'b010;
										assign node3684 = (inp[9]) ? node3692 : node3685;
											assign node3685 = (inp[4]) ? node3689 : node3686;
												assign node3686 = (inp[3]) ? 3'b001 : 3'b011;
												assign node3689 = (inp[3]) ? 3'b011 : 3'b001;
											assign node3692 = (inp[4]) ? 3'b010 : 3'b000;
								assign node3695 = (inp[3]) ? node3719 : node3696;
									assign node3696 = (inp[4]) ? node3704 : node3697;
										assign node3697 = (inp[9]) ? node3701 : node3698;
											assign node3698 = (inp[7]) ? 3'b001 : 3'b000;
											assign node3701 = (inp[7]) ? 3'b000 : 3'b001;
										assign node3704 = (inp[11]) ? node3712 : node3705;
											assign node3705 = (inp[9]) ? node3709 : node3706;
												assign node3706 = (inp[7]) ? 3'b011 : 3'b010;
												assign node3709 = (inp[7]) ? 3'b010 : 3'b011;
											assign node3712 = (inp[7]) ? node3716 : node3713;
												assign node3713 = (inp[9]) ? 3'b011 : 3'b010;
												assign node3716 = (inp[9]) ? 3'b010 : 3'b011;
									assign node3719 = (inp[4]) ? node3727 : node3720;
										assign node3720 = (inp[9]) ? node3724 : node3721;
											assign node3721 = (inp[7]) ? 3'b011 : 3'b010;
											assign node3724 = (inp[7]) ? 3'b010 : 3'b011;
										assign node3727 = (inp[11]) ? node3735 : node3728;
											assign node3728 = (inp[7]) ? node3732 : node3729;
												assign node3729 = (inp[9]) ? 3'b001 : 3'b000;
												assign node3732 = (inp[9]) ? 3'b000 : 3'b001;
											assign node3735 = (inp[7]) ? node3739 : node3736;
												assign node3736 = (inp[9]) ? 3'b001 : 3'b000;
												assign node3739 = (inp[9]) ? 3'b000 : 3'b001;
						assign node3742 = (inp[2]) ? node3774 : node3743;
							assign node3743 = (inp[7]) ? node3759 : node3744;
								assign node3744 = (inp[9]) ? node3752 : node3745;
									assign node3745 = (inp[8]) ? node3749 : node3746;
										assign node3746 = (inp[4]) ? 3'b010 : 3'b001;
										assign node3749 = (inp[4]) ? 3'b000 : 3'b010;
									assign node3752 = (inp[8]) ? node3756 : node3753;
										assign node3753 = (inp[4]) ? 3'b011 : 3'b000;
										assign node3756 = (inp[4]) ? 3'b001 : 3'b011;
								assign node3759 = (inp[9]) ? node3767 : node3760;
									assign node3760 = (inp[8]) ? node3764 : node3761;
										assign node3761 = (inp[4]) ? 3'b011 : 3'b000;
										assign node3764 = (inp[4]) ? 3'b001 : 3'b011;
									assign node3767 = (inp[8]) ? node3771 : node3768;
										assign node3768 = (inp[4]) ? 3'b010 : 3'b001;
										assign node3771 = (inp[4]) ? 3'b000 : 3'b010;
							assign node3774 = (inp[7]) ? node3806 : node3775;
								assign node3775 = (inp[9]) ? node3791 : node3776;
									assign node3776 = (inp[3]) ? node3786 : node3777;
										assign node3777 = (inp[11]) ? node3781 : node3778;
											assign node3778 = (inp[8]) ? 3'b010 : 3'b000;
											assign node3781 = (inp[4]) ? node3783 : 3'b000;
												assign node3783 = (inp[8]) ? 3'b000 : 3'b010;
										assign node3786 = (inp[8]) ? 3'b010 : node3787;
											assign node3787 = (inp[4]) ? 3'b010 : 3'b000;
									assign node3791 = (inp[11]) ? node3799 : node3792;
										assign node3792 = (inp[4]) ? node3796 : node3793;
											assign node3793 = (inp[8]) ? 3'b011 : 3'b001;
											assign node3796 = (inp[8]) ? 3'b001 : 3'b011;
										assign node3799 = (inp[4]) ? node3803 : node3800;
											assign node3800 = (inp[8]) ? 3'b011 : 3'b001;
											assign node3803 = (inp[8]) ? 3'b001 : 3'b011;
								assign node3806 = (inp[9]) ? node3814 : node3807;
									assign node3807 = (inp[8]) ? node3811 : node3808;
										assign node3808 = (inp[4]) ? 3'b011 : 3'b001;
										assign node3811 = (inp[4]) ? 3'b001 : 3'b011;
									assign node3814 = (inp[11]) ? node3820 : node3815;
										assign node3815 = (inp[4]) ? node3817 : 3'b010;
											assign node3817 = (inp[8]) ? 3'b000 : 3'b010;
										assign node3820 = (inp[8]) ? node3824 : node3821;
											assign node3821 = (inp[4]) ? 3'b010 : 3'b000;
											assign node3824 = (inp[4]) ? 3'b000 : 3'b010;

endmodule