module dtc_split33_bm30 (
	input  wire [14-1:0] inp,
	output wire [8-1:0] outp
);

	wire [8-1:0] node1;
	wire [8-1:0] node2;
	wire [8-1:0] node3;
	wire [8-1:0] node4;
	wire [8-1:0] node5;
	wire [8-1:0] node6;
	wire [8-1:0] node7;
	wire [8-1:0] node9;
	wire [8-1:0] node10;
	wire [8-1:0] node14;
	wire [8-1:0] node15;
	wire [8-1:0] node16;
	wire [8-1:0] node20;
	wire [8-1:0] node21;
	wire [8-1:0] node23;
	wire [8-1:0] node26;
	wire [8-1:0] node28;
	wire [8-1:0] node31;
	wire [8-1:0] node32;
	wire [8-1:0] node33;
	wire [8-1:0] node34;
	wire [8-1:0] node38;
	wire [8-1:0] node40;
	wire [8-1:0] node41;
	wire [8-1:0] node44;
	wire [8-1:0] node47;
	wire [8-1:0] node48;
	wire [8-1:0] node50;
	wire [8-1:0] node51;
	wire [8-1:0] node54;
	wire [8-1:0] node57;
	wire [8-1:0] node59;
	wire [8-1:0] node60;
	wire [8-1:0] node61;
	wire [8-1:0] node64;
	wire [8-1:0] node67;
	wire [8-1:0] node68;
	wire [8-1:0] node71;
	wire [8-1:0] node74;
	wire [8-1:0] node75;
	wire [8-1:0] node76;
	wire [8-1:0] node77;
	wire [8-1:0] node79;
	wire [8-1:0] node82;
	wire [8-1:0] node83;
	wire [8-1:0] node84;
	wire [8-1:0] node88;
	wire [8-1:0] node90;
	wire [8-1:0] node93;
	wire [8-1:0] node94;
	wire [8-1:0] node95;
	wire [8-1:0] node96;
	wire [8-1:0] node97;
	wire [8-1:0] node102;
	wire [8-1:0] node103;
	wire [8-1:0] node104;
	wire [8-1:0] node108;
	wire [8-1:0] node111;
	wire [8-1:0] node112;
	wire [8-1:0] node113;
	wire [8-1:0] node116;
	wire [8-1:0] node117;
	wire [8-1:0] node123;
	wire [8-1:0] node124;
	wire [8-1:0] node125;
	wire [8-1:0] node126;
	wire [8-1:0] node129;
	wire [8-1:0] node130;
	wire [8-1:0] node131;
	wire [8-1:0] node132;
	wire [8-1:0] node136;
	wire [8-1:0] node139;
	wire [8-1:0] node141;
	wire [8-1:0] node142;
	wire [8-1:0] node146;
	wire [8-1:0] node147;
	wire [8-1:0] node148;
	wire [8-1:0] node149;
	wire [8-1:0] node151;
	wire [8-1:0] node154;
	wire [8-1:0] node156;
	wire [8-1:0] node159;
	wire [8-1:0] node160;
	wire [8-1:0] node162;
	wire [8-1:0] node163;
	wire [8-1:0] node167;
	wire [8-1:0] node168;
	wire [8-1:0] node169;
	wire [8-1:0] node174;
	wire [8-1:0] node175;
	wire [8-1:0] node176;
	wire [8-1:0] node178;
	wire [8-1:0] node181;
	wire [8-1:0] node183;
	wire [8-1:0] node186;
	wire [8-1:0] node187;
	wire [8-1:0] node189;
	wire [8-1:0] node192;
	wire [8-1:0] node193;
	wire [8-1:0] node194;
	wire [8-1:0] node197;
	wire [8-1:0] node201;
	wire [8-1:0] node202;
	wire [8-1:0] node203;
	wire [8-1:0] node204;
	wire [8-1:0] node205;
	wire [8-1:0] node208;
	wire [8-1:0] node211;
	wire [8-1:0] node212;
	wire [8-1:0] node215;
	wire [8-1:0] node218;
	wire [8-1:0] node219;
	wire [8-1:0] node220;
	wire [8-1:0] node221;
	wire [8-1:0] node224;
	wire [8-1:0] node227;
	wire [8-1:0] node228;
	wire [8-1:0] node229;
	wire [8-1:0] node233;
	wire [8-1:0] node234;
	wire [8-1:0] node237;
	wire [8-1:0] node240;
	wire [8-1:0] node241;
	wire [8-1:0] node243;
	wire [8-1:0] node244;
	wire [8-1:0] node248;
	wire [8-1:0] node249;
	wire [8-1:0] node251;
	wire [8-1:0] node254;
	wire [8-1:0] node255;
	wire [8-1:0] node258;
	wire [8-1:0] node260;
	wire [8-1:0] node263;
	wire [8-1:0] node264;
	wire [8-1:0] node265;
	wire [8-1:0] node266;
	wire [8-1:0] node267;
	wire [8-1:0] node271;
	wire [8-1:0] node272;
	wire [8-1:0] node273;
	wire [8-1:0] node276;
	wire [8-1:0] node280;
	wire [8-1:0] node281;
	wire [8-1:0] node282;
	wire [8-1:0] node286;
	wire [8-1:0] node287;
	wire [8-1:0] node291;
	wire [8-1:0] node292;
	wire [8-1:0] node293;
	wire [8-1:0] node294;
	wire [8-1:0] node295;
	wire [8-1:0] node298;
	wire [8-1:0] node301;
	wire [8-1:0] node304;
	wire [8-1:0] node305;
	wire [8-1:0] node306;
	wire [8-1:0] node310;
	wire [8-1:0] node311;
	wire [8-1:0] node315;
	wire [8-1:0] node316;
	wire [8-1:0] node317;
	wire [8-1:0] node319;
	wire [8-1:0] node320;
	wire [8-1:0] node321;
	wire [8-1:0] node326;
	wire [8-1:0] node329;
	wire [8-1:0] node332;
	wire [8-1:0] node333;
	wire [8-1:0] node334;
	wire [8-1:0] node335;
	wire [8-1:0] node336;
	wire [8-1:0] node337;
	wire [8-1:0] node338;
	wire [8-1:0] node339;
	wire [8-1:0] node342;
	wire [8-1:0] node345;
	wire [8-1:0] node346;
	wire [8-1:0] node349;
	wire [8-1:0] node350;
	wire [8-1:0] node354;
	wire [8-1:0] node355;
	wire [8-1:0] node356;
	wire [8-1:0] node357;
	wire [8-1:0] node361;
	wire [8-1:0] node362;
	wire [8-1:0] node364;
	wire [8-1:0] node366;
	wire [8-1:0] node370;
	wire [8-1:0] node372;
	wire [8-1:0] node373;
	wire [8-1:0] node374;
	wire [8-1:0] node375;
	wire [8-1:0] node379;
	wire [8-1:0] node383;
	wire [8-1:0] node384;
	wire [8-1:0] node386;
	wire [8-1:0] node387;
	wire [8-1:0] node391;
	wire [8-1:0] node392;
	wire [8-1:0] node395;
	wire [8-1:0] node398;
	wire [8-1:0] node399;
	wire [8-1:0] node400;
	wire [8-1:0] node401;
	wire [8-1:0] node402;
	wire [8-1:0] node403;
	wire [8-1:0] node406;
	wire [8-1:0] node410;
	wire [8-1:0] node411;
	wire [8-1:0] node415;
	wire [8-1:0] node416;
	wire [8-1:0] node420;
	wire [8-1:0] node421;
	wire [8-1:0] node422;
	wire [8-1:0] node423;
	wire [8-1:0] node424;
	wire [8-1:0] node427;
	wire [8-1:0] node430;
	wire [8-1:0] node432;
	wire [8-1:0] node433;
	wire [8-1:0] node437;
	wire [8-1:0] node438;
	wire [8-1:0] node439;
	wire [8-1:0] node441;
	wire [8-1:0] node446;
	wire [8-1:0] node447;
	wire [8-1:0] node448;
	wire [8-1:0] node450;
	wire [8-1:0] node452;
	wire [8-1:0] node454;
	wire [8-1:0] node457;
	wire [8-1:0] node458;
	wire [8-1:0] node461;
	wire [8-1:0] node463;
	wire [8-1:0] node466;
	wire [8-1:0] node467;
	wire [8-1:0] node470;
	wire [8-1:0] node472;
	wire [8-1:0] node475;
	wire [8-1:0] node476;
	wire [8-1:0] node477;
	wire [8-1:0] node478;
	wire [8-1:0] node479;
	wire [8-1:0] node480;
	wire [8-1:0] node481;
	wire [8-1:0] node483;
	wire [8-1:0] node487;
	wire [8-1:0] node488;
	wire [8-1:0] node490;
	wire [8-1:0] node493;
	wire [8-1:0] node496;
	wire [8-1:0] node497;
	wire [8-1:0] node500;
	wire [8-1:0] node501;
	wire [8-1:0] node502;
	wire [8-1:0] node505;
	wire [8-1:0] node508;
	wire [8-1:0] node511;
	wire [8-1:0] node512;
	wire [8-1:0] node513;
	wire [8-1:0] node515;
	wire [8-1:0] node518;
	wire [8-1:0] node520;
	wire [8-1:0] node521;
	wire [8-1:0] node525;
	wire [8-1:0] node526;
	wire [8-1:0] node528;
	wire [8-1:0] node529;
	wire [8-1:0] node533;
	wire [8-1:0] node535;
	wire [8-1:0] node538;
	wire [8-1:0] node539;
	wire [8-1:0] node540;
	wire [8-1:0] node541;
	wire [8-1:0] node543;
	wire [8-1:0] node545;
	wire [8-1:0] node548;
	wire [8-1:0] node551;
	wire [8-1:0] node552;
	wire [8-1:0] node554;
	wire [8-1:0] node557;
	wire [8-1:0] node559;
	wire [8-1:0] node562;
	wire [8-1:0] node563;
	wire [8-1:0] node564;
	wire [8-1:0] node565;
	wire [8-1:0] node566;
	wire [8-1:0] node567;
	wire [8-1:0] node572;
	wire [8-1:0] node573;
	wire [8-1:0] node577;
	wire [8-1:0] node579;
	wire [8-1:0] node582;
	wire [8-1:0] node583;
	wire [8-1:0] node584;
	wire [8-1:0] node585;
	wire [8-1:0] node588;
	wire [8-1:0] node592;
	wire [8-1:0] node593;
	wire [8-1:0] node596;
	wire [8-1:0] node599;
	wire [8-1:0] node600;
	wire [8-1:0] node601;
	wire [8-1:0] node602;
	wire [8-1:0] node603;
	wire [8-1:0] node604;
	wire [8-1:0] node605;
	wire [8-1:0] node608;
	wire [8-1:0] node611;
	wire [8-1:0] node614;
	wire [8-1:0] node616;
	wire [8-1:0] node619;
	wire [8-1:0] node620;
	wire [8-1:0] node621;
	wire [8-1:0] node625;
	wire [8-1:0] node626;
	wire [8-1:0] node627;
	wire [8-1:0] node631;
	wire [8-1:0] node633;
	wire [8-1:0] node634;
	wire [8-1:0] node638;
	wire [8-1:0] node639;
	wire [8-1:0] node640;
	wire [8-1:0] node642;
	wire [8-1:0] node646;
	wire [8-1:0] node647;
	wire [8-1:0] node650;
	wire [8-1:0] node651;
	wire [8-1:0] node655;
	wire [8-1:0] node656;
	wire [8-1:0] node657;
	wire [8-1:0] node658;
	wire [8-1:0] node659;
	wire [8-1:0] node661;
	wire [8-1:0] node662;
	wire [8-1:0] node667;
	wire [8-1:0] node668;
	wire [8-1:0] node671;
	wire [8-1:0] node674;
	wire [8-1:0] node675;
	wire [8-1:0] node676;
	wire [8-1:0] node677;
	wire [8-1:0] node679;
	wire [8-1:0] node684;
	wire [8-1:0] node685;
	wire [8-1:0] node687;
	wire [8-1:0] node691;
	wire [8-1:0] node692;
	wire [8-1:0] node693;
	wire [8-1:0] node694;
	wire [8-1:0] node697;
	wire [8-1:0] node700;
	wire [8-1:0] node701;
	wire [8-1:0] node703;
	wire [8-1:0] node704;
	wire [8-1:0] node708;
	wire [8-1:0] node709;
	wire [8-1:0] node713;
	wire [8-1:0] node714;
	wire [8-1:0] node716;
	wire [8-1:0] node719;
	wire [8-1:0] node721;
	wire [8-1:0] node724;
	wire [8-1:0] node725;
	wire [8-1:0] node726;
	wire [8-1:0] node727;
	wire [8-1:0] node728;
	wire [8-1:0] node729;
	wire [8-1:0] node730;
	wire [8-1:0] node732;
	wire [8-1:0] node735;
	wire [8-1:0] node736;
	wire [8-1:0] node740;
	wire [8-1:0] node742;
	wire [8-1:0] node744;
	wire [8-1:0] node747;
	wire [8-1:0] node748;
	wire [8-1:0] node749;
	wire [8-1:0] node751;
	wire [8-1:0] node755;
	wire [8-1:0] node757;
	wire [8-1:0] node759;
	wire [8-1:0] node762;
	wire [8-1:0] node763;
	wire [8-1:0] node764;
	wire [8-1:0] node765;
	wire [8-1:0] node768;
	wire [8-1:0] node770;
	wire [8-1:0] node772;
	wire [8-1:0] node775;
	wire [8-1:0] node777;
	wire [8-1:0] node779;
	wire [8-1:0] node782;
	wire [8-1:0] node783;
	wire [8-1:0] node784;
	wire [8-1:0] node785;
	wire [8-1:0] node789;
	wire [8-1:0] node790;
	wire [8-1:0] node793;
	wire [8-1:0] node796;
	wire [8-1:0] node797;
	wire [8-1:0] node799;
	wire [8-1:0] node802;
	wire [8-1:0] node805;
	wire [8-1:0] node806;
	wire [8-1:0] node807;
	wire [8-1:0] node808;
	wire [8-1:0] node809;
	wire [8-1:0] node811;
	wire [8-1:0] node814;
	wire [8-1:0] node816;
	wire [8-1:0] node819;
	wire [8-1:0] node820;
	wire [8-1:0] node821;
	wire [8-1:0] node825;
	wire [8-1:0] node827;
	wire [8-1:0] node830;
	wire [8-1:0] node831;
	wire [8-1:0] node832;
	wire [8-1:0] node833;
	wire [8-1:0] node836;
	wire [8-1:0] node839;
	wire [8-1:0] node840;
	wire [8-1:0] node844;
	wire [8-1:0] node845;
	wire [8-1:0] node847;
	wire [8-1:0] node851;
	wire [8-1:0] node852;
	wire [8-1:0] node853;
	wire [8-1:0] node854;
	wire [8-1:0] node856;
	wire [8-1:0] node859;
	wire [8-1:0] node860;
	wire [8-1:0] node864;
	wire [8-1:0] node865;
	wire [8-1:0] node866;
	wire [8-1:0] node870;
	wire [8-1:0] node872;
	wire [8-1:0] node875;
	wire [8-1:0] node876;
	wire [8-1:0] node877;
	wire [8-1:0] node880;
	wire [8-1:0] node882;
	wire [8-1:0] node885;
	wire [8-1:0] node886;
	wire [8-1:0] node887;
	wire [8-1:0] node891;
	wire [8-1:0] node892;
	wire [8-1:0] node895;
	wire [8-1:0] node898;
	wire [8-1:0] node899;
	wire [8-1:0] node900;
	wire [8-1:0] node901;
	wire [8-1:0] node902;
	wire [8-1:0] node903;
	wire [8-1:0] node907;
	wire [8-1:0] node908;
	wire [8-1:0] node909;
	wire [8-1:0] node910;
	wire [8-1:0] node916;
	wire [8-1:0] node917;
	wire [8-1:0] node918;
	wire [8-1:0] node919;
	wire [8-1:0] node923;
	wire [8-1:0] node926;
	wire [8-1:0] node927;
	wire [8-1:0] node931;
	wire [8-1:0] node932;
	wire [8-1:0] node933;
	wire [8-1:0] node934;
	wire [8-1:0] node936;
	wire [8-1:0] node937;
	wire [8-1:0] node941;
	wire [8-1:0] node942;
	wire [8-1:0] node945;
	wire [8-1:0] node948;
	wire [8-1:0] node949;
	wire [8-1:0] node950;
	wire [8-1:0] node954;
	wire [8-1:0] node956;
	wire [8-1:0] node957;
	wire [8-1:0] node960;
	wire [8-1:0] node963;
	wire [8-1:0] node964;
	wire [8-1:0] node965;
	wire [8-1:0] node966;
	wire [8-1:0] node970;
	wire [8-1:0] node971;
	wire [8-1:0] node974;
	wire [8-1:0] node977;
	wire [8-1:0] node978;
	wire [8-1:0] node979;
	wire [8-1:0] node980;
	wire [8-1:0] node984;
	wire [8-1:0] node987;
	wire [8-1:0] node989;
	wire [8-1:0] node991;
	wire [8-1:0] node994;
	wire [8-1:0] node995;
	wire [8-1:0] node996;
	wire [8-1:0] node997;
	wire [8-1:0] node998;
	wire [8-1:0] node999;
	wire [8-1:0] node1000;
	wire [8-1:0] node1005;
	wire [8-1:0] node1008;
	wire [8-1:0] node1009;
	wire [8-1:0] node1011;
	wire [8-1:0] node1014;
	wire [8-1:0] node1015;
	wire [8-1:0] node1019;
	wire [8-1:0] node1020;
	wire [8-1:0] node1021;
	wire [8-1:0] node1022;
	wire [8-1:0] node1026;
	wire [8-1:0] node1028;
	wire [8-1:0] node1031;
	wire [8-1:0] node1032;
	wire [8-1:0] node1035;
	wire [8-1:0] node1038;
	wire [8-1:0] node1039;
	wire [8-1:0] node1040;
	wire [8-1:0] node1041;
	wire [8-1:0] node1042;
	wire [8-1:0] node1045;
	wire [8-1:0] node1048;
	wire [8-1:0] node1049;
	wire [8-1:0] node1050;
	wire [8-1:0] node1054;
	wire [8-1:0] node1057;
	wire [8-1:0] node1058;
	wire [8-1:0] node1059;
	wire [8-1:0] node1063;
	wire [8-1:0] node1064;
	wire [8-1:0] node1066;
	wire [8-1:0] node1069;
	wire [8-1:0] node1070;
	wire [8-1:0] node1074;
	wire [8-1:0] node1075;
	wire [8-1:0] node1076;
	wire [8-1:0] node1077;
	wire [8-1:0] node1079;
	wire [8-1:0] node1082;
	wire [8-1:0] node1085;
	wire [8-1:0] node1086;
	wire [8-1:0] node1089;
	wire [8-1:0] node1090;
	wire [8-1:0] node1094;
	wire [8-1:0] node1095;
	wire [8-1:0] node1096;
	wire [8-1:0] node1099;
	wire [8-1:0] node1102;
	wire [8-1:0] node1105;
	wire [8-1:0] node1106;
	wire [8-1:0] node1107;
	wire [8-1:0] node1108;
	wire [8-1:0] node1109;
	wire [8-1:0] node1110;
	wire [8-1:0] node1111;
	wire [8-1:0] node1112;
	wire [8-1:0] node1115;
	wire [8-1:0] node1118;
	wire [8-1:0] node1121;
	wire [8-1:0] node1122;
	wire [8-1:0] node1123;
	wire [8-1:0] node1127;
	wire [8-1:0] node1129;
	wire [8-1:0] node1132;
	wire [8-1:0] node1133;
	wire [8-1:0] node1134;
	wire [8-1:0] node1135;
	wire [8-1:0] node1136;
	wire [8-1:0] node1137;
	wire [8-1:0] node1141;
	wire [8-1:0] node1142;
	wire [8-1:0] node1147;
	wire [8-1:0] node1148;
	wire [8-1:0] node1149;
	wire [8-1:0] node1150;
	wire [8-1:0] node1153;
	wire [8-1:0] node1157;
	wire [8-1:0] node1160;
	wire [8-1:0] node1161;
	wire [8-1:0] node1162;
	wire [8-1:0] node1163;
	wire [8-1:0] node1167;
	wire [8-1:0] node1168;
	wire [8-1:0] node1170;
	wire [8-1:0] node1174;
	wire [8-1:0] node1175;
	wire [8-1:0] node1176;
	wire [8-1:0] node1177;
	wire [8-1:0] node1181;
	wire [8-1:0] node1184;
	wire [8-1:0] node1185;
	wire [8-1:0] node1189;
	wire [8-1:0] node1190;
	wire [8-1:0] node1191;
	wire [8-1:0] node1192;
	wire [8-1:0] node1194;
	wire [8-1:0] node1197;
	wire [8-1:0] node1199;
	wire [8-1:0] node1202;
	wire [8-1:0] node1203;
	wire [8-1:0] node1204;
	wire [8-1:0] node1205;
	wire [8-1:0] node1209;
	wire [8-1:0] node1210;
	wire [8-1:0] node1213;
	wire [8-1:0] node1216;
	wire [8-1:0] node1217;
	wire [8-1:0] node1218;
	wire [8-1:0] node1221;
	wire [8-1:0] node1224;
	wire [8-1:0] node1225;
	wire [8-1:0] node1226;
	wire [8-1:0] node1230;
	wire [8-1:0] node1233;
	wire [8-1:0] node1234;
	wire [8-1:0] node1235;
	wire [8-1:0] node1236;
	wire [8-1:0] node1238;
	wire [8-1:0] node1242;
	wire [8-1:0] node1243;
	wire [8-1:0] node1245;
	wire [8-1:0] node1249;
	wire [8-1:0] node1250;
	wire [8-1:0] node1252;
	wire [8-1:0] node1256;
	wire [8-1:0] node1257;
	wire [8-1:0] node1258;
	wire [8-1:0] node1259;
	wire [8-1:0] node1260;
	wire [8-1:0] node1261;
	wire [8-1:0] node1263;
	wire [8-1:0] node1264;
	wire [8-1:0] node1266;
	wire [8-1:0] node1270;
	wire [8-1:0] node1272;
	wire [8-1:0] node1274;
	wire [8-1:0] node1277;
	wire [8-1:0] node1278;
	wire [8-1:0] node1279;
	wire [8-1:0] node1282;
	wire [8-1:0] node1284;
	wire [8-1:0] node1287;
	wire [8-1:0] node1288;
	wire [8-1:0] node1289;
	wire [8-1:0] node1293;
	wire [8-1:0] node1296;
	wire [8-1:0] node1297;
	wire [8-1:0] node1298;
	wire [8-1:0] node1299;
	wire [8-1:0] node1302;
	wire [8-1:0] node1304;
	wire [8-1:0] node1307;
	wire [8-1:0] node1308;
	wire [8-1:0] node1310;
	wire [8-1:0] node1313;
	wire [8-1:0] node1315;
	wire [8-1:0] node1316;
	wire [8-1:0] node1320;
	wire [8-1:0] node1321;
	wire [8-1:0] node1322;
	wire [8-1:0] node1325;
	wire [8-1:0] node1328;
	wire [8-1:0] node1329;
	wire [8-1:0] node1333;
	wire [8-1:0] node1334;
	wire [8-1:0] node1335;
	wire [8-1:0] node1336;
	wire [8-1:0] node1337;
	wire [8-1:0] node1340;
	wire [8-1:0] node1343;
	wire [8-1:0] node1344;
	wire [8-1:0] node1346;
	wire [8-1:0] node1349;
	wire [8-1:0] node1350;
	wire [8-1:0] node1353;
	wire [8-1:0] node1356;
	wire [8-1:0] node1357;
	wire [8-1:0] node1359;
	wire [8-1:0] node1360;
	wire [8-1:0] node1364;
	wire [8-1:0] node1365;
	wire [8-1:0] node1366;
	wire [8-1:0] node1369;
	wire [8-1:0] node1372;
	wire [8-1:0] node1373;
	wire [8-1:0] node1375;
	wire [8-1:0] node1378;
	wire [8-1:0] node1379;
	wire [8-1:0] node1382;
	wire [8-1:0] node1385;
	wire [8-1:0] node1386;
	wire [8-1:0] node1387;
	wire [8-1:0] node1388;
	wire [8-1:0] node1389;
	wire [8-1:0] node1392;
	wire [8-1:0] node1396;
	wire [8-1:0] node1397;
	wire [8-1:0] node1399;
	wire [8-1:0] node1400;
	wire [8-1:0] node1404;
	wire [8-1:0] node1406;
	wire [8-1:0] node1407;
	wire [8-1:0] node1410;
	wire [8-1:0] node1411;
	wire [8-1:0] node1415;
	wire [8-1:0] node1416;
	wire [8-1:0] node1417;
	wire [8-1:0] node1418;
	wire [8-1:0] node1422;
	wire [8-1:0] node1423;
	wire [8-1:0] node1426;
	wire [8-1:0] node1428;
	wire [8-1:0] node1431;
	wire [8-1:0] node1432;
	wire [8-1:0] node1433;
	wire [8-1:0] node1434;
	wire [8-1:0] node1437;
	wire [8-1:0] node1440;
	wire [8-1:0] node1441;
	wire [8-1:0] node1445;
	wire [8-1:0] node1446;
	wire [8-1:0] node1449;
	wire [8-1:0] node1452;
	wire [8-1:0] node1453;
	wire [8-1:0] node1454;
	wire [8-1:0] node1455;
	wire [8-1:0] node1456;
	wire [8-1:0] node1458;
	wire [8-1:0] node1461;
	wire [8-1:0] node1462;
	wire [8-1:0] node1464;
	wire [8-1:0] node1468;
	wire [8-1:0] node1469;
	wire [8-1:0] node1470;
	wire [8-1:0] node1473;
	wire [8-1:0] node1476;
	wire [8-1:0] node1477;
	wire [8-1:0] node1480;
	wire [8-1:0] node1481;
	wire [8-1:0] node1484;
	wire [8-1:0] node1485;
	wire [8-1:0] node1489;
	wire [8-1:0] node1490;
	wire [8-1:0] node1491;
	wire [8-1:0] node1492;
	wire [8-1:0] node1494;
	wire [8-1:0] node1495;
	wire [8-1:0] node1499;
	wire [8-1:0] node1502;
	wire [8-1:0] node1503;
	wire [8-1:0] node1506;
	wire [8-1:0] node1507;
	wire [8-1:0] node1508;
	wire [8-1:0] node1513;
	wire [8-1:0] node1514;
	wire [8-1:0] node1515;
	wire [8-1:0] node1517;
	wire [8-1:0] node1518;
	wire [8-1:0] node1522;
	wire [8-1:0] node1523;
	wire [8-1:0] node1527;
	wire [8-1:0] node1528;
	wire [8-1:0] node1529;
	wire [8-1:0] node1532;
	wire [8-1:0] node1535;
	wire [8-1:0] node1536;
	wire [8-1:0] node1539;
	wire [8-1:0] node1542;
	wire [8-1:0] node1543;
	wire [8-1:0] node1544;
	wire [8-1:0] node1545;
	wire [8-1:0] node1546;
	wire [8-1:0] node1549;
	wire [8-1:0] node1550;
	wire [8-1:0] node1553;
	wire [8-1:0] node1556;
	wire [8-1:0] node1557;
	wire [8-1:0] node1558;
	wire [8-1:0] node1561;
	wire [8-1:0] node1564;
	wire [8-1:0] node1565;
	wire [8-1:0] node1569;
	wire [8-1:0] node1570;
	wire [8-1:0] node1571;
	wire [8-1:0] node1572;
	wire [8-1:0] node1576;
	wire [8-1:0] node1579;
	wire [8-1:0] node1580;
	wire [8-1:0] node1581;
	wire [8-1:0] node1582;
	wire [8-1:0] node1586;
	wire [8-1:0] node1587;
	wire [8-1:0] node1591;
	wire [8-1:0] node1594;
	wire [8-1:0] node1595;
	wire [8-1:0] node1596;
	wire [8-1:0] node1597;
	wire [8-1:0] node1598;
	wire [8-1:0] node1602;
	wire [8-1:0] node1604;
	wire [8-1:0] node1607;
	wire [8-1:0] node1608;
	wire [8-1:0] node1609;
	wire [8-1:0] node1612;
	wire [8-1:0] node1615;
	wire [8-1:0] node1616;
	wire [8-1:0] node1620;
	wire [8-1:0] node1621;
	wire [8-1:0] node1622;
	wire [8-1:0] node1624;
	wire [8-1:0] node1627;
	wire [8-1:0] node1629;
	wire [8-1:0] node1632;
	wire [8-1:0] node1633;
	wire [8-1:0] node1634;
	wire [8-1:0] node1637;
	wire [8-1:0] node1638;
	wire [8-1:0] node1641;
	wire [8-1:0] node1644;
	wire [8-1:0] node1645;
	wire [8-1:0] node1648;
	wire [8-1:0] node1651;
	wire [8-1:0] node1652;
	wire [8-1:0] node1653;
	wire [8-1:0] node1654;
	wire [8-1:0] node1655;
	wire [8-1:0] node1656;
	wire [8-1:0] node1657;
	wire [8-1:0] node1658;
	wire [8-1:0] node1659;
	wire [8-1:0] node1663;
	wire [8-1:0] node1664;
	wire [8-1:0] node1668;
	wire [8-1:0] node1670;
	wire [8-1:0] node1673;
	wire [8-1:0] node1674;
	wire [8-1:0] node1675;
	wire [8-1:0] node1678;
	wire [8-1:0] node1679;
	wire [8-1:0] node1680;
	wire [8-1:0] node1684;
	wire [8-1:0] node1687;
	wire [8-1:0] node1688;
	wire [8-1:0] node1690;
	wire [8-1:0] node1693;
	wire [8-1:0] node1694;
	wire [8-1:0] node1697;
	wire [8-1:0] node1700;
	wire [8-1:0] node1701;
	wire [8-1:0] node1702;
	wire [8-1:0] node1704;
	wire [8-1:0] node1706;
	wire [8-1:0] node1707;
	wire [8-1:0] node1711;
	wire [8-1:0] node1712;
	wire [8-1:0] node1714;
	wire [8-1:0] node1717;
	wire [8-1:0] node1718;
	wire [8-1:0] node1720;
	wire [8-1:0] node1723;
	wire [8-1:0] node1725;
	wire [8-1:0] node1728;
	wire [8-1:0] node1729;
	wire [8-1:0] node1730;
	wire [8-1:0] node1731;
	wire [8-1:0] node1735;
	wire [8-1:0] node1736;
	wire [8-1:0] node1738;
	wire [8-1:0] node1742;
	wire [8-1:0] node1743;
	wire [8-1:0] node1746;
	wire [8-1:0] node1747;
	wire [8-1:0] node1749;
	wire [8-1:0] node1753;
	wire [8-1:0] node1754;
	wire [8-1:0] node1755;
	wire [8-1:0] node1756;
	wire [8-1:0] node1758;
	wire [8-1:0] node1759;
	wire [8-1:0] node1762;
	wire [8-1:0] node1765;
	wire [8-1:0] node1766;
	wire [8-1:0] node1768;
	wire [8-1:0] node1771;
	wire [8-1:0] node1774;
	wire [8-1:0] node1775;
	wire [8-1:0] node1776;
	wire [8-1:0] node1780;
	wire [8-1:0] node1781;
	wire [8-1:0] node1782;
	wire [8-1:0] node1786;
	wire [8-1:0] node1787;
	wire [8-1:0] node1791;
	wire [8-1:0] node1792;
	wire [8-1:0] node1793;
	wire [8-1:0] node1794;
	wire [8-1:0] node1797;
	wire [8-1:0] node1798;
	wire [8-1:0] node1799;
	wire [8-1:0] node1802;
	wire [8-1:0] node1805;
	wire [8-1:0] node1807;
	wire [8-1:0] node1810;
	wire [8-1:0] node1811;
	wire [8-1:0] node1812;
	wire [8-1:0] node1814;
	wire [8-1:0] node1817;
	wire [8-1:0] node1820;
	wire [8-1:0] node1822;
	wire [8-1:0] node1825;
	wire [8-1:0] node1826;
	wire [8-1:0] node1827;
	wire [8-1:0] node1830;
	wire [8-1:0] node1832;
	wire [8-1:0] node1835;
	wire [8-1:0] node1836;
	wire [8-1:0] node1837;
	wire [8-1:0] node1839;
	wire [8-1:0] node1843;
	wire [8-1:0] node1844;
	wire [8-1:0] node1846;
	wire [8-1:0] node1849;
	wire [8-1:0] node1850;
	wire [8-1:0] node1854;
	wire [8-1:0] node1855;
	wire [8-1:0] node1857;
	wire [8-1:0] node1859;
	wire [8-1:0] node1862;
	wire [8-1:0] node1863;
	wire [8-1:0] node1864;
	wire [8-1:0] node1865;
	wire [8-1:0] node1866;
	wire [8-1:0] node1869;
	wire [8-1:0] node1870;
	wire [8-1:0] node1874;
	wire [8-1:0] node1875;
	wire [8-1:0] node1879;
	wire [8-1:0] node1880;
	wire [8-1:0] node1881;
	wire [8-1:0] node1882;
	wire [8-1:0] node1886;
	wire [8-1:0] node1889;
	wire [8-1:0] node1890;
	wire [8-1:0] node1894;
	wire [8-1:0] node1895;
	wire [8-1:0] node1896;
	wire [8-1:0] node1898;
	wire [8-1:0] node1901;
	wire [8-1:0] node1904;
	wire [8-1:0] node1905;
	wire [8-1:0] node1909;
	wire [8-1:0] node1910;
	wire [8-1:0] node1911;
	wire [8-1:0] node1912;
	wire [8-1:0] node1913;
	wire [8-1:0] node1914;
	wire [8-1:0] node1915;
	wire [8-1:0] node1916;
	wire [8-1:0] node1919;
	wire [8-1:0] node1922;
	wire [8-1:0] node1923;
	wire [8-1:0] node1925;
	wire [8-1:0] node1928;
	wire [8-1:0] node1931;
	wire [8-1:0] node1932;
	wire [8-1:0] node1934;
	wire [8-1:0] node1937;
	wire [8-1:0] node1938;
	wire [8-1:0] node1939;
	wire [8-1:0] node1942;
	wire [8-1:0] node1943;
	wire [8-1:0] node1947;
	wire [8-1:0] node1950;
	wire [8-1:0] node1951;
	wire [8-1:0] node1952;
	wire [8-1:0] node1953;
	wire [8-1:0] node1958;
	wire [8-1:0] node1959;
	wire [8-1:0] node1960;
	wire [8-1:0] node1963;
	wire [8-1:0] node1964;
	wire [8-1:0] node1965;
	wire [8-1:0] node1970;
	wire [8-1:0] node1971;
	wire [8-1:0] node1974;
	wire [8-1:0] node1977;
	wire [8-1:0] node1978;
	wire [8-1:0] node1979;
	wire [8-1:0] node1980;
	wire [8-1:0] node1983;
	wire [8-1:0] node1984;
	wire [8-1:0] node1988;
	wire [8-1:0] node1989;
	wire [8-1:0] node1992;
	wire [8-1:0] node1995;
	wire [8-1:0] node1996;
	wire [8-1:0] node1997;
	wire [8-1:0] node1998;
	wire [8-1:0] node2000;
	wire [8-1:0] node2002;
	wire [8-1:0] node2005;
	wire [8-1:0] node2008;
	wire [8-1:0] node2011;
	wire [8-1:0] node2012;
	wire [8-1:0] node2015;
	wire [8-1:0] node2016;
	wire [8-1:0] node2019;
	wire [8-1:0] node2022;
	wire [8-1:0] node2023;
	wire [8-1:0] node2024;
	wire [8-1:0] node2025;
	wire [8-1:0] node2027;
	wire [8-1:0] node2028;
	wire [8-1:0] node2031;
	wire [8-1:0] node2032;
	wire [8-1:0] node2036;
	wire [8-1:0] node2037;
	wire [8-1:0] node2039;
	wire [8-1:0] node2041;
	wire [8-1:0] node2044;
	wire [8-1:0] node2045;
	wire [8-1:0] node2046;
	wire [8-1:0] node2050;
	wire [8-1:0] node2051;
	wire [8-1:0] node2055;
	wire [8-1:0] node2056;
	wire [8-1:0] node2057;
	wire [8-1:0] node2059;
	wire [8-1:0] node2062;
	wire [8-1:0] node2064;
	wire [8-1:0] node2067;
	wire [8-1:0] node2068;
	wire [8-1:0] node2071;
	wire [8-1:0] node2073;
	wire [8-1:0] node2076;
	wire [8-1:0] node2077;
	wire [8-1:0] node2078;
	wire [8-1:0] node2080;
	wire [8-1:0] node2081;
	wire [8-1:0] node2084;
	wire [8-1:0] node2085;
	wire [8-1:0] node2088;
	wire [8-1:0] node2091;
	wire [8-1:0] node2092;
	wire [8-1:0] node2093;
	wire [8-1:0] node2096;
	wire [8-1:0] node2099;
	wire [8-1:0] node2100;
	wire [8-1:0] node2102;
	wire [8-1:0] node2105;
	wire [8-1:0] node2108;
	wire [8-1:0] node2109;
	wire [8-1:0] node2110;
	wire [8-1:0] node2111;
	wire [8-1:0] node2113;
	wire [8-1:0] node2117;
	wire [8-1:0] node2120;
	wire [8-1:0] node2121;
	wire [8-1:0] node2122;
	wire [8-1:0] node2126;
	wire [8-1:0] node2127;
	wire [8-1:0] node2130;
	wire [8-1:0] node2133;
	wire [8-1:0] node2134;
	wire [8-1:0] node2135;
	wire [8-1:0] node2136;
	wire [8-1:0] node2137;
	wire [8-1:0] node2138;
	wire [8-1:0] node2139;
	wire [8-1:0] node2140;
	wire [8-1:0] node2144;
	wire [8-1:0] node2147;
	wire [8-1:0] node2149;
	wire [8-1:0] node2152;
	wire [8-1:0] node2153;
	wire [8-1:0] node2154;
	wire [8-1:0] node2159;
	wire [8-1:0] node2160;
	wire [8-1:0] node2161;
	wire [8-1:0] node2162;
	wire [8-1:0] node2165;
	wire [8-1:0] node2166;
	wire [8-1:0] node2169;
	wire [8-1:0] node2171;
	wire [8-1:0] node2174;
	wire [8-1:0] node2177;
	wire [8-1:0] node2178;
	wire [8-1:0] node2179;
	wire [8-1:0] node2182;
	wire [8-1:0] node2185;
	wire [8-1:0] node2188;
	wire [8-1:0] node2189;
	wire [8-1:0] node2190;
	wire [8-1:0] node2191;
	wire [8-1:0] node2193;
	wire [8-1:0] node2197;
	wire [8-1:0] node2198;
	wire [8-1:0] node2201;
	wire [8-1:0] node2204;
	wire [8-1:0] node2205;
	wire [8-1:0] node2207;
	wire [8-1:0] node2208;
	wire [8-1:0] node2212;
	wire [8-1:0] node2214;
	wire [8-1:0] node2217;
	wire [8-1:0] node2218;
	wire [8-1:0] node2219;
	wire [8-1:0] node2220;
	wire [8-1:0] node2221;
	wire [8-1:0] node2222;
	wire [8-1:0] node2223;
	wire [8-1:0] node2226;
	wire [8-1:0] node2229;
	wire [8-1:0] node2232;
	wire [8-1:0] node2233;
	wire [8-1:0] node2234;
	wire [8-1:0] node2238;
	wire [8-1:0] node2241;
	wire [8-1:0] node2242;
	wire [8-1:0] node2243;
	wire [8-1:0] node2245;
	wire [8-1:0] node2248;
	wire [8-1:0] node2251;
	wire [8-1:0] node2253;
	wire [8-1:0] node2256;
	wire [8-1:0] node2257;
	wire [8-1:0] node2260;
	wire [8-1:0] node2262;
	wire [8-1:0] node2265;
	wire [8-1:0] node2266;
	wire [8-1:0] node2267;
	wire [8-1:0] node2268;
	wire [8-1:0] node2269;
	wire [8-1:0] node2273;
	wire [8-1:0] node2274;
	wire [8-1:0] node2275;
	wire [8-1:0] node2278;
	wire [8-1:0] node2279;
	wire [8-1:0] node2283;
	wire [8-1:0] node2284;
	wire [8-1:0] node2288;
	wire [8-1:0] node2289;
	wire [8-1:0] node2291;
	wire [8-1:0] node2293;
	wire [8-1:0] node2296;
	wire [8-1:0] node2297;
	wire [8-1:0] node2299;
	wire [8-1:0] node2302;
	wire [8-1:0] node2305;
	wire [8-1:0] node2308;
	wire [8-1:0] node2309;
	wire [8-1:0] node2310;
	wire [8-1:0] node2311;
	wire [8-1:0] node2312;
	wire [8-1:0] node2313;
	wire [8-1:0] node2314;
	wire [8-1:0] node2315;
	wire [8-1:0] node2316;
	wire [8-1:0] node2317;
	wire [8-1:0] node2319;
	wire [8-1:0] node2322;
	wire [8-1:0] node2324;
	wire [8-1:0] node2327;
	wire [8-1:0] node2329;
	wire [8-1:0] node2331;
	wire [8-1:0] node2334;
	wire [8-1:0] node2335;
	wire [8-1:0] node2336;
	wire [8-1:0] node2338;
	wire [8-1:0] node2340;
	wire [8-1:0] node2343;
	wire [8-1:0] node2344;
	wire [8-1:0] node2346;
	wire [8-1:0] node2349;
	wire [8-1:0] node2351;
	wire [8-1:0] node2354;
	wire [8-1:0] node2355;
	wire [8-1:0] node2358;
	wire [8-1:0] node2360;
	wire [8-1:0] node2363;
	wire [8-1:0] node2364;
	wire [8-1:0] node2365;
	wire [8-1:0] node2366;
	wire [8-1:0] node2369;
	wire [8-1:0] node2370;
	wire [8-1:0] node2371;
	wire [8-1:0] node2375;
	wire [8-1:0] node2378;
	wire [8-1:0] node2379;
	wire [8-1:0] node2380;
	wire [8-1:0] node2384;
	wire [8-1:0] node2386;
	wire [8-1:0] node2389;
	wire [8-1:0] node2390;
	wire [8-1:0] node2392;
	wire [8-1:0] node2393;
	wire [8-1:0] node2396;
	wire [8-1:0] node2399;
	wire [8-1:0] node2400;
	wire [8-1:0] node2402;
	wire [8-1:0] node2405;
	wire [8-1:0] node2408;
	wire [8-1:0] node2409;
	wire [8-1:0] node2410;
	wire [8-1:0] node2411;
	wire [8-1:0] node2412;
	wire [8-1:0] node2414;
	wire [8-1:0] node2417;
	wire [8-1:0] node2419;
	wire [8-1:0] node2422;
	wire [8-1:0] node2423;
	wire [8-1:0] node2425;
	wire [8-1:0] node2429;
	wire [8-1:0] node2430;
	wire [8-1:0] node2431;
	wire [8-1:0] node2433;
	wire [8-1:0] node2436;
	wire [8-1:0] node2437;
	wire [8-1:0] node2441;
	wire [8-1:0] node2442;
	wire [8-1:0] node2445;
	wire [8-1:0] node2446;
	wire [8-1:0] node2450;
	wire [8-1:0] node2451;
	wire [8-1:0] node2452;
	wire [8-1:0] node2454;
	wire [8-1:0] node2455;
	wire [8-1:0] node2456;
	wire [8-1:0] node2461;
	wire [8-1:0] node2462;
	wire [8-1:0] node2463;
	wire [8-1:0] node2466;
	wire [8-1:0] node2469;
	wire [8-1:0] node2470;
	wire [8-1:0] node2474;
	wire [8-1:0] node2475;
	wire [8-1:0] node2476;
	wire [8-1:0] node2479;
	wire [8-1:0] node2481;
	wire [8-1:0] node2484;
	wire [8-1:0] node2485;
	wire [8-1:0] node2487;
	wire [8-1:0] node2490;
	wire [8-1:0] node2491;
	wire [8-1:0] node2493;
	wire [8-1:0] node2494;
	wire [8-1:0] node2498;
	wire [8-1:0] node2501;
	wire [8-1:0] node2502;
	wire [8-1:0] node2503;
	wire [8-1:0] node2504;
	wire [8-1:0] node2505;
	wire [8-1:0] node2506;
	wire [8-1:0] node2509;
	wire [8-1:0] node2510;
	wire [8-1:0] node2514;
	wire [8-1:0] node2515;
	wire [8-1:0] node2517;
	wire [8-1:0] node2521;
	wire [8-1:0] node2522;
	wire [8-1:0] node2523;
	wire [8-1:0] node2524;
	wire [8-1:0] node2528;
	wire [8-1:0] node2529;
	wire [8-1:0] node2532;
	wire [8-1:0] node2535;
	wire [8-1:0] node2536;
	wire [8-1:0] node2538;
	wire [8-1:0] node2540;
	wire [8-1:0] node2543;
	wire [8-1:0] node2544;
	wire [8-1:0] node2548;
	wire [8-1:0] node2549;
	wire [8-1:0] node2550;
	wire [8-1:0] node2551;
	wire [8-1:0] node2552;
	wire [8-1:0] node2554;
	wire [8-1:0] node2556;
	wire [8-1:0] node2560;
	wire [8-1:0] node2561;
	wire [8-1:0] node2563;
	wire [8-1:0] node2566;
	wire [8-1:0] node2569;
	wire [8-1:0] node2570;
	wire [8-1:0] node2571;
	wire [8-1:0] node2574;
	wire [8-1:0] node2577;
	wire [8-1:0] node2580;
	wire [8-1:0] node2581;
	wire [8-1:0] node2582;
	wire [8-1:0] node2583;
	wire [8-1:0] node2586;
	wire [8-1:0] node2589;
	wire [8-1:0] node2592;
	wire [8-1:0] node2593;
	wire [8-1:0] node2594;
	wire [8-1:0] node2598;
	wire [8-1:0] node2601;
	wire [8-1:0] node2602;
	wire [8-1:0] node2603;
	wire [8-1:0] node2604;
	wire [8-1:0] node2605;
	wire [8-1:0] node2609;
	wire [8-1:0] node2612;
	wire [8-1:0] node2613;
	wire [8-1:0] node2614;
	wire [8-1:0] node2617;
	wire [8-1:0] node2618;
	wire [8-1:0] node2620;
	wire [8-1:0] node2624;
	wire [8-1:0] node2625;
	wire [8-1:0] node2627;
	wire [8-1:0] node2629;
	wire [8-1:0] node2632;
	wire [8-1:0] node2633;
	wire [8-1:0] node2635;
	wire [8-1:0] node2638;
	wire [8-1:0] node2641;
	wire [8-1:0] node2642;
	wire [8-1:0] node2643;
	wire [8-1:0] node2644;
	wire [8-1:0] node2645;
	wire [8-1:0] node2646;
	wire [8-1:0] node2650;
	wire [8-1:0] node2651;
	wire [8-1:0] node2655;
	wire [8-1:0] node2657;
	wire [8-1:0] node2660;
	wire [8-1:0] node2662;
	wire [8-1:0] node2663;
	wire [8-1:0] node2665;
	wire [8-1:0] node2669;
	wire [8-1:0] node2670;
	wire [8-1:0] node2671;
	wire [8-1:0] node2672;
	wire [8-1:0] node2673;
	wire [8-1:0] node2674;
	wire [8-1:0] node2680;
	wire [8-1:0] node2682;
	wire [8-1:0] node2685;
	wire [8-1:0] node2686;
	wire [8-1:0] node2687;
	wire [8-1:0] node2688;
	wire [8-1:0] node2692;
	wire [8-1:0] node2695;
	wire [8-1:0] node2697;
	wire [8-1:0] node2700;
	wire [8-1:0] node2701;
	wire [8-1:0] node2702;
	wire [8-1:0] node2703;
	wire [8-1:0] node2704;
	wire [8-1:0] node2705;
	wire [8-1:0] node2706;
	wire [8-1:0] node2709;
	wire [8-1:0] node2712;
	wire [8-1:0] node2713;
	wire [8-1:0] node2714;
	wire [8-1:0] node2718;
	wire [8-1:0] node2721;
	wire [8-1:0] node2722;
	wire [8-1:0] node2725;
	wire [8-1:0] node2727;
	wire [8-1:0] node2730;
	wire [8-1:0] node2731;
	wire [8-1:0] node2732;
	wire [8-1:0] node2733;
	wire [8-1:0] node2736;
	wire [8-1:0] node2737;
	wire [8-1:0] node2740;
	wire [8-1:0] node2741;
	wire [8-1:0] node2744;
	wire [8-1:0] node2747;
	wire [8-1:0] node2748;
	wire [8-1:0] node2749;
	wire [8-1:0] node2752;
	wire [8-1:0] node2755;
	wire [8-1:0] node2758;
	wire [8-1:0] node2759;
	wire [8-1:0] node2760;
	wire [8-1:0] node2761;
	wire [8-1:0] node2764;
	wire [8-1:0] node2765;
	wire [8-1:0] node2767;
	wire [8-1:0] node2771;
	wire [8-1:0] node2773;
	wire [8-1:0] node2775;
	wire [8-1:0] node2776;
	wire [8-1:0] node2779;
	wire [8-1:0] node2782;
	wire [8-1:0] node2783;
	wire [8-1:0] node2784;
	wire [8-1:0] node2787;
	wire [8-1:0] node2789;
	wire [8-1:0] node2790;
	wire [8-1:0] node2794;
	wire [8-1:0] node2797;
	wire [8-1:0] node2798;
	wire [8-1:0] node2799;
	wire [8-1:0] node2800;
	wire [8-1:0] node2803;
	wire [8-1:0] node2804;
	wire [8-1:0] node2806;
	wire [8-1:0] node2809;
	wire [8-1:0] node2812;
	wire [8-1:0] node2813;
	wire [8-1:0] node2814;
	wire [8-1:0] node2818;
	wire [8-1:0] node2820;
	wire [8-1:0] node2821;
	wire [8-1:0] node2825;
	wire [8-1:0] node2826;
	wire [8-1:0] node2827;
	wire [8-1:0] node2829;
	wire [8-1:0] node2832;
	wire [8-1:0] node2834;
	wire [8-1:0] node2837;
	wire [8-1:0] node2838;
	wire [8-1:0] node2842;
	wire [8-1:0] node2843;
	wire [8-1:0] node2844;
	wire [8-1:0] node2845;
	wire [8-1:0] node2846;
	wire [8-1:0] node2847;
	wire [8-1:0] node2848;
	wire [8-1:0] node2851;
	wire [8-1:0] node2854;
	wire [8-1:0] node2856;
	wire [8-1:0] node2859;
	wire [8-1:0] node2860;
	wire [8-1:0] node2862;
	wire [8-1:0] node2864;
	wire [8-1:0] node2867;
	wire [8-1:0] node2869;
	wire [8-1:0] node2870;
	wire [8-1:0] node2874;
	wire [8-1:0] node2875;
	wire [8-1:0] node2876;
	wire [8-1:0] node2878;
	wire [8-1:0] node2881;
	wire [8-1:0] node2882;
	wire [8-1:0] node2884;
	wire [8-1:0] node2887;
	wire [8-1:0] node2890;
	wire [8-1:0] node2891;
	wire [8-1:0] node2893;
	wire [8-1:0] node2896;
	wire [8-1:0] node2898;
	wire [8-1:0] node2901;
	wire [8-1:0] node2902;
	wire [8-1:0] node2903;
	wire [8-1:0] node2904;
	wire [8-1:0] node2906;
	wire [8-1:0] node2909;
	wire [8-1:0] node2912;
	wire [8-1:0] node2913;
	wire [8-1:0] node2914;
	wire [8-1:0] node2915;
	wire [8-1:0] node2919;
	wire [8-1:0] node2922;
	wire [8-1:0] node2923;
	wire [8-1:0] node2925;
	wire [8-1:0] node2929;
	wire [8-1:0] node2930;
	wire [8-1:0] node2931;
	wire [8-1:0] node2932;
	wire [8-1:0] node2936;
	wire [8-1:0] node2938;
	wire [8-1:0] node2941;
	wire [8-1:0] node2944;
	wire [8-1:0] node2945;
	wire [8-1:0] node2946;
	wire [8-1:0] node2947;
	wire [8-1:0] node2948;
	wire [8-1:0] node2950;
	wire [8-1:0] node2953;
	wire [8-1:0] node2954;
	wire [8-1:0] node2956;
	wire [8-1:0] node2959;
	wire [8-1:0] node2962;
	wire [8-1:0] node2963;
	wire [8-1:0] node2964;
	wire [8-1:0] node2968;
	wire [8-1:0] node2969;
	wire [8-1:0] node2971;
	wire [8-1:0] node2974;
	wire [8-1:0] node2977;
	wire [8-1:0] node2978;
	wire [8-1:0] node2979;
	wire [8-1:0] node2980;
	wire [8-1:0] node2984;
	wire [8-1:0] node2987;
	wire [8-1:0] node2988;
	wire [8-1:0] node2990;
	wire [8-1:0] node2993;
	wire [8-1:0] node2994;
	wire [8-1:0] node2997;
	wire [8-1:0] node2999;
	wire [8-1:0] node3002;
	wire [8-1:0] node3003;
	wire [8-1:0] node3004;
	wire [8-1:0] node3005;
	wire [8-1:0] node3008;
	wire [8-1:0] node3009;
	wire [8-1:0] node3010;
	wire [8-1:0] node3011;
	wire [8-1:0] node3015;
	wire [8-1:0] node3018;
	wire [8-1:0] node3021;
	wire [8-1:0] node3022;
	wire [8-1:0] node3024;
	wire [8-1:0] node3027;
	wire [8-1:0] node3028;
	wire [8-1:0] node3029;
	wire [8-1:0] node3032;
	wire [8-1:0] node3035;
	wire [8-1:0] node3038;
	wire [8-1:0] node3039;
	wire [8-1:0] node3041;
	wire [8-1:0] node3042;
	wire [8-1:0] node3046;
	wire [8-1:0] node3047;
	wire [8-1:0] node3048;
	wire [8-1:0] node3051;
	wire [8-1:0] node3054;
	wire [8-1:0] node3055;
	wire [8-1:0] node3058;
	wire [8-1:0] node3061;
	wire [8-1:0] node3062;
	wire [8-1:0] node3063;
	wire [8-1:0] node3064;
	wire [8-1:0] node3065;
	wire [8-1:0] node3066;
	wire [8-1:0] node3067;
	wire [8-1:0] node3069;
	wire [8-1:0] node3072;
	wire [8-1:0] node3073;
	wire [8-1:0] node3074;
	wire [8-1:0] node3078;
	wire [8-1:0] node3081;
	wire [8-1:0] node3082;
	wire [8-1:0] node3083;
	wire [8-1:0] node3084;
	wire [8-1:0] node3088;
	wire [8-1:0] node3089;
	wire [8-1:0] node3090;
	wire [8-1:0] node3094;
	wire [8-1:0] node3097;
	wire [8-1:0] node3098;
	wire [8-1:0] node3099;
	wire [8-1:0] node3103;
	wire [8-1:0] node3105;
	wire [8-1:0] node3108;
	wire [8-1:0] node3109;
	wire [8-1:0] node3111;
	wire [8-1:0] node3112;
	wire [8-1:0] node3114;
	wire [8-1:0] node3117;
	wire [8-1:0] node3118;
	wire [8-1:0] node3122;
	wire [8-1:0] node3123;
	wire [8-1:0] node3124;
	wire [8-1:0] node3125;
	wire [8-1:0] node3129;
	wire [8-1:0] node3131;
	wire [8-1:0] node3134;
	wire [8-1:0] node3135;
	wire [8-1:0] node3136;
	wire [8-1:0] node3140;
	wire [8-1:0] node3142;
	wire [8-1:0] node3145;
	wire [8-1:0] node3146;
	wire [8-1:0] node3147;
	wire [8-1:0] node3148;
	wire [8-1:0] node3152;
	wire [8-1:0] node3153;
	wire [8-1:0] node3154;
	wire [8-1:0] node3158;
	wire [8-1:0] node3160;
	wire [8-1:0] node3163;
	wire [8-1:0] node3164;
	wire [8-1:0] node3165;
	wire [8-1:0] node3168;
	wire [8-1:0] node3170;
	wire [8-1:0] node3173;
	wire [8-1:0] node3174;
	wire [8-1:0] node3175;
	wire [8-1:0] node3179;
	wire [8-1:0] node3182;
	wire [8-1:0] node3183;
	wire [8-1:0] node3184;
	wire [8-1:0] node3185;
	wire [8-1:0] node3186;
	wire [8-1:0] node3187;
	wire [8-1:0] node3188;
	wire [8-1:0] node3189;
	wire [8-1:0] node3192;
	wire [8-1:0] node3195;
	wire [8-1:0] node3197;
	wire [8-1:0] node3199;
	wire [8-1:0] node3202;
	wire [8-1:0] node3203;
	wire [8-1:0] node3207;
	wire [8-1:0] node3208;
	wire [8-1:0] node3209;
	wire [8-1:0] node3210;
	wire [8-1:0] node3214;
	wire [8-1:0] node3217;
	wire [8-1:0] node3218;
	wire [8-1:0] node3221;
	wire [8-1:0] node3223;
	wire [8-1:0] node3226;
	wire [8-1:0] node3227;
	wire [8-1:0] node3228;
	wire [8-1:0] node3232;
	wire [8-1:0] node3233;
	wire [8-1:0] node3234;
	wire [8-1:0] node3236;
	wire [8-1:0] node3239;
	wire [8-1:0] node3242;
	wire [8-1:0] node3243;
	wire [8-1:0] node3246;
	wire [8-1:0] node3249;
	wire [8-1:0] node3250;
	wire [8-1:0] node3251;
	wire [8-1:0] node3252;
	wire [8-1:0] node3253;
	wire [8-1:0] node3256;
	wire [8-1:0] node3259;
	wire [8-1:0] node3260;
	wire [8-1:0] node3264;
	wire [8-1:0] node3265;
	wire [8-1:0] node3268;
	wire [8-1:0] node3269;
	wire [8-1:0] node3273;
	wire [8-1:0] node3274;
	wire [8-1:0] node3275;
	wire [8-1:0] node3276;
	wire [8-1:0] node3280;
	wire [8-1:0] node3282;
	wire [8-1:0] node3283;
	wire [8-1:0] node3286;
	wire [8-1:0] node3289;
	wire [8-1:0] node3290;
	wire [8-1:0] node3293;
	wire [8-1:0] node3294;
	wire [8-1:0] node3298;
	wire [8-1:0] node3299;
	wire [8-1:0] node3300;
	wire [8-1:0] node3301;
	wire [8-1:0] node3302;
	wire [8-1:0] node3305;
	wire [8-1:0] node3307;
	wire [8-1:0] node3310;
	wire [8-1:0] node3311;
	wire [8-1:0] node3314;
	wire [8-1:0] node3316;
	wire [8-1:0] node3319;
	wire [8-1:0] node3320;
	wire [8-1:0] node3321;
	wire [8-1:0] node3324;
	wire [8-1:0] node3327;
	wire [8-1:0] node3328;
	wire [8-1:0] node3329;
	wire [8-1:0] node3332;
	wire [8-1:0] node3335;
	wire [8-1:0] node3336;
	wire [8-1:0] node3339;
	wire [8-1:0] node3342;
	wire [8-1:0] node3343;
	wire [8-1:0] node3344;
	wire [8-1:0] node3345;
	wire [8-1:0] node3348;
	wire [8-1:0] node3350;
	wire [8-1:0] node3353;
	wire [8-1:0] node3354;
	wire [8-1:0] node3357;
	wire [8-1:0] node3358;
	wire [8-1:0] node3361;
	wire [8-1:0] node3363;
	wire [8-1:0] node3366;
	wire [8-1:0] node3367;
	wire [8-1:0] node3368;
	wire [8-1:0] node3370;
	wire [8-1:0] node3373;
	wire [8-1:0] node3375;
	wire [8-1:0] node3378;
	wire [8-1:0] node3380;
	wire [8-1:0] node3381;
	wire [8-1:0] node3384;
	wire [8-1:0] node3387;
	wire [8-1:0] node3388;
	wire [8-1:0] node3389;
	wire [8-1:0] node3390;
	wire [8-1:0] node3391;
	wire [8-1:0] node3392;
	wire [8-1:0] node3393;
	wire [8-1:0] node3394;
	wire [8-1:0] node3397;
	wire [8-1:0] node3400;
	wire [8-1:0] node3401;
	wire [8-1:0] node3404;
	wire [8-1:0] node3407;
	wire [8-1:0] node3408;
	wire [8-1:0] node3410;
	wire [8-1:0] node3413;
	wire [8-1:0] node3414;
	wire [8-1:0] node3415;
	wire [8-1:0] node3417;
	wire [8-1:0] node3421;
	wire [8-1:0] node3424;
	wire [8-1:0] node3425;
	wire [8-1:0] node3426;
	wire [8-1:0] node3428;
	wire [8-1:0] node3431;
	wire [8-1:0] node3432;
	wire [8-1:0] node3435;
	wire [8-1:0] node3437;
	wire [8-1:0] node3440;
	wire [8-1:0] node3441;
	wire [8-1:0] node3442;
	wire [8-1:0] node3445;
	wire [8-1:0] node3448;
	wire [8-1:0] node3449;
	wire [8-1:0] node3452;
	wire [8-1:0] node3455;
	wire [8-1:0] node3456;
	wire [8-1:0] node3457;
	wire [8-1:0] node3458;
	wire [8-1:0] node3459;
	wire [8-1:0] node3461;
	wire [8-1:0] node3465;
	wire [8-1:0] node3468;
	wire [8-1:0] node3469;
	wire [8-1:0] node3470;
	wire [8-1:0] node3471;
	wire [8-1:0] node3475;
	wire [8-1:0] node3476;
	wire [8-1:0] node3480;
	wire [8-1:0] node3481;
	wire [8-1:0] node3482;
	wire [8-1:0] node3483;
	wire [8-1:0] node3488;
	wire [8-1:0] node3490;
	wire [8-1:0] node3493;
	wire [8-1:0] node3494;
	wire [8-1:0] node3495;
	wire [8-1:0] node3496;
	wire [8-1:0] node3499;
	wire [8-1:0] node3502;
	wire [8-1:0] node3503;
	wire [8-1:0] node3506;
	wire [8-1:0] node3509;
	wire [8-1:0] node3510;
	wire [8-1:0] node3511;
	wire [8-1:0] node3514;
	wire [8-1:0] node3517;
	wire [8-1:0] node3518;
	wire [8-1:0] node3519;
	wire [8-1:0] node3523;
	wire [8-1:0] node3525;
	wire [8-1:0] node3528;
	wire [8-1:0] node3529;
	wire [8-1:0] node3530;
	wire [8-1:0] node3531;
	wire [8-1:0] node3532;
	wire [8-1:0] node3533;
	wire [8-1:0] node3534;
	wire [8-1:0] node3537;
	wire [8-1:0] node3540;
	wire [8-1:0] node3541;
	wire [8-1:0] node3545;
	wire [8-1:0] node3547;
	wire [8-1:0] node3549;
	wire [8-1:0] node3552;
	wire [8-1:0] node3553;
	wire [8-1:0] node3554;
	wire [8-1:0] node3555;
	wire [8-1:0] node3560;
	wire [8-1:0] node3561;
	wire [8-1:0] node3562;
	wire [8-1:0] node3566;
	wire [8-1:0] node3569;
	wire [8-1:0] node3570;
	wire [8-1:0] node3571;
	wire [8-1:0] node3572;
	wire [8-1:0] node3575;
	wire [8-1:0] node3578;
	wire [8-1:0] node3580;
	wire [8-1:0] node3583;
	wire [8-1:0] node3584;
	wire [8-1:0] node3585;
	wire [8-1:0] node3588;
	wire [8-1:0] node3590;
	wire [8-1:0] node3592;
	wire [8-1:0] node3595;
	wire [8-1:0] node3596;
	wire [8-1:0] node3597;
	wire [8-1:0] node3602;
	wire [8-1:0] node3603;
	wire [8-1:0] node3604;
	wire [8-1:0] node3605;
	wire [8-1:0] node3607;
	wire [8-1:0] node3608;
	wire [8-1:0] node3612;
	wire [8-1:0] node3613;
	wire [8-1:0] node3615;
	wire [8-1:0] node3618;
	wire [8-1:0] node3621;
	wire [8-1:0] node3622;
	wire [8-1:0] node3624;
	wire [8-1:0] node3625;
	wire [8-1:0] node3629;
	wire [8-1:0] node3631;
	wire [8-1:0] node3634;
	wire [8-1:0] node3635;
	wire [8-1:0] node3636;
	wire [8-1:0] node3637;
	wire [8-1:0] node3640;
	wire [8-1:0] node3642;
	wire [8-1:0] node3645;
	wire [8-1:0] node3648;
	wire [8-1:0] node3649;
	wire [8-1:0] node3650;
	wire [8-1:0] node3653;
	wire [8-1:0] node3654;
	wire [8-1:0] node3655;
	wire [8-1:0] node3660;
	wire [8-1:0] node3661;
	wire [8-1:0] node3665;
	wire [8-1:0] node3666;
	wire [8-1:0] node3667;
	wire [8-1:0] node3668;
	wire [8-1:0] node3669;
	wire [8-1:0] node3670;
	wire [8-1:0] node3671;
	wire [8-1:0] node3675;
	wire [8-1:0] node3678;
	wire [8-1:0] node3679;
	wire [8-1:0] node3683;
	wire [8-1:0] node3684;
	wire [8-1:0] node3685;
	wire [8-1:0] node3686;
	wire [8-1:0] node3690;
	wire [8-1:0] node3692;
	wire [8-1:0] node3695;
	wire [8-1:0] node3696;
	wire [8-1:0] node3697;
	wire [8-1:0] node3702;
	wire [8-1:0] node3703;
	wire [8-1:0] node3704;
	wire [8-1:0] node3705;
	wire [8-1:0] node3707;
	wire [8-1:0] node3710;
	wire [8-1:0] node3712;
	wire [8-1:0] node3715;
	wire [8-1:0] node3716;
	wire [8-1:0] node3717;
	wire [8-1:0] node3720;
	wire [8-1:0] node3723;
	wire [8-1:0] node3725;
	wire [8-1:0] node3728;
	wire [8-1:0] node3729;
	wire [8-1:0] node3730;
	wire [8-1:0] node3732;
	wire [8-1:0] node3736;
	wire [8-1:0] node3738;
	wire [8-1:0] node3741;
	wire [8-1:0] node3742;
	wire [8-1:0] node3743;
	wire [8-1:0] node3744;
	wire [8-1:0] node3745;
	wire [8-1:0] node3746;
	wire [8-1:0] node3748;
	wire [8-1:0] node3751;
	wire [8-1:0] node3754;
	wire [8-1:0] node3757;
	wire [8-1:0] node3758;
	wire [8-1:0] node3761;
	wire [8-1:0] node3764;
	wire [8-1:0] node3765;
	wire [8-1:0] node3766;
	wire [8-1:0] node3767;
	wire [8-1:0] node3770;
	wire [8-1:0] node3773;
	wire [8-1:0] node3774;
	wire [8-1:0] node3776;
	wire [8-1:0] node3780;
	wire [8-1:0] node3781;
	wire [8-1:0] node3782;
	wire [8-1:0] node3784;
	wire [8-1:0] node3789;
	wire [8-1:0] node3790;
	wire [8-1:0] node3791;
	wire [8-1:0] node3792;
	wire [8-1:0] node3793;
	wire [8-1:0] node3796;
	wire [8-1:0] node3799;
	wire [8-1:0] node3802;
	wire [8-1:0] node3803;
	wire [8-1:0] node3804;
	wire [8-1:0] node3808;
	wire [8-1:0] node3811;
	wire [8-1:0] node3812;
	wire [8-1:0] node3813;
	wire [8-1:0] node3816;
	wire [8-1:0] node3819;
	wire [8-1:0] node3822;
	wire [8-1:0] node3823;
	wire [8-1:0] node3824;
	wire [8-1:0] node3825;
	wire [8-1:0] node3827;
	wire [8-1:0] node3828;
	wire [8-1:0] node3829;
	wire [8-1:0] node3830;
	wire [8-1:0] node3832;
	wire [8-1:0] node3835;
	wire [8-1:0] node3838;
	wire [8-1:0] node3839;
	wire [8-1:0] node3840;
	wire [8-1:0] node3842;
	wire [8-1:0] node3846;
	wire [8-1:0] node3847;
	wire [8-1:0] node3849;
	wire [8-1:0] node3852;
	wire [8-1:0] node3855;
	wire [8-1:0] node3856;
	wire [8-1:0] node3857;
	wire [8-1:0] node3858;
	wire [8-1:0] node3861;
	wire [8-1:0] node3863;
	wire [8-1:0] node3866;
	wire [8-1:0] node3867;
	wire [8-1:0] node3870;
	wire [8-1:0] node3871;
	wire [8-1:0] node3873;
	wire [8-1:0] node3876;
	wire [8-1:0] node3879;
	wire [8-1:0] node3880;
	wire [8-1:0] node3881;
	wire [8-1:0] node3884;
	wire [8-1:0] node3887;
	wire [8-1:0] node3888;
	wire [8-1:0] node3890;
	wire [8-1:0] node3893;
	wire [8-1:0] node3894;
	wire [8-1:0] node3896;
	wire [8-1:0] node3899;
	wire [8-1:0] node3902;
	wire [8-1:0] node3903;
	wire [8-1:0] node3904;
	wire [8-1:0] node3905;
	wire [8-1:0] node3907;
	wire [8-1:0] node3908;
	wire [8-1:0] node3912;
	wire [8-1:0] node3913;
	wire [8-1:0] node3915;
	wire [8-1:0] node3918;
	wire [8-1:0] node3919;
	wire [8-1:0] node3923;
	wire [8-1:0] node3924;
	wire [8-1:0] node3925;
	wire [8-1:0] node3926;
	wire [8-1:0] node3927;
	wire [8-1:0] node3931;
	wire [8-1:0] node3932;
	wire [8-1:0] node3935;
	wire [8-1:0] node3938;
	wire [8-1:0] node3939;
	wire [8-1:0] node3942;
	wire [8-1:0] node3943;
	wire [8-1:0] node3947;
	wire [8-1:0] node3948;
	wire [8-1:0] node3951;
	wire [8-1:0] node3954;
	wire [8-1:0] node3955;
	wire [8-1:0] node3956;
	wire [8-1:0] node3957;
	wire [8-1:0] node3958;
	wire [8-1:0] node3962;
	wire [8-1:0] node3963;
	wire [8-1:0] node3964;
	wire [8-1:0] node3967;
	wire [8-1:0] node3971;
	wire [8-1:0] node3972;
	wire [8-1:0] node3973;
	wire [8-1:0] node3977;
	wire [8-1:0] node3978;
	wire [8-1:0] node3979;
	wire [8-1:0] node3980;
	wire [8-1:0] node3984;
	wire [8-1:0] node3988;
	wire [8-1:0] node3989;
	wire [8-1:0] node3990;
	wire [8-1:0] node3991;
	wire [8-1:0] node3992;
	wire [8-1:0] node3996;
	wire [8-1:0] node3999;
	wire [8-1:0] node4000;
	wire [8-1:0] node4001;
	wire [8-1:0] node4002;
	wire [8-1:0] node4005;
	wire [8-1:0] node4008;
	wire [8-1:0] node4012;
	wire [8-1:0] node4013;
	wire [8-1:0] node4014;
	wire [8-1:0] node4015;
	wire [8-1:0] node4017;
	wire [8-1:0] node4020;
	wire [8-1:0] node4021;
	wire [8-1:0] node4025;
	wire [8-1:0] node4026;
	wire [8-1:0] node4028;
	wire [8-1:0] node4031;
	wire [8-1:0] node4032;
	wire [8-1:0] node4035;
	wire [8-1:0] node4038;
	wire [8-1:0] node4041;
	wire [8-1:0] node4042;
	wire [8-1:0] node4044;
	wire [8-1:0] node4045;
	wire [8-1:0] node4046;
	wire [8-1:0] node4047;
	wire [8-1:0] node4049;
	wire [8-1:0] node4052;
	wire [8-1:0] node4053;
	wire [8-1:0] node4055;
	wire [8-1:0] node4059;
	wire [8-1:0] node4060;
	wire [8-1:0] node4063;
	wire [8-1:0] node4064;
	wire [8-1:0] node4066;
	wire [8-1:0] node4069;
	wire [8-1:0] node4072;
	wire [8-1:0] node4073;
	wire [8-1:0] node4074;
	wire [8-1:0] node4075;
	wire [8-1:0] node4078;
	wire [8-1:0] node4079;
	wire [8-1:0] node4083;
	wire [8-1:0] node4084;
	wire [8-1:0] node4087;
	wire [8-1:0] node4089;
	wire [8-1:0] node4090;
	wire [8-1:0] node4094;
	wire [8-1:0] node4095;
	wire [8-1:0] node4097;
	wire [8-1:0] node4100;
	wire [8-1:0] node4101;
	wire [8-1:0] node4103;
	wire [8-1:0] node4106;
	wire [8-1:0] node4108;
	wire [8-1:0] node4111;
	wire [8-1:0] node4112;
	wire [8-1:0] node4113;
	wire [8-1:0] node4114;
	wire [8-1:0] node4116;
	wire [8-1:0] node4118;
	wire [8-1:0] node4121;
	wire [8-1:0] node4122;
	wire [8-1:0] node4125;
	wire [8-1:0] node4126;
	wire [8-1:0] node4129;
	wire [8-1:0] node4131;
	wire [8-1:0] node4134;
	wire [8-1:0] node4135;
	wire [8-1:0] node4136;
	wire [8-1:0] node4137;
	wire [8-1:0] node4138;
	wire [8-1:0] node4142;
	wire [8-1:0] node4144;
	wire [8-1:0] node4147;
	wire [8-1:0] node4150;
	wire [8-1:0] node4151;
	wire [8-1:0] node4152;
	wire [8-1:0] node4153;
	wire [8-1:0] node4158;
	wire [8-1:0] node4159;
	wire [8-1:0] node4160;
	wire [8-1:0] node4164;
	wire [8-1:0] node4167;
	wire [8-1:0] node4168;
	wire [8-1:0] node4169;
	wire [8-1:0] node4170;
	wire [8-1:0] node4172;
	wire [8-1:0] node4174;
	wire [8-1:0] node4177;
	wire [8-1:0] node4178;
	wire [8-1:0] node4181;
	wire [8-1:0] node4184;
	wire [8-1:0] node4185;
	wire [8-1:0] node4186;
	wire [8-1:0] node4188;
	wire [8-1:0] node4191;
	wire [8-1:0] node4194;
	wire [8-1:0] node4195;
	wire [8-1:0] node4196;
	wire [8-1:0] node4199;
	wire [8-1:0] node4203;
	wire [8-1:0] node4204;
	wire [8-1:0] node4205;
	wire [8-1:0] node4206;
	wire [8-1:0] node4207;
	wire [8-1:0] node4208;
	wire [8-1:0] node4212;
	wire [8-1:0] node4214;
	wire [8-1:0] node4217;
	wire [8-1:0] node4219;
	wire [8-1:0] node4222;
	wire [8-1:0] node4225;
	wire [8-1:0] node4226;
	wire [8-1:0] node4227;
	wire [8-1:0] node4228;
	wire [8-1:0] node4230;
	wire [8-1:0] node4233;
	wire [8-1:0] node4236;
	wire [8-1:0] node4239;
	wire [8-1:0] node4242;
	wire [8-1:0] node4243;
	wire [8-1:0] node4245;
	wire [8-1:0] node4246;
	wire [8-1:0] node4247;
	wire [8-1:0] node4248;
	wire [8-1:0] node4249;
	wire [8-1:0] node4251;
	wire [8-1:0] node4252;
	wire [8-1:0] node4256;
	wire [8-1:0] node4257;
	wire [8-1:0] node4258;
	wire [8-1:0] node4260;
	wire [8-1:0] node4265;
	wire [8-1:0] node4266;
	wire [8-1:0] node4267;
	wire [8-1:0] node4270;
	wire [8-1:0] node4273;
	wire [8-1:0] node4275;
	wire [8-1:0] node4277;
	wire [8-1:0] node4280;
	wire [8-1:0] node4281;
	wire [8-1:0] node4282;
	wire [8-1:0] node4286;
	wire [8-1:0] node4287;
	wire [8-1:0] node4288;
	wire [8-1:0] node4292;
	wire [8-1:0] node4293;
	wire [8-1:0] node4295;
	wire [8-1:0] node4299;
	wire [8-1:0] node4300;
	wire [8-1:0] node4301;
	wire [8-1:0] node4302;
	wire [8-1:0] node4303;
	wire [8-1:0] node4304;
	wire [8-1:0] node4307;
	wire [8-1:0] node4309;
	wire [8-1:0] node4312;
	wire [8-1:0] node4313;
	wire [8-1:0] node4317;
	wire [8-1:0] node4318;
	wire [8-1:0] node4319;
	wire [8-1:0] node4322;
	wire [8-1:0] node4323;
	wire [8-1:0] node4327;
	wire [8-1:0] node4330;
	wire [8-1:0] node4331;
	wire [8-1:0] node4332;
	wire [8-1:0] node4334;
	wire [8-1:0] node4335;
	wire [8-1:0] node4339;
	wire [8-1:0] node4341;
	wire [8-1:0] node4344;
	wire [8-1:0] node4345;
	wire [8-1:0] node4346;
	wire [8-1:0] node4350;
	wire [8-1:0] node4352;
	wire [8-1:0] node4355;
	wire [8-1:0] node4356;
	wire [8-1:0] node4357;
	wire [8-1:0] node4358;
	wire [8-1:0] node4361;
	wire [8-1:0] node4363;
	wire [8-1:0] node4364;
	wire [8-1:0] node4367;
	wire [8-1:0] node4370;
	wire [8-1:0] node4371;
	wire [8-1:0] node4375;
	wire [8-1:0] node4376;
	wire [8-1:0] node4377;
	wire [8-1:0] node4379;
	wire [8-1:0] node4382;
	wire [8-1:0] node4383;
	wire [8-1:0] node4385;
	wire [8-1:0] node4388;
	wire [8-1:0] node4391;
	wire [8-1:0] node4393;
	wire [8-1:0] node4396;
	wire [8-1:0] node4397;
	wire [8-1:0] node4398;
	wire [8-1:0] node4399;
	wire [8-1:0] node4401;
	wire [8-1:0] node4402;
	wire [8-1:0] node4406;
	wire [8-1:0] node4407;
	wire [8-1:0] node4408;
	wire [8-1:0] node4410;
	wire [8-1:0] node4413;
	wire [8-1:0] node4415;
	wire [8-1:0] node4416;
	wire [8-1:0] node4417;
	wire [8-1:0] node4421;
	wire [8-1:0] node4424;
	wire [8-1:0] node4425;
	wire [8-1:0] node4427;
	wire [8-1:0] node4428;
	wire [8-1:0] node4432;
	wire [8-1:0] node4434;
	wire [8-1:0] node4435;
	wire [8-1:0] node4439;
	wire [8-1:0] node4440;
	wire [8-1:0] node4441;
	wire [8-1:0] node4443;
	wire [8-1:0] node4446;
	wire [8-1:0] node4447;
	wire [8-1:0] node4448;
	wire [8-1:0] node4451;
	wire [8-1:0] node4453;
	wire [8-1:0] node4456;
	wire [8-1:0] node4458;
	wire [8-1:0] node4460;
	wire [8-1:0] node4463;
	wire [8-1:0] node4464;
	wire [8-1:0] node4465;
	wire [8-1:0] node4468;
	wire [8-1:0] node4471;
	wire [8-1:0] node4472;
	wire [8-1:0] node4475;
	wire [8-1:0] node4478;
	wire [8-1:0] node4479;
	wire [8-1:0] node4480;
	wire [8-1:0] node4481;
	wire [8-1:0] node4482;
	wire [8-1:0] node4484;
	wire [8-1:0] node4486;
	wire [8-1:0] node4489;
	wire [8-1:0] node4490;
	wire [8-1:0] node4493;
	wire [8-1:0] node4494;
	wire [8-1:0] node4498;
	wire [8-1:0] node4499;
	wire [8-1:0] node4500;
	wire [8-1:0] node4502;
	wire [8-1:0] node4505;
	wire [8-1:0] node4506;
	wire [8-1:0] node4509;
	wire [8-1:0] node4512;
	wire [8-1:0] node4513;
	wire [8-1:0] node4514;
	wire [8-1:0] node4516;
	wire [8-1:0] node4520;
	wire [8-1:0] node4522;
	wire [8-1:0] node4523;
	wire [8-1:0] node4527;
	wire [8-1:0] node4528;
	wire [8-1:0] node4529;
	wire [8-1:0] node4531;
	wire [8-1:0] node4532;
	wire [8-1:0] node4536;
	wire [8-1:0] node4537;
	wire [8-1:0] node4539;
	wire [8-1:0] node4542;
	wire [8-1:0] node4544;
	wire [8-1:0] node4545;
	wire [8-1:0] node4549;
	wire [8-1:0] node4550;
	wire [8-1:0] node4552;
	wire [8-1:0] node4553;
	wire [8-1:0] node4557;
	wire [8-1:0] node4558;
	wire [8-1:0] node4561;
	wire [8-1:0] node4563;
	wire [8-1:0] node4565;
	wire [8-1:0] node4568;
	wire [8-1:0] node4569;
	wire [8-1:0] node4570;
	wire [8-1:0] node4571;
	wire [8-1:0] node4574;
	wire [8-1:0] node4577;
	wire [8-1:0] node4578;
	wire [8-1:0] node4582;
	wire [8-1:0] node4583;
	wire [8-1:0] node4584;
	wire [8-1:0] node4587;
	wire [8-1:0] node4590;
	wire [8-1:0] node4591;
	wire [8-1:0] node4594;

	assign outp = (inp[4]) ? node2308 : node1;
		assign node1 = (inp[13]) ? node1105 : node2;
			assign node2 = (inp[7]) ? node332 : node3;
				assign node3 = (inp[11]) ? node123 : node4;
					assign node4 = (inp[5]) ? node74 : node5;
						assign node5 = (inp[1]) ? node31 : node6;
							assign node6 = (inp[8]) ? node14 : node7;
								assign node7 = (inp[2]) ? node9 : 8'b01111111;
									assign node9 = (inp[6]) ? 8'b00101111 : node10;
										assign node10 = (inp[0]) ? 8'b01111111 : 8'b00101111;
								assign node14 = (inp[2]) ? node20 : node15;
									assign node15 = (inp[10]) ? 8'b00111011 : node16;
										assign node16 = (inp[0]) ? 8'b01111111 : 8'b00111011;
									assign node20 = (inp[6]) ? node26 : node21;
										assign node21 = (inp[0]) ? node23 : 8'b00101011;
											assign node23 = (inp[10]) ? 8'b00111011 : 8'b01111111;
										assign node26 = (inp[12]) ? node28 : 8'b00101011;
											assign node28 = (inp[10]) ? 8'b00101011 : 8'b00101111;
							assign node31 = (inp[2]) ? node47 : node32;
								assign node32 = (inp[8]) ? node38 : node33;
									assign node33 = (inp[3]) ? 8'b00111110 : node34;
										assign node34 = (inp[0]) ? 8'b01111111 : 8'b00111110;
									assign node38 = (inp[0]) ? node40 : 8'b00111010;
										assign node40 = (inp[10]) ? node44 : node41;
											assign node41 = (inp[3]) ? 8'b00111110 : 8'b01111111;
											assign node44 = (inp[3]) ? 8'b00111010 : 8'b00111011;
								assign node47 = (inp[8]) ? node57 : node48;
									assign node48 = (inp[0]) ? node50 : 8'b00101110;
										assign node50 = (inp[3]) ? node54 : node51;
											assign node51 = (inp[6]) ? 8'b00101111 : 8'b01111111;
											assign node54 = (inp[6]) ? 8'b00101110 : 8'b00111110;
									assign node57 = (inp[0]) ? node59 : 8'b00101010;
										assign node59 = (inp[6]) ? node67 : node60;
											assign node60 = (inp[3]) ? node64 : node61;
												assign node61 = (inp[10]) ? 8'b00111011 : 8'b01111111;
												assign node64 = (inp[10]) ? 8'b00111010 : 8'b00111110;
											assign node67 = (inp[10]) ? node71 : node68;
												assign node68 = (inp[3]) ? 8'b00101110 : 8'b00101111;
												assign node71 = (inp[3]) ? 8'b00101010 : 8'b00101011;
						assign node74 = (inp[0]) ? 8'b01111111 : node75;
							assign node75 = (inp[2]) ? node93 : node76;
								assign node76 = (inp[8]) ? node82 : node77;
									assign node77 = (inp[1]) ? node79 : 8'b01111111;
										assign node79 = (inp[3]) ? 8'b01111111 : 8'b00111110;
									assign node82 = (inp[10]) ? node88 : node83;
										assign node83 = (inp[3]) ? 8'b00111011 : node84;
											assign node84 = (inp[1]) ? 8'b00111010 : 8'b00111011;
										assign node88 = (inp[1]) ? node90 : 8'b01111111;
											assign node90 = (inp[3]) ? 8'b01111111 : 8'b00111110;
								assign node93 = (inp[6]) ? node111 : node94;
									assign node94 = (inp[8]) ? node102 : node95;
										assign node95 = (inp[9]) ? 8'b00101111 : node96;
											assign node96 = (inp[3]) ? 8'b00101111 : node97;
												assign node97 = (inp[1]) ? 8'b00101110 : 8'b00101111;
										assign node102 = (inp[10]) ? node108 : node103;
											assign node103 = (inp[3]) ? 8'b00101011 : node104;
												assign node104 = (inp[1]) ? 8'b00101010 : 8'b00101011;
											assign node108 = (inp[3]) ? 8'b00101111 : 8'b00101110;
									assign node111 = (inp[3]) ? 8'b01111111 : node112;
										assign node112 = (inp[1]) ? node116 : node113;
											assign node113 = (inp[10]) ? 8'b01111111 : 8'b00111011;
											assign node116 = (inp[10]) ? 8'b00111110 : node117;
												assign node117 = (inp[12]) ? 8'b00111110 : 8'b00111010;
					assign node123 = (inp[8]) ? node201 : node124;
						assign node124 = (inp[1]) ? node146 : node125;
							assign node125 = (inp[2]) ? node129 : node126;
								assign node126 = (inp[12]) ? 8'b01111111 : 8'b00101111;
								assign node129 = (inp[12]) ? node139 : node130;
									assign node130 = (inp[5]) ? node136 : node131;
										assign node131 = (inp[6]) ? 8'b00111110 : node132;
											assign node132 = (inp[3]) ? 8'b00101110 : 8'b00111110;
										assign node136 = (inp[6]) ? 8'b00101110 : 8'b00111110;
									assign node139 = (inp[5]) ? node141 : 8'b00101111;
										assign node141 = (inp[0]) ? 8'b00111110 : node142;
											assign node142 = (inp[6]) ? 8'b00111110 : 8'b00101111;
							assign node146 = (inp[12]) ? node174 : node147;
								assign node147 = (inp[2]) ? node159 : node148;
									assign node148 = (inp[0]) ? node154 : node149;
										assign node149 = (inp[5]) ? node151 : 8'b00101110;
											assign node151 = (inp[3]) ? 8'b00101011 : 8'b00101110;
										assign node154 = (inp[3]) ? node156 : 8'b00101011;
											assign node156 = (inp[5]) ? 8'b00101011 : 8'b00101110;
									assign node159 = (inp[5]) ? node167 : node160;
										assign node160 = (inp[0]) ? node162 : 8'b00111011;
											assign node162 = (inp[6]) ? 8'b00111011 : node163;
												assign node163 = (inp[3]) ? 8'b00101011 : 8'b00101010;
										assign node167 = (inp[3]) ? 8'b00101010 : node168;
											assign node168 = (inp[0]) ? 8'b00101010 : node169;
												assign node169 = (inp[6]) ? 8'b00101011 : 8'b00111011;
								assign node174 = (inp[2]) ? node186 : node175;
									assign node175 = (inp[0]) ? node181 : node176;
										assign node176 = (inp[3]) ? node178 : 8'b00111110;
											assign node178 = (inp[5]) ? 8'b00111011 : 8'b00111110;
										assign node181 = (inp[3]) ? node183 : 8'b00111011;
											assign node183 = (inp[5]) ? 8'b00111011 : 8'b00111110;
									assign node186 = (inp[0]) ? node192 : node187;
										assign node187 = (inp[5]) ? node189 : 8'b00101110;
											assign node189 = (inp[6]) ? 8'b00111011 : 8'b00101011;
										assign node192 = (inp[5]) ? 8'b00111010 : node193;
											assign node193 = (inp[6]) ? node197 : node194;
												assign node194 = (inp[3]) ? 8'b00111011 : 8'b00111010;
												assign node197 = (inp[3]) ? 8'b00101110 : 8'b00101011;
						assign node201 = (inp[5]) ? node263 : node202;
							assign node202 = (inp[0]) ? node218 : node203;
								assign node203 = (inp[1]) ? node211 : node204;
									assign node204 = (inp[12]) ? node208 : node205;
										assign node205 = (inp[2]) ? 8'b00111010 : 8'b00101011;
										assign node208 = (inp[2]) ? 8'b00101011 : 8'b00111011;
									assign node211 = (inp[12]) ? node215 : node212;
										assign node212 = (inp[2]) ? 8'b00011111 : 8'b00101010;
										assign node215 = (inp[2]) ? 8'b00101010 : 8'b00111010;
								assign node218 = (inp[10]) ? node240 : node219;
									assign node219 = (inp[2]) ? node227 : node220;
										assign node220 = (inp[1]) ? node224 : node221;
											assign node221 = (inp[12]) ? 8'b00011111 : 8'b00001111;
											assign node224 = (inp[12]) ? 8'b00011110 : 8'b00001110;
										assign node227 = (inp[1]) ? node233 : node228;
											assign node228 = (inp[3]) ? 8'b00001111 : node229;
												assign node229 = (inp[6]) ? 8'b00011110 : 8'b00001110;
											assign node233 = (inp[6]) ? node237 : node234;
												assign node234 = (inp[3]) ? 8'b00001011 : 8'b00001010;
												assign node237 = (inp[3]) ? 8'b00001110 : 8'b00001011;
									assign node240 = (inp[1]) ? node248 : node241;
										assign node241 = (inp[2]) ? node243 : 8'b00101011;
											assign node243 = (inp[6]) ? 8'b00111010 : node244;
												assign node244 = (inp[12]) ? 8'b00111010 : 8'b00101010;
										assign node248 = (inp[3]) ? node254 : node249;
											assign node249 = (inp[12]) ? node251 : 8'b00001111;
												assign node251 = (inp[2]) ? 8'b00001111 : 8'b00011111;
											assign node254 = (inp[2]) ? node258 : node255;
												assign node255 = (inp[12]) ? 8'b00111010 : 8'b00101010;
												assign node258 = (inp[12]) ? node260 : 8'b00011111;
													assign node260 = (inp[6]) ? 8'b00101010 : 8'b00011111;
							assign node263 = (inp[2]) ? node291 : node264;
								assign node264 = (inp[12]) ? node280 : node265;
									assign node265 = (inp[1]) ? node271 : node266;
										assign node266 = (inp[10]) ? 8'b00001111 : node267;
											assign node267 = (inp[0]) ? 8'b00001111 : 8'b00101011;
										assign node271 = (inp[0]) ? 8'b00001011 : node272;
											assign node272 = (inp[3]) ? node276 : node273;
												assign node273 = (inp[9]) ? 8'b00001110 : 8'b00101010;
												assign node276 = (inp[10]) ? 8'b00001011 : 8'b00001111;
									assign node280 = (inp[1]) ? node286 : node281;
										assign node281 = (inp[0]) ? 8'b00011111 : node282;
											assign node282 = (inp[10]) ? 8'b00011111 : 8'b00111011;
										assign node286 = (inp[0]) ? 8'b00011011 : node287;
											assign node287 = (inp[10]) ? 8'b00011011 : 8'b00111010;
								assign node291 = (inp[1]) ? node315 : node292;
									assign node292 = (inp[10]) ? node304 : node293;
										assign node293 = (inp[0]) ? node301 : node294;
											assign node294 = (inp[12]) ? node298 : node295;
												assign node295 = (inp[6]) ? 8'b00101010 : 8'b00111010;
												assign node298 = (inp[6]) ? 8'b00111010 : 8'b00101011;
											assign node301 = (inp[12]) ? 8'b00011110 : 8'b00001110;
										assign node304 = (inp[12]) ? node310 : node305;
											assign node305 = (inp[6]) ? 8'b00001110 : node306;
												assign node306 = (inp[0]) ? 8'b00001110 : 8'b00011110;
											assign node310 = (inp[0]) ? 8'b00011110 : node311;
												assign node311 = (inp[6]) ? 8'b00011110 : 8'b00001111;
									assign node315 = (inp[0]) ? node329 : node316;
										assign node316 = (inp[9]) ? node326 : node317;
											assign node317 = (inp[3]) ? node319 : 8'b00001110;
												assign node319 = (inp[10]) ? 8'b00011010 : node320;
													assign node320 = (inp[12]) ? 8'b00011110 : node321;
														assign node321 = (inp[6]) ? 8'b00001110 : 8'b00011110;
											assign node326 = (inp[12]) ? 8'b00011011 : 8'b00001011;
										assign node329 = (inp[12]) ? 8'b00011010 : 8'b00001010;
				assign node332 = (inp[9]) ? node724 : node333;
					assign node333 = (inp[11]) ? node475 : node334;
						assign node334 = (inp[10]) ? node398 : node335;
							assign node335 = (inp[0]) ? node383 : node336;
								assign node336 = (inp[8]) ? node354 : node337;
									assign node337 = (inp[1]) ? node345 : node338;
										assign node338 = (inp[2]) ? node342 : node339;
											assign node339 = (inp[6]) ? 8'b00101111 : 8'b01111111;
											assign node342 = (inp[3]) ? 8'b00101110 : 8'b00101111;
										assign node345 = (inp[2]) ? node349 : node346;
											assign node346 = (inp[6]) ? 8'b00101110 : 8'b00111110;
											assign node349 = (inp[3]) ? 8'b01111111 : node350;
												assign node350 = (inp[5]) ? 8'b00111110 : 8'b00101110;
									assign node354 = (inp[3]) ? node370 : node355;
										assign node355 = (inp[1]) ? node361 : node356;
											assign node356 = (inp[2]) ? 8'b00101011 : node357;
												assign node357 = (inp[6]) ? 8'b00101011 : 8'b00111011;
											assign node361 = (inp[12]) ? 8'b00101010 : node362;
												assign node362 = (inp[5]) ? node364 : 8'b00111010;
													assign node364 = (inp[6]) ? node366 : 8'b00101010;
														assign node366 = (inp[2]) ? 8'b00111010 : 8'b00101010;
										assign node370 = (inp[5]) ? node372 : 8'b00101010;
											assign node372 = (inp[1]) ? 8'b00111011 : node373;
												assign node373 = (inp[12]) ? node379 : node374;
													assign node374 = (inp[2]) ? 8'b00111010 : node375;
														assign node375 = (inp[6]) ? 8'b00101010 : 8'b00111010;
													assign node379 = (inp[6]) ? 8'b00111010 : 8'b00101010;
								assign node383 = (inp[3]) ? node391 : node384;
									assign node384 = (inp[6]) ? node386 : 8'b01111111;
										assign node386 = (inp[1]) ? 8'b00101111 : node387;
											assign node387 = (inp[5]) ? 8'b01111111 : 8'b00101111;
									assign node391 = (inp[5]) ? node395 : node392;
										assign node392 = (inp[6]) ? 8'b00101110 : 8'b00111110;
										assign node395 = (inp[1]) ? 8'b01111111 : 8'b00111110;
							assign node398 = (inp[5]) ? node420 : node399;
								assign node399 = (inp[6]) ? node415 : node400;
									assign node400 = (inp[3]) ? node410 : node401;
										assign node401 = (inp[0]) ? 8'b00111011 : node402;
											assign node402 = (inp[1]) ? node406 : node403;
												assign node403 = (inp[2]) ? 8'b00101011 : 8'b00111011;
												assign node406 = (inp[2]) ? 8'b00101010 : 8'b00111010;
										assign node410 = (inp[0]) ? 8'b00111010 : node411;
											assign node411 = (inp[2]) ? 8'b00101010 : 8'b00111010;
									assign node415 = (inp[3]) ? 8'b00101010 : node416;
										assign node416 = (inp[0]) ? 8'b00101011 : 8'b00101010;
								assign node420 = (inp[8]) ? node446 : node421;
									assign node421 = (inp[3]) ? node437 : node422;
										assign node422 = (inp[0]) ? node430 : node423;
											assign node423 = (inp[1]) ? node427 : node424;
												assign node424 = (inp[6]) ? 8'b00111011 : 8'b00101011;
												assign node427 = (inp[2]) ? 8'b00101010 : 8'b00111010;
											assign node430 = (inp[1]) ? node432 : 8'b00101011;
												assign node432 = (inp[2]) ? 8'b00111011 : node433;
													assign node433 = (inp[6]) ? 8'b00101011 : 8'b00111011;
										assign node437 = (inp[1]) ? 8'b00111011 : node438;
											assign node438 = (inp[12]) ? 8'b00111010 : node439;
												assign node439 = (inp[6]) ? node441 : 8'b00111010;
													assign node441 = (inp[2]) ? 8'b00111010 : 8'b00101010;
									assign node446 = (inp[0]) ? node466 : node447;
										assign node447 = (inp[12]) ? node457 : node448;
											assign node448 = (inp[1]) ? node450 : 8'b00101110;
												assign node450 = (inp[3]) ? node452 : 8'b00101110;
													assign node452 = (inp[6]) ? node454 : 8'b00101111;
														assign node454 = (inp[2]) ? 8'b01111111 : 8'b00101111;
											assign node457 = (inp[1]) ? node461 : node458;
												assign node458 = (inp[3]) ? 8'b00111110 : 8'b01111111;
												assign node461 = (inp[6]) ? node463 : 8'b00101111;
													assign node463 = (inp[2]) ? 8'b00111110 : 8'b00101110;
										assign node466 = (inp[2]) ? node470 : node467;
											assign node467 = (inp[3]) ? 8'b01111111 : 8'b00101111;
											assign node470 = (inp[3]) ? node472 : 8'b01111111;
												assign node472 = (inp[1]) ? 8'b01111111 : 8'b00111110;
						assign node475 = (inp[8]) ? node599 : node476;
							assign node476 = (inp[10]) ? node538 : node477;
								assign node477 = (inp[0]) ? node511 : node478;
									assign node478 = (inp[3]) ? node496 : node479;
										assign node479 = (inp[1]) ? node487 : node480;
											assign node480 = (inp[2]) ? 8'b00111110 : node481;
												assign node481 = (inp[6]) ? node483 : 8'b01111111;
													assign node483 = (inp[12]) ? 8'b00101111 : 8'b00111110;
											assign node487 = (inp[6]) ? node493 : node488;
												assign node488 = (inp[12]) ? node490 : 8'b00101110;
													assign node490 = (inp[2]) ? 8'b00101110 : 8'b00111110;
												assign node493 = (inp[12]) ? 8'b00101110 : 8'b00111011;
										assign node496 = (inp[1]) ? node500 : node497;
											assign node497 = (inp[12]) ? 8'b00101110 : 8'b00111011;
											assign node500 = (inp[6]) ? node508 : node501;
												assign node501 = (inp[5]) ? node505 : node502;
													assign node502 = (inp[12]) ? 8'b00111110 : 8'b00101110;
													assign node505 = (inp[2]) ? 8'b00111010 : 8'b00111011;
												assign node508 = (inp[12]) ? 8'b00111010 : 8'b00111011;
									assign node511 = (inp[1]) ? node525 : node512;
										assign node512 = (inp[5]) ? node518 : node513;
											assign node513 = (inp[6]) ? node515 : 8'b00111011;
												assign node515 = (inp[3]) ? 8'b00101110 : 8'b00101111;
											assign node518 = (inp[3]) ? node520 : 8'b00111110;
												assign node520 = (inp[2]) ? 8'b00111011 : node521;
													assign node521 = (inp[6]) ? 8'b00111011 : 8'b00101110;
										assign node525 = (inp[2]) ? node533 : node526;
											assign node526 = (inp[3]) ? node528 : 8'b00101011;
												assign node528 = (inp[6]) ? 8'b00111011 : node529;
													assign node529 = (inp[5]) ? 8'b00101011 : 8'b00101110;
											assign node533 = (inp[3]) ? node535 : 8'b00111010;
												assign node535 = (inp[12]) ? 8'b00101110 : 8'b00101010;
								assign node538 = (inp[12]) ? node562 : node539;
									assign node539 = (inp[3]) ? node551 : node540;
										assign node540 = (inp[1]) ? node548 : node541;
											assign node541 = (inp[5]) ? node543 : 8'b00111010;
												assign node543 = (inp[6]) ? node545 : 8'b00101011;
													assign node545 = (inp[2]) ? 8'b00101010 : 8'b00111010;
											assign node548 = (inp[0]) ? 8'b00011110 : 8'b00011111;
										assign node551 = (inp[6]) ? node557 : node552;
											assign node552 = (inp[2]) ? node554 : 8'b00101010;
												assign node554 = (inp[0]) ? 8'b00001111 : 8'b00011111;
											assign node557 = (inp[5]) ? node559 : 8'b00011111;
												assign node559 = (inp[2]) ? 8'b00001110 : 8'b00011111;
									assign node562 = (inp[0]) ? node582 : node563;
										assign node563 = (inp[1]) ? node577 : node564;
											assign node564 = (inp[3]) ? node572 : node565;
												assign node565 = (inp[5]) ? 8'b00111011 : node566;
													assign node566 = (inp[2]) ? 8'b00101011 : node567;
														assign node567 = (inp[6]) ? 8'b00101011 : 8'b00111011;
												assign node572 = (inp[6]) ? 8'b00101010 : node573;
													assign node573 = (inp[2]) ? 8'b00101010 : 8'b00111010;
											assign node577 = (inp[5]) ? node579 : 8'b00101010;
												assign node579 = (inp[3]) ? 8'b00001111 : 8'b00101010;
										assign node582 = (inp[2]) ? node592 : node583;
											assign node583 = (inp[5]) ? 8'b00001111 : node584;
												assign node584 = (inp[3]) ? node588 : node585;
													assign node585 = (inp[6]) ? 8'b00101011 : 8'b00111011;
													assign node588 = (inp[6]) ? 8'b00101010 : 8'b00111010;
											assign node592 = (inp[5]) ? node596 : node593;
												assign node593 = (inp[6]) ? 8'b00101010 : 8'b00011111;
												assign node596 = (inp[1]) ? 8'b00011110 : 8'b00111010;
							assign node599 = (inp[5]) ? node655 : node600;
								assign node600 = (inp[2]) ? node638 : node601;
									assign node601 = (inp[0]) ? node619 : node602;
										assign node602 = (inp[1]) ? node614 : node603;
											assign node603 = (inp[3]) ? node611 : node604;
												assign node604 = (inp[12]) ? node608 : node605;
													assign node605 = (inp[6]) ? 8'b00111010 : 8'b00101011;
													assign node608 = (inp[6]) ? 8'b00101011 : 8'b00111011;
												assign node611 = (inp[12]) ? 8'b00111010 : 8'b00011111;
											assign node614 = (inp[12]) ? node616 : 8'b00101010;
												assign node616 = (inp[6]) ? 8'b00101010 : 8'b00111010;
										assign node619 = (inp[10]) ? node625 : node620;
											assign node620 = (inp[12]) ? 8'b00011011 : node621;
												assign node621 = (inp[3]) ? 8'b00011011 : 8'b00001011;
											assign node625 = (inp[6]) ? node631 : node626;
												assign node626 = (inp[1]) ? 8'b00111010 : node627;
													assign node627 = (inp[12]) ? 8'b00111011 : 8'b00101011;
												assign node631 = (inp[12]) ? node633 : 8'b00011111;
													assign node633 = (inp[3]) ? 8'b00101010 : node634;
														assign node634 = (inp[1]) ? 8'b00001111 : 8'b00101011;
									assign node638 = (inp[12]) ? node646 : node639;
										assign node639 = (inp[3]) ? 8'b00011111 : node640;
											assign node640 = (inp[0]) ? node642 : 8'b00111010;
												assign node642 = (inp[6]) ? 8'b00011110 : 8'b00001110;
										assign node646 = (inp[3]) ? node650 : node647;
											assign node647 = (inp[6]) ? 8'b00001111 : 8'b00011110;
											assign node650 = (inp[6]) ? 8'b00101010 : node651;
												assign node651 = (inp[0]) ? 8'b00011111 : 8'b00101010;
								assign node655 = (inp[3]) ? node691 : node656;
									assign node656 = (inp[10]) ? node674 : node657;
										assign node657 = (inp[0]) ? node667 : node658;
											assign node658 = (inp[1]) ? 8'b00011111 : node659;
												assign node659 = (inp[6]) ? node661 : 8'b00101011;
													assign node661 = (inp[12]) ? 8'b00111010 : node662;
														assign node662 = (inp[2]) ? 8'b00101010 : 8'b00111010;
											assign node667 = (inp[1]) ? node671 : node668;
												assign node668 = (inp[2]) ? 8'b00001110 : 8'b00001111;
												assign node671 = (inp[2]) ? 8'b00001010 : 8'b00011010;
										assign node674 = (inp[0]) ? node684 : node675;
											assign node675 = (inp[12]) ? 8'b00011110 : node676;
												assign node676 = (inp[1]) ? 8'b00001110 : node677;
													assign node677 = (inp[2]) ? node679 : 8'b00011110;
														assign node679 = (inp[6]) ? 8'b00001110 : 8'b00011110;
											assign node684 = (inp[1]) ? 8'b00001011 : node685;
												assign node685 = (inp[12]) ? node687 : 8'b00001111;
													assign node687 = (inp[2]) ? 8'b00011110 : 8'b00011111;
									assign node691 = (inp[10]) ? node713 : node692;
										assign node692 = (inp[0]) ? node700 : node693;
											assign node693 = (inp[6]) ? node697 : node694;
												assign node694 = (inp[2]) ? 8'b00101010 : 8'b00001111;
												assign node697 = (inp[1]) ? 8'b00011110 : 8'b00011111;
											assign node700 = (inp[2]) ? node708 : node701;
												assign node701 = (inp[6]) ? node703 : 8'b00011011;
													assign node703 = (inp[12]) ? 8'b00001110 : node704;
														assign node704 = (inp[1]) ? 8'b00011010 : 8'b00011011;
												assign node708 = (inp[12]) ? 8'b00011010 : node709;
													assign node709 = (inp[1]) ? 8'b00001010 : 8'b00001011;
										assign node713 = (inp[6]) ? node719 : node714;
											assign node714 = (inp[0]) ? node716 : 8'b00011011;
												assign node716 = (inp[1]) ? 8'b00011010 : 8'b00011011;
											assign node719 = (inp[0]) ? node721 : 8'b00001011;
												assign node721 = (inp[12]) ? 8'b00011010 : 8'b00001011;
					assign node724 = (inp[8]) ? node898 : node725;
						assign node725 = (inp[10]) ? node805 : node726;
							assign node726 = (inp[11]) ? node762 : node727;
								assign node727 = (inp[3]) ? node747 : node728;
									assign node728 = (inp[0]) ? node740 : node729;
										assign node729 = (inp[1]) ? node735 : node730;
											assign node730 = (inp[2]) ? node732 : 8'b00011111;
												assign node732 = (inp[6]) ? 8'b00011111 : 8'b00001111;
											assign node735 = (inp[5]) ? 8'b00011110 : node736;
												assign node736 = (inp[2]) ? 8'b00001110 : 8'b00011110;
										assign node740 = (inp[6]) ? node742 : 8'b00011111;
											assign node742 = (inp[5]) ? node744 : 8'b00001111;
												assign node744 = (inp[2]) ? 8'b00011111 : 8'b00001111;
									assign node747 = (inp[6]) ? node755 : node748;
										assign node748 = (inp[0]) ? 8'b00011110 : node749;
											assign node749 = (inp[2]) ? node751 : 8'b00011110;
												assign node751 = (inp[5]) ? 8'b00001111 : 8'b00001110;
										assign node755 = (inp[5]) ? node757 : 8'b00001110;
											assign node757 = (inp[2]) ? node759 : 8'b00001110;
												assign node759 = (inp[12]) ? 8'b00011110 : 8'b00011111;
								assign node762 = (inp[1]) ? node782 : node763;
									assign node763 = (inp[5]) ? node775 : node764;
										assign node764 = (inp[2]) ? node768 : node765;
											assign node765 = (inp[3]) ? 8'b00011110 : 8'b00001111;
											assign node768 = (inp[3]) ? node770 : 8'b00011110;
												assign node770 = (inp[0]) ? node772 : 8'b00011011;
													assign node772 = (inp[12]) ? 8'b00011011 : 8'b00001011;
										assign node775 = (inp[0]) ? node777 : 8'b00001110;
											assign node777 = (inp[6]) ? node779 : 8'b00011111;
												assign node779 = (inp[12]) ? 8'b00001110 : 8'b00011110;
									assign node782 = (inp[2]) ? node796 : node783;
										assign node783 = (inp[0]) ? node789 : node784;
											assign node784 = (inp[3]) ? 8'b00001011 : node785;
												assign node785 = (inp[5]) ? 8'b00001110 : 8'b00011110;
											assign node789 = (inp[6]) ? node793 : node790;
												assign node790 = (inp[12]) ? 8'b00011011 : 8'b00001011;
												assign node793 = (inp[12]) ? 8'b00001011 : 8'b00011011;
										assign node796 = (inp[5]) ? node802 : node797;
											assign node797 = (inp[12]) ? node799 : 8'b00011011;
												assign node799 = (inp[6]) ? 8'b00001110 : 8'b00011011;
											assign node802 = (inp[12]) ? 8'b00011010 : 8'b00001010;
							assign node805 = (inp[3]) ? node851 : node806;
								assign node806 = (inp[1]) ? node830 : node807;
									assign node807 = (inp[6]) ? node819 : node808;
										assign node808 = (inp[11]) ? node814 : node809;
											assign node809 = (inp[2]) ? node811 : 8'b00011011;
												assign node811 = (inp[0]) ? 8'b00011011 : 8'b00001011;
											assign node814 = (inp[12]) ? node816 : 8'b00001011;
												assign node816 = (inp[0]) ? 8'b00011010 : 8'b00011011;
										assign node819 = (inp[12]) ? node825 : node820;
											assign node820 = (inp[11]) ? 8'b00011010 : node821;
												assign node821 = (inp[0]) ? 8'b00001011 : 8'b00011011;
											assign node825 = (inp[2]) ? node827 : 8'b00001011;
												assign node827 = (inp[5]) ? 8'b00011011 : 8'b00001011;
									assign node830 = (inp[0]) ? node844 : node831;
										assign node831 = (inp[6]) ? node839 : node832;
											assign node832 = (inp[2]) ? node836 : node833;
												assign node833 = (inp[11]) ? 8'b00001010 : 8'b00011010;
												assign node836 = (inp[12]) ? 8'b00000010 : 8'b10000010;
											assign node839 = (inp[12]) ? 8'b00000010 : node840;
												assign node840 = (inp[2]) ? 8'b10100101 : 8'b11110111;
										assign node844 = (inp[11]) ? 8'b10100101 : node845;
											assign node845 = (inp[2]) ? node847 : 8'b10011001;
												assign node847 = (inp[6]) ? 8'b10000001 : 8'b10010001;
								assign node851 = (inp[11]) ? node875 : node852;
									assign node852 = (inp[2]) ? node864 : node853;
										assign node853 = (inp[6]) ? node859 : node854;
											assign node854 = (inp[5]) ? node856 : 8'b00011010;
												assign node856 = (inp[1]) ? 8'b10011001 : 8'b00011010;
											assign node859 = (inp[1]) ? 8'b10000001 : node860;
												assign node860 = (inp[5]) ? 8'b10000010 : 8'b00000010;
										assign node864 = (inp[0]) ? node870 : node865;
											assign node865 = (inp[6]) ? 8'b10010000 : node866;
												assign node866 = (inp[12]) ? 8'b00000010 : 8'b10000010;
											assign node870 = (inp[6]) ? node872 : 8'b10010000;
												assign node872 = (inp[1]) ? 8'b10010001 : 8'b10000010;
									assign node875 = (inp[12]) ? node885 : node876;
										assign node876 = (inp[6]) ? node880 : node877;
											assign node877 = (inp[0]) ? 8'b00001010 : 8'b11110111;
											assign node880 = (inp[5]) ? node882 : 8'b11110111;
												assign node882 = (inp[2]) ? 8'b10100101 : 8'b11110111;
										assign node885 = (inp[5]) ? node891 : node886;
											assign node886 = (inp[6]) ? 8'b00000010 : node887;
												assign node887 = (inp[0]) ? 8'b00011010 : 8'b00000010;
											assign node891 = (inp[2]) ? node895 : node892;
												assign node892 = (inp[6]) ? 8'b10100101 : 8'b11111101;
												assign node895 = (inp[1]) ? 8'b10110100 : 8'b11110101;
						assign node898 = (inp[0]) ? node994 : node899;
							assign node899 = (inp[5]) ? node931 : node900;
								assign node900 = (inp[12]) ? node916 : node901;
									assign node901 = (inp[11]) ? node907 : node902;
										assign node902 = (inp[2]) ? 8'b10000010 : node903;
											assign node903 = (inp[6]) ? 8'b10000010 : 8'b00011010;
										assign node907 = (inp[3]) ? 8'b11110111 : node908;
											assign node908 = (inp[2]) ? 8'b11110111 : node909;
												assign node909 = (inp[6]) ? 8'b00011010 : node910;
													assign node910 = (inp[1]) ? 8'b00001010 : 8'b00001011;
									assign node916 = (inp[2]) ? node926 : node917;
										assign node917 = (inp[6]) ? node923 : node918;
											assign node918 = (inp[1]) ? 8'b00011010 : node919;
												assign node919 = (inp[3]) ? 8'b00011010 : 8'b00011011;
											assign node923 = (inp[3]) ? 8'b00000010 : 8'b00001011;
										assign node926 = (inp[1]) ? 8'b00000010 : node927;
											assign node927 = (inp[3]) ? 8'b00000010 : 8'b00001011;
								assign node931 = (inp[10]) ? node963 : node932;
									assign node932 = (inp[1]) ? node948 : node933;
										assign node933 = (inp[3]) ? node941 : node934;
											assign node934 = (inp[11]) ? node936 : 8'b00011011;
												assign node936 = (inp[2]) ? 8'b00011010 : node937;
													assign node937 = (inp[12]) ? 8'b00001011 : 8'b00011010;
											assign node941 = (inp[6]) ? node945 : node942;
												assign node942 = (inp[2]) ? 8'b00000010 : 8'b00011010;
												assign node945 = (inp[2]) ? 8'b10010000 : 8'b11110111;
										assign node948 = (inp[11]) ? node954 : node949;
											assign node949 = (inp[3]) ? 8'b10000001 : node950;
												assign node950 = (inp[12]) ? 8'b10010000 : 8'b10000010;
											assign node954 = (inp[2]) ? node956 : 8'b00001010;
												assign node956 = (inp[3]) ? node960 : node957;
													assign node957 = (inp[12]) ? 8'b11110101 : 8'b11110111;
													assign node960 = (inp[12]) ? 8'b10100101 : 8'b10110100;
									assign node963 = (inp[11]) ? node977 : node964;
										assign node964 = (inp[1]) ? node970 : node965;
											assign node965 = (inp[3]) ? 8'b10011100 : node966;
												assign node966 = (inp[2]) ? 8'b10011101 : 8'b10001101;
											assign node970 = (inp[6]) ? node974 : node971;
												assign node971 = (inp[3]) ? 8'b10000101 : 8'b10000100;
												assign node974 = (inp[12]) ? 8'b10010100 : 8'b10010101;
										assign node977 = (inp[2]) ? node987 : node978;
											assign node978 = (inp[12]) ? node984 : node979;
												assign node979 = (inp[6]) ? 8'b10111100 : node980;
													assign node980 = (inp[1]) ? 8'b10101100 : 8'b10101101;
												assign node984 = (inp[1]) ? 8'b10111100 : 8'b11111101;
											assign node987 = (inp[12]) ? node989 : 8'b10110001;
												assign node989 = (inp[1]) ? node991 : 8'b10100100;
													assign node991 = (inp[3]) ? 8'b10100001 : 8'b10100100;
							assign node994 = (inp[11]) ? node1038 : node995;
								assign node995 = (inp[6]) ? node1019 : node996;
									assign node996 = (inp[3]) ? node1008 : node997;
										assign node997 = (inp[2]) ? node1005 : node998;
											assign node998 = (inp[1]) ? 8'b10011001 : node999;
												assign node999 = (inp[5]) ? 8'b10011101 : node1000;
													assign node1000 = (inp[10]) ? 8'b00011011 : 8'b10011101;
											assign node1005 = (inp[1]) ? 8'b10010101 : 8'b10011101;
										assign node1008 = (inp[2]) ? node1014 : node1009;
											assign node1009 = (inp[1]) ? node1011 : 8'b10011100;
												assign node1011 = (inp[10]) ? 8'b00011010 : 8'b10011100;
											assign node1014 = (inp[12]) ? 8'b10010100 : node1015;
												assign node1015 = (inp[5]) ? 8'b10010101 : 8'b10010000;
									assign node1019 = (inp[5]) ? node1031 : node1020;
										assign node1020 = (inp[3]) ? node1026 : node1021;
											assign node1021 = (inp[1]) ? 8'b10000001 : node1022;
												assign node1022 = (inp[10]) ? 8'b00001011 : 8'b10001101;
											assign node1026 = (inp[10]) ? node1028 : 8'b10000100;
												assign node1028 = (inp[12]) ? 8'b00000010 : 8'b10000010;
										assign node1031 = (inp[1]) ? node1035 : node1032;
											assign node1032 = (inp[3]) ? 8'b10000100 : 8'b10001101;
											assign node1035 = (inp[2]) ? 8'b10010101 : 8'b10000101;
								assign node1038 = (inp[1]) ? node1074 : node1039;
									assign node1039 = (inp[3]) ? node1057 : node1040;
										assign node1040 = (inp[2]) ? node1048 : node1041;
											assign node1041 = (inp[6]) ? node1045 : node1042;
												assign node1042 = (inp[12]) ? 8'b11111101 : 8'b00001011;
												assign node1045 = (inp[12]) ? 8'b10101101 : 8'b10111100;
											assign node1048 = (inp[12]) ? node1054 : node1049;
												assign node1049 = (inp[10]) ? 8'b10101100 : node1050;
													assign node1050 = (inp[6]) ? 8'b10111100 : 8'b10101100;
												assign node1054 = (inp[5]) ? 8'b10111100 : 8'b00011010;
										assign node1057 = (inp[10]) ? node1063 : node1058;
											assign node1058 = (inp[12]) ? 8'b10110001 : node1059;
												assign node1059 = (inp[6]) ? 8'b10110001 : 8'b10100001;
											assign node1063 = (inp[12]) ? node1069 : node1064;
												assign node1064 = (inp[2]) ? node1066 : 8'b10110001;
													assign node1066 = (inp[6]) ? 8'b11110111 : 8'b10100101;
												assign node1069 = (inp[5]) ? 8'b10111100 : node1070;
													assign node1070 = (inp[6]) ? 8'b00000010 : 8'b00011010;
									assign node1074 = (inp[5]) ? node1094 : node1075;
										assign node1075 = (inp[6]) ? node1085 : node1076;
											assign node1076 = (inp[2]) ? node1082 : node1077;
												assign node1077 = (inp[3]) ? node1079 : 8'b10101101;
													assign node1079 = (inp[12]) ? 8'b10111100 : 8'b10101100;
												assign node1082 = (inp[10]) ? 8'b11110101 : 8'b10110001;
											assign node1085 = (inp[12]) ? node1089 : node1086;
												assign node1086 = (inp[3]) ? 8'b11110111 : 8'b10110100;
												assign node1089 = (inp[10]) ? 8'b00000010 : node1090;
													assign node1090 = (inp[3]) ? 8'b10100100 : 8'b10100001;
										assign node1094 = (inp[2]) ? node1102 : node1095;
											assign node1095 = (inp[6]) ? node1099 : node1096;
												assign node1096 = (inp[12]) ? 8'b10111001 : 8'b10101001;
												assign node1099 = (inp[12]) ? 8'b10100001 : 8'b10110000;
											assign node1102 = (inp[12]) ? 8'b10110000 : 8'b10100000;
			assign node1105 = (inp[5]) ? node1651 : node1106;
				assign node1106 = (inp[0]) ? node1256 : node1107;
					assign node1107 = (inp[8]) ? node1189 : node1108;
						assign node1108 = (inp[7]) ? node1132 : node1109;
							assign node1109 = (inp[1]) ? node1121 : node1110;
								assign node1110 = (inp[12]) ? node1118 : node1111;
									assign node1111 = (inp[11]) ? node1115 : node1112;
										assign node1112 = (inp[2]) ? 8'b00001111 : 8'b00011111;
										assign node1115 = (inp[2]) ? 8'b00011110 : 8'b00001111;
									assign node1118 = (inp[2]) ? 8'b00001111 : 8'b00011111;
								assign node1121 = (inp[2]) ? node1127 : node1122;
									assign node1122 = (inp[12]) ? 8'b00011110 : node1123;
										assign node1123 = (inp[11]) ? 8'b00001110 : 8'b00011110;
									assign node1127 = (inp[11]) ? node1129 : 8'b00001110;
										assign node1129 = (inp[12]) ? 8'b00001110 : 8'b00011011;
							assign node1132 = (inp[10]) ? node1160 : node1133;
								assign node1133 = (inp[11]) ? node1147 : node1134;
									assign node1134 = (inp[1]) ? 8'b00001110 : node1135;
										assign node1135 = (inp[3]) ? node1141 : node1136;
											assign node1136 = (inp[2]) ? 8'b00001111 : node1137;
												assign node1137 = (inp[6]) ? 8'b00001111 : 8'b00011111;
											assign node1141 = (inp[6]) ? 8'b00001110 : node1142;
												assign node1142 = (inp[12]) ? 8'b00011110 : 8'b00001110;
									assign node1147 = (inp[12]) ? node1157 : node1148;
										assign node1148 = (inp[3]) ? 8'b00011011 : node1149;
											assign node1149 = (inp[2]) ? node1153 : node1150;
												assign node1150 = (inp[1]) ? 8'b00001110 : 8'b00011110;
												assign node1153 = (inp[1]) ? 8'b00011011 : 8'b00011110;
										assign node1157 = (inp[3]) ? 8'b00001110 : 8'b00001111;
								assign node1160 = (inp[12]) ? node1174 : node1161;
									assign node1161 = (inp[11]) ? node1167 : node1162;
										assign node1162 = (inp[3]) ? 8'b10000010 : node1163;
											assign node1163 = (inp[1]) ? 8'b10000010 : 8'b00001011;
										assign node1167 = (inp[6]) ? 8'b11110111 : node1168;
											assign node1168 = (inp[2]) ? node1170 : 8'b00001010;
												assign node1170 = (inp[9]) ? 8'b11110111 : 8'b00011010;
									assign node1174 = (inp[6]) ? node1184 : node1175;
										assign node1175 = (inp[2]) ? node1181 : node1176;
											assign node1176 = (inp[3]) ? 8'b00011010 : node1177;
												assign node1177 = (inp[9]) ? 8'b00011011 : 8'b00011010;
											assign node1181 = (inp[3]) ? 8'b00000010 : 8'b00001011;
										assign node1184 = (inp[3]) ? 8'b00000010 : node1185;
											assign node1185 = (inp[1]) ? 8'b00000010 : 8'b00001011;
						assign node1189 = (inp[1]) ? node1233 : node1190;
							assign node1190 = (inp[7]) ? node1202 : node1191;
								assign node1191 = (inp[2]) ? node1197 : node1192;
									assign node1192 = (inp[11]) ? node1194 : 8'b00011011;
										assign node1194 = (inp[12]) ? 8'b00011011 : 8'b00001011;
									assign node1197 = (inp[11]) ? node1199 : 8'b00001011;
										assign node1199 = (inp[12]) ? 8'b00001011 : 8'b00011010;
								assign node1202 = (inp[3]) ? node1216 : node1203;
									assign node1203 = (inp[11]) ? node1209 : node1204;
										assign node1204 = (inp[2]) ? 8'b00001011 : node1205;
											assign node1205 = (inp[6]) ? 8'b00001011 : 8'b00011011;
										assign node1209 = (inp[12]) ? node1213 : node1210;
											assign node1210 = (inp[2]) ? 8'b00011010 : 8'b00001011;
											assign node1213 = (inp[2]) ? 8'b00001011 : 8'b00011011;
									assign node1216 = (inp[11]) ? node1224 : node1217;
										assign node1217 = (inp[2]) ? node1221 : node1218;
											assign node1218 = (inp[6]) ? 8'b10000010 : 8'b00011010;
											assign node1221 = (inp[12]) ? 8'b00000010 : 8'b10000010;
										assign node1224 = (inp[12]) ? node1230 : node1225;
											assign node1225 = (inp[2]) ? 8'b11110111 : node1226;
												assign node1226 = (inp[10]) ? 8'b00001010 : 8'b11110111;
											assign node1230 = (inp[2]) ? 8'b00000010 : 8'b00011010;
							assign node1233 = (inp[12]) ? node1249 : node1234;
								assign node1234 = (inp[11]) ? node1242 : node1235;
									assign node1235 = (inp[2]) ? 8'b10000010 : node1236;
										assign node1236 = (inp[6]) ? node1238 : 8'b00011010;
											assign node1238 = (inp[7]) ? 8'b10000010 : 8'b00011010;
									assign node1242 = (inp[2]) ? 8'b11110111 : node1243;
										assign node1243 = (inp[6]) ? node1245 : 8'b00001010;
											assign node1245 = (inp[7]) ? 8'b11110111 : 8'b00001010;
								assign node1249 = (inp[2]) ? 8'b00000010 : node1250;
									assign node1250 = (inp[6]) ? node1252 : 8'b00011010;
										assign node1252 = (inp[7]) ? 8'b00000010 : 8'b00011010;
					assign node1256 = (inp[9]) ? node1452 : node1257;
						assign node1257 = (inp[11]) ? node1333 : node1258;
							assign node1258 = (inp[6]) ? node1296 : node1259;
								assign node1259 = (inp[3]) ? node1277 : node1260;
									assign node1260 = (inp[7]) ? node1270 : node1261;
										assign node1261 = (inp[8]) ? node1263 : 8'b11111101;
											assign node1263 = (inp[10]) ? 8'b10111001 : node1264;
												assign node1264 = (inp[2]) ? node1266 : 8'b11111101;
													assign node1266 = (inp[1]) ? 8'b11110101 : 8'b11111101;
										assign node1270 = (inp[10]) ? node1272 : 8'b11111101;
											assign node1272 = (inp[1]) ? node1274 : 8'b10111001;
												assign node1274 = (inp[2]) ? 8'b10110001 : 8'b10111001;
									assign node1277 = (inp[10]) ? node1287 : node1278;
										assign node1278 = (inp[1]) ? node1282 : node1279;
											assign node1279 = (inp[12]) ? 8'b10110100 : 8'b11111101;
											assign node1282 = (inp[12]) ? node1284 : 8'b10111100;
												assign node1284 = (inp[2]) ? 8'b10110100 : 8'b10111100;
										assign node1287 = (inp[2]) ? node1293 : node1288;
											assign node1288 = (inp[7]) ? 8'b10111000 : node1289;
												assign node1289 = (inp[1]) ? 8'b10111000 : 8'b10111001;
											assign node1293 = (inp[1]) ? 8'b10111100 : 8'b10110000;
								assign node1296 = (inp[10]) ? node1320 : node1297;
									assign node1297 = (inp[3]) ? node1307 : node1298;
										assign node1298 = (inp[2]) ? node1302 : node1299;
											assign node1299 = (inp[7]) ? 8'b10101101 : 8'b11111101;
											assign node1302 = (inp[1]) ? node1304 : 8'b10101101;
												assign node1304 = (inp[8]) ? 8'b10100101 : 8'b10101101;
										assign node1307 = (inp[1]) ? node1313 : node1308;
											assign node1308 = (inp[8]) ? node1310 : 8'b11111101;
												assign node1310 = (inp[7]) ? 8'b10100100 : 8'b10101101;
											assign node1313 = (inp[8]) ? node1315 : 8'b10101100;
												assign node1315 = (inp[2]) ? 8'b10100100 : node1316;
													assign node1316 = (inp[7]) ? 8'b10100100 : 8'b10111100;
									assign node1320 = (inp[7]) ? node1328 : node1321;
										assign node1321 = (inp[2]) ? node1325 : node1322;
											assign node1322 = (inp[1]) ? 8'b10111100 : 8'b10111001;
											assign node1325 = (inp[8]) ? 8'b10101001 : 8'b10101101;
										assign node1328 = (inp[3]) ? 8'b10100000 : node1329;
											assign node1329 = (inp[1]) ? 8'b10100001 : 8'b10101001;
							assign node1333 = (inp[8]) ? node1385 : node1334;
								assign node1334 = (inp[7]) ? node1356 : node1335;
									assign node1335 = (inp[1]) ? node1343 : node1336;
										assign node1336 = (inp[2]) ? node1340 : node1337;
											assign node1337 = (inp[12]) ? 8'b11111101 : 8'b10101101;
											assign node1340 = (inp[3]) ? 8'b10101100 : 8'b10111100;
										assign node1343 = (inp[3]) ? node1349 : node1344;
											assign node1344 = (inp[12]) ? node1346 : 8'b10101001;
												assign node1346 = (inp[2]) ? 8'b10101001 : 8'b10111001;
											assign node1349 = (inp[2]) ? node1353 : node1350;
												assign node1350 = (inp[10]) ? 8'b10101100 : 8'b10111100;
												assign node1353 = (inp[12]) ? 8'b10111001 : 8'b10101001;
									assign node1356 = (inp[10]) ? node1364 : node1357;
										assign node1357 = (inp[1]) ? node1359 : 8'b10101101;
											assign node1359 = (inp[3]) ? 8'b10101100 : node1360;
												assign node1360 = (inp[2]) ? 8'b10111000 : 8'b10101001;
										assign node1364 = (inp[1]) ? node1372 : node1365;
											assign node1365 = (inp[12]) ? node1369 : node1366;
												assign node1366 = (inp[2]) ? 8'b10000101 : 8'b10101000;
												assign node1369 = (inp[6]) ? 8'b10101001 : 8'b10111000;
											assign node1372 = (inp[12]) ? node1378 : node1373;
												assign node1373 = (inp[3]) ? node1375 : 8'b10010100;
													assign node1375 = (inp[6]) ? 8'b10010101 : 8'b10000101;
												assign node1378 = (inp[3]) ? node1382 : node1379;
													assign node1379 = (inp[6]) ? 8'b10000101 : 8'b10011101;
													assign node1382 = (inp[6]) ? 8'b10100000 : 8'b10111000;
								assign node1385 = (inp[1]) ? node1415 : node1386;
									assign node1386 = (inp[10]) ? node1396 : node1387;
										assign node1387 = (inp[7]) ? 8'b10011100 : node1388;
											assign node1388 = (inp[12]) ? node1392 : node1389;
												assign node1389 = (inp[3]) ? 8'b10001100 : 8'b10011100;
												assign node1392 = (inp[2]) ? 8'b10001101 : 8'b10011101;
										assign node1396 = (inp[7]) ? node1404 : node1397;
											assign node1397 = (inp[2]) ? node1399 : 8'b10111001;
												assign node1399 = (inp[12]) ? 8'b10111000 : node1400;
													assign node1400 = (inp[6]) ? 8'b10111000 : 8'b10101000;
											assign node1404 = (inp[3]) ? node1406 : 8'b10111000;
												assign node1406 = (inp[2]) ? node1410 : node1407;
													assign node1407 = (inp[6]) ? 8'b10010101 : 8'b10101000;
													assign node1410 = (inp[6]) ? 8'b10100000 : node1411;
														assign node1411 = (inp[12]) ? 8'b10010101 : 8'b10000101;
									assign node1415 = (inp[2]) ? node1431 : node1416;
										assign node1416 = (inp[10]) ? node1422 : node1417;
											assign node1417 = (inp[3]) ? 8'b10001100 : node1418;
												assign node1418 = (inp[12]) ? 8'b10011001 : 8'b10001001;
											assign node1422 = (inp[6]) ? node1426 : node1423;
												assign node1423 = (inp[3]) ? 8'b10111000 : 8'b10011101;
												assign node1426 = (inp[7]) ? node1428 : 8'b10011101;
													assign node1428 = (inp[12]) ? 8'b10000101 : 8'b10010101;
										assign node1431 = (inp[10]) ? node1445 : node1432;
											assign node1432 = (inp[3]) ? node1440 : node1433;
												assign node1433 = (inp[12]) ? node1437 : node1434;
													assign node1434 = (inp[7]) ? 8'b10010000 : 8'b10000000;
													assign node1437 = (inp[6]) ? 8'b10000001 : 8'b10010000;
												assign node1440 = (inp[12]) ? 8'b10010001 : node1441;
													assign node1441 = (inp[6]) ? 8'b10010001 : 8'b10000001;
											assign node1445 = (inp[3]) ? node1449 : node1446;
												assign node1446 = (inp[6]) ? 8'b10000101 : 8'b10000100;
												assign node1449 = (inp[6]) ? 8'b10100000 : 8'b10010101;
						assign node1452 = (inp[8]) ? node1542 : node1453;
							assign node1453 = (inp[7]) ? node1489 : node1454;
								assign node1454 = (inp[11]) ? node1468 : node1455;
									assign node1455 = (inp[2]) ? node1461 : node1456;
										assign node1456 = (inp[3]) ? node1458 : 8'b00011111;
											assign node1458 = (inp[1]) ? 8'b00011110 : 8'b00011111;
										assign node1461 = (inp[6]) ? 8'b00001111 : node1462;
											assign node1462 = (inp[1]) ? node1464 : 8'b00011111;
												assign node1464 = (inp[10]) ? 8'b00011111 : 8'b00011110;
									assign node1468 = (inp[1]) ? node1476 : node1469;
										assign node1469 = (inp[2]) ? node1473 : node1470;
											assign node1470 = (inp[12]) ? 8'b00011111 : 8'b00001111;
											assign node1473 = (inp[6]) ? 8'b00001111 : 8'b00001110;
										assign node1476 = (inp[3]) ? node1480 : node1477;
											assign node1477 = (inp[12]) ? 8'b00011011 : 8'b00001011;
											assign node1480 = (inp[2]) ? node1484 : node1481;
												assign node1481 = (inp[12]) ? 8'b00011110 : 8'b00001110;
												assign node1484 = (inp[12]) ? 8'b00001110 : node1485;
													assign node1485 = (inp[10]) ? 8'b00011011 : 8'b00001011;
								assign node1489 = (inp[10]) ? node1513 : node1490;
									assign node1490 = (inp[3]) ? node1502 : node1491;
										assign node1491 = (inp[6]) ? node1499 : node1492;
											assign node1492 = (inp[11]) ? node1494 : 8'b00011111;
												assign node1494 = (inp[2]) ? 8'b00001110 : node1495;
													assign node1495 = (inp[12]) ? 8'b00011111 : 8'b00001111;
											assign node1499 = (inp[11]) ? 8'b00001011 : 8'b00001111;
										assign node1502 = (inp[11]) ? node1506 : node1503;
											assign node1503 = (inp[6]) ? 8'b00001110 : 8'b00011110;
											assign node1506 = (inp[12]) ? 8'b00011110 : node1507;
												assign node1507 = (inp[6]) ? 8'b00011011 : node1508;
													assign node1508 = (inp[2]) ? 8'b00001011 : 8'b00001110;
									assign node1513 = (inp[1]) ? node1527 : node1514;
										assign node1514 = (inp[3]) ? node1522 : node1515;
											assign node1515 = (inp[11]) ? node1517 : 8'b00001011;
												assign node1517 = (inp[12]) ? 8'b00011011 : node1518;
													assign node1518 = (inp[6]) ? 8'b00011010 : 8'b00001010;
											assign node1522 = (inp[2]) ? 8'b10010000 : node1523;
												assign node1523 = (inp[6]) ? 8'b10000010 : 8'b00011010;
										assign node1527 = (inp[11]) ? node1535 : node1528;
											assign node1528 = (inp[3]) ? node1532 : node1529;
												assign node1529 = (inp[6]) ? 8'b10000001 : 8'b10010001;
												assign node1532 = (inp[6]) ? 8'b00000010 : 8'b10010000;
											assign node1535 = (inp[3]) ? node1539 : node1536;
												assign node1536 = (inp[2]) ? 8'b10110100 : 8'b11111101;
												assign node1539 = (inp[6]) ? 8'b11110111 : 8'b00011010;
							assign node1542 = (inp[10]) ? node1594 : node1543;
								assign node1543 = (inp[11]) ? node1569 : node1544;
									assign node1544 = (inp[6]) ? node1556 : node1545;
										assign node1545 = (inp[3]) ? node1549 : node1546;
											assign node1546 = (inp[1]) ? 8'b10010101 : 8'b10011101;
											assign node1549 = (inp[7]) ? node1553 : node1550;
												assign node1550 = (inp[1]) ? 8'b10011100 : 8'b10011101;
												assign node1553 = (inp[2]) ? 8'b10010100 : 8'b10011100;
										assign node1556 = (inp[7]) ? node1564 : node1557;
											assign node1557 = (inp[2]) ? node1561 : node1558;
												assign node1558 = (inp[1]) ? 8'b10011100 : 8'b10011101;
												assign node1561 = (inp[3]) ? 8'b10001101 : 8'b10000101;
											assign node1564 = (inp[3]) ? 8'b10000100 : node1565;
												assign node1565 = (inp[1]) ? 8'b10000101 : 8'b10001101;
									assign node1569 = (inp[12]) ? node1579 : node1570;
										assign node1570 = (inp[6]) ? node1576 : node1571;
											assign node1571 = (inp[3]) ? 8'b10101100 : node1572;
												assign node1572 = (inp[1]) ? 8'b10100000 : 8'b10101100;
											assign node1576 = (inp[1]) ? 8'b10110000 : 8'b10111100;
										assign node1579 = (inp[6]) ? node1591 : node1580;
											assign node1580 = (inp[2]) ? node1586 : node1581;
												assign node1581 = (inp[3]) ? 8'b10111100 : node1582;
													assign node1582 = (inp[1]) ? 8'b10111001 : 8'b11111101;
												assign node1586 = (inp[7]) ? 8'b10110001 : node1587;
													assign node1587 = (inp[3]) ? 8'b10111100 : 8'b10110000;
											assign node1591 = (inp[7]) ? 8'b10100100 : 8'b10101101;
								assign node1594 = (inp[1]) ? node1620 : node1595;
									assign node1595 = (inp[7]) ? node1607 : node1596;
										assign node1596 = (inp[2]) ? node1602 : node1597;
											assign node1597 = (inp[12]) ? 8'b00011011 : node1598;
												assign node1598 = (inp[6]) ? 8'b00011011 : 8'b00001011;
											assign node1602 = (inp[12]) ? node1604 : 8'b00001010;
												assign node1604 = (inp[6]) ? 8'b00001011 : 8'b00011011;
										assign node1607 = (inp[6]) ? node1615 : node1608;
											assign node1608 = (inp[3]) ? node1612 : node1609;
												assign node1609 = (inp[11]) ? 8'b00011010 : 8'b00011011;
												assign node1612 = (inp[2]) ? 8'b11110101 : 8'b00011010;
											assign node1615 = (inp[3]) ? 8'b00000010 : node1616;
												assign node1616 = (inp[12]) ? 8'b00001011 : 8'b00011010;
									assign node1620 = (inp[3]) ? node1632 : node1621;
										assign node1621 = (inp[11]) ? node1627 : node1622;
											assign node1622 = (inp[2]) ? node1624 : 8'b10011001;
												assign node1624 = (inp[6]) ? 8'b10000001 : 8'b10010001;
											assign node1627 = (inp[7]) ? node1629 : 8'b11111101;
												assign node1629 = (inp[12]) ? 8'b10110100 : 8'b10100100;
										assign node1632 = (inp[2]) ? node1644 : node1633;
											assign node1633 = (inp[7]) ? node1637 : node1634;
												assign node1634 = (inp[11]) ? 8'b00001010 : 8'b00011010;
												assign node1637 = (inp[12]) ? node1641 : node1638;
													assign node1638 = (inp[11]) ? 8'b11110111 : 8'b10000010;
													assign node1641 = (inp[6]) ? 8'b00000010 : 8'b00011010;
											assign node1644 = (inp[6]) ? node1648 : node1645;
												assign node1645 = (inp[11]) ? 8'b11110101 : 8'b10010000;
												assign node1648 = (inp[12]) ? 8'b00000010 : 8'b10000010;
				assign node1651 = (inp[11]) ? node1909 : node1652;
					assign node1652 = (inp[0]) ? node1854 : node1653;
						assign node1653 = (inp[9]) ? node1753 : node1654;
							assign node1654 = (inp[8]) ? node1700 : node1655;
								assign node1655 = (inp[7]) ? node1673 : node1656;
									assign node1656 = (inp[3]) ? node1668 : node1657;
										assign node1657 = (inp[1]) ? node1663 : node1658;
											assign node1658 = (inp[6]) ? 8'b00011111 : node1659;
												assign node1659 = (inp[10]) ? 8'b00001111 : 8'b00011111;
											assign node1663 = (inp[6]) ? 8'b00011110 : node1664;
												assign node1664 = (inp[2]) ? 8'b00001110 : 8'b00011110;
										assign node1668 = (inp[2]) ? node1670 : 8'b00011111;
											assign node1670 = (inp[6]) ? 8'b00011111 : 8'b00001111;
									assign node1673 = (inp[10]) ? node1687 : node1674;
										assign node1674 = (inp[3]) ? node1678 : node1675;
											assign node1675 = (inp[1]) ? 8'b00011110 : 8'b00011111;
											assign node1678 = (inp[1]) ? node1684 : node1679;
												assign node1679 = (inp[6]) ? 8'b00001110 : node1680;
													assign node1680 = (inp[2]) ? 8'b00001110 : 8'b00011110;
												assign node1684 = (inp[6]) ? 8'b00001111 : 8'b00011111;
										assign node1687 = (inp[1]) ? node1693 : node1688;
											assign node1688 = (inp[6]) ? node1690 : 8'b00011010;
												assign node1690 = (inp[2]) ? 8'b00011011 : 8'b00001011;
											assign node1693 = (inp[6]) ? node1697 : node1694;
												assign node1694 = (inp[12]) ? 8'b00000010 : 8'b00011010;
												assign node1697 = (inp[3]) ? 8'b10000001 : 8'b10010000;
								assign node1700 = (inp[10]) ? node1728 : node1701;
									assign node1701 = (inp[1]) ? node1711 : node1702;
										assign node1702 = (inp[7]) ? node1704 : 8'b00011011;
											assign node1704 = (inp[3]) ? node1706 : 8'b00001011;
												assign node1706 = (inp[6]) ? 8'b10000010 : node1707;
													assign node1707 = (inp[12]) ? 8'b00000010 : 8'b00011010;
										assign node1711 = (inp[3]) ? node1717 : node1712;
											assign node1712 = (inp[2]) ? node1714 : 8'b00011010;
												assign node1714 = (inp[6]) ? 8'b10010000 : 8'b00000010;
											assign node1717 = (inp[7]) ? node1723 : node1718;
												assign node1718 = (inp[2]) ? node1720 : 8'b10011001;
													assign node1720 = (inp[6]) ? 8'b10010001 : 8'b10000001;
												assign node1723 = (inp[12]) ? node1725 : 8'b10000001;
													assign node1725 = (inp[2]) ? 8'b10010001 : 8'b10000001;
									assign node1728 = (inp[6]) ? node1742 : node1729;
										assign node1729 = (inp[2]) ? node1735 : node1730;
											assign node1730 = (inp[12]) ? 8'b10011101 : node1731;
												assign node1731 = (inp[3]) ? 8'b10011101 : 8'b10011100;
											assign node1735 = (inp[1]) ? 8'b10000100 : node1736;
												assign node1736 = (inp[3]) ? node1738 : 8'b10001101;
													assign node1738 = (inp[7]) ? 8'b10000100 : 8'b10001101;
										assign node1742 = (inp[7]) ? node1746 : node1743;
											assign node1743 = (inp[3]) ? 8'b10010101 : 8'b10011101;
											assign node1746 = (inp[2]) ? 8'b10010100 : node1747;
												assign node1747 = (inp[1]) ? node1749 : 8'b10000100;
													assign node1749 = (inp[3]) ? 8'b10000101 : 8'b10000100;
							assign node1753 = (inp[7]) ? node1791 : node1754;
								assign node1754 = (inp[6]) ? node1774 : node1755;
									assign node1755 = (inp[2]) ? node1765 : node1756;
										assign node1756 = (inp[8]) ? node1758 : 8'b11111101;
											assign node1758 = (inp[10]) ? node1762 : node1759;
												assign node1759 = (inp[3]) ? 8'b10111001 : 8'b10111000;
												assign node1762 = (inp[3]) ? 8'b11111101 : 8'b10111100;
										assign node1765 = (inp[3]) ? node1771 : node1766;
											assign node1766 = (inp[8]) ? node1768 : 8'b10101100;
												assign node1768 = (inp[10]) ? 8'b10101101 : 8'b10101001;
											assign node1771 = (inp[8]) ? 8'b10100101 : 8'b10101101;
									assign node1774 = (inp[1]) ? node1780 : node1775;
										assign node1775 = (inp[10]) ? 8'b11111101 : node1776;
											assign node1776 = (inp[8]) ? 8'b10111001 : 8'b11111101;
										assign node1780 = (inp[3]) ? node1786 : node1781;
											assign node1781 = (inp[2]) ? 8'b10110000 : node1782;
												assign node1782 = (inp[10]) ? 8'b10111100 : 8'b10111000;
											assign node1786 = (inp[12]) ? 8'b10110001 : node1787;
												assign node1787 = (inp[8]) ? 8'b11110101 : 8'b11111101;
								assign node1791 = (inp[10]) ? node1825 : node1792;
									assign node1792 = (inp[8]) ? node1810 : node1793;
										assign node1793 = (inp[2]) ? node1797 : node1794;
											assign node1794 = (inp[6]) ? 8'b10101101 : 8'b11111101;
											assign node1797 = (inp[6]) ? node1805 : node1798;
												assign node1798 = (inp[1]) ? node1802 : node1799;
													assign node1799 = (inp[3]) ? 8'b10101100 : 8'b10101101;
													assign node1802 = (inp[3]) ? 8'b10101101 : 8'b10101100;
												assign node1805 = (inp[1]) ? node1807 : 8'b10111100;
													assign node1807 = (inp[3]) ? 8'b11111101 : 8'b10111100;
										assign node1810 = (inp[1]) ? node1820 : node1811;
											assign node1811 = (inp[3]) ? node1817 : node1812;
												assign node1812 = (inp[12]) ? node1814 : 8'b10101001;
													assign node1814 = (inp[6]) ? 8'b10111001 : 8'b10101001;
												assign node1817 = (inp[6]) ? 8'b10100000 : 8'b10111000;
											assign node1820 = (inp[2]) ? node1822 : 8'b10111001;
												assign node1822 = (inp[3]) ? 8'b10100001 : 8'b10110000;
									assign node1825 = (inp[8]) ? node1835 : node1826;
										assign node1826 = (inp[6]) ? node1830 : node1827;
											assign node1827 = (inp[2]) ? 8'b10100000 : 8'b10111000;
											assign node1830 = (inp[2]) ? node1832 : 8'b10100001;
												assign node1832 = (inp[3]) ? 8'b10110001 : 8'b10111001;
										assign node1835 = (inp[2]) ? node1843 : node1836;
											assign node1836 = (inp[6]) ? 8'b10100101 : node1837;
												assign node1837 = (inp[3]) ? node1839 : 8'b10111100;
													assign node1839 = (inp[1]) ? 8'b11111101 : 8'b10111100;
											assign node1843 = (inp[6]) ? node1849 : node1844;
												assign node1844 = (inp[3]) ? node1846 : 8'b10100100;
													assign node1846 = (inp[1]) ? 8'b10100101 : 8'b10100100;
												assign node1849 = (inp[3]) ? 8'b10110100 : node1850;
													assign node1850 = (inp[12]) ? 8'b11111101 : 8'b10110100;
						assign node1854 = (inp[7]) ? node1862 : node1855;
							assign node1855 = (inp[8]) ? node1857 : 8'b11111101;
								assign node1857 = (inp[1]) ? node1859 : 8'b11111101;
									assign node1859 = (inp[2]) ? 8'b11110101 : 8'b11111101;
							assign node1862 = (inp[2]) ? node1894 : node1863;
								assign node1863 = (inp[6]) ? node1879 : node1864;
									assign node1864 = (inp[8]) ? node1874 : node1865;
										assign node1865 = (inp[10]) ? node1869 : node1866;
											assign node1866 = (inp[1]) ? 8'b11111101 : 8'b10111100;
											assign node1869 = (inp[1]) ? 8'b10111001 : node1870;
												assign node1870 = (inp[3]) ? 8'b10111000 : 8'b10111001;
										assign node1874 = (inp[1]) ? 8'b11111101 : node1875;
											assign node1875 = (inp[3]) ? 8'b10111100 : 8'b11111101;
									assign node1879 = (inp[1]) ? node1889 : node1880;
										assign node1880 = (inp[3]) ? node1886 : node1881;
											assign node1881 = (inp[8]) ? 8'b10101101 : node1882;
												assign node1882 = (inp[10]) ? 8'b10101001 : 8'b10101101;
											assign node1886 = (inp[8]) ? 8'b10100100 : 8'b10101100;
										assign node1889 = (inp[8]) ? 8'b10100101 : node1890;
											assign node1890 = (inp[10]) ? 8'b10100001 : 8'b10101101;
								assign node1894 = (inp[1]) ? node1904 : node1895;
									assign node1895 = (inp[3]) ? node1901 : node1896;
										assign node1896 = (inp[10]) ? node1898 : 8'b11111101;
											assign node1898 = (inp[8]) ? 8'b11111101 : 8'b10111001;
										assign node1901 = (inp[8]) ? 8'b10110100 : 8'b10111100;
									assign node1904 = (inp[8]) ? 8'b11110101 : node1905;
										assign node1905 = (inp[10]) ? 8'b10110001 : 8'b11111101;
					assign node1909 = (inp[8]) ? node2133 : node1910;
						assign node1910 = (inp[9]) ? node2022 : node1911;
							assign node1911 = (inp[0]) ? node1977 : node1912;
								assign node1912 = (inp[10]) ? node1950 : node1913;
									assign node1913 = (inp[1]) ? node1931 : node1914;
										assign node1914 = (inp[2]) ? node1922 : node1915;
											assign node1915 = (inp[7]) ? node1919 : node1916;
												assign node1916 = (inp[12]) ? 8'b00011111 : 8'b00001111;
												assign node1919 = (inp[3]) ? 8'b00011011 : 8'b00011110;
											assign node1922 = (inp[6]) ? node1928 : node1923;
												assign node1923 = (inp[7]) ? node1925 : 8'b00001111;
													assign node1925 = (inp[3]) ? 8'b00001110 : 8'b00001111;
												assign node1928 = (inp[12]) ? 8'b00011110 : 8'b00001110;
										assign node1931 = (inp[6]) ? node1937 : node1932;
											assign node1932 = (inp[3]) ? node1934 : 8'b00001110;
												assign node1934 = (inp[2]) ? 8'b00011010 : 8'b00001011;
											assign node1937 = (inp[2]) ? node1947 : node1938;
												assign node1938 = (inp[7]) ? node1942 : node1939;
													assign node1939 = (inp[12]) ? 8'b00011110 : 8'b00001110;
													assign node1942 = (inp[12]) ? 8'b00001011 : node1943;
														assign node1943 = (inp[3]) ? 8'b00011010 : 8'b00011011;
												assign node1947 = (inp[12]) ? 8'b00011011 : 8'b00001011;
									assign node1950 = (inp[7]) ? node1958 : node1951;
										assign node1951 = (inp[1]) ? 8'b00011011 : node1952;
											assign node1952 = (inp[2]) ? 8'b00011110 : node1953;
												assign node1953 = (inp[6]) ? 8'b00001111 : 8'b00011111;
										assign node1958 = (inp[3]) ? node1970 : node1959;
											assign node1959 = (inp[1]) ? node1963 : node1960;
												assign node1960 = (inp[6]) ? 8'b00011010 : 8'b00001011;
												assign node1963 = (inp[12]) ? 8'b00000010 : node1964;
													assign node1964 = (inp[6]) ? 8'b11110111 : node1965;
														assign node1965 = (inp[2]) ? 8'b11110111 : 8'b00001010;
											assign node1970 = (inp[1]) ? node1974 : node1971;
												assign node1971 = (inp[12]) ? 8'b00000010 : 8'b11110111;
												assign node1974 = (inp[6]) ? 8'b10100101 : 8'b10110100;
								assign node1977 = (inp[12]) ? node1995 : node1978;
									assign node1978 = (inp[2]) ? node1988 : node1979;
										assign node1979 = (inp[7]) ? node1983 : node1980;
											assign node1980 = (inp[6]) ? 8'b10101101 : 8'b10101001;
											assign node1983 = (inp[6]) ? 8'b10111000 : node1984;
												assign node1984 = (inp[3]) ? 8'b10101000 : 8'b10101001;
										assign node1988 = (inp[10]) ? node1992 : node1989;
											assign node1989 = (inp[1]) ? 8'b10101000 : 8'b10101001;
											assign node1992 = (inp[7]) ? 8'b10000100 : 8'b10101100;
									assign node1995 = (inp[2]) ? node2011 : node1996;
										assign node1996 = (inp[6]) ? node2008 : node1997;
											assign node1997 = (inp[1]) ? node2005 : node1998;
												assign node1998 = (inp[7]) ? node2000 : 8'b11111101;
													assign node2000 = (inp[10]) ? node2002 : 8'b11111101;
														assign node2002 = (inp[3]) ? 8'b10111000 : 8'b10111001;
												assign node2005 = (inp[7]) ? 8'b10011101 : 8'b10111001;
											assign node2008 = (inp[1]) ? 8'b10000101 : 8'b10101101;
										assign node2011 = (inp[7]) ? node2015 : node2012;
											assign node2012 = (inp[1]) ? 8'b10111000 : 8'b10111100;
											assign node2015 = (inp[1]) ? node2019 : node2016;
												assign node2016 = (inp[6]) ? 8'b10111000 : 8'b10111001;
												assign node2019 = (inp[10]) ? 8'b10010100 : 8'b10111000;
							assign node2022 = (inp[12]) ? node2076 : node2023;
								assign node2023 = (inp[0]) ? node2055 : node2024;
									assign node2024 = (inp[7]) ? node2036 : node2025;
										assign node2025 = (inp[1]) ? node2027 : 8'b10101100;
											assign node2027 = (inp[2]) ? node2031 : node2028;
												assign node2028 = (inp[3]) ? 8'b10101001 : 8'b10101100;
												assign node2031 = (inp[3]) ? 8'b10111000 : node2032;
													assign node2032 = (inp[6]) ? 8'b10101001 : 8'b10111001;
										assign node2036 = (inp[10]) ? node2044 : node2037;
											assign node2037 = (inp[1]) ? node2039 : 8'b10111001;
												assign node2039 = (inp[6]) ? node2041 : 8'b10101001;
													assign node2041 = (inp[3]) ? 8'b10101000 : 8'b10101001;
											assign node2044 = (inp[1]) ? node2050 : node2045;
												assign node2045 = (inp[6]) ? 8'b10101000 : node2046;
													assign node2046 = (inp[2]) ? 8'b10010101 : 8'b10101000;
												assign node2050 = (inp[6]) ? 8'b10010100 : node2051;
													assign node2051 = (inp[3]) ? 8'b10001101 : 8'b10010101;
									assign node2055 = (inp[2]) ? node2067 : node2056;
										assign node2056 = (inp[1]) ? node2062 : node2057;
											assign node2057 = (inp[3]) ? node2059 : 8'b10101001;
												assign node2059 = (inp[7]) ? 8'b10101100 : 8'b10101101;
											assign node2062 = (inp[6]) ? node2064 : 8'b10101001;
												assign node2064 = (inp[10]) ? 8'b10101001 : 8'b10111000;
										assign node2067 = (inp[1]) ? node2071 : node2068;
											assign node2068 = (inp[3]) ? 8'b10101100 : 8'b10101000;
											assign node2071 = (inp[7]) ? node2073 : 8'b10101000;
												assign node2073 = (inp[10]) ? 8'b10000100 : 8'b10101000;
								assign node2076 = (inp[2]) ? node2108 : node2077;
									assign node2077 = (inp[1]) ? node2091 : node2078;
										assign node2078 = (inp[7]) ? node2080 : 8'b11111101;
											assign node2080 = (inp[6]) ? node2084 : node2081;
												assign node2081 = (inp[10]) ? 8'b10111001 : 8'b11111101;
												assign node2084 = (inp[10]) ? node2088 : node2085;
													assign node2085 = (inp[0]) ? 8'b10101101 : 8'b10101100;
													assign node2088 = (inp[3]) ? 8'b10100000 : 8'b10101001;
										assign node2091 = (inp[3]) ? node2099 : node2092;
											assign node2092 = (inp[0]) ? node2096 : node2093;
												assign node2093 = (inp[10]) ? 8'b10111000 : 8'b10111100;
												assign node2096 = (inp[7]) ? 8'b10000101 : 8'b10111001;
											assign node2099 = (inp[10]) ? node2105 : node2100;
												assign node2100 = (inp[6]) ? node2102 : 8'b10111001;
													assign node2102 = (inp[0]) ? 8'b10111001 : 8'b10101001;
												assign node2105 = (inp[7]) ? 8'b10011101 : 8'b10111001;
									assign node2108 = (inp[6]) ? node2120 : node2109;
										assign node2109 = (inp[0]) ? node2117 : node2110;
											assign node2110 = (inp[1]) ? 8'b10101100 : node2111;
												assign node2111 = (inp[7]) ? node2113 : 8'b10101101;
													assign node2113 = (inp[10]) ? 8'b10101001 : 8'b10101101;
											assign node2117 = (inp[1]) ? 8'b10111000 : 8'b10111100;
										assign node2120 = (inp[1]) ? node2126 : node2121;
											assign node2121 = (inp[0]) ? 8'b10111100 : node2122;
												assign node2122 = (inp[10]) ? 8'b10111000 : 8'b10111100;
											assign node2126 = (inp[10]) ? node2130 : node2127;
												assign node2127 = (inp[7]) ? 8'b10111000 : 8'b10111001;
												assign node2130 = (inp[3]) ? 8'b10111000 : 8'b10010100;
						assign node2133 = (inp[1]) ? node2217 : node2134;
							assign node2134 = (inp[0]) ? node2188 : node2135;
								assign node2135 = (inp[10]) ? node2159 : node2136;
									assign node2136 = (inp[9]) ? node2152 : node2137;
										assign node2137 = (inp[3]) ? node2147 : node2138;
											assign node2138 = (inp[2]) ? node2144 : node2139;
												assign node2139 = (inp[7]) ? 8'b00001011 : node2140;
													assign node2140 = (inp[12]) ? 8'b00011011 : 8'b00001011;
												assign node2144 = (inp[6]) ? 8'b00011010 : 8'b00001011;
											assign node2147 = (inp[7]) ? node2149 : 8'b00001011;
												assign node2149 = (inp[6]) ? 8'b00000010 : 8'b11110111;
										assign node2152 = (inp[7]) ? 8'b10010101 : node2153;
											assign node2153 = (inp[2]) ? 8'b10111000 : node2154;
												assign node2154 = (inp[12]) ? 8'b10111001 : 8'b10101001;
									assign node2159 = (inp[9]) ? node2177 : node2160;
										assign node2160 = (inp[12]) ? node2174 : node2161;
											assign node2161 = (inp[2]) ? node2165 : node2162;
												assign node2162 = (inp[7]) ? 8'b10101100 : 8'b10101101;
												assign node2165 = (inp[3]) ? node2169 : node2166;
													assign node2166 = (inp[6]) ? 8'b10101100 : 8'b10111100;
													assign node2169 = (inp[7]) ? node2171 : 8'b10101100;
														assign node2171 = (inp[6]) ? 8'b10100001 : 8'b10110001;
											assign node2174 = (inp[2]) ? 8'b10101101 : 8'b11111101;
										assign node2177 = (inp[7]) ? node2185 : node2178;
											assign node2178 = (inp[2]) ? node2182 : node2179;
												assign node2179 = (inp[12]) ? 8'b10011101 : 8'b10001101;
												assign node2182 = (inp[6]) ? 8'b10001100 : 8'b10011100;
											assign node2185 = (inp[12]) ? 8'b10001101 : 8'b10010001;
								assign node2188 = (inp[12]) ? node2204 : node2189;
									assign node2189 = (inp[3]) ? node2197 : node2190;
										assign node2190 = (inp[2]) ? 8'b10001100 : node2191;
											assign node2191 = (inp[7]) ? node2193 : 8'b10001101;
												assign node2193 = (inp[6]) ? 8'b10011100 : 8'b10001101;
										assign node2197 = (inp[7]) ? node2201 : node2198;
											assign node2198 = (inp[10]) ? 8'b10001100 : 8'b10001101;
											assign node2201 = (inp[2]) ? 8'b10000001 : 8'b10010001;
									assign node2204 = (inp[2]) ? node2212 : node2205;
										assign node2205 = (inp[7]) ? node2207 : 8'b10011101;
											assign node2207 = (inp[3]) ? 8'b10000100 : node2208;
												assign node2208 = (inp[6]) ? 8'b10001101 : 8'b10011101;
										assign node2212 = (inp[3]) ? node2214 : 8'b10011100;
											assign node2214 = (inp[7]) ? 8'b10010001 : 8'b10011100;
							assign node2217 = (inp[2]) ? node2265 : node2218;
								assign node2218 = (inp[0]) ? node2256 : node2219;
									assign node2219 = (inp[3]) ? node2241 : node2220;
										assign node2220 = (inp[9]) ? node2232 : node2221;
											assign node2221 = (inp[10]) ? node2229 : node2222;
												assign node2222 = (inp[6]) ? node2226 : node2223;
													assign node2223 = (inp[12]) ? 8'b00011010 : 8'b00001010;
													assign node2226 = (inp[7]) ? 8'b00000010 : 8'b00001010;
												assign node2229 = (inp[7]) ? 8'b10100100 : 8'b10101100;
											assign node2232 = (inp[7]) ? node2238 : node2233;
												assign node2233 = (inp[10]) ? 8'b10011100 : node2234;
													assign node2234 = (inp[6]) ? 8'b10111000 : 8'b10101000;
												assign node2238 = (inp[12]) ? 8'b10100000 : 8'b10010101;
										assign node2241 = (inp[9]) ? node2251 : node2242;
											assign node2242 = (inp[12]) ? node2248 : node2243;
												assign node2243 = (inp[6]) ? node2245 : 8'b10101101;
													assign node2245 = (inp[10]) ? 8'b10110000 : 8'b10110100;
												assign node2248 = (inp[10]) ? 8'b10111001 : 8'b11111101;
											assign node2251 = (inp[6]) ? node2253 : 8'b10001001;
												assign node2253 = (inp[12]) ? 8'b10000101 : 8'b10001101;
									assign node2256 = (inp[7]) ? node2260 : node2257;
										assign node2257 = (inp[12]) ? 8'b10011001 : 8'b10001001;
										assign node2260 = (inp[12]) ? node2262 : 8'b10010000;
											assign node2262 = (inp[6]) ? 8'b10000001 : 8'b10011001;
								assign node2265 = (inp[0]) ? node2305 : node2266;
									assign node2266 = (inp[9]) ? node2288 : node2267;
										assign node2267 = (inp[10]) ? node2273 : node2268;
											assign node2268 = (inp[12]) ? 8'b00000010 : node2269;
												assign node2269 = (inp[7]) ? 8'b10100101 : 8'b10100100;
											assign node2273 = (inp[3]) ? node2283 : node2274;
												assign node2274 = (inp[7]) ? node2278 : node2275;
													assign node2275 = (inp[12]) ? 8'b10100100 : 8'b10110001;
													assign node2278 = (inp[12]) ? 8'b10110001 : node2279;
														assign node2279 = (inp[6]) ? 8'b10100001 : 8'b10110001;
												assign node2283 = (inp[12]) ? 8'b10100001 : node2284;
													assign node2284 = (inp[7]) ? 8'b10100000 : 8'b10110000;
										assign node2288 = (inp[10]) ? node2296 : node2289;
											assign node2289 = (inp[3]) ? node2291 : 8'b10000101;
												assign node2291 = (inp[7]) ? node2293 : 8'b10010100;
													assign node2293 = (inp[12]) ? 8'b10000101 : 8'b10010100;
											assign node2296 = (inp[12]) ? node2302 : node2297;
												assign node2297 = (inp[6]) ? node2299 : 8'b10010001;
													assign node2299 = (inp[7]) ? 8'b10000001 : 8'b10000000;
												assign node2302 = (inp[6]) ? 8'b10010000 : 8'b10000100;
									assign node2305 = (inp[12]) ? 8'b10010000 : 8'b10000000;
		assign node2308 = (inp[7]) ? node3822 : node2309;
			assign node2309 = (inp[13]) ? node3061 : node2310;
				assign node2310 = (inp[9]) ? node2700 : node2311;
					assign node2311 = (inp[8]) ? node2501 : node2312;
						assign node2312 = (inp[10]) ? node2408 : node2313;
							assign node2313 = (inp[1]) ? node2363 : node2314;
								assign node2314 = (inp[3]) ? node2334 : node2315;
									assign node2315 = (inp[12]) ? node2327 : node2316;
										assign node2316 = (inp[11]) ? node2322 : node2317;
											assign node2317 = (inp[6]) ? node2319 : 8'b10000010;
												assign node2319 = (inp[5]) ? 8'b10010000 : 8'b00011010;
											assign node2322 = (inp[2]) ? node2324 : 8'b11110111;
												assign node2324 = (inp[0]) ? 8'b10100101 : 8'b11110111;
										assign node2327 = (inp[6]) ? node2329 : 8'b00000010;
											assign node2329 = (inp[2]) ? node2331 : 8'b00011010;
												assign node2331 = (inp[5]) ? 8'b10010000 : 8'b00000010;
									assign node2334 = (inp[12]) ? node2354 : node2335;
										assign node2335 = (inp[11]) ? node2343 : node2336;
											assign node2336 = (inp[6]) ? node2338 : 8'b00001011;
												assign node2338 = (inp[0]) ? node2340 : 8'b00011011;
													assign node2340 = (inp[2]) ? 8'b00001011 : 8'b00011011;
											assign node2343 = (inp[6]) ? node2349 : node2344;
												assign node2344 = (inp[2]) ? node2346 : 8'b00011010;
													assign node2346 = (inp[0]) ? 8'b00001010 : 8'b00011010;
												assign node2349 = (inp[2]) ? node2351 : 8'b00001011;
													assign node2351 = (inp[5]) ? 8'b00001010 : 8'b00011010;
										assign node2354 = (inp[6]) ? node2358 : node2355;
											assign node2355 = (inp[2]) ? 8'b00011011 : 8'b00001011;
											assign node2358 = (inp[2]) ? node2360 : 8'b00011011;
												assign node2360 = (inp[5]) ? 8'b00011011 : 8'b00001011;
								assign node2363 = (inp[11]) ? node2389 : node2364;
									assign node2364 = (inp[6]) ? node2378 : node2365;
										assign node2365 = (inp[0]) ? node2369 : node2366;
											assign node2366 = (inp[12]) ? 8'b00000010 : 8'b10000010;
											assign node2369 = (inp[2]) ? node2375 : node2370;
												assign node2370 = (inp[5]) ? 8'b10000001 : node2371;
													assign node2371 = (inp[3]) ? 8'b00000010 : 8'b10000001;
												assign node2375 = (inp[5]) ? 8'b10010001 : 8'b10010000;
										assign node2378 = (inp[2]) ? node2384 : node2379;
											assign node2379 = (inp[0]) ? 8'b10011001 : node2380;
												assign node2380 = (inp[3]) ? 8'b10011001 : 8'b00011010;
											assign node2384 = (inp[5]) ? node2386 : 8'b00000010;
												assign node2386 = (inp[12]) ? 8'b10010001 : 8'b10010000;
									assign node2389 = (inp[12]) ? node2399 : node2390;
										assign node2390 = (inp[2]) ? node2392 : 8'b11110111;
											assign node2392 = (inp[3]) ? node2396 : node2393;
												assign node2393 = (inp[5]) ? 8'b10100101 : 8'b10110100;
												assign node2396 = (inp[6]) ? 8'b11110111 : 8'b10100101;
										assign node2399 = (inp[5]) ? node2405 : node2400;
											assign node2400 = (inp[0]) ? node2402 : 8'b00000010;
												assign node2402 = (inp[6]) ? 8'b00011010 : 8'b10100101;
											assign node2405 = (inp[2]) ? 8'b10110100 : 8'b11111101;
							assign node2408 = (inp[11]) ? node2450 : node2409;
								assign node2409 = (inp[3]) ? node2429 : node2410;
									assign node2410 = (inp[6]) ? node2422 : node2411;
										assign node2411 = (inp[2]) ? node2417 : node2412;
											assign node2412 = (inp[1]) ? node2414 : 8'b00001110;
												assign node2414 = (inp[0]) ? 8'b00001111 : 8'b00001110;
											assign node2417 = (inp[0]) ? node2419 : 8'b00001110;
												assign node2419 = (inp[1]) ? 8'b00011111 : 8'b00011110;
										assign node2422 = (inp[2]) ? 8'b00001110 : node2423;
											assign node2423 = (inp[1]) ? node2425 : 8'b00011110;
												assign node2425 = (inp[0]) ? 8'b00011111 : 8'b00011110;
									assign node2429 = (inp[1]) ? node2441 : node2430;
										assign node2430 = (inp[6]) ? node2436 : node2431;
											assign node2431 = (inp[2]) ? node2433 : 8'b00001111;
												assign node2433 = (inp[0]) ? 8'b00011111 : 8'b00001111;
											assign node2436 = (inp[5]) ? 8'b00011111 : node2437;
												assign node2437 = (inp[2]) ? 8'b00001111 : 8'b00011111;
										assign node2441 = (inp[5]) ? node2445 : node2442;
											assign node2442 = (inp[2]) ? 8'b00001110 : 8'b00011110;
											assign node2445 = (inp[6]) ? 8'b00011111 : node2446;
												assign node2446 = (inp[0]) ? 8'b00011111 : 8'b00001111;
								assign node2450 = (inp[1]) ? node2474 : node2451;
									assign node2451 = (inp[12]) ? node2461 : node2452;
										assign node2452 = (inp[6]) ? node2454 : 8'b00011011;
											assign node2454 = (inp[5]) ? 8'b00001110 : node2455;
												assign node2455 = (inp[2]) ? 8'b00011011 : node2456;
													assign node2456 = (inp[3]) ? 8'b00001111 : 8'b00001110;
										assign node2461 = (inp[6]) ? node2469 : node2462;
											assign node2462 = (inp[5]) ? node2466 : node2463;
												assign node2463 = (inp[2]) ? 8'b00011110 : 8'b00001110;
												assign node2466 = (inp[3]) ? 8'b00001111 : 8'b00001110;
											assign node2469 = (inp[0]) ? 8'b00011110 : node2470;
												assign node2470 = (inp[2]) ? 8'b00001110 : 8'b00011110;
									assign node2474 = (inp[0]) ? node2484 : node2475;
										assign node2475 = (inp[12]) ? node2479 : node2476;
											assign node2476 = (inp[6]) ? 8'b00001011 : 8'b00011010;
											assign node2479 = (inp[5]) ? node2481 : 8'b00001110;
												assign node2481 = (inp[6]) ? 8'b00011110 : 8'b00001110;
										assign node2484 = (inp[2]) ? node2490 : node2485;
											assign node2485 = (inp[12]) ? node2487 : 8'b00011010;
												assign node2487 = (inp[6]) ? 8'b00011011 : 8'b00001011;
											assign node2490 = (inp[3]) ? node2498 : node2491;
												assign node2491 = (inp[12]) ? node2493 : 8'b00001010;
													assign node2493 = (inp[5]) ? 8'b00011010 : node2494;
														assign node2494 = (inp[6]) ? 8'b00001011 : 8'b00011010;
												assign node2498 = (inp[12]) ? 8'b00001110 : 8'b00001011;
						assign node2501 = (inp[11]) ? node2601 : node2502;
							assign node2502 = (inp[0]) ? node2548 : node2503;
								assign node2503 = (inp[6]) ? node2521 : node2504;
									assign node2504 = (inp[3]) ? node2514 : node2505;
										assign node2505 = (inp[10]) ? node2509 : node2506;
											assign node2506 = (inp[12]) ? 8'b00000010 : 8'b10000010;
											assign node2509 = (inp[5]) ? 8'b10000100 : node2510;
												assign node2510 = (inp[12]) ? 8'b00000010 : 8'b10000010;
										assign node2514 = (inp[1]) ? 8'b10000010 : node2515;
											assign node2515 = (inp[10]) ? node2517 : 8'b00001011;
												assign node2517 = (inp[12]) ? 8'b00001011 : 8'b10001101;
									assign node2521 = (inp[5]) ? node2535 : node2522;
										assign node2522 = (inp[2]) ? node2528 : node2523;
											assign node2523 = (inp[1]) ? 8'b00011010 : node2524;
												assign node2524 = (inp[3]) ? 8'b00011011 : 8'b00011010;
											assign node2528 = (inp[1]) ? node2532 : node2529;
												assign node2529 = (inp[3]) ? 8'b00001011 : 8'b00000010;
												assign node2532 = (inp[3]) ? 8'b10000010 : 8'b00000010;
										assign node2535 = (inp[10]) ? node2543 : node2536;
											assign node2536 = (inp[2]) ? node2538 : 8'b00011010;
												assign node2538 = (inp[3]) ? node2540 : 8'b10010000;
													assign node2540 = (inp[1]) ? 8'b10010001 : 8'b00011011;
											assign node2543 = (inp[2]) ? 8'b10010101 : node2544;
												assign node2544 = (inp[3]) ? 8'b10011101 : 8'b10011100;
								assign node2548 = (inp[5]) ? node2580 : node2549;
									assign node2549 = (inp[10]) ? node2569 : node2550;
										assign node2550 = (inp[2]) ? node2560 : node2551;
											assign node2551 = (inp[6]) ? 8'b10011101 : node2552;
												assign node2552 = (inp[12]) ? node2554 : 8'b10001101;
													assign node2554 = (inp[1]) ? node2556 : 8'b10000100;
														assign node2556 = (inp[3]) ? 8'b10000100 : 8'b10000101;
											assign node2560 = (inp[6]) ? node2566 : node2561;
												assign node2561 = (inp[1]) ? node2563 : 8'b10010100;
													assign node2563 = (inp[3]) ? 8'b10010100 : 8'b10010101;
												assign node2566 = (inp[3]) ? 8'b10000100 : 8'b10000101;
										assign node2569 = (inp[6]) ? node2577 : node2570;
											assign node2570 = (inp[1]) ? node2574 : node2571;
												assign node2571 = (inp[2]) ? 8'b10010000 : 8'b00000010;
												assign node2574 = (inp[2]) ? 8'b10010001 : 8'b10000001;
											assign node2577 = (inp[12]) ? 8'b00000010 : 8'b00011010;
									assign node2580 = (inp[6]) ? node2592 : node2581;
										assign node2581 = (inp[2]) ? node2589 : node2582;
											assign node2582 = (inp[3]) ? node2586 : node2583;
												assign node2583 = (inp[1]) ? 8'b10000101 : 8'b10000100;
												assign node2586 = (inp[1]) ? 8'b10000101 : 8'b10001101;
											assign node2589 = (inp[1]) ? 8'b10010101 : 8'b10010100;
										assign node2592 = (inp[2]) ? node2598 : node2593;
											assign node2593 = (inp[12]) ? 8'b10011101 : node2594;
												assign node2594 = (inp[3]) ? 8'b10011101 : 8'b10011100;
											assign node2598 = (inp[1]) ? 8'b10010101 : 8'b10011101;
							assign node2601 = (inp[0]) ? node2641 : node2602;
								assign node2602 = (inp[5]) ? node2612 : node2603;
									assign node2603 = (inp[12]) ? node2609 : node2604;
										assign node2604 = (inp[1]) ? 8'b11110111 : node2605;
											assign node2605 = (inp[3]) ? 8'b00011010 : 8'b11110111;
										assign node2609 = (inp[6]) ? 8'b00011011 : 8'b00000010;
									assign node2612 = (inp[3]) ? node2624 : node2613;
										assign node2613 = (inp[2]) ? node2617 : node2614;
											assign node2614 = (inp[1]) ? 8'b00001010 : 8'b10100100;
											assign node2617 = (inp[10]) ? 8'b10110001 : node2618;
												assign node2618 = (inp[6]) ? node2620 : 8'b11110111;
													assign node2620 = (inp[12]) ? 8'b11110101 : 8'b10100101;
										assign node2624 = (inp[1]) ? node2632 : node2625;
											assign node2625 = (inp[10]) ? node2627 : 8'b00011010;
												assign node2627 = (inp[6]) ? node2629 : 8'b10111100;
													assign node2629 = (inp[2]) ? 8'b10111100 : 8'b11111101;
											assign node2632 = (inp[2]) ? node2638 : node2633;
												assign node2633 = (inp[10]) ? node2635 : 8'b11111101;
													assign node2635 = (inp[6]) ? 8'b10111001 : 8'b10100001;
												assign node2638 = (inp[10]) ? 8'b10110000 : 8'b10110100;
								assign node2641 = (inp[1]) ? node2669 : node2642;
									assign node2642 = (inp[3]) ? node2660 : node2643;
										assign node2643 = (inp[2]) ? node2655 : node2644;
											assign node2644 = (inp[6]) ? node2650 : node2645;
												assign node2645 = (inp[12]) ? 8'b10100100 : node2646;
													assign node2646 = (inp[10]) ? 8'b11110111 : 8'b10110001;
												assign node2650 = (inp[10]) ? 8'b00011010 : node2651;
													assign node2651 = (inp[12]) ? 8'b10111100 : 8'b10101100;
											assign node2655 = (inp[10]) ? node2657 : 8'b10110001;
												assign node2657 = (inp[12]) ? 8'b10110001 : 8'b10100001;
										assign node2660 = (inp[5]) ? node2662 : 8'b00001011;
											assign node2662 = (inp[2]) ? 8'b10101100 : node2663;
												assign node2663 = (inp[6]) ? node2665 : 8'b10101101;
													assign node2665 = (inp[12]) ? 8'b11111101 : 8'b10101101;
									assign node2669 = (inp[5]) ? node2685 : node2670;
										assign node2670 = (inp[10]) ? node2680 : node2671;
											assign node2671 = (inp[6]) ? 8'b10111100 : node2672;
												assign node2672 = (inp[3]) ? 8'b10110001 : node2673;
													assign node2673 = (inp[12]) ? 8'b10110000 : node2674;
														assign node2674 = (inp[2]) ? 8'b10100000 : 8'b10110000;
											assign node2680 = (inp[6]) ? node2682 : 8'b10100101;
												assign node2682 = (inp[12]) ? 8'b10100101 : 8'b10110100;
										assign node2685 = (inp[3]) ? node2695 : node2686;
											assign node2686 = (inp[2]) ? node2692 : node2687;
												assign node2687 = (inp[6]) ? 8'b10101001 : node2688;
													assign node2688 = (inp[12]) ? 8'b10100001 : 8'b10110000;
												assign node2692 = (inp[12]) ? 8'b10110000 : 8'b10100000;
											assign node2695 = (inp[6]) ? node2697 : 8'b10110000;
												assign node2697 = (inp[12]) ? 8'b10110000 : 8'b10100000;
					assign node2700 = (inp[11]) ? node2842 : node2701;
						assign node2701 = (inp[5]) ? node2797 : node2702;
							assign node2702 = (inp[0]) ? node2730 : node2703;
								assign node2703 = (inp[2]) ? node2721 : node2704;
									assign node2704 = (inp[6]) ? node2712 : node2705;
										assign node2705 = (inp[8]) ? node2709 : node2706;
											assign node2706 = (inp[12]) ? 8'b00101110 : 8'b00101010;
											assign node2709 = (inp[12]) ? 8'b00101011 : 8'b00101010;
										assign node2712 = (inp[3]) ? node2718 : node2713;
											assign node2713 = (inp[8]) ? 8'b00111010 : node2714;
												assign node2714 = (inp[10]) ? 8'b00111110 : 8'b00111010;
											assign node2718 = (inp[1]) ? 8'b00111110 : 8'b00111011;
									assign node2721 = (inp[8]) ? node2725 : node2722;
										assign node2722 = (inp[10]) ? 8'b00101110 : 8'b00101010;
										assign node2725 = (inp[3]) ? node2727 : 8'b00101010;
											assign node2727 = (inp[1]) ? 8'b00101010 : 8'b00101011;
								assign node2730 = (inp[8]) ? node2758 : node2731;
									assign node2731 = (inp[10]) ? node2747 : node2732;
										assign node2732 = (inp[3]) ? node2736 : node2733;
											assign node2733 = (inp[1]) ? 8'b00101011 : 8'b00101010;
											assign node2736 = (inp[1]) ? node2740 : node2737;
												assign node2737 = (inp[6]) ? 8'b00111011 : 8'b00101011;
												assign node2740 = (inp[6]) ? node2744 : node2741;
													assign node2741 = (inp[2]) ? 8'b00111010 : 8'b00101010;
													assign node2744 = (inp[2]) ? 8'b00101010 : 8'b00111010;
										assign node2747 = (inp[2]) ? node2755 : node2748;
											assign node2748 = (inp[6]) ? node2752 : node2749;
												assign node2749 = (inp[12]) ? 8'b00101111 : 8'b00101110;
												assign node2752 = (inp[3]) ? 8'b00111110 : 8'b01111111;
											assign node2755 = (inp[6]) ? 8'b00101110 : 8'b00111110;
									assign node2758 = (inp[10]) ? node2782 : node2759;
										assign node2759 = (inp[12]) ? node2771 : node2760;
											assign node2760 = (inp[1]) ? node2764 : node2761;
												assign node2761 = (inp[2]) ? 8'b00101111 : 8'b01111111;
												assign node2764 = (inp[3]) ? 8'b00101110 : node2765;
													assign node2765 = (inp[2]) ? node2767 : 8'b00101111;
														assign node2767 = (inp[6]) ? 8'b00101111 : 8'b01111111;
											assign node2771 = (inp[3]) ? node2773 : 8'b00111110;
												assign node2773 = (inp[1]) ? node2775 : 8'b00101111;
													assign node2775 = (inp[6]) ? node2779 : node2776;
														assign node2776 = (inp[2]) ? 8'b00111110 : 8'b00101110;
														assign node2779 = (inp[2]) ? 8'b00101110 : 8'b00111110;
										assign node2782 = (inp[3]) ? node2794 : node2783;
											assign node2783 = (inp[1]) ? node2787 : node2784;
												assign node2784 = (inp[2]) ? 8'b00111010 : 8'b00101010;
												assign node2787 = (inp[12]) ? node2789 : 8'b00101011;
													assign node2789 = (inp[2]) ? 8'b00111011 : node2790;
														assign node2790 = (inp[6]) ? 8'b00111011 : 8'b00101011;
											assign node2794 = (inp[1]) ? 8'b00111010 : 8'b00111011;
							assign node2797 = (inp[6]) ? node2825 : node2798;
								assign node2798 = (inp[10]) ? node2812 : node2799;
									assign node2799 = (inp[0]) ? node2803 : node2800;
										assign node2800 = (inp[3]) ? 8'b00101011 : 8'b00101010;
										assign node2803 = (inp[8]) ? node2809 : node2804;
											assign node2804 = (inp[2]) ? node2806 : 8'b00101011;
												assign node2806 = (inp[1]) ? 8'b00111011 : 8'b00111010;
											assign node2809 = (inp[2]) ? 8'b01111111 : 8'b00101111;
									assign node2812 = (inp[2]) ? node2818 : node2813;
										assign node2813 = (inp[3]) ? 8'b00101111 : node2814;
											assign node2814 = (inp[1]) ? 8'b00101111 : 8'b00101110;
										assign node2818 = (inp[0]) ? node2820 : 8'b00101110;
											assign node2820 = (inp[12]) ? 8'b01111111 : node2821;
												assign node2821 = (inp[3]) ? 8'b01111111 : 8'b00111110;
								assign node2825 = (inp[3]) ? node2837 : node2826;
									assign node2826 = (inp[10]) ? node2832 : node2827;
										assign node2827 = (inp[0]) ? node2829 : 8'b00111010;
											assign node2829 = (inp[8]) ? 8'b01111111 : 8'b00111011;
										assign node2832 = (inp[1]) ? node2834 : 8'b00111110;
											assign node2834 = (inp[0]) ? 8'b01111111 : 8'b00111110;
									assign node2837 = (inp[10]) ? 8'b01111111 : node2838;
										assign node2838 = (inp[8]) ? 8'b01111111 : 8'b00111011;
						assign node2842 = (inp[8]) ? node2944 : node2843;
							assign node2843 = (inp[10]) ? node2901 : node2844;
								assign node2844 = (inp[1]) ? node2874 : node2845;
									assign node2845 = (inp[3]) ? node2859 : node2846;
										assign node2846 = (inp[2]) ? node2854 : node2847;
											assign node2847 = (inp[6]) ? node2851 : node2848;
												assign node2848 = (inp[12]) ? 8'b00101010 : 8'b00011111;
												assign node2851 = (inp[12]) ? 8'b00111010 : 8'b00101010;
											assign node2854 = (inp[12]) ? node2856 : 8'b00011111;
												assign node2856 = (inp[5]) ? 8'b00011111 : 8'b00101010;
										assign node2859 = (inp[12]) ? node2867 : node2860;
											assign node2860 = (inp[6]) ? node2862 : 8'b00111010;
												assign node2862 = (inp[2]) ? node2864 : 8'b00101011;
													assign node2864 = (inp[5]) ? 8'b00101010 : 8'b00111010;
											assign node2867 = (inp[0]) ? node2869 : 8'b00101011;
												assign node2869 = (inp[5]) ? 8'b00111010 : node2870;
													assign node2870 = (inp[6]) ? 8'b00111011 : 8'b00101011;
									assign node2874 = (inp[12]) ? node2890 : node2875;
										assign node2875 = (inp[0]) ? node2881 : node2876;
											assign node2876 = (inp[6]) ? node2878 : 8'b00011111;
												assign node2878 = (inp[2]) ? 8'b00001111 : 8'b00101010;
											assign node2881 = (inp[5]) ? node2887 : node2882;
												assign node2882 = (inp[2]) ? node2884 : 8'b00011110;
													assign node2884 = (inp[6]) ? 8'b00011110 : 8'b00001110;
												assign node2887 = (inp[2]) ? 8'b00001110 : 8'b00001111;
										assign node2890 = (inp[5]) ? node2896 : node2891;
											assign node2891 = (inp[6]) ? node2893 : 8'b00101010;
												assign node2893 = (inp[2]) ? 8'b00101010 : 8'b00111010;
											assign node2896 = (inp[2]) ? node2898 : 8'b00111010;
												assign node2898 = (inp[3]) ? 8'b00011110 : 8'b00011111;
								assign node2901 = (inp[2]) ? node2929 : node2902;
									assign node2902 = (inp[1]) ? node2912 : node2903;
										assign node2903 = (inp[3]) ? node2909 : node2904;
											assign node2904 = (inp[6]) ? node2906 : 8'b00101110;
												assign node2906 = (inp[0]) ? 8'b00111110 : 8'b00101110;
											assign node2909 = (inp[12]) ? 8'b00101111 : 8'b00111110;
										assign node2912 = (inp[0]) ? node2922 : node2913;
											assign node2913 = (inp[6]) ? node2919 : node2914;
												assign node2914 = (inp[12]) ? 8'b00101110 : node2915;
													assign node2915 = (inp[5]) ? 8'b00111010 : 8'b00111011;
												assign node2919 = (inp[12]) ? 8'b00111110 : 8'b00101110;
											assign node2922 = (inp[3]) ? 8'b00111110 : node2923;
												assign node2923 = (inp[6]) ? node2925 : 8'b00111010;
													assign node2925 = (inp[5]) ? 8'b00111011 : 8'b00101011;
									assign node2929 = (inp[3]) ? node2941 : node2930;
										assign node2930 = (inp[1]) ? node2936 : node2931;
											assign node2931 = (inp[0]) ? 8'b00111011 : node2932;
												assign node2932 = (inp[5]) ? 8'b00101011 : 8'b00111011;
											assign node2936 = (inp[5]) ? node2938 : 8'b00111010;
												assign node2938 = (inp[6]) ? 8'b00111011 : 8'b00101110;
										assign node2941 = (inp[12]) ? 8'b00111010 : 8'b00111110;
							assign node2944 = (inp[0]) ? node3002 : node2945;
								assign node2945 = (inp[12]) ? node2977 : node2946;
									assign node2946 = (inp[6]) ? node2962 : node2947;
										assign node2947 = (inp[3]) ? node2953 : node2948;
											assign node2948 = (inp[5]) ? node2950 : 8'b00011111;
												assign node2950 = (inp[10]) ? 8'b00011011 : 8'b00011111;
											assign node2953 = (inp[1]) ? node2959 : node2954;
												assign node2954 = (inp[5]) ? node2956 : 8'b00111010;
													assign node2956 = (inp[10]) ? 8'b00011110 : 8'b00111010;
												assign node2959 = (inp[5]) ? 8'b00011010 : 8'b00011111;
										assign node2962 = (inp[2]) ? node2968 : node2963;
											assign node2963 = (inp[1]) ? 8'b00101010 : node2964;
												assign node2964 = (inp[5]) ? 8'b00001110 : 8'b00101011;
											assign node2968 = (inp[3]) ? node2974 : node2969;
												assign node2969 = (inp[5]) ? node2971 : 8'b00011111;
													assign node2971 = (inp[10]) ? 8'b00001011 : 8'b00001111;
												assign node2974 = (inp[1]) ? 8'b00001110 : 8'b00101010;
									assign node2977 = (inp[5]) ? node2987 : node2978;
										assign node2978 = (inp[3]) ? node2984 : node2979;
											assign node2979 = (inp[2]) ? 8'b00101010 : node2980;
												assign node2980 = (inp[1]) ? 8'b00101010 : 8'b00111010;
											assign node2984 = (inp[1]) ? 8'b00101010 : 8'b00101011;
										assign node2987 = (inp[6]) ? node2993 : node2988;
											assign node2988 = (inp[3]) ? node2990 : 8'b00101010;
												assign node2990 = (inp[10]) ? 8'b00001011 : 8'b00101011;
											assign node2993 = (inp[3]) ? node2997 : node2994;
												assign node2994 = (inp[10]) ? 8'b00011011 : 8'b00011111;
												assign node2997 = (inp[1]) ? node2999 : 8'b00111010;
													assign node2999 = (inp[2]) ? 8'b00011110 : 8'b00011111;
								assign node3002 = (inp[12]) ? node3038 : node3003;
									assign node3003 = (inp[10]) ? node3021 : node3004;
										assign node3004 = (inp[1]) ? node3008 : node3005;
											assign node3005 = (inp[2]) ? 8'b00001011 : 8'b00011011;
											assign node3008 = (inp[5]) ? node3018 : node3009;
												assign node3009 = (inp[3]) ? node3015 : node3010;
													assign node3010 = (inp[6]) ? 8'b00011010 : node3011;
														assign node3011 = (inp[2]) ? 8'b00001010 : 8'b00011010;
													assign node3015 = (inp[2]) ? 8'b00001011 : 8'b00001110;
												assign node3018 = (inp[6]) ? 8'b00001011 : 8'b00011010;
										assign node3021 = (inp[5]) ? node3027 : node3022;
											assign node3022 = (inp[3]) ? node3024 : 8'b00011110;
												assign node3024 = (inp[2]) ? 8'b00001111 : 8'b00011111;
											assign node3027 = (inp[2]) ? node3035 : node3028;
												assign node3028 = (inp[6]) ? node3032 : node3029;
													assign node3029 = (inp[1]) ? 8'b00011010 : 8'b00011110;
													assign node3032 = (inp[3]) ? 8'b00001111 : 8'b00001110;
												assign node3035 = (inp[1]) ? 8'b00001010 : 8'b00001011;
									assign node3038 = (inp[10]) ? node3046 : node3039;
										assign node3039 = (inp[1]) ? node3041 : 8'b00011110;
											assign node3041 = (inp[2]) ? 8'b00011010 : node3042;
												assign node3042 = (inp[3]) ? 8'b00011110 : 8'b00001011;
										assign node3046 = (inp[5]) ? node3054 : node3047;
											assign node3047 = (inp[2]) ? node3051 : node3048;
												assign node3048 = (inp[6]) ? 8'b00111010 : 8'b00101010;
												assign node3051 = (inp[6]) ? 8'b00001111 : 8'b00011110;
											assign node3054 = (inp[2]) ? node3058 : node3055;
												assign node3055 = (inp[6]) ? 8'b00011011 : 8'b00001011;
												assign node3058 = (inp[1]) ? 8'b00011010 : 8'b00011011;
				assign node3061 = (inp[0]) ? node3387 : node3062;
					assign node3062 = (inp[5]) ? node3182 : node3063;
						assign node3063 = (inp[12]) ? node3145 : node3064;
							assign node3064 = (inp[11]) ? node3108 : node3065;
								assign node3065 = (inp[10]) ? node3081 : node3066;
									assign node3066 = (inp[6]) ? node3072 : node3067;
										assign node3067 = (inp[3]) ? node3069 : 8'b10000010;
											assign node3069 = (inp[1]) ? 8'b10000010 : 8'b00001011;
										assign node3072 = (inp[2]) ? node3078 : node3073;
											assign node3073 = (inp[8]) ? 8'b00011010 : node3074;
												assign node3074 = (inp[9]) ? 8'b00011010 : 8'b00011011;
											assign node3078 = (inp[9]) ? 8'b10000010 : 8'b00001011;
									assign node3081 = (inp[8]) ? node3097 : node3082;
										assign node3082 = (inp[3]) ? node3088 : node3083;
											assign node3083 = (inp[2]) ? 8'b00001110 : node3084;
												assign node3084 = (inp[6]) ? 8'b00011110 : 8'b00001110;
											assign node3088 = (inp[1]) ? node3094 : node3089;
												assign node3089 = (inp[2]) ? 8'b00001111 : node3090;
													assign node3090 = (inp[6]) ? 8'b00011111 : 8'b00001111;
												assign node3094 = (inp[2]) ? 8'b00001110 : 8'b00011110;
										assign node3097 = (inp[3]) ? node3103 : node3098;
											assign node3098 = (inp[2]) ? 8'b10000010 : node3099;
												assign node3099 = (inp[9]) ? 8'b10000010 : 8'b00011010;
											assign node3103 = (inp[6]) ? node3105 : 8'b00001011;
												assign node3105 = (inp[1]) ? 8'b00011010 : 8'b00011011;
								assign node3108 = (inp[6]) ? node3122 : node3109;
									assign node3109 = (inp[10]) ? node3111 : 8'b11110111;
										assign node3111 = (inp[8]) ? node3117 : node3112;
											assign node3112 = (inp[9]) ? node3114 : 8'b00011011;
												assign node3114 = (inp[1]) ? 8'b00011011 : 8'b00011110;
											assign node3117 = (inp[1]) ? 8'b11110111 : node3118;
												assign node3118 = (inp[3]) ? 8'b00011010 : 8'b11110111;
									assign node3122 = (inp[2]) ? node3134 : node3123;
										assign node3123 = (inp[1]) ? node3129 : node3124;
											assign node3124 = (inp[3]) ? 8'b00001011 : node3125;
												assign node3125 = (inp[8]) ? 8'b00001010 : 8'b00001110;
											assign node3129 = (inp[10]) ? node3131 : 8'b00001010;
												assign node3131 = (inp[8]) ? 8'b00001010 : 8'b00001110;
										assign node3134 = (inp[8]) ? node3140 : node3135;
											assign node3135 = (inp[3]) ? 8'b00011010 : node3136;
												assign node3136 = (inp[10]) ? 8'b00011011 : 8'b11110111;
											assign node3140 = (inp[3]) ? node3142 : 8'b11110111;
												assign node3142 = (inp[1]) ? 8'b11110111 : 8'b00011010;
							assign node3145 = (inp[10]) ? node3163 : node3146;
								assign node3146 = (inp[3]) ? node3152 : node3147;
									assign node3147 = (inp[2]) ? 8'b00000010 : node3148;
										assign node3148 = (inp[6]) ? 8'b00011010 : 8'b00000010;
									assign node3152 = (inp[1]) ? node3158 : node3153;
										assign node3153 = (inp[2]) ? 8'b00001011 : node3154;
											assign node3154 = (inp[6]) ? 8'b00011011 : 8'b00001011;
										assign node3158 = (inp[6]) ? node3160 : 8'b00000010;
											assign node3160 = (inp[2]) ? 8'b00000010 : 8'b00011010;
								assign node3163 = (inp[8]) ? node3173 : node3164;
									assign node3164 = (inp[1]) ? node3168 : node3165;
										assign node3165 = (inp[3]) ? 8'b00001111 : 8'b00001110;
										assign node3168 = (inp[6]) ? node3170 : 8'b00001110;
											assign node3170 = (inp[2]) ? 8'b00001110 : 8'b00011110;
									assign node3173 = (inp[6]) ? node3179 : node3174;
										assign node3174 = (inp[1]) ? 8'b00000010 : node3175;
											assign node3175 = (inp[3]) ? 8'b00001011 : 8'b00000010;
										assign node3179 = (inp[2]) ? 8'b00000010 : 8'b00011010;
						assign node3182 = (inp[9]) ? node3298 : node3183;
							assign node3183 = (inp[8]) ? node3249 : node3184;
								assign node3184 = (inp[10]) ? node3226 : node3185;
									assign node3185 = (inp[1]) ? node3207 : node3186;
										assign node3186 = (inp[3]) ? node3202 : node3187;
											assign node3187 = (inp[11]) ? node3195 : node3188;
												assign node3188 = (inp[2]) ? node3192 : node3189;
													assign node3189 = (inp[6]) ? 8'b00011010 : 8'b00000010;
													assign node3192 = (inp[12]) ? 8'b10010000 : 8'b10000010;
												assign node3195 = (inp[12]) ? node3197 : 8'b11110111;
													assign node3197 = (inp[2]) ? node3199 : 8'b00011010;
														assign node3199 = (inp[6]) ? 8'b11110101 : 8'b00000010;
											assign node3202 = (inp[11]) ? 8'b00011010 : node3203;
												assign node3203 = (inp[6]) ? 8'b00011011 : 8'b00001011;
										assign node3207 = (inp[11]) ? node3217 : node3208;
											assign node3208 = (inp[3]) ? node3214 : node3209;
												assign node3209 = (inp[6]) ? 8'b10010000 : node3210;
													assign node3210 = (inp[12]) ? 8'b00000010 : 8'b10000010;
												assign node3214 = (inp[6]) ? 8'b10011001 : 8'b10000001;
											assign node3217 = (inp[3]) ? node3221 : node3218;
												assign node3218 = (inp[2]) ? 8'b11110101 : 8'b00001010;
												assign node3221 = (inp[6]) ? node3223 : 8'b10110100;
													assign node3223 = (inp[12]) ? 8'b10110100 : 8'b10100100;
									assign node3226 = (inp[11]) ? node3232 : node3227;
										assign node3227 = (inp[6]) ? 8'b00011110 : node3228;
											assign node3228 = (inp[3]) ? 8'b00001111 : 8'b00001110;
										assign node3232 = (inp[12]) ? node3242 : node3233;
											assign node3233 = (inp[6]) ? node3239 : node3234;
												assign node3234 = (inp[1]) ? node3236 : 8'b00011110;
													assign node3236 = (inp[3]) ? 8'b00011010 : 8'b00011011;
												assign node3239 = (inp[2]) ? 8'b00001011 : 8'b00001110;
											assign node3242 = (inp[6]) ? node3246 : node3243;
												assign node3243 = (inp[1]) ? 8'b00001011 : 8'b00001111;
												assign node3246 = (inp[3]) ? 8'b00011111 : 8'b00011011;
								assign node3249 = (inp[11]) ? node3273 : node3250;
									assign node3250 = (inp[10]) ? node3264 : node3251;
										assign node3251 = (inp[6]) ? node3259 : node3252;
											assign node3252 = (inp[1]) ? node3256 : node3253;
												assign node3253 = (inp[3]) ? 8'b00001011 : 8'b10000010;
												assign node3256 = (inp[3]) ? 8'b10000001 : 8'b10000010;
											assign node3259 = (inp[2]) ? 8'b10010000 : node3260;
												assign node3260 = (inp[3]) ? 8'b00011011 : 8'b00011010;
										assign node3264 = (inp[6]) ? node3268 : node3265;
											assign node3265 = (inp[3]) ? 8'b10000101 : 8'b10000100;
											assign node3268 = (inp[2]) ? 8'b10010100 : node3269;
												assign node3269 = (inp[3]) ? 8'b10011101 : 8'b10011100;
									assign node3273 = (inp[1]) ? node3289 : node3274;
										assign node3274 = (inp[3]) ? node3280 : node3275;
											assign node3275 = (inp[12]) ? 8'b10100100 : node3276;
												assign node3276 = (inp[10]) ? 8'b10110001 : 8'b10100101;
											assign node3280 = (inp[10]) ? node3282 : 8'b00001010;
												assign node3282 = (inp[6]) ? node3286 : node3283;
													assign node3283 = (inp[12]) ? 8'b10101101 : 8'b10111100;
													assign node3286 = (inp[12]) ? 8'b11111101 : 8'b10101101;
										assign node3289 = (inp[10]) ? node3293 : node3290;
											assign node3290 = (inp[6]) ? 8'b10100100 : 8'b10100101;
											assign node3293 = (inp[12]) ? 8'b10100001 : node3294;
												assign node3294 = (inp[3]) ? 8'b10110000 : 8'b10110001;
							assign node3298 = (inp[6]) ? node3342 : node3299;
								assign node3299 = (inp[8]) ? node3319 : node3300;
									assign node3300 = (inp[10]) ? node3310 : node3301;
										assign node3301 = (inp[11]) ? node3305 : node3302;
											assign node3302 = (inp[3]) ? 8'b10101001 : 8'b10100000;
											assign node3305 = (inp[12]) ? node3307 : 8'b10010101;
												assign node3307 = (inp[2]) ? 8'b10000101 : 8'b10100000;
										assign node3310 = (inp[3]) ? node3314 : node3311;
											assign node3311 = (inp[11]) ? 8'b10111001 : 8'b10101100;
											assign node3314 = (inp[11]) ? node3316 : 8'b10101101;
												assign node3316 = (inp[1]) ? 8'b10101001 : 8'b10101101;
									assign node3319 = (inp[11]) ? node3327 : node3320;
										assign node3320 = (inp[3]) ? node3324 : node3321;
											assign node3321 = (inp[10]) ? 8'b10100100 : 8'b10100000;
											assign node3324 = (inp[12]) ? 8'b10100101 : 8'b10100001;
										assign node3327 = (inp[12]) ? node3335 : node3328;
											assign node3328 = (inp[3]) ? node3332 : node3329;
												assign node3329 = (inp[10]) ? 8'b10010001 : 8'b10010101;
												assign node3332 = (inp[1]) ? 8'b10010000 : 8'b10011100;
											assign node3335 = (inp[3]) ? node3339 : node3336;
												assign node3336 = (inp[10]) ? 8'b10000100 : 8'b10100000;
												assign node3339 = (inp[10]) ? 8'b10000001 : 8'b10101001;
								assign node3342 = (inp[10]) ? node3366 : node3343;
									assign node3343 = (inp[11]) ? node3353 : node3344;
										assign node3344 = (inp[3]) ? node3348 : node3345;
											assign node3345 = (inp[2]) ? 8'b10110000 : 8'b10111000;
											assign node3348 = (inp[1]) ? node3350 : 8'b10111001;
												assign node3350 = (inp[2]) ? 8'b10110001 : 8'b10111001;
										assign node3353 = (inp[1]) ? node3357 : node3354;
											assign node3354 = (inp[12]) ? 8'b10111000 : 8'b10101000;
											assign node3357 = (inp[12]) ? node3361 : node3358;
												assign node3358 = (inp[3]) ? 8'b10000100 : 8'b10101000;
												assign node3361 = (inp[2]) ? node3363 : 8'b10011101;
													assign node3363 = (inp[3]) ? 8'b10010100 : 8'b10010101;
									assign node3366 = (inp[3]) ? node3378 : node3367;
										assign node3367 = (inp[1]) ? node3373 : node3368;
											assign node3368 = (inp[11]) ? node3370 : 8'b10111100;
												assign node3370 = (inp[2]) ? 8'b10101001 : 8'b10101100;
											assign node3373 = (inp[8]) ? node3375 : 8'b10111100;
												assign node3375 = (inp[2]) ? 8'b10110100 : 8'b10111100;
										assign node3378 = (inp[11]) ? node3380 : 8'b11111101;
											assign node3380 = (inp[1]) ? node3384 : node3381;
												assign node3381 = (inp[2]) ? 8'b10101100 : 8'b11111101;
												assign node3384 = (inp[2]) ? 8'b10010000 : 8'b10011001;
					assign node3387 = (inp[5]) ? node3665 : node3388;
						assign node3388 = (inp[9]) ? node3528 : node3389;
							assign node3389 = (inp[10]) ? node3455 : node3390;
								assign node3390 = (inp[11]) ? node3424 : node3391;
									assign node3391 = (inp[8]) ? node3407 : node3392;
										assign node3392 = (inp[3]) ? node3400 : node3393;
											assign node3393 = (inp[1]) ? node3397 : node3394;
												assign node3394 = (inp[6]) ? 8'b10100000 : 8'b10110000;
												assign node3397 = (inp[2]) ? 8'b10110001 : 8'b10100001;
											assign node3400 = (inp[1]) ? node3404 : node3401;
												assign node3401 = (inp[6]) ? 8'b10101001 : 8'b10111001;
												assign node3404 = (inp[6]) ? 8'b10111000 : 8'b10110000;
										assign node3407 = (inp[2]) ? node3413 : node3408;
											assign node3408 = (inp[6]) ? node3410 : 8'b10100100;
												assign node3410 = (inp[3]) ? 8'b11111101 : 8'b10111100;
											assign node3413 = (inp[6]) ? node3421 : node3414;
												assign node3414 = (inp[12]) ? 8'b11110101 : node3415;
													assign node3415 = (inp[1]) ? node3417 : 8'b10110100;
														assign node3417 = (inp[3]) ? 8'b10110100 : 8'b11110101;
												assign node3421 = (inp[1]) ? 8'b10100101 : 8'b10100100;
									assign node3424 = (inp[6]) ? node3440 : node3425;
										assign node3425 = (inp[8]) ? node3431 : node3426;
											assign node3426 = (inp[2]) ? node3428 : 8'b10111000;
												assign node3428 = (inp[12]) ? 8'b10010101 : 8'b10000101;
											assign node3431 = (inp[2]) ? node3435 : node3432;
												assign node3432 = (inp[1]) ? 8'b10000001 : 8'b10000100;
												assign node3435 = (inp[12]) ? node3437 : 8'b10000001;
													assign node3437 = (inp[1]) ? 8'b10010000 : 8'b10010001;
										assign node3440 = (inp[2]) ? node3448 : node3441;
											assign node3441 = (inp[12]) ? node3445 : node3442;
												assign node3442 = (inp[3]) ? 8'b10001101 : 8'b10101000;
												assign node3445 = (inp[8]) ? 8'b10011001 : 8'b10011101;
											assign node3448 = (inp[12]) ? node3452 : node3449;
												assign node3449 = (inp[3]) ? 8'b10111000 : 8'b10010100;
												assign node3452 = (inp[8]) ? 8'b10000100 : 8'b10100000;
								assign node3455 = (inp[8]) ? node3493 : node3456;
									assign node3456 = (inp[11]) ? node3468 : node3457;
										assign node3457 = (inp[2]) ? node3465 : node3458;
											assign node3458 = (inp[6]) ? 8'b10111100 : node3459;
												assign node3459 = (inp[3]) ? node3461 : 8'b10101101;
													assign node3461 = (inp[1]) ? 8'b10101100 : 8'b10101101;
											assign node3465 = (inp[3]) ? 8'b11111101 : 8'b10101100;
										assign node3468 = (inp[3]) ? node3480 : node3469;
											assign node3469 = (inp[12]) ? node3475 : node3470;
												assign node3470 = (inp[1]) ? 8'b10111000 : node3471;
													assign node3471 = (inp[2]) ? 8'b10101001 : 8'b10111001;
												assign node3475 = (inp[2]) ? 8'b10111001 : node3476;
													assign node3476 = (inp[6]) ? 8'b10111001 : 8'b10101001;
											assign node3480 = (inp[12]) ? node3488 : node3481;
												assign node3481 = (inp[2]) ? 8'b10111001 : node3482;
													assign node3482 = (inp[6]) ? 8'b10101100 : node3483;
														assign node3483 = (inp[1]) ? 8'b10111001 : 8'b10111100;
												assign node3488 = (inp[6]) ? node3490 : 8'b10101100;
													assign node3490 = (inp[2]) ? 8'b10101101 : 8'b11111101;
									assign node3493 = (inp[12]) ? node3509 : node3494;
										assign node3494 = (inp[11]) ? node3502 : node3495;
											assign node3495 = (inp[6]) ? node3499 : node3496;
												assign node3496 = (inp[3]) ? 8'b10110000 : 8'b10110001;
												assign node3499 = (inp[1]) ? 8'b10111001 : 8'b10111000;
											assign node3502 = (inp[1]) ? node3506 : node3503;
												assign node3503 = (inp[3]) ? 8'b10111000 : 8'b10010101;
												assign node3506 = (inp[6]) ? 8'b10010101 : 8'b10010100;
										assign node3509 = (inp[3]) ? node3517 : node3510;
											assign node3510 = (inp[2]) ? node3514 : node3511;
												assign node3511 = (inp[1]) ? 8'b10100001 : 8'b10100000;
												assign node3514 = (inp[1]) ? 8'b10100001 : 8'b10010101;
											assign node3517 = (inp[1]) ? node3523 : node3518;
												assign node3518 = (inp[11]) ? 8'b10101001 : node3519;
													assign node3519 = (inp[6]) ? 8'b10111001 : 8'b10101001;
												assign node3523 = (inp[2]) ? node3525 : 8'b10111000;
													assign node3525 = (inp[6]) ? 8'b10100000 : 8'b10110000;
							assign node3528 = (inp[8]) ? node3602 : node3529;
								assign node3529 = (inp[10]) ? node3569 : node3530;
									assign node3530 = (inp[1]) ? node3552 : node3531;
										assign node3531 = (inp[3]) ? node3545 : node3532;
											assign node3532 = (inp[2]) ? node3540 : node3533;
												assign node3533 = (inp[6]) ? node3537 : node3534;
													assign node3534 = (inp[12]) ? 8'b00000010 : 8'b10000010;
													assign node3537 = (inp[11]) ? 8'b00001010 : 8'b00011010;
												assign node3540 = (inp[11]) ? 8'b11110111 : node3541;
													assign node3541 = (inp[12]) ? 8'b10010000 : 8'b10000010;
											assign node3545 = (inp[11]) ? node3547 : 8'b00011011;
												assign node3547 = (inp[2]) ? node3549 : 8'b00001011;
													assign node3549 = (inp[12]) ? 8'b00011010 : 8'b00001010;
										assign node3552 = (inp[3]) ? node3560 : node3553;
											assign node3553 = (inp[11]) ? 8'b10100101 : node3554;
												assign node3554 = (inp[6]) ? 8'b10000001 : node3555;
													assign node3555 = (inp[2]) ? 8'b10010001 : 8'b10000001;
											assign node3560 = (inp[2]) ? node3566 : node3561;
												assign node3561 = (inp[6]) ? 8'b00011010 : node3562;
													assign node3562 = (inp[11]) ? 8'b00000010 : 8'b10000010;
												assign node3566 = (inp[6]) ? 8'b11110111 : 8'b10010000;
									assign node3569 = (inp[1]) ? node3583 : node3570;
										assign node3570 = (inp[3]) ? node3578 : node3571;
											assign node3571 = (inp[2]) ? node3575 : node3572;
												assign node3572 = (inp[6]) ? 8'b00011110 : 8'b00001110;
												assign node3575 = (inp[6]) ? 8'b00001110 : 8'b00011110;
											assign node3578 = (inp[12]) ? node3580 : 8'b00011110;
												assign node3580 = (inp[6]) ? 8'b00011111 : 8'b00001111;
										assign node3583 = (inp[3]) ? node3595 : node3584;
											assign node3584 = (inp[11]) ? node3588 : node3585;
												assign node3585 = (inp[6]) ? 8'b00011111 : 8'b00001111;
												assign node3588 = (inp[12]) ? node3590 : 8'b00001011;
													assign node3590 = (inp[6]) ? node3592 : 8'b00001011;
														assign node3592 = (inp[2]) ? 8'b00001011 : 8'b00011011;
											assign node3595 = (inp[11]) ? 8'b00001110 : node3596;
												assign node3596 = (inp[2]) ? 8'b00011110 : node3597;
													assign node3597 = (inp[6]) ? 8'b00011110 : 8'b00001110;
								assign node3602 = (inp[11]) ? node3634 : node3603;
									assign node3603 = (inp[10]) ? node3621 : node3604;
										assign node3604 = (inp[6]) ? node3612 : node3605;
											assign node3605 = (inp[2]) ? node3607 : 8'b10000100;
												assign node3607 = (inp[3]) ? 8'b10010100 : node3608;
													assign node3608 = (inp[1]) ? 8'b10010101 : 8'b10010100;
											assign node3612 = (inp[2]) ? node3618 : node3613;
												assign node3613 = (inp[3]) ? node3615 : 8'b10011101;
													assign node3615 = (inp[1]) ? 8'b10011100 : 8'b10011101;
												assign node3618 = (inp[12]) ? 8'b10001101 : 8'b10000100;
										assign node3621 = (inp[3]) ? node3629 : node3622;
											assign node3622 = (inp[1]) ? node3624 : 8'b10000010;
												assign node3624 = (inp[6]) ? 8'b10011001 : node3625;
													assign node3625 = (inp[2]) ? 8'b10010001 : 8'b10000001;
											assign node3629 = (inp[6]) ? node3631 : 8'b00011011;
												assign node3631 = (inp[12]) ? 8'b00000010 : 8'b10000010;
									assign node3634 = (inp[6]) ? node3648 : node3635;
										assign node3635 = (inp[10]) ? node3645 : node3636;
											assign node3636 = (inp[3]) ? node3640 : node3637;
												assign node3637 = (inp[1]) ? 8'b10110000 : 8'b10110001;
												assign node3640 = (inp[2]) ? node3642 : 8'b10100100;
													assign node3642 = (inp[12]) ? 8'b10110001 : 8'b10100001;
											assign node3645 = (inp[1]) ? 8'b10100100 : 8'b10100101;
										assign node3648 = (inp[2]) ? node3660 : node3649;
											assign node3649 = (inp[12]) ? node3653 : node3650;
												assign node3650 = (inp[3]) ? 8'b00001010 : 8'b10101101;
												assign node3653 = (inp[10]) ? 8'b11111101 : node3654;
													assign node3654 = (inp[3]) ? 8'b11111101 : node3655;
														assign node3655 = (inp[1]) ? 8'b10111001 : 8'b10111100;
											assign node3660 = (inp[10]) ? 8'b00000010 : node3661;
												assign node3661 = (inp[12]) ? 8'b10100100 : 8'b10111100;
						assign node3665 = (inp[11]) ? node3741 : node3666;
							assign node3666 = (inp[3]) ? node3702 : node3667;
								assign node3667 = (inp[1]) ? node3683 : node3668;
									assign node3668 = (inp[8]) ? node3678 : node3669;
										assign node3669 = (inp[10]) ? node3675 : node3670;
											assign node3670 = (inp[2]) ? 8'b10110000 : node3671;
												assign node3671 = (inp[6]) ? 8'b10111000 : 8'b10100000;
											assign node3675 = (inp[2]) ? 8'b10111100 : 8'b10101100;
										assign node3678 = (inp[2]) ? 8'b10110100 : node3679;
											assign node3679 = (inp[6]) ? 8'b10111100 : 8'b10100100;
									assign node3683 = (inp[6]) ? node3695 : node3684;
										assign node3684 = (inp[2]) ? node3690 : node3685;
											assign node3685 = (inp[8]) ? 8'b10100101 : node3686;
												assign node3686 = (inp[10]) ? 8'b10101101 : 8'b10100001;
											assign node3690 = (inp[10]) ? node3692 : 8'b10110001;
												assign node3692 = (inp[12]) ? 8'b11111101 : 8'b11110101;
										assign node3695 = (inp[2]) ? 8'b11110101 : node3696;
											assign node3696 = (inp[8]) ? 8'b11111101 : node3697;
												assign node3697 = (inp[12]) ? 8'b11111101 : 8'b10111001;
								assign node3702 = (inp[6]) ? node3728 : node3703;
									assign node3703 = (inp[2]) ? node3715 : node3704;
										assign node3704 = (inp[10]) ? node3710 : node3705;
											assign node3705 = (inp[1]) ? node3707 : 8'b10101001;
												assign node3707 = (inp[8]) ? 8'b10100101 : 8'b10100001;
											assign node3710 = (inp[8]) ? node3712 : 8'b10101101;
												assign node3712 = (inp[1]) ? 8'b10100101 : 8'b10101101;
										assign node3715 = (inp[10]) ? node3723 : node3716;
											assign node3716 = (inp[8]) ? node3720 : node3717;
												assign node3717 = (inp[9]) ? 8'b10110001 : 8'b10111001;
												assign node3720 = (inp[1]) ? 8'b11110101 : 8'b11111101;
											assign node3723 = (inp[8]) ? node3725 : 8'b11111101;
												assign node3725 = (inp[1]) ? 8'b11110101 : 8'b11111101;
									assign node3728 = (inp[8]) ? node3736 : node3729;
										assign node3729 = (inp[10]) ? 8'b11111101 : node3730;
											assign node3730 = (inp[1]) ? node3732 : 8'b10111001;
												assign node3732 = (inp[12]) ? 8'b10111001 : 8'b10110001;
										assign node3736 = (inp[2]) ? node3738 : 8'b11111101;
											assign node3738 = (inp[1]) ? 8'b11110101 : 8'b11111101;
							assign node3741 = (inp[8]) ? node3789 : node3742;
								assign node3742 = (inp[10]) ? node3764 : node3743;
									assign node3743 = (inp[1]) ? node3757 : node3744;
										assign node3744 = (inp[3]) ? node3754 : node3745;
											assign node3745 = (inp[2]) ? node3751 : node3746;
												assign node3746 = (inp[12]) ? node3748 : 8'b10010101;
													assign node3748 = (inp[9]) ? 8'b10111000 : 8'b10100000;
												assign node3751 = (inp[6]) ? 8'b10000101 : 8'b10010101;
											assign node3754 = (inp[12]) ? 8'b10111000 : 8'b10101000;
										assign node3757 = (inp[2]) ? node3761 : node3758;
											assign node3758 = (inp[12]) ? 8'b10011101 : 8'b10010100;
											assign node3761 = (inp[12]) ? 8'b10010100 : 8'b10000100;
									assign node3764 = (inp[1]) ? node3780 : node3765;
										assign node3765 = (inp[12]) ? node3773 : node3766;
											assign node3766 = (inp[2]) ? node3770 : node3767;
												assign node3767 = (inp[3]) ? 8'b10111100 : 8'b10101100;
												assign node3770 = (inp[3]) ? 8'b10101100 : 8'b10101001;
											assign node3773 = (inp[6]) ? 8'b11111101 : node3774;
												assign node3774 = (inp[2]) ? node3776 : 8'b10101100;
													assign node3776 = (inp[3]) ? 8'b10111100 : 8'b10111001;
										assign node3780 = (inp[2]) ? 8'b10111000 : node3781;
											assign node3781 = (inp[9]) ? 8'b10111000 : node3782;
												assign node3782 = (inp[12]) ? node3784 : 8'b10101001;
													assign node3784 = (inp[6]) ? 8'b10111001 : 8'b10101001;
								assign node3789 = (inp[1]) ? node3811 : node3790;
									assign node3790 = (inp[3]) ? node3802 : node3791;
										assign node3791 = (inp[2]) ? node3799 : node3792;
											assign node3792 = (inp[6]) ? node3796 : node3793;
												assign node3793 = (inp[12]) ? 8'b10000100 : 8'b10010001;
												assign node3796 = (inp[12]) ? 8'b10011100 : 8'b10001100;
											assign node3799 = (inp[12]) ? 8'b10010001 : 8'b10000001;
										assign node3802 = (inp[12]) ? node3808 : node3803;
											assign node3803 = (inp[2]) ? 8'b10001100 : node3804;
												assign node3804 = (inp[6]) ? 8'b10001101 : 8'b10011100;
											assign node3808 = (inp[2]) ? 8'b10011100 : 8'b10011101;
									assign node3811 = (inp[2]) ? node3819 : node3812;
										assign node3812 = (inp[6]) ? node3816 : node3813;
											assign node3813 = (inp[12]) ? 8'b10000001 : 8'b10010000;
											assign node3816 = (inp[12]) ? 8'b10011001 : 8'b10001001;
										assign node3819 = (inp[12]) ? 8'b10010000 : 8'b10000000;
			assign node3822 = (inp[12]) ? node4242 : node3823;
				assign node3823 = (inp[11]) ? node4041 : node3824;
					assign node3824 = (inp[0]) ? node3902 : node3825;
						assign node3825 = (inp[5]) ? node3827 : 8'b10000010;
							assign node3827 = (inp[6]) ? node3855 : node3828;
								assign node3828 = (inp[8]) ? node3838 : node3829;
									assign node3829 = (inp[9]) ? node3835 : node3830;
										assign node3830 = (inp[1]) ? node3832 : 8'b10000010;
											assign node3832 = (inp[3]) ? 8'b10000001 : 8'b10000010;
										assign node3835 = (inp[13]) ? 8'b10100000 : 8'b10000010;
									assign node3838 = (inp[10]) ? node3846 : node3839;
										assign node3839 = (inp[9]) ? 8'b10100000 : node3840;
											assign node3840 = (inp[3]) ? node3842 : 8'b10000010;
												assign node3842 = (inp[1]) ? 8'b10000001 : 8'b10000010;
										assign node3846 = (inp[13]) ? node3852 : node3847;
											assign node3847 = (inp[3]) ? node3849 : 8'b10000100;
												assign node3849 = (inp[1]) ? 8'b10000101 : 8'b10000100;
											assign node3852 = (inp[9]) ? 8'b10100100 : 8'b10000100;
								assign node3855 = (inp[2]) ? node3879 : node3856;
									assign node3856 = (inp[10]) ? node3866 : node3857;
										assign node3857 = (inp[3]) ? node3861 : node3858;
											assign node3858 = (inp[1]) ? 8'b10000010 : 8'b10100000;
											assign node3861 = (inp[13]) ? node3863 : 8'b10000001;
												assign node3863 = (inp[9]) ? 8'b10100001 : 8'b10000001;
										assign node3866 = (inp[8]) ? node3870 : node3867;
											assign node3867 = (inp[9]) ? 8'b10000001 : 8'b10000010;
											assign node3870 = (inp[9]) ? node3876 : node3871;
												assign node3871 = (inp[13]) ? node3873 : 8'b10000100;
													assign node3873 = (inp[3]) ? 8'b10000101 : 8'b10000100;
												assign node3876 = (inp[13]) ? 8'b10100100 : 8'b10000101;
									assign node3879 = (inp[9]) ? node3887 : node3880;
										assign node3880 = (inp[8]) ? node3884 : node3881;
											assign node3881 = (inp[3]) ? 8'b10010001 : 8'b10010000;
											assign node3884 = (inp[10]) ? 8'b10010100 : 8'b10010001;
										assign node3887 = (inp[13]) ? node3893 : node3888;
											assign node3888 = (inp[3]) ? node3890 : 8'b10010000;
												assign node3890 = (inp[1]) ? 8'b10010001 : 8'b10010000;
											assign node3893 = (inp[3]) ? node3899 : node3894;
												assign node3894 = (inp[8]) ? node3896 : 8'b10110000;
													assign node3896 = (inp[10]) ? 8'b10110100 : 8'b10110000;
												assign node3899 = (inp[1]) ? 8'b10110001 : 8'b10110000;
						assign node3902 = (inp[8]) ? node3954 : node3903;
							assign node3903 = (inp[1]) ? node3923 : node3904;
								assign node3904 = (inp[13]) ? node3912 : node3905;
									assign node3905 = (inp[2]) ? node3907 : 8'b10000010;
										assign node3907 = (inp[5]) ? 8'b10010000 : node3908;
											assign node3908 = (inp[6]) ? 8'b10000010 : 8'b10010000;
									assign node3912 = (inp[2]) ? node3918 : node3913;
										assign node3913 = (inp[9]) ? node3915 : 8'b10100000;
											assign node3915 = (inp[5]) ? 8'b10100000 : 8'b10000010;
										assign node3918 = (inp[5]) ? 8'b10110000 : node3919;
											assign node3919 = (inp[3]) ? 8'b10110000 : 8'b10010000;
								assign node3923 = (inp[5]) ? node3947 : node3924;
									assign node3924 = (inp[3]) ? node3938 : node3925;
										assign node3925 = (inp[13]) ? node3931 : node3926;
											assign node3926 = (inp[6]) ? 8'b10000001 : node3927;
												assign node3927 = (inp[2]) ? 8'b10010001 : 8'b10000001;
											assign node3931 = (inp[9]) ? node3935 : node3932;
												assign node3932 = (inp[2]) ? 8'b10110001 : 8'b10100001;
												assign node3935 = (inp[2]) ? 8'b10010001 : 8'b10000001;
										assign node3938 = (inp[6]) ? node3942 : node3939;
											assign node3939 = (inp[2]) ? 8'b10010000 : 8'b10000010;
											assign node3942 = (inp[9]) ? 8'b10000010 : node3943;
												assign node3943 = (inp[2]) ? 8'b10000010 : 8'b10100000;
									assign node3947 = (inp[13]) ? node3951 : node3948;
										assign node3948 = (inp[2]) ? 8'b10010001 : 8'b10000001;
										assign node3951 = (inp[2]) ? 8'b10110001 : 8'b10100001;
							assign node3954 = (inp[13]) ? node3988 : node3955;
								assign node3955 = (inp[2]) ? node3971 : node3956;
									assign node3956 = (inp[1]) ? node3962 : node3957;
										assign node3957 = (inp[5]) ? 8'b10000100 : node3958;
											assign node3958 = (inp[10]) ? 8'b10000010 : 8'b10000100;
										assign node3962 = (inp[5]) ? 8'b10000101 : node3963;
											assign node3963 = (inp[10]) ? node3967 : node3964;
												assign node3964 = (inp[9]) ? 8'b10000100 : 8'b10000101;
												assign node3967 = (inp[3]) ? 8'b10000010 : 8'b10000001;
									assign node3971 = (inp[1]) ? node3977 : node3972;
										assign node3972 = (inp[5]) ? 8'b10010100 : node3973;
											assign node3973 = (inp[6]) ? 8'b10000100 : 8'b10010100;
										assign node3977 = (inp[5]) ? 8'b10010101 : node3978;
											assign node3978 = (inp[3]) ? node3984 : node3979;
												assign node3979 = (inp[10]) ? 8'b10010001 : node3980;
													assign node3980 = (inp[9]) ? 8'b10000101 : 8'b10010101;
												assign node3984 = (inp[6]) ? 8'b10000100 : 8'b10010100;
								assign node3988 = (inp[2]) ? node4012 : node3989;
									assign node3989 = (inp[1]) ? node3999 : node3990;
										assign node3990 = (inp[10]) ? node3996 : node3991;
											assign node3991 = (inp[5]) ? 8'b10100100 : node3992;
												assign node3992 = (inp[9]) ? 8'b10000100 : 8'b10100100;
											assign node3996 = (inp[5]) ? 8'b10100100 : 8'b10100000;
										assign node3999 = (inp[5]) ? 8'b10100101 : node4000;
											assign node4000 = (inp[9]) ? node4008 : node4001;
												assign node4001 = (inp[3]) ? node4005 : node4002;
													assign node4002 = (inp[10]) ? 8'b10100001 : 8'b10100101;
													assign node4005 = (inp[10]) ? 8'b10100000 : 8'b10100100;
												assign node4008 = (inp[10]) ? 8'b10000010 : 8'b10000100;
									assign node4012 = (inp[5]) ? node4038 : node4013;
										assign node4013 = (inp[6]) ? node4025 : node4014;
											assign node4014 = (inp[10]) ? node4020 : node4015;
												assign node4015 = (inp[9]) ? node4017 : 8'b10110100;
													assign node4017 = (inp[3]) ? 8'b10010100 : 8'b10010101;
												assign node4020 = (inp[9]) ? 8'b10010000 : node4021;
													assign node4021 = (inp[1]) ? 8'b10110001 : 8'b10110000;
											assign node4025 = (inp[9]) ? node4031 : node4026;
												assign node4026 = (inp[10]) ? node4028 : 8'b10100100;
													assign node4028 = (inp[3]) ? 8'b10100000 : 8'b10100001;
												assign node4031 = (inp[3]) ? node4035 : node4032;
													assign node4032 = (inp[10]) ? 8'b10000001 : 8'b10000101;
													assign node4035 = (inp[10]) ? 8'b10000010 : 8'b10000100;
										assign node4038 = (inp[1]) ? 8'b11110101 : 8'b10110100;
					assign node4041 = (inp[0]) ? node4111 : node4042;
						assign node4042 = (inp[5]) ? node4044 : 8'b11110111;
							assign node4044 = (inp[6]) ? node4072 : node4045;
								assign node4045 = (inp[1]) ? node4059 : node4046;
									assign node4046 = (inp[13]) ? node4052 : node4047;
										assign node4047 = (inp[10]) ? node4049 : 8'b11110111;
											assign node4049 = (inp[3]) ? 8'b11110111 : 8'b10110001;
										assign node4052 = (inp[9]) ? 8'b10010101 : node4053;
											assign node4053 = (inp[8]) ? node4055 : 8'b11110111;
												assign node4055 = (inp[10]) ? 8'b10110001 : 8'b11110111;
									assign node4059 = (inp[3]) ? node4063 : node4060;
										assign node4060 = (inp[8]) ? 8'b10110001 : 8'b11110111;
										assign node4063 = (inp[9]) ? node4069 : node4064;
											assign node4064 = (inp[10]) ? node4066 : 8'b10110100;
												assign node4066 = (inp[8]) ? 8'b10110000 : 8'b10110100;
											assign node4069 = (inp[13]) ? 8'b10010100 : 8'b10110100;
								assign node4072 = (inp[2]) ? node4094 : node4073;
									assign node4073 = (inp[9]) ? node4083 : node4074;
										assign node4074 = (inp[3]) ? node4078 : node4075;
											assign node4075 = (inp[8]) ? 8'b10110001 : 8'b11110111;
											assign node4078 = (inp[1]) ? 8'b10110100 : node4079;
												assign node4079 = (inp[10]) ? 8'b10110001 : 8'b11110111;
										assign node4083 = (inp[13]) ? node4087 : node4084;
											assign node4084 = (inp[1]) ? 8'b10110100 : 8'b11110111;
											assign node4087 = (inp[10]) ? node4089 : 8'b10010101;
												assign node4089 = (inp[3]) ? 8'b10010000 : node4090;
													assign node4090 = (inp[8]) ? 8'b10010001 : 8'b10010101;
									assign node4094 = (inp[3]) ? node4100 : node4095;
										assign node4095 = (inp[8]) ? node4097 : 8'b10100101;
											assign node4097 = (inp[10]) ? 8'b10100001 : 8'b10100101;
										assign node4100 = (inp[1]) ? node4106 : node4101;
											assign node4101 = (inp[9]) ? node4103 : 8'b10100101;
												assign node4103 = (inp[13]) ? 8'b10000101 : 8'b10100101;
											assign node4106 = (inp[9]) ? node4108 : 8'b10100100;
												assign node4108 = (inp[13]) ? 8'b10000100 : 8'b10100100;
						assign node4111 = (inp[2]) ? node4167 : node4112;
							assign node4112 = (inp[13]) ? node4134 : node4113;
								assign node4113 = (inp[8]) ? node4121 : node4114;
									assign node4114 = (inp[1]) ? node4116 : 8'b11110111;
										assign node4116 = (inp[3]) ? node4118 : 8'b10110100;
											assign node4118 = (inp[5]) ? 8'b10110100 : 8'b11110111;
									assign node4121 = (inp[10]) ? node4125 : node4122;
										assign node4122 = (inp[1]) ? 8'b10110000 : 8'b10110001;
										assign node4125 = (inp[3]) ? node4129 : node4126;
											assign node4126 = (inp[5]) ? 8'b10110000 : 8'b10110100;
											assign node4129 = (inp[5]) ? node4131 : 8'b11110111;
												assign node4131 = (inp[6]) ? 8'b10110001 : 8'b10110000;
								assign node4134 = (inp[8]) ? node4150 : node4135;
									assign node4135 = (inp[5]) ? node4147 : node4136;
										assign node4136 = (inp[9]) ? node4142 : node4137;
											assign node4137 = (inp[3]) ? 8'b10010101 : node4138;
												assign node4138 = (inp[6]) ? 8'b10010100 : 8'b10010101;
											assign node4142 = (inp[1]) ? node4144 : 8'b11110111;
												assign node4144 = (inp[3]) ? 8'b11110111 : 8'b10110100;
										assign node4147 = (inp[1]) ? 8'b10010100 : 8'b10010101;
									assign node4150 = (inp[1]) ? node4158 : node4151;
										assign node4151 = (inp[9]) ? 8'b10110001 : node4152;
											assign node4152 = (inp[5]) ? 8'b10010001 : node4153;
												assign node4153 = (inp[10]) ? 8'b10010101 : 8'b10010001;
										assign node4158 = (inp[3]) ? node4164 : node4159;
											assign node4159 = (inp[6]) ? 8'b10010000 : node4160;
												assign node4160 = (inp[5]) ? 8'b10010000 : 8'b10010100;
											assign node4164 = (inp[5]) ? 8'b10010000 : 8'b10110001;
							assign node4167 = (inp[1]) ? node4203 : node4168;
								assign node4168 = (inp[8]) ? node4184 : node4169;
									assign node4169 = (inp[6]) ? node4177 : node4170;
										assign node4170 = (inp[13]) ? node4172 : 8'b10100101;
											assign node4172 = (inp[9]) ? node4174 : 8'b10000101;
												assign node4174 = (inp[3]) ? 8'b10000101 : 8'b10100101;
										assign node4177 = (inp[5]) ? node4181 : node4178;
											assign node4178 = (inp[9]) ? 8'b11110111 : 8'b10010101;
											assign node4181 = (inp[13]) ? 8'b10000101 : 8'b10100101;
									assign node4184 = (inp[13]) ? node4194 : node4185;
										assign node4185 = (inp[9]) ? node4191 : node4186;
											assign node4186 = (inp[6]) ? node4188 : 8'b10100001;
												assign node4188 = (inp[5]) ? 8'b10100001 : 8'b10110001;
											assign node4191 = (inp[10]) ? 8'b10100101 : 8'b10100001;
										assign node4194 = (inp[5]) ? 8'b10000001 : node4195;
											assign node4195 = (inp[9]) ? node4199 : node4196;
												assign node4196 = (inp[6]) ? 8'b10010001 : 8'b10000001;
												assign node4199 = (inp[10]) ? 8'b10100101 : 8'b10110001;
								assign node4203 = (inp[13]) ? node4225 : node4204;
									assign node4204 = (inp[5]) ? node4222 : node4205;
										assign node4205 = (inp[3]) ? node4217 : node4206;
											assign node4206 = (inp[6]) ? node4212 : node4207;
												assign node4207 = (inp[10]) ? 8'b10100100 : node4208;
													assign node4208 = (inp[8]) ? 8'b10100000 : 8'b10100100;
												assign node4212 = (inp[8]) ? node4214 : 8'b10110100;
													assign node4214 = (inp[9]) ? 8'b10110000 : 8'b10110100;
											assign node4217 = (inp[6]) ? node4219 : 8'b10100101;
												assign node4219 = (inp[8]) ? 8'b10110001 : 8'b11110111;
										assign node4222 = (inp[8]) ? 8'b10100000 : 8'b10100100;
									assign node4225 = (inp[5]) ? node4239 : node4226;
										assign node4226 = (inp[3]) ? node4236 : node4227;
											assign node4227 = (inp[9]) ? node4233 : node4228;
												assign node4228 = (inp[8]) ? node4230 : 8'b10010100;
													assign node4230 = (inp[10]) ? 8'b10000100 : 8'b10000000;
												assign node4233 = (inp[6]) ? 8'b10110100 : 8'b10100100;
											assign node4236 = (inp[9]) ? 8'b10100101 : 8'b10000101;
										assign node4239 = (inp[8]) ? 8'b10000000 : 8'b10000100;
				assign node4242 = (inp[5]) ? node4396 : node4243;
					assign node4243 = (inp[0]) ? node4245 : 8'b00000010;
						assign node4245 = (inp[1]) ? node4299 : node4246;
							assign node4246 = (inp[10]) ? node4280 : node4247;
								assign node4247 = (inp[8]) ? node4265 : node4248;
									assign node4248 = (inp[13]) ? node4256 : node4249;
										assign node4249 = (inp[2]) ? node4251 : 8'b00000010;
											assign node4251 = (inp[6]) ? 8'b00000010 : node4252;
												assign node4252 = (inp[11]) ? 8'b11110101 : 8'b10010000;
										assign node4256 = (inp[9]) ? 8'b00000010 : node4257;
											assign node4257 = (inp[6]) ? 8'b10100000 : node4258;
												assign node4258 = (inp[2]) ? node4260 : 8'b10100000;
													assign node4260 = (inp[11]) ? 8'b10010101 : 8'b10110000;
									assign node4265 = (inp[11]) ? node4273 : node4266;
										assign node4266 = (inp[9]) ? node4270 : node4267;
											assign node4267 = (inp[13]) ? 8'b10100100 : 8'b10010100;
											assign node4270 = (inp[2]) ? 8'b10010100 : 8'b10000100;
										assign node4273 = (inp[13]) ? node4275 : 8'b10100100;
											assign node4275 = (inp[9]) ? node4277 : 8'b10000100;
												assign node4277 = (inp[6]) ? 8'b10100100 : 8'b10110001;
								assign node4280 = (inp[13]) ? node4286 : node4281;
									assign node4281 = (inp[6]) ? 8'b00000010 : node4282;
										assign node4282 = (inp[2]) ? 8'b10010000 : 8'b00000010;
									assign node4286 = (inp[9]) ? node4292 : node4287;
										assign node4287 = (inp[6]) ? 8'b10100000 : node4288;
											assign node4288 = (inp[2]) ? 8'b10010101 : 8'b10100000;
										assign node4292 = (inp[6]) ? 8'b00000010 : node4293;
											assign node4293 = (inp[2]) ? node4295 : 8'b00000010;
												assign node4295 = (inp[11]) ? 8'b11110101 : 8'b10010000;
							assign node4299 = (inp[3]) ? node4355 : node4300;
								assign node4300 = (inp[11]) ? node4330 : node4301;
									assign node4301 = (inp[8]) ? node4317 : node4302;
										assign node4302 = (inp[9]) ? node4312 : node4303;
											assign node4303 = (inp[13]) ? node4307 : node4304;
												assign node4304 = (inp[2]) ? 8'b10010001 : 8'b10000001;
												assign node4307 = (inp[2]) ? node4309 : 8'b10100001;
													assign node4309 = (inp[6]) ? 8'b10100001 : 8'b10110001;
											assign node4312 = (inp[6]) ? 8'b10000001 : node4313;
												assign node4313 = (inp[2]) ? 8'b10010001 : 8'b10000001;
										assign node4317 = (inp[10]) ? node4327 : node4318;
											assign node4318 = (inp[2]) ? node4322 : node4319;
												assign node4319 = (inp[9]) ? 8'b10000101 : 8'b10100101;
												assign node4322 = (inp[6]) ? 8'b10000101 : node4323;
													assign node4323 = (inp[9]) ? 8'b10010101 : 8'b11110101;
											assign node4327 = (inp[6]) ? 8'b10000001 : 8'b10010001;
									assign node4330 = (inp[2]) ? node4344 : node4331;
										assign node4331 = (inp[10]) ? node4339 : node4332;
											assign node4332 = (inp[8]) ? node4334 : 8'b10100101;
												assign node4334 = (inp[6]) ? 8'b10100001 : node4335;
													assign node4335 = (inp[9]) ? 8'b10100001 : 8'b10000001;
											assign node4339 = (inp[13]) ? node4341 : 8'b10100101;
												assign node4341 = (inp[9]) ? 8'b10100101 : 8'b10000101;
										assign node4344 = (inp[6]) ? node4350 : node4345;
											assign node4345 = (inp[10]) ? 8'b10110100 : node4346;
												assign node4346 = (inp[8]) ? 8'b10110000 : 8'b10110100;
											assign node4350 = (inp[8]) ? node4352 : 8'b10100101;
												assign node4352 = (inp[13]) ? 8'b10000101 : 8'b10100101;
								assign node4355 = (inp[2]) ? node4375 : node4356;
									assign node4356 = (inp[10]) ? node4370 : node4357;
										assign node4357 = (inp[8]) ? node4361 : node4358;
											assign node4358 = (inp[11]) ? 8'b10100000 : 8'b00000010;
											assign node4361 = (inp[13]) ? node4363 : 8'b10100100;
												assign node4363 = (inp[11]) ? node4367 : node4364;
													assign node4364 = (inp[6]) ? 8'b10000100 : 8'b10100100;
													assign node4367 = (inp[9]) ? 8'b10100100 : 8'b10000100;
										assign node4370 = (inp[9]) ? 8'b00000010 : node4371;
											assign node4371 = (inp[13]) ? 8'b10100000 : 8'b00000010;
									assign node4375 = (inp[6]) ? node4391 : node4376;
										assign node4376 = (inp[11]) ? node4382 : node4377;
											assign node4377 = (inp[8]) ? node4379 : 8'b10010000;
												assign node4379 = (inp[9]) ? 8'b10010100 : 8'b10010000;
											assign node4382 = (inp[10]) ? node4388 : node4383;
												assign node4383 = (inp[13]) ? node4385 : 8'b10110001;
													assign node4385 = (inp[9]) ? 8'b10110001 : 8'b10010001;
												assign node4388 = (inp[8]) ? 8'b11110101 : 8'b10010101;
										assign node4391 = (inp[8]) ? node4393 : 8'b00000010;
											assign node4393 = (inp[10]) ? 8'b10100000 : 8'b10100100;
					assign node4396 = (inp[2]) ? node4478 : node4397;
						assign node4397 = (inp[1]) ? node4439 : node4398;
							assign node4398 = (inp[8]) ? node4406 : node4399;
								assign node4399 = (inp[13]) ? node4401 : 8'b00000010;
									assign node4401 = (inp[0]) ? 8'b10100000 : node4402;
										assign node4402 = (inp[9]) ? 8'b10100000 : 8'b00000010;
								assign node4406 = (inp[10]) ? node4424 : node4407;
									assign node4407 = (inp[0]) ? node4413 : node4408;
										assign node4408 = (inp[3]) ? node4410 : 8'b00000010;
											assign node4410 = (inp[6]) ? 8'b00000010 : 8'b10100000;
										assign node4413 = (inp[3]) ? node4415 : 8'b10000100;
											assign node4415 = (inp[9]) ? node4421 : node4416;
												assign node4416 = (inp[11]) ? 8'b10100100 : node4417;
													assign node4417 = (inp[13]) ? 8'b10100100 : 8'b10000100;
												assign node4421 = (inp[6]) ? 8'b10000100 : 8'b10100100;
									assign node4424 = (inp[11]) ? node4432 : node4425;
										assign node4425 = (inp[13]) ? node4427 : 8'b10000100;
											assign node4427 = (inp[0]) ? 8'b10100100 : node4428;
												assign node4428 = (inp[9]) ? 8'b10100100 : 8'b10000100;
										assign node4432 = (inp[13]) ? node4434 : 8'b10100100;
											assign node4434 = (inp[9]) ? 8'b10000100 : node4435;
												assign node4435 = (inp[0]) ? 8'b10000100 : 8'b10100100;
							assign node4439 = (inp[0]) ? node4463 : node4440;
								assign node4440 = (inp[3]) ? node4446 : node4441;
									assign node4441 = (inp[10]) ? node4443 : 8'b00000010;
										assign node4443 = (inp[8]) ? 8'b10100100 : 8'b00000010;
									assign node4446 = (inp[11]) ? node4456 : node4447;
										assign node4447 = (inp[8]) ? node4451 : node4448;
											assign node4448 = (inp[9]) ? 8'b10100001 : 8'b10000001;
											assign node4451 = (inp[10]) ? node4453 : 8'b10000001;
												assign node4453 = (inp[13]) ? 8'b10100101 : 8'b10000101;
										assign node4456 = (inp[10]) ? node4458 : 8'b10100101;
											assign node4458 = (inp[13]) ? node4460 : 8'b10100101;
												assign node4460 = (inp[8]) ? 8'b10000001 : 8'b10000101;
								assign node4463 = (inp[13]) ? node4471 : node4464;
									assign node4464 = (inp[11]) ? node4468 : node4465;
										assign node4465 = (inp[8]) ? 8'b10000101 : 8'b10000001;
										assign node4468 = (inp[8]) ? 8'b10100001 : 8'b10100101;
									assign node4471 = (inp[11]) ? node4475 : node4472;
										assign node4472 = (inp[8]) ? 8'b10100101 : 8'b10100001;
										assign node4475 = (inp[8]) ? 8'b10000001 : 8'b10000101;
						assign node4478 = (inp[0]) ? node4568 : node4479;
							assign node4479 = (inp[6]) ? node4527 : node4480;
								assign node4480 = (inp[1]) ? node4498 : node4481;
									assign node4481 = (inp[9]) ? node4489 : node4482;
										assign node4482 = (inp[10]) ? node4484 : 8'b00000010;
											assign node4484 = (inp[8]) ? node4486 : 8'b00000010;
												assign node4486 = (inp[3]) ? 8'b10000100 : 8'b10100100;
										assign node4489 = (inp[10]) ? node4493 : node4490;
											assign node4490 = (inp[13]) ? 8'b10100000 : 8'b00000010;
											assign node4493 = (inp[13]) ? 8'b10100000 : node4494;
												assign node4494 = (inp[11]) ? 8'b10100100 : 8'b10000100;
									assign node4498 = (inp[3]) ? node4512 : node4499;
										assign node4499 = (inp[10]) ? node4505 : node4500;
											assign node4500 = (inp[9]) ? node4502 : 8'b00000010;
												assign node4502 = (inp[13]) ? 8'b10100000 : 8'b00000010;
											assign node4505 = (inp[11]) ? node4509 : node4506;
												assign node4506 = (inp[13]) ? 8'b10100100 : 8'b10000100;
												assign node4509 = (inp[13]) ? 8'b10000100 : 8'b10100100;
										assign node4512 = (inp[11]) ? node4520 : node4513;
											assign node4513 = (inp[13]) ? 8'b10100001 : node4514;
												assign node4514 = (inp[10]) ? node4516 : 8'b10000001;
													assign node4516 = (inp[8]) ? 8'b10000101 : 8'b10000001;
											assign node4520 = (inp[8]) ? node4522 : 8'b10100101;
												assign node4522 = (inp[9]) ? 8'b10000001 : node4523;
													assign node4523 = (inp[10]) ? 8'b10100001 : 8'b10100101;
								assign node4527 = (inp[11]) ? node4549 : node4528;
									assign node4528 = (inp[8]) ? node4536 : node4529;
										assign node4529 = (inp[13]) ? node4531 : 8'b10010000;
											assign node4531 = (inp[1]) ? 8'b10010001 : node4532;
												assign node4532 = (inp[9]) ? 8'b10110000 : 8'b10010000;
										assign node4536 = (inp[10]) ? node4542 : node4537;
											assign node4537 = (inp[1]) ? node4539 : 8'b10110000;
												assign node4539 = (inp[3]) ? 8'b10010001 : 8'b10010000;
											assign node4542 = (inp[1]) ? node4544 : 8'b10010100;
												assign node4544 = (inp[13]) ? 8'b11110101 : node4545;
													assign node4545 = (inp[9]) ? 8'b10010101 : 8'b10010100;
									assign node4549 = (inp[9]) ? node4557 : node4550;
										assign node4550 = (inp[8]) ? node4552 : 8'b11110101;
											assign node4552 = (inp[10]) ? 8'b10110001 : node4553;
												assign node4553 = (inp[3]) ? 8'b10110100 : 8'b11110101;
										assign node4557 = (inp[1]) ? node4561 : node4558;
											assign node4558 = (inp[13]) ? 8'b10010001 : 8'b10110001;
											assign node4561 = (inp[13]) ? node4563 : 8'b10110100;
												assign node4563 = (inp[3]) ? node4565 : 8'b10010101;
													assign node4565 = (inp[10]) ? 8'b10010000 : 8'b10010100;
							assign node4568 = (inp[11]) ? node4582 : node4569;
								assign node4569 = (inp[13]) ? node4577 : node4570;
									assign node4570 = (inp[8]) ? node4574 : node4571;
										assign node4571 = (inp[1]) ? 8'b10010001 : 8'b10010000;
										assign node4574 = (inp[1]) ? 8'b10010101 : 8'b10010100;
									assign node4577 = (inp[8]) ? 8'b11110101 : node4578;
										assign node4578 = (inp[1]) ? 8'b10110001 : 8'b10110000;
								assign node4582 = (inp[1]) ? node4590 : node4583;
									assign node4583 = (inp[13]) ? node4587 : node4584;
										assign node4584 = (inp[8]) ? 8'b10110001 : 8'b11110101;
										assign node4587 = (inp[8]) ? 8'b10010001 : 8'b10010101;
									assign node4590 = (inp[13]) ? node4594 : node4591;
										assign node4591 = (inp[8]) ? 8'b10110000 : 8'b10110100;
										assign node4594 = (inp[8]) ? 8'b10010000 : 8'b10010100;

endmodule