module dtc_split125_bm13 (
	input  wire [11-1:0] inp,
	output wire [1-1:0] outp
);

	wire [1-1:0] node1;
	wire [1-1:0] node2;
	wire [1-1:0] node3;
	wire [1-1:0] node5;
	wire [1-1:0] node7;
	wire [1-1:0] node9;
	wire [1-1:0] node10;
	wire [1-1:0] node12;
	wire [1-1:0] node16;
	wire [1-1:0] node17;
	wire [1-1:0] node19;
	wire [1-1:0] node21;
	wire [1-1:0] node22;
	wire [1-1:0] node26;
	wire [1-1:0] node27;
	wire [1-1:0] node29;
	wire [1-1:0] node31;
	wire [1-1:0] node32;
	wire [1-1:0] node36;
	wire [1-1:0] node37;
	wire [1-1:0] node41;
	wire [1-1:0] node42;
	wire [1-1:0] node43;
	wire [1-1:0] node45;
	wire [1-1:0] node48;
	wire [1-1:0] node49;
	wire [1-1:0] node51;
	wire [1-1:0] node54;
	wire [1-1:0] node55;
	wire [1-1:0] node59;
	wire [1-1:0] node60;
	wire [1-1:0] node62;
	wire [1-1:0] node63;
	wire [1-1:0] node65;
	wire [1-1:0] node67;
	wire [1-1:0] node68;
	wire [1-1:0] node73;
	wire [1-1:0] node74;
	wire [1-1:0] node75;
	wire [1-1:0] node80;
	wire [1-1:0] node81;
	wire [1-1:0] node82;
	wire [1-1:0] node83;
	wire [1-1:0] node85;
	wire [1-1:0] node87;
	wire [1-1:0] node90;
	wire [1-1:0] node91;
	wire [1-1:0] node93;
	wire [1-1:0] node97;
	wire [1-1:0] node98;
	wire [1-1:0] node99;
	wire [1-1:0] node101;
	wire [1-1:0] node103;
	wire [1-1:0] node104;
	wire [1-1:0] node108;
	wire [1-1:0] node109;
	wire [1-1:0] node111;
	wire [1-1:0] node115;
	wire [1-1:0] node116;
	wire [1-1:0] node117;
	wire [1-1:0] node119;
	wire [1-1:0] node120;
	wire [1-1:0] node126;
	wire [1-1:0] node127;
	wire [1-1:0] node128;
	wire [1-1:0] node129;
	wire [1-1:0] node131;
	wire [1-1:0] node134;
	wire [1-1:0] node135;
	wire [1-1:0] node136;
	wire [1-1:0] node137;
	wire [1-1:0] node143;
	wire [1-1:0] node144;
	wire [1-1:0] node145;

	assign outp = (inp[8]) ? node80 : node1;
		assign node1 = (inp[3]) ? node41 : node2;
			assign node2 = (inp[4]) ? node16 : node3;
				assign node3 = (inp[10]) ? node5 : 1'b1;
					assign node5 = (inp[6]) ? node7 : 1'b1;
						assign node7 = (inp[5]) ? node9 : 1'b1;
							assign node9 = (inp[7]) ? 1'b0 : node10;
								assign node10 = (inp[9]) ? node12 : 1'b1;
									assign node12 = (inp[1]) ? 1'b0 : 1'b1;
				assign node16 = (inp[0]) ? node26 : node17;
					assign node17 = (inp[7]) ? node19 : 1'b1;
						assign node19 = (inp[5]) ? node21 : 1'b1;
							assign node21 = (inp[1]) ? 1'b0 : node22;
								assign node22 = (inp[10]) ? 1'b0 : 1'b1;
					assign node26 = (inp[5]) ? node36 : node27;
						assign node27 = (inp[6]) ? node29 : 1'b1;
							assign node29 = (inp[1]) ? node31 : 1'b1;
								assign node31 = (inp[2]) ? 1'b0 : node32;
									assign node32 = (inp[9]) ? 1'b0 : 1'b1;
						assign node36 = (inp[9]) ? 1'b0 : node37;
							assign node37 = (inp[6]) ? 1'b1 : 1'b0;
			assign node41 = (inp[1]) ? node59 : node42;
				assign node42 = (inp[5]) ? node48 : node43;
					assign node43 = (inp[2]) ? node45 : 1'b1;
						assign node45 = (inp[7]) ? 1'b0 : 1'b1;
					assign node48 = (inp[0]) ? node54 : node49;
						assign node49 = (inp[4]) ? node51 : 1'b1;
							assign node51 = (inp[7]) ? 1'b0 : 1'b1;
						assign node54 = (inp[7]) ? 1'b0 : node55;
							assign node55 = (inp[2]) ? 1'b0 : 1'b1;
				assign node59 = (inp[10]) ? node73 : node60;
					assign node60 = (inp[0]) ? node62 : 1'b1;
						assign node62 = (inp[9]) ? 1'b0 : node63;
							assign node63 = (inp[4]) ? node65 : 1'b1;
								assign node65 = (inp[5]) ? node67 : 1'b1;
									assign node67 = (inp[2]) ? 1'b0 : node68;
										assign node68 = (inp[7]) ? 1'b0 : 1'b1;
					assign node73 = (inp[7]) ? 1'b0 : node74;
						assign node74 = (inp[6]) ? 1'b0 : node75;
							assign node75 = (inp[0]) ? 1'b0 : 1'b1;
		assign node80 = (inp[4]) ? node126 : node81;
			assign node81 = (inp[3]) ? node97 : node82;
				assign node82 = (inp[7]) ? node90 : node83;
					assign node83 = (inp[5]) ? node85 : 1'b1;
						assign node85 = (inp[9]) ? node87 : 1'b1;
							assign node87 = (inp[2]) ? 1'b0 : 1'b1;
					assign node90 = (inp[9]) ? 1'b0 : node91;
						assign node91 = (inp[10]) ? node93 : 1'b1;
							assign node93 = (inp[1]) ? 1'b1 : 1'b0;
				assign node97 = (inp[2]) ? node115 : node98;
					assign node98 = (inp[9]) ? node108 : node99;
						assign node99 = (inp[5]) ? node101 : 1'b1;
							assign node101 = (inp[10]) ? node103 : 1'b1;
								assign node103 = (inp[7]) ? 1'b0 : node104;
									assign node104 = (inp[1]) ? 1'b0 : 1'b1;
						assign node108 = (inp[6]) ? 1'b0 : node109;
							assign node109 = (inp[1]) ? node111 : 1'b1;
								assign node111 = (inp[7]) ? 1'b0 : 1'b1;
					assign node115 = (inp[5]) ? 1'b0 : node116;
						assign node116 = (inp[1]) ? 1'b0 : node117;
							assign node117 = (inp[10]) ? node119 : 1'b1;
								assign node119 = (inp[9]) ? 1'b0 : node120;
									assign node120 = (inp[0]) ? 1'b0 : 1'b1;
			assign node126 = (inp[10]) ? 1'b0 : node127;
				assign node127 = (inp[9]) ? node143 : node128;
					assign node128 = (inp[6]) ? node134 : node129;
						assign node129 = (inp[5]) ? node131 : 1'b1;
							assign node131 = (inp[3]) ? 1'b0 : 1'b1;
						assign node134 = (inp[0]) ? 1'b0 : node135;
							assign node135 = (inp[5]) ? 1'b1 : node136;
								assign node136 = (inp[2]) ? 1'b0 : node137;
									assign node137 = (inp[7]) ? 1'b0 : 1'b1;
					assign node143 = (inp[1]) ? 1'b0 : node144;
						assign node144 = (inp[5]) ? 1'b0 : node145;
							assign node145 = (inp[3]) ? 1'b0 : 1'b1;

endmodule