module dtc_split66_bm62 (
	input  wire [16-1:0] inp,
	output wire [4-1:0] outp
);

	wire [4-1:0] node1;
	wire [4-1:0] node2;
	wire [4-1:0] node3;
	wire [4-1:0] node4;
	wire [4-1:0] node5;
	wire [4-1:0] node6;
	wire [4-1:0] node7;
	wire [4-1:0] node8;
	wire [4-1:0] node9;
	wire [4-1:0] node10;
	wire [4-1:0] node11;
	wire [4-1:0] node12;
	wire [4-1:0] node13;
	wire [4-1:0] node14;
	wire [4-1:0] node17;
	wire [4-1:0] node20;
	wire [4-1:0] node23;
	wire [4-1:0] node24;
	wire [4-1:0] node25;
	wire [4-1:0] node26;
	wire [4-1:0] node30;
	wire [4-1:0] node31;
	wire [4-1:0] node36;
	wire [4-1:0] node37;
	wire [4-1:0] node38;
	wire [4-1:0] node39;
	wire [4-1:0] node41;
	wire [4-1:0] node44;
	wire [4-1:0] node47;
	wire [4-1:0] node49;
	wire [4-1:0] node52;
	wire [4-1:0] node53;
	wire [4-1:0] node55;
	wire [4-1:0] node58;
	wire [4-1:0] node59;
	wire [4-1:0] node60;
	wire [4-1:0] node63;
	wire [4-1:0] node66;
	wire [4-1:0] node67;
	wire [4-1:0] node71;
	wire [4-1:0] node72;
	wire [4-1:0] node73;
	wire [4-1:0] node74;
	wire [4-1:0] node75;
	wire [4-1:0] node76;
	wire [4-1:0] node80;
	wire [4-1:0] node81;
	wire [4-1:0] node85;
	wire [4-1:0] node88;
	wire [4-1:0] node89;
	wire [4-1:0] node90;
	wire [4-1:0] node93;
	wire [4-1:0] node95;
	wire [4-1:0] node98;
	wire [4-1:0] node100;
	wire [4-1:0] node101;
	wire [4-1:0] node105;
	wire [4-1:0] node106;
	wire [4-1:0] node107;
	wire [4-1:0] node108;
	wire [4-1:0] node109;
	wire [4-1:0] node112;
	wire [4-1:0] node116;
	wire [4-1:0] node117;
	wire [4-1:0] node119;
	wire [4-1:0] node122;
	wire [4-1:0] node125;
	wire [4-1:0] node126;
	wire [4-1:0] node127;
	wire [4-1:0] node129;
	wire [4-1:0] node132;
	wire [4-1:0] node134;
	wire [4-1:0] node137;
	wire [4-1:0] node138;
	wire [4-1:0] node140;
	wire [4-1:0] node143;
	wire [4-1:0] node144;
	wire [4-1:0] node147;
	wire [4-1:0] node150;
	wire [4-1:0] node151;
	wire [4-1:0] node152;
	wire [4-1:0] node153;
	wire [4-1:0] node154;
	wire [4-1:0] node155;
	wire [4-1:0] node158;
	wire [4-1:0] node162;
	wire [4-1:0] node163;
	wire [4-1:0] node164;
	wire [4-1:0] node166;
	wire [4-1:0] node169;
	wire [4-1:0] node172;
	wire [4-1:0] node173;
	wire [4-1:0] node174;
	wire [4-1:0] node177;
	wire [4-1:0] node180;
	wire [4-1:0] node181;
	wire [4-1:0] node185;
	wire [4-1:0] node186;
	wire [4-1:0] node187;
	wire [4-1:0] node188;
	wire [4-1:0] node190;
	wire [4-1:0] node193;
	wire [4-1:0] node194;
	wire [4-1:0] node197;
	wire [4-1:0] node200;
	wire [4-1:0] node203;
	wire [4-1:0] node204;
	wire [4-1:0] node205;
	wire [4-1:0] node208;
	wire [4-1:0] node211;
	wire [4-1:0] node213;
	wire [4-1:0] node214;
	wire [4-1:0] node218;
	wire [4-1:0] node219;
	wire [4-1:0] node220;
	wire [4-1:0] node221;
	wire [4-1:0] node222;
	wire [4-1:0] node225;
	wire [4-1:0] node228;
	wire [4-1:0] node229;
	wire [4-1:0] node232;
	wire [4-1:0] node235;
	wire [4-1:0] node236;
	wire [4-1:0] node239;
	wire [4-1:0] node242;
	wire [4-1:0] node243;
	wire [4-1:0] node244;
	wire [4-1:0] node247;
	wire [4-1:0] node250;
	wire [4-1:0] node251;
	wire [4-1:0] node252;
	wire [4-1:0] node253;
	wire [4-1:0] node256;
	wire [4-1:0] node259;
	wire [4-1:0] node260;
	wire [4-1:0] node263;
	wire [4-1:0] node266;
	wire [4-1:0] node267;
	wire [4-1:0] node268;
	wire [4-1:0] node272;
	wire [4-1:0] node275;
	wire [4-1:0] node276;
	wire [4-1:0] node277;
	wire [4-1:0] node278;
	wire [4-1:0] node279;
	wire [4-1:0] node280;
	wire [4-1:0] node282;
	wire [4-1:0] node285;
	wire [4-1:0] node286;
	wire [4-1:0] node290;
	wire [4-1:0] node292;
	wire [4-1:0] node293;
	wire [4-1:0] node294;
	wire [4-1:0] node297;
	wire [4-1:0] node300;
	wire [4-1:0] node301;
	wire [4-1:0] node305;
	wire [4-1:0] node306;
	wire [4-1:0] node307;
	wire [4-1:0] node308;
	wire [4-1:0] node311;
	wire [4-1:0] node314;
	wire [4-1:0] node315;
	wire [4-1:0] node319;
	wire [4-1:0] node320;
	wire [4-1:0] node321;
	wire [4-1:0] node325;
	wire [4-1:0] node326;
	wire [4-1:0] node329;
	wire [4-1:0] node332;
	wire [4-1:0] node333;
	wire [4-1:0] node334;
	wire [4-1:0] node335;
	wire [4-1:0] node336;
	wire [4-1:0] node337;
	wire [4-1:0] node340;
	wire [4-1:0] node344;
	wire [4-1:0] node345;
	wire [4-1:0] node348;
	wire [4-1:0] node351;
	wire [4-1:0] node352;
	wire [4-1:0] node353;
	wire [4-1:0] node356;
	wire [4-1:0] node359;
	wire [4-1:0] node360;
	wire [4-1:0] node363;
	wire [4-1:0] node366;
	wire [4-1:0] node367;
	wire [4-1:0] node368;
	wire [4-1:0] node370;
	wire [4-1:0] node373;
	wire [4-1:0] node375;
	wire [4-1:0] node378;
	wire [4-1:0] node379;
	wire [4-1:0] node380;
	wire [4-1:0] node383;
	wire [4-1:0] node386;
	wire [4-1:0] node387;
	wire [4-1:0] node388;
	wire [4-1:0] node392;
	wire [4-1:0] node394;
	wire [4-1:0] node397;
	wire [4-1:0] node398;
	wire [4-1:0] node399;
	wire [4-1:0] node400;
	wire [4-1:0] node401;
	wire [4-1:0] node402;
	wire [4-1:0] node404;
	wire [4-1:0] node407;
	wire [4-1:0] node408;
	wire [4-1:0] node411;
	wire [4-1:0] node414;
	wire [4-1:0] node415;
	wire [4-1:0] node419;
	wire [4-1:0] node420;
	wire [4-1:0] node422;
	wire [4-1:0] node425;
	wire [4-1:0] node426;
	wire [4-1:0] node429;
	wire [4-1:0] node432;
	wire [4-1:0] node433;
	wire [4-1:0] node434;
	wire [4-1:0] node436;
	wire [4-1:0] node438;
	wire [4-1:0] node441;
	wire [4-1:0] node442;
	wire [4-1:0] node444;
	wire [4-1:0] node447;
	wire [4-1:0] node448;
	wire [4-1:0] node451;
	wire [4-1:0] node454;
	wire [4-1:0] node455;
	wire [4-1:0] node456;
	wire [4-1:0] node459;
	wire [4-1:0] node462;
	wire [4-1:0] node463;
	wire [4-1:0] node464;
	wire [4-1:0] node467;
	wire [4-1:0] node470;
	wire [4-1:0] node473;
	wire [4-1:0] node474;
	wire [4-1:0] node475;
	wire [4-1:0] node476;
	wire [4-1:0] node477;
	wire [4-1:0] node480;
	wire [4-1:0] node484;
	wire [4-1:0] node485;
	wire [4-1:0] node486;
	wire [4-1:0] node489;
	wire [4-1:0] node492;
	wire [4-1:0] node493;
	wire [4-1:0] node496;
	wire [4-1:0] node499;
	wire [4-1:0] node500;
	wire [4-1:0] node501;
	wire [4-1:0] node504;
	wire [4-1:0] node507;
	wire [4-1:0] node508;
	wire [4-1:0] node509;
	wire [4-1:0] node512;
	wire [4-1:0] node515;
	wire [4-1:0] node517;
	wire [4-1:0] node519;
	wire [4-1:0] node522;
	wire [4-1:0] node523;
	wire [4-1:0] node524;
	wire [4-1:0] node525;
	wire [4-1:0] node526;
	wire [4-1:0] node527;
	wire [4-1:0] node528;
	wire [4-1:0] node530;
	wire [4-1:0] node534;
	wire [4-1:0] node535;
	wire [4-1:0] node537;
	wire [4-1:0] node540;
	wire [4-1:0] node542;
	wire [4-1:0] node545;
	wire [4-1:0] node546;
	wire [4-1:0] node547;
	wire [4-1:0] node550;
	wire [4-1:0] node553;
	wire [4-1:0] node555;
	wire [4-1:0] node556;
	wire [4-1:0] node557;
	wire [4-1:0] node560;
	wire [4-1:0] node564;
	wire [4-1:0] node565;
	wire [4-1:0] node566;
	wire [4-1:0] node567;
	wire [4-1:0] node569;
	wire [4-1:0] node572;
	wire [4-1:0] node574;
	wire [4-1:0] node577;
	wire [4-1:0] node578;
	wire [4-1:0] node580;
	wire [4-1:0] node583;
	wire [4-1:0] node585;
	wire [4-1:0] node588;
	wire [4-1:0] node589;
	wire [4-1:0] node590;
	wire [4-1:0] node591;
	wire [4-1:0] node595;
	wire [4-1:0] node598;
	wire [4-1:0] node599;
	wire [4-1:0] node602;
	wire [4-1:0] node605;
	wire [4-1:0] node606;
	wire [4-1:0] node607;
	wire [4-1:0] node608;
	wire [4-1:0] node609;
	wire [4-1:0] node610;
	wire [4-1:0] node613;
	wire [4-1:0] node616;
	wire [4-1:0] node617;
	wire [4-1:0] node618;
	wire [4-1:0] node621;
	wire [4-1:0] node625;
	wire [4-1:0] node626;
	wire [4-1:0] node627;
	wire [4-1:0] node630;
	wire [4-1:0] node633;
	wire [4-1:0] node634;
	wire [4-1:0] node635;
	wire [4-1:0] node638;
	wire [4-1:0] node641;
	wire [4-1:0] node642;
	wire [4-1:0] node645;
	wire [4-1:0] node648;
	wire [4-1:0] node649;
	wire [4-1:0] node650;
	wire [4-1:0] node651;
	wire [4-1:0] node654;
	wire [4-1:0] node657;
	wire [4-1:0] node659;
	wire [4-1:0] node662;
	wire [4-1:0] node663;
	wire [4-1:0] node664;
	wire [4-1:0] node667;
	wire [4-1:0] node669;
	wire [4-1:0] node672;
	wire [4-1:0] node673;
	wire [4-1:0] node675;
	wire [4-1:0] node678;
	wire [4-1:0] node679;
	wire [4-1:0] node683;
	wire [4-1:0] node684;
	wire [4-1:0] node685;
	wire [4-1:0] node686;
	wire [4-1:0] node687;
	wire [4-1:0] node690;
	wire [4-1:0] node693;
	wire [4-1:0] node694;
	wire [4-1:0] node697;
	wire [4-1:0] node698;
	wire [4-1:0] node702;
	wire [4-1:0] node703;
	wire [4-1:0] node704;
	wire [4-1:0] node706;
	wire [4-1:0] node709;
	wire [4-1:0] node710;
	wire [4-1:0] node714;
	wire [4-1:0] node715;
	wire [4-1:0] node717;
	wire [4-1:0] node720;
	wire [4-1:0] node723;
	wire [4-1:0] node724;
	wire [4-1:0] node725;
	wire [4-1:0] node726;
	wire [4-1:0] node729;
	wire [4-1:0] node732;
	wire [4-1:0] node733;
	wire [4-1:0] node734;
	wire [4-1:0] node737;
	wire [4-1:0] node741;
	wire [4-1:0] node742;
	wire [4-1:0] node744;
	wire [4-1:0] node745;
	wire [4-1:0] node749;
	wire [4-1:0] node750;
	wire [4-1:0] node752;
	wire [4-1:0] node755;
	wire [4-1:0] node757;
	wire [4-1:0] node760;
	wire [4-1:0] node761;
	wire [4-1:0] node762;
	wire [4-1:0] node763;
	wire [4-1:0] node764;
	wire [4-1:0] node765;
	wire [4-1:0] node768;
	wire [4-1:0] node771;
	wire [4-1:0] node772;
	wire [4-1:0] node774;
	wire [4-1:0] node775;
	wire [4-1:0] node778;
	wire [4-1:0] node781;
	wire [4-1:0] node782;
	wire [4-1:0] node785;
	wire [4-1:0] node788;
	wire [4-1:0] node789;
	wire [4-1:0] node790;
	wire [4-1:0] node791;
	wire [4-1:0] node794;
	wire [4-1:0] node797;
	wire [4-1:0] node798;
	wire [4-1:0] node801;
	wire [4-1:0] node804;
	wire [4-1:0] node805;
	wire [4-1:0] node806;
	wire [4-1:0] node809;
	wire [4-1:0] node812;
	wire [4-1:0] node813;
	wire [4-1:0] node814;
	wire [4-1:0] node817;
	wire [4-1:0] node820;
	wire [4-1:0] node821;
	wire [4-1:0] node825;
	wire [4-1:0] node826;
	wire [4-1:0] node827;
	wire [4-1:0] node828;
	wire [4-1:0] node831;
	wire [4-1:0] node833;
	wire [4-1:0] node836;
	wire [4-1:0] node837;
	wire [4-1:0] node838;
	wire [4-1:0] node840;
	wire [4-1:0] node843;
	wire [4-1:0] node846;
	wire [4-1:0] node848;
	wire [4-1:0] node849;
	wire [4-1:0] node852;
	wire [4-1:0] node855;
	wire [4-1:0] node856;
	wire [4-1:0] node857;
	wire [4-1:0] node859;
	wire [4-1:0] node863;
	wire [4-1:0] node864;
	wire [4-1:0] node866;
	wire [4-1:0] node870;
	wire [4-1:0] node871;
	wire [4-1:0] node872;
	wire [4-1:0] node873;
	wire [4-1:0] node874;
	wire [4-1:0] node876;
	wire [4-1:0] node879;
	wire [4-1:0] node880;
	wire [4-1:0] node883;
	wire [4-1:0] node886;
	wire [4-1:0] node887;
	wire [4-1:0] node889;
	wire [4-1:0] node890;
	wire [4-1:0] node894;
	wire [4-1:0] node895;
	wire [4-1:0] node899;
	wire [4-1:0] node900;
	wire [4-1:0] node901;
	wire [4-1:0] node903;
	wire [4-1:0] node906;
	wire [4-1:0] node908;
	wire [4-1:0] node911;
	wire [4-1:0] node912;
	wire [4-1:0] node914;
	wire [4-1:0] node917;
	wire [4-1:0] node919;
	wire [4-1:0] node922;
	wire [4-1:0] node923;
	wire [4-1:0] node924;
	wire [4-1:0] node925;
	wire [4-1:0] node926;
	wire [4-1:0] node929;
	wire [4-1:0] node932;
	wire [4-1:0] node933;
	wire [4-1:0] node936;
	wire [4-1:0] node939;
	wire [4-1:0] node940;
	wire [4-1:0] node941;
	wire [4-1:0] node943;
	wire [4-1:0] node946;
	wire [4-1:0] node949;
	wire [4-1:0] node950;
	wire [4-1:0] node954;
	wire [4-1:0] node955;
	wire [4-1:0] node956;
	wire [4-1:0] node959;
	wire [4-1:0] node960;
	wire [4-1:0] node964;
	wire [4-1:0] node965;
	wire [4-1:0] node966;
	wire [4-1:0] node970;
	wire [4-1:0] node971;
	wire [4-1:0] node975;
	wire [4-1:0] node976;
	wire [4-1:0] node977;
	wire [4-1:0] node978;
	wire [4-1:0] node979;
	wire [4-1:0] node980;
	wire [4-1:0] node981;
	wire [4-1:0] node984;
	wire [4-1:0] node987;
	wire [4-1:0] node988;
	wire [4-1:0] node989;
	wire [4-1:0] node992;
	wire [4-1:0] node995;
	wire [4-1:0] node996;
	wire [4-1:0] node999;
	wire [4-1:0] node1002;
	wire [4-1:0] node1003;
	wire [4-1:0] node1004;
	wire [4-1:0] node1005;
	wire [4-1:0] node1006;
	wire [4-1:0] node1009;
	wire [4-1:0] node1012;
	wire [4-1:0] node1013;
	wire [4-1:0] node1016;
	wire [4-1:0] node1019;
	wire [4-1:0] node1020;
	wire [4-1:0] node1021;
	wire [4-1:0] node1023;
	wire [4-1:0] node1027;
	wire [4-1:0] node1028;
	wire [4-1:0] node1029;
	wire [4-1:0] node1032;
	wire [4-1:0] node1036;
	wire [4-1:0] node1037;
	wire [4-1:0] node1039;
	wire [4-1:0] node1040;
	wire [4-1:0] node1042;
	wire [4-1:0] node1045;
	wire [4-1:0] node1046;
	wire [4-1:0] node1049;
	wire [4-1:0] node1052;
	wire [4-1:0] node1054;
	wire [4-1:0] node1056;
	wire [4-1:0] node1059;
	wire [4-1:0] node1060;
	wire [4-1:0] node1061;
	wire [4-1:0] node1062;
	wire [4-1:0] node1063;
	wire [4-1:0] node1066;
	wire [4-1:0] node1069;
	wire [4-1:0] node1070;
	wire [4-1:0] node1071;
	wire [4-1:0] node1074;
	wire [4-1:0] node1077;
	wire [4-1:0] node1078;
	wire [4-1:0] node1081;
	wire [4-1:0] node1084;
	wire [4-1:0] node1085;
	wire [4-1:0] node1086;
	wire [4-1:0] node1088;
	wire [4-1:0] node1091;
	wire [4-1:0] node1092;
	wire [4-1:0] node1093;
	wire [4-1:0] node1097;
	wire [4-1:0] node1098;
	wire [4-1:0] node1102;
	wire [4-1:0] node1103;
	wire [4-1:0] node1104;
	wire [4-1:0] node1105;
	wire [4-1:0] node1109;
	wire [4-1:0] node1111;
	wire [4-1:0] node1114;
	wire [4-1:0] node1115;
	wire [4-1:0] node1117;
	wire [4-1:0] node1121;
	wire [4-1:0] node1122;
	wire [4-1:0] node1123;
	wire [4-1:0] node1124;
	wire [4-1:0] node1125;
	wire [4-1:0] node1127;
	wire [4-1:0] node1131;
	wire [4-1:0] node1132;
	wire [4-1:0] node1133;
	wire [4-1:0] node1137;
	wire [4-1:0] node1138;
	wire [4-1:0] node1141;
	wire [4-1:0] node1144;
	wire [4-1:0] node1145;
	wire [4-1:0] node1146;
	wire [4-1:0] node1149;
	wire [4-1:0] node1153;
	wire [4-1:0] node1154;
	wire [4-1:0] node1155;
	wire [4-1:0] node1156;
	wire [4-1:0] node1157;
	wire [4-1:0] node1161;
	wire [4-1:0] node1163;
	wire [4-1:0] node1166;
	wire [4-1:0] node1167;
	wire [4-1:0] node1171;
	wire [4-1:0] node1172;
	wire [4-1:0] node1173;
	wire [4-1:0] node1176;
	wire [4-1:0] node1179;
	wire [4-1:0] node1180;
	wire [4-1:0] node1183;
	wire [4-1:0] node1186;
	wire [4-1:0] node1187;
	wire [4-1:0] node1188;
	wire [4-1:0] node1189;
	wire [4-1:0] node1190;
	wire [4-1:0] node1191;
	wire [4-1:0] node1192;
	wire [4-1:0] node1193;
	wire [4-1:0] node1196;
	wire [4-1:0] node1199;
	wire [4-1:0] node1200;
	wire [4-1:0] node1204;
	wire [4-1:0] node1205;
	wire [4-1:0] node1206;
	wire [4-1:0] node1210;
	wire [4-1:0] node1211;
	wire [4-1:0] node1214;
	wire [4-1:0] node1217;
	wire [4-1:0] node1218;
	wire [4-1:0] node1220;
	wire [4-1:0] node1223;
	wire [4-1:0] node1225;
	wire [4-1:0] node1226;
	wire [4-1:0] node1230;
	wire [4-1:0] node1231;
	wire [4-1:0] node1232;
	wire [4-1:0] node1234;
	wire [4-1:0] node1235;
	wire [4-1:0] node1238;
	wire [4-1:0] node1241;
	wire [4-1:0] node1242;
	wire [4-1:0] node1245;
	wire [4-1:0] node1248;
	wire [4-1:0] node1249;
	wire [4-1:0] node1250;
	wire [4-1:0] node1253;
	wire [4-1:0] node1256;
	wire [4-1:0] node1258;
	wire [4-1:0] node1261;
	wire [4-1:0] node1262;
	wire [4-1:0] node1263;
	wire [4-1:0] node1264;
	wire [4-1:0] node1265;
	wire [4-1:0] node1268;
	wire [4-1:0] node1271;
	wire [4-1:0] node1273;
	wire [4-1:0] node1276;
	wire [4-1:0] node1278;
	wire [4-1:0] node1279;
	wire [4-1:0] node1282;
	wire [4-1:0] node1285;
	wire [4-1:0] node1286;
	wire [4-1:0] node1287;
	wire [4-1:0] node1289;
	wire [4-1:0] node1290;
	wire [4-1:0] node1293;
	wire [4-1:0] node1296;
	wire [4-1:0] node1298;
	wire [4-1:0] node1299;
	wire [4-1:0] node1302;
	wire [4-1:0] node1305;
	wire [4-1:0] node1306;
	wire [4-1:0] node1308;
	wire [4-1:0] node1309;
	wire [4-1:0] node1314;
	wire [4-1:0] node1315;
	wire [4-1:0] node1316;
	wire [4-1:0] node1317;
	wire [4-1:0] node1318;
	wire [4-1:0] node1319;
	wire [4-1:0] node1321;
	wire [4-1:0] node1324;
	wire [4-1:0] node1327;
	wire [4-1:0] node1330;
	wire [4-1:0] node1331;
	wire [4-1:0] node1332;
	wire [4-1:0] node1335;
	wire [4-1:0] node1338;
	wire [4-1:0] node1339;
	wire [4-1:0] node1342;
	wire [4-1:0] node1345;
	wire [4-1:0] node1346;
	wire [4-1:0] node1347;
	wire [4-1:0] node1348;
	wire [4-1:0] node1351;
	wire [4-1:0] node1354;
	wire [4-1:0] node1355;
	wire [4-1:0] node1358;
	wire [4-1:0] node1361;
	wire [4-1:0] node1363;
	wire [4-1:0] node1365;
	wire [4-1:0] node1368;
	wire [4-1:0] node1369;
	wire [4-1:0] node1370;
	wire [4-1:0] node1371;
	wire [4-1:0] node1373;
	wire [4-1:0] node1375;
	wire [4-1:0] node1378;
	wire [4-1:0] node1379;
	wire [4-1:0] node1382;
	wire [4-1:0] node1385;
	wire [4-1:0] node1386;
	wire [4-1:0] node1389;
	wire [4-1:0] node1392;
	wire [4-1:0] node1393;
	wire [4-1:0] node1395;
	wire [4-1:0] node1396;
	wire [4-1:0] node1399;
	wire [4-1:0] node1402;
	wire [4-1:0] node1403;
	wire [4-1:0] node1404;
	wire [4-1:0] node1407;
	wire [4-1:0] node1410;
	wire [4-1:0] node1411;
	wire [4-1:0] node1414;
	wire [4-1:0] node1417;
	wire [4-1:0] node1418;
	wire [4-1:0] node1419;
	wire [4-1:0] node1420;
	wire [4-1:0] node1421;
	wire [4-1:0] node1422;
	wire [4-1:0] node1423;
	wire [4-1:0] node1424;
	wire [4-1:0] node1425;
	wire [4-1:0] node1428;
	wire [4-1:0] node1431;
	wire [4-1:0] node1432;
	wire [4-1:0] node1436;
	wire [4-1:0] node1438;
	wire [4-1:0] node1439;
	wire [4-1:0] node1442;
	wire [4-1:0] node1445;
	wire [4-1:0] node1446;
	wire [4-1:0] node1447;
	wire [4-1:0] node1448;
	wire [4-1:0] node1452;
	wire [4-1:0] node1453;
	wire [4-1:0] node1456;
	wire [4-1:0] node1459;
	wire [4-1:0] node1460;
	wire [4-1:0] node1462;
	wire [4-1:0] node1465;
	wire [4-1:0] node1466;
	wire [4-1:0] node1469;
	wire [4-1:0] node1472;
	wire [4-1:0] node1473;
	wire [4-1:0] node1474;
	wire [4-1:0] node1475;
	wire [4-1:0] node1478;
	wire [4-1:0] node1479;
	wire [4-1:0] node1482;
	wire [4-1:0] node1485;
	wire [4-1:0] node1486;
	wire [4-1:0] node1488;
	wire [4-1:0] node1492;
	wire [4-1:0] node1493;
	wire [4-1:0] node1494;
	wire [4-1:0] node1496;
	wire [4-1:0] node1499;
	wire [4-1:0] node1502;
	wire [4-1:0] node1503;
	wire [4-1:0] node1505;
	wire [4-1:0] node1508;
	wire [4-1:0] node1511;
	wire [4-1:0] node1512;
	wire [4-1:0] node1513;
	wire [4-1:0] node1514;
	wire [4-1:0] node1515;
	wire [4-1:0] node1518;
	wire [4-1:0] node1521;
	wire [4-1:0] node1522;
	wire [4-1:0] node1526;
	wire [4-1:0] node1527;
	wire [4-1:0] node1528;
	wire [4-1:0] node1529;
	wire [4-1:0] node1532;
	wire [4-1:0] node1535;
	wire [4-1:0] node1536;
	wire [4-1:0] node1539;
	wire [4-1:0] node1542;
	wire [4-1:0] node1543;
	wire [4-1:0] node1544;
	wire [4-1:0] node1547;
	wire [4-1:0] node1550;
	wire [4-1:0] node1552;
	wire [4-1:0] node1555;
	wire [4-1:0] node1556;
	wire [4-1:0] node1557;
	wire [4-1:0] node1558;
	wire [4-1:0] node1561;
	wire [4-1:0] node1563;
	wire [4-1:0] node1566;
	wire [4-1:0] node1568;
	wire [4-1:0] node1569;
	wire [4-1:0] node1572;
	wire [4-1:0] node1575;
	wire [4-1:0] node1576;
	wire [4-1:0] node1579;
	wire [4-1:0] node1581;
	wire [4-1:0] node1583;
	wire [4-1:0] node1586;
	wire [4-1:0] node1587;
	wire [4-1:0] node1588;
	wire [4-1:0] node1589;
	wire [4-1:0] node1590;
	wire [4-1:0] node1591;
	wire [4-1:0] node1593;
	wire [4-1:0] node1596;
	wire [4-1:0] node1597;
	wire [4-1:0] node1600;
	wire [4-1:0] node1604;
	wire [4-1:0] node1605;
	wire [4-1:0] node1606;
	wire [4-1:0] node1607;
	wire [4-1:0] node1610;
	wire [4-1:0] node1613;
	wire [4-1:0] node1614;
	wire [4-1:0] node1618;
	wire [4-1:0] node1619;
	wire [4-1:0] node1620;
	wire [4-1:0] node1625;
	wire [4-1:0] node1626;
	wire [4-1:0] node1627;
	wire [4-1:0] node1628;
	wire [4-1:0] node1631;
	wire [4-1:0] node1634;
	wire [4-1:0] node1636;
	wire [4-1:0] node1637;
	wire [4-1:0] node1640;
	wire [4-1:0] node1643;
	wire [4-1:0] node1644;
	wire [4-1:0] node1646;
	wire [4-1:0] node1649;
	wire [4-1:0] node1650;
	wire [4-1:0] node1651;
	wire [4-1:0] node1654;
	wire [4-1:0] node1658;
	wire [4-1:0] node1659;
	wire [4-1:0] node1660;
	wire [4-1:0] node1661;
	wire [4-1:0] node1663;
	wire [4-1:0] node1667;
	wire [4-1:0] node1668;
	wire [4-1:0] node1670;
	wire [4-1:0] node1671;
	wire [4-1:0] node1674;
	wire [4-1:0] node1677;
	wire [4-1:0] node1679;
	wire [4-1:0] node1680;
	wire [4-1:0] node1683;
	wire [4-1:0] node1686;
	wire [4-1:0] node1687;
	wire [4-1:0] node1688;
	wire [4-1:0] node1690;
	wire [4-1:0] node1693;
	wire [4-1:0] node1694;
	wire [4-1:0] node1697;
	wire [4-1:0] node1700;
	wire [4-1:0] node1701;
	wire [4-1:0] node1702;
	wire [4-1:0] node1706;
	wire [4-1:0] node1707;
	wire [4-1:0] node1708;
	wire [4-1:0] node1711;
	wire [4-1:0] node1715;
	wire [4-1:0] node1716;
	wire [4-1:0] node1717;
	wire [4-1:0] node1718;
	wire [4-1:0] node1719;
	wire [4-1:0] node1720;
	wire [4-1:0] node1721;
	wire [4-1:0] node1723;
	wire [4-1:0] node1727;
	wire [4-1:0] node1728;
	wire [4-1:0] node1730;
	wire [4-1:0] node1733;
	wire [4-1:0] node1734;
	wire [4-1:0] node1737;
	wire [4-1:0] node1740;
	wire [4-1:0] node1741;
	wire [4-1:0] node1743;
	wire [4-1:0] node1746;
	wire [4-1:0] node1748;
	wire [4-1:0] node1749;
	wire [4-1:0] node1752;
	wire [4-1:0] node1755;
	wire [4-1:0] node1756;
	wire [4-1:0] node1757;
	wire [4-1:0] node1758;
	wire [4-1:0] node1762;
	wire [4-1:0] node1764;
	wire [4-1:0] node1766;
	wire [4-1:0] node1769;
	wire [4-1:0] node1770;
	wire [4-1:0] node1772;
	wire [4-1:0] node1773;
	wire [4-1:0] node1776;
	wire [4-1:0] node1779;
	wire [4-1:0] node1780;
	wire [4-1:0] node1782;
	wire [4-1:0] node1785;
	wire [4-1:0] node1786;
	wire [4-1:0] node1790;
	wire [4-1:0] node1791;
	wire [4-1:0] node1792;
	wire [4-1:0] node1793;
	wire [4-1:0] node1797;
	wire [4-1:0] node1798;
	wire [4-1:0] node1799;
	wire [4-1:0] node1802;
	wire [4-1:0] node1805;
	wire [4-1:0] node1807;
	wire [4-1:0] node1810;
	wire [4-1:0] node1811;
	wire [4-1:0] node1812;
	wire [4-1:0] node1813;
	wire [4-1:0] node1816;
	wire [4-1:0] node1819;
	wire [4-1:0] node1820;
	wire [4-1:0] node1823;
	wire [4-1:0] node1824;
	wire [4-1:0] node1828;
	wire [4-1:0] node1829;
	wire [4-1:0] node1830;
	wire [4-1:0] node1833;
	wire [4-1:0] node1836;
	wire [4-1:0] node1837;
	wire [4-1:0] node1840;
	wire [4-1:0] node1843;
	wire [4-1:0] node1844;
	wire [4-1:0] node1845;
	wire [4-1:0] node1846;
	wire [4-1:0] node1847;
	wire [4-1:0] node1849;
	wire [4-1:0] node1852;
	wire [4-1:0] node1853;
	wire [4-1:0] node1857;
	wire [4-1:0] node1858;
	wire [4-1:0] node1859;
	wire [4-1:0] node1860;
	wire [4-1:0] node1863;
	wire [4-1:0] node1866;
	wire [4-1:0] node1867;
	wire [4-1:0] node1870;
	wire [4-1:0] node1873;
	wire [4-1:0] node1875;
	wire [4-1:0] node1878;
	wire [4-1:0] node1879;
	wire [4-1:0] node1880;
	wire [4-1:0] node1881;
	wire [4-1:0] node1885;
	wire [4-1:0] node1886;
	wire [4-1:0] node1889;
	wire [4-1:0] node1892;
	wire [4-1:0] node1893;
	wire [4-1:0] node1894;
	wire [4-1:0] node1897;
	wire [4-1:0] node1900;
	wire [4-1:0] node1901;
	wire [4-1:0] node1905;
	wire [4-1:0] node1906;
	wire [4-1:0] node1907;
	wire [4-1:0] node1908;
	wire [4-1:0] node1910;
	wire [4-1:0] node1913;
	wire [4-1:0] node1915;
	wire [4-1:0] node1918;
	wire [4-1:0] node1919;
	wire [4-1:0] node1920;
	wire [4-1:0] node1925;
	wire [4-1:0] node1926;
	wire [4-1:0] node1927;
	wire [4-1:0] node1928;
	wire [4-1:0] node1932;
	wire [4-1:0] node1933;
	wire [4-1:0] node1936;
	wire [4-1:0] node1939;
	wire [4-1:0] node1940;
	wire [4-1:0] node1943;
	wire [4-1:0] node1945;
	wire [4-1:0] node1948;
	wire [4-1:0] node1949;
	wire [4-1:0] node1950;
	wire [4-1:0] node1951;
	wire [4-1:0] node1952;
	wire [4-1:0] node1953;
	wire [4-1:0] node1954;
	wire [4-1:0] node1955;
	wire [4-1:0] node1956;
	wire [4-1:0] node1958;
	wire [4-1:0] node1961;
	wire [4-1:0] node1963;
	wire [4-1:0] node1966;
	wire [4-1:0] node1968;
	wire [4-1:0] node1970;
	wire [4-1:0] node1972;
	wire [4-1:0] node1975;
	wire [4-1:0] node1976;
	wire [4-1:0] node1977;
	wire [4-1:0] node1978;
	wire [4-1:0] node1981;
	wire [4-1:0] node1984;
	wire [4-1:0] node1986;
	wire [4-1:0] node1989;
	wire [4-1:0] node1990;
	wire [4-1:0] node1992;
	wire [4-1:0] node1994;
	wire [4-1:0] node1997;
	wire [4-1:0] node1998;
	wire [4-1:0] node1999;
	wire [4-1:0] node2002;
	wire [4-1:0] node2005;
	wire [4-1:0] node2007;
	wire [4-1:0] node2010;
	wire [4-1:0] node2011;
	wire [4-1:0] node2012;
	wire [4-1:0] node2013;
	wire [4-1:0] node2014;
	wire [4-1:0] node2015;
	wire [4-1:0] node2020;
	wire [4-1:0] node2021;
	wire [4-1:0] node2023;
	wire [4-1:0] node2026;
	wire [4-1:0] node2028;
	wire [4-1:0] node2031;
	wire [4-1:0] node2033;
	wire [4-1:0] node2034;
	wire [4-1:0] node2037;
	wire [4-1:0] node2040;
	wire [4-1:0] node2041;
	wire [4-1:0] node2042;
	wire [4-1:0] node2043;
	wire [4-1:0] node2047;
	wire [4-1:0] node2048;
	wire [4-1:0] node2051;
	wire [4-1:0] node2054;
	wire [4-1:0] node2055;
	wire [4-1:0] node2056;
	wire [4-1:0] node2058;
	wire [4-1:0] node2061;
	wire [4-1:0] node2064;
	wire [4-1:0] node2065;
	wire [4-1:0] node2066;
	wire [4-1:0] node2069;
	wire [4-1:0] node2072;
	wire [4-1:0] node2073;
	wire [4-1:0] node2076;
	wire [4-1:0] node2079;
	wire [4-1:0] node2080;
	wire [4-1:0] node2081;
	wire [4-1:0] node2082;
	wire [4-1:0] node2083;
	wire [4-1:0] node2086;
	wire [4-1:0] node2088;
	wire [4-1:0] node2091;
	wire [4-1:0] node2092;
	wire [4-1:0] node2093;
	wire [4-1:0] node2096;
	wire [4-1:0] node2100;
	wire [4-1:0] node2101;
	wire [4-1:0] node2102;
	wire [4-1:0] node2103;
	wire [4-1:0] node2106;
	wire [4-1:0] node2109;
	wire [4-1:0] node2111;
	wire [4-1:0] node2114;
	wire [4-1:0] node2115;
	wire [4-1:0] node2117;
	wire [4-1:0] node2120;
	wire [4-1:0] node2121;
	wire [4-1:0] node2122;
	wire [4-1:0] node2125;
	wire [4-1:0] node2128;
	wire [4-1:0] node2130;
	wire [4-1:0] node2133;
	wire [4-1:0] node2134;
	wire [4-1:0] node2135;
	wire [4-1:0] node2136;
	wire [4-1:0] node2137;
	wire [4-1:0] node2139;
	wire [4-1:0] node2142;
	wire [4-1:0] node2143;
	wire [4-1:0] node2146;
	wire [4-1:0] node2149;
	wire [4-1:0] node2152;
	wire [4-1:0] node2153;
	wire [4-1:0] node2154;
	wire [4-1:0] node2156;
	wire [4-1:0] node2159;
	wire [4-1:0] node2161;
	wire [4-1:0] node2164;
	wire [4-1:0] node2166;
	wire [4-1:0] node2169;
	wire [4-1:0] node2170;
	wire [4-1:0] node2171;
	wire [4-1:0] node2172;
	wire [4-1:0] node2173;
	wire [4-1:0] node2176;
	wire [4-1:0] node2179;
	wire [4-1:0] node2180;
	wire [4-1:0] node2183;
	wire [4-1:0] node2186;
	wire [4-1:0] node2188;
	wire [4-1:0] node2191;
	wire [4-1:0] node2192;
	wire [4-1:0] node2193;
	wire [4-1:0] node2195;
	wire [4-1:0] node2198;
	wire [4-1:0] node2199;
	wire [4-1:0] node2202;
	wire [4-1:0] node2205;
	wire [4-1:0] node2206;
	wire [4-1:0] node2209;
	wire [4-1:0] node2212;
	wire [4-1:0] node2213;
	wire [4-1:0] node2214;
	wire [4-1:0] node2215;
	wire [4-1:0] node2216;
	wire [4-1:0] node2219;
	wire [4-1:0] node2221;
	wire [4-1:0] node2224;
	wire [4-1:0] node2225;
	wire [4-1:0] node2226;
	wire [4-1:0] node2229;
	wire [4-1:0] node2232;
	wire [4-1:0] node2233;
	wire [4-1:0] node2234;
	wire [4-1:0] node2237;
	wire [4-1:0] node2240;
	wire [4-1:0] node2241;
	wire [4-1:0] node2244;
	wire [4-1:0] node2247;
	wire [4-1:0] node2248;
	wire [4-1:0] node2249;
	wire [4-1:0] node2252;
	wire [4-1:0] node2254;
	wire [4-1:0] node2257;
	wire [4-1:0] node2258;
	wire [4-1:0] node2259;
	wire [4-1:0] node2262;
	wire [4-1:0] node2265;
	wire [4-1:0] node2266;
	wire [4-1:0] node2267;
	wire [4-1:0] node2270;
	wire [4-1:0] node2273;
	wire [4-1:0] node2274;
	wire [4-1:0] node2278;
	wire [4-1:0] node2279;
	wire [4-1:0] node2280;
	wire [4-1:0] node2281;
	wire [4-1:0] node2284;
	wire [4-1:0] node2286;
	wire [4-1:0] node2289;
	wire [4-1:0] node2290;
	wire [4-1:0] node2291;
	wire [4-1:0] node2294;
	wire [4-1:0] node2297;
	wire [4-1:0] node2298;
	wire [4-1:0] node2301;
	wire [4-1:0] node2304;
	wire [4-1:0] node2305;
	wire [4-1:0] node2306;
	wire [4-1:0] node2309;
	wire [4-1:0] node2311;
	wire [4-1:0] node2314;
	wire [4-1:0] node2315;
	wire [4-1:0] node2316;
	wire [4-1:0] node2319;
	wire [4-1:0] node2322;
	wire [4-1:0] node2323;
	wire [4-1:0] node2325;
	wire [4-1:0] node2328;
	wire [4-1:0] node2329;
	wire [4-1:0] node2332;
	wire [4-1:0] node2335;
	wire [4-1:0] node2336;
	wire [4-1:0] node2337;
	wire [4-1:0] node2338;
	wire [4-1:0] node2339;
	wire [4-1:0] node2340;
	wire [4-1:0] node2341;
	wire [4-1:0] node2342;
	wire [4-1:0] node2344;
	wire [4-1:0] node2348;
	wire [4-1:0] node2349;
	wire [4-1:0] node2352;
	wire [4-1:0] node2355;
	wire [4-1:0] node2356;
	wire [4-1:0] node2357;
	wire [4-1:0] node2361;
	wire [4-1:0] node2362;
	wire [4-1:0] node2364;
	wire [4-1:0] node2368;
	wire [4-1:0] node2369;
	wire [4-1:0] node2370;
	wire [4-1:0] node2371;
	wire [4-1:0] node2375;
	wire [4-1:0] node2376;
	wire [4-1:0] node2378;
	wire [4-1:0] node2382;
	wire [4-1:0] node2383;
	wire [4-1:0] node2385;
	wire [4-1:0] node2386;
	wire [4-1:0] node2389;
	wire [4-1:0] node2392;
	wire [4-1:0] node2393;
	wire [4-1:0] node2396;
	wire [4-1:0] node2397;
	wire [4-1:0] node2401;
	wire [4-1:0] node2402;
	wire [4-1:0] node2403;
	wire [4-1:0] node2404;
	wire [4-1:0] node2407;
	wire [4-1:0] node2408;
	wire [4-1:0] node2412;
	wire [4-1:0] node2413;
	wire [4-1:0] node2415;
	wire [4-1:0] node2418;
	wire [4-1:0] node2419;
	wire [4-1:0] node2423;
	wire [4-1:0] node2424;
	wire [4-1:0] node2425;
	wire [4-1:0] node2428;
	wire [4-1:0] node2430;
	wire [4-1:0] node2433;
	wire [4-1:0] node2434;
	wire [4-1:0] node2435;
	wire [4-1:0] node2440;
	wire [4-1:0] node2441;
	wire [4-1:0] node2442;
	wire [4-1:0] node2443;
	wire [4-1:0] node2444;
	wire [4-1:0] node2445;
	wire [4-1:0] node2447;
	wire [4-1:0] node2450;
	wire [4-1:0] node2452;
	wire [4-1:0] node2455;
	wire [4-1:0] node2456;
	wire [4-1:0] node2460;
	wire [4-1:0] node2462;
	wire [4-1:0] node2463;
	wire [4-1:0] node2464;
	wire [4-1:0] node2469;
	wire [4-1:0] node2470;
	wire [4-1:0] node2472;
	wire [4-1:0] node2475;
	wire [4-1:0] node2476;
	wire [4-1:0] node2478;
	wire [4-1:0] node2479;
	wire [4-1:0] node2482;
	wire [4-1:0] node2485;
	wire [4-1:0] node2486;
	wire [4-1:0] node2490;
	wire [4-1:0] node2491;
	wire [4-1:0] node2492;
	wire [4-1:0] node2493;
	wire [4-1:0] node2494;
	wire [4-1:0] node2497;
	wire [4-1:0] node2500;
	wire [4-1:0] node2501;
	wire [4-1:0] node2502;
	wire [4-1:0] node2506;
	wire [4-1:0] node2509;
	wire [4-1:0] node2510;
	wire [4-1:0] node2511;
	wire [4-1:0] node2515;
	wire [4-1:0] node2517;
	wire [4-1:0] node2520;
	wire [4-1:0] node2521;
	wire [4-1:0] node2522;
	wire [4-1:0] node2523;
	wire [4-1:0] node2524;
	wire [4-1:0] node2529;
	wire [4-1:0] node2530;
	wire [4-1:0] node2533;
	wire [4-1:0] node2536;
	wire [4-1:0] node2537;
	wire [4-1:0] node2538;
	wire [4-1:0] node2539;
	wire [4-1:0] node2542;
	wire [4-1:0] node2546;
	wire [4-1:0] node2547;
	wire [4-1:0] node2548;
	wire [4-1:0] node2552;
	wire [4-1:0] node2553;
	wire [4-1:0] node2556;
	wire [4-1:0] node2559;
	wire [4-1:0] node2560;
	wire [4-1:0] node2561;
	wire [4-1:0] node2562;
	wire [4-1:0] node2563;
	wire [4-1:0] node2564;
	wire [4-1:0] node2567;
	wire [4-1:0] node2570;
	wire [4-1:0] node2572;
	wire [4-1:0] node2574;
	wire [4-1:0] node2575;
	wire [4-1:0] node2578;
	wire [4-1:0] node2581;
	wire [4-1:0] node2582;
	wire [4-1:0] node2584;
	wire [4-1:0] node2587;
	wire [4-1:0] node2588;
	wire [4-1:0] node2589;
	wire [4-1:0] node2592;
	wire [4-1:0] node2595;
	wire [4-1:0] node2596;
	wire [4-1:0] node2600;
	wire [4-1:0] node2601;
	wire [4-1:0] node2602;
	wire [4-1:0] node2603;
	wire [4-1:0] node2605;
	wire [4-1:0] node2606;
	wire [4-1:0] node2609;
	wire [4-1:0] node2612;
	wire [4-1:0] node2613;
	wire [4-1:0] node2614;
	wire [4-1:0] node2617;
	wire [4-1:0] node2620;
	wire [4-1:0] node2621;
	wire [4-1:0] node2624;
	wire [4-1:0] node2627;
	wire [4-1:0] node2628;
	wire [4-1:0] node2629;
	wire [4-1:0] node2632;
	wire [4-1:0] node2635;
	wire [4-1:0] node2636;
	wire [4-1:0] node2637;
	wire [4-1:0] node2640;
	wire [4-1:0] node2644;
	wire [4-1:0] node2645;
	wire [4-1:0] node2646;
	wire [4-1:0] node2647;
	wire [4-1:0] node2649;
	wire [4-1:0] node2652;
	wire [4-1:0] node2655;
	wire [4-1:0] node2656;
	wire [4-1:0] node2659;
	wire [4-1:0] node2662;
	wire [4-1:0] node2663;
	wire [4-1:0] node2664;
	wire [4-1:0] node2667;
	wire [4-1:0] node2670;
	wire [4-1:0] node2671;
	wire [4-1:0] node2674;
	wire [4-1:0] node2677;
	wire [4-1:0] node2678;
	wire [4-1:0] node2679;
	wire [4-1:0] node2680;
	wire [4-1:0] node2681;
	wire [4-1:0] node2682;
	wire [4-1:0] node2685;
	wire [4-1:0] node2688;
	wire [4-1:0] node2689;
	wire [4-1:0] node2692;
	wire [4-1:0] node2695;
	wire [4-1:0] node2696;
	wire [4-1:0] node2697;
	wire [4-1:0] node2700;
	wire [4-1:0] node2704;
	wire [4-1:0] node2705;
	wire [4-1:0] node2707;
	wire [4-1:0] node2709;
	wire [4-1:0] node2712;
	wire [4-1:0] node2713;
	wire [4-1:0] node2717;
	wire [4-1:0] node2718;
	wire [4-1:0] node2719;
	wire [4-1:0] node2720;
	wire [4-1:0] node2724;
	wire [4-1:0] node2725;
	wire [4-1:0] node2729;
	wire [4-1:0] node2730;
	wire [4-1:0] node2731;
	wire [4-1:0] node2735;
	wire [4-1:0] node2736;
	wire [4-1:0] node2740;
	wire [4-1:0] node2741;
	wire [4-1:0] node2742;
	wire [4-1:0] node2743;
	wire [4-1:0] node2744;
	wire [4-1:0] node2745;
	wire [4-1:0] node2746;
	wire [4-1:0] node2747;
	wire [4-1:0] node2750;
	wire [4-1:0] node2753;
	wire [4-1:0] node2754;
	wire [4-1:0] node2755;
	wire [4-1:0] node2756;
	wire [4-1:0] node2759;
	wire [4-1:0] node2762;
	wire [4-1:0] node2763;
	wire [4-1:0] node2767;
	wire [4-1:0] node2768;
	wire [4-1:0] node2769;
	wire [4-1:0] node2772;
	wire [4-1:0] node2776;
	wire [4-1:0] node2777;
	wire [4-1:0] node2778;
	wire [4-1:0] node2780;
	wire [4-1:0] node2783;
	wire [4-1:0] node2785;
	wire [4-1:0] node2788;
	wire [4-1:0] node2789;
	wire [4-1:0] node2792;
	wire [4-1:0] node2794;
	wire [4-1:0] node2797;
	wire [4-1:0] node2798;
	wire [4-1:0] node2799;
	wire [4-1:0] node2800;
	wire [4-1:0] node2802;
	wire [4-1:0] node2805;
	wire [4-1:0] node2808;
	wire [4-1:0] node2810;
	wire [4-1:0] node2812;
	wire [4-1:0] node2815;
	wire [4-1:0] node2816;
	wire [4-1:0] node2817;
	wire [4-1:0] node2819;
	wire [4-1:0] node2820;
	wire [4-1:0] node2825;
	wire [4-1:0] node2826;
	wire [4-1:0] node2827;
	wire [4-1:0] node2831;
	wire [4-1:0] node2832;
	wire [4-1:0] node2836;
	wire [4-1:0] node2837;
	wire [4-1:0] node2838;
	wire [4-1:0] node2839;
	wire [4-1:0] node2840;
	wire [4-1:0] node2843;
	wire [4-1:0] node2846;
	wire [4-1:0] node2847;
	wire [4-1:0] node2848;
	wire [4-1:0] node2852;
	wire [4-1:0] node2853;
	wire [4-1:0] node2856;
	wire [4-1:0] node2859;
	wire [4-1:0] node2860;
	wire [4-1:0] node2861;
	wire [4-1:0] node2862;
	wire [4-1:0] node2865;
	wire [4-1:0] node2868;
	wire [4-1:0] node2870;
	wire [4-1:0] node2873;
	wire [4-1:0] node2875;
	wire [4-1:0] node2877;
	wire [4-1:0] node2880;
	wire [4-1:0] node2881;
	wire [4-1:0] node2882;
	wire [4-1:0] node2883;
	wire [4-1:0] node2884;
	wire [4-1:0] node2885;
	wire [4-1:0] node2888;
	wire [4-1:0] node2892;
	wire [4-1:0] node2893;
	wire [4-1:0] node2896;
	wire [4-1:0] node2899;
	wire [4-1:0] node2900;
	wire [4-1:0] node2902;
	wire [4-1:0] node2904;
	wire [4-1:0] node2907;
	wire [4-1:0] node2908;
	wire [4-1:0] node2912;
	wire [4-1:0] node2913;
	wire [4-1:0] node2914;
	wire [4-1:0] node2916;
	wire [4-1:0] node2919;
	wire [4-1:0] node2921;
	wire [4-1:0] node2924;
	wire [4-1:0] node2926;
	wire [4-1:0] node2929;
	wire [4-1:0] node2930;
	wire [4-1:0] node2931;
	wire [4-1:0] node2932;
	wire [4-1:0] node2933;
	wire [4-1:0] node2936;
	wire [4-1:0] node2937;
	wire [4-1:0] node2941;
	wire [4-1:0] node2942;
	wire [4-1:0] node2943;
	wire [4-1:0] node2944;
	wire [4-1:0] node2945;
	wire [4-1:0] node2949;
	wire [4-1:0] node2950;
	wire [4-1:0] node2953;
	wire [4-1:0] node2956;
	wire [4-1:0] node2957;
	wire [4-1:0] node2960;
	wire [4-1:0] node2963;
	wire [4-1:0] node2964;
	wire [4-1:0] node2967;
	wire [4-1:0] node2970;
	wire [4-1:0] node2971;
	wire [4-1:0] node2972;
	wire [4-1:0] node2973;
	wire [4-1:0] node2974;
	wire [4-1:0] node2977;
	wire [4-1:0] node2980;
	wire [4-1:0] node2981;
	wire [4-1:0] node2985;
	wire [4-1:0] node2987;
	wire [4-1:0] node2990;
	wire [4-1:0] node2991;
	wire [4-1:0] node2994;
	wire [4-1:0] node2997;
	wire [4-1:0] node2998;
	wire [4-1:0] node2999;
	wire [4-1:0] node3000;
	wire [4-1:0] node3001;
	wire [4-1:0] node3004;
	wire [4-1:0] node3007;
	wire [4-1:0] node3008;
	wire [4-1:0] node3011;
	wire [4-1:0] node3014;
	wire [4-1:0] node3015;
	wire [4-1:0] node3017;
	wire [4-1:0] node3018;
	wire [4-1:0] node3021;
	wire [4-1:0] node3024;
	wire [4-1:0] node3025;
	wire [4-1:0] node3028;
	wire [4-1:0] node3031;
	wire [4-1:0] node3032;
	wire [4-1:0] node3033;
	wire [4-1:0] node3034;
	wire [4-1:0] node3037;
	wire [4-1:0] node3040;
	wire [4-1:0] node3041;
	wire [4-1:0] node3044;
	wire [4-1:0] node3047;
	wire [4-1:0] node3048;
	wire [4-1:0] node3049;
	wire [4-1:0] node3050;
	wire [4-1:0] node3051;
	wire [4-1:0] node3054;
	wire [4-1:0] node3057;
	wire [4-1:0] node3058;
	wire [4-1:0] node3062;
	wire [4-1:0] node3063;
	wire [4-1:0] node3066;
	wire [4-1:0] node3069;
	wire [4-1:0] node3070;
	wire [4-1:0] node3073;
	wire [4-1:0] node3076;
	wire [4-1:0] node3077;
	wire [4-1:0] node3078;
	wire [4-1:0] node3079;
	wire [4-1:0] node3080;
	wire [4-1:0] node3081;
	wire [4-1:0] node3082;
	wire [4-1:0] node3084;
	wire [4-1:0] node3087;
	wire [4-1:0] node3089;
	wire [4-1:0] node3092;
	wire [4-1:0] node3093;
	wire [4-1:0] node3096;
	wire [4-1:0] node3097;
	wire [4-1:0] node3099;
	wire [4-1:0] node3103;
	wire [4-1:0] node3104;
	wire [4-1:0] node3107;
	wire [4-1:0] node3108;
	wire [4-1:0] node3110;
	wire [4-1:0] node3113;
	wire [4-1:0] node3115;
	wire [4-1:0] node3118;
	wire [4-1:0] node3119;
	wire [4-1:0] node3120;
	wire [4-1:0] node3121;
	wire [4-1:0] node3124;
	wire [4-1:0] node3127;
	wire [4-1:0] node3128;
	wire [4-1:0] node3129;
	wire [4-1:0] node3132;
	wire [4-1:0] node3133;
	wire [4-1:0] node3138;
	wire [4-1:0] node3139;
	wire [4-1:0] node3140;
	wire [4-1:0] node3142;
	wire [4-1:0] node3143;
	wire [4-1:0] node3147;
	wire [4-1:0] node3148;
	wire [4-1:0] node3152;
	wire [4-1:0] node3153;
	wire [4-1:0] node3154;
	wire [4-1:0] node3155;
	wire [4-1:0] node3158;
	wire [4-1:0] node3161;
	wire [4-1:0] node3162;
	wire [4-1:0] node3166;
	wire [4-1:0] node3167;
	wire [4-1:0] node3168;
	wire [4-1:0] node3171;
	wire [4-1:0] node3175;
	wire [4-1:0] node3176;
	wire [4-1:0] node3177;
	wire [4-1:0] node3178;
	wire [4-1:0] node3179;
	wire [4-1:0] node3181;
	wire [4-1:0] node3184;
	wire [4-1:0] node3186;
	wire [4-1:0] node3189;
	wire [4-1:0] node3190;
	wire [4-1:0] node3193;
	wire [4-1:0] node3195;
	wire [4-1:0] node3198;
	wire [4-1:0] node3199;
	wire [4-1:0] node3200;
	wire [4-1:0] node3202;
	wire [4-1:0] node3205;
	wire [4-1:0] node3206;
	wire [4-1:0] node3210;
	wire [4-1:0] node3211;
	wire [4-1:0] node3212;
	wire [4-1:0] node3216;
	wire [4-1:0] node3217;
	wire [4-1:0] node3221;
	wire [4-1:0] node3222;
	wire [4-1:0] node3223;
	wire [4-1:0] node3224;
	wire [4-1:0] node3228;
	wire [4-1:0] node3230;
	wire [4-1:0] node3231;
	wire [4-1:0] node3234;
	wire [4-1:0] node3237;
	wire [4-1:0] node3238;
	wire [4-1:0] node3239;
	wire [4-1:0] node3241;
	wire [4-1:0] node3244;
	wire [4-1:0] node3245;
	wire [4-1:0] node3248;
	wire [4-1:0] node3251;
	wire [4-1:0] node3252;
	wire [4-1:0] node3253;
	wire [4-1:0] node3256;
	wire [4-1:0] node3259;
	wire [4-1:0] node3260;
	wire [4-1:0] node3264;
	wire [4-1:0] node3265;
	wire [4-1:0] node3266;
	wire [4-1:0] node3267;
	wire [4-1:0] node3268;
	wire [4-1:0] node3271;
	wire [4-1:0] node3273;
	wire [4-1:0] node3276;
	wire [4-1:0] node3277;
	wire [4-1:0] node3280;
	wire [4-1:0] node3282;
	wire [4-1:0] node3285;
	wire [4-1:0] node3286;
	wire [4-1:0] node3287;
	wire [4-1:0] node3288;
	wire [4-1:0] node3291;
	wire [4-1:0] node3294;
	wire [4-1:0] node3296;
	wire [4-1:0] node3299;
	wire [4-1:0] node3300;
	wire [4-1:0] node3303;
	wire [4-1:0] node3305;
	wire [4-1:0] node3308;
	wire [4-1:0] node3309;
	wire [4-1:0] node3310;
	wire [4-1:0] node3311;
	wire [4-1:0] node3313;
	wire [4-1:0] node3314;
	wire [4-1:0] node3317;
	wire [4-1:0] node3320;
	wire [4-1:0] node3321;
	wire [4-1:0] node3323;
	wire [4-1:0] node3324;
	wire [4-1:0] node3328;
	wire [4-1:0] node3329;
	wire [4-1:0] node3330;
	wire [4-1:0] node3333;
	wire [4-1:0] node3337;
	wire [4-1:0] node3338;
	wire [4-1:0] node3339;
	wire [4-1:0] node3340;
	wire [4-1:0] node3344;
	wire [4-1:0] node3346;
	wire [4-1:0] node3348;
	wire [4-1:0] node3351;
	wire [4-1:0] node3352;
	wire [4-1:0] node3355;
	wire [4-1:0] node3358;
	wire [4-1:0] node3359;
	wire [4-1:0] node3360;
	wire [4-1:0] node3361;
	wire [4-1:0] node3362;
	wire [4-1:0] node3363;
	wire [4-1:0] node3366;
	wire [4-1:0] node3369;
	wire [4-1:0] node3371;
	wire [4-1:0] node3374;
	wire [4-1:0] node3375;
	wire [4-1:0] node3376;
	wire [4-1:0] node3379;
	wire [4-1:0] node3382;
	wire [4-1:0] node3383;
	wire [4-1:0] node3386;
	wire [4-1:0] node3389;
	wire [4-1:0] node3390;
	wire [4-1:0] node3392;
	wire [4-1:0] node3395;
	wire [4-1:0] node3397;
	wire [4-1:0] node3400;
	wire [4-1:0] node3401;
	wire [4-1:0] node3402;
	wire [4-1:0] node3403;
	wire [4-1:0] node3405;
	wire [4-1:0] node3409;
	wire [4-1:0] node3410;
	wire [4-1:0] node3412;
	wire [4-1:0] node3415;
	wire [4-1:0] node3416;
	wire [4-1:0] node3420;
	wire [4-1:0] node3421;
	wire [4-1:0] node3424;
	wire [4-1:0] node3427;
	wire [4-1:0] node3428;
	wire [4-1:0] node3429;
	wire [4-1:0] node3430;
	wire [4-1:0] node3431;
	wire [4-1:0] node3432;
	wire [4-1:0] node3433;
	wire [4-1:0] node3434;
	wire [4-1:0] node3435;
	wire [4-1:0] node3436;
	wire [4-1:0] node3439;
	wire [4-1:0] node3442;
	wire [4-1:0] node3443;
	wire [4-1:0] node3444;
	wire [4-1:0] node3445;
	wire [4-1:0] node3448;
	wire [4-1:0] node3452;
	wire [4-1:0] node3453;
	wire [4-1:0] node3456;
	wire [4-1:0] node3459;
	wire [4-1:0] node3460;
	wire [4-1:0] node3462;
	wire [4-1:0] node3465;
	wire [4-1:0] node3467;
	wire [4-1:0] node3468;
	wire [4-1:0] node3471;
	wire [4-1:0] node3474;
	wire [4-1:0] node3475;
	wire [4-1:0] node3476;
	wire [4-1:0] node3477;
	wire [4-1:0] node3479;
	wire [4-1:0] node3482;
	wire [4-1:0] node3484;
	wire [4-1:0] node3485;
	wire [4-1:0] node3489;
	wire [4-1:0] node3490;
	wire [4-1:0] node3491;
	wire [4-1:0] node3495;
	wire [4-1:0] node3496;
	wire [4-1:0] node3500;
	wire [4-1:0] node3501;
	wire [4-1:0] node3502;
	wire [4-1:0] node3503;
	wire [4-1:0] node3506;
	wire [4-1:0] node3509;
	wire [4-1:0] node3510;
	wire [4-1:0] node3513;
	wire [4-1:0] node3516;
	wire [4-1:0] node3517;
	wire [4-1:0] node3518;
	wire [4-1:0] node3522;
	wire [4-1:0] node3523;
	wire [4-1:0] node3524;
	wire [4-1:0] node3528;
	wire [4-1:0] node3529;
	wire [4-1:0] node3533;
	wire [4-1:0] node3534;
	wire [4-1:0] node3535;
	wire [4-1:0] node3536;
	wire [4-1:0] node3537;
	wire [4-1:0] node3538;
	wire [4-1:0] node3540;
	wire [4-1:0] node3543;
	wire [4-1:0] node3544;
	wire [4-1:0] node3547;
	wire [4-1:0] node3550;
	wire [4-1:0] node3551;
	wire [4-1:0] node3554;
	wire [4-1:0] node3557;
	wire [4-1:0] node3558;
	wire [4-1:0] node3559;
	wire [4-1:0] node3562;
	wire [4-1:0] node3564;
	wire [4-1:0] node3567;
	wire [4-1:0] node3568;
	wire [4-1:0] node3571;
	wire [4-1:0] node3573;
	wire [4-1:0] node3576;
	wire [4-1:0] node3577;
	wire [4-1:0] node3578;
	wire [4-1:0] node3579;
	wire [4-1:0] node3583;
	wire [4-1:0] node3584;
	wire [4-1:0] node3585;
	wire [4-1:0] node3588;
	wire [4-1:0] node3591;
	wire [4-1:0] node3594;
	wire [4-1:0] node3595;
	wire [4-1:0] node3597;
	wire [4-1:0] node3600;
	wire [4-1:0] node3601;
	wire [4-1:0] node3602;
	wire [4-1:0] node3606;
	wire [4-1:0] node3609;
	wire [4-1:0] node3610;
	wire [4-1:0] node3611;
	wire [4-1:0] node3612;
	wire [4-1:0] node3613;
	wire [4-1:0] node3615;
	wire [4-1:0] node3619;
	wire [4-1:0] node3620;
	wire [4-1:0] node3622;
	wire [4-1:0] node3626;
	wire [4-1:0] node3627;
	wire [4-1:0] node3628;
	wire [4-1:0] node3629;
	wire [4-1:0] node3632;
	wire [4-1:0] node3636;
	wire [4-1:0] node3637;
	wire [4-1:0] node3641;
	wire [4-1:0] node3642;
	wire [4-1:0] node3643;
	wire [4-1:0] node3645;
	wire [4-1:0] node3648;
	wire [4-1:0] node3650;
	wire [4-1:0] node3652;
	wire [4-1:0] node3655;
	wire [4-1:0] node3656;
	wire [4-1:0] node3657;
	wire [4-1:0] node3661;
	wire [4-1:0] node3662;
	wire [4-1:0] node3663;
	wire [4-1:0] node3667;
	wire [4-1:0] node3670;
	wire [4-1:0] node3671;
	wire [4-1:0] node3672;
	wire [4-1:0] node3673;
	wire [4-1:0] node3674;
	wire [4-1:0] node3675;
	wire [4-1:0] node3677;
	wire [4-1:0] node3681;
	wire [4-1:0] node3682;
	wire [4-1:0] node3684;
	wire [4-1:0] node3687;
	wire [4-1:0] node3690;
	wire [4-1:0] node3691;
	wire [4-1:0] node3692;
	wire [4-1:0] node3695;
	wire [4-1:0] node3698;
	wire [4-1:0] node3699;
	wire [4-1:0] node3701;
	wire [4-1:0] node3702;
	wire [4-1:0] node3705;
	wire [4-1:0] node3708;
	wire [4-1:0] node3709;
	wire [4-1:0] node3712;
	wire [4-1:0] node3715;
	wire [4-1:0] node3716;
	wire [4-1:0] node3717;
	wire [4-1:0] node3718;
	wire [4-1:0] node3719;
	wire [4-1:0] node3721;
	wire [4-1:0] node3724;
	wire [4-1:0] node3727;
	wire [4-1:0] node3729;
	wire [4-1:0] node3731;
	wire [4-1:0] node3734;
	wire [4-1:0] node3735;
	wire [4-1:0] node3736;
	wire [4-1:0] node3739;
	wire [4-1:0] node3740;
	wire [4-1:0] node3744;
	wire [4-1:0] node3747;
	wire [4-1:0] node3748;
	wire [4-1:0] node3749;
	wire [4-1:0] node3750;
	wire [4-1:0] node3753;
	wire [4-1:0] node3756;
	wire [4-1:0] node3757;
	wire [4-1:0] node3760;
	wire [4-1:0] node3763;
	wire [4-1:0] node3764;
	wire [4-1:0] node3765;
	wire [4-1:0] node3768;
	wire [4-1:0] node3771;
	wire [4-1:0] node3772;
	wire [4-1:0] node3775;
	wire [4-1:0] node3778;
	wire [4-1:0] node3779;
	wire [4-1:0] node3780;
	wire [4-1:0] node3781;
	wire [4-1:0] node3782;
	wire [4-1:0] node3785;
	wire [4-1:0] node3788;
	wire [4-1:0] node3790;
	wire [4-1:0] node3791;
	wire [4-1:0] node3794;
	wire [4-1:0] node3797;
	wire [4-1:0] node3798;
	wire [4-1:0] node3799;
	wire [4-1:0] node3802;
	wire [4-1:0] node3804;
	wire [4-1:0] node3807;
	wire [4-1:0] node3808;
	wire [4-1:0] node3811;
	wire [4-1:0] node3813;
	wire [4-1:0] node3816;
	wire [4-1:0] node3817;
	wire [4-1:0] node3818;
	wire [4-1:0] node3819;
	wire [4-1:0] node3820;
	wire [4-1:0] node3824;
	wire [4-1:0] node3826;
	wire [4-1:0] node3829;
	wire [4-1:0] node3830;
	wire [4-1:0] node3831;
	wire [4-1:0] node3835;
	wire [4-1:0] node3837;
	wire [4-1:0] node3838;
	wire [4-1:0] node3841;
	wire [4-1:0] node3844;
	wire [4-1:0] node3845;
	wire [4-1:0] node3846;
	wire [4-1:0] node3848;
	wire [4-1:0] node3849;
	wire [4-1:0] node3853;
	wire [4-1:0] node3856;
	wire [4-1:0] node3857;
	wire [4-1:0] node3859;
	wire [4-1:0] node3860;
	wire [4-1:0] node3864;
	wire [4-1:0] node3865;
	wire [4-1:0] node3867;
	wire [4-1:0] node3870;
	wire [4-1:0] node3873;
	wire [4-1:0] node3874;
	wire [4-1:0] node3875;
	wire [4-1:0] node3876;
	wire [4-1:0] node3877;
	wire [4-1:0] node3878;
	wire [4-1:0] node3879;
	wire [4-1:0] node3882;
	wire [4-1:0] node3884;
	wire [4-1:0] node3887;
	wire [4-1:0] node3888;
	wire [4-1:0] node3890;
	wire [4-1:0] node3893;
	wire [4-1:0] node3895;
	wire [4-1:0] node3898;
	wire [4-1:0] node3899;
	wire [4-1:0] node3900;
	wire [4-1:0] node3903;
	wire [4-1:0] node3906;
	wire [4-1:0] node3907;
	wire [4-1:0] node3908;
	wire [4-1:0] node3911;
	wire [4-1:0] node3914;
	wire [4-1:0] node3915;
	wire [4-1:0] node3918;
	wire [4-1:0] node3921;
	wire [4-1:0] node3922;
	wire [4-1:0] node3923;
	wire [4-1:0] node3924;
	wire [4-1:0] node3925;
	wire [4-1:0] node3926;
	wire [4-1:0] node3929;
	wire [4-1:0] node3932;
	wire [4-1:0] node3933;
	wire [4-1:0] node3937;
	wire [4-1:0] node3938;
	wire [4-1:0] node3941;
	wire [4-1:0] node3944;
	wire [4-1:0] node3945;
	wire [4-1:0] node3946;
	wire [4-1:0] node3949;
	wire [4-1:0] node3952;
	wire [4-1:0] node3953;
	wire [4-1:0] node3957;
	wire [4-1:0] node3958;
	wire [4-1:0] node3959;
	wire [4-1:0] node3962;
	wire [4-1:0] node3964;
	wire [4-1:0] node3967;
	wire [4-1:0] node3968;
	wire [4-1:0] node3970;
	wire [4-1:0] node3973;
	wire [4-1:0] node3974;
	wire [4-1:0] node3977;
	wire [4-1:0] node3980;
	wire [4-1:0] node3981;
	wire [4-1:0] node3982;
	wire [4-1:0] node3983;
	wire [4-1:0] node3984;
	wire [4-1:0] node3987;
	wire [4-1:0] node3989;
	wire [4-1:0] node3991;
	wire [4-1:0] node3994;
	wire [4-1:0] node3995;
	wire [4-1:0] node3996;
	wire [4-1:0] node3997;
	wire [4-1:0] node4001;
	wire [4-1:0] node4004;
	wire [4-1:0] node4006;
	wire [4-1:0] node4007;
	wire [4-1:0] node4011;
	wire [4-1:0] node4012;
	wire [4-1:0] node4013;
	wire [4-1:0] node4015;
	wire [4-1:0] node4018;
	wire [4-1:0] node4019;
	wire [4-1:0] node4022;
	wire [4-1:0] node4025;
	wire [4-1:0] node4026;
	wire [4-1:0] node4028;
	wire [4-1:0] node4029;
	wire [4-1:0] node4032;
	wire [4-1:0] node4035;
	wire [4-1:0] node4036;
	wire [4-1:0] node4040;
	wire [4-1:0] node4041;
	wire [4-1:0] node4042;
	wire [4-1:0] node4043;
	wire [4-1:0] node4044;
	wire [4-1:0] node4048;
	wire [4-1:0] node4049;
	wire [4-1:0] node4052;
	wire [4-1:0] node4055;
	wire [4-1:0] node4057;
	wire [4-1:0] node4058;
	wire [4-1:0] node4060;
	wire [4-1:0] node4063;
	wire [4-1:0] node4066;
	wire [4-1:0] node4067;
	wire [4-1:0] node4068;
	wire [4-1:0] node4069;
	wire [4-1:0] node4071;
	wire [4-1:0] node4074;
	wire [4-1:0] node4076;
	wire [4-1:0] node4079;
	wire [4-1:0] node4081;
	wire [4-1:0] node4083;
	wire [4-1:0] node4086;
	wire [4-1:0] node4087;
	wire [4-1:0] node4089;
	wire [4-1:0] node4090;
	wire [4-1:0] node4093;
	wire [4-1:0] node4096;
	wire [4-1:0] node4097;
	wire [4-1:0] node4100;
	wire [4-1:0] node4103;
	wire [4-1:0] node4104;
	wire [4-1:0] node4105;
	wire [4-1:0] node4106;
	wire [4-1:0] node4107;
	wire [4-1:0] node4109;
	wire [4-1:0] node4112;
	wire [4-1:0] node4114;
	wire [4-1:0] node4117;
	wire [4-1:0] node4118;
	wire [4-1:0] node4120;
	wire [4-1:0] node4123;
	wire [4-1:0] node4125;
	wire [4-1:0] node4128;
	wire [4-1:0] node4129;
	wire [4-1:0] node4131;
	wire [4-1:0] node4132;
	wire [4-1:0] node4135;
	wire [4-1:0] node4137;
	wire [4-1:0] node4140;
	wire [4-1:0] node4141;
	wire [4-1:0] node4143;
	wire [4-1:0] node4145;
	wire [4-1:0] node4148;
	wire [4-1:0] node4149;
	wire [4-1:0] node4152;
	wire [4-1:0] node4154;
	wire [4-1:0] node4157;
	wire [4-1:0] node4158;
	wire [4-1:0] node4159;
	wire [4-1:0] node4160;
	wire [4-1:0] node4162;
	wire [4-1:0] node4165;
	wire [4-1:0] node4167;
	wire [4-1:0] node4170;
	wire [4-1:0] node4171;
	wire [4-1:0] node4173;
	wire [4-1:0] node4176;
	wire [4-1:0] node4178;
	wire [4-1:0] node4181;
	wire [4-1:0] node4182;
	wire [4-1:0] node4183;
	wire [4-1:0] node4184;
	wire [4-1:0] node4188;
	wire [4-1:0] node4189;
	wire [4-1:0] node4193;
	wire [4-1:0] node4194;
	wire [4-1:0] node4195;
	wire [4-1:0] node4199;
	wire [4-1:0] node4200;
	wire [4-1:0] node4204;
	wire [4-1:0] node4205;
	wire [4-1:0] node4206;
	wire [4-1:0] node4207;
	wire [4-1:0] node4208;
	wire [4-1:0] node4209;
	wire [4-1:0] node4210;
	wire [4-1:0] node4211;
	wire [4-1:0] node4212;
	wire [4-1:0] node4216;
	wire [4-1:0] node4217;
	wire [4-1:0] node4220;
	wire [4-1:0] node4223;
	wire [4-1:0] node4224;
	wire [4-1:0] node4225;
	wire [4-1:0] node4226;
	wire [4-1:0] node4231;
	wire [4-1:0] node4232;
	wire [4-1:0] node4234;
	wire [4-1:0] node4237;
	wire [4-1:0] node4239;
	wire [4-1:0] node4242;
	wire [4-1:0] node4243;
	wire [4-1:0] node4244;
	wire [4-1:0] node4246;
	wire [4-1:0] node4249;
	wire [4-1:0] node4251;
	wire [4-1:0] node4254;
	wire [4-1:0] node4255;
	wire [4-1:0] node4257;
	wire [4-1:0] node4260;
	wire [4-1:0] node4261;
	wire [4-1:0] node4262;
	wire [4-1:0] node4265;
	wire [4-1:0] node4268;
	wire [4-1:0] node4269;
	wire [4-1:0] node4272;
	wire [4-1:0] node4275;
	wire [4-1:0] node4276;
	wire [4-1:0] node4277;
	wire [4-1:0] node4278;
	wire [4-1:0] node4279;
	wire [4-1:0] node4280;
	wire [4-1:0] node4285;
	wire [4-1:0] node4286;
	wire [4-1:0] node4287;
	wire [4-1:0] node4290;
	wire [4-1:0] node4293;
	wire [4-1:0] node4294;
	wire [4-1:0] node4297;
	wire [4-1:0] node4300;
	wire [4-1:0] node4301;
	wire [4-1:0] node4302;
	wire [4-1:0] node4303;
	wire [4-1:0] node4306;
	wire [4-1:0] node4310;
	wire [4-1:0] node4312;
	wire [4-1:0] node4315;
	wire [4-1:0] node4316;
	wire [4-1:0] node4317;
	wire [4-1:0] node4320;
	wire [4-1:0] node4321;
	wire [4-1:0] node4322;
	wire [4-1:0] node4325;
	wire [4-1:0] node4328;
	wire [4-1:0] node4329;
	wire [4-1:0] node4332;
	wire [4-1:0] node4335;
	wire [4-1:0] node4336;
	wire [4-1:0] node4339;
	wire [4-1:0] node4340;
	wire [4-1:0] node4343;
	wire [4-1:0] node4345;
	wire [4-1:0] node4348;
	wire [4-1:0] node4349;
	wire [4-1:0] node4350;
	wire [4-1:0] node4351;
	wire [4-1:0] node4352;
	wire [4-1:0] node4353;
	wire [4-1:0] node4356;
	wire [4-1:0] node4359;
	wire [4-1:0] node4360;
	wire [4-1:0] node4363;
	wire [4-1:0] node4366;
	wire [4-1:0] node4367;
	wire [4-1:0] node4368;
	wire [4-1:0] node4372;
	wire [4-1:0] node4373;
	wire [4-1:0] node4376;
	wire [4-1:0] node4379;
	wire [4-1:0] node4380;
	wire [4-1:0] node4381;
	wire [4-1:0] node4383;
	wire [4-1:0] node4384;
	wire [4-1:0] node4388;
	wire [4-1:0] node4389;
	wire [4-1:0] node4392;
	wire [4-1:0] node4395;
	wire [4-1:0] node4397;
	wire [4-1:0] node4398;
	wire [4-1:0] node4399;
	wire [4-1:0] node4404;
	wire [4-1:0] node4405;
	wire [4-1:0] node4406;
	wire [4-1:0] node4407;
	wire [4-1:0] node4408;
	wire [4-1:0] node4411;
	wire [4-1:0] node4414;
	wire [4-1:0] node4415;
	wire [4-1:0] node4419;
	wire [4-1:0] node4420;
	wire [4-1:0] node4423;
	wire [4-1:0] node4424;
	wire [4-1:0] node4428;
	wire [4-1:0] node4429;
	wire [4-1:0] node4430;
	wire [4-1:0] node4431;
	wire [4-1:0] node4432;
	wire [4-1:0] node4436;
	wire [4-1:0] node4438;
	wire [4-1:0] node4441;
	wire [4-1:0] node4442;
	wire [4-1:0] node4443;
	wire [4-1:0] node4446;
	wire [4-1:0] node4449;
	wire [4-1:0] node4450;
	wire [4-1:0] node4454;
	wire [4-1:0] node4455;
	wire [4-1:0] node4456;
	wire [4-1:0] node4459;
	wire [4-1:0] node4460;
	wire [4-1:0] node4464;
	wire [4-1:0] node4465;
	wire [4-1:0] node4468;
	wire [4-1:0] node4470;
	wire [4-1:0] node4473;
	wire [4-1:0] node4474;
	wire [4-1:0] node4475;
	wire [4-1:0] node4476;
	wire [4-1:0] node4477;
	wire [4-1:0] node4478;
	wire [4-1:0] node4479;
	wire [4-1:0] node4482;
	wire [4-1:0] node4485;
	wire [4-1:0] node4486;
	wire [4-1:0] node4489;
	wire [4-1:0] node4492;
	wire [4-1:0] node4493;
	wire [4-1:0] node4494;
	wire [4-1:0] node4497;
	wire [4-1:0] node4501;
	wire [4-1:0] node4502;
	wire [4-1:0] node4503;
	wire [4-1:0] node4504;
	wire [4-1:0] node4505;
	wire [4-1:0] node4509;
	wire [4-1:0] node4511;
	wire [4-1:0] node4514;
	wire [4-1:0] node4515;
	wire [4-1:0] node4518;
	wire [4-1:0] node4521;
	wire [4-1:0] node4522;
	wire [4-1:0] node4523;
	wire [4-1:0] node4524;
	wire [4-1:0] node4528;
	wire [4-1:0] node4529;
	wire [4-1:0] node4532;
	wire [4-1:0] node4535;
	wire [4-1:0] node4536;
	wire [4-1:0] node4537;
	wire [4-1:0] node4540;
	wire [4-1:0] node4543;
	wire [4-1:0] node4544;
	wire [4-1:0] node4547;
	wire [4-1:0] node4550;
	wire [4-1:0] node4551;
	wire [4-1:0] node4552;
	wire [4-1:0] node4553;
	wire [4-1:0] node4554;
	wire [4-1:0] node4556;
	wire [4-1:0] node4560;
	wire [4-1:0] node4561;
	wire [4-1:0] node4563;
	wire [4-1:0] node4566;
	wire [4-1:0] node4568;
	wire [4-1:0] node4571;
	wire [4-1:0] node4572;
	wire [4-1:0] node4573;
	wire [4-1:0] node4577;
	wire [4-1:0] node4578;
	wire [4-1:0] node4580;
	wire [4-1:0] node4584;
	wire [4-1:0] node4585;
	wire [4-1:0] node4586;
	wire [4-1:0] node4587;
	wire [4-1:0] node4592;
	wire [4-1:0] node4593;
	wire [4-1:0] node4594;
	wire [4-1:0] node4598;
	wire [4-1:0] node4599;
	wire [4-1:0] node4603;
	wire [4-1:0] node4604;
	wire [4-1:0] node4605;
	wire [4-1:0] node4606;
	wire [4-1:0] node4607;
	wire [4-1:0] node4608;
	wire [4-1:0] node4610;
	wire [4-1:0] node4613;
	wire [4-1:0] node4614;
	wire [4-1:0] node4617;
	wire [4-1:0] node4620;
	wire [4-1:0] node4621;
	wire [4-1:0] node4624;
	wire [4-1:0] node4627;
	wire [4-1:0] node4628;
	wire [4-1:0] node4630;
	wire [4-1:0] node4631;
	wire [4-1:0] node4634;
	wire [4-1:0] node4637;
	wire [4-1:0] node4638;
	wire [4-1:0] node4639;
	wire [4-1:0] node4642;
	wire [4-1:0] node4646;
	wire [4-1:0] node4647;
	wire [4-1:0] node4648;
	wire [4-1:0] node4649;
	wire [4-1:0] node4650;
	wire [4-1:0] node4653;
	wire [4-1:0] node4657;
	wire [4-1:0] node4658;
	wire [4-1:0] node4659;
	wire [4-1:0] node4663;
	wire [4-1:0] node4664;
	wire [4-1:0] node4667;
	wire [4-1:0] node4670;
	wire [4-1:0] node4671;
	wire [4-1:0] node4673;
	wire [4-1:0] node4675;
	wire [4-1:0] node4678;
	wire [4-1:0] node4679;
	wire [4-1:0] node4680;
	wire [4-1:0] node4683;
	wire [4-1:0] node4687;
	wire [4-1:0] node4688;
	wire [4-1:0] node4689;
	wire [4-1:0] node4690;
	wire [4-1:0] node4693;
	wire [4-1:0] node4695;
	wire [4-1:0] node4696;
	wire [4-1:0] node4699;
	wire [4-1:0] node4702;
	wire [4-1:0] node4703;
	wire [4-1:0] node4704;
	wire [4-1:0] node4707;
	wire [4-1:0] node4709;
	wire [4-1:0] node4712;
	wire [4-1:0] node4713;
	wire [4-1:0] node4715;
	wire [4-1:0] node4719;
	wire [4-1:0] node4720;
	wire [4-1:0] node4721;
	wire [4-1:0] node4723;
	wire [4-1:0] node4726;
	wire [4-1:0] node4727;
	wire [4-1:0] node4730;
	wire [4-1:0] node4731;
	wire [4-1:0] node4734;
	wire [4-1:0] node4737;
	wire [4-1:0] node4738;
	wire [4-1:0] node4739;
	wire [4-1:0] node4742;
	wire [4-1:0] node4745;
	wire [4-1:0] node4746;
	wire [4-1:0] node4750;
	wire [4-1:0] node4751;
	wire [4-1:0] node4752;
	wire [4-1:0] node4753;
	wire [4-1:0] node4754;
	wire [4-1:0] node4755;
	wire [4-1:0] node4756;
	wire [4-1:0] node4757;
	wire [4-1:0] node4759;
	wire [4-1:0] node4763;
	wire [4-1:0] node4764;
	wire [4-1:0] node4767;
	wire [4-1:0] node4770;
	wire [4-1:0] node4771;
	wire [4-1:0] node4773;
	wire [4-1:0] node4774;
	wire [4-1:0] node4777;
	wire [4-1:0] node4780;
	wire [4-1:0] node4782;
	wire [4-1:0] node4783;
	wire [4-1:0] node4786;
	wire [4-1:0] node4789;
	wire [4-1:0] node4790;
	wire [4-1:0] node4791;
	wire [4-1:0] node4794;
	wire [4-1:0] node4797;
	wire [4-1:0] node4798;
	wire [4-1:0] node4800;
	wire [4-1:0] node4801;
	wire [4-1:0] node4804;
	wire [4-1:0] node4807;
	wire [4-1:0] node4808;
	wire [4-1:0] node4809;
	wire [4-1:0] node4812;
	wire [4-1:0] node4815;
	wire [4-1:0] node4816;
	wire [4-1:0] node4820;
	wire [4-1:0] node4821;
	wire [4-1:0] node4822;
	wire [4-1:0] node4823;
	wire [4-1:0] node4824;
	wire [4-1:0] node4825;
	wire [4-1:0] node4828;
	wire [4-1:0] node4831;
	wire [4-1:0] node4832;
	wire [4-1:0] node4835;
	wire [4-1:0] node4838;
	wire [4-1:0] node4839;
	wire [4-1:0] node4841;
	wire [4-1:0] node4844;
	wire [4-1:0] node4845;
	wire [4-1:0] node4849;
	wire [4-1:0] node4850;
	wire [4-1:0] node4851;
	wire [4-1:0] node4854;
	wire [4-1:0] node4857;
	wire [4-1:0] node4858;
	wire [4-1:0] node4859;
	wire [4-1:0] node4863;
	wire [4-1:0] node4864;
	wire [4-1:0] node4868;
	wire [4-1:0] node4869;
	wire [4-1:0] node4870;
	wire [4-1:0] node4871;
	wire [4-1:0] node4875;
	wire [4-1:0] node4876;
	wire [4-1:0] node4879;
	wire [4-1:0] node4882;
	wire [4-1:0] node4883;
	wire [4-1:0] node4886;
	wire [4-1:0] node4889;
	wire [4-1:0] node4890;
	wire [4-1:0] node4891;
	wire [4-1:0] node4892;
	wire [4-1:0] node4893;
	wire [4-1:0] node4895;
	wire [4-1:0] node4898;
	wire [4-1:0] node4900;
	wire [4-1:0] node4903;
	wire [4-1:0] node4904;
	wire [4-1:0] node4907;
	wire [4-1:0] node4909;
	wire [4-1:0] node4912;
	wire [4-1:0] node4913;
	wire [4-1:0] node4914;
	wire [4-1:0] node4918;
	wire [4-1:0] node4919;
	wire [4-1:0] node4923;
	wire [4-1:0] node4924;
	wire [4-1:0] node4925;
	wire [4-1:0] node4926;
	wire [4-1:0] node4928;
	wire [4-1:0] node4931;
	wire [4-1:0] node4933;
	wire [4-1:0] node4936;
	wire [4-1:0] node4937;
	wire [4-1:0] node4939;
	wire [4-1:0] node4942;
	wire [4-1:0] node4944;
	wire [4-1:0] node4947;
	wire [4-1:0] node4948;
	wire [4-1:0] node4950;
	wire [4-1:0] node4951;
	wire [4-1:0] node4952;
	wire [4-1:0] node4956;
	wire [4-1:0] node4957;
	wire [4-1:0] node4961;
	wire [4-1:0] node4962;
	wire [4-1:0] node4966;
	wire [4-1:0] node4967;
	wire [4-1:0] node4968;
	wire [4-1:0] node4969;
	wire [4-1:0] node4970;
	wire [4-1:0] node4973;
	wire [4-1:0] node4975;
	wire [4-1:0] node4978;
	wire [4-1:0] node4979;
	wire [4-1:0] node4980;
	wire [4-1:0] node4981;
	wire [4-1:0] node4984;
	wire [4-1:0] node4987;
	wire [4-1:0] node4989;
	wire [4-1:0] node4992;
	wire [4-1:0] node4993;
	wire [4-1:0] node4996;
	wire [4-1:0] node4999;
	wire [4-1:0] node5000;
	wire [4-1:0] node5001;
	wire [4-1:0] node5002;
	wire [4-1:0] node5003;
	wire [4-1:0] node5006;
	wire [4-1:0] node5009;
	wire [4-1:0] node5010;
	wire [4-1:0] node5013;
	wire [4-1:0] node5016;
	wire [4-1:0] node5017;
	wire [4-1:0] node5020;
	wire [4-1:0] node5023;
	wire [4-1:0] node5024;
	wire [4-1:0] node5027;
	wire [4-1:0] node5029;
	wire [4-1:0] node5032;
	wire [4-1:0] node5033;
	wire [4-1:0] node5034;
	wire [4-1:0] node5035;
	wire [4-1:0] node5037;
	wire [4-1:0] node5040;
	wire [4-1:0] node5041;
	wire [4-1:0] node5042;
	wire [4-1:0] node5043;
	wire [4-1:0] node5046;
	wire [4-1:0] node5049;
	wire [4-1:0] node5050;
	wire [4-1:0] node5053;
	wire [4-1:0] node5056;
	wire [4-1:0] node5057;
	wire [4-1:0] node5060;
	wire [4-1:0] node5063;
	wire [4-1:0] node5064;
	wire [4-1:0] node5065;
	wire [4-1:0] node5068;
	wire [4-1:0] node5071;
	wire [4-1:0] node5072;
	wire [4-1:0] node5074;
	wire [4-1:0] node5077;
	wire [4-1:0] node5078;
	wire [4-1:0] node5082;
	wire [4-1:0] node5083;
	wire [4-1:0] node5084;
	wire [4-1:0] node5085;
	wire [4-1:0] node5088;
	wire [4-1:0] node5091;
	wire [4-1:0] node5092;
	wire [4-1:0] node5095;
	wire [4-1:0] node5098;
	wire [4-1:0] node5099;
	wire [4-1:0] node5100;
	wire [4-1:0] node5103;
	wire [4-1:0] node5106;
	wire [4-1:0] node5107;
	wire [4-1:0] node5108;
	wire [4-1:0] node5111;
	wire [4-1:0] node5115;
	wire [4-1:0] node5116;
	wire [4-1:0] node5117;
	wire [4-1:0] node5118;
	wire [4-1:0] node5119;
	wire [4-1:0] node5120;
	wire [4-1:0] node5121;
	wire [4-1:0] node5122;
	wire [4-1:0] node5123;
	wire [4-1:0] node5124;
	wire [4-1:0] node5128;
	wire [4-1:0] node5129;
	wire [4-1:0] node5133;
	wire [4-1:0] node5134;
	wire [4-1:0] node5135;
	wire [4-1:0] node5138;
	wire [4-1:0] node5141;
	wire [4-1:0] node5142;
	wire [4-1:0] node5145;
	wire [4-1:0] node5146;
	wire [4-1:0] node5150;
	wire [4-1:0] node5151;
	wire [4-1:0] node5152;
	wire [4-1:0] node5153;
	wire [4-1:0] node5154;
	wire [4-1:0] node5157;
	wire [4-1:0] node5160;
	wire [4-1:0] node5161;
	wire [4-1:0] node5164;
	wire [4-1:0] node5167;
	wire [4-1:0] node5168;
	wire [4-1:0] node5171;
	wire [4-1:0] node5174;
	wire [4-1:0] node5175;
	wire [4-1:0] node5176;
	wire [4-1:0] node5177;
	wire [4-1:0] node5180;
	wire [4-1:0] node5184;
	wire [4-1:0] node5185;
	wire [4-1:0] node5187;
	wire [4-1:0] node5190;
	wire [4-1:0] node5191;
	wire [4-1:0] node5195;
	wire [4-1:0] node5196;
	wire [4-1:0] node5197;
	wire [4-1:0] node5198;
	wire [4-1:0] node5199;
	wire [4-1:0] node5202;
	wire [4-1:0] node5205;
	wire [4-1:0] node5206;
	wire [4-1:0] node5207;
	wire [4-1:0] node5211;
	wire [4-1:0] node5213;
	wire [4-1:0] node5216;
	wire [4-1:0] node5217;
	wire [4-1:0] node5219;
	wire [4-1:0] node5220;
	wire [4-1:0] node5223;
	wire [4-1:0] node5226;
	wire [4-1:0] node5227;
	wire [4-1:0] node5230;
	wire [4-1:0] node5233;
	wire [4-1:0] node5234;
	wire [4-1:0] node5235;
	wire [4-1:0] node5237;
	wire [4-1:0] node5240;
	wire [4-1:0] node5241;
	wire [4-1:0] node5245;
	wire [4-1:0] node5246;
	wire [4-1:0] node5249;
	wire [4-1:0] node5252;
	wire [4-1:0] node5253;
	wire [4-1:0] node5254;
	wire [4-1:0] node5255;
	wire [4-1:0] node5256;
	wire [4-1:0] node5257;
	wire [4-1:0] node5261;
	wire [4-1:0] node5262;
	wire [4-1:0] node5266;
	wire [4-1:0] node5267;
	wire [4-1:0] node5268;
	wire [4-1:0] node5269;
	wire [4-1:0] node5272;
	wire [4-1:0] node5276;
	wire [4-1:0] node5277;
	wire [4-1:0] node5280;
	wire [4-1:0] node5283;
	wire [4-1:0] node5284;
	wire [4-1:0] node5285;
	wire [4-1:0] node5286;
	wire [4-1:0] node5289;
	wire [4-1:0] node5292;
	wire [4-1:0] node5293;
	wire [4-1:0] node5294;
	wire [4-1:0] node5297;
	wire [4-1:0] node5301;
	wire [4-1:0] node5302;
	wire [4-1:0] node5303;
	wire [4-1:0] node5304;
	wire [4-1:0] node5307;
	wire [4-1:0] node5310;
	wire [4-1:0] node5311;
	wire [4-1:0] node5315;
	wire [4-1:0] node5317;
	wire [4-1:0] node5320;
	wire [4-1:0] node5321;
	wire [4-1:0] node5322;
	wire [4-1:0] node5323;
	wire [4-1:0] node5324;
	wire [4-1:0] node5327;
	wire [4-1:0] node5330;
	wire [4-1:0] node5331;
	wire [4-1:0] node5335;
	wire [4-1:0] node5336;
	wire [4-1:0] node5339;
	wire [4-1:0] node5342;
	wire [4-1:0] node5343;
	wire [4-1:0] node5344;
	wire [4-1:0] node5345;
	wire [4-1:0] node5346;
	wire [4-1:0] node5350;
	wire [4-1:0] node5351;
	wire [4-1:0] node5356;
	wire [4-1:0] node5357;
	wire [4-1:0] node5359;
	wire [4-1:0] node5362;
	wire [4-1:0] node5363;
	wire [4-1:0] node5366;
	wire [4-1:0] node5369;
	wire [4-1:0] node5370;
	wire [4-1:0] node5371;
	wire [4-1:0] node5372;
	wire [4-1:0] node5373;
	wire [4-1:0] node5374;
	wire [4-1:0] node5375;
	wire [4-1:0] node5378;
	wire [4-1:0] node5381;
	wire [4-1:0] node5382;
	wire [4-1:0] node5384;
	wire [4-1:0] node5388;
	wire [4-1:0] node5390;
	wire [4-1:0] node5393;
	wire [4-1:0] node5394;
	wire [4-1:0] node5395;
	wire [4-1:0] node5398;
	wire [4-1:0] node5399;
	wire [4-1:0] node5400;
	wire [4-1:0] node5405;
	wire [4-1:0] node5406;
	wire [4-1:0] node5407;
	wire [4-1:0] node5409;
	wire [4-1:0] node5412;
	wire [4-1:0] node5414;
	wire [4-1:0] node5417;
	wire [4-1:0] node5419;
	wire [4-1:0] node5421;
	wire [4-1:0] node5424;
	wire [4-1:0] node5425;
	wire [4-1:0] node5426;
	wire [4-1:0] node5427;
	wire [4-1:0] node5430;
	wire [4-1:0] node5431;
	wire [4-1:0] node5435;
	wire [4-1:0] node5436;
	wire [4-1:0] node5438;
	wire [4-1:0] node5441;
	wire [4-1:0] node5444;
	wire [4-1:0] node5445;
	wire [4-1:0] node5446;
	wire [4-1:0] node5448;
	wire [4-1:0] node5451;
	wire [4-1:0] node5452;
	wire [4-1:0] node5453;
	wire [4-1:0] node5457;
	wire [4-1:0] node5460;
	wire [4-1:0] node5461;
	wire [4-1:0] node5462;
	wire [4-1:0] node5466;
	wire [4-1:0] node5467;
	wire [4-1:0] node5468;
	wire [4-1:0] node5472;
	wire [4-1:0] node5475;
	wire [4-1:0] node5476;
	wire [4-1:0] node5477;
	wire [4-1:0] node5478;
	wire [4-1:0] node5479;
	wire [4-1:0] node5480;
	wire [4-1:0] node5483;
	wire [4-1:0] node5486;
	wire [4-1:0] node5487;
	wire [4-1:0] node5490;
	wire [4-1:0] node5493;
	wire [4-1:0] node5494;
	wire [4-1:0] node5497;
	wire [4-1:0] node5500;
	wire [4-1:0] node5501;
	wire [4-1:0] node5502;
	wire [4-1:0] node5503;
	wire [4-1:0] node5507;
	wire [4-1:0] node5508;
	wire [4-1:0] node5512;
	wire [4-1:0] node5513;
	wire [4-1:0] node5514;
	wire [4-1:0] node5518;
	wire [4-1:0] node5519;
	wire [4-1:0] node5523;
	wire [4-1:0] node5524;
	wire [4-1:0] node5525;
	wire [4-1:0] node5526;
	wire [4-1:0] node5527;
	wire [4-1:0] node5528;
	wire [4-1:0] node5531;
	wire [4-1:0] node5534;
	wire [4-1:0] node5535;
	wire [4-1:0] node5540;
	wire [4-1:0] node5541;
	wire [4-1:0] node5542;
	wire [4-1:0] node5543;
	wire [4-1:0] node5546;
	wire [4-1:0] node5550;
	wire [4-1:0] node5551;
	wire [4-1:0] node5554;
	wire [4-1:0] node5557;
	wire [4-1:0] node5558;
	wire [4-1:0] node5559;
	wire [4-1:0] node5560;
	wire [4-1:0] node5564;
	wire [4-1:0] node5565;
	wire [4-1:0] node5569;
	wire [4-1:0] node5570;
	wire [4-1:0] node5571;
	wire [4-1:0] node5575;
	wire [4-1:0] node5577;
	wire [4-1:0] node5580;
	wire [4-1:0] node5581;
	wire [4-1:0] node5582;
	wire [4-1:0] node5583;
	wire [4-1:0] node5584;
	wire [4-1:0] node5585;
	wire [4-1:0] node5586;
	wire [4-1:0] node5587;
	wire [4-1:0] node5592;
	wire [4-1:0] node5593;
	wire [4-1:0] node5594;
	wire [4-1:0] node5598;
	wire [4-1:0] node5599;
	wire [4-1:0] node5603;
	wire [4-1:0] node5604;
	wire [4-1:0] node5605;
	wire [4-1:0] node5606;
	wire [4-1:0] node5610;
	wire [4-1:0] node5611;
	wire [4-1:0] node5615;
	wire [4-1:0] node5616;
	wire [4-1:0] node5617;
	wire [4-1:0] node5621;
	wire [4-1:0] node5622;
	wire [4-1:0] node5626;
	wire [4-1:0] node5627;
	wire [4-1:0] node5629;
	wire [4-1:0] node5630;
	wire [4-1:0] node5634;
	wire [4-1:0] node5635;
	wire [4-1:0] node5636;
	wire [4-1:0] node5640;
	wire [4-1:0] node5641;
	wire [4-1:0] node5645;
	wire [4-1:0] node5646;
	wire [4-1:0] node5647;
	wire [4-1:0] node5648;
	wire [4-1:0] node5649;
	wire [4-1:0] node5653;
	wire [4-1:0] node5654;
	wire [4-1:0] node5658;
	wire [4-1:0] node5659;
	wire [4-1:0] node5660;
	wire [4-1:0] node5664;
	wire [4-1:0] node5665;
	wire [4-1:0] node5669;
	wire [4-1:0] node5670;
	wire [4-1:0] node5671;
	wire [4-1:0] node5672;
	wire [4-1:0] node5673;
	wire [4-1:0] node5674;
	wire [4-1:0] node5677;
	wire [4-1:0] node5680;
	wire [4-1:0] node5681;
	wire [4-1:0] node5685;
	wire [4-1:0] node5687;
	wire [4-1:0] node5690;
	wire [4-1:0] node5691;
	wire [4-1:0] node5692;
	wire [4-1:0] node5695;
	wire [4-1:0] node5698;
	wire [4-1:0] node5700;
	wire [4-1:0] node5703;
	wire [4-1:0] node5704;
	wire [4-1:0] node5705;
	wire [4-1:0] node5707;
	wire [4-1:0] node5708;
	wire [4-1:0] node5711;
	wire [4-1:0] node5714;
	wire [4-1:0] node5716;
	wire [4-1:0] node5719;
	wire [4-1:0] node5721;
	wire [4-1:0] node5722;
	wire [4-1:0] node5725;
	wire [4-1:0] node5728;
	wire [4-1:0] node5729;
	wire [4-1:0] node5730;
	wire [4-1:0] node5731;
	wire [4-1:0] node5732;
	wire [4-1:0] node5733;
	wire [4-1:0] node5734;
	wire [4-1:0] node5738;
	wire [4-1:0] node5739;
	wire [4-1:0] node5743;
	wire [4-1:0] node5744;
	wire [4-1:0] node5747;
	wire [4-1:0] node5748;
	wire [4-1:0] node5752;
	wire [4-1:0] node5753;
	wire [4-1:0] node5754;
	wire [4-1:0] node5756;
	wire [4-1:0] node5757;
	wire [4-1:0] node5761;
	wire [4-1:0] node5762;
	wire [4-1:0] node5763;
	wire [4-1:0] node5767;
	wire [4-1:0] node5770;
	wire [4-1:0] node5771;
	wire [4-1:0] node5774;
	wire [4-1:0] node5775;
	wire [4-1:0] node5779;
	wire [4-1:0] node5780;
	wire [4-1:0] node5781;
	wire [4-1:0] node5783;
	wire [4-1:0] node5784;
	wire [4-1:0] node5788;
	wire [4-1:0] node5789;
	wire [4-1:0] node5790;
	wire [4-1:0] node5794;
	wire [4-1:0] node5797;
	wire [4-1:0] node5798;
	wire [4-1:0] node5799;
	wire [4-1:0] node5800;
	wire [4-1:0] node5801;
	wire [4-1:0] node5805;
	wire [4-1:0] node5806;
	wire [4-1:0] node5809;
	wire [4-1:0] node5812;
	wire [4-1:0] node5813;
	wire [4-1:0] node5817;
	wire [4-1:0] node5818;
	wire [4-1:0] node5821;
	wire [4-1:0] node5824;
	wire [4-1:0] node5825;
	wire [4-1:0] node5826;
	wire [4-1:0] node5827;
	wire [4-1:0] node5828;
	wire [4-1:0] node5829;
	wire [4-1:0] node5830;
	wire [4-1:0] node5833;
	wire [4-1:0] node5836;
	wire [4-1:0] node5837;
	wire [4-1:0] node5841;
	wire [4-1:0] node5842;
	wire [4-1:0] node5845;
	wire [4-1:0] node5846;
	wire [4-1:0] node5849;
	wire [4-1:0] node5852;
	wire [4-1:0] node5853;
	wire [4-1:0] node5854;
	wire [4-1:0] node5855;
	wire [4-1:0] node5859;
	wire [4-1:0] node5862;
	wire [4-1:0] node5863;
	wire [4-1:0] node5864;
	wire [4-1:0] node5868;
	wire [4-1:0] node5869;
	wire [4-1:0] node5872;
	wire [4-1:0] node5875;
	wire [4-1:0] node5876;
	wire [4-1:0] node5877;
	wire [4-1:0] node5879;
	wire [4-1:0] node5882;
	wire [4-1:0] node5884;
	wire [4-1:0] node5887;
	wire [4-1:0] node5888;
	wire [4-1:0] node5889;
	wire [4-1:0] node5892;
	wire [4-1:0] node5895;
	wire [4-1:0] node5898;
	wire [4-1:0] node5899;
	wire [4-1:0] node5900;
	wire [4-1:0] node5902;
	wire [4-1:0] node5903;
	wire [4-1:0] node5906;
	wire [4-1:0] node5909;
	wire [4-1:0] node5910;
	wire [4-1:0] node5911;
	wire [4-1:0] node5912;
	wire [4-1:0] node5915;
	wire [4-1:0] node5919;
	wire [4-1:0] node5922;
	wire [4-1:0] node5923;
	wire [4-1:0] node5924;
	wire [4-1:0] node5925;
	wire [4-1:0] node5927;
	wire [4-1:0] node5930;
	wire [4-1:0] node5933;
	wire [4-1:0] node5934;
	wire [4-1:0] node5935;
	wire [4-1:0] node5938;
	wire [4-1:0] node5942;
	wire [4-1:0] node5943;
	wire [4-1:0] node5944;
	wire [4-1:0] node5946;
	wire [4-1:0] node5950;
	wire [4-1:0] node5951;
	wire [4-1:0] node5952;
	wire [4-1:0] node5956;
	wire [4-1:0] node5957;
	wire [4-1:0] node5960;
	wire [4-1:0] node5963;
	wire [4-1:0] node5964;
	wire [4-1:0] node5965;
	wire [4-1:0] node5966;
	wire [4-1:0] node5967;
	wire [4-1:0] node5968;
	wire [4-1:0] node5969;
	wire [4-1:0] node5970;
	wire [4-1:0] node5971;
	wire [4-1:0] node5974;
	wire [4-1:0] node5977;
	wire [4-1:0] node5978;
	wire [4-1:0] node5981;
	wire [4-1:0] node5984;
	wire [4-1:0] node5985;
	wire [4-1:0] node5986;
	wire [4-1:0] node5989;
	wire [4-1:0] node5992;
	wire [4-1:0] node5993;
	wire [4-1:0] node5994;
	wire [4-1:0] node5998;
	wire [4-1:0] node6000;
	wire [4-1:0] node6003;
	wire [4-1:0] node6004;
	wire [4-1:0] node6005;
	wire [4-1:0] node6008;
	wire [4-1:0] node6011;
	wire [4-1:0] node6012;
	wire [4-1:0] node6015;
	wire [4-1:0] node6018;
	wire [4-1:0] node6019;
	wire [4-1:0] node6020;
	wire [4-1:0] node6021;
	wire [4-1:0] node6024;
	wire [4-1:0] node6027;
	wire [4-1:0] node6028;
	wire [4-1:0] node6030;
	wire [4-1:0] node6033;
	wire [4-1:0] node6034;
	wire [4-1:0] node6037;
	wire [4-1:0] node6040;
	wire [4-1:0] node6041;
	wire [4-1:0] node6042;
	wire [4-1:0] node6043;
	wire [4-1:0] node6046;
	wire [4-1:0] node6049;
	wire [4-1:0] node6051;
	wire [4-1:0] node6052;
	wire [4-1:0] node6055;
	wire [4-1:0] node6058;
	wire [4-1:0] node6059;
	wire [4-1:0] node6060;
	wire [4-1:0] node6061;
	wire [4-1:0] node6065;
	wire [4-1:0] node6068;
	wire [4-1:0] node6069;
	wire [4-1:0] node6072;
	wire [4-1:0] node6075;
	wire [4-1:0] node6076;
	wire [4-1:0] node6077;
	wire [4-1:0] node6078;
	wire [4-1:0] node6080;
	wire [4-1:0] node6081;
	wire [4-1:0] node6084;
	wire [4-1:0] node6087;
	wire [4-1:0] node6088;
	wire [4-1:0] node6090;
	wire [4-1:0] node6093;
	wire [4-1:0] node6094;
	wire [4-1:0] node6097;
	wire [4-1:0] node6100;
	wire [4-1:0] node6101;
	wire [4-1:0] node6102;
	wire [4-1:0] node6105;
	wire [4-1:0] node6108;
	wire [4-1:0] node6109;
	wire [4-1:0] node6110;
	wire [4-1:0] node6114;
	wire [4-1:0] node6115;
	wire [4-1:0] node6118;
	wire [4-1:0] node6121;
	wire [4-1:0] node6122;
	wire [4-1:0] node6123;
	wire [4-1:0] node6124;
	wire [4-1:0] node6125;
	wire [4-1:0] node6127;
	wire [4-1:0] node6131;
	wire [4-1:0] node6133;
	wire [4-1:0] node6136;
	wire [4-1:0] node6137;
	wire [4-1:0] node6140;
	wire [4-1:0] node6143;
	wire [4-1:0] node6144;
	wire [4-1:0] node6145;
	wire [4-1:0] node6146;
	wire [4-1:0] node6150;
	wire [4-1:0] node6151;
	wire [4-1:0] node6155;
	wire [4-1:0] node6157;
	wire [4-1:0] node6160;
	wire [4-1:0] node6161;
	wire [4-1:0] node6162;
	wire [4-1:0] node6163;
	wire [4-1:0] node6164;
	wire [4-1:0] node6165;
	wire [4-1:0] node6166;
	wire [4-1:0] node6167;
	wire [4-1:0] node6170;
	wire [4-1:0] node6174;
	wire [4-1:0] node6176;
	wire [4-1:0] node6177;
	wire [4-1:0] node6180;
	wire [4-1:0] node6183;
	wire [4-1:0] node6184;
	wire [4-1:0] node6186;
	wire [4-1:0] node6187;
	wire [4-1:0] node6191;
	wire [4-1:0] node6192;
	wire [4-1:0] node6195;
	wire [4-1:0] node6198;
	wire [4-1:0] node6199;
	wire [4-1:0] node6200;
	wire [4-1:0] node6201;
	wire [4-1:0] node6205;
	wire [4-1:0] node6206;
	wire [4-1:0] node6210;
	wire [4-1:0] node6211;
	wire [4-1:0] node6212;
	wire [4-1:0] node6215;
	wire [4-1:0] node6218;
	wire [4-1:0] node6221;
	wire [4-1:0] node6222;
	wire [4-1:0] node6223;
	wire [4-1:0] node6224;
	wire [4-1:0] node6225;
	wire [4-1:0] node6228;
	wire [4-1:0] node6231;
	wire [4-1:0] node6233;
	wire [4-1:0] node6236;
	wire [4-1:0] node6237;
	wire [4-1:0] node6238;
	wire [4-1:0] node6239;
	wire [4-1:0] node6243;
	wire [4-1:0] node6245;
	wire [4-1:0] node6248;
	wire [4-1:0] node6249;
	wire [4-1:0] node6250;
	wire [4-1:0] node6255;
	wire [4-1:0] node6256;
	wire [4-1:0] node6257;
	wire [4-1:0] node6259;
	wire [4-1:0] node6262;
	wire [4-1:0] node6263;
	wire [4-1:0] node6266;
	wire [4-1:0] node6269;
	wire [4-1:0] node6270;
	wire [4-1:0] node6272;
	wire [4-1:0] node6275;
	wire [4-1:0] node6276;
	wire [4-1:0] node6277;
	wire [4-1:0] node6281;
	wire [4-1:0] node6282;
	wire [4-1:0] node6286;
	wire [4-1:0] node6287;
	wire [4-1:0] node6288;
	wire [4-1:0] node6289;
	wire [4-1:0] node6290;
	wire [4-1:0] node6291;
	wire [4-1:0] node6293;
	wire [4-1:0] node6296;
	wire [4-1:0] node6297;
	wire [4-1:0] node6301;
	wire [4-1:0] node6302;
	wire [4-1:0] node6303;
	wire [4-1:0] node6306;
	wire [4-1:0] node6309;
	wire [4-1:0] node6311;
	wire [4-1:0] node6314;
	wire [4-1:0] node6315;
	wire [4-1:0] node6316;
	wire [4-1:0] node6317;
	wire [4-1:0] node6322;
	wire [4-1:0] node6323;
	wire [4-1:0] node6326;
	wire [4-1:0] node6329;
	wire [4-1:0] node6330;
	wire [4-1:0] node6331;
	wire [4-1:0] node6332;
	wire [4-1:0] node6335;
	wire [4-1:0] node6338;
	wire [4-1:0] node6339;
	wire [4-1:0] node6340;
	wire [4-1:0] node6343;
	wire [4-1:0] node6347;
	wire [4-1:0] node6350;
	wire [4-1:0] node6351;
	wire [4-1:0] node6352;
	wire [4-1:0] node6353;
	wire [4-1:0] node6354;
	wire [4-1:0] node6357;
	wire [4-1:0] node6360;
	wire [4-1:0] node6362;
	wire [4-1:0] node6363;
	wire [4-1:0] node6367;
	wire [4-1:0] node6368;
	wire [4-1:0] node6369;
	wire [4-1:0] node6373;
	wire [4-1:0] node6375;
	wire [4-1:0] node6376;
	wire [4-1:0] node6379;
	wire [4-1:0] node6382;
	wire [4-1:0] node6383;
	wire [4-1:0] node6384;
	wire [4-1:0] node6386;
	wire [4-1:0] node6388;
	wire [4-1:0] node6391;
	wire [4-1:0] node6392;
	wire [4-1:0] node6393;
	wire [4-1:0] node6398;
	wire [4-1:0] node6399;
	wire [4-1:0] node6400;
	wire [4-1:0] node6401;
	wire [4-1:0] node6404;
	wire [4-1:0] node6407;
	wire [4-1:0] node6409;
	wire [4-1:0] node6412;
	wire [4-1:0] node6414;
	wire [4-1:0] node6417;
	wire [4-1:0] node6418;
	wire [4-1:0] node6419;
	wire [4-1:0] node6420;
	wire [4-1:0] node6421;
	wire [4-1:0] node6422;
	wire [4-1:0] node6423;
	wire [4-1:0] node6424;
	wire [4-1:0] node6427;
	wire [4-1:0] node6431;
	wire [4-1:0] node6432;
	wire [4-1:0] node6433;
	wire [4-1:0] node6434;
	wire [4-1:0] node6437;
	wire [4-1:0] node6441;
	wire [4-1:0] node6442;
	wire [4-1:0] node6446;
	wire [4-1:0] node6447;
	wire [4-1:0] node6449;
	wire [4-1:0] node6452;
	wire [4-1:0] node6453;
	wire [4-1:0] node6454;
	wire [4-1:0] node6457;
	wire [4-1:0] node6460;
	wire [4-1:0] node6462;
	wire [4-1:0] node6465;
	wire [4-1:0] node6466;
	wire [4-1:0] node6467;
	wire [4-1:0] node6468;
	wire [4-1:0] node6469;
	wire [4-1:0] node6472;
	wire [4-1:0] node6475;
	wire [4-1:0] node6476;
	wire [4-1:0] node6477;
	wire [4-1:0] node6481;
	wire [4-1:0] node6483;
	wire [4-1:0] node6486;
	wire [4-1:0] node6487;
	wire [4-1:0] node6491;
	wire [4-1:0] node6492;
	wire [4-1:0] node6495;
	wire [4-1:0] node6498;
	wire [4-1:0] node6499;
	wire [4-1:0] node6500;
	wire [4-1:0] node6501;
	wire [4-1:0] node6502;
	wire [4-1:0] node6506;
	wire [4-1:0] node6507;
	wire [4-1:0] node6511;
	wire [4-1:0] node6512;
	wire [4-1:0] node6513;
	wire [4-1:0] node6517;
	wire [4-1:0] node6518;
	wire [4-1:0] node6522;
	wire [4-1:0] node6523;
	wire [4-1:0] node6524;
	wire [4-1:0] node6525;
	wire [4-1:0] node6526;
	wire [4-1:0] node6529;
	wire [4-1:0] node6533;
	wire [4-1:0] node6534;
	wire [4-1:0] node6536;
	wire [4-1:0] node6540;
	wire [4-1:0] node6541;
	wire [4-1:0] node6542;
	wire [4-1:0] node6543;
	wire [4-1:0] node6548;
	wire [4-1:0] node6549;
	wire [4-1:0] node6550;
	wire [4-1:0] node6554;
	wire [4-1:0] node6555;
	wire [4-1:0] node6559;
	wire [4-1:0] node6560;
	wire [4-1:0] node6561;
	wire [4-1:0] node6562;
	wire [4-1:0] node6563;
	wire [4-1:0] node6564;
	wire [4-1:0] node6566;
	wire [4-1:0] node6567;
	wire [4-1:0] node6570;
	wire [4-1:0] node6573;
	wire [4-1:0] node6574;
	wire [4-1:0] node6577;
	wire [4-1:0] node6580;
	wire [4-1:0] node6581;
	wire [4-1:0] node6582;
	wire [4-1:0] node6583;
	wire [4-1:0] node6587;
	wire [4-1:0] node6589;
	wire [4-1:0] node6592;
	wire [4-1:0] node6595;
	wire [4-1:0] node6596;
	wire [4-1:0] node6597;
	wire [4-1:0] node6600;
	wire [4-1:0] node6601;
	wire [4-1:0] node6605;
	wire [4-1:0] node6606;
	wire [4-1:0] node6607;
	wire [4-1:0] node6611;
	wire [4-1:0] node6612;
	wire [4-1:0] node6616;
	wire [4-1:0] node6617;
	wire [4-1:0] node6618;
	wire [4-1:0] node6620;
	wire [4-1:0] node6621;
	wire [4-1:0] node6625;
	wire [4-1:0] node6626;
	wire [4-1:0] node6627;
	wire [4-1:0] node6628;
	wire [4-1:0] node6633;
	wire [4-1:0] node6634;
	wire [4-1:0] node6635;
	wire [4-1:0] node6640;
	wire [4-1:0] node6641;
	wire [4-1:0] node6642;
	wire [4-1:0] node6644;
	wire [4-1:0] node6645;
	wire [4-1:0] node6648;
	wire [4-1:0] node6651;
	wire [4-1:0] node6652;
	wire [4-1:0] node6655;
	wire [4-1:0] node6658;
	wire [4-1:0] node6659;
	wire [4-1:0] node6660;
	wire [4-1:0] node6661;
	wire [4-1:0] node6664;
	wire [4-1:0] node6667;
	wire [4-1:0] node6668;
	wire [4-1:0] node6671;
	wire [4-1:0] node6674;
	wire [4-1:0] node6676;
	wire [4-1:0] node6677;
	wire [4-1:0] node6680;
	wire [4-1:0] node6683;
	wire [4-1:0] node6684;
	wire [4-1:0] node6685;
	wire [4-1:0] node6686;
	wire [4-1:0] node6687;
	wire [4-1:0] node6688;
	wire [4-1:0] node6689;
	wire [4-1:0] node6692;
	wire [4-1:0] node6695;
	wire [4-1:0] node6697;
	wire [4-1:0] node6700;
	wire [4-1:0] node6703;
	wire [4-1:0] node6704;
	wire [4-1:0] node6705;
	wire [4-1:0] node6708;
	wire [4-1:0] node6712;
	wire [4-1:0] node6713;
	wire [4-1:0] node6714;
	wire [4-1:0] node6715;
	wire [4-1:0] node6717;
	wire [4-1:0] node6721;
	wire [4-1:0] node6722;
	wire [4-1:0] node6725;
	wire [4-1:0] node6728;
	wire [4-1:0] node6729;
	wire [4-1:0] node6731;
	wire [4-1:0] node6734;
	wire [4-1:0] node6735;
	wire [4-1:0] node6738;
	wire [4-1:0] node6741;
	wire [4-1:0] node6742;
	wire [4-1:0] node6743;
	wire [4-1:0] node6744;
	wire [4-1:0] node6745;
	wire [4-1:0] node6748;
	wire [4-1:0] node6751;
	wire [4-1:0] node6752;
	wire [4-1:0] node6755;
	wire [4-1:0] node6758;
	wire [4-1:0] node6759;
	wire [4-1:0] node6760;
	wire [4-1:0] node6763;
	wire [4-1:0] node6766;
	wire [4-1:0] node6767;
	wire [4-1:0] node6771;
	wire [4-1:0] node6772;
	wire [4-1:0] node6773;
	wire [4-1:0] node6774;
	wire [4-1:0] node6777;
	wire [4-1:0] node6780;
	wire [4-1:0] node6782;
	wire [4-1:0] node6785;
	wire [4-1:0] node6786;
	wire [4-1:0] node6789;
	wire [4-1:0] node6792;
	wire [4-1:0] node6793;
	wire [4-1:0] node6794;
	wire [4-1:0] node6795;
	wire [4-1:0] node6796;
	wire [4-1:0] node6797;
	wire [4-1:0] node6798;
	wire [4-1:0] node6799;
	wire [4-1:0] node6800;
	wire [4-1:0] node6801;
	wire [4-1:0] node6802;
	wire [4-1:0] node6803;
	wire [4-1:0] node6806;
	wire [4-1:0] node6809;
	wire [4-1:0] node6810;
	wire [4-1:0] node6813;
	wire [4-1:0] node6816;
	wire [4-1:0] node6817;
	wire [4-1:0] node6818;
	wire [4-1:0] node6819;
	wire [4-1:0] node6824;
	wire [4-1:0] node6825;
	wire [4-1:0] node6828;
	wire [4-1:0] node6831;
	wire [4-1:0] node6832;
	wire [4-1:0] node6833;
	wire [4-1:0] node6834;
	wire [4-1:0] node6837;
	wire [4-1:0] node6840;
	wire [4-1:0] node6841;
	wire [4-1:0] node6844;
	wire [4-1:0] node6847;
	wire [4-1:0] node6848;
	wire [4-1:0] node6850;
	wire [4-1:0] node6853;
	wire [4-1:0] node6854;
	wire [4-1:0] node6857;
	wire [4-1:0] node6860;
	wire [4-1:0] node6861;
	wire [4-1:0] node6862;
	wire [4-1:0] node6864;
	wire [4-1:0] node6865;
	wire [4-1:0] node6869;
	wire [4-1:0] node6870;
	wire [4-1:0] node6872;
	wire [4-1:0] node6875;
	wire [4-1:0] node6876;
	wire [4-1:0] node6879;
	wire [4-1:0] node6882;
	wire [4-1:0] node6883;
	wire [4-1:0] node6884;
	wire [4-1:0] node6885;
	wire [4-1:0] node6886;
	wire [4-1:0] node6890;
	wire [4-1:0] node6891;
	wire [4-1:0] node6895;
	wire [4-1:0] node6896;
	wire [4-1:0] node6899;
	wire [4-1:0] node6902;
	wire [4-1:0] node6903;
	wire [4-1:0] node6905;
	wire [4-1:0] node6906;
	wire [4-1:0] node6910;
	wire [4-1:0] node6912;
	wire [4-1:0] node6914;
	wire [4-1:0] node6917;
	wire [4-1:0] node6918;
	wire [4-1:0] node6919;
	wire [4-1:0] node6920;
	wire [4-1:0] node6921;
	wire [4-1:0] node6922;
	wire [4-1:0] node6925;
	wire [4-1:0] node6929;
	wire [4-1:0] node6930;
	wire [4-1:0] node6931;
	wire [4-1:0] node6934;
	wire [4-1:0] node6937;
	wire [4-1:0] node6938;
	wire [4-1:0] node6940;
	wire [4-1:0] node6943;
	wire [4-1:0] node6944;
	wire [4-1:0] node6948;
	wire [4-1:0] node6949;
	wire [4-1:0] node6950;
	wire [4-1:0] node6952;
	wire [4-1:0] node6955;
	wire [4-1:0] node6957;
	wire [4-1:0] node6960;
	wire [4-1:0] node6961;
	wire [4-1:0] node6962;
	wire [4-1:0] node6965;
	wire [4-1:0] node6968;
	wire [4-1:0] node6969;
	wire [4-1:0] node6973;
	wire [4-1:0] node6974;
	wire [4-1:0] node6975;
	wire [4-1:0] node6976;
	wire [4-1:0] node6977;
	wire [4-1:0] node6979;
	wire [4-1:0] node6982;
	wire [4-1:0] node6983;
	wire [4-1:0] node6986;
	wire [4-1:0] node6989;
	wire [4-1:0] node6991;
	wire [4-1:0] node6994;
	wire [4-1:0] node6995;
	wire [4-1:0] node6996;
	wire [4-1:0] node7000;
	wire [4-1:0] node7001;
	wire [4-1:0] node7004;
	wire [4-1:0] node7007;
	wire [4-1:0] node7008;
	wire [4-1:0] node7009;
	wire [4-1:0] node7010;
	wire [4-1:0] node7014;
	wire [4-1:0] node7015;
	wire [4-1:0] node7019;
	wire [4-1:0] node7020;
	wire [4-1:0] node7021;
	wire [4-1:0] node7024;
	wire [4-1:0] node7027;
	wire [4-1:0] node7028;
	wire [4-1:0] node7032;
	wire [4-1:0] node7033;
	wire [4-1:0] node7034;
	wire [4-1:0] node7035;
	wire [4-1:0] node7036;
	wire [4-1:0] node7038;
	wire [4-1:0] node7040;
	wire [4-1:0] node7043;
	wire [4-1:0] node7044;
	wire [4-1:0] node7045;
	wire [4-1:0] node7048;
	wire [4-1:0] node7051;
	wire [4-1:0] node7052;
	wire [4-1:0] node7055;
	wire [4-1:0] node7058;
	wire [4-1:0] node7059;
	wire [4-1:0] node7060;
	wire [4-1:0] node7061;
	wire [4-1:0] node7065;
	wire [4-1:0] node7066;
	wire [4-1:0] node7069;
	wire [4-1:0] node7072;
	wire [4-1:0] node7073;
	wire [4-1:0] node7074;
	wire [4-1:0] node7075;
	wire [4-1:0] node7079;
	wire [4-1:0] node7080;
	wire [4-1:0] node7084;
	wire [4-1:0] node7085;
	wire [4-1:0] node7087;
	wire [4-1:0] node7090;
	wire [4-1:0] node7091;
	wire [4-1:0] node7095;
	wire [4-1:0] node7096;
	wire [4-1:0] node7097;
	wire [4-1:0] node7098;
	wire [4-1:0] node7099;
	wire [4-1:0] node7102;
	wire [4-1:0] node7105;
	wire [4-1:0] node7106;
	wire [4-1:0] node7109;
	wire [4-1:0] node7112;
	wire [4-1:0] node7114;
	wire [4-1:0] node7115;
	wire [4-1:0] node7116;
	wire [4-1:0] node7120;
	wire [4-1:0] node7121;
	wire [4-1:0] node7124;
	wire [4-1:0] node7127;
	wire [4-1:0] node7128;
	wire [4-1:0] node7129;
	wire [4-1:0] node7130;
	wire [4-1:0] node7134;
	wire [4-1:0] node7135;
	wire [4-1:0] node7136;
	wire [4-1:0] node7140;
	wire [4-1:0] node7141;
	wire [4-1:0] node7144;
	wire [4-1:0] node7147;
	wire [4-1:0] node7148;
	wire [4-1:0] node7149;
	wire [4-1:0] node7153;
	wire [4-1:0] node7154;
	wire [4-1:0] node7158;
	wire [4-1:0] node7159;
	wire [4-1:0] node7160;
	wire [4-1:0] node7161;
	wire [4-1:0] node7162;
	wire [4-1:0] node7165;
	wire [4-1:0] node7168;
	wire [4-1:0] node7170;
	wire [4-1:0] node7173;
	wire [4-1:0] node7174;
	wire [4-1:0] node7175;
	wire [4-1:0] node7176;
	wire [4-1:0] node7177;
	wire [4-1:0] node7180;
	wire [4-1:0] node7183;
	wire [4-1:0] node7184;
	wire [4-1:0] node7188;
	wire [4-1:0] node7190;
	wire [4-1:0] node7193;
	wire [4-1:0] node7194;
	wire [4-1:0] node7195;
	wire [4-1:0] node7197;
	wire [4-1:0] node7200;
	wire [4-1:0] node7201;
	wire [4-1:0] node7205;
	wire [4-1:0] node7206;
	wire [4-1:0] node7209;
	wire [4-1:0] node7211;
	wire [4-1:0] node7214;
	wire [4-1:0] node7215;
	wire [4-1:0] node7216;
	wire [4-1:0] node7217;
	wire [4-1:0] node7220;
	wire [4-1:0] node7223;
	wire [4-1:0] node7224;
	wire [4-1:0] node7227;
	wire [4-1:0] node7228;
	wire [4-1:0] node7232;
	wire [4-1:0] node7233;
	wire [4-1:0] node7234;
	wire [4-1:0] node7235;
	wire [4-1:0] node7238;
	wire [4-1:0] node7241;
	wire [4-1:0] node7242;
	wire [4-1:0] node7245;
	wire [4-1:0] node7248;
	wire [4-1:0] node7249;
	wire [4-1:0] node7251;
	wire [4-1:0] node7252;
	wire [4-1:0] node7255;
	wire [4-1:0] node7258;
	wire [4-1:0] node7259;
	wire [4-1:0] node7263;
	wire [4-1:0] node7264;
	wire [4-1:0] node7265;
	wire [4-1:0] node7266;
	wire [4-1:0] node7267;
	wire [4-1:0] node7268;
	wire [4-1:0] node7269;
	wire [4-1:0] node7273;
	wire [4-1:0] node7274;
	wire [4-1:0] node7277;
	wire [4-1:0] node7280;
	wire [4-1:0] node7281;
	wire [4-1:0] node7283;
	wire [4-1:0] node7285;
	wire [4-1:0] node7288;
	wire [4-1:0] node7289;
	wire [4-1:0] node7292;
	wire [4-1:0] node7295;
	wire [4-1:0] node7296;
	wire [4-1:0] node7297;
	wire [4-1:0] node7300;
	wire [4-1:0] node7303;
	wire [4-1:0] node7304;
	wire [4-1:0] node7305;
	wire [4-1:0] node7306;
	wire [4-1:0] node7308;
	wire [4-1:0] node7312;
	wire [4-1:0] node7313;
	wire [4-1:0] node7314;
	wire [4-1:0] node7318;
	wire [4-1:0] node7320;
	wire [4-1:0] node7323;
	wire [4-1:0] node7324;
	wire [4-1:0] node7325;
	wire [4-1:0] node7329;
	wire [4-1:0] node7331;
	wire [4-1:0] node7334;
	wire [4-1:0] node7335;
	wire [4-1:0] node7336;
	wire [4-1:0] node7337;
	wire [4-1:0] node7340;
	wire [4-1:0] node7343;
	wire [4-1:0] node7344;
	wire [4-1:0] node7345;
	wire [4-1:0] node7347;
	wire [4-1:0] node7350;
	wire [4-1:0] node7352;
	wire [4-1:0] node7355;
	wire [4-1:0] node7356;
	wire [4-1:0] node7359;
	wire [4-1:0] node7362;
	wire [4-1:0] node7363;
	wire [4-1:0] node7364;
	wire [4-1:0] node7367;
	wire [4-1:0] node7370;
	wire [4-1:0] node7371;
	wire [4-1:0] node7372;
	wire [4-1:0] node7375;
	wire [4-1:0] node7378;
	wire [4-1:0] node7379;
	wire [4-1:0] node7380;
	wire [4-1:0] node7383;
	wire [4-1:0] node7386;
	wire [4-1:0] node7387;
	wire [4-1:0] node7388;
	wire [4-1:0] node7392;
	wire [4-1:0] node7394;
	wire [4-1:0] node7397;
	wire [4-1:0] node7398;
	wire [4-1:0] node7399;
	wire [4-1:0] node7400;
	wire [4-1:0] node7401;
	wire [4-1:0] node7402;
	wire [4-1:0] node7403;
	wire [4-1:0] node7406;
	wire [4-1:0] node7407;
	wire [4-1:0] node7411;
	wire [4-1:0] node7413;
	wire [4-1:0] node7416;
	wire [4-1:0] node7417;
	wire [4-1:0] node7418;
	wire [4-1:0] node7420;
	wire [4-1:0] node7423;
	wire [4-1:0] node7425;
	wire [4-1:0] node7428;
	wire [4-1:0] node7431;
	wire [4-1:0] node7432;
	wire [4-1:0] node7433;
	wire [4-1:0] node7434;
	wire [4-1:0] node7438;
	wire [4-1:0] node7439;
	wire [4-1:0] node7442;
	wire [4-1:0] node7443;
	wire [4-1:0] node7447;
	wire [4-1:0] node7448;
	wire [4-1:0] node7449;
	wire [4-1:0] node7452;
	wire [4-1:0] node7455;
	wire [4-1:0] node7456;
	wire [4-1:0] node7459;
	wire [4-1:0] node7462;
	wire [4-1:0] node7463;
	wire [4-1:0] node7464;
	wire [4-1:0] node7465;
	wire [4-1:0] node7468;
	wire [4-1:0] node7471;
	wire [4-1:0] node7472;
	wire [4-1:0] node7475;
	wire [4-1:0] node7478;
	wire [4-1:0] node7479;
	wire [4-1:0] node7480;
	wire [4-1:0] node7483;
	wire [4-1:0] node7486;
	wire [4-1:0] node7487;
	wire [4-1:0] node7488;
	wire [4-1:0] node7492;
	wire [4-1:0] node7493;
	wire [4-1:0] node7494;
	wire [4-1:0] node7499;
	wire [4-1:0] node7500;
	wire [4-1:0] node7501;
	wire [4-1:0] node7502;
	wire [4-1:0] node7503;
	wire [4-1:0] node7504;
	wire [4-1:0] node7507;
	wire [4-1:0] node7510;
	wire [4-1:0] node7511;
	wire [4-1:0] node7514;
	wire [4-1:0] node7517;
	wire [4-1:0] node7518;
	wire [4-1:0] node7520;
	wire [4-1:0] node7523;
	wire [4-1:0] node7525;
	wire [4-1:0] node7526;
	wire [4-1:0] node7529;
	wire [4-1:0] node7532;
	wire [4-1:0] node7533;
	wire [4-1:0] node7534;
	wire [4-1:0] node7535;
	wire [4-1:0] node7538;
	wire [4-1:0] node7541;
	wire [4-1:0] node7542;
	wire [4-1:0] node7543;
	wire [4-1:0] node7546;
	wire [4-1:0] node7549;
	wire [4-1:0] node7552;
	wire [4-1:0] node7553;
	wire [4-1:0] node7554;
	wire [4-1:0] node7555;
	wire [4-1:0] node7558;
	wire [4-1:0] node7562;
	wire [4-1:0] node7563;
	wire [4-1:0] node7564;
	wire [4-1:0] node7568;
	wire [4-1:0] node7569;
	wire [4-1:0] node7573;
	wire [4-1:0] node7574;
	wire [4-1:0] node7575;
	wire [4-1:0] node7576;
	wire [4-1:0] node7577;
	wire [4-1:0] node7580;
	wire [4-1:0] node7584;
	wire [4-1:0] node7585;
	wire [4-1:0] node7586;
	wire [4-1:0] node7589;
	wire [4-1:0] node7592;
	wire [4-1:0] node7593;
	wire [4-1:0] node7596;
	wire [4-1:0] node7599;
	wire [4-1:0] node7600;
	wire [4-1:0] node7601;
	wire [4-1:0] node7602;
	wire [4-1:0] node7606;
	wire [4-1:0] node7607;
	wire [4-1:0] node7608;
	wire [4-1:0] node7611;
	wire [4-1:0] node7615;
	wire [4-1:0] node7616;
	wire [4-1:0] node7619;
	wire [4-1:0] node7622;
	wire [4-1:0] node7623;
	wire [4-1:0] node7624;
	wire [4-1:0] node7625;
	wire [4-1:0] node7626;
	wire [4-1:0] node7627;
	wire [4-1:0] node7628;
	wire [4-1:0] node7629;
	wire [4-1:0] node7630;
	wire [4-1:0] node7631;
	wire [4-1:0] node7634;
	wire [4-1:0] node7637;
	wire [4-1:0] node7638;
	wire [4-1:0] node7642;
	wire [4-1:0] node7643;
	wire [4-1:0] node7644;
	wire [4-1:0] node7647;
	wire [4-1:0] node7651;
	wire [4-1:0] node7652;
	wire [4-1:0] node7653;
	wire [4-1:0] node7654;
	wire [4-1:0] node7657;
	wire [4-1:0] node7660;
	wire [4-1:0] node7663;
	wire [4-1:0] node7664;
	wire [4-1:0] node7667;
	wire [4-1:0] node7670;
	wire [4-1:0] node7671;
	wire [4-1:0] node7672;
	wire [4-1:0] node7673;
	wire [4-1:0] node7674;
	wire [4-1:0] node7677;
	wire [4-1:0] node7680;
	wire [4-1:0] node7683;
	wire [4-1:0] node7684;
	wire [4-1:0] node7688;
	wire [4-1:0] node7689;
	wire [4-1:0] node7692;
	wire [4-1:0] node7693;
	wire [4-1:0] node7696;
	wire [4-1:0] node7699;
	wire [4-1:0] node7700;
	wire [4-1:0] node7701;
	wire [4-1:0] node7702;
	wire [4-1:0] node7703;
	wire [4-1:0] node7704;
	wire [4-1:0] node7708;
	wire [4-1:0] node7709;
	wire [4-1:0] node7712;
	wire [4-1:0] node7715;
	wire [4-1:0] node7716;
	wire [4-1:0] node7717;
	wire [4-1:0] node7720;
	wire [4-1:0] node7724;
	wire [4-1:0] node7725;
	wire [4-1:0] node7726;
	wire [4-1:0] node7728;
	wire [4-1:0] node7733;
	wire [4-1:0] node7734;
	wire [4-1:0] node7735;
	wire [4-1:0] node7737;
	wire [4-1:0] node7740;
	wire [4-1:0] node7742;
	wire [4-1:0] node7745;
	wire [4-1:0] node7746;
	wire [4-1:0] node7748;
	wire [4-1:0] node7749;
	wire [4-1:0] node7753;
	wire [4-1:0] node7754;
	wire [4-1:0] node7755;
	wire [4-1:0] node7758;
	wire [4-1:0] node7762;
	wire [4-1:0] node7763;
	wire [4-1:0] node7764;
	wire [4-1:0] node7765;
	wire [4-1:0] node7766;
	wire [4-1:0] node7767;
	wire [4-1:0] node7768;
	wire [4-1:0] node7771;
	wire [4-1:0] node7775;
	wire [4-1:0] node7776;
	wire [4-1:0] node7779;
	wire [4-1:0] node7782;
	wire [4-1:0] node7783;
	wire [4-1:0] node7784;
	wire [4-1:0] node7785;
	wire [4-1:0] node7789;
	wire [4-1:0] node7792;
	wire [4-1:0] node7793;
	wire [4-1:0] node7795;
	wire [4-1:0] node7798;
	wire [4-1:0] node7799;
	wire [4-1:0] node7802;
	wire [4-1:0] node7805;
	wire [4-1:0] node7806;
	wire [4-1:0] node7807;
	wire [4-1:0] node7808;
	wire [4-1:0] node7809;
	wire [4-1:0] node7814;
	wire [4-1:0] node7815;
	wire [4-1:0] node7818;
	wire [4-1:0] node7821;
	wire [4-1:0] node7822;
	wire [4-1:0] node7823;
	wire [4-1:0] node7827;
	wire [4-1:0] node7828;
	wire [4-1:0] node7830;
	wire [4-1:0] node7833;
	wire [4-1:0] node7834;
	wire [4-1:0] node7837;
	wire [4-1:0] node7840;
	wire [4-1:0] node7841;
	wire [4-1:0] node7842;
	wire [4-1:0] node7843;
	wire [4-1:0] node7844;
	wire [4-1:0] node7846;
	wire [4-1:0] node7849;
	wire [4-1:0] node7852;
	wire [4-1:0] node7855;
	wire [4-1:0] node7856;
	wire [4-1:0] node7857;
	wire [4-1:0] node7860;
	wire [4-1:0] node7861;
	wire [4-1:0] node7864;
	wire [4-1:0] node7867;
	wire [4-1:0] node7870;
	wire [4-1:0] node7871;
	wire [4-1:0] node7872;
	wire [4-1:0] node7874;
	wire [4-1:0] node7876;
	wire [4-1:0] node7880;
	wire [4-1:0] node7881;
	wire [4-1:0] node7882;
	wire [4-1:0] node7885;
	wire [4-1:0] node7888;
	wire [4-1:0] node7890;
	wire [4-1:0] node7893;
	wire [4-1:0] node7894;
	wire [4-1:0] node7895;
	wire [4-1:0] node7896;
	wire [4-1:0] node7897;
	wire [4-1:0] node7898;
	wire [4-1:0] node7899;
	wire [4-1:0] node7900;
	wire [4-1:0] node7903;
	wire [4-1:0] node7906;
	wire [4-1:0] node7907;
	wire [4-1:0] node7910;
	wire [4-1:0] node7913;
	wire [4-1:0] node7914;
	wire [4-1:0] node7915;
	wire [4-1:0] node7918;
	wire [4-1:0] node7922;
	wire [4-1:0] node7923;
	wire [4-1:0] node7924;
	wire [4-1:0] node7927;
	wire [4-1:0] node7929;
	wire [4-1:0] node7932;
	wire [4-1:0] node7933;
	wire [4-1:0] node7934;
	wire [4-1:0] node7937;
	wire [4-1:0] node7941;
	wire [4-1:0] node7942;
	wire [4-1:0] node7943;
	wire [4-1:0] node7944;
	wire [4-1:0] node7945;
	wire [4-1:0] node7950;
	wire [4-1:0] node7951;
	wire [4-1:0] node7954;
	wire [4-1:0] node7957;
	wire [4-1:0] node7958;
	wire [4-1:0] node7960;
	wire [4-1:0] node7961;
	wire [4-1:0] node7965;
	wire [4-1:0] node7968;
	wire [4-1:0] node7969;
	wire [4-1:0] node7970;
	wire [4-1:0] node7971;
	wire [4-1:0] node7973;
	wire [4-1:0] node7974;
	wire [4-1:0] node7978;
	wire [4-1:0] node7980;
	wire [4-1:0] node7983;
	wire [4-1:0] node7984;
	wire [4-1:0] node7986;
	wire [4-1:0] node7989;
	wire [4-1:0] node7990;
	wire [4-1:0] node7994;
	wire [4-1:0] node7995;
	wire [4-1:0] node7996;
	wire [4-1:0] node7999;
	wire [4-1:0] node8000;
	wire [4-1:0] node8003;
	wire [4-1:0] node8006;
	wire [4-1:0] node8007;
	wire [4-1:0] node8008;
	wire [4-1:0] node8011;
	wire [4-1:0] node8012;
	wire [4-1:0] node8016;
	wire [4-1:0] node8017;
	wire [4-1:0] node8021;
	wire [4-1:0] node8022;
	wire [4-1:0] node8023;
	wire [4-1:0] node8024;
	wire [4-1:0] node8025;
	wire [4-1:0] node8027;
	wire [4-1:0] node8028;
	wire [4-1:0] node8032;
	wire [4-1:0] node8033;
	wire [4-1:0] node8036;
	wire [4-1:0] node8037;
	wire [4-1:0] node8040;
	wire [4-1:0] node8043;
	wire [4-1:0] node8044;
	wire [4-1:0] node8046;
	wire [4-1:0] node8047;
	wire [4-1:0] node8050;
	wire [4-1:0] node8053;
	wire [4-1:0] node8056;
	wire [4-1:0] node8057;
	wire [4-1:0] node8058;
	wire [4-1:0] node8059;
	wire [4-1:0] node8063;
	wire [4-1:0] node8064;
	wire [4-1:0] node8067;
	wire [4-1:0] node8070;
	wire [4-1:0] node8071;
	wire [4-1:0] node8072;
	wire [4-1:0] node8075;
	wire [4-1:0] node8078;
	wire [4-1:0] node8079;
	wire [4-1:0] node8083;
	wire [4-1:0] node8084;
	wire [4-1:0] node8085;
	wire [4-1:0] node8086;
	wire [4-1:0] node8087;
	wire [4-1:0] node8089;
	wire [4-1:0] node8092;
	wire [4-1:0] node8093;
	wire [4-1:0] node8096;
	wire [4-1:0] node8099;
	wire [4-1:0] node8100;
	wire [4-1:0] node8103;
	wire [4-1:0] node8106;
	wire [4-1:0] node8107;
	wire [4-1:0] node8108;
	wire [4-1:0] node8109;
	wire [4-1:0] node8113;
	wire [4-1:0] node8114;
	wire [4-1:0] node8117;
	wire [4-1:0] node8120;
	wire [4-1:0] node8122;
	wire [4-1:0] node8123;
	wire [4-1:0] node8127;
	wire [4-1:0] node8128;
	wire [4-1:0] node8129;
	wire [4-1:0] node8130;
	wire [4-1:0] node8131;
	wire [4-1:0] node8134;
	wire [4-1:0] node8137;
	wire [4-1:0] node8138;
	wire [4-1:0] node8141;
	wire [4-1:0] node8144;
	wire [4-1:0] node8145;
	wire [4-1:0] node8149;
	wire [4-1:0] node8150;
	wire [4-1:0] node8151;
	wire [4-1:0] node8154;
	wire [4-1:0] node8157;
	wire [4-1:0] node8159;
	wire [4-1:0] node8162;
	wire [4-1:0] node8163;
	wire [4-1:0] node8164;
	wire [4-1:0] node8165;
	wire [4-1:0] node8166;
	wire [4-1:0] node8167;
	wire [4-1:0] node8168;
	wire [4-1:0] node8169;
	wire [4-1:0] node8170;
	wire [4-1:0] node8174;
	wire [4-1:0] node8176;
	wire [4-1:0] node8180;
	wire [4-1:0] node8181;
	wire [4-1:0] node8182;
	wire [4-1:0] node8183;
	wire [4-1:0] node8186;
	wire [4-1:0] node8189;
	wire [4-1:0] node8190;
	wire [4-1:0] node8194;
	wire [4-1:0] node8196;
	wire [4-1:0] node8199;
	wire [4-1:0] node8200;
	wire [4-1:0] node8201;
	wire [4-1:0] node8203;
	wire [4-1:0] node8205;
	wire [4-1:0] node8208;
	wire [4-1:0] node8209;
	wire [4-1:0] node8212;
	wire [4-1:0] node8215;
	wire [4-1:0] node8216;
	wire [4-1:0] node8217;
	wire [4-1:0] node8218;
	wire [4-1:0] node8222;
	wire [4-1:0] node8225;
	wire [4-1:0] node8226;
	wire [4-1:0] node8229;
	wire [4-1:0] node8232;
	wire [4-1:0] node8233;
	wire [4-1:0] node8234;
	wire [4-1:0] node8235;
	wire [4-1:0] node8236;
	wire [4-1:0] node8237;
	wire [4-1:0] node8240;
	wire [4-1:0] node8243;
	wire [4-1:0] node8244;
	wire [4-1:0] node8247;
	wire [4-1:0] node8250;
	wire [4-1:0] node8251;
	wire [4-1:0] node8252;
	wire [4-1:0] node8256;
	wire [4-1:0] node8258;
	wire [4-1:0] node8261;
	wire [4-1:0] node8262;
	wire [4-1:0] node8263;
	wire [4-1:0] node8265;
	wire [4-1:0] node8269;
	wire [4-1:0] node8270;
	wire [4-1:0] node8273;
	wire [4-1:0] node8274;
	wire [4-1:0] node8278;
	wire [4-1:0] node8279;
	wire [4-1:0] node8280;
	wire [4-1:0] node8282;
	wire [4-1:0] node8285;
	wire [4-1:0] node8286;
	wire [4-1:0] node8287;
	wire [4-1:0] node8290;
	wire [4-1:0] node8294;
	wire [4-1:0] node8295;
	wire [4-1:0] node8296;
	wire [4-1:0] node8298;
	wire [4-1:0] node8301;
	wire [4-1:0] node8302;
	wire [4-1:0] node8306;
	wire [4-1:0] node8307;
	wire [4-1:0] node8308;
	wire [4-1:0] node8311;
	wire [4-1:0] node8315;
	wire [4-1:0] node8316;
	wire [4-1:0] node8317;
	wire [4-1:0] node8318;
	wire [4-1:0] node8319;
	wire [4-1:0] node8321;
	wire [4-1:0] node8324;
	wire [4-1:0] node8326;
	wire [4-1:0] node8329;
	wire [4-1:0] node8330;
	wire [4-1:0] node8331;
	wire [4-1:0] node8333;
	wire [4-1:0] node8336;
	wire [4-1:0] node8337;
	wire [4-1:0] node8340;
	wire [4-1:0] node8343;
	wire [4-1:0] node8345;
	wire [4-1:0] node8348;
	wire [4-1:0] node8349;
	wire [4-1:0] node8350;
	wire [4-1:0] node8351;
	wire [4-1:0] node8352;
	wire [4-1:0] node8355;
	wire [4-1:0] node8358;
	wire [4-1:0] node8360;
	wire [4-1:0] node8363;
	wire [4-1:0] node8364;
	wire [4-1:0] node8367;
	wire [4-1:0] node8370;
	wire [4-1:0] node8371;
	wire [4-1:0] node8375;
	wire [4-1:0] node8376;
	wire [4-1:0] node8377;
	wire [4-1:0] node8378;
	wire [4-1:0] node8379;
	wire [4-1:0] node8380;
	wire [4-1:0] node8385;
	wire [4-1:0] node8386;
	wire [4-1:0] node8387;
	wire [4-1:0] node8390;
	wire [4-1:0] node8394;
	wire [4-1:0] node8395;
	wire [4-1:0] node8396;
	wire [4-1:0] node8397;
	wire [4-1:0] node8400;
	wire [4-1:0] node8404;
	wire [4-1:0] node8405;
	wire [4-1:0] node8409;
	wire [4-1:0] node8410;
	wire [4-1:0] node8411;
	wire [4-1:0] node8412;
	wire [4-1:0] node8415;
	wire [4-1:0] node8418;
	wire [4-1:0] node8419;
	wire [4-1:0] node8422;
	wire [4-1:0] node8425;
	wire [4-1:0] node8426;
	wire [4-1:0] node8427;
	wire [4-1:0] node8430;
	wire [4-1:0] node8433;
	wire [4-1:0] node8434;
	wire [4-1:0] node8438;
	wire [4-1:0] node8439;
	wire [4-1:0] node8440;
	wire [4-1:0] node8441;
	wire [4-1:0] node8442;
	wire [4-1:0] node8443;
	wire [4-1:0] node8444;
	wire [4-1:0] node8448;
	wire [4-1:0] node8450;
	wire [4-1:0] node8451;
	wire [4-1:0] node8454;
	wire [4-1:0] node8457;
	wire [4-1:0] node8458;
	wire [4-1:0] node8460;
	wire [4-1:0] node8461;
	wire [4-1:0] node8465;
	wire [4-1:0] node8466;
	wire [4-1:0] node8467;
	wire [4-1:0] node8470;
	wire [4-1:0] node8473;
	wire [4-1:0] node8475;
	wire [4-1:0] node8478;
	wire [4-1:0] node8479;
	wire [4-1:0] node8480;
	wire [4-1:0] node8481;
	wire [4-1:0] node8485;
	wire [4-1:0] node8486;
	wire [4-1:0] node8489;
	wire [4-1:0] node8492;
	wire [4-1:0] node8493;
	wire [4-1:0] node8495;
	wire [4-1:0] node8498;
	wire [4-1:0] node8499;
	wire [4-1:0] node8502;
	wire [4-1:0] node8505;
	wire [4-1:0] node8506;
	wire [4-1:0] node8507;
	wire [4-1:0] node8508;
	wire [4-1:0] node8509;
	wire [4-1:0] node8510;
	wire [4-1:0] node8514;
	wire [4-1:0] node8515;
	wire [4-1:0] node8518;
	wire [4-1:0] node8521;
	wire [4-1:0] node8522;
	wire [4-1:0] node8523;
	wire [4-1:0] node8527;
	wire [4-1:0] node8529;
	wire [4-1:0] node8532;
	wire [4-1:0] node8533;
	wire [4-1:0] node8535;
	wire [4-1:0] node8536;
	wire [4-1:0] node8540;
	wire [4-1:0] node8541;
	wire [4-1:0] node8544;
	wire [4-1:0] node8547;
	wire [4-1:0] node8548;
	wire [4-1:0] node8549;
	wire [4-1:0] node8550;
	wire [4-1:0] node8552;
	wire [4-1:0] node8555;
	wire [4-1:0] node8556;
	wire [4-1:0] node8559;
	wire [4-1:0] node8562;
	wire [4-1:0] node8563;
	wire [4-1:0] node8566;
	wire [4-1:0] node8569;
	wire [4-1:0] node8570;
	wire [4-1:0] node8573;
	wire [4-1:0] node8574;
	wire [4-1:0] node8577;
	wire [4-1:0] node8580;
	wire [4-1:0] node8581;
	wire [4-1:0] node8582;
	wire [4-1:0] node8583;
	wire [4-1:0] node8584;
	wire [4-1:0] node8585;
	wire [4-1:0] node8586;
	wire [4-1:0] node8589;
	wire [4-1:0] node8592;
	wire [4-1:0] node8593;
	wire [4-1:0] node8596;
	wire [4-1:0] node8599;
	wire [4-1:0] node8600;
	wire [4-1:0] node8602;
	wire [4-1:0] node8606;
	wire [4-1:0] node8607;
	wire [4-1:0] node8608;
	wire [4-1:0] node8609;
	wire [4-1:0] node8612;
	wire [4-1:0] node8615;
	wire [4-1:0] node8618;
	wire [4-1:0] node8619;
	wire [4-1:0] node8622;
	wire [4-1:0] node8625;
	wire [4-1:0] node8626;
	wire [4-1:0] node8627;
	wire [4-1:0] node8628;
	wire [4-1:0] node8631;
	wire [4-1:0] node8633;
	wire [4-1:0] node8636;
	wire [4-1:0] node8637;
	wire [4-1:0] node8638;
	wire [4-1:0] node8643;
	wire [4-1:0] node8644;
	wire [4-1:0] node8645;
	wire [4-1:0] node8646;
	wire [4-1:0] node8650;
	wire [4-1:0] node8651;
	wire [4-1:0] node8655;
	wire [4-1:0] node8657;
	wire [4-1:0] node8659;
	wire [4-1:0] node8662;
	wire [4-1:0] node8663;
	wire [4-1:0] node8664;
	wire [4-1:0] node8665;
	wire [4-1:0] node8666;
	wire [4-1:0] node8667;
	wire [4-1:0] node8671;
	wire [4-1:0] node8674;
	wire [4-1:0] node8675;
	wire [4-1:0] node8676;
	wire [4-1:0] node8681;
	wire [4-1:0] node8682;
	wire [4-1:0] node8683;
	wire [4-1:0] node8687;
	wire [4-1:0] node8689;
	wire [4-1:0] node8690;
	wire [4-1:0] node8694;
	wire [4-1:0] node8695;
	wire [4-1:0] node8696;
	wire [4-1:0] node8698;
	wire [4-1:0] node8701;
	wire [4-1:0] node8702;
	wire [4-1:0] node8705;
	wire [4-1:0] node8708;
	wire [4-1:0] node8709;
	wire [4-1:0] node8710;
	wire [4-1:0] node8711;
	wire [4-1:0] node8714;
	wire [4-1:0] node8718;
	wire [4-1:0] node8719;
	wire [4-1:0] node8722;
	wire [4-1:0] node8725;
	wire [4-1:0] node8726;
	wire [4-1:0] node8727;
	wire [4-1:0] node8728;
	wire [4-1:0] node8729;
	wire [4-1:0] node8730;
	wire [4-1:0] node8731;
	wire [4-1:0] node8732;
	wire [4-1:0] node8733;
	wire [4-1:0] node8734;
	wire [4-1:0] node8736;
	wire [4-1:0] node8739;
	wire [4-1:0] node8740;
	wire [4-1:0] node8743;
	wire [4-1:0] node8746;
	wire [4-1:0] node8747;
	wire [4-1:0] node8751;
	wire [4-1:0] node8752;
	wire [4-1:0] node8753;
	wire [4-1:0] node8757;
	wire [4-1:0] node8758;
	wire [4-1:0] node8759;
	wire [4-1:0] node8762;
	wire [4-1:0] node8766;
	wire [4-1:0] node8767;
	wire [4-1:0] node8768;
	wire [4-1:0] node8769;
	wire [4-1:0] node8771;
	wire [4-1:0] node8775;
	wire [4-1:0] node8776;
	wire [4-1:0] node8779;
	wire [4-1:0] node8782;
	wire [4-1:0] node8783;
	wire [4-1:0] node8784;
	wire [4-1:0] node8786;
	wire [4-1:0] node8790;
	wire [4-1:0] node8791;
	wire [4-1:0] node8792;
	wire [4-1:0] node8795;
	wire [4-1:0] node8798;
	wire [4-1:0] node8800;
	wire [4-1:0] node8803;
	wire [4-1:0] node8804;
	wire [4-1:0] node8805;
	wire [4-1:0] node8806;
	wire [4-1:0] node8807;
	wire [4-1:0] node8809;
	wire [4-1:0] node8812;
	wire [4-1:0] node8814;
	wire [4-1:0] node8817;
	wire [4-1:0] node8818;
	wire [4-1:0] node8822;
	wire [4-1:0] node8823;
	wire [4-1:0] node8824;
	wire [4-1:0] node8825;
	wire [4-1:0] node8828;
	wire [4-1:0] node8831;
	wire [4-1:0] node8832;
	wire [4-1:0] node8835;
	wire [4-1:0] node8838;
	wire [4-1:0] node8839;
	wire [4-1:0] node8842;
	wire [4-1:0] node8845;
	wire [4-1:0] node8846;
	wire [4-1:0] node8847;
	wire [4-1:0] node8848;
	wire [4-1:0] node8850;
	wire [4-1:0] node8854;
	wire [4-1:0] node8855;
	wire [4-1:0] node8858;
	wire [4-1:0] node8861;
	wire [4-1:0] node8862;
	wire [4-1:0] node8863;
	wire [4-1:0] node8866;
	wire [4-1:0] node8870;
	wire [4-1:0] node8871;
	wire [4-1:0] node8872;
	wire [4-1:0] node8873;
	wire [4-1:0] node8875;
	wire [4-1:0] node8877;
	wire [4-1:0] node8879;
	wire [4-1:0] node8882;
	wire [4-1:0] node8884;
	wire [4-1:0] node8885;
	wire [4-1:0] node8888;
	wire [4-1:0] node8891;
	wire [4-1:0] node8892;
	wire [4-1:0] node8893;
	wire [4-1:0] node8894;
	wire [4-1:0] node8897;
	wire [4-1:0] node8900;
	wire [4-1:0] node8901;
	wire [4-1:0] node8904;
	wire [4-1:0] node8907;
	wire [4-1:0] node8908;
	wire [4-1:0] node8910;
	wire [4-1:0] node8913;
	wire [4-1:0] node8914;
	wire [4-1:0] node8916;
	wire [4-1:0] node8920;
	wire [4-1:0] node8921;
	wire [4-1:0] node8922;
	wire [4-1:0] node8923;
	wire [4-1:0] node8927;
	wire [4-1:0] node8928;
	wire [4-1:0] node8930;
	wire [4-1:0] node8931;
	wire [4-1:0] node8934;
	wire [4-1:0] node8937;
	wire [4-1:0] node8939;
	wire [4-1:0] node8942;
	wire [4-1:0] node8943;
	wire [4-1:0] node8944;
	wire [4-1:0] node8945;
	wire [4-1:0] node8948;
	wire [4-1:0] node8949;
	wire [4-1:0] node8953;
	wire [4-1:0] node8954;
	wire [4-1:0] node8955;
	wire [4-1:0] node8960;
	wire [4-1:0] node8961;
	wire [4-1:0] node8962;
	wire [4-1:0] node8963;
	wire [4-1:0] node8967;
	wire [4-1:0] node8968;
	wire [4-1:0] node8971;
	wire [4-1:0] node8974;
	wire [4-1:0] node8976;
	wire [4-1:0] node8979;
	wire [4-1:0] node8980;
	wire [4-1:0] node8981;
	wire [4-1:0] node8982;
	wire [4-1:0] node8983;
	wire [4-1:0] node8984;
	wire [4-1:0] node8986;
	wire [4-1:0] node8989;
	wire [4-1:0] node8990;
	wire [4-1:0] node8991;
	wire [4-1:0] node8994;
	wire [4-1:0] node8998;
	wire [4-1:0] node8999;
	wire [4-1:0] node9000;
	wire [4-1:0] node9003;
	wire [4-1:0] node9006;
	wire [4-1:0] node9007;
	wire [4-1:0] node9008;
	wire [4-1:0] node9011;
	wire [4-1:0] node9015;
	wire [4-1:0] node9016;
	wire [4-1:0] node9017;
	wire [4-1:0] node9018;
	wire [4-1:0] node9020;
	wire [4-1:0] node9023;
	wire [4-1:0] node9026;
	wire [4-1:0] node9027;
	wire [4-1:0] node9029;
	wire [4-1:0] node9032;
	wire [4-1:0] node9035;
	wire [4-1:0] node9036;
	wire [4-1:0] node9037;
	wire [4-1:0] node9038;
	wire [4-1:0] node9042;
	wire [4-1:0] node9043;
	wire [4-1:0] node9047;
	wire [4-1:0] node9049;
	wire [4-1:0] node9052;
	wire [4-1:0] node9053;
	wire [4-1:0] node9054;
	wire [4-1:0] node9055;
	wire [4-1:0] node9056;
	wire [4-1:0] node9058;
	wire [4-1:0] node9061;
	wire [4-1:0] node9062;
	wire [4-1:0] node9066;
	wire [4-1:0] node9067;
	wire [4-1:0] node9068;
	wire [4-1:0] node9071;
	wire [4-1:0] node9075;
	wire [4-1:0] node9076;
	wire [4-1:0] node9077;
	wire [4-1:0] node9081;
	wire [4-1:0] node9083;
	wire [4-1:0] node9084;
	wire [4-1:0] node9087;
	wire [4-1:0] node9090;
	wire [4-1:0] node9091;
	wire [4-1:0] node9092;
	wire [4-1:0] node9093;
	wire [4-1:0] node9096;
	wire [4-1:0] node9098;
	wire [4-1:0] node9101;
	wire [4-1:0] node9104;
	wire [4-1:0] node9106;
	wire [4-1:0] node9107;
	wire [4-1:0] node9110;
	wire [4-1:0] node9111;
	wire [4-1:0] node9115;
	wire [4-1:0] node9116;
	wire [4-1:0] node9117;
	wire [4-1:0] node9118;
	wire [4-1:0] node9119;
	wire [4-1:0] node9123;
	wire [4-1:0] node9124;
	wire [4-1:0] node9125;
	wire [4-1:0] node9128;
	wire [4-1:0] node9131;
	wire [4-1:0] node9133;
	wire [4-1:0] node9136;
	wire [4-1:0] node9137;
	wire [4-1:0] node9139;
	wire [4-1:0] node9141;
	wire [4-1:0] node9144;
	wire [4-1:0] node9145;
	wire [4-1:0] node9149;
	wire [4-1:0] node9150;
	wire [4-1:0] node9151;
	wire [4-1:0] node9152;
	wire [4-1:0] node9153;
	wire [4-1:0] node9156;
	wire [4-1:0] node9159;
	wire [4-1:0] node9160;
	wire [4-1:0] node9163;
	wire [4-1:0] node9166;
	wire [4-1:0] node9167;
	wire [4-1:0] node9169;
	wire [4-1:0] node9172;
	wire [4-1:0] node9175;
	wire [4-1:0] node9176;
	wire [4-1:0] node9177;
	wire [4-1:0] node9180;
	wire [4-1:0] node9182;
	wire [4-1:0] node9185;
	wire [4-1:0] node9186;
	wire [4-1:0] node9187;
	wire [4-1:0] node9191;
	wire [4-1:0] node9192;
	wire [4-1:0] node9195;
	wire [4-1:0] node9198;
	wire [4-1:0] node9199;
	wire [4-1:0] node9200;
	wire [4-1:0] node9201;
	wire [4-1:0] node9202;
	wire [4-1:0] node9203;
	wire [4-1:0] node9204;
	wire [4-1:0] node9205;
	wire [4-1:0] node9209;
	wire [4-1:0] node9210;
	wire [4-1:0] node9211;
	wire [4-1:0] node9214;
	wire [4-1:0] node9217;
	wire [4-1:0] node9218;
	wire [4-1:0] node9222;
	wire [4-1:0] node9224;
	wire [4-1:0] node9226;
	wire [4-1:0] node9227;
	wire [4-1:0] node9231;
	wire [4-1:0] node9232;
	wire [4-1:0] node9233;
	wire [4-1:0] node9235;
	wire [4-1:0] node9238;
	wire [4-1:0] node9240;
	wire [4-1:0] node9243;
	wire [4-1:0] node9244;
	wire [4-1:0] node9247;
	wire [4-1:0] node9249;
	wire [4-1:0] node9252;
	wire [4-1:0] node9253;
	wire [4-1:0] node9254;
	wire [4-1:0] node9255;
	wire [4-1:0] node9257;
	wire [4-1:0] node9260;
	wire [4-1:0] node9262;
	wire [4-1:0] node9265;
	wire [4-1:0] node9266;
	wire [4-1:0] node9268;
	wire [4-1:0] node9272;
	wire [4-1:0] node9273;
	wire [4-1:0] node9274;
	wire [4-1:0] node9276;
	wire [4-1:0] node9279;
	wire [4-1:0] node9280;
	wire [4-1:0] node9284;
	wire [4-1:0] node9285;
	wire [4-1:0] node9286;
	wire [4-1:0] node9290;
	wire [4-1:0] node9291;
	wire [4-1:0] node9295;
	wire [4-1:0] node9296;
	wire [4-1:0] node9297;
	wire [4-1:0] node9298;
	wire [4-1:0] node9299;
	wire [4-1:0] node9301;
	wire [4-1:0] node9304;
	wire [4-1:0] node9306;
	wire [4-1:0] node9308;
	wire [4-1:0] node9311;
	wire [4-1:0] node9312;
	wire [4-1:0] node9313;
	wire [4-1:0] node9314;
	wire [4-1:0] node9317;
	wire [4-1:0] node9321;
	wire [4-1:0] node9322;
	wire [4-1:0] node9326;
	wire [4-1:0] node9327;
	wire [4-1:0] node9328;
	wire [4-1:0] node9330;
	wire [4-1:0] node9333;
	wire [4-1:0] node9334;
	wire [4-1:0] node9335;
	wire [4-1:0] node9338;
	wire [4-1:0] node9341;
	wire [4-1:0] node9342;
	wire [4-1:0] node9346;
	wire [4-1:0] node9347;
	wire [4-1:0] node9348;
	wire [4-1:0] node9349;
	wire [4-1:0] node9354;
	wire [4-1:0] node9355;
	wire [4-1:0] node9359;
	wire [4-1:0] node9360;
	wire [4-1:0] node9361;
	wire [4-1:0] node9362;
	wire [4-1:0] node9363;
	wire [4-1:0] node9365;
	wire [4-1:0] node9368;
	wire [4-1:0] node9371;
	wire [4-1:0] node9372;
	wire [4-1:0] node9375;
	wire [4-1:0] node9377;
	wire [4-1:0] node9380;
	wire [4-1:0] node9381;
	wire [4-1:0] node9382;
	wire [4-1:0] node9383;
	wire [4-1:0] node9387;
	wire [4-1:0] node9388;
	wire [4-1:0] node9392;
	wire [4-1:0] node9393;
	wire [4-1:0] node9394;
	wire [4-1:0] node9397;
	wire [4-1:0] node9401;
	wire [4-1:0] node9402;
	wire [4-1:0] node9403;
	wire [4-1:0] node9404;
	wire [4-1:0] node9406;
	wire [4-1:0] node9409;
	wire [4-1:0] node9411;
	wire [4-1:0] node9414;
	wire [4-1:0] node9417;
	wire [4-1:0] node9418;
	wire [4-1:0] node9419;
	wire [4-1:0] node9423;
	wire [4-1:0] node9424;
	wire [4-1:0] node9425;
	wire [4-1:0] node9430;
	wire [4-1:0] node9431;
	wire [4-1:0] node9432;
	wire [4-1:0] node9433;
	wire [4-1:0] node9434;
	wire [4-1:0] node9435;
	wire [4-1:0] node9436;
	wire [4-1:0] node9440;
	wire [4-1:0] node9441;
	wire [4-1:0] node9444;
	wire [4-1:0] node9447;
	wire [4-1:0] node9448;
	wire [4-1:0] node9449;
	wire [4-1:0] node9450;
	wire [4-1:0] node9453;
	wire [4-1:0] node9457;
	wire [4-1:0] node9458;
	wire [4-1:0] node9460;
	wire [4-1:0] node9464;
	wire [4-1:0] node9465;
	wire [4-1:0] node9466;
	wire [4-1:0] node9468;
	wire [4-1:0] node9471;
	wire [4-1:0] node9472;
	wire [4-1:0] node9476;
	wire [4-1:0] node9477;
	wire [4-1:0] node9480;
	wire [4-1:0] node9481;
	wire [4-1:0] node9484;
	wire [4-1:0] node9487;
	wire [4-1:0] node9488;
	wire [4-1:0] node9489;
	wire [4-1:0] node9490;
	wire [4-1:0] node9491;
	wire [4-1:0] node9494;
	wire [4-1:0] node9497;
	wire [4-1:0] node9498;
	wire [4-1:0] node9501;
	wire [4-1:0] node9504;
	wire [4-1:0] node9506;
	wire [4-1:0] node9507;
	wire [4-1:0] node9510;
	wire [4-1:0] node9513;
	wire [4-1:0] node9514;
	wire [4-1:0] node9515;
	wire [4-1:0] node9516;
	wire [4-1:0] node9519;
	wire [4-1:0] node9522;
	wire [4-1:0] node9523;
	wire [4-1:0] node9524;
	wire [4-1:0] node9528;
	wire [4-1:0] node9531;
	wire [4-1:0] node9532;
	wire [4-1:0] node9533;
	wire [4-1:0] node9536;
	wire [4-1:0] node9539;
	wire [4-1:0] node9540;
	wire [4-1:0] node9543;
	wire [4-1:0] node9546;
	wire [4-1:0] node9547;
	wire [4-1:0] node9548;
	wire [4-1:0] node9549;
	wire [4-1:0] node9550;
	wire [4-1:0] node9551;
	wire [4-1:0] node9554;
	wire [4-1:0] node9557;
	wire [4-1:0] node9559;
	wire [4-1:0] node9562;
	wire [4-1:0] node9563;
	wire [4-1:0] node9565;
	wire [4-1:0] node9568;
	wire [4-1:0] node9569;
	wire [4-1:0] node9572;
	wire [4-1:0] node9575;
	wire [4-1:0] node9576;
	wire [4-1:0] node9577;
	wire [4-1:0] node9578;
	wire [4-1:0] node9581;
	wire [4-1:0] node9584;
	wire [4-1:0] node9585;
	wire [4-1:0] node9587;
	wire [4-1:0] node9591;
	wire [4-1:0] node9592;
	wire [4-1:0] node9593;
	wire [4-1:0] node9596;
	wire [4-1:0] node9599;
	wire [4-1:0] node9600;
	wire [4-1:0] node9603;
	wire [4-1:0] node9606;
	wire [4-1:0] node9607;
	wire [4-1:0] node9608;
	wire [4-1:0] node9610;
	wire [4-1:0] node9611;
	wire [4-1:0] node9614;
	wire [4-1:0] node9617;
	wire [4-1:0] node9618;
	wire [4-1:0] node9620;
	wire [4-1:0] node9621;
	wire [4-1:0] node9624;
	wire [4-1:0] node9627;
	wire [4-1:0] node9628;
	wire [4-1:0] node9631;
	wire [4-1:0] node9634;
	wire [4-1:0] node9635;
	wire [4-1:0] node9637;
	wire [4-1:0] node9638;
	wire [4-1:0] node9641;
	wire [4-1:0] node9644;
	wire [4-1:0] node9647;
	wire [4-1:0] node9648;
	wire [4-1:0] node9649;
	wire [4-1:0] node9650;
	wire [4-1:0] node9651;
	wire [4-1:0] node9652;
	wire [4-1:0] node9653;
	wire [4-1:0] node9654;
	wire [4-1:0] node9655;
	wire [4-1:0] node9658;
	wire [4-1:0] node9661;
	wire [4-1:0] node9662;
	wire [4-1:0] node9665;
	wire [4-1:0] node9668;
	wire [4-1:0] node9669;
	wire [4-1:0] node9670;
	wire [4-1:0] node9673;
	wire [4-1:0] node9676;
	wire [4-1:0] node9677;
	wire [4-1:0] node9679;
	wire [4-1:0] node9683;
	wire [4-1:0] node9684;
	wire [4-1:0] node9685;
	wire [4-1:0] node9688;
	wire [4-1:0] node9690;
	wire [4-1:0] node9693;
	wire [4-1:0] node9694;
	wire [4-1:0] node9695;
	wire [4-1:0] node9698;
	wire [4-1:0] node9701;
	wire [4-1:0] node9702;
	wire [4-1:0] node9705;
	wire [4-1:0] node9708;
	wire [4-1:0] node9709;
	wire [4-1:0] node9710;
	wire [4-1:0] node9711;
	wire [4-1:0] node9714;
	wire [4-1:0] node9717;
	wire [4-1:0] node9718;
	wire [4-1:0] node9720;
	wire [4-1:0] node9723;
	wire [4-1:0] node9725;
	wire [4-1:0] node9727;
	wire [4-1:0] node9730;
	wire [4-1:0] node9731;
	wire [4-1:0] node9732;
	wire [4-1:0] node9736;
	wire [4-1:0] node9737;
	wire [4-1:0] node9739;
	wire [4-1:0] node9742;
	wire [4-1:0] node9743;
	wire [4-1:0] node9744;
	wire [4-1:0] node9747;
	wire [4-1:0] node9750;
	wire [4-1:0] node9751;
	wire [4-1:0] node9754;
	wire [4-1:0] node9757;
	wire [4-1:0] node9758;
	wire [4-1:0] node9759;
	wire [4-1:0] node9760;
	wire [4-1:0] node9761;
	wire [4-1:0] node9762;
	wire [4-1:0] node9765;
	wire [4-1:0] node9766;
	wire [4-1:0] node9770;
	wire [4-1:0] node9772;
	wire [4-1:0] node9775;
	wire [4-1:0] node9777;
	wire [4-1:0] node9778;
	wire [4-1:0] node9779;
	wire [4-1:0] node9783;
	wire [4-1:0] node9784;
	wire [4-1:0] node9787;
	wire [4-1:0] node9790;
	wire [4-1:0] node9791;
	wire [4-1:0] node9792;
	wire [4-1:0] node9793;
	wire [4-1:0] node9794;
	wire [4-1:0] node9798;
	wire [4-1:0] node9800;
	wire [4-1:0] node9803;
	wire [4-1:0] node9804;
	wire [4-1:0] node9805;
	wire [4-1:0] node9808;
	wire [4-1:0] node9812;
	wire [4-1:0] node9813;
	wire [4-1:0] node9814;
	wire [4-1:0] node9815;
	wire [4-1:0] node9820;
	wire [4-1:0] node9822;
	wire [4-1:0] node9823;
	wire [4-1:0] node9826;
	wire [4-1:0] node9829;
	wire [4-1:0] node9830;
	wire [4-1:0] node9831;
	wire [4-1:0] node9832;
	wire [4-1:0] node9833;
	wire [4-1:0] node9835;
	wire [4-1:0] node9838;
	wire [4-1:0] node9839;
	wire [4-1:0] node9842;
	wire [4-1:0] node9845;
	wire [4-1:0] node9846;
	wire [4-1:0] node9848;
	wire [4-1:0] node9852;
	wire [4-1:0] node9853;
	wire [4-1:0] node9854;
	wire [4-1:0] node9855;
	wire [4-1:0] node9858;
	wire [4-1:0] node9861;
	wire [4-1:0] node9862;
	wire [4-1:0] node9866;
	wire [4-1:0] node9867;
	wire [4-1:0] node9871;
	wire [4-1:0] node9872;
	wire [4-1:0] node9873;
	wire [4-1:0] node9874;
	wire [4-1:0] node9876;
	wire [4-1:0] node9880;
	wire [4-1:0] node9883;
	wire [4-1:0] node9884;
	wire [4-1:0] node9886;
	wire [4-1:0] node9887;
	wire [4-1:0] node9890;
	wire [4-1:0] node9893;
	wire [4-1:0] node9894;
	wire [4-1:0] node9896;
	wire [4-1:0] node9899;
	wire [4-1:0] node9901;
	wire [4-1:0] node9904;
	wire [4-1:0] node9905;
	wire [4-1:0] node9906;
	wire [4-1:0] node9907;
	wire [4-1:0] node9908;
	wire [4-1:0] node9909;
	wire [4-1:0] node9910;
	wire [4-1:0] node9912;
	wire [4-1:0] node9915;
	wire [4-1:0] node9917;
	wire [4-1:0] node9920;
	wire [4-1:0] node9922;
	wire [4-1:0] node9923;
	wire [4-1:0] node9927;
	wire [4-1:0] node9928;
	wire [4-1:0] node9930;
	wire [4-1:0] node9933;
	wire [4-1:0] node9935;
	wire [4-1:0] node9937;
	wire [4-1:0] node9940;
	wire [4-1:0] node9941;
	wire [4-1:0] node9942;
	wire [4-1:0] node9944;
	wire [4-1:0] node9945;
	wire [4-1:0] node9949;
	wire [4-1:0] node9950;
	wire [4-1:0] node9951;
	wire [4-1:0] node9955;
	wire [4-1:0] node9957;
	wire [4-1:0] node9960;
	wire [4-1:0] node9961;
	wire [4-1:0] node9962;
	wire [4-1:0] node9965;
	wire [4-1:0] node9966;
	wire [4-1:0] node9970;
	wire [4-1:0] node9972;
	wire [4-1:0] node9975;
	wire [4-1:0] node9976;
	wire [4-1:0] node9977;
	wire [4-1:0] node9978;
	wire [4-1:0] node9979;
	wire [4-1:0] node9980;
	wire [4-1:0] node9983;
	wire [4-1:0] node9986;
	wire [4-1:0] node9989;
	wire [4-1:0] node9990;
	wire [4-1:0] node9991;
	wire [4-1:0] node9994;
	wire [4-1:0] node9997;
	wire [4-1:0] node9998;
	wire [4-1:0] node10001;
	wire [4-1:0] node10004;
	wire [4-1:0] node10005;
	wire [4-1:0] node10006;
	wire [4-1:0] node10007;
	wire [4-1:0] node10011;
	wire [4-1:0] node10014;
	wire [4-1:0] node10015;
	wire [4-1:0] node10019;
	wire [4-1:0] node10020;
	wire [4-1:0] node10021;
	wire [4-1:0] node10022;
	wire [4-1:0] node10023;
	wire [4-1:0] node10026;
	wire [4-1:0] node10029;
	wire [4-1:0] node10030;
	wire [4-1:0] node10034;
	wire [4-1:0] node10036;
	wire [4-1:0] node10039;
	wire [4-1:0] node10040;
	wire [4-1:0] node10041;
	wire [4-1:0] node10042;
	wire [4-1:0] node10047;
	wire [4-1:0] node10048;
	wire [4-1:0] node10051;
	wire [4-1:0] node10054;
	wire [4-1:0] node10055;
	wire [4-1:0] node10056;
	wire [4-1:0] node10057;
	wire [4-1:0] node10058;
	wire [4-1:0] node10059;
	wire [4-1:0] node10060;
	wire [4-1:0] node10063;
	wire [4-1:0] node10066;
	wire [4-1:0] node10068;
	wire [4-1:0] node10071;
	wire [4-1:0] node10073;
	wire [4-1:0] node10076;
	wire [4-1:0] node10077;
	wire [4-1:0] node10078;
	wire [4-1:0] node10079;
	wire [4-1:0] node10082;
	wire [4-1:0] node10086;
	wire [4-1:0] node10088;
	wire [4-1:0] node10089;
	wire [4-1:0] node10093;
	wire [4-1:0] node10094;
	wire [4-1:0] node10095;
	wire [4-1:0] node10096;
	wire [4-1:0] node10099;
	wire [4-1:0] node10100;
	wire [4-1:0] node10103;
	wire [4-1:0] node10106;
	wire [4-1:0] node10108;
	wire [4-1:0] node10110;
	wire [4-1:0] node10113;
	wire [4-1:0] node10114;
	wire [4-1:0] node10115;
	wire [4-1:0] node10116;
	wire [4-1:0] node10119;
	wire [4-1:0] node10122;
	wire [4-1:0] node10123;
	wire [4-1:0] node10127;
	wire [4-1:0] node10128;
	wire [4-1:0] node10130;
	wire [4-1:0] node10133;
	wire [4-1:0] node10135;
	wire [4-1:0] node10138;
	wire [4-1:0] node10139;
	wire [4-1:0] node10140;
	wire [4-1:0] node10141;
	wire [4-1:0] node10142;
	wire [4-1:0] node10143;
	wire [4-1:0] node10147;
	wire [4-1:0] node10149;
	wire [4-1:0] node10152;
	wire [4-1:0] node10153;
	wire [4-1:0] node10154;
	wire [4-1:0] node10158;
	wire [4-1:0] node10159;
	wire [4-1:0] node10162;
	wire [4-1:0] node10165;
	wire [4-1:0] node10166;
	wire [4-1:0] node10167;
	wire [4-1:0] node10168;
	wire [4-1:0] node10172;
	wire [4-1:0] node10175;
	wire [4-1:0] node10176;
	wire [4-1:0] node10177;
	wire [4-1:0] node10182;
	wire [4-1:0] node10183;
	wire [4-1:0] node10184;
	wire [4-1:0] node10186;
	wire [4-1:0] node10188;
	wire [4-1:0] node10191;
	wire [4-1:0] node10192;
	wire [4-1:0] node10193;
	wire [4-1:0] node10196;
	wire [4-1:0] node10200;
	wire [4-1:0] node10201;
	wire [4-1:0] node10202;
	wire [4-1:0] node10204;
	wire [4-1:0] node10207;
	wire [4-1:0] node10209;
	wire [4-1:0] node10212;
	wire [4-1:0] node10214;
	wire [4-1:0] node10217;
	wire [4-1:0] node10218;
	wire [4-1:0] node10219;
	wire [4-1:0] node10220;
	wire [4-1:0] node10221;
	wire [4-1:0] node10222;
	wire [4-1:0] node10223;
	wire [4-1:0] node10224;
	wire [4-1:0] node10227;
	wire [4-1:0] node10230;
	wire [4-1:0] node10232;
	wire [4-1:0] node10233;
	wire [4-1:0] node10236;
	wire [4-1:0] node10239;
	wire [4-1:0] node10240;
	wire [4-1:0] node10241;
	wire [4-1:0] node10244;
	wire [4-1:0] node10247;
	wire [4-1:0] node10248;
	wire [4-1:0] node10249;
	wire [4-1:0] node10253;
	wire [4-1:0] node10255;
	wire [4-1:0] node10258;
	wire [4-1:0] node10259;
	wire [4-1:0] node10260;
	wire [4-1:0] node10261;
	wire [4-1:0] node10264;
	wire [4-1:0] node10267;
	wire [4-1:0] node10268;
	wire [4-1:0] node10269;
	wire [4-1:0] node10272;
	wire [4-1:0] node10275;
	wire [4-1:0] node10277;
	wire [4-1:0] node10280;
	wire [4-1:0] node10281;
	wire [4-1:0] node10282;
	wire [4-1:0] node10286;
	wire [4-1:0] node10287;
	wire [4-1:0] node10290;
	wire [4-1:0] node10293;
	wire [4-1:0] node10294;
	wire [4-1:0] node10295;
	wire [4-1:0] node10296;
	wire [4-1:0] node10297;
	wire [4-1:0] node10301;
	wire [4-1:0] node10302;
	wire [4-1:0] node10303;
	wire [4-1:0] node10307;
	wire [4-1:0] node10308;
	wire [4-1:0] node10312;
	wire [4-1:0] node10313;
	wire [4-1:0] node10315;
	wire [4-1:0] node10318;
	wire [4-1:0] node10319;
	wire [4-1:0] node10320;
	wire [4-1:0] node10324;
	wire [4-1:0] node10327;
	wire [4-1:0] node10328;
	wire [4-1:0] node10329;
	wire [4-1:0] node10330;
	wire [4-1:0] node10332;
	wire [4-1:0] node10335;
	wire [4-1:0] node10336;
	wire [4-1:0] node10339;
	wire [4-1:0] node10342;
	wire [4-1:0] node10343;
	wire [4-1:0] node10347;
	wire [4-1:0] node10348;
	wire [4-1:0] node10351;
	wire [4-1:0] node10352;
	wire [4-1:0] node10354;
	wire [4-1:0] node10358;
	wire [4-1:0] node10359;
	wire [4-1:0] node10360;
	wire [4-1:0] node10361;
	wire [4-1:0] node10362;
	wire [4-1:0] node10363;
	wire [4-1:0] node10366;
	wire [4-1:0] node10368;
	wire [4-1:0] node10371;
	wire [4-1:0] node10372;
	wire [4-1:0] node10376;
	wire [4-1:0] node10377;
	wire [4-1:0] node10379;
	wire [4-1:0] node10381;
	wire [4-1:0] node10384;
	wire [4-1:0] node10385;
	wire [4-1:0] node10388;
	wire [4-1:0] node10391;
	wire [4-1:0] node10392;
	wire [4-1:0] node10393;
	wire [4-1:0] node10394;
	wire [4-1:0] node10396;
	wire [4-1:0] node10400;
	wire [4-1:0] node10402;
	wire [4-1:0] node10405;
	wire [4-1:0] node10406;
	wire [4-1:0] node10407;
	wire [4-1:0] node10408;
	wire [4-1:0] node10411;
	wire [4-1:0] node10414;
	wire [4-1:0] node10415;
	wire [4-1:0] node10419;
	wire [4-1:0] node10421;
	wire [4-1:0] node10424;
	wire [4-1:0] node10425;
	wire [4-1:0] node10426;
	wire [4-1:0] node10427;
	wire [4-1:0] node10428;
	wire [4-1:0] node10429;
	wire [4-1:0] node10432;
	wire [4-1:0] node10435;
	wire [4-1:0] node10436;
	wire [4-1:0] node10440;
	wire [4-1:0] node10441;
	wire [4-1:0] node10444;
	wire [4-1:0] node10447;
	wire [4-1:0] node10448;
	wire [4-1:0] node10450;
	wire [4-1:0] node10453;
	wire [4-1:0] node10454;
	wire [4-1:0] node10457;
	wire [4-1:0] node10460;
	wire [4-1:0] node10461;
	wire [4-1:0] node10462;
	wire [4-1:0] node10464;
	wire [4-1:0] node10466;
	wire [4-1:0] node10469;
	wire [4-1:0] node10470;
	wire [4-1:0] node10471;
	wire [4-1:0] node10475;
	wire [4-1:0] node10478;
	wire [4-1:0] node10479;
	wire [4-1:0] node10482;
	wire [4-1:0] node10485;
	wire [4-1:0] node10486;
	wire [4-1:0] node10487;
	wire [4-1:0] node10488;
	wire [4-1:0] node10489;
	wire [4-1:0] node10490;
	wire [4-1:0] node10492;
	wire [4-1:0] node10493;
	wire [4-1:0] node10496;
	wire [4-1:0] node10499;
	wire [4-1:0] node10500;
	wire [4-1:0] node10503;
	wire [4-1:0] node10506;
	wire [4-1:0] node10507;
	wire [4-1:0] node10510;
	wire [4-1:0] node10512;
	wire [4-1:0] node10515;
	wire [4-1:0] node10516;
	wire [4-1:0] node10517;
	wire [4-1:0] node10520;
	wire [4-1:0] node10522;
	wire [4-1:0] node10525;
	wire [4-1:0] node10527;
	wire [4-1:0] node10528;
	wire [4-1:0] node10531;
	wire [4-1:0] node10532;
	wire [4-1:0] node10536;
	wire [4-1:0] node10537;
	wire [4-1:0] node10538;
	wire [4-1:0] node10539;
	wire [4-1:0] node10540;
	wire [4-1:0] node10544;
	wire [4-1:0] node10545;
	wire [4-1:0] node10548;
	wire [4-1:0] node10551;
	wire [4-1:0] node10552;
	wire [4-1:0] node10553;
	wire [4-1:0] node10556;
	wire [4-1:0] node10559;
	wire [4-1:0] node10560;
	wire [4-1:0] node10564;
	wire [4-1:0] node10565;
	wire [4-1:0] node10566;
	wire [4-1:0] node10567;
	wire [4-1:0] node10570;
	wire [4-1:0] node10573;
	wire [4-1:0] node10575;
	wire [4-1:0] node10577;
	wire [4-1:0] node10580;
	wire [4-1:0] node10581;
	wire [4-1:0] node10582;
	wire [4-1:0] node10587;
	wire [4-1:0] node10588;
	wire [4-1:0] node10589;
	wire [4-1:0] node10590;
	wire [4-1:0] node10591;
	wire [4-1:0] node10592;
	wire [4-1:0] node10595;
	wire [4-1:0] node10598;
	wire [4-1:0] node10600;
	wire [4-1:0] node10601;
	wire [4-1:0] node10604;
	wire [4-1:0] node10607;
	wire [4-1:0] node10608;
	wire [4-1:0] node10609;
	wire [4-1:0] node10613;
	wire [4-1:0] node10616;
	wire [4-1:0] node10617;
	wire [4-1:0] node10618;
	wire [4-1:0] node10619;
	wire [4-1:0] node10622;
	wire [4-1:0] node10625;
	wire [4-1:0] node10626;
	wire [4-1:0] node10629;
	wire [4-1:0] node10632;
	wire [4-1:0] node10633;
	wire [4-1:0] node10634;
	wire [4-1:0] node10637;
	wire [4-1:0] node10640;
	wire [4-1:0] node10641;
	wire [4-1:0] node10644;
	wire [4-1:0] node10647;
	wire [4-1:0] node10648;
	wire [4-1:0] node10649;
	wire [4-1:0] node10650;
	wire [4-1:0] node10652;
	wire [4-1:0] node10653;
	wire [4-1:0] node10657;
	wire [4-1:0] node10659;
	wire [4-1:0] node10660;
	wire [4-1:0] node10663;
	wire [4-1:0] node10666;
	wire [4-1:0] node10667;
	wire [4-1:0] node10669;
	wire [4-1:0] node10672;
	wire [4-1:0] node10673;
	wire [4-1:0] node10676;
	wire [4-1:0] node10677;
	wire [4-1:0] node10681;
	wire [4-1:0] node10682;
	wire [4-1:0] node10683;
	wire [4-1:0] node10684;
	wire [4-1:0] node10685;
	wire [4-1:0] node10690;
	wire [4-1:0] node10691;
	wire [4-1:0] node10694;
	wire [4-1:0] node10697;
	wire [4-1:0] node10698;
	wire [4-1:0] node10699;
	wire [4-1:0] node10702;
	wire [4-1:0] node10705;
	wire [4-1:0] node10706;
	wire [4-1:0] node10707;
	wire [4-1:0] node10710;
	wire [4-1:0] node10714;
	wire [4-1:0] node10715;
	wire [4-1:0] node10716;
	wire [4-1:0] node10717;
	wire [4-1:0] node10718;
	wire [4-1:0] node10719;
	wire [4-1:0] node10720;
	wire [4-1:0] node10721;
	wire [4-1:0] node10722;
	wire [4-1:0] node10723;
	wire [4-1:0] node10726;
	wire [4-1:0] node10728;
	wire [4-1:0] node10731;
	wire [4-1:0] node10732;
	wire [4-1:0] node10735;
	wire [4-1:0] node10737;
	wire [4-1:0] node10740;
	wire [4-1:0] node10741;
	wire [4-1:0] node10742;
	wire [4-1:0] node10743;
	wire [4-1:0] node10746;
	wire [4-1:0] node10749;
	wire [4-1:0] node10750;
	wire [4-1:0] node10753;
	wire [4-1:0] node10756;
	wire [4-1:0] node10757;
	wire [4-1:0] node10758;
	wire [4-1:0] node10762;
	wire [4-1:0] node10764;
	wire [4-1:0] node10766;
	wire [4-1:0] node10769;
	wire [4-1:0] node10770;
	wire [4-1:0] node10771;
	wire [4-1:0] node10772;
	wire [4-1:0] node10773;
	wire [4-1:0] node10777;
	wire [4-1:0] node10778;
	wire [4-1:0] node10781;
	wire [4-1:0] node10784;
	wire [4-1:0] node10785;
	wire [4-1:0] node10786;
	wire [4-1:0] node10789;
	wire [4-1:0] node10792;
	wire [4-1:0] node10793;
	wire [4-1:0] node10796;
	wire [4-1:0] node10799;
	wire [4-1:0] node10800;
	wire [4-1:0] node10801;
	wire [4-1:0] node10802;
	wire [4-1:0] node10805;
	wire [4-1:0] node10808;
	wire [4-1:0] node10809;
	wire [4-1:0] node10811;
	wire [4-1:0] node10814;
	wire [4-1:0] node10815;
	wire [4-1:0] node10818;
	wire [4-1:0] node10821;
	wire [4-1:0] node10822;
	wire [4-1:0] node10823;
	wire [4-1:0] node10826;
	wire [4-1:0] node10829;
	wire [4-1:0] node10831;
	wire [4-1:0] node10834;
	wire [4-1:0] node10835;
	wire [4-1:0] node10836;
	wire [4-1:0] node10837;
	wire [4-1:0] node10838;
	wire [4-1:0] node10839;
	wire [4-1:0] node10841;
	wire [4-1:0] node10844;
	wire [4-1:0] node10845;
	wire [4-1:0] node10849;
	wire [4-1:0] node10850;
	wire [4-1:0] node10854;
	wire [4-1:0] node10855;
	wire [4-1:0] node10857;
	wire [4-1:0] node10860;
	wire [4-1:0] node10862;
	wire [4-1:0] node10864;
	wire [4-1:0] node10867;
	wire [4-1:0] node10868;
	wire [4-1:0] node10870;
	wire [4-1:0] node10872;
	wire [4-1:0] node10875;
	wire [4-1:0] node10876;
	wire [4-1:0] node10878;
	wire [4-1:0] node10881;
	wire [4-1:0] node10882;
	wire [4-1:0] node10886;
	wire [4-1:0] node10887;
	wire [4-1:0] node10888;
	wire [4-1:0] node10889;
	wire [4-1:0] node10890;
	wire [4-1:0] node10891;
	wire [4-1:0] node10896;
	wire [4-1:0] node10898;
	wire [4-1:0] node10899;
	wire [4-1:0] node10903;
	wire [4-1:0] node10904;
	wire [4-1:0] node10905;
	wire [4-1:0] node10908;
	wire [4-1:0] node10911;
	wire [4-1:0] node10912;
	wire [4-1:0] node10915;
	wire [4-1:0] node10916;
	wire [4-1:0] node10920;
	wire [4-1:0] node10921;
	wire [4-1:0] node10922;
	wire [4-1:0] node10924;
	wire [4-1:0] node10927;
	wire [4-1:0] node10928;
	wire [4-1:0] node10929;
	wire [4-1:0] node10933;
	wire [4-1:0] node10936;
	wire [4-1:0] node10937;
	wire [4-1:0] node10939;
	wire [4-1:0] node10942;
	wire [4-1:0] node10943;
	wire [4-1:0] node10944;
	wire [4-1:0] node10947;
	wire [4-1:0] node10950;
	wire [4-1:0] node10951;
	wire [4-1:0] node10954;
	wire [4-1:0] node10957;
	wire [4-1:0] node10958;
	wire [4-1:0] node10959;
	wire [4-1:0] node10960;
	wire [4-1:0] node10961;
	wire [4-1:0] node10964;
	wire [4-1:0] node10967;
	wire [4-1:0] node10968;
	wire [4-1:0] node10969;
	wire [4-1:0] node10970;
	wire [4-1:0] node10973;
	wire [4-1:0] node10975;
	wire [4-1:0] node10978;
	wire [4-1:0] node10979;
	wire [4-1:0] node10982;
	wire [4-1:0] node10985;
	wire [4-1:0] node10986;
	wire [4-1:0] node10987;
	wire [4-1:0] node10990;
	wire [4-1:0] node10993;
	wire [4-1:0] node10994;
	wire [4-1:0] node10995;
	wire [4-1:0] node10999;
	wire [4-1:0] node11002;
	wire [4-1:0] node11003;
	wire [4-1:0] node11004;
	wire [4-1:0] node11005;
	wire [4-1:0] node11008;
	wire [4-1:0] node11011;
	wire [4-1:0] node11012;
	wire [4-1:0] node11014;
	wire [4-1:0] node11015;
	wire [4-1:0] node11018;
	wire [4-1:0] node11021;
	wire [4-1:0] node11022;
	wire [4-1:0] node11024;
	wire [4-1:0] node11027;
	wire [4-1:0] node11029;
	wire [4-1:0] node11032;
	wire [4-1:0] node11033;
	wire [4-1:0] node11034;
	wire [4-1:0] node11037;
	wire [4-1:0] node11039;
	wire [4-1:0] node11042;
	wire [4-1:0] node11043;
	wire [4-1:0] node11045;
	wire [4-1:0] node11048;
	wire [4-1:0] node11050;
	wire [4-1:0] node11053;
	wire [4-1:0] node11054;
	wire [4-1:0] node11055;
	wire [4-1:0] node11056;
	wire [4-1:0] node11057;
	wire [4-1:0] node11058;
	wire [4-1:0] node11061;
	wire [4-1:0] node11064;
	wire [4-1:0] node11065;
	wire [4-1:0] node11068;
	wire [4-1:0] node11071;
	wire [4-1:0] node11072;
	wire [4-1:0] node11074;
	wire [4-1:0] node11076;
	wire [4-1:0] node11079;
	wire [4-1:0] node11080;
	wire [4-1:0] node11084;
	wire [4-1:0] node11085;
	wire [4-1:0] node11086;
	wire [4-1:0] node11089;
	wire [4-1:0] node11092;
	wire [4-1:0] node11093;
	wire [4-1:0] node11095;
	wire [4-1:0] node11098;
	wire [4-1:0] node11099;
	wire [4-1:0] node11102;
	wire [4-1:0] node11105;
	wire [4-1:0] node11106;
	wire [4-1:0] node11107;
	wire [4-1:0] node11108;
	wire [4-1:0] node11109;
	wire [4-1:0] node11112;
	wire [4-1:0] node11116;
	wire [4-1:0] node11117;
	wire [4-1:0] node11118;
	wire [4-1:0] node11122;
	wire [4-1:0] node11123;
	wire [4-1:0] node11126;
	wire [4-1:0] node11129;
	wire [4-1:0] node11130;
	wire [4-1:0] node11133;
	wire [4-1:0] node11136;
	wire [4-1:0] node11137;
	wire [4-1:0] node11138;
	wire [4-1:0] node11139;
	wire [4-1:0] node11140;
	wire [4-1:0] node11141;
	wire [4-1:0] node11142;
	wire [4-1:0] node11143;
	wire [4-1:0] node11146;
	wire [4-1:0] node11147;
	wire [4-1:0] node11152;
	wire [4-1:0] node11153;
	wire [4-1:0] node11155;
	wire [4-1:0] node11158;
	wire [4-1:0] node11159;
	wire [4-1:0] node11163;
	wire [4-1:0] node11164;
	wire [4-1:0] node11165;
	wire [4-1:0] node11166;
	wire [4-1:0] node11170;
	wire [4-1:0] node11171;
	wire [4-1:0] node11175;
	wire [4-1:0] node11176;
	wire [4-1:0] node11178;
	wire [4-1:0] node11179;
	wire [4-1:0] node11183;
	wire [4-1:0] node11184;
	wire [4-1:0] node11185;
	wire [4-1:0] node11189;
	wire [4-1:0] node11190;
	wire [4-1:0] node11193;
	wire [4-1:0] node11196;
	wire [4-1:0] node11197;
	wire [4-1:0] node11198;
	wire [4-1:0] node11199;
	wire [4-1:0] node11200;
	wire [4-1:0] node11204;
	wire [4-1:0] node11205;
	wire [4-1:0] node11207;
	wire [4-1:0] node11210;
	wire [4-1:0] node11211;
	wire [4-1:0] node11215;
	wire [4-1:0] node11216;
	wire [4-1:0] node11217;
	wire [4-1:0] node11220;
	wire [4-1:0] node11222;
	wire [4-1:0] node11225;
	wire [4-1:0] node11226;
	wire [4-1:0] node11229;
	wire [4-1:0] node11232;
	wire [4-1:0] node11233;
	wire [4-1:0] node11234;
	wire [4-1:0] node11236;
	wire [4-1:0] node11237;
	wire [4-1:0] node11241;
	wire [4-1:0] node11242;
	wire [4-1:0] node11244;
	wire [4-1:0] node11247;
	wire [4-1:0] node11250;
	wire [4-1:0] node11251;
	wire [4-1:0] node11253;
	wire [4-1:0] node11254;
	wire [4-1:0] node11258;
	wire [4-1:0] node11259;
	wire [4-1:0] node11261;
	wire [4-1:0] node11264;
	wire [4-1:0] node11265;
	wire [4-1:0] node11268;
	wire [4-1:0] node11271;
	wire [4-1:0] node11272;
	wire [4-1:0] node11273;
	wire [4-1:0] node11274;
	wire [4-1:0] node11275;
	wire [4-1:0] node11277;
	wire [4-1:0] node11279;
	wire [4-1:0] node11282;
	wire [4-1:0] node11283;
	wire [4-1:0] node11284;
	wire [4-1:0] node11287;
	wire [4-1:0] node11290;
	wire [4-1:0] node11292;
	wire [4-1:0] node11295;
	wire [4-1:0] node11296;
	wire [4-1:0] node11297;
	wire [4-1:0] node11298;
	wire [4-1:0] node11301;
	wire [4-1:0] node11304;
	wire [4-1:0] node11305;
	wire [4-1:0] node11308;
	wire [4-1:0] node11311;
	wire [4-1:0] node11312;
	wire [4-1:0] node11315;
	wire [4-1:0] node11318;
	wire [4-1:0] node11319;
	wire [4-1:0] node11320;
	wire [4-1:0] node11321;
	wire [4-1:0] node11323;
	wire [4-1:0] node11326;
	wire [4-1:0] node11328;
	wire [4-1:0] node11331;
	wire [4-1:0] node11332;
	wire [4-1:0] node11333;
	wire [4-1:0] node11338;
	wire [4-1:0] node11339;
	wire [4-1:0] node11340;
	wire [4-1:0] node11341;
	wire [4-1:0] node11345;
	wire [4-1:0] node11346;
	wire [4-1:0] node11349;
	wire [4-1:0] node11352;
	wire [4-1:0] node11354;
	wire [4-1:0] node11357;
	wire [4-1:0] node11358;
	wire [4-1:0] node11359;
	wire [4-1:0] node11360;
	wire [4-1:0] node11361;
	wire [4-1:0] node11362;
	wire [4-1:0] node11366;
	wire [4-1:0] node11368;
	wire [4-1:0] node11371;
	wire [4-1:0] node11373;
	wire [4-1:0] node11374;
	wire [4-1:0] node11378;
	wire [4-1:0] node11379;
	wire [4-1:0] node11381;
	wire [4-1:0] node11382;
	wire [4-1:0] node11385;
	wire [4-1:0] node11388;
	wire [4-1:0] node11389;
	wire [4-1:0] node11390;
	wire [4-1:0] node11393;
	wire [4-1:0] node11397;
	wire [4-1:0] node11398;
	wire [4-1:0] node11399;
	wire [4-1:0] node11400;
	wire [4-1:0] node11404;
	wire [4-1:0] node11405;
	wire [4-1:0] node11408;
	wire [4-1:0] node11411;
	wire [4-1:0] node11412;
	wire [4-1:0] node11413;
	wire [4-1:0] node11414;
	wire [4-1:0] node11418;
	wire [4-1:0] node11419;
	wire [4-1:0] node11423;
	wire [4-1:0] node11425;
	wire [4-1:0] node11426;
	wire [4-1:0] node11429;
	wire [4-1:0] node11432;
	wire [4-1:0] node11433;
	wire [4-1:0] node11434;
	wire [4-1:0] node11435;
	wire [4-1:0] node11436;
	wire [4-1:0] node11437;
	wire [4-1:0] node11438;
	wire [4-1:0] node11442;
	wire [4-1:0] node11443;
	wire [4-1:0] node11446;
	wire [4-1:0] node11449;
	wire [4-1:0] node11450;
	wire [4-1:0] node11451;
	wire [4-1:0] node11452;
	wire [4-1:0] node11456;
	wire [4-1:0] node11459;
	wire [4-1:0] node11461;
	wire [4-1:0] node11463;
	wire [4-1:0] node11466;
	wire [4-1:0] node11467;
	wire [4-1:0] node11468;
	wire [4-1:0] node11470;
	wire [4-1:0] node11473;
	wire [4-1:0] node11474;
	wire [4-1:0] node11477;
	wire [4-1:0] node11480;
	wire [4-1:0] node11481;
	wire [4-1:0] node11482;
	wire [4-1:0] node11484;
	wire [4-1:0] node11487;
	wire [4-1:0] node11488;
	wire [4-1:0] node11492;
	wire [4-1:0] node11493;
	wire [4-1:0] node11496;
	wire [4-1:0] node11499;
	wire [4-1:0] node11500;
	wire [4-1:0] node11501;
	wire [4-1:0] node11502;
	wire [4-1:0] node11504;
	wire [4-1:0] node11507;
	wire [4-1:0] node11508;
	wire [4-1:0] node11509;
	wire [4-1:0] node11512;
	wire [4-1:0] node11515;
	wire [4-1:0] node11516;
	wire [4-1:0] node11519;
	wire [4-1:0] node11522;
	wire [4-1:0] node11523;
	wire [4-1:0] node11524;
	wire [4-1:0] node11527;
	wire [4-1:0] node11530;
	wire [4-1:0] node11531;
	wire [4-1:0] node11534;
	wire [4-1:0] node11535;
	wire [4-1:0] node11539;
	wire [4-1:0] node11540;
	wire [4-1:0] node11541;
	wire [4-1:0] node11542;
	wire [4-1:0] node11543;
	wire [4-1:0] node11546;
	wire [4-1:0] node11550;
	wire [4-1:0] node11552;
	wire [4-1:0] node11555;
	wire [4-1:0] node11556;
	wire [4-1:0] node11559;
	wire [4-1:0] node11562;
	wire [4-1:0] node11563;
	wire [4-1:0] node11564;
	wire [4-1:0] node11565;
	wire [4-1:0] node11566;
	wire [4-1:0] node11567;
	wire [4-1:0] node11569;
	wire [4-1:0] node11572;
	wire [4-1:0] node11573;
	wire [4-1:0] node11576;
	wire [4-1:0] node11579;
	wire [4-1:0] node11580;
	wire [4-1:0] node11581;
	wire [4-1:0] node11584;
	wire [4-1:0] node11588;
	wire [4-1:0] node11589;
	wire [4-1:0] node11590;
	wire [4-1:0] node11591;
	wire [4-1:0] node11594;
	wire [4-1:0] node11598;
	wire [4-1:0] node11600;
	wire [4-1:0] node11603;
	wire [4-1:0] node11604;
	wire [4-1:0] node11605;
	wire [4-1:0] node11606;
	wire [4-1:0] node11610;
	wire [4-1:0] node11611;
	wire [4-1:0] node11612;
	wire [4-1:0] node11615;
	wire [4-1:0] node11619;
	wire [4-1:0] node11620;
	wire [4-1:0] node11621;
	wire [4-1:0] node11624;
	wire [4-1:0] node11627;
	wire [4-1:0] node11628;
	wire [4-1:0] node11631;
	wire [4-1:0] node11634;
	wire [4-1:0] node11635;
	wire [4-1:0] node11636;
	wire [4-1:0] node11637;
	wire [4-1:0] node11639;
	wire [4-1:0] node11640;
	wire [4-1:0] node11644;
	wire [4-1:0] node11645;
	wire [4-1:0] node11648;
	wire [4-1:0] node11651;
	wire [4-1:0] node11652;
	wire [4-1:0] node11653;
	wire [4-1:0] node11656;
	wire [4-1:0] node11659;
	wire [4-1:0] node11660;
	wire [4-1:0] node11663;
	wire [4-1:0] node11666;
	wire [4-1:0] node11667;
	wire [4-1:0] node11668;
	wire [4-1:0] node11669;
	wire [4-1:0] node11672;
	wire [4-1:0] node11675;
	wire [4-1:0] node11676;
	wire [4-1:0] node11679;
	wire [4-1:0] node11682;
	wire [4-1:0] node11683;
	wire [4-1:0] node11684;
	wire [4-1:0] node11685;
	wire [4-1:0] node11689;
	wire [4-1:0] node11690;
	wire [4-1:0] node11694;
	wire [4-1:0] node11695;
	wire [4-1:0] node11696;
	wire [4-1:0] node11700;
	wire [4-1:0] node11702;
	wire [4-1:0] node11705;
	wire [4-1:0] node11706;
	wire [4-1:0] node11707;
	wire [4-1:0] node11708;
	wire [4-1:0] node11709;
	wire [4-1:0] node11710;
	wire [4-1:0] node11711;
	wire [4-1:0] node11712;
	wire [4-1:0] node11713;
	wire [4-1:0] node11716;
	wire [4-1:0] node11719;
	wire [4-1:0] node11720;
	wire [4-1:0] node11723;
	wire [4-1:0] node11726;
	wire [4-1:0] node11727;
	wire [4-1:0] node11728;
	wire [4-1:0] node11732;
	wire [4-1:0] node11733;
	wire [4-1:0] node11737;
	wire [4-1:0] node11738;
	wire [4-1:0] node11739;
	wire [4-1:0] node11740;
	wire [4-1:0] node11741;
	wire [4-1:0] node11745;
	wire [4-1:0] node11746;
	wire [4-1:0] node11750;
	wire [4-1:0] node11751;
	wire [4-1:0] node11755;
	wire [4-1:0] node11756;
	wire [4-1:0] node11759;
	wire [4-1:0] node11762;
	wire [4-1:0] node11763;
	wire [4-1:0] node11764;
	wire [4-1:0] node11766;
	wire [4-1:0] node11767;
	wire [4-1:0] node11768;
	wire [4-1:0] node11772;
	wire [4-1:0] node11773;
	wire [4-1:0] node11776;
	wire [4-1:0] node11779;
	wire [4-1:0] node11780;
	wire [4-1:0] node11782;
	wire [4-1:0] node11785;
	wire [4-1:0] node11788;
	wire [4-1:0] node11789;
	wire [4-1:0] node11790;
	wire [4-1:0] node11791;
	wire [4-1:0] node11794;
	wire [4-1:0] node11797;
	wire [4-1:0] node11798;
	wire [4-1:0] node11801;
	wire [4-1:0] node11804;
	wire [4-1:0] node11805;
	wire [4-1:0] node11807;
	wire [4-1:0] node11808;
	wire [4-1:0] node11811;
	wire [4-1:0] node11814;
	wire [4-1:0] node11815;
	wire [4-1:0] node11816;
	wire [4-1:0] node11820;
	wire [4-1:0] node11823;
	wire [4-1:0] node11824;
	wire [4-1:0] node11825;
	wire [4-1:0] node11826;
	wire [4-1:0] node11827;
	wire [4-1:0] node11828;
	wire [4-1:0] node11831;
	wire [4-1:0] node11833;
	wire [4-1:0] node11836;
	wire [4-1:0] node11837;
	wire [4-1:0] node11839;
	wire [4-1:0] node11842;
	wire [4-1:0] node11843;
	wire [4-1:0] node11847;
	wire [4-1:0] node11848;
	wire [4-1:0] node11849;
	wire [4-1:0] node11852;
	wire [4-1:0] node11853;
	wire [4-1:0] node11857;
	wire [4-1:0] node11858;
	wire [4-1:0] node11861;
	wire [4-1:0] node11864;
	wire [4-1:0] node11865;
	wire [4-1:0] node11866;
	wire [4-1:0] node11869;
	wire [4-1:0] node11870;
	wire [4-1:0] node11872;
	wire [4-1:0] node11876;
	wire [4-1:0] node11877;
	wire [4-1:0] node11878;
	wire [4-1:0] node11879;
	wire [4-1:0] node11883;
	wire [4-1:0] node11884;
	wire [4-1:0] node11887;
	wire [4-1:0] node11890;
	wire [4-1:0] node11891;
	wire [4-1:0] node11894;
	wire [4-1:0] node11896;
	wire [4-1:0] node11899;
	wire [4-1:0] node11900;
	wire [4-1:0] node11901;
	wire [4-1:0] node11902;
	wire [4-1:0] node11904;
	wire [4-1:0] node11906;
	wire [4-1:0] node11909;
	wire [4-1:0] node11910;
	wire [4-1:0] node11911;
	wire [4-1:0] node11914;
	wire [4-1:0] node11917;
	wire [4-1:0] node11919;
	wire [4-1:0] node11922;
	wire [4-1:0] node11923;
	wire [4-1:0] node11924;
	wire [4-1:0] node11926;
	wire [4-1:0] node11930;
	wire [4-1:0] node11931;
	wire [4-1:0] node11932;
	wire [4-1:0] node11937;
	wire [4-1:0] node11938;
	wire [4-1:0] node11939;
	wire [4-1:0] node11940;
	wire [4-1:0] node11941;
	wire [4-1:0] node11945;
	wire [4-1:0] node11946;
	wire [4-1:0] node11950;
	wire [4-1:0] node11951;
	wire [4-1:0] node11954;
	wire [4-1:0] node11956;
	wire [4-1:0] node11959;
	wire [4-1:0] node11960;
	wire [4-1:0] node11962;
	wire [4-1:0] node11965;
	wire [4-1:0] node11966;
	wire [4-1:0] node11969;
	wire [4-1:0] node11972;
	wire [4-1:0] node11973;
	wire [4-1:0] node11974;
	wire [4-1:0] node11975;
	wire [4-1:0] node11976;
	wire [4-1:0] node11977;
	wire [4-1:0] node11978;
	wire [4-1:0] node11982;
	wire [4-1:0] node11983;
	wire [4-1:0] node11986;
	wire [4-1:0] node11987;
	wire [4-1:0] node11991;
	wire [4-1:0] node11992;
	wire [4-1:0] node11993;
	wire [4-1:0] node11996;
	wire [4-1:0] node11999;
	wire [4-1:0] node12001;
	wire [4-1:0] node12004;
	wire [4-1:0] node12005;
	wire [4-1:0] node12006;
	wire [4-1:0] node12009;
	wire [4-1:0] node12011;
	wire [4-1:0] node12014;
	wire [4-1:0] node12015;
	wire [4-1:0] node12016;
	wire [4-1:0] node12020;
	wire [4-1:0] node12021;
	wire [4-1:0] node12024;
	wire [4-1:0] node12027;
	wire [4-1:0] node12028;
	wire [4-1:0] node12029;
	wire [4-1:0] node12030;
	wire [4-1:0] node12031;
	wire [4-1:0] node12035;
	wire [4-1:0] node12037;
	wire [4-1:0] node12040;
	wire [4-1:0] node12041;
	wire [4-1:0] node12042;
	wire [4-1:0] node12045;
	wire [4-1:0] node12048;
	wire [4-1:0] node12049;
	wire [4-1:0] node12052;
	wire [4-1:0] node12055;
	wire [4-1:0] node12056;
	wire [4-1:0] node12057;
	wire [4-1:0] node12059;
	wire [4-1:0] node12062;
	wire [4-1:0] node12064;
	wire [4-1:0] node12067;
	wire [4-1:0] node12068;
	wire [4-1:0] node12069;
	wire [4-1:0] node12072;
	wire [4-1:0] node12075;
	wire [4-1:0] node12076;
	wire [4-1:0] node12078;
	wire [4-1:0] node12081;
	wire [4-1:0] node12084;
	wire [4-1:0] node12085;
	wire [4-1:0] node12086;
	wire [4-1:0] node12087;
	wire [4-1:0] node12088;
	wire [4-1:0] node12089;
	wire [4-1:0] node12090;
	wire [4-1:0] node12094;
	wire [4-1:0] node12096;
	wire [4-1:0] node12099;
	wire [4-1:0] node12100;
	wire [4-1:0] node12103;
	wire [4-1:0] node12106;
	wire [4-1:0] node12107;
	wire [4-1:0] node12108;
	wire [4-1:0] node12112;
	wire [4-1:0] node12113;
	wire [4-1:0] node12116;
	wire [4-1:0] node12119;
	wire [4-1:0] node12120;
	wire [4-1:0] node12121;
	wire [4-1:0] node12124;
	wire [4-1:0] node12126;
	wire [4-1:0] node12129;
	wire [4-1:0] node12130;
	wire [4-1:0] node12131;
	wire [4-1:0] node12134;
	wire [4-1:0] node12137;
	wire [4-1:0] node12138;
	wire [4-1:0] node12141;
	wire [4-1:0] node12144;
	wire [4-1:0] node12145;
	wire [4-1:0] node12146;
	wire [4-1:0] node12147;
	wire [4-1:0] node12148;
	wire [4-1:0] node12151;
	wire [4-1:0] node12154;
	wire [4-1:0] node12156;
	wire [4-1:0] node12158;
	wire [4-1:0] node12161;
	wire [4-1:0] node12162;
	wire [4-1:0] node12165;
	wire [4-1:0] node12168;
	wire [4-1:0] node12169;
	wire [4-1:0] node12170;
	wire [4-1:0] node12171;
	wire [4-1:0] node12174;
	wire [4-1:0] node12177;
	wire [4-1:0] node12178;
	wire [4-1:0] node12181;
	wire [4-1:0] node12184;
	wire [4-1:0] node12185;
	wire [4-1:0] node12186;
	wire [4-1:0] node12189;
	wire [4-1:0] node12193;
	wire [4-1:0] node12194;
	wire [4-1:0] node12195;
	wire [4-1:0] node12196;
	wire [4-1:0] node12197;
	wire [4-1:0] node12198;
	wire [4-1:0] node12199;
	wire [4-1:0] node12200;
	wire [4-1:0] node12203;
	wire [4-1:0] node12206;
	wire [4-1:0] node12209;
	wire [4-1:0] node12210;
	wire [4-1:0] node12211;
	wire [4-1:0] node12212;
	wire [4-1:0] node12215;
	wire [4-1:0] node12218;
	wire [4-1:0] node12219;
	wire [4-1:0] node12222;
	wire [4-1:0] node12225;
	wire [4-1:0] node12226;
	wire [4-1:0] node12228;
	wire [4-1:0] node12231;
	wire [4-1:0] node12232;
	wire [4-1:0] node12235;
	wire [4-1:0] node12238;
	wire [4-1:0] node12239;
	wire [4-1:0] node12240;
	wire [4-1:0] node12241;
	wire [4-1:0] node12244;
	wire [4-1:0] node12247;
	wire [4-1:0] node12248;
	wire [4-1:0] node12249;
	wire [4-1:0] node12254;
	wire [4-1:0] node12255;
	wire [4-1:0] node12256;
	wire [4-1:0] node12259;
	wire [4-1:0] node12261;
	wire [4-1:0] node12264;
	wire [4-1:0] node12265;
	wire [4-1:0] node12266;
	wire [4-1:0] node12271;
	wire [4-1:0] node12272;
	wire [4-1:0] node12273;
	wire [4-1:0] node12274;
	wire [4-1:0] node12276;
	wire [4-1:0] node12277;
	wire [4-1:0] node12280;
	wire [4-1:0] node12283;
	wire [4-1:0] node12284;
	wire [4-1:0] node12285;
	wire [4-1:0] node12289;
	wire [4-1:0] node12290;
	wire [4-1:0] node12294;
	wire [4-1:0] node12295;
	wire [4-1:0] node12296;
	wire [4-1:0] node12297;
	wire [4-1:0] node12302;
	wire [4-1:0] node12304;
	wire [4-1:0] node12307;
	wire [4-1:0] node12308;
	wire [4-1:0] node12309;
	wire [4-1:0] node12310;
	wire [4-1:0] node12311;
	wire [4-1:0] node12314;
	wire [4-1:0] node12318;
	wire [4-1:0] node12320;
	wire [4-1:0] node12323;
	wire [4-1:0] node12324;
	wire [4-1:0] node12326;
	wire [4-1:0] node12329;
	wire [4-1:0] node12330;
	wire [4-1:0] node12333;
	wire [4-1:0] node12336;
	wire [4-1:0] node12337;
	wire [4-1:0] node12338;
	wire [4-1:0] node12339;
	wire [4-1:0] node12340;
	wire [4-1:0] node12342;
	wire [4-1:0] node12343;
	wire [4-1:0] node12346;
	wire [4-1:0] node12349;
	wire [4-1:0] node12350;
	wire [4-1:0] node12353;
	wire [4-1:0] node12356;
	wire [4-1:0] node12357;
	wire [4-1:0] node12358;
	wire [4-1:0] node12359;
	wire [4-1:0] node12363;
	wire [4-1:0] node12365;
	wire [4-1:0] node12368;
	wire [4-1:0] node12370;
	wire [4-1:0] node12372;
	wire [4-1:0] node12375;
	wire [4-1:0] node12376;
	wire [4-1:0] node12377;
	wire [4-1:0] node12378;
	wire [4-1:0] node12381;
	wire [4-1:0] node12385;
	wire [4-1:0] node12386;
	wire [4-1:0] node12388;
	wire [4-1:0] node12391;
	wire [4-1:0] node12392;
	wire [4-1:0] node12394;
	wire [4-1:0] node12398;
	wire [4-1:0] node12399;
	wire [4-1:0] node12400;
	wire [4-1:0] node12401;
	wire [4-1:0] node12402;
	wire [4-1:0] node12404;
	wire [4-1:0] node12407;
	wire [4-1:0] node12408;
	wire [4-1:0] node12412;
	wire [4-1:0] node12414;
	wire [4-1:0] node12417;
	wire [4-1:0] node12418;
	wire [4-1:0] node12419;
	wire [4-1:0] node12420;
	wire [4-1:0] node12424;
	wire [4-1:0] node12425;
	wire [4-1:0] node12428;
	wire [4-1:0] node12431;
	wire [4-1:0] node12432;
	wire [4-1:0] node12434;
	wire [4-1:0] node12437;
	wire [4-1:0] node12439;
	wire [4-1:0] node12442;
	wire [4-1:0] node12443;
	wire [4-1:0] node12445;
	wire [4-1:0] node12448;
	wire [4-1:0] node12449;
	wire [4-1:0] node12450;
	wire [4-1:0] node12451;
	wire [4-1:0] node12456;
	wire [4-1:0] node12457;
	wire [4-1:0] node12458;
	wire [4-1:0] node12461;
	wire [4-1:0] node12465;
	wire [4-1:0] node12466;
	wire [4-1:0] node12467;
	wire [4-1:0] node12468;
	wire [4-1:0] node12469;
	wire [4-1:0] node12470;
	wire [4-1:0] node12471;
	wire [4-1:0] node12474;
	wire [4-1:0] node12478;
	wire [4-1:0] node12479;
	wire [4-1:0] node12480;
	wire [4-1:0] node12484;
	wire [4-1:0] node12487;
	wire [4-1:0] node12488;
	wire [4-1:0] node12489;
	wire [4-1:0] node12490;
	wire [4-1:0] node12492;
	wire [4-1:0] node12495;
	wire [4-1:0] node12496;
	wire [4-1:0] node12499;
	wire [4-1:0] node12502;
	wire [4-1:0] node12503;
	wire [4-1:0] node12506;
	wire [4-1:0] node12508;
	wire [4-1:0] node12511;
	wire [4-1:0] node12512;
	wire [4-1:0] node12513;
	wire [4-1:0] node12516;
	wire [4-1:0] node12519;
	wire [4-1:0] node12520;
	wire [4-1:0] node12522;
	wire [4-1:0] node12526;
	wire [4-1:0] node12527;
	wire [4-1:0] node12528;
	wire [4-1:0] node12529;
	wire [4-1:0] node12531;
	wire [4-1:0] node12534;
	wire [4-1:0] node12536;
	wire [4-1:0] node12539;
	wire [4-1:0] node12541;
	wire [4-1:0] node12542;
	wire [4-1:0] node12545;
	wire [4-1:0] node12548;
	wire [4-1:0] node12549;
	wire [4-1:0] node12550;
	wire [4-1:0] node12552;
	wire [4-1:0] node12553;
	wire [4-1:0] node12556;
	wire [4-1:0] node12559;
	wire [4-1:0] node12560;
	wire [4-1:0] node12562;
	wire [4-1:0] node12566;
	wire [4-1:0] node12567;
	wire [4-1:0] node12569;
	wire [4-1:0] node12570;
	wire [4-1:0] node12573;
	wire [4-1:0] node12576;
	wire [4-1:0] node12578;
	wire [4-1:0] node12580;
	wire [4-1:0] node12583;
	wire [4-1:0] node12584;
	wire [4-1:0] node12585;
	wire [4-1:0] node12586;
	wire [4-1:0] node12587;
	wire [4-1:0] node12588;
	wire [4-1:0] node12591;
	wire [4-1:0] node12594;
	wire [4-1:0] node12597;
	wire [4-1:0] node12598;
	wire [4-1:0] node12599;
	wire [4-1:0] node12600;
	wire [4-1:0] node12603;
	wire [4-1:0] node12606;
	wire [4-1:0] node12608;
	wire [4-1:0] node12611;
	wire [4-1:0] node12612;
	wire [4-1:0] node12613;
	wire [4-1:0] node12616;
	wire [4-1:0] node12620;
	wire [4-1:0] node12621;
	wire [4-1:0] node12622;
	wire [4-1:0] node12623;
	wire [4-1:0] node12626;
	wire [4-1:0] node12629;
	wire [4-1:0] node12630;
	wire [4-1:0] node12632;
	wire [4-1:0] node12635;
	wire [4-1:0] node12637;
	wire [4-1:0] node12640;
	wire [4-1:0] node12641;
	wire [4-1:0] node12643;
	wire [4-1:0] node12644;
	wire [4-1:0] node12647;
	wire [4-1:0] node12650;
	wire [4-1:0] node12651;
	wire [4-1:0] node12653;
	wire [4-1:0] node12656;
	wire [4-1:0] node12658;
	wire [4-1:0] node12661;
	wire [4-1:0] node12662;
	wire [4-1:0] node12663;
	wire [4-1:0] node12665;
	wire [4-1:0] node12668;
	wire [4-1:0] node12669;
	wire [4-1:0] node12671;
	wire [4-1:0] node12675;
	wire [4-1:0] node12676;
	wire [4-1:0] node12677;
	wire [4-1:0] node12678;
	wire [4-1:0] node12679;
	wire [4-1:0] node12683;
	wire [4-1:0] node12684;
	wire [4-1:0] node12688;
	wire [4-1:0] node12689;
	wire [4-1:0] node12692;
	wire [4-1:0] node12695;
	wire [4-1:0] node12696;
	wire [4-1:0] node12697;
	wire [4-1:0] node12700;
	wire [4-1:0] node12703;
	wire [4-1:0] node12704;
	wire [4-1:0] node12707;
	wire [4-1:0] node12710;
	wire [4-1:0] node12711;
	wire [4-1:0] node12712;
	wire [4-1:0] node12713;
	wire [4-1:0] node12714;
	wire [4-1:0] node12715;
	wire [4-1:0] node12716;
	wire [4-1:0] node12717;
	wire [4-1:0] node12718;
	wire [4-1:0] node12720;
	wire [4-1:0] node12721;
	wire [4-1:0] node12724;
	wire [4-1:0] node12727;
	wire [4-1:0] node12728;
	wire [4-1:0] node12731;
	wire [4-1:0] node12734;
	wire [4-1:0] node12735;
	wire [4-1:0] node12736;
	wire [4-1:0] node12737;
	wire [4-1:0] node12740;
	wire [4-1:0] node12743;
	wire [4-1:0] node12745;
	wire [4-1:0] node12748;
	wire [4-1:0] node12751;
	wire [4-1:0] node12752;
	wire [4-1:0] node12753;
	wire [4-1:0] node12755;
	wire [4-1:0] node12756;
	wire [4-1:0] node12760;
	wire [4-1:0] node12761;
	wire [4-1:0] node12762;
	wire [4-1:0] node12765;
	wire [4-1:0] node12768;
	wire [4-1:0] node12770;
	wire [4-1:0] node12773;
	wire [4-1:0] node12774;
	wire [4-1:0] node12775;
	wire [4-1:0] node12777;
	wire [4-1:0] node12780;
	wire [4-1:0] node12781;
	wire [4-1:0] node12785;
	wire [4-1:0] node12786;
	wire [4-1:0] node12787;
	wire [4-1:0] node12790;
	wire [4-1:0] node12793;
	wire [4-1:0] node12794;
	wire [4-1:0] node12797;
	wire [4-1:0] node12800;
	wire [4-1:0] node12801;
	wire [4-1:0] node12802;
	wire [4-1:0] node12803;
	wire [4-1:0] node12806;
	wire [4-1:0] node12807;
	wire [4-1:0] node12810;
	wire [4-1:0] node12811;
	wire [4-1:0] node12814;
	wire [4-1:0] node12817;
	wire [4-1:0] node12818;
	wire [4-1:0] node12820;
	wire [4-1:0] node12822;
	wire [4-1:0] node12825;
	wire [4-1:0] node12826;
	wire [4-1:0] node12828;
	wire [4-1:0] node12832;
	wire [4-1:0] node12833;
	wire [4-1:0] node12834;
	wire [4-1:0] node12835;
	wire [4-1:0] node12838;
	wire [4-1:0] node12839;
	wire [4-1:0] node12842;
	wire [4-1:0] node12845;
	wire [4-1:0] node12846;
	wire [4-1:0] node12847;
	wire [4-1:0] node12850;
	wire [4-1:0] node12853;
	wire [4-1:0] node12854;
	wire [4-1:0] node12857;
	wire [4-1:0] node12860;
	wire [4-1:0] node12861;
	wire [4-1:0] node12862;
	wire [4-1:0] node12863;
	wire [4-1:0] node12868;
	wire [4-1:0] node12870;
	wire [4-1:0] node12871;
	wire [4-1:0] node12875;
	wire [4-1:0] node12876;
	wire [4-1:0] node12877;
	wire [4-1:0] node12878;
	wire [4-1:0] node12879;
	wire [4-1:0] node12880;
	wire [4-1:0] node12881;
	wire [4-1:0] node12884;
	wire [4-1:0] node12887;
	wire [4-1:0] node12890;
	wire [4-1:0] node12891;
	wire [4-1:0] node12895;
	wire [4-1:0] node12896;
	wire [4-1:0] node12897;
	wire [4-1:0] node12900;
	wire [4-1:0] node12903;
	wire [4-1:0] node12904;
	wire [4-1:0] node12905;
	wire [4-1:0] node12909;
	wire [4-1:0] node12910;
	wire [4-1:0] node12913;
	wire [4-1:0] node12916;
	wire [4-1:0] node12917;
	wire [4-1:0] node12918;
	wire [4-1:0] node12920;
	wire [4-1:0] node12923;
	wire [4-1:0] node12924;
	wire [4-1:0] node12928;
	wire [4-1:0] node12929;
	wire [4-1:0] node12930;
	wire [4-1:0] node12933;
	wire [4-1:0] node12934;
	wire [4-1:0] node12938;
	wire [4-1:0] node12941;
	wire [4-1:0] node12942;
	wire [4-1:0] node12943;
	wire [4-1:0] node12944;
	wire [4-1:0] node12945;
	wire [4-1:0] node12949;
	wire [4-1:0] node12950;
	wire [4-1:0] node12952;
	wire [4-1:0] node12955;
	wire [4-1:0] node12956;
	wire [4-1:0] node12960;
	wire [4-1:0] node12961;
	wire [4-1:0] node12962;
	wire [4-1:0] node12964;
	wire [4-1:0] node12968;
	wire [4-1:0] node12969;
	wire [4-1:0] node12971;
	wire [4-1:0] node12974;
	wire [4-1:0] node12975;
	wire [4-1:0] node12979;
	wire [4-1:0] node12980;
	wire [4-1:0] node12981;
	wire [4-1:0] node12982;
	wire [4-1:0] node12983;
	wire [4-1:0] node12986;
	wire [4-1:0] node12990;
	wire [4-1:0] node12991;
	wire [4-1:0] node12993;
	wire [4-1:0] node12996;
	wire [4-1:0] node12997;
	wire [4-1:0] node13001;
	wire [4-1:0] node13002;
	wire [4-1:0] node13003;
	wire [4-1:0] node13004;
	wire [4-1:0] node13008;
	wire [4-1:0] node13011;
	wire [4-1:0] node13012;
	wire [4-1:0] node13014;
	wire [4-1:0] node13017;
	wire [4-1:0] node13019;
	wire [4-1:0] node13022;
	wire [4-1:0] node13023;
	wire [4-1:0] node13024;
	wire [4-1:0] node13025;
	wire [4-1:0] node13026;
	wire [4-1:0] node13027;
	wire [4-1:0] node13029;
	wire [4-1:0] node13030;
	wire [4-1:0] node13033;
	wire [4-1:0] node13036;
	wire [4-1:0] node13038;
	wire [4-1:0] node13041;
	wire [4-1:0] node13042;
	wire [4-1:0] node13043;
	wire [4-1:0] node13045;
	wire [4-1:0] node13048;
	wire [4-1:0] node13049;
	wire [4-1:0] node13053;
	wire [4-1:0] node13054;
	wire [4-1:0] node13055;
	wire [4-1:0] node13058;
	wire [4-1:0] node13061;
	wire [4-1:0] node13062;
	wire [4-1:0] node13065;
	wire [4-1:0] node13068;
	wire [4-1:0] node13069;
	wire [4-1:0] node13070;
	wire [4-1:0] node13071;
	wire [4-1:0] node13072;
	wire [4-1:0] node13075;
	wire [4-1:0] node13078;
	wire [4-1:0] node13081;
	wire [4-1:0] node13082;
	wire [4-1:0] node13084;
	wire [4-1:0] node13088;
	wire [4-1:0] node13089;
	wire [4-1:0] node13090;
	wire [4-1:0] node13093;
	wire [4-1:0] node13094;
	wire [4-1:0] node13097;
	wire [4-1:0] node13100;
	wire [4-1:0] node13102;
	wire [4-1:0] node13104;
	wire [4-1:0] node13107;
	wire [4-1:0] node13108;
	wire [4-1:0] node13109;
	wire [4-1:0] node13110;
	wire [4-1:0] node13111;
	wire [4-1:0] node13112;
	wire [4-1:0] node13115;
	wire [4-1:0] node13118;
	wire [4-1:0] node13120;
	wire [4-1:0] node13123;
	wire [4-1:0] node13124;
	wire [4-1:0] node13125;
	wire [4-1:0] node13129;
	wire [4-1:0] node13131;
	wire [4-1:0] node13134;
	wire [4-1:0] node13135;
	wire [4-1:0] node13136;
	wire [4-1:0] node13139;
	wire [4-1:0] node13141;
	wire [4-1:0] node13144;
	wire [4-1:0] node13145;
	wire [4-1:0] node13148;
	wire [4-1:0] node13149;
	wire [4-1:0] node13152;
	wire [4-1:0] node13155;
	wire [4-1:0] node13156;
	wire [4-1:0] node13157;
	wire [4-1:0] node13158;
	wire [4-1:0] node13161;
	wire [4-1:0] node13162;
	wire [4-1:0] node13165;
	wire [4-1:0] node13168;
	wire [4-1:0] node13169;
	wire [4-1:0] node13172;
	wire [4-1:0] node13173;
	wire [4-1:0] node13176;
	wire [4-1:0] node13179;
	wire [4-1:0] node13180;
	wire [4-1:0] node13181;
	wire [4-1:0] node13183;
	wire [4-1:0] node13186;
	wire [4-1:0] node13187;
	wire [4-1:0] node13191;
	wire [4-1:0] node13193;
	wire [4-1:0] node13195;
	wire [4-1:0] node13198;
	wire [4-1:0] node13199;
	wire [4-1:0] node13200;
	wire [4-1:0] node13201;
	wire [4-1:0] node13202;
	wire [4-1:0] node13203;
	wire [4-1:0] node13204;
	wire [4-1:0] node13207;
	wire [4-1:0] node13211;
	wire [4-1:0] node13212;
	wire [4-1:0] node13215;
	wire [4-1:0] node13218;
	wire [4-1:0] node13220;
	wire [4-1:0] node13221;
	wire [4-1:0] node13224;
	wire [4-1:0] node13225;
	wire [4-1:0] node13228;
	wire [4-1:0] node13231;
	wire [4-1:0] node13232;
	wire [4-1:0] node13233;
	wire [4-1:0] node13234;
	wire [4-1:0] node13235;
	wire [4-1:0] node13239;
	wire [4-1:0] node13240;
	wire [4-1:0] node13243;
	wire [4-1:0] node13246;
	wire [4-1:0] node13248;
	wire [4-1:0] node13251;
	wire [4-1:0] node13252;
	wire [4-1:0] node13253;
	wire [4-1:0] node13256;
	wire [4-1:0] node13259;
	wire [4-1:0] node13261;
	wire [4-1:0] node13264;
	wire [4-1:0] node13265;
	wire [4-1:0] node13266;
	wire [4-1:0] node13267;
	wire [4-1:0] node13268;
	wire [4-1:0] node13269;
	wire [4-1:0] node13272;
	wire [4-1:0] node13275;
	wire [4-1:0] node13278;
	wire [4-1:0] node13279;
	wire [4-1:0] node13283;
	wire [4-1:0] node13284;
	wire [4-1:0] node13285;
	wire [4-1:0] node13286;
	wire [4-1:0] node13289;
	wire [4-1:0] node13292;
	wire [4-1:0] node13293;
	wire [4-1:0] node13297;
	wire [4-1:0] node13298;
	wire [4-1:0] node13302;
	wire [4-1:0] node13303;
	wire [4-1:0] node13304;
	wire [4-1:0] node13305;
	wire [4-1:0] node13307;
	wire [4-1:0] node13310;
	wire [4-1:0] node13311;
	wire [4-1:0] node13314;
	wire [4-1:0] node13317;
	wire [4-1:0] node13319;
	wire [4-1:0] node13320;
	wire [4-1:0] node13323;
	wire [4-1:0] node13326;
	wire [4-1:0] node13327;
	wire [4-1:0] node13328;
	wire [4-1:0] node13329;
	wire [4-1:0] node13332;
	wire [4-1:0] node13336;
	wire [4-1:0] node13337;
	wire [4-1:0] node13340;
	wire [4-1:0] node13343;
	wire [4-1:0] node13344;
	wire [4-1:0] node13345;
	wire [4-1:0] node13346;
	wire [4-1:0] node13347;
	wire [4-1:0] node13348;
	wire [4-1:0] node13349;
	wire [4-1:0] node13350;
	wire [4-1:0] node13352;
	wire [4-1:0] node13355;
	wire [4-1:0] node13358;
	wire [4-1:0] node13361;
	wire [4-1:0] node13362;
	wire [4-1:0] node13363;
	wire [4-1:0] node13366;
	wire [4-1:0] node13367;
	wire [4-1:0] node13370;
	wire [4-1:0] node13373;
	wire [4-1:0] node13374;
	wire [4-1:0] node13375;
	wire [4-1:0] node13380;
	wire [4-1:0] node13381;
	wire [4-1:0] node13382;
	wire [4-1:0] node13383;
	wire [4-1:0] node13384;
	wire [4-1:0] node13387;
	wire [4-1:0] node13391;
	wire [4-1:0] node13393;
	wire [4-1:0] node13394;
	wire [4-1:0] node13397;
	wire [4-1:0] node13400;
	wire [4-1:0] node13401;
	wire [4-1:0] node13402;
	wire [4-1:0] node13403;
	wire [4-1:0] node13407;
	wire [4-1:0] node13408;
	wire [4-1:0] node13412;
	wire [4-1:0] node13413;
	wire [4-1:0] node13414;
	wire [4-1:0] node13418;
	wire [4-1:0] node13421;
	wire [4-1:0] node13422;
	wire [4-1:0] node13423;
	wire [4-1:0] node13424;
	wire [4-1:0] node13425;
	wire [4-1:0] node13426;
	wire [4-1:0] node13432;
	wire [4-1:0] node13433;
	wire [4-1:0] node13435;
	wire [4-1:0] node13437;
	wire [4-1:0] node13440;
	wire [4-1:0] node13442;
	wire [4-1:0] node13443;
	wire [4-1:0] node13446;
	wire [4-1:0] node13449;
	wire [4-1:0] node13450;
	wire [4-1:0] node13451;
	wire [4-1:0] node13452;
	wire [4-1:0] node13453;
	wire [4-1:0] node13457;
	wire [4-1:0] node13460;
	wire [4-1:0] node13461;
	wire [4-1:0] node13463;
	wire [4-1:0] node13466;
	wire [4-1:0] node13467;
	wire [4-1:0] node13470;
	wire [4-1:0] node13473;
	wire [4-1:0] node13474;
	wire [4-1:0] node13475;
	wire [4-1:0] node13478;
	wire [4-1:0] node13479;
	wire [4-1:0] node13482;
	wire [4-1:0] node13485;
	wire [4-1:0] node13488;
	wire [4-1:0] node13489;
	wire [4-1:0] node13490;
	wire [4-1:0] node13491;
	wire [4-1:0] node13492;
	wire [4-1:0] node13493;
	wire [4-1:0] node13494;
	wire [4-1:0] node13499;
	wire [4-1:0] node13500;
	wire [4-1:0] node13501;
	wire [4-1:0] node13504;
	wire [4-1:0] node13507;
	wire [4-1:0] node13509;
	wire [4-1:0] node13512;
	wire [4-1:0] node13513;
	wire [4-1:0] node13514;
	wire [4-1:0] node13515;
	wire [4-1:0] node13520;
	wire [4-1:0] node13521;
	wire [4-1:0] node13524;
	wire [4-1:0] node13525;
	wire [4-1:0] node13529;
	wire [4-1:0] node13530;
	wire [4-1:0] node13531;
	wire [4-1:0] node13532;
	wire [4-1:0] node13534;
	wire [4-1:0] node13538;
	wire [4-1:0] node13539;
	wire [4-1:0] node13540;
	wire [4-1:0] node13543;
	wire [4-1:0] node13546;
	wire [4-1:0] node13548;
	wire [4-1:0] node13551;
	wire [4-1:0] node13552;
	wire [4-1:0] node13554;
	wire [4-1:0] node13555;
	wire [4-1:0] node13558;
	wire [4-1:0] node13561;
	wire [4-1:0] node13562;
	wire [4-1:0] node13563;
	wire [4-1:0] node13567;
	wire [4-1:0] node13569;
	wire [4-1:0] node13572;
	wire [4-1:0] node13573;
	wire [4-1:0] node13574;
	wire [4-1:0] node13575;
	wire [4-1:0] node13577;
	wire [4-1:0] node13578;
	wire [4-1:0] node13581;
	wire [4-1:0] node13584;
	wire [4-1:0] node13585;
	wire [4-1:0] node13586;
	wire [4-1:0] node13589;
	wire [4-1:0] node13592;
	wire [4-1:0] node13593;
	wire [4-1:0] node13596;
	wire [4-1:0] node13599;
	wire [4-1:0] node13600;
	wire [4-1:0] node13601;
	wire [4-1:0] node13604;
	wire [4-1:0] node13605;
	wire [4-1:0] node13608;
	wire [4-1:0] node13611;
	wire [4-1:0] node13612;
	wire [4-1:0] node13614;
	wire [4-1:0] node13617;
	wire [4-1:0] node13618;
	wire [4-1:0] node13621;
	wire [4-1:0] node13624;
	wire [4-1:0] node13625;
	wire [4-1:0] node13626;
	wire [4-1:0] node13627;
	wire [4-1:0] node13628;
	wire [4-1:0] node13632;
	wire [4-1:0] node13633;
	wire [4-1:0] node13637;
	wire [4-1:0] node13640;
	wire [4-1:0] node13641;
	wire [4-1:0] node13642;
	wire [4-1:0] node13644;
	wire [4-1:0] node13647;
	wire [4-1:0] node13648;
	wire [4-1:0] node13651;
	wire [4-1:0] node13654;
	wire [4-1:0] node13656;
	wire [4-1:0] node13659;
	wire [4-1:0] node13660;
	wire [4-1:0] node13661;
	wire [4-1:0] node13662;
	wire [4-1:0] node13663;
	wire [4-1:0] node13664;
	wire [4-1:0] node13665;
	wire [4-1:0] node13666;
	wire [4-1:0] node13669;
	wire [4-1:0] node13672;
	wire [4-1:0] node13673;
	wire [4-1:0] node13677;
	wire [4-1:0] node13679;
	wire [4-1:0] node13681;
	wire [4-1:0] node13684;
	wire [4-1:0] node13685;
	wire [4-1:0] node13687;
	wire [4-1:0] node13690;
	wire [4-1:0] node13691;
	wire [4-1:0] node13694;
	wire [4-1:0] node13697;
	wire [4-1:0] node13698;
	wire [4-1:0] node13699;
	wire [4-1:0] node13700;
	wire [4-1:0] node13701;
	wire [4-1:0] node13704;
	wire [4-1:0] node13707;
	wire [4-1:0] node13709;
	wire [4-1:0] node13712;
	wire [4-1:0] node13713;
	wire [4-1:0] node13716;
	wire [4-1:0] node13719;
	wire [4-1:0] node13720;
	wire [4-1:0] node13721;
	wire [4-1:0] node13722;
	wire [4-1:0] node13725;
	wire [4-1:0] node13728;
	wire [4-1:0] node13730;
	wire [4-1:0] node13733;
	wire [4-1:0] node13734;
	wire [4-1:0] node13736;
	wire [4-1:0] node13740;
	wire [4-1:0] node13741;
	wire [4-1:0] node13742;
	wire [4-1:0] node13743;
	wire [4-1:0] node13744;
	wire [4-1:0] node13747;
	wire [4-1:0] node13750;
	wire [4-1:0] node13751;
	wire [4-1:0] node13752;
	wire [4-1:0] node13755;
	wire [4-1:0] node13758;
	wire [4-1:0] node13759;
	wire [4-1:0] node13763;
	wire [4-1:0] node13765;
	wire [4-1:0] node13766;
	wire [4-1:0] node13769;
	wire [4-1:0] node13772;
	wire [4-1:0] node13773;
	wire [4-1:0] node13774;
	wire [4-1:0] node13776;
	wire [4-1:0] node13779;
	wire [4-1:0] node13782;
	wire [4-1:0] node13783;
	wire [4-1:0] node13784;
	wire [4-1:0] node13785;
	wire [4-1:0] node13788;
	wire [4-1:0] node13791;
	wire [4-1:0] node13792;
	wire [4-1:0] node13795;
	wire [4-1:0] node13798;
	wire [4-1:0] node13799;
	wire [4-1:0] node13801;
	wire [4-1:0] node13804;
	wire [4-1:0] node13807;
	wire [4-1:0] node13808;
	wire [4-1:0] node13809;
	wire [4-1:0] node13810;
	wire [4-1:0] node13811;
	wire [4-1:0] node13812;
	wire [4-1:0] node13815;
	wire [4-1:0] node13818;
	wire [4-1:0] node13819;
	wire [4-1:0] node13820;
	wire [4-1:0] node13824;
	wire [4-1:0] node13825;
	wire [4-1:0] node13828;
	wire [4-1:0] node13831;
	wire [4-1:0] node13832;
	wire [4-1:0] node13833;
	wire [4-1:0] node13834;
	wire [4-1:0] node13837;
	wire [4-1:0] node13840;
	wire [4-1:0] node13841;
	wire [4-1:0] node13844;
	wire [4-1:0] node13847;
	wire [4-1:0] node13848;
	wire [4-1:0] node13851;
	wire [4-1:0] node13854;
	wire [4-1:0] node13855;
	wire [4-1:0] node13856;
	wire [4-1:0] node13858;
	wire [4-1:0] node13861;
	wire [4-1:0] node13862;
	wire [4-1:0] node13864;
	wire [4-1:0] node13867;
	wire [4-1:0] node13869;
	wire [4-1:0] node13872;
	wire [4-1:0] node13873;
	wire [4-1:0] node13874;
	wire [4-1:0] node13878;
	wire [4-1:0] node13879;
	wire [4-1:0] node13880;
	wire [4-1:0] node13883;
	wire [4-1:0] node13886;
	wire [4-1:0] node13887;
	wire [4-1:0] node13891;
	wire [4-1:0] node13892;
	wire [4-1:0] node13893;
	wire [4-1:0] node13894;
	wire [4-1:0] node13895;
	wire [4-1:0] node13898;
	wire [4-1:0] node13899;
	wire [4-1:0] node13902;
	wire [4-1:0] node13905;
	wire [4-1:0] node13906;
	wire [4-1:0] node13909;
	wire [4-1:0] node13912;
	wire [4-1:0] node13913;
	wire [4-1:0] node13914;
	wire [4-1:0] node13915;
	wire [4-1:0] node13918;
	wire [4-1:0] node13922;
	wire [4-1:0] node13923;
	wire [4-1:0] node13925;
	wire [4-1:0] node13928;
	wire [4-1:0] node13931;
	wire [4-1:0] node13932;
	wire [4-1:0] node13933;
	wire [4-1:0] node13935;
	wire [4-1:0] node13938;
	wire [4-1:0] node13939;
	wire [4-1:0] node13940;
	wire [4-1:0] node13945;
	wire [4-1:0] node13946;
	wire [4-1:0] node13947;
	wire [4-1:0] node13949;
	wire [4-1:0] node13952;
	wire [4-1:0] node13953;
	wire [4-1:0] node13956;
	wire [4-1:0] node13959;
	wire [4-1:0] node13960;
	wire [4-1:0] node13961;
	wire [4-1:0] node13965;
	wire [4-1:0] node13968;
	wire [4-1:0] node13969;
	wire [4-1:0] node13970;
	wire [4-1:0] node13971;
	wire [4-1:0] node13972;
	wire [4-1:0] node13973;
	wire [4-1:0] node13974;
	wire [4-1:0] node13975;
	wire [4-1:0] node13976;
	wire [4-1:0] node13979;
	wire [4-1:0] node13982;
	wire [4-1:0] node13983;
	wire [4-1:0] node13987;
	wire [4-1:0] node13988;
	wire [4-1:0] node13989;
	wire [4-1:0] node13990;
	wire [4-1:0] node13995;
	wire [4-1:0] node13996;
	wire [4-1:0] node13997;
	wire [4-1:0] node14002;
	wire [4-1:0] node14003;
	wire [4-1:0] node14004;
	wire [4-1:0] node14006;
	wire [4-1:0] node14007;
	wire [4-1:0] node14010;
	wire [4-1:0] node14013;
	wire [4-1:0] node14014;
	wire [4-1:0] node14016;
	wire [4-1:0] node14019;
	wire [4-1:0] node14021;
	wire [4-1:0] node14024;
	wire [4-1:0] node14025;
	wire [4-1:0] node14026;
	wire [4-1:0] node14027;
	wire [4-1:0] node14030;
	wire [4-1:0] node14033;
	wire [4-1:0] node14034;
	wire [4-1:0] node14038;
	wire [4-1:0] node14039;
	wire [4-1:0] node14043;
	wire [4-1:0] node14044;
	wire [4-1:0] node14045;
	wire [4-1:0] node14046;
	wire [4-1:0] node14048;
	wire [4-1:0] node14051;
	wire [4-1:0] node14052;
	wire [4-1:0] node14054;
	wire [4-1:0] node14058;
	wire [4-1:0] node14059;
	wire [4-1:0] node14060;
	wire [4-1:0] node14063;
	wire [4-1:0] node14066;
	wire [4-1:0] node14067;
	wire [4-1:0] node14071;
	wire [4-1:0] node14072;
	wire [4-1:0] node14073;
	wire [4-1:0] node14074;
	wire [4-1:0] node14077;
	wire [4-1:0] node14080;
	wire [4-1:0] node14081;
	wire [4-1:0] node14082;
	wire [4-1:0] node14085;
	wire [4-1:0] node14088;
	wire [4-1:0] node14089;
	wire [4-1:0] node14092;
	wire [4-1:0] node14095;
	wire [4-1:0] node14096;
	wire [4-1:0] node14097;
	wire [4-1:0] node14100;
	wire [4-1:0] node14103;
	wire [4-1:0] node14104;
	wire [4-1:0] node14105;
	wire [4-1:0] node14108;
	wire [4-1:0] node14111;
	wire [4-1:0] node14113;
	wire [4-1:0] node14116;
	wire [4-1:0] node14117;
	wire [4-1:0] node14118;
	wire [4-1:0] node14119;
	wire [4-1:0] node14120;
	wire [4-1:0] node14123;
	wire [4-1:0] node14125;
	wire [4-1:0] node14128;
	wire [4-1:0] node14129;
	wire [4-1:0] node14130;
	wire [4-1:0] node14134;
	wire [4-1:0] node14135;
	wire [4-1:0] node14138;
	wire [4-1:0] node14141;
	wire [4-1:0] node14142;
	wire [4-1:0] node14143;
	wire [4-1:0] node14145;
	wire [4-1:0] node14148;
	wire [4-1:0] node14149;
	wire [4-1:0] node14153;
	wire [4-1:0] node14154;
	wire [4-1:0] node14157;
	wire [4-1:0] node14158;
	wire [4-1:0] node14161;
	wire [4-1:0] node14164;
	wire [4-1:0] node14165;
	wire [4-1:0] node14166;
	wire [4-1:0] node14168;
	wire [4-1:0] node14171;
	wire [4-1:0] node14172;
	wire [4-1:0] node14174;
	wire [4-1:0] node14177;
	wire [4-1:0] node14178;
	wire [4-1:0] node14182;
	wire [4-1:0] node14183;
	wire [4-1:0] node14184;
	wire [4-1:0] node14186;
	wire [4-1:0] node14189;
	wire [4-1:0] node14191;
	wire [4-1:0] node14194;
	wire [4-1:0] node14195;
	wire [4-1:0] node14196;
	wire [4-1:0] node14200;
	wire [4-1:0] node14201;
	wire [4-1:0] node14205;
	wire [4-1:0] node14206;
	wire [4-1:0] node14207;
	wire [4-1:0] node14208;
	wire [4-1:0] node14209;
	wire [4-1:0] node14210;
	wire [4-1:0] node14213;
	wire [4-1:0] node14216;
	wire [4-1:0] node14217;
	wire [4-1:0] node14218;
	wire [4-1:0] node14221;
	wire [4-1:0] node14224;
	wire [4-1:0] node14226;
	wire [4-1:0] node14229;
	wire [4-1:0] node14230;
	wire [4-1:0] node14231;
	wire [4-1:0] node14232;
	wire [4-1:0] node14234;
	wire [4-1:0] node14237;
	wire [4-1:0] node14240;
	wire [4-1:0] node14241;
	wire [4-1:0] node14245;
	wire [4-1:0] node14246;
	wire [4-1:0] node14248;
	wire [4-1:0] node14249;
	wire [4-1:0] node14252;
	wire [4-1:0] node14255;
	wire [4-1:0] node14256;
	wire [4-1:0] node14257;
	wire [4-1:0] node14260;
	wire [4-1:0] node14263;
	wire [4-1:0] node14265;
	wire [4-1:0] node14268;
	wire [4-1:0] node14269;
	wire [4-1:0] node14270;
	wire [4-1:0] node14271;
	wire [4-1:0] node14273;
	wire [4-1:0] node14276;
	wire [4-1:0] node14279;
	wire [4-1:0] node14280;
	wire [4-1:0] node14283;
	wire [4-1:0] node14285;
	wire [4-1:0] node14288;
	wire [4-1:0] node14289;
	wire [4-1:0] node14290;
	wire [4-1:0] node14291;
	wire [4-1:0] node14294;
	wire [4-1:0] node14297;
	wire [4-1:0] node14299;
	wire [4-1:0] node14302;
	wire [4-1:0] node14303;
	wire [4-1:0] node14304;
	wire [4-1:0] node14307;
	wire [4-1:0] node14310;
	wire [4-1:0] node14311;
	wire [4-1:0] node14312;
	wire [4-1:0] node14315;
	wire [4-1:0] node14318;
	wire [4-1:0] node14319;
	wire [4-1:0] node14322;
	wire [4-1:0] node14325;
	wire [4-1:0] node14326;
	wire [4-1:0] node14327;
	wire [4-1:0] node14328;
	wire [4-1:0] node14329;
	wire [4-1:0] node14330;
	wire [4-1:0] node14332;
	wire [4-1:0] node14335;
	wire [4-1:0] node14337;
	wire [4-1:0] node14340;
	wire [4-1:0] node14342;
	wire [4-1:0] node14345;
	wire [4-1:0] node14346;
	wire [4-1:0] node14347;
	wire [4-1:0] node14350;
	wire [4-1:0] node14353;
	wire [4-1:0] node14354;
	wire [4-1:0] node14355;
	wire [4-1:0] node14359;
	wire [4-1:0] node14361;
	wire [4-1:0] node14364;
	wire [4-1:0] node14365;
	wire [4-1:0] node14366;
	wire [4-1:0] node14367;
	wire [4-1:0] node14370;
	wire [4-1:0] node14373;
	wire [4-1:0] node14375;
	wire [4-1:0] node14378;
	wire [4-1:0] node14379;
	wire [4-1:0] node14380;
	wire [4-1:0] node14383;
	wire [4-1:0] node14386;
	wire [4-1:0] node14387;
	wire [4-1:0] node14391;
	wire [4-1:0] node14392;
	wire [4-1:0] node14393;
	wire [4-1:0] node14394;
	wire [4-1:0] node14396;
	wire [4-1:0] node14399;
	wire [4-1:0] node14400;
	wire [4-1:0] node14402;
	wire [4-1:0] node14405;
	wire [4-1:0] node14406;
	wire [4-1:0] node14409;
	wire [4-1:0] node14412;
	wire [4-1:0] node14413;
	wire [4-1:0] node14414;
	wire [4-1:0] node14417;
	wire [4-1:0] node14420;
	wire [4-1:0] node14421;
	wire [4-1:0] node14422;
	wire [4-1:0] node14425;
	wire [4-1:0] node14429;
	wire [4-1:0] node14430;
	wire [4-1:0] node14431;
	wire [4-1:0] node14434;
	wire [4-1:0] node14435;
	wire [4-1:0] node14436;
	wire [4-1:0] node14440;
	wire [4-1:0] node14441;
	wire [4-1:0] node14445;
	wire [4-1:0] node14446;
	wire [4-1:0] node14447;
	wire [4-1:0] node14450;
	wire [4-1:0] node14453;
	wire [4-1:0] node14456;
	wire [4-1:0] node14457;
	wire [4-1:0] node14458;
	wire [4-1:0] node14459;
	wire [4-1:0] node14460;
	wire [4-1:0] node14461;
	wire [4-1:0] node14462;
	wire [4-1:0] node14464;
	wire [4-1:0] node14467;
	wire [4-1:0] node14469;
	wire [4-1:0] node14471;
	wire [4-1:0] node14474;
	wire [4-1:0] node14475;
	wire [4-1:0] node14476;
	wire [4-1:0] node14480;
	wire [4-1:0] node14483;
	wire [4-1:0] node14484;
	wire [4-1:0] node14485;
	wire [4-1:0] node14486;
	wire [4-1:0] node14489;
	wire [4-1:0] node14492;
	wire [4-1:0] node14493;
	wire [4-1:0] node14495;
	wire [4-1:0] node14499;
	wire [4-1:0] node14500;
	wire [4-1:0] node14501;
	wire [4-1:0] node14503;
	wire [4-1:0] node14507;
	wire [4-1:0] node14508;
	wire [4-1:0] node14509;
	wire [4-1:0] node14512;
	wire [4-1:0] node14516;
	wire [4-1:0] node14517;
	wire [4-1:0] node14518;
	wire [4-1:0] node14519;
	wire [4-1:0] node14522;
	wire [4-1:0] node14524;
	wire [4-1:0] node14527;
	wire [4-1:0] node14528;
	wire [4-1:0] node14529;
	wire [4-1:0] node14533;
	wire [4-1:0] node14536;
	wire [4-1:0] node14537;
	wire [4-1:0] node14538;
	wire [4-1:0] node14539;
	wire [4-1:0] node14543;
	wire [4-1:0] node14544;
	wire [4-1:0] node14547;
	wire [4-1:0] node14550;
	wire [4-1:0] node14551;
	wire [4-1:0] node14552;
	wire [4-1:0] node14555;
	wire [4-1:0] node14558;
	wire [4-1:0] node14559;
	wire [4-1:0] node14561;
	wire [4-1:0] node14564;
	wire [4-1:0] node14565;
	wire [4-1:0] node14569;
	wire [4-1:0] node14570;
	wire [4-1:0] node14571;
	wire [4-1:0] node14572;
	wire [4-1:0] node14574;
	wire [4-1:0] node14576;
	wire [4-1:0] node14579;
	wire [4-1:0] node14580;
	wire [4-1:0] node14582;
	wire [4-1:0] node14585;
	wire [4-1:0] node14588;
	wire [4-1:0] node14589;
	wire [4-1:0] node14590;
	wire [4-1:0] node14591;
	wire [4-1:0] node14595;
	wire [4-1:0] node14596;
	wire [4-1:0] node14600;
	wire [4-1:0] node14601;
	wire [4-1:0] node14603;
	wire [4-1:0] node14604;
	wire [4-1:0] node14608;
	wire [4-1:0] node14611;
	wire [4-1:0] node14612;
	wire [4-1:0] node14613;
	wire [4-1:0] node14614;
	wire [4-1:0] node14615;
	wire [4-1:0] node14619;
	wire [4-1:0] node14622;
	wire [4-1:0] node14623;
	wire [4-1:0] node14626;
	wire [4-1:0] node14627;
	wire [4-1:0] node14631;
	wire [4-1:0] node14632;
	wire [4-1:0] node14633;
	wire [4-1:0] node14634;
	wire [4-1:0] node14635;
	wire [4-1:0] node14638;
	wire [4-1:0] node14643;
	wire [4-1:0] node14644;
	wire [4-1:0] node14646;
	wire [4-1:0] node14647;
	wire [4-1:0] node14650;
	wire [4-1:0] node14654;
	wire [4-1:0] node14655;
	wire [4-1:0] node14656;
	wire [4-1:0] node14657;
	wire [4-1:0] node14658;
	wire [4-1:0] node14659;
	wire [4-1:0] node14660;
	wire [4-1:0] node14662;
	wire [4-1:0] node14665;
	wire [4-1:0] node14666;
	wire [4-1:0] node14670;
	wire [4-1:0] node14671;
	wire [4-1:0] node14674;
	wire [4-1:0] node14677;
	wire [4-1:0] node14678;
	wire [4-1:0] node14679;
	wire [4-1:0] node14680;
	wire [4-1:0] node14684;
	wire [4-1:0] node14685;
	wire [4-1:0] node14689;
	wire [4-1:0] node14690;
	wire [4-1:0] node14693;
	wire [4-1:0] node14696;
	wire [4-1:0] node14697;
	wire [4-1:0] node14698;
	wire [4-1:0] node14700;
	wire [4-1:0] node14701;
	wire [4-1:0] node14704;
	wire [4-1:0] node14707;
	wire [4-1:0] node14708;
	wire [4-1:0] node14711;
	wire [4-1:0] node14714;
	wire [4-1:0] node14715;
	wire [4-1:0] node14716;
	wire [4-1:0] node14718;
	wire [4-1:0] node14721;
	wire [4-1:0] node14724;
	wire [4-1:0] node14725;
	wire [4-1:0] node14727;
	wire [4-1:0] node14731;
	wire [4-1:0] node14732;
	wire [4-1:0] node14733;
	wire [4-1:0] node14734;
	wire [4-1:0] node14735;
	wire [4-1:0] node14736;
	wire [4-1:0] node14741;
	wire [4-1:0] node14743;
	wire [4-1:0] node14745;
	wire [4-1:0] node14748;
	wire [4-1:0] node14749;
	wire [4-1:0] node14751;
	wire [4-1:0] node14752;
	wire [4-1:0] node14756;
	wire [4-1:0] node14757;
	wire [4-1:0] node14758;
	wire [4-1:0] node14762;
	wire [4-1:0] node14763;
	wire [4-1:0] node14767;
	wire [4-1:0] node14768;
	wire [4-1:0] node14769;
	wire [4-1:0] node14770;
	wire [4-1:0] node14771;
	wire [4-1:0] node14776;
	wire [4-1:0] node14777;
	wire [4-1:0] node14780;
	wire [4-1:0] node14783;
	wire [4-1:0] node14784;
	wire [4-1:0] node14785;
	wire [4-1:0] node14786;
	wire [4-1:0] node14790;
	wire [4-1:0] node14793;
	wire [4-1:0] node14794;
	wire [4-1:0] node14795;
	wire [4-1:0] node14798;
	wire [4-1:0] node14802;
	wire [4-1:0] node14803;
	wire [4-1:0] node14804;
	wire [4-1:0] node14805;
	wire [4-1:0] node14806;
	wire [4-1:0] node14807;
	wire [4-1:0] node14810;
	wire [4-1:0] node14812;
	wire [4-1:0] node14815;
	wire [4-1:0] node14816;
	wire [4-1:0] node14820;
	wire [4-1:0] node14821;
	wire [4-1:0] node14822;
	wire [4-1:0] node14826;
	wire [4-1:0] node14827;
	wire [4-1:0] node14830;
	wire [4-1:0] node14833;
	wire [4-1:0] node14834;
	wire [4-1:0] node14835;
	wire [4-1:0] node14836;
	wire [4-1:0] node14840;
	wire [4-1:0] node14841;
	wire [4-1:0] node14844;
	wire [4-1:0] node14847;
	wire [4-1:0] node14848;
	wire [4-1:0] node14849;
	wire [4-1:0] node14852;
	wire [4-1:0] node14855;
	wire [4-1:0] node14856;
	wire [4-1:0] node14860;
	wire [4-1:0] node14861;
	wire [4-1:0] node14862;
	wire [4-1:0] node14863;
	wire [4-1:0] node14864;
	wire [4-1:0] node14868;
	wire [4-1:0] node14869;
	wire [4-1:0] node14873;
	wire [4-1:0] node14874;
	wire [4-1:0] node14875;
	wire [4-1:0] node14879;
	wire [4-1:0] node14880;
	wire [4-1:0] node14884;
	wire [4-1:0] node14885;
	wire [4-1:0] node14886;
	wire [4-1:0] node14887;
	wire [4-1:0] node14891;
	wire [4-1:0] node14892;
	wire [4-1:0] node14893;
	wire [4-1:0] node14898;
	wire [4-1:0] node14899;
	wire [4-1:0] node14900;
	wire [4-1:0] node14901;
	wire [4-1:0] node14904;
	wire [4-1:0] node14908;
	wire [4-1:0] node14909;
	wire [4-1:0] node14910;
	wire [4-1:0] node14913;
	wire [4-1:0] node14916;
	wire [4-1:0] node14917;
	wire [4-1:0] node14920;
	wire [4-1:0] node14923;
	wire [4-1:0] node14924;
	wire [4-1:0] node14925;
	wire [4-1:0] node14926;
	wire [4-1:0] node14927;
	wire [4-1:0] node14928;
	wire [4-1:0] node14929;
	wire [4-1:0] node14930;
	wire [4-1:0] node14931;
	wire [4-1:0] node14932;
	wire [4-1:0] node14933;
	wire [4-1:0] node14934;
	wire [4-1:0] node14936;
	wire [4-1:0] node14939;
	wire [4-1:0] node14941;
	wire [4-1:0] node14944;
	wire [4-1:0] node14945;
	wire [4-1:0] node14947;
	wire [4-1:0] node14950;
	wire [4-1:0] node14951;
	wire [4-1:0] node14955;
	wire [4-1:0] node14956;
	wire [4-1:0] node14957;
	wire [4-1:0] node14958;
	wire [4-1:0] node14961;
	wire [4-1:0] node14963;
	wire [4-1:0] node14966;
	wire [4-1:0] node14967;
	wire [4-1:0] node14971;
	wire [4-1:0] node14972;
	wire [4-1:0] node14973;
	wire [4-1:0] node14974;
	wire [4-1:0] node14978;
	wire [4-1:0] node14981;
	wire [4-1:0] node14982;
	wire [4-1:0] node14983;
	wire [4-1:0] node14986;
	wire [4-1:0] node14990;
	wire [4-1:0] node14991;
	wire [4-1:0] node14992;
	wire [4-1:0] node14993;
	wire [4-1:0] node14995;
	wire [4-1:0] node14996;
	wire [4-1:0] node14999;
	wire [4-1:0] node15002;
	wire [4-1:0] node15003;
	wire [4-1:0] node15006;
	wire [4-1:0] node15009;
	wire [4-1:0] node15010;
	wire [4-1:0] node15012;
	wire [4-1:0] node15015;
	wire [4-1:0] node15016;
	wire [4-1:0] node15017;
	wire [4-1:0] node15021;
	wire [4-1:0] node15023;
	wire [4-1:0] node15026;
	wire [4-1:0] node15027;
	wire [4-1:0] node15028;
	wire [4-1:0] node15029;
	wire [4-1:0] node15032;
	wire [4-1:0] node15036;
	wire [4-1:0] node15037;
	wire [4-1:0] node15038;
	wire [4-1:0] node15039;
	wire [4-1:0] node15042;
	wire [4-1:0] node15046;
	wire [4-1:0] node15047;
	wire [4-1:0] node15050;
	wire [4-1:0] node15051;
	wire [4-1:0] node15055;
	wire [4-1:0] node15056;
	wire [4-1:0] node15057;
	wire [4-1:0] node15058;
	wire [4-1:0] node15059;
	wire [4-1:0] node15061;
	wire [4-1:0] node15064;
	wire [4-1:0] node15065;
	wire [4-1:0] node15068;
	wire [4-1:0] node15071;
	wire [4-1:0] node15072;
	wire [4-1:0] node15075;
	wire [4-1:0] node15076;
	wire [4-1:0] node15078;
	wire [4-1:0] node15082;
	wire [4-1:0] node15083;
	wire [4-1:0] node15084;
	wire [4-1:0] node15085;
	wire [4-1:0] node15086;
	wire [4-1:0] node15089;
	wire [4-1:0] node15092;
	wire [4-1:0] node15093;
	wire [4-1:0] node15097;
	wire [4-1:0] node15098;
	wire [4-1:0] node15101;
	wire [4-1:0] node15102;
	wire [4-1:0] node15105;
	wire [4-1:0] node15108;
	wire [4-1:0] node15109;
	wire [4-1:0] node15110;
	wire [4-1:0] node15111;
	wire [4-1:0] node15116;
	wire [4-1:0] node15118;
	wire [4-1:0] node15119;
	wire [4-1:0] node15123;
	wire [4-1:0] node15124;
	wire [4-1:0] node15125;
	wire [4-1:0] node15126;
	wire [4-1:0] node15127;
	wire [4-1:0] node15131;
	wire [4-1:0] node15133;
	wire [4-1:0] node15134;
	wire [4-1:0] node15137;
	wire [4-1:0] node15140;
	wire [4-1:0] node15141;
	wire [4-1:0] node15142;
	wire [4-1:0] node15145;
	wire [4-1:0] node15149;
	wire [4-1:0] node15150;
	wire [4-1:0] node15151;
	wire [4-1:0] node15152;
	wire [4-1:0] node15153;
	wire [4-1:0] node15156;
	wire [4-1:0] node15160;
	wire [4-1:0] node15161;
	wire [4-1:0] node15162;
	wire [4-1:0] node15165;
	wire [4-1:0] node15168;
	wire [4-1:0] node15171;
	wire [4-1:0] node15172;
	wire [4-1:0] node15173;
	wire [4-1:0] node15175;
	wire [4-1:0] node15178;
	wire [4-1:0] node15179;
	wire [4-1:0] node15183;
	wire [4-1:0] node15185;
	wire [4-1:0] node15187;
	wire [4-1:0] node15190;
	wire [4-1:0] node15191;
	wire [4-1:0] node15192;
	wire [4-1:0] node15193;
	wire [4-1:0] node15194;
	wire [4-1:0] node15195;
	wire [4-1:0] node15196;
	wire [4-1:0] node15197;
	wire [4-1:0] node15201;
	wire [4-1:0] node15202;
	wire [4-1:0] node15205;
	wire [4-1:0] node15208;
	wire [4-1:0] node15209;
	wire [4-1:0] node15212;
	wire [4-1:0] node15215;
	wire [4-1:0] node15216;
	wire [4-1:0] node15218;
	wire [4-1:0] node15219;
	wire [4-1:0] node15222;
	wire [4-1:0] node15225;
	wire [4-1:0] node15226;
	wire [4-1:0] node15227;
	wire [4-1:0] node15232;
	wire [4-1:0] node15233;
	wire [4-1:0] node15234;
	wire [4-1:0] node15236;
	wire [4-1:0] node15239;
	wire [4-1:0] node15240;
	wire [4-1:0] node15243;
	wire [4-1:0] node15246;
	wire [4-1:0] node15248;
	wire [4-1:0] node15249;
	wire [4-1:0] node15250;
	wire [4-1:0] node15253;
	wire [4-1:0] node15256;
	wire [4-1:0] node15257;
	wire [4-1:0] node15260;
	wire [4-1:0] node15263;
	wire [4-1:0] node15264;
	wire [4-1:0] node15265;
	wire [4-1:0] node15266;
	wire [4-1:0] node15267;
	wire [4-1:0] node15270;
	wire [4-1:0] node15273;
	wire [4-1:0] node15275;
	wire [4-1:0] node15276;
	wire [4-1:0] node15279;
	wire [4-1:0] node15282;
	wire [4-1:0] node15283;
	wire [4-1:0] node15284;
	wire [4-1:0] node15285;
	wire [4-1:0] node15288;
	wire [4-1:0] node15292;
	wire [4-1:0] node15293;
	wire [4-1:0] node15294;
	wire [4-1:0] node15297;
	wire [4-1:0] node15301;
	wire [4-1:0] node15302;
	wire [4-1:0] node15303;
	wire [4-1:0] node15304;
	wire [4-1:0] node15308;
	wire [4-1:0] node15309;
	wire [4-1:0] node15313;
	wire [4-1:0] node15314;
	wire [4-1:0] node15315;
	wire [4-1:0] node15316;
	wire [4-1:0] node15319;
	wire [4-1:0] node15322;
	wire [4-1:0] node15323;
	wire [4-1:0] node15326;
	wire [4-1:0] node15329;
	wire [4-1:0] node15330;
	wire [4-1:0] node15331;
	wire [4-1:0] node15334;
	wire [4-1:0] node15337;
	wire [4-1:0] node15338;
	wire [4-1:0] node15341;
	wire [4-1:0] node15344;
	wire [4-1:0] node15345;
	wire [4-1:0] node15346;
	wire [4-1:0] node15347;
	wire [4-1:0] node15349;
	wire [4-1:0] node15352;
	wire [4-1:0] node15353;
	wire [4-1:0] node15355;
	wire [4-1:0] node15358;
	wire [4-1:0] node15359;
	wire [4-1:0] node15362;
	wire [4-1:0] node15365;
	wire [4-1:0] node15366;
	wire [4-1:0] node15367;
	wire [4-1:0] node15368;
	wire [4-1:0] node15370;
	wire [4-1:0] node15373;
	wire [4-1:0] node15376;
	wire [4-1:0] node15377;
	wire [4-1:0] node15381;
	wire [4-1:0] node15382;
	wire [4-1:0] node15383;
	wire [4-1:0] node15385;
	wire [4-1:0] node15388;
	wire [4-1:0] node15390;
	wire [4-1:0] node15393;
	wire [4-1:0] node15394;
	wire [4-1:0] node15395;
	wire [4-1:0] node15400;
	wire [4-1:0] node15401;
	wire [4-1:0] node15402;
	wire [4-1:0] node15403;
	wire [4-1:0] node15404;
	wire [4-1:0] node15406;
	wire [4-1:0] node15409;
	wire [4-1:0] node15412;
	wire [4-1:0] node15415;
	wire [4-1:0] node15416;
	wire [4-1:0] node15417;
	wire [4-1:0] node15418;
	wire [4-1:0] node15421;
	wire [4-1:0] node15424;
	wire [4-1:0] node15425;
	wire [4-1:0] node15428;
	wire [4-1:0] node15431;
	wire [4-1:0] node15433;
	wire [4-1:0] node15434;
	wire [4-1:0] node15437;
	wire [4-1:0] node15440;
	wire [4-1:0] node15441;
	wire [4-1:0] node15442;
	wire [4-1:0] node15444;
	wire [4-1:0] node15445;
	wire [4-1:0] node15449;
	wire [4-1:0] node15451;
	wire [4-1:0] node15453;
	wire [4-1:0] node15456;
	wire [4-1:0] node15457;
	wire [4-1:0] node15458;
	wire [4-1:0] node15462;
	wire [4-1:0] node15463;
	wire [4-1:0] node15465;
	wire [4-1:0] node15468;
	wire [4-1:0] node15469;
	wire [4-1:0] node15473;
	wire [4-1:0] node15474;
	wire [4-1:0] node15475;
	wire [4-1:0] node15476;
	wire [4-1:0] node15477;
	wire [4-1:0] node15478;
	wire [4-1:0] node15479;
	wire [4-1:0] node15482;
	wire [4-1:0] node15485;
	wire [4-1:0] node15486;
	wire [4-1:0] node15489;
	wire [4-1:0] node15492;
	wire [4-1:0] node15493;
	wire [4-1:0] node15496;
	wire [4-1:0] node15499;
	wire [4-1:0] node15500;
	wire [4-1:0] node15501;
	wire [4-1:0] node15502;
	wire [4-1:0] node15505;
	wire [4-1:0] node15508;
	wire [4-1:0] node15509;
	wire [4-1:0] node15512;
	wire [4-1:0] node15515;
	wire [4-1:0] node15516;
	wire [4-1:0] node15517;
	wire [4-1:0] node15518;
	wire [4-1:0] node15521;
	wire [4-1:0] node15524;
	wire [4-1:0] node15526;
	wire [4-1:0] node15529;
	wire [4-1:0] node15530;
	wire [4-1:0] node15531;
	wire [4-1:0] node15535;
	wire [4-1:0] node15536;
	wire [4-1:0] node15537;
	wire [4-1:0] node15541;
	wire [4-1:0] node15543;
	wire [4-1:0] node15546;
	wire [4-1:0] node15547;
	wire [4-1:0] node15548;
	wire [4-1:0] node15549;
	wire [4-1:0] node15550;
	wire [4-1:0] node15551;
	wire [4-1:0] node15554;
	wire [4-1:0] node15557;
	wire [4-1:0] node15558;
	wire [4-1:0] node15561;
	wire [4-1:0] node15564;
	wire [4-1:0] node15565;
	wire [4-1:0] node15567;
	wire [4-1:0] node15568;
	wire [4-1:0] node15571;
	wire [4-1:0] node15574;
	wire [4-1:0] node15575;
	wire [4-1:0] node15578;
	wire [4-1:0] node15581;
	wire [4-1:0] node15582;
	wire [4-1:0] node15584;
	wire [4-1:0] node15585;
	wire [4-1:0] node15588;
	wire [4-1:0] node15591;
	wire [4-1:0] node15592;
	wire [4-1:0] node15595;
	wire [4-1:0] node15598;
	wire [4-1:0] node15599;
	wire [4-1:0] node15600;
	wire [4-1:0] node15601;
	wire [4-1:0] node15602;
	wire [4-1:0] node15605;
	wire [4-1:0] node15608;
	wire [4-1:0] node15609;
	wire [4-1:0] node15612;
	wire [4-1:0] node15615;
	wire [4-1:0] node15616;
	wire [4-1:0] node15619;
	wire [4-1:0] node15622;
	wire [4-1:0] node15623;
	wire [4-1:0] node15625;
	wire [4-1:0] node15627;
	wire [4-1:0] node15630;
	wire [4-1:0] node15631;
	wire [4-1:0] node15634;
	wire [4-1:0] node15637;
	wire [4-1:0] node15638;
	wire [4-1:0] node15639;
	wire [4-1:0] node15640;
	wire [4-1:0] node15641;
	wire [4-1:0] node15644;
	wire [4-1:0] node15647;
	wire [4-1:0] node15648;
	wire [4-1:0] node15649;
	wire [4-1:0] node15650;
	wire [4-1:0] node15654;
	wire [4-1:0] node15655;
	wire [4-1:0] node15659;
	wire [4-1:0] node15660;
	wire [4-1:0] node15663;
	wire [4-1:0] node15666;
	wire [4-1:0] node15667;
	wire [4-1:0] node15668;
	wire [4-1:0] node15671;
	wire [4-1:0] node15674;
	wire [4-1:0] node15675;
	wire [4-1:0] node15678;
	wire [4-1:0] node15681;
	wire [4-1:0] node15682;
	wire [4-1:0] node15683;
	wire [4-1:0] node15684;
	wire [4-1:0] node15685;
	wire [4-1:0] node15686;
	wire [4-1:0] node15689;
	wire [4-1:0] node15692;
	wire [4-1:0] node15693;
	wire [4-1:0] node15696;
	wire [4-1:0] node15699;
	wire [4-1:0] node15700;
	wire [4-1:0] node15701;
	wire [4-1:0] node15705;
	wire [4-1:0] node15706;
	wire [4-1:0] node15709;
	wire [4-1:0] node15712;
	wire [4-1:0] node15713;
	wire [4-1:0] node15714;
	wire [4-1:0] node15717;
	wire [4-1:0] node15718;
	wire [4-1:0] node15719;
	wire [4-1:0] node15724;
	wire [4-1:0] node15725;
	wire [4-1:0] node15726;
	wire [4-1:0] node15729;
	wire [4-1:0] node15733;
	wire [4-1:0] node15734;
	wire [4-1:0] node15735;
	wire [4-1:0] node15736;
	wire [4-1:0] node15739;
	wire [4-1:0] node15742;
	wire [4-1:0] node15743;
	wire [4-1:0] node15746;
	wire [4-1:0] node15749;
	wire [4-1:0] node15750;
	wire [4-1:0] node15751;
	wire [4-1:0] node15752;
	wire [4-1:0] node15753;
	wire [4-1:0] node15756;
	wire [4-1:0] node15760;
	wire [4-1:0] node15762;
	wire [4-1:0] node15765;
	wire [4-1:0] node15766;
	wire [4-1:0] node15769;
	wire [4-1:0] node15772;
	wire [4-1:0] node15773;
	wire [4-1:0] node15774;
	wire [4-1:0] node15775;
	wire [4-1:0] node15776;
	wire [4-1:0] node15777;
	wire [4-1:0] node15778;
	wire [4-1:0] node15780;
	wire [4-1:0] node15781;
	wire [4-1:0] node15784;
	wire [4-1:0] node15787;
	wire [4-1:0] node15788;
	wire [4-1:0] node15789;
	wire [4-1:0] node15790;
	wire [4-1:0] node15794;
	wire [4-1:0] node15795;
	wire [4-1:0] node15800;
	wire [4-1:0] node15801;
	wire [4-1:0] node15802;
	wire [4-1:0] node15803;
	wire [4-1:0] node15804;
	wire [4-1:0] node15808;
	wire [4-1:0] node15811;
	wire [4-1:0] node15813;
	wire [4-1:0] node15816;
	wire [4-1:0] node15818;
	wire [4-1:0] node15821;
	wire [4-1:0] node15822;
	wire [4-1:0] node15823;
	wire [4-1:0] node15824;
	wire [4-1:0] node15825;
	wire [4-1:0] node15827;
	wire [4-1:0] node15831;
	wire [4-1:0] node15834;
	wire [4-1:0] node15835;
	wire [4-1:0] node15838;
	wire [4-1:0] node15839;
	wire [4-1:0] node15842;
	wire [4-1:0] node15845;
	wire [4-1:0] node15846;
	wire [4-1:0] node15847;
	wire [4-1:0] node15848;
	wire [4-1:0] node15849;
	wire [4-1:0] node15854;
	wire [4-1:0] node15856;
	wire [4-1:0] node15859;
	wire [4-1:0] node15860;
	wire [4-1:0] node15861;
	wire [4-1:0] node15862;
	wire [4-1:0] node15866;
	wire [4-1:0] node15869;
	wire [4-1:0] node15870;
	wire [4-1:0] node15873;
	wire [4-1:0] node15876;
	wire [4-1:0] node15877;
	wire [4-1:0] node15878;
	wire [4-1:0] node15879;
	wire [4-1:0] node15880;
	wire [4-1:0] node15881;
	wire [4-1:0] node15883;
	wire [4-1:0] node15887;
	wire [4-1:0] node15888;
	wire [4-1:0] node15891;
	wire [4-1:0] node15894;
	wire [4-1:0] node15895;
	wire [4-1:0] node15896;
	wire [4-1:0] node15897;
	wire [4-1:0] node15902;
	wire [4-1:0] node15904;
	wire [4-1:0] node15907;
	wire [4-1:0] node15908;
	wire [4-1:0] node15909;
	wire [4-1:0] node15912;
	wire [4-1:0] node15915;
	wire [4-1:0] node15916;
	wire [4-1:0] node15918;
	wire [4-1:0] node15920;
	wire [4-1:0] node15923;
	wire [4-1:0] node15924;
	wire [4-1:0] node15927;
	wire [4-1:0] node15930;
	wire [4-1:0] node15931;
	wire [4-1:0] node15932;
	wire [4-1:0] node15933;
	wire [4-1:0] node15934;
	wire [4-1:0] node15936;
	wire [4-1:0] node15939;
	wire [4-1:0] node15940;
	wire [4-1:0] node15944;
	wire [4-1:0] node15945;
	wire [4-1:0] node15947;
	wire [4-1:0] node15950;
	wire [4-1:0] node15951;
	wire [4-1:0] node15955;
	wire [4-1:0] node15956;
	wire [4-1:0] node15957;
	wire [4-1:0] node15958;
	wire [4-1:0] node15961;
	wire [4-1:0] node15965;
	wire [4-1:0] node15966;
	wire [4-1:0] node15969;
	wire [4-1:0] node15970;
	wire [4-1:0] node15973;
	wire [4-1:0] node15976;
	wire [4-1:0] node15977;
	wire [4-1:0] node15978;
	wire [4-1:0] node15979;
	wire [4-1:0] node15982;
	wire [4-1:0] node15985;
	wire [4-1:0] node15986;
	wire [4-1:0] node15987;
	wire [4-1:0] node15990;
	wire [4-1:0] node15994;
	wire [4-1:0] node15995;
	wire [4-1:0] node15997;
	wire [4-1:0] node15998;
	wire [4-1:0] node16002;
	wire [4-1:0] node16004;
	wire [4-1:0] node16007;
	wire [4-1:0] node16008;
	wire [4-1:0] node16009;
	wire [4-1:0] node16010;
	wire [4-1:0] node16011;
	wire [4-1:0] node16012;
	wire [4-1:0] node16013;
	wire [4-1:0] node16016;
	wire [4-1:0] node16019;
	wire [4-1:0] node16020;
	wire [4-1:0] node16021;
	wire [4-1:0] node16025;
	wire [4-1:0] node16026;
	wire [4-1:0] node16029;
	wire [4-1:0] node16032;
	wire [4-1:0] node16033;
	wire [4-1:0] node16034;
	wire [4-1:0] node16037;
	wire [4-1:0] node16040;
	wire [4-1:0] node16041;
	wire [4-1:0] node16044;
	wire [4-1:0] node16047;
	wire [4-1:0] node16048;
	wire [4-1:0] node16049;
	wire [4-1:0] node16050;
	wire [4-1:0] node16053;
	wire [4-1:0] node16056;
	wire [4-1:0] node16057;
	wire [4-1:0] node16058;
	wire [4-1:0] node16061;
	wire [4-1:0] node16065;
	wire [4-1:0] node16066;
	wire [4-1:0] node16068;
	wire [4-1:0] node16069;
	wire [4-1:0] node16073;
	wire [4-1:0] node16074;
	wire [4-1:0] node16075;
	wire [4-1:0] node16078;
	wire [4-1:0] node16081;
	wire [4-1:0] node16083;
	wire [4-1:0] node16086;
	wire [4-1:0] node16087;
	wire [4-1:0] node16088;
	wire [4-1:0] node16089;
	wire [4-1:0] node16090;
	wire [4-1:0] node16091;
	wire [4-1:0] node16094;
	wire [4-1:0] node16097;
	wire [4-1:0] node16098;
	wire [4-1:0] node16101;
	wire [4-1:0] node16104;
	wire [4-1:0] node16106;
	wire [4-1:0] node16109;
	wire [4-1:0] node16110;
	wire [4-1:0] node16111;
	wire [4-1:0] node16113;
	wire [4-1:0] node16116;
	wire [4-1:0] node16117;
	wire [4-1:0] node16120;
	wire [4-1:0] node16123;
	wire [4-1:0] node16124;
	wire [4-1:0] node16127;
	wire [4-1:0] node16130;
	wire [4-1:0] node16131;
	wire [4-1:0] node16133;
	wire [4-1:0] node16134;
	wire [4-1:0] node16135;
	wire [4-1:0] node16139;
	wire [4-1:0] node16141;
	wire [4-1:0] node16144;
	wire [4-1:0] node16145;
	wire [4-1:0] node16146;
	wire [4-1:0] node16147;
	wire [4-1:0] node16150;
	wire [4-1:0] node16153;
	wire [4-1:0] node16154;
	wire [4-1:0] node16157;
	wire [4-1:0] node16160;
	wire [4-1:0] node16161;
	wire [4-1:0] node16164;
	wire [4-1:0] node16167;
	wire [4-1:0] node16168;
	wire [4-1:0] node16169;
	wire [4-1:0] node16170;
	wire [4-1:0] node16171;
	wire [4-1:0] node16172;
	wire [4-1:0] node16173;
	wire [4-1:0] node16176;
	wire [4-1:0] node16179;
	wire [4-1:0] node16181;
	wire [4-1:0] node16184;
	wire [4-1:0] node16185;
	wire [4-1:0] node16186;
	wire [4-1:0] node16189;
	wire [4-1:0] node16192;
	wire [4-1:0] node16194;
	wire [4-1:0] node16197;
	wire [4-1:0] node16198;
	wire [4-1:0] node16199;
	wire [4-1:0] node16201;
	wire [4-1:0] node16205;
	wire [4-1:0] node16206;
	wire [4-1:0] node16207;
	wire [4-1:0] node16210;
	wire [4-1:0] node16213;
	wire [4-1:0] node16214;
	wire [4-1:0] node16217;
	wire [4-1:0] node16220;
	wire [4-1:0] node16221;
	wire [4-1:0] node16222;
	wire [4-1:0] node16223;
	wire [4-1:0] node16224;
	wire [4-1:0] node16229;
	wire [4-1:0] node16231;
	wire [4-1:0] node16234;
	wire [4-1:0] node16235;
	wire [4-1:0] node16237;
	wire [4-1:0] node16240;
	wire [4-1:0] node16241;
	wire [4-1:0] node16242;
	wire [4-1:0] node16246;
	wire [4-1:0] node16247;
	wire [4-1:0] node16251;
	wire [4-1:0] node16252;
	wire [4-1:0] node16253;
	wire [4-1:0] node16255;
	wire [4-1:0] node16258;
	wire [4-1:0] node16259;
	wire [4-1:0] node16262;
	wire [4-1:0] node16265;
	wire [4-1:0] node16266;
	wire [4-1:0] node16267;
	wire [4-1:0] node16268;
	wire [4-1:0] node16271;
	wire [4-1:0] node16274;
	wire [4-1:0] node16275;
	wire [4-1:0] node16278;
	wire [4-1:0] node16281;
	wire [4-1:0] node16282;
	wire [4-1:0] node16284;
	wire [4-1:0] node16285;
	wire [4-1:0] node16288;
	wire [4-1:0] node16291;
	wire [4-1:0] node16292;
	wire [4-1:0] node16293;
	wire [4-1:0] node16297;
	wire [4-1:0] node16299;
	wire [4-1:0] node16302;
	wire [4-1:0] node16303;
	wire [4-1:0] node16304;
	wire [4-1:0] node16305;
	wire [4-1:0] node16306;
	wire [4-1:0] node16307;
	wire [4-1:0] node16308;
	wire [4-1:0] node16310;
	wire [4-1:0] node16311;
	wire [4-1:0] node16314;
	wire [4-1:0] node16317;
	wire [4-1:0] node16320;
	wire [4-1:0] node16321;
	wire [4-1:0] node16323;
	wire [4-1:0] node16324;
	wire [4-1:0] node16327;
	wire [4-1:0] node16330;
	wire [4-1:0] node16331;
	wire [4-1:0] node16332;
	wire [4-1:0] node16335;
	wire [4-1:0] node16339;
	wire [4-1:0] node16340;
	wire [4-1:0] node16341;
	wire [4-1:0] node16342;
	wire [4-1:0] node16343;
	wire [4-1:0] node16346;
	wire [4-1:0] node16350;
	wire [4-1:0] node16351;
	wire [4-1:0] node16352;
	wire [4-1:0] node16355;
	wire [4-1:0] node16358;
	wire [4-1:0] node16359;
	wire [4-1:0] node16363;
	wire [4-1:0] node16364;
	wire [4-1:0] node16366;
	wire [4-1:0] node16369;
	wire [4-1:0] node16370;
	wire [4-1:0] node16372;
	wire [4-1:0] node16375;
	wire [4-1:0] node16377;
	wire [4-1:0] node16380;
	wire [4-1:0] node16381;
	wire [4-1:0] node16382;
	wire [4-1:0] node16383;
	wire [4-1:0] node16384;
	wire [4-1:0] node16387;
	wire [4-1:0] node16390;
	wire [4-1:0] node16391;
	wire [4-1:0] node16394;
	wire [4-1:0] node16397;
	wire [4-1:0] node16398;
	wire [4-1:0] node16399;
	wire [4-1:0] node16403;
	wire [4-1:0] node16404;
	wire [4-1:0] node16407;
	wire [4-1:0] node16410;
	wire [4-1:0] node16411;
	wire [4-1:0] node16412;
	wire [4-1:0] node16413;
	wire [4-1:0] node16416;
	wire [4-1:0] node16417;
	wire [4-1:0] node16420;
	wire [4-1:0] node16423;
	wire [4-1:0] node16424;
	wire [4-1:0] node16426;
	wire [4-1:0] node16429;
	wire [4-1:0] node16430;
	wire [4-1:0] node16433;
	wire [4-1:0] node16436;
	wire [4-1:0] node16437;
	wire [4-1:0] node16438;
	wire [4-1:0] node16439;
	wire [4-1:0] node16442;
	wire [4-1:0] node16445;
	wire [4-1:0] node16446;
	wire [4-1:0] node16450;
	wire [4-1:0] node16451;
	wire [4-1:0] node16453;
	wire [4-1:0] node16457;
	wire [4-1:0] node16458;
	wire [4-1:0] node16459;
	wire [4-1:0] node16460;
	wire [4-1:0] node16461;
	wire [4-1:0] node16463;
	wire [4-1:0] node16464;
	wire [4-1:0] node16467;
	wire [4-1:0] node16470;
	wire [4-1:0] node16471;
	wire [4-1:0] node16472;
	wire [4-1:0] node16476;
	wire [4-1:0] node16477;
	wire [4-1:0] node16481;
	wire [4-1:0] node16482;
	wire [4-1:0] node16483;
	wire [4-1:0] node16486;
	wire [4-1:0] node16487;
	wire [4-1:0] node16490;
	wire [4-1:0] node16493;
	wire [4-1:0] node16494;
	wire [4-1:0] node16495;
	wire [4-1:0] node16499;
	wire [4-1:0] node16500;
	wire [4-1:0] node16503;
	wire [4-1:0] node16506;
	wire [4-1:0] node16507;
	wire [4-1:0] node16508;
	wire [4-1:0] node16509;
	wire [4-1:0] node16511;
	wire [4-1:0] node16515;
	wire [4-1:0] node16516;
	wire [4-1:0] node16520;
	wire [4-1:0] node16521;
	wire [4-1:0] node16522;
	wire [4-1:0] node16524;
	wire [4-1:0] node16527;
	wire [4-1:0] node16529;
	wire [4-1:0] node16532;
	wire [4-1:0] node16533;
	wire [4-1:0] node16536;
	wire [4-1:0] node16539;
	wire [4-1:0] node16540;
	wire [4-1:0] node16541;
	wire [4-1:0] node16543;
	wire [4-1:0] node16545;
	wire [4-1:0] node16548;
	wire [4-1:0] node16549;
	wire [4-1:0] node16551;
	wire [4-1:0] node16554;
	wire [4-1:0] node16555;
	wire [4-1:0] node16558;
	wire [4-1:0] node16561;
	wire [4-1:0] node16562;
	wire [4-1:0] node16563;
	wire [4-1:0] node16564;
	wire [4-1:0] node16565;
	wire [4-1:0] node16568;
	wire [4-1:0] node16572;
	wire [4-1:0] node16573;
	wire [4-1:0] node16574;
	wire [4-1:0] node16577;
	wire [4-1:0] node16581;
	wire [4-1:0] node16582;
	wire [4-1:0] node16583;
	wire [4-1:0] node16587;
	wire [4-1:0] node16588;
	wire [4-1:0] node16591;
	wire [4-1:0] node16594;
	wire [4-1:0] node16595;
	wire [4-1:0] node16596;
	wire [4-1:0] node16597;
	wire [4-1:0] node16598;
	wire [4-1:0] node16599;
	wire [4-1:0] node16600;
	wire [4-1:0] node16603;
	wire [4-1:0] node16606;
	wire [4-1:0] node16607;
	wire [4-1:0] node16610;
	wire [4-1:0] node16613;
	wire [4-1:0] node16614;
	wire [4-1:0] node16617;
	wire [4-1:0] node16620;
	wire [4-1:0] node16621;
	wire [4-1:0] node16622;
	wire [4-1:0] node16625;
	wire [4-1:0] node16628;
	wire [4-1:0] node16629;
	wire [4-1:0] node16632;
	wire [4-1:0] node16635;
	wire [4-1:0] node16636;
	wire [4-1:0] node16637;
	wire [4-1:0] node16638;
	wire [4-1:0] node16641;
	wire [4-1:0] node16644;
	wire [4-1:0] node16645;
	wire [4-1:0] node16646;
	wire [4-1:0] node16650;
	wire [4-1:0] node16651;
	wire [4-1:0] node16655;
	wire [4-1:0] node16656;
	wire [4-1:0] node16659;
	wire [4-1:0] node16662;
	wire [4-1:0] node16663;
	wire [4-1:0] node16664;
	wire [4-1:0] node16665;
	wire [4-1:0] node16666;
	wire [4-1:0] node16669;
	wire [4-1:0] node16672;
	wire [4-1:0] node16673;
	wire [4-1:0] node16677;
	wire [4-1:0] node16678;
	wire [4-1:0] node16680;
	wire [4-1:0] node16681;
	wire [4-1:0] node16684;
	wire [4-1:0] node16687;
	wire [4-1:0] node16688;
	wire [4-1:0] node16690;
	wire [4-1:0] node16693;
	wire [4-1:0] node16696;
	wire [4-1:0] node16697;
	wire [4-1:0] node16698;
	wire [4-1:0] node16699;
	wire [4-1:0] node16702;
	wire [4-1:0] node16703;
	wire [4-1:0] node16707;
	wire [4-1:0] node16708;
	wire [4-1:0] node16711;
	wire [4-1:0] node16714;
	wire [4-1:0] node16715;
	wire [4-1:0] node16718;
	wire [4-1:0] node16721;
	wire [4-1:0] node16722;
	wire [4-1:0] node16723;
	wire [4-1:0] node16724;
	wire [4-1:0] node16725;
	wire [4-1:0] node16726;
	wire [4-1:0] node16727;
	wire [4-1:0] node16728;
	wire [4-1:0] node16729;
	wire [4-1:0] node16730;
	wire [4-1:0] node16733;
	wire [4-1:0] node16736;
	wire [4-1:0] node16739;
	wire [4-1:0] node16740;
	wire [4-1:0] node16741;
	wire [4-1:0] node16744;
	wire [4-1:0] node16748;
	wire [4-1:0] node16749;
	wire [4-1:0] node16750;
	wire [4-1:0] node16753;
	wire [4-1:0] node16755;
	wire [4-1:0] node16758;
	wire [4-1:0] node16759;
	wire [4-1:0] node16760;
	wire [4-1:0] node16763;
	wire [4-1:0] node16766;
	wire [4-1:0] node16767;
	wire [4-1:0] node16770;
	wire [4-1:0] node16773;
	wire [4-1:0] node16774;
	wire [4-1:0] node16775;
	wire [4-1:0] node16776;
	wire [4-1:0] node16779;
	wire [4-1:0] node16782;
	wire [4-1:0] node16784;
	wire [4-1:0] node16785;
	wire [4-1:0] node16789;
	wire [4-1:0] node16790;
	wire [4-1:0] node16791;
	wire [4-1:0] node16794;
	wire [4-1:0] node16797;
	wire [4-1:0] node16798;
	wire [4-1:0] node16800;
	wire [4-1:0] node16803;
	wire [4-1:0] node16804;
	wire [4-1:0] node16808;
	wire [4-1:0] node16809;
	wire [4-1:0] node16810;
	wire [4-1:0] node16811;
	wire [4-1:0] node16812;
	wire [4-1:0] node16815;
	wire [4-1:0] node16818;
	wire [4-1:0] node16819;
	wire [4-1:0] node16820;
	wire [4-1:0] node16823;
	wire [4-1:0] node16826;
	wire [4-1:0] node16827;
	wire [4-1:0] node16830;
	wire [4-1:0] node16833;
	wire [4-1:0] node16834;
	wire [4-1:0] node16835;
	wire [4-1:0] node16837;
	wire [4-1:0] node16840;
	wire [4-1:0] node16841;
	wire [4-1:0] node16844;
	wire [4-1:0] node16847;
	wire [4-1:0] node16848;
	wire [4-1:0] node16850;
	wire [4-1:0] node16853;
	wire [4-1:0] node16854;
	wire [4-1:0] node16855;
	wire [4-1:0] node16858;
	wire [4-1:0] node16861;
	wire [4-1:0] node16863;
	wire [4-1:0] node16866;
	wire [4-1:0] node16867;
	wire [4-1:0] node16868;
	wire [4-1:0] node16869;
	wire [4-1:0] node16870;
	wire [4-1:0] node16873;
	wire [4-1:0] node16876;
	wire [4-1:0] node16877;
	wire [4-1:0] node16878;
	wire [4-1:0] node16882;
	wire [4-1:0] node16883;
	wire [4-1:0] node16887;
	wire [4-1:0] node16889;
	wire [4-1:0] node16890;
	wire [4-1:0] node16893;
	wire [4-1:0] node16896;
	wire [4-1:0] node16897;
	wire [4-1:0] node16898;
	wire [4-1:0] node16899;
	wire [4-1:0] node16903;
	wire [4-1:0] node16904;
	wire [4-1:0] node16907;
	wire [4-1:0] node16910;
	wire [4-1:0] node16911;
	wire [4-1:0] node16912;
	wire [4-1:0] node16913;
	wire [4-1:0] node16918;
	wire [4-1:0] node16919;
	wire [4-1:0] node16920;
	wire [4-1:0] node16924;
	wire [4-1:0] node16925;
	wire [4-1:0] node16929;
	wire [4-1:0] node16930;
	wire [4-1:0] node16931;
	wire [4-1:0] node16932;
	wire [4-1:0] node16933;
	wire [4-1:0] node16934;
	wire [4-1:0] node16935;
	wire [4-1:0] node16939;
	wire [4-1:0] node16940;
	wire [4-1:0] node16943;
	wire [4-1:0] node16946;
	wire [4-1:0] node16947;
	wire [4-1:0] node16948;
	wire [4-1:0] node16949;
	wire [4-1:0] node16953;
	wire [4-1:0] node16954;
	wire [4-1:0] node16958;
	wire [4-1:0] node16959;
	wire [4-1:0] node16960;
	wire [4-1:0] node16963;
	wire [4-1:0] node16966;
	wire [4-1:0] node16967;
	wire [4-1:0] node16971;
	wire [4-1:0] node16972;
	wire [4-1:0] node16973;
	wire [4-1:0] node16974;
	wire [4-1:0] node16977;
	wire [4-1:0] node16980;
	wire [4-1:0] node16982;
	wire [4-1:0] node16985;
	wire [4-1:0] node16986;
	wire [4-1:0] node16987;
	wire [4-1:0] node16990;
	wire [4-1:0] node16993;
	wire [4-1:0] node16994;
	wire [4-1:0] node16995;
	wire [4-1:0] node16998;
	wire [4-1:0] node17001;
	wire [4-1:0] node17002;
	wire [4-1:0] node17005;
	wire [4-1:0] node17008;
	wire [4-1:0] node17009;
	wire [4-1:0] node17010;
	wire [4-1:0] node17011;
	wire [4-1:0] node17014;
	wire [4-1:0] node17017;
	wire [4-1:0] node17018;
	wire [4-1:0] node17021;
	wire [4-1:0] node17024;
	wire [4-1:0] node17025;
	wire [4-1:0] node17026;
	wire [4-1:0] node17028;
	wire [4-1:0] node17032;
	wire [4-1:0] node17033;
	wire [4-1:0] node17036;
	wire [4-1:0] node17039;
	wire [4-1:0] node17040;
	wire [4-1:0] node17041;
	wire [4-1:0] node17042;
	wire [4-1:0] node17043;
	wire [4-1:0] node17046;
	wire [4-1:0] node17049;
	wire [4-1:0] node17050;
	wire [4-1:0] node17053;
	wire [4-1:0] node17056;
	wire [4-1:0] node17057;
	wire [4-1:0] node17058;
	wire [4-1:0] node17061;
	wire [4-1:0] node17064;
	wire [4-1:0] node17065;
	wire [4-1:0] node17068;
	wire [4-1:0] node17071;
	wire [4-1:0] node17072;
	wire [4-1:0] node17073;
	wire [4-1:0] node17074;
	wire [4-1:0] node17077;
	wire [4-1:0] node17080;
	wire [4-1:0] node17081;
	wire [4-1:0] node17084;
	wire [4-1:0] node17087;
	wire [4-1:0] node17088;
	wire [4-1:0] node17089;
	wire [4-1:0] node17092;
	wire [4-1:0] node17095;
	wire [4-1:0] node17096;
	wire [4-1:0] node17099;
	wire [4-1:0] node17102;
	wire [4-1:0] node17103;
	wire [4-1:0] node17104;
	wire [4-1:0] node17105;
	wire [4-1:0] node17106;
	wire [4-1:0] node17107;
	wire [4-1:0] node17108;
	wire [4-1:0] node17111;
	wire [4-1:0] node17113;
	wire [4-1:0] node17116;
	wire [4-1:0] node17117;
	wire [4-1:0] node17118;
	wire [4-1:0] node17121;
	wire [4-1:0] node17124;
	wire [4-1:0] node17126;
	wire [4-1:0] node17129;
	wire [4-1:0] node17130;
	wire [4-1:0] node17131;
	wire [4-1:0] node17134;
	wire [4-1:0] node17136;
	wire [4-1:0] node17139;
	wire [4-1:0] node17140;
	wire [4-1:0] node17141;
	wire [4-1:0] node17144;
	wire [4-1:0] node17147;
	wire [4-1:0] node17149;
	wire [4-1:0] node17150;
	wire [4-1:0] node17153;
	wire [4-1:0] node17156;
	wire [4-1:0] node17157;
	wire [4-1:0] node17158;
	wire [4-1:0] node17159;
	wire [4-1:0] node17160;
	wire [4-1:0] node17163;
	wire [4-1:0] node17166;
	wire [4-1:0] node17168;
	wire [4-1:0] node17170;
	wire [4-1:0] node17173;
	wire [4-1:0] node17174;
	wire [4-1:0] node17175;
	wire [4-1:0] node17178;
	wire [4-1:0] node17181;
	wire [4-1:0] node17182;
	wire [4-1:0] node17183;
	wire [4-1:0] node17187;
	wire [4-1:0] node17188;
	wire [4-1:0] node17191;
	wire [4-1:0] node17194;
	wire [4-1:0] node17195;
	wire [4-1:0] node17196;
	wire [4-1:0] node17199;
	wire [4-1:0] node17201;
	wire [4-1:0] node17204;
	wire [4-1:0] node17205;
	wire [4-1:0] node17206;
	wire [4-1:0] node17209;
	wire [4-1:0] node17212;
	wire [4-1:0] node17213;
	wire [4-1:0] node17217;
	wire [4-1:0] node17218;
	wire [4-1:0] node17219;
	wire [4-1:0] node17220;
	wire [4-1:0] node17221;
	wire [4-1:0] node17223;
	wire [4-1:0] node17224;
	wire [4-1:0] node17228;
	wire [4-1:0] node17229;
	wire [4-1:0] node17230;
	wire [4-1:0] node17233;
	wire [4-1:0] node17237;
	wire [4-1:0] node17238;
	wire [4-1:0] node17239;
	wire [4-1:0] node17240;
	wire [4-1:0] node17243;
	wire [4-1:0] node17246;
	wire [4-1:0] node17247;
	wire [4-1:0] node17251;
	wire [4-1:0] node17252;
	wire [4-1:0] node17256;
	wire [4-1:0] node17257;
	wire [4-1:0] node17258;
	wire [4-1:0] node17259;
	wire [4-1:0] node17260;
	wire [4-1:0] node17263;
	wire [4-1:0] node17266;
	wire [4-1:0] node17267;
	wire [4-1:0] node17270;
	wire [4-1:0] node17273;
	wire [4-1:0] node17275;
	wire [4-1:0] node17276;
	wire [4-1:0] node17280;
	wire [4-1:0] node17281;
	wire [4-1:0] node17282;
	wire [4-1:0] node17283;
	wire [4-1:0] node17286;
	wire [4-1:0] node17290;
	wire [4-1:0] node17292;
	wire [4-1:0] node17293;
	wire [4-1:0] node17297;
	wire [4-1:0] node17298;
	wire [4-1:0] node17299;
	wire [4-1:0] node17300;
	wire [4-1:0] node17303;
	wire [4-1:0] node17304;
	wire [4-1:0] node17306;
	wire [4-1:0] node17310;
	wire [4-1:0] node17311;
	wire [4-1:0] node17312;
	wire [4-1:0] node17313;
	wire [4-1:0] node17316;
	wire [4-1:0] node17320;
	wire [4-1:0] node17322;
	wire [4-1:0] node17324;
	wire [4-1:0] node17327;
	wire [4-1:0] node17328;
	wire [4-1:0] node17330;
	wire [4-1:0] node17332;
	wire [4-1:0] node17334;
	wire [4-1:0] node17337;
	wire [4-1:0] node17338;
	wire [4-1:0] node17339;
	wire [4-1:0] node17342;
	wire [4-1:0] node17345;
	wire [4-1:0] node17346;
	wire [4-1:0] node17349;
	wire [4-1:0] node17352;
	wire [4-1:0] node17353;
	wire [4-1:0] node17354;
	wire [4-1:0] node17355;
	wire [4-1:0] node17356;
	wire [4-1:0] node17357;
	wire [4-1:0] node17358;
	wire [4-1:0] node17360;
	wire [4-1:0] node17363;
	wire [4-1:0] node17364;
	wire [4-1:0] node17368;
	wire [4-1:0] node17370;
	wire [4-1:0] node17371;
	wire [4-1:0] node17374;
	wire [4-1:0] node17377;
	wire [4-1:0] node17378;
	wire [4-1:0] node17379;
	wire [4-1:0] node17380;
	wire [4-1:0] node17383;
	wire [4-1:0] node17387;
	wire [4-1:0] node17389;
	wire [4-1:0] node17390;
	wire [4-1:0] node17393;
	wire [4-1:0] node17396;
	wire [4-1:0] node17397;
	wire [4-1:0] node17398;
	wire [4-1:0] node17399;
	wire [4-1:0] node17401;
	wire [4-1:0] node17404;
	wire [4-1:0] node17405;
	wire [4-1:0] node17409;
	wire [4-1:0] node17410;
	wire [4-1:0] node17413;
	wire [4-1:0] node17414;
	wire [4-1:0] node17417;
	wire [4-1:0] node17420;
	wire [4-1:0] node17421;
	wire [4-1:0] node17422;
	wire [4-1:0] node17426;
	wire [4-1:0] node17428;
	wire [4-1:0] node17430;
	wire [4-1:0] node17433;
	wire [4-1:0] node17434;
	wire [4-1:0] node17435;
	wire [4-1:0] node17436;
	wire [4-1:0] node17437;
	wire [4-1:0] node17438;
	wire [4-1:0] node17441;
	wire [4-1:0] node17445;
	wire [4-1:0] node17447;
	wire [4-1:0] node17448;
	wire [4-1:0] node17451;
	wire [4-1:0] node17454;
	wire [4-1:0] node17455;
	wire [4-1:0] node17457;
	wire [4-1:0] node17458;
	wire [4-1:0] node17461;
	wire [4-1:0] node17464;
	wire [4-1:0] node17465;
	wire [4-1:0] node17468;
	wire [4-1:0] node17469;
	wire [4-1:0] node17472;
	wire [4-1:0] node17475;
	wire [4-1:0] node17476;
	wire [4-1:0] node17477;
	wire [4-1:0] node17478;
	wire [4-1:0] node17479;
	wire [4-1:0] node17484;
	wire [4-1:0] node17486;
	wire [4-1:0] node17487;
	wire [4-1:0] node17490;
	wire [4-1:0] node17493;
	wire [4-1:0] node17494;
	wire [4-1:0] node17495;
	wire [4-1:0] node17499;
	wire [4-1:0] node17502;
	wire [4-1:0] node17503;
	wire [4-1:0] node17504;
	wire [4-1:0] node17505;
	wire [4-1:0] node17506;
	wire [4-1:0] node17507;
	wire [4-1:0] node17508;
	wire [4-1:0] node17511;
	wire [4-1:0] node17514;
	wire [4-1:0] node17516;
	wire [4-1:0] node17519;
	wire [4-1:0] node17521;
	wire [4-1:0] node17524;
	wire [4-1:0] node17525;
	wire [4-1:0] node17526;
	wire [4-1:0] node17527;
	wire [4-1:0] node17531;
	wire [4-1:0] node17534;
	wire [4-1:0] node17535;
	wire [4-1:0] node17538;
	wire [4-1:0] node17539;
	wire [4-1:0] node17542;
	wire [4-1:0] node17545;
	wire [4-1:0] node17546;
	wire [4-1:0] node17547;
	wire [4-1:0] node17548;
	wire [4-1:0] node17551;
	wire [4-1:0] node17554;
	wire [4-1:0] node17555;
	wire [4-1:0] node17558;
	wire [4-1:0] node17561;
	wire [4-1:0] node17562;
	wire [4-1:0] node17564;
	wire [4-1:0] node17566;
	wire [4-1:0] node17569;
	wire [4-1:0] node17570;
	wire [4-1:0] node17572;
	wire [4-1:0] node17575;
	wire [4-1:0] node17578;
	wire [4-1:0] node17579;
	wire [4-1:0] node17580;
	wire [4-1:0] node17581;
	wire [4-1:0] node17582;
	wire [4-1:0] node17585;
	wire [4-1:0] node17588;
	wire [4-1:0] node17589;
	wire [4-1:0] node17592;
	wire [4-1:0] node17593;
	wire [4-1:0] node17597;
	wire [4-1:0] node17598;
	wire [4-1:0] node17599;
	wire [4-1:0] node17600;
	wire [4-1:0] node17603;
	wire [4-1:0] node17607;
	wire [4-1:0] node17609;
	wire [4-1:0] node17612;
	wire [4-1:0] node17613;
	wire [4-1:0] node17614;
	wire [4-1:0] node17615;
	wire [4-1:0] node17618;
	wire [4-1:0] node17619;
	wire [4-1:0] node17623;
	wire [4-1:0] node17624;
	wire [4-1:0] node17627;
	wire [4-1:0] node17630;
	wire [4-1:0] node17631;
	wire [4-1:0] node17632;
	wire [4-1:0] node17635;
	wire [4-1:0] node17638;
	wire [4-1:0] node17641;
	wire [4-1:0] node17642;
	wire [4-1:0] node17643;
	wire [4-1:0] node17644;
	wire [4-1:0] node17645;
	wire [4-1:0] node17646;
	wire [4-1:0] node17647;
	wire [4-1:0] node17649;
	wire [4-1:0] node17650;
	wire [4-1:0] node17653;
	wire [4-1:0] node17656;
	wire [4-1:0] node17657;
	wire [4-1:0] node17658;
	wire [4-1:0] node17662;
	wire [4-1:0] node17664;
	wire [4-1:0] node17667;
	wire [4-1:0] node17668;
	wire [4-1:0] node17669;
	wire [4-1:0] node17670;
	wire [4-1:0] node17674;
	wire [4-1:0] node17675;
	wire [4-1:0] node17679;
	wire [4-1:0] node17680;
	wire [4-1:0] node17681;
	wire [4-1:0] node17684;
	wire [4-1:0] node17687;
	wire [4-1:0] node17689;
	wire [4-1:0] node17690;
	wire [4-1:0] node17694;
	wire [4-1:0] node17695;
	wire [4-1:0] node17696;
	wire [4-1:0] node17697;
	wire [4-1:0] node17698;
	wire [4-1:0] node17701;
	wire [4-1:0] node17702;
	wire [4-1:0] node17705;
	wire [4-1:0] node17708;
	wire [4-1:0] node17709;
	wire [4-1:0] node17713;
	wire [4-1:0] node17714;
	wire [4-1:0] node17717;
	wire [4-1:0] node17719;
	wire [4-1:0] node17720;
	wire [4-1:0] node17724;
	wire [4-1:0] node17725;
	wire [4-1:0] node17726;
	wire [4-1:0] node17727;
	wire [4-1:0] node17730;
	wire [4-1:0] node17733;
	wire [4-1:0] node17734;
	wire [4-1:0] node17738;
	wire [4-1:0] node17739;
	wire [4-1:0] node17740;
	wire [4-1:0] node17741;
	wire [4-1:0] node17746;
	wire [4-1:0] node17747;
	wire [4-1:0] node17750;
	wire [4-1:0] node17753;
	wire [4-1:0] node17754;
	wire [4-1:0] node17755;
	wire [4-1:0] node17756;
	wire [4-1:0] node17757;
	wire [4-1:0] node17758;
	wire [4-1:0] node17759;
	wire [4-1:0] node17763;
	wire [4-1:0] node17764;
	wire [4-1:0] node17768;
	wire [4-1:0] node17769;
	wire [4-1:0] node17770;
	wire [4-1:0] node17774;
	wire [4-1:0] node17775;
	wire [4-1:0] node17778;
	wire [4-1:0] node17781;
	wire [4-1:0] node17782;
	wire [4-1:0] node17784;
	wire [4-1:0] node17785;
	wire [4-1:0] node17789;
	wire [4-1:0] node17791;
	wire [4-1:0] node17792;
	wire [4-1:0] node17796;
	wire [4-1:0] node17797;
	wire [4-1:0] node17798;
	wire [4-1:0] node17799;
	wire [4-1:0] node17800;
	wire [4-1:0] node17804;
	wire [4-1:0] node17806;
	wire [4-1:0] node17809;
	wire [4-1:0] node17810;
	wire [4-1:0] node17814;
	wire [4-1:0] node17815;
	wire [4-1:0] node17817;
	wire [4-1:0] node17818;
	wire [4-1:0] node17821;
	wire [4-1:0] node17824;
	wire [4-1:0] node17825;
	wire [4-1:0] node17826;
	wire [4-1:0] node17830;
	wire [4-1:0] node17831;
	wire [4-1:0] node17835;
	wire [4-1:0] node17836;
	wire [4-1:0] node17837;
	wire [4-1:0] node17838;
	wire [4-1:0] node17841;
	wire [4-1:0] node17844;
	wire [4-1:0] node17846;
	wire [4-1:0] node17847;
	wire [4-1:0] node17851;
	wire [4-1:0] node17852;
	wire [4-1:0] node17853;
	wire [4-1:0] node17854;
	wire [4-1:0] node17857;
	wire [4-1:0] node17858;
	wire [4-1:0] node17861;
	wire [4-1:0] node17864;
	wire [4-1:0] node17865;
	wire [4-1:0] node17868;
	wire [4-1:0] node17871;
	wire [4-1:0] node17872;
	wire [4-1:0] node17873;
	wire [4-1:0] node17875;
	wire [4-1:0] node17879;
	wire [4-1:0] node17881;
	wire [4-1:0] node17884;
	wire [4-1:0] node17885;
	wire [4-1:0] node17886;
	wire [4-1:0] node17887;
	wire [4-1:0] node17888;
	wire [4-1:0] node17889;
	wire [4-1:0] node17892;
	wire [4-1:0] node17895;
	wire [4-1:0] node17896;
	wire [4-1:0] node17897;
	wire [4-1:0] node17900;
	wire [4-1:0] node17903;
	wire [4-1:0] node17904;
	wire [4-1:0] node17907;
	wire [4-1:0] node17910;
	wire [4-1:0] node17911;
	wire [4-1:0] node17913;
	wire [4-1:0] node17916;
	wire [4-1:0] node17917;
	wire [4-1:0] node17918;
	wire [4-1:0] node17921;
	wire [4-1:0] node17925;
	wire [4-1:0] node17926;
	wire [4-1:0] node17927;
	wire [4-1:0] node17928;
	wire [4-1:0] node17929;
	wire [4-1:0] node17933;
	wire [4-1:0] node17934;
	wire [4-1:0] node17937;
	wire [4-1:0] node17940;
	wire [4-1:0] node17941;
	wire [4-1:0] node17942;
	wire [4-1:0] node17943;
	wire [4-1:0] node17947;
	wire [4-1:0] node17949;
	wire [4-1:0] node17952;
	wire [4-1:0] node17954;
	wire [4-1:0] node17955;
	wire [4-1:0] node17959;
	wire [4-1:0] node17960;
	wire [4-1:0] node17961;
	wire [4-1:0] node17962;
	wire [4-1:0] node17965;
	wire [4-1:0] node17968;
	wire [4-1:0] node17969;
	wire [4-1:0] node17971;
	wire [4-1:0] node17975;
	wire [4-1:0] node17976;
	wire [4-1:0] node17977;
	wire [4-1:0] node17980;
	wire [4-1:0] node17983;
	wire [4-1:0] node17984;
	wire [4-1:0] node17987;
	wire [4-1:0] node17990;
	wire [4-1:0] node17991;
	wire [4-1:0] node17992;
	wire [4-1:0] node17993;
	wire [4-1:0] node17994;
	wire [4-1:0] node17996;
	wire [4-1:0] node17999;
	wire [4-1:0] node18000;
	wire [4-1:0] node18003;
	wire [4-1:0] node18006;
	wire [4-1:0] node18007;
	wire [4-1:0] node18008;
	wire [4-1:0] node18012;
	wire [4-1:0] node18015;
	wire [4-1:0] node18016;
	wire [4-1:0] node18017;
	wire [4-1:0] node18018;
	wire [4-1:0] node18022;
	wire [4-1:0] node18023;
	wire [4-1:0] node18026;
	wire [4-1:0] node18029;
	wire [4-1:0] node18031;
	wire [4-1:0] node18032;
	wire [4-1:0] node18033;
	wire [4-1:0] node18036;
	wire [4-1:0] node18039;
	wire [4-1:0] node18041;
	wire [4-1:0] node18044;
	wire [4-1:0] node18045;
	wire [4-1:0] node18046;
	wire [4-1:0] node18047;
	wire [4-1:0] node18049;
	wire [4-1:0] node18052;
	wire [4-1:0] node18053;
	wire [4-1:0] node18057;
	wire [4-1:0] node18060;
	wire [4-1:0] node18061;
	wire [4-1:0] node18062;
	wire [4-1:0] node18064;
	wire [4-1:0] node18065;
	wire [4-1:0] node18068;
	wire [4-1:0] node18071;
	wire [4-1:0] node18072;
	wire [4-1:0] node18075;
	wire [4-1:0] node18078;
	wire [4-1:0] node18079;
	wire [4-1:0] node18080;
	wire [4-1:0] node18083;
	wire [4-1:0] node18086;
	wire [4-1:0] node18087;
	wire [4-1:0] node18090;
	wire [4-1:0] node18093;
	wire [4-1:0] node18094;
	wire [4-1:0] node18095;
	wire [4-1:0] node18096;
	wire [4-1:0] node18097;
	wire [4-1:0] node18098;
	wire [4-1:0] node18099;
	wire [4-1:0] node18100;
	wire [4-1:0] node18103;
	wire [4-1:0] node18106;
	wire [4-1:0] node18109;
	wire [4-1:0] node18110;
	wire [4-1:0] node18111;
	wire [4-1:0] node18112;
	wire [4-1:0] node18117;
	wire [4-1:0] node18118;
	wire [4-1:0] node18119;
	wire [4-1:0] node18122;
	wire [4-1:0] node18125;
	wire [4-1:0] node18128;
	wire [4-1:0] node18129;
	wire [4-1:0] node18130;
	wire [4-1:0] node18132;
	wire [4-1:0] node18135;
	wire [4-1:0] node18136;
	wire [4-1:0] node18139;
	wire [4-1:0] node18140;
	wire [4-1:0] node18144;
	wire [4-1:0] node18145;
	wire [4-1:0] node18146;
	wire [4-1:0] node18148;
	wire [4-1:0] node18152;
	wire [4-1:0] node18154;
	wire [4-1:0] node18155;
	wire [4-1:0] node18159;
	wire [4-1:0] node18160;
	wire [4-1:0] node18161;
	wire [4-1:0] node18162;
	wire [4-1:0] node18163;
	wire [4-1:0] node18164;
	wire [4-1:0] node18169;
	wire [4-1:0] node18170;
	wire [4-1:0] node18172;
	wire [4-1:0] node18175;
	wire [4-1:0] node18177;
	wire [4-1:0] node18180;
	wire [4-1:0] node18181;
	wire [4-1:0] node18182;
	wire [4-1:0] node18184;
	wire [4-1:0] node18188;
	wire [4-1:0] node18190;
	wire [4-1:0] node18193;
	wire [4-1:0] node18194;
	wire [4-1:0] node18195;
	wire [4-1:0] node18196;
	wire [4-1:0] node18197;
	wire [4-1:0] node18200;
	wire [4-1:0] node18204;
	wire [4-1:0] node18206;
	wire [4-1:0] node18209;
	wire [4-1:0] node18210;
	wire [4-1:0] node18212;
	wire [4-1:0] node18213;
	wire [4-1:0] node18216;
	wire [4-1:0] node18219;
	wire [4-1:0] node18220;
	wire [4-1:0] node18221;
	wire [4-1:0] node18224;
	wire [4-1:0] node18227;
	wire [4-1:0] node18228;
	wire [4-1:0] node18231;
	wire [4-1:0] node18234;
	wire [4-1:0] node18235;
	wire [4-1:0] node18236;
	wire [4-1:0] node18237;
	wire [4-1:0] node18239;
	wire [4-1:0] node18240;
	wire [4-1:0] node18241;
	wire [4-1:0] node18244;
	wire [4-1:0] node18248;
	wire [4-1:0] node18249;
	wire [4-1:0] node18250;
	wire [4-1:0] node18251;
	wire [4-1:0] node18256;
	wire [4-1:0] node18257;
	wire [4-1:0] node18261;
	wire [4-1:0] node18262;
	wire [4-1:0] node18263;
	wire [4-1:0] node18264;
	wire [4-1:0] node18265;
	wire [4-1:0] node18269;
	wire [4-1:0] node18270;
	wire [4-1:0] node18274;
	wire [4-1:0] node18275;
	wire [4-1:0] node18278;
	wire [4-1:0] node18279;
	wire [4-1:0] node18282;
	wire [4-1:0] node18285;
	wire [4-1:0] node18286;
	wire [4-1:0] node18287;
	wire [4-1:0] node18288;
	wire [4-1:0] node18291;
	wire [4-1:0] node18295;
	wire [4-1:0] node18296;
	wire [4-1:0] node18297;
	wire [4-1:0] node18300;
	wire [4-1:0] node18304;
	wire [4-1:0] node18305;
	wire [4-1:0] node18306;
	wire [4-1:0] node18307;
	wire [4-1:0] node18308;
	wire [4-1:0] node18311;
	wire [4-1:0] node18312;
	wire [4-1:0] node18315;
	wire [4-1:0] node18318;
	wire [4-1:0] node18319;
	wire [4-1:0] node18321;
	wire [4-1:0] node18324;
	wire [4-1:0] node18325;
	wire [4-1:0] node18328;
	wire [4-1:0] node18331;
	wire [4-1:0] node18332;
	wire [4-1:0] node18333;
	wire [4-1:0] node18334;
	wire [4-1:0] node18337;
	wire [4-1:0] node18340;
	wire [4-1:0] node18343;
	wire [4-1:0] node18344;
	wire [4-1:0] node18347;
	wire [4-1:0] node18350;
	wire [4-1:0] node18351;
	wire [4-1:0] node18352;
	wire [4-1:0] node18354;
	wire [4-1:0] node18357;
	wire [4-1:0] node18358;
	wire [4-1:0] node18359;
	wire [4-1:0] node18362;
	wire [4-1:0] node18366;
	wire [4-1:0] node18367;
	wire [4-1:0] node18369;
	wire [4-1:0] node18372;
	wire [4-1:0] node18373;
	wire [4-1:0] node18374;
	wire [4-1:0] node18379;
	wire [4-1:0] node18380;
	wire [4-1:0] node18381;
	wire [4-1:0] node18382;
	wire [4-1:0] node18383;
	wire [4-1:0] node18384;
	wire [4-1:0] node18385;
	wire [4-1:0] node18386;
	wire [4-1:0] node18390;
	wire [4-1:0] node18393;
	wire [4-1:0] node18394;
	wire [4-1:0] node18395;
	wire [4-1:0] node18398;
	wire [4-1:0] node18401;
	wire [4-1:0] node18403;
	wire [4-1:0] node18406;
	wire [4-1:0] node18407;
	wire [4-1:0] node18408;
	wire [4-1:0] node18410;
	wire [4-1:0] node18414;
	wire [4-1:0] node18416;
	wire [4-1:0] node18417;
	wire [4-1:0] node18420;
	wire [4-1:0] node18423;
	wire [4-1:0] node18424;
	wire [4-1:0] node18425;
	wire [4-1:0] node18426;
	wire [4-1:0] node18427;
	wire [4-1:0] node18432;
	wire [4-1:0] node18433;
	wire [4-1:0] node18434;
	wire [4-1:0] node18437;
	wire [4-1:0] node18440;
	wire [4-1:0] node18441;
	wire [4-1:0] node18445;
	wire [4-1:0] node18446;
	wire [4-1:0] node18447;
	wire [4-1:0] node18448;
	wire [4-1:0] node18453;
	wire [4-1:0] node18454;
	wire [4-1:0] node18455;
	wire [4-1:0] node18458;
	wire [4-1:0] node18461;
	wire [4-1:0] node18462;
	wire [4-1:0] node18465;
	wire [4-1:0] node18468;
	wire [4-1:0] node18469;
	wire [4-1:0] node18470;
	wire [4-1:0] node18471;
	wire [4-1:0] node18472;
	wire [4-1:0] node18475;
	wire [4-1:0] node18478;
	wire [4-1:0] node18479;
	wire [4-1:0] node18482;
	wire [4-1:0] node18485;
	wire [4-1:0] node18486;
	wire [4-1:0] node18487;
	wire [4-1:0] node18490;
	wire [4-1:0] node18494;
	wire [4-1:0] node18495;
	wire [4-1:0] node18496;
	wire [4-1:0] node18497;
	wire [4-1:0] node18500;
	wire [4-1:0] node18503;
	wire [4-1:0] node18504;
	wire [4-1:0] node18507;
	wire [4-1:0] node18510;
	wire [4-1:0] node18511;
	wire [4-1:0] node18512;
	wire [4-1:0] node18514;
	wire [4-1:0] node18518;
	wire [4-1:0] node18519;
	wire [4-1:0] node18522;
	wire [4-1:0] node18525;
	wire [4-1:0] node18526;
	wire [4-1:0] node18527;
	wire [4-1:0] node18528;
	wire [4-1:0] node18529;
	wire [4-1:0] node18530;
	wire [4-1:0] node18531;
	wire [4-1:0] node18535;
	wire [4-1:0] node18538;
	wire [4-1:0] node18539;
	wire [4-1:0] node18543;
	wire [4-1:0] node18544;
	wire [4-1:0] node18546;
	wire [4-1:0] node18547;
	wire [4-1:0] node18550;
	wire [4-1:0] node18553;
	wire [4-1:0] node18554;
	wire [4-1:0] node18555;
	wire [4-1:0] node18558;
	wire [4-1:0] node18562;
	wire [4-1:0] node18563;
	wire [4-1:0] node18564;
	wire [4-1:0] node18566;
	wire [4-1:0] node18567;
	wire [4-1:0] node18571;
	wire [4-1:0] node18572;
	wire [4-1:0] node18575;
	wire [4-1:0] node18576;
	wire [4-1:0] node18580;
	wire [4-1:0] node18581;
	wire [4-1:0] node18582;
	wire [4-1:0] node18583;
	wire [4-1:0] node18587;
	wire [4-1:0] node18588;
	wire [4-1:0] node18591;
	wire [4-1:0] node18594;
	wire [4-1:0] node18595;
	wire [4-1:0] node18596;
	wire [4-1:0] node18601;
	wire [4-1:0] node18602;
	wire [4-1:0] node18603;
	wire [4-1:0] node18604;
	wire [4-1:0] node18605;
	wire [4-1:0] node18606;
	wire [4-1:0] node18609;
	wire [4-1:0] node18613;
	wire [4-1:0] node18614;
	wire [4-1:0] node18617;
	wire [4-1:0] node18620;
	wire [4-1:0] node18621;
	wire [4-1:0] node18622;
	wire [4-1:0] node18623;
	wire [4-1:0] node18626;
	wire [4-1:0] node18629;
	wire [4-1:0] node18632;
	wire [4-1:0] node18633;
	wire [4-1:0] node18635;
	wire [4-1:0] node18639;
	wire [4-1:0] node18640;
	wire [4-1:0] node18641;
	wire [4-1:0] node18644;
	wire [4-1:0] node18645;
	wire [4-1:0] node18647;
	wire [4-1:0] node18651;
	wire [4-1:0] node18652;
	wire [4-1:0] node18653;
	wire [4-1:0] node18655;
	wire [4-1:0] node18658;
	wire [4-1:0] node18659;
	wire [4-1:0] node18662;
	wire [4-1:0] node18665;
	wire [4-1:0] node18668;
	wire [4-1:0] node18669;
	wire [4-1:0] node18670;
	wire [4-1:0] node18671;
	wire [4-1:0] node18672;
	wire [4-1:0] node18673;
	wire [4-1:0] node18674;
	wire [4-1:0] node18675;
	wire [4-1:0] node18676;
	wire [4-1:0] node18677;
	wire [4-1:0] node18680;
	wire [4-1:0] node18682;
	wire [4-1:0] node18685;
	wire [4-1:0] node18686;
	wire [4-1:0] node18688;
	wire [4-1:0] node18691;
	wire [4-1:0] node18693;
	wire [4-1:0] node18694;
	wire [4-1:0] node18697;
	wire [4-1:0] node18700;
	wire [4-1:0] node18701;
	wire [4-1:0] node18702;
	wire [4-1:0] node18705;
	wire [4-1:0] node18707;
	wire [4-1:0] node18710;
	wire [4-1:0] node18711;
	wire [4-1:0] node18712;
	wire [4-1:0] node18716;
	wire [4-1:0] node18717;
	wire [4-1:0] node18720;
	wire [4-1:0] node18723;
	wire [4-1:0] node18724;
	wire [4-1:0] node18725;
	wire [4-1:0] node18726;
	wire [4-1:0] node18729;
	wire [4-1:0] node18732;
	wire [4-1:0] node18733;
	wire [4-1:0] node18735;
	wire [4-1:0] node18736;
	wire [4-1:0] node18739;
	wire [4-1:0] node18742;
	wire [4-1:0] node18743;
	wire [4-1:0] node18746;
	wire [4-1:0] node18749;
	wire [4-1:0] node18750;
	wire [4-1:0] node18751;
	wire [4-1:0] node18754;
	wire [4-1:0] node18757;
	wire [4-1:0] node18758;
	wire [4-1:0] node18759;
	wire [4-1:0] node18762;
	wire [4-1:0] node18765;
	wire [4-1:0] node18767;
	wire [4-1:0] node18768;
	wire [4-1:0] node18771;
	wire [4-1:0] node18774;
	wire [4-1:0] node18775;
	wire [4-1:0] node18776;
	wire [4-1:0] node18777;
	wire [4-1:0] node18778;
	wire [4-1:0] node18781;
	wire [4-1:0] node18784;
	wire [4-1:0] node18785;
	wire [4-1:0] node18786;
	wire [4-1:0] node18788;
	wire [4-1:0] node18792;
	wire [4-1:0] node18793;
	wire [4-1:0] node18796;
	wire [4-1:0] node18799;
	wire [4-1:0] node18800;
	wire [4-1:0] node18801;
	wire [4-1:0] node18804;
	wire [4-1:0] node18807;
	wire [4-1:0] node18808;
	wire [4-1:0] node18809;
	wire [4-1:0] node18812;
	wire [4-1:0] node18815;
	wire [4-1:0] node18816;
	wire [4-1:0] node18819;
	wire [4-1:0] node18822;
	wire [4-1:0] node18823;
	wire [4-1:0] node18824;
	wire [4-1:0] node18825;
	wire [4-1:0] node18826;
	wire [4-1:0] node18828;
	wire [4-1:0] node18832;
	wire [4-1:0] node18834;
	wire [4-1:0] node18837;
	wire [4-1:0] node18838;
	wire [4-1:0] node18840;
	wire [4-1:0] node18843;
	wire [4-1:0] node18844;
	wire [4-1:0] node18845;
	wire [4-1:0] node18848;
	wire [4-1:0] node18852;
	wire [4-1:0] node18853;
	wire [4-1:0] node18854;
	wire [4-1:0] node18855;
	wire [4-1:0] node18857;
	wire [4-1:0] node18860;
	wire [4-1:0] node18861;
	wire [4-1:0] node18865;
	wire [4-1:0] node18868;
	wire [4-1:0] node18869;
	wire [4-1:0] node18870;
	wire [4-1:0] node18871;
	wire [4-1:0] node18875;
	wire [4-1:0] node18876;
	wire [4-1:0] node18880;
	wire [4-1:0] node18881;
	wire [4-1:0] node18883;
	wire [4-1:0] node18886;
	wire [4-1:0] node18889;
	wire [4-1:0] node18890;
	wire [4-1:0] node18891;
	wire [4-1:0] node18892;
	wire [4-1:0] node18893;
	wire [4-1:0] node18894;
	wire [4-1:0] node18895;
	wire [4-1:0] node18897;
	wire [4-1:0] node18900;
	wire [4-1:0] node18901;
	wire [4-1:0] node18904;
	wire [4-1:0] node18907;
	wire [4-1:0] node18908;
	wire [4-1:0] node18911;
	wire [4-1:0] node18914;
	wire [4-1:0] node18915;
	wire [4-1:0] node18916;
	wire [4-1:0] node18919;
	wire [4-1:0] node18922;
	wire [4-1:0] node18923;
	wire [4-1:0] node18926;
	wire [4-1:0] node18928;
	wire [4-1:0] node18931;
	wire [4-1:0] node18932;
	wire [4-1:0] node18933;
	wire [4-1:0] node18934;
	wire [4-1:0] node18935;
	wire [4-1:0] node18939;
	wire [4-1:0] node18940;
	wire [4-1:0] node18944;
	wire [4-1:0] node18945;
	wire [4-1:0] node18946;
	wire [4-1:0] node18949;
	wire [4-1:0] node18952;
	wire [4-1:0] node18954;
	wire [4-1:0] node18957;
	wire [4-1:0] node18958;
	wire [4-1:0] node18959;
	wire [4-1:0] node18962;
	wire [4-1:0] node18965;
	wire [4-1:0] node18966;
	wire [4-1:0] node18969;
	wire [4-1:0] node18972;
	wire [4-1:0] node18973;
	wire [4-1:0] node18974;
	wire [4-1:0] node18975;
	wire [4-1:0] node18977;
	wire [4-1:0] node18978;
	wire [4-1:0] node18982;
	wire [4-1:0] node18983;
	wire [4-1:0] node18984;
	wire [4-1:0] node18988;
	wire [4-1:0] node18989;
	wire [4-1:0] node18992;
	wire [4-1:0] node18995;
	wire [4-1:0] node18996;
	wire [4-1:0] node18997;
	wire [4-1:0] node18999;
	wire [4-1:0] node19002;
	wire [4-1:0] node19003;
	wire [4-1:0] node19007;
	wire [4-1:0] node19009;
	wire [4-1:0] node19012;
	wire [4-1:0] node19013;
	wire [4-1:0] node19014;
	wire [4-1:0] node19015;
	wire [4-1:0] node19018;
	wire [4-1:0] node19021;
	wire [4-1:0] node19022;
	wire [4-1:0] node19024;
	wire [4-1:0] node19027;
	wire [4-1:0] node19028;
	wire [4-1:0] node19032;
	wire [4-1:0] node19033;
	wire [4-1:0] node19034;
	wire [4-1:0] node19037;
	wire [4-1:0] node19040;
	wire [4-1:0] node19041;
	wire [4-1:0] node19042;
	wire [4-1:0] node19046;
	wire [4-1:0] node19049;
	wire [4-1:0] node19050;
	wire [4-1:0] node19051;
	wire [4-1:0] node19052;
	wire [4-1:0] node19053;
	wire [4-1:0] node19054;
	wire [4-1:0] node19055;
	wire [4-1:0] node19059;
	wire [4-1:0] node19060;
	wire [4-1:0] node19063;
	wire [4-1:0] node19066;
	wire [4-1:0] node19067;
	wire [4-1:0] node19070;
	wire [4-1:0] node19073;
	wire [4-1:0] node19074;
	wire [4-1:0] node19075;
	wire [4-1:0] node19078;
	wire [4-1:0] node19081;
	wire [4-1:0] node19083;
	wire [4-1:0] node19086;
	wire [4-1:0] node19087;
	wire [4-1:0] node19088;
	wire [4-1:0] node19089;
	wire [4-1:0] node19094;
	wire [4-1:0] node19095;
	wire [4-1:0] node19098;
	wire [4-1:0] node19101;
	wire [4-1:0] node19102;
	wire [4-1:0] node19103;
	wire [4-1:0] node19104;
	wire [4-1:0] node19107;
	wire [4-1:0] node19109;
	wire [4-1:0] node19112;
	wire [4-1:0] node19113;
	wire [4-1:0] node19115;
	wire [4-1:0] node19116;
	wire [4-1:0] node19120;
	wire [4-1:0] node19121;
	wire [4-1:0] node19122;
	wire [4-1:0] node19125;
	wire [4-1:0] node19128;
	wire [4-1:0] node19130;
	wire [4-1:0] node19133;
	wire [4-1:0] node19134;
	wire [4-1:0] node19137;
	wire [4-1:0] node19138;
	wire [4-1:0] node19140;
	wire [4-1:0] node19143;
	wire [4-1:0] node19144;
	wire [4-1:0] node19148;
	wire [4-1:0] node19149;
	wire [4-1:0] node19150;
	wire [4-1:0] node19151;
	wire [4-1:0] node19152;
	wire [4-1:0] node19153;
	wire [4-1:0] node19154;
	wire [4-1:0] node19157;
	wire [4-1:0] node19159;
	wire [4-1:0] node19162;
	wire [4-1:0] node19163;
	wire [4-1:0] node19166;
	wire [4-1:0] node19168;
	wire [4-1:0] node19171;
	wire [4-1:0] node19172;
	wire [4-1:0] node19173;
	wire [4-1:0] node19174;
	wire [4-1:0] node19177;
	wire [4-1:0] node19180;
	wire [4-1:0] node19181;
	wire [4-1:0] node19185;
	wire [4-1:0] node19186;
	wire [4-1:0] node19189;
	wire [4-1:0] node19190;
	wire [4-1:0] node19191;
	wire [4-1:0] node19194;
	wire [4-1:0] node19197;
	wire [4-1:0] node19198;
	wire [4-1:0] node19201;
	wire [4-1:0] node19204;
	wire [4-1:0] node19205;
	wire [4-1:0] node19206;
	wire [4-1:0] node19207;
	wire [4-1:0] node19208;
	wire [4-1:0] node19211;
	wire [4-1:0] node19215;
	wire [4-1:0] node19216;
	wire [4-1:0] node19218;
	wire [4-1:0] node19219;
	wire [4-1:0] node19223;
	wire [4-1:0] node19224;
	wire [4-1:0] node19227;
	wire [4-1:0] node19230;
	wire [4-1:0] node19231;
	wire [4-1:0] node19232;
	wire [4-1:0] node19235;
	wire [4-1:0] node19237;
	wire [4-1:0] node19240;
	wire [4-1:0] node19241;
	wire [4-1:0] node19243;
	wire [4-1:0] node19244;
	wire [4-1:0] node19247;
	wire [4-1:0] node19250;
	wire [4-1:0] node19251;
	wire [4-1:0] node19255;
	wire [4-1:0] node19256;
	wire [4-1:0] node19257;
	wire [4-1:0] node19258;
	wire [4-1:0] node19260;
	wire [4-1:0] node19262;
	wire [4-1:0] node19263;
	wire [4-1:0] node19267;
	wire [4-1:0] node19268;
	wire [4-1:0] node19269;
	wire [4-1:0] node19272;
	wire [4-1:0] node19275;
	wire [4-1:0] node19276;
	wire [4-1:0] node19277;
	wire [4-1:0] node19282;
	wire [4-1:0] node19283;
	wire [4-1:0] node19284;
	wire [4-1:0] node19286;
	wire [4-1:0] node19287;
	wire [4-1:0] node19290;
	wire [4-1:0] node19293;
	wire [4-1:0] node19295;
	wire [4-1:0] node19298;
	wire [4-1:0] node19299;
	wire [4-1:0] node19300;
	wire [4-1:0] node19301;
	wire [4-1:0] node19307;
	wire [4-1:0] node19308;
	wire [4-1:0] node19309;
	wire [4-1:0] node19310;
	wire [4-1:0] node19314;
	wire [4-1:0] node19315;
	wire [4-1:0] node19317;
	wire [4-1:0] node19318;
	wire [4-1:0] node19321;
	wire [4-1:0] node19324;
	wire [4-1:0] node19325;
	wire [4-1:0] node19326;
	wire [4-1:0] node19330;
	wire [4-1:0] node19331;
	wire [4-1:0] node19335;
	wire [4-1:0] node19336;
	wire [4-1:0] node19337;
	wire [4-1:0] node19339;
	wire [4-1:0] node19342;
	wire [4-1:0] node19343;
	wire [4-1:0] node19346;
	wire [4-1:0] node19347;
	wire [4-1:0] node19351;
	wire [4-1:0] node19352;
	wire [4-1:0] node19354;
	wire [4-1:0] node19355;
	wire [4-1:0] node19358;
	wire [4-1:0] node19361;
	wire [4-1:0] node19363;
	wire [4-1:0] node19366;
	wire [4-1:0] node19367;
	wire [4-1:0] node19368;
	wire [4-1:0] node19369;
	wire [4-1:0] node19370;
	wire [4-1:0] node19371;
	wire [4-1:0] node19372;
	wire [4-1:0] node19373;
	wire [4-1:0] node19376;
	wire [4-1:0] node19379;
	wire [4-1:0] node19382;
	wire [4-1:0] node19384;
	wire [4-1:0] node19387;
	wire [4-1:0] node19388;
	wire [4-1:0] node19389;
	wire [4-1:0] node19390;
	wire [4-1:0] node19393;
	wire [4-1:0] node19397;
	wire [4-1:0] node19399;
	wire [4-1:0] node19400;
	wire [4-1:0] node19403;
	wire [4-1:0] node19406;
	wire [4-1:0] node19407;
	wire [4-1:0] node19408;
	wire [4-1:0] node19409;
	wire [4-1:0] node19412;
	wire [4-1:0] node19413;
	wire [4-1:0] node19417;
	wire [4-1:0] node19418;
	wire [4-1:0] node19421;
	wire [4-1:0] node19424;
	wire [4-1:0] node19425;
	wire [4-1:0] node19426;
	wire [4-1:0] node19429;
	wire [4-1:0] node19430;
	wire [4-1:0] node19434;
	wire [4-1:0] node19435;
	wire [4-1:0] node19438;
	wire [4-1:0] node19441;
	wire [4-1:0] node19442;
	wire [4-1:0] node19443;
	wire [4-1:0] node19444;
	wire [4-1:0] node19445;
	wire [4-1:0] node19446;
	wire [4-1:0] node19449;
	wire [4-1:0] node19452;
	wire [4-1:0] node19453;
	wire [4-1:0] node19457;
	wire [4-1:0] node19459;
	wire [4-1:0] node19460;
	wire [4-1:0] node19463;
	wire [4-1:0] node19466;
	wire [4-1:0] node19467;
	wire [4-1:0] node19468;
	wire [4-1:0] node19469;
	wire [4-1:0] node19473;
	wire [4-1:0] node19474;
	wire [4-1:0] node19477;
	wire [4-1:0] node19480;
	wire [4-1:0] node19482;
	wire [4-1:0] node19483;
	wire [4-1:0] node19487;
	wire [4-1:0] node19488;
	wire [4-1:0] node19489;
	wire [4-1:0] node19491;
	wire [4-1:0] node19492;
	wire [4-1:0] node19495;
	wire [4-1:0] node19498;
	wire [4-1:0] node19499;
	wire [4-1:0] node19503;
	wire [4-1:0] node19504;
	wire [4-1:0] node19505;
	wire [4-1:0] node19507;
	wire [4-1:0] node19510;
	wire [4-1:0] node19512;
	wire [4-1:0] node19515;
	wire [4-1:0] node19517;
	wire [4-1:0] node19520;
	wire [4-1:0] node19521;
	wire [4-1:0] node19522;
	wire [4-1:0] node19523;
	wire [4-1:0] node19524;
	wire [4-1:0] node19527;
	wire [4-1:0] node19529;
	wire [4-1:0] node19531;
	wire [4-1:0] node19534;
	wire [4-1:0] node19535;
	wire [4-1:0] node19537;
	wire [4-1:0] node19538;
	wire [4-1:0] node19541;
	wire [4-1:0] node19544;
	wire [4-1:0] node19545;
	wire [4-1:0] node19546;
	wire [4-1:0] node19549;
	wire [4-1:0] node19553;
	wire [4-1:0] node19554;
	wire [4-1:0] node19555;
	wire [4-1:0] node19557;
	wire [4-1:0] node19558;
	wire [4-1:0] node19562;
	wire [4-1:0] node19563;
	wire [4-1:0] node19566;
	wire [4-1:0] node19569;
	wire [4-1:0] node19570;
	wire [4-1:0] node19572;
	wire [4-1:0] node19573;
	wire [4-1:0] node19577;
	wire [4-1:0] node19578;
	wire [4-1:0] node19582;
	wire [4-1:0] node19583;
	wire [4-1:0] node19584;
	wire [4-1:0] node19585;
	wire [4-1:0] node19588;
	wire [4-1:0] node19590;
	wire [4-1:0] node19591;
	wire [4-1:0] node19594;
	wire [4-1:0] node19597;
	wire [4-1:0] node19598;
	wire [4-1:0] node19599;
	wire [4-1:0] node19601;
	wire [4-1:0] node19604;
	wire [4-1:0] node19607;
	wire [4-1:0] node19608;
	wire [4-1:0] node19611;
	wire [4-1:0] node19614;
	wire [4-1:0] node19615;
	wire [4-1:0] node19616;
	wire [4-1:0] node19618;
	wire [4-1:0] node19619;
	wire [4-1:0] node19623;
	wire [4-1:0] node19624;
	wire [4-1:0] node19625;
	wire [4-1:0] node19629;
	wire [4-1:0] node19632;
	wire [4-1:0] node19633;
	wire [4-1:0] node19634;
	wire [4-1:0] node19635;
	wire [4-1:0] node19639;
	wire [4-1:0] node19642;
	wire [4-1:0] node19643;
	wire [4-1:0] node19646;
	wire [4-1:0] node19647;
	wire [4-1:0] node19650;
	wire [4-1:0] node19653;
	wire [4-1:0] node19654;
	wire [4-1:0] node19655;
	wire [4-1:0] node19656;
	wire [4-1:0] node19657;
	wire [4-1:0] node19658;
	wire [4-1:0] node19659;
	wire [4-1:0] node19660;
	wire [4-1:0] node19661;
	wire [4-1:0] node19665;
	wire [4-1:0] node19666;
	wire [4-1:0] node19669;
	wire [4-1:0] node19671;
	wire [4-1:0] node19674;
	wire [4-1:0] node19675;
	wire [4-1:0] node19676;
	wire [4-1:0] node19679;
	wire [4-1:0] node19682;
	wire [4-1:0] node19683;
	wire [4-1:0] node19684;
	wire [4-1:0] node19687;
	wire [4-1:0] node19690;
	wire [4-1:0] node19691;
	wire [4-1:0] node19695;
	wire [4-1:0] node19696;
	wire [4-1:0] node19697;
	wire [4-1:0] node19698;
	wire [4-1:0] node19701;
	wire [4-1:0] node19705;
	wire [4-1:0] node19706;
	wire [4-1:0] node19708;
	wire [4-1:0] node19709;
	wire [4-1:0] node19712;
	wire [4-1:0] node19715;
	wire [4-1:0] node19716;
	wire [4-1:0] node19720;
	wire [4-1:0] node19721;
	wire [4-1:0] node19722;
	wire [4-1:0] node19723;
	wire [4-1:0] node19724;
	wire [4-1:0] node19727;
	wire [4-1:0] node19730;
	wire [4-1:0] node19731;
	wire [4-1:0] node19734;
	wire [4-1:0] node19737;
	wire [4-1:0] node19738;
	wire [4-1:0] node19739;
	wire [4-1:0] node19742;
	wire [4-1:0] node19745;
	wire [4-1:0] node19747;
	wire [4-1:0] node19750;
	wire [4-1:0] node19751;
	wire [4-1:0] node19752;
	wire [4-1:0] node19753;
	wire [4-1:0] node19756;
	wire [4-1:0] node19759;
	wire [4-1:0] node19760;
	wire [4-1:0] node19763;
	wire [4-1:0] node19766;
	wire [4-1:0] node19767;
	wire [4-1:0] node19768;
	wire [4-1:0] node19771;
	wire [4-1:0] node19775;
	wire [4-1:0] node19776;
	wire [4-1:0] node19777;
	wire [4-1:0] node19778;
	wire [4-1:0] node19779;
	wire [4-1:0] node19780;
	wire [4-1:0] node19785;
	wire [4-1:0] node19786;
	wire [4-1:0] node19787;
	wire [4-1:0] node19790;
	wire [4-1:0] node19793;
	wire [4-1:0] node19795;
	wire [4-1:0] node19796;
	wire [4-1:0] node19799;
	wire [4-1:0] node19802;
	wire [4-1:0] node19803;
	wire [4-1:0] node19804;
	wire [4-1:0] node19805;
	wire [4-1:0] node19809;
	wire [4-1:0] node19810;
	wire [4-1:0] node19811;
	wire [4-1:0] node19814;
	wire [4-1:0] node19817;
	wire [4-1:0] node19820;
	wire [4-1:0] node19821;
	wire [4-1:0] node19822;
	wire [4-1:0] node19826;
	wire [4-1:0] node19827;
	wire [4-1:0] node19828;
	wire [4-1:0] node19832;
	wire [4-1:0] node19833;
	wire [4-1:0] node19836;
	wire [4-1:0] node19839;
	wire [4-1:0] node19840;
	wire [4-1:0] node19841;
	wire [4-1:0] node19842;
	wire [4-1:0] node19843;
	wire [4-1:0] node19845;
	wire [4-1:0] node19848;
	wire [4-1:0] node19851;
	wire [4-1:0] node19853;
	wire [4-1:0] node19856;
	wire [4-1:0] node19857;
	wire [4-1:0] node19859;
	wire [4-1:0] node19861;
	wire [4-1:0] node19864;
	wire [4-1:0] node19865;
	wire [4-1:0] node19867;
	wire [4-1:0] node19870;
	wire [4-1:0] node19871;
	wire [4-1:0] node19874;
	wire [4-1:0] node19877;
	wire [4-1:0] node19878;
	wire [4-1:0] node19879;
	wire [4-1:0] node19880;
	wire [4-1:0] node19881;
	wire [4-1:0] node19885;
	wire [4-1:0] node19886;
	wire [4-1:0] node19890;
	wire [4-1:0] node19891;
	wire [4-1:0] node19894;
	wire [4-1:0] node19897;
	wire [4-1:0] node19898;
	wire [4-1:0] node19900;
	wire [4-1:0] node19901;
	wire [4-1:0] node19905;
	wire [4-1:0] node19907;
	wire [4-1:0] node19908;
	wire [4-1:0] node19912;
	wire [4-1:0] node19913;
	wire [4-1:0] node19914;
	wire [4-1:0] node19915;
	wire [4-1:0] node19916;
	wire [4-1:0] node19917;
	wire [4-1:0] node19919;
	wire [4-1:0] node19921;
	wire [4-1:0] node19924;
	wire [4-1:0] node19925;
	wire [4-1:0] node19926;
	wire [4-1:0] node19929;
	wire [4-1:0] node19933;
	wire [4-1:0] node19934;
	wire [4-1:0] node19935;
	wire [4-1:0] node19939;
	wire [4-1:0] node19941;
	wire [4-1:0] node19944;
	wire [4-1:0] node19945;
	wire [4-1:0] node19946;
	wire [4-1:0] node19947;
	wire [4-1:0] node19950;
	wire [4-1:0] node19953;
	wire [4-1:0] node19955;
	wire [4-1:0] node19958;
	wire [4-1:0] node19959;
	wire [4-1:0] node19960;
	wire [4-1:0] node19963;
	wire [4-1:0] node19966;
	wire [4-1:0] node19967;
	wire [4-1:0] node19970;
	wire [4-1:0] node19973;
	wire [4-1:0] node19974;
	wire [4-1:0] node19975;
	wire [4-1:0] node19976;
	wire [4-1:0] node19977;
	wire [4-1:0] node19980;
	wire [4-1:0] node19983;
	wire [4-1:0] node19985;
	wire [4-1:0] node19988;
	wire [4-1:0] node19989;
	wire [4-1:0] node19990;
	wire [4-1:0] node19991;
	wire [4-1:0] node19994;
	wire [4-1:0] node19997;
	wire [4-1:0] node19998;
	wire [4-1:0] node20001;
	wire [4-1:0] node20004;
	wire [4-1:0] node20005;
	wire [4-1:0] node20007;
	wire [4-1:0] node20011;
	wire [4-1:0] node20012;
	wire [4-1:0] node20013;
	wire [4-1:0] node20014;
	wire [4-1:0] node20018;
	wire [4-1:0] node20021;
	wire [4-1:0] node20022;
	wire [4-1:0] node20024;
	wire [4-1:0] node20025;
	wire [4-1:0] node20028;
	wire [4-1:0] node20031;
	wire [4-1:0] node20032;
	wire [4-1:0] node20036;
	wire [4-1:0] node20037;
	wire [4-1:0] node20038;
	wire [4-1:0] node20039;
	wire [4-1:0] node20040;
	wire [4-1:0] node20041;
	wire [4-1:0] node20044;
	wire [4-1:0] node20047;
	wire [4-1:0] node20048;
	wire [4-1:0] node20051;
	wire [4-1:0] node20054;
	wire [4-1:0] node20055;
	wire [4-1:0] node20056;
	wire [4-1:0] node20059;
	wire [4-1:0] node20062;
	wire [4-1:0] node20064;
	wire [4-1:0] node20067;
	wire [4-1:0] node20068;
	wire [4-1:0] node20069;
	wire [4-1:0] node20070;
	wire [4-1:0] node20073;
	wire [4-1:0] node20076;
	wire [4-1:0] node20078;
	wire [4-1:0] node20080;
	wire [4-1:0] node20083;
	wire [4-1:0] node20084;
	wire [4-1:0] node20085;
	wire [4-1:0] node20088;
	wire [4-1:0] node20091;
	wire [4-1:0] node20092;
	wire [4-1:0] node20094;
	wire [4-1:0] node20097;
	wire [4-1:0] node20098;
	wire [4-1:0] node20101;
	wire [4-1:0] node20104;
	wire [4-1:0] node20105;
	wire [4-1:0] node20106;
	wire [4-1:0] node20107;
	wire [4-1:0] node20108;
	wire [4-1:0] node20111;
	wire [4-1:0] node20114;
	wire [4-1:0] node20116;
	wire [4-1:0] node20117;
	wire [4-1:0] node20120;
	wire [4-1:0] node20123;
	wire [4-1:0] node20124;
	wire [4-1:0] node20125;
	wire [4-1:0] node20128;
	wire [4-1:0] node20131;
	wire [4-1:0] node20132;
	wire [4-1:0] node20135;
	wire [4-1:0] node20138;
	wire [4-1:0] node20139;
	wire [4-1:0] node20140;
	wire [4-1:0] node20141;
	wire [4-1:0] node20144;
	wire [4-1:0] node20147;
	wire [4-1:0] node20149;
	wire [4-1:0] node20152;
	wire [4-1:0] node20153;
	wire [4-1:0] node20154;
	wire [4-1:0] node20155;
	wire [4-1:0] node20158;
	wire [4-1:0] node20161;
	wire [4-1:0] node20163;
	wire [4-1:0] node20166;
	wire [4-1:0] node20168;
	wire [4-1:0] node20171;
	wire [4-1:0] node20172;
	wire [4-1:0] node20173;
	wire [4-1:0] node20174;
	wire [4-1:0] node20175;
	wire [4-1:0] node20176;
	wire [4-1:0] node20177;
	wire [4-1:0] node20178;
	wire [4-1:0] node20181;
	wire [4-1:0] node20184;
	wire [4-1:0] node20185;
	wire [4-1:0] node20188;
	wire [4-1:0] node20191;
	wire [4-1:0] node20192;
	wire [4-1:0] node20194;
	wire [4-1:0] node20197;
	wire [4-1:0] node20199;
	wire [4-1:0] node20200;
	wire [4-1:0] node20203;
	wire [4-1:0] node20206;
	wire [4-1:0] node20207;
	wire [4-1:0] node20208;
	wire [4-1:0] node20209;
	wire [4-1:0] node20211;
	wire [4-1:0] node20214;
	wire [4-1:0] node20215;
	wire [4-1:0] node20218;
	wire [4-1:0] node20221;
	wire [4-1:0] node20222;
	wire [4-1:0] node20224;
	wire [4-1:0] node20227;
	wire [4-1:0] node20228;
	wire [4-1:0] node20232;
	wire [4-1:0] node20233;
	wire [4-1:0] node20235;
	wire [4-1:0] node20237;
	wire [4-1:0] node20240;
	wire [4-1:0] node20241;
	wire [4-1:0] node20245;
	wire [4-1:0] node20246;
	wire [4-1:0] node20247;
	wire [4-1:0] node20248;
	wire [4-1:0] node20249;
	wire [4-1:0] node20250;
	wire [4-1:0] node20253;
	wire [4-1:0] node20256;
	wire [4-1:0] node20258;
	wire [4-1:0] node20261;
	wire [4-1:0] node20263;
	wire [4-1:0] node20264;
	wire [4-1:0] node20267;
	wire [4-1:0] node20270;
	wire [4-1:0] node20271;
	wire [4-1:0] node20273;
	wire [4-1:0] node20276;
	wire [4-1:0] node20277;
	wire [4-1:0] node20278;
	wire [4-1:0] node20281;
	wire [4-1:0] node20284;
	wire [4-1:0] node20285;
	wire [4-1:0] node20288;
	wire [4-1:0] node20291;
	wire [4-1:0] node20292;
	wire [4-1:0] node20293;
	wire [4-1:0] node20294;
	wire [4-1:0] node20296;
	wire [4-1:0] node20300;
	wire [4-1:0] node20301;
	wire [4-1:0] node20302;
	wire [4-1:0] node20305;
	wire [4-1:0] node20308;
	wire [4-1:0] node20309;
	wire [4-1:0] node20313;
	wire [4-1:0] node20314;
	wire [4-1:0] node20315;
	wire [4-1:0] node20317;
	wire [4-1:0] node20320;
	wire [4-1:0] node20321;
	wire [4-1:0] node20324;
	wire [4-1:0] node20327;
	wire [4-1:0] node20329;
	wire [4-1:0] node20330;
	wire [4-1:0] node20334;
	wire [4-1:0] node20335;
	wire [4-1:0] node20336;
	wire [4-1:0] node20337;
	wire [4-1:0] node20338;
	wire [4-1:0] node20339;
	wire [4-1:0] node20343;
	wire [4-1:0] node20344;
	wire [4-1:0] node20345;
	wire [4-1:0] node20349;
	wire [4-1:0] node20351;
	wire [4-1:0] node20354;
	wire [4-1:0] node20355;
	wire [4-1:0] node20356;
	wire [4-1:0] node20360;
	wire [4-1:0] node20362;
	wire [4-1:0] node20364;
	wire [4-1:0] node20367;
	wire [4-1:0] node20368;
	wire [4-1:0] node20369;
	wire [4-1:0] node20370;
	wire [4-1:0] node20371;
	wire [4-1:0] node20375;
	wire [4-1:0] node20376;
	wire [4-1:0] node20380;
	wire [4-1:0] node20382;
	wire [4-1:0] node20385;
	wire [4-1:0] node20386;
	wire [4-1:0] node20387;
	wire [4-1:0] node20391;
	wire [4-1:0] node20392;
	wire [4-1:0] node20395;
	wire [4-1:0] node20398;
	wire [4-1:0] node20399;
	wire [4-1:0] node20400;
	wire [4-1:0] node20401;
	wire [4-1:0] node20402;
	wire [4-1:0] node20405;
	wire [4-1:0] node20408;
	wire [4-1:0] node20411;
	wire [4-1:0] node20413;
	wire [4-1:0] node20414;
	wire [4-1:0] node20416;
	wire [4-1:0] node20419;
	wire [4-1:0] node20420;
	wire [4-1:0] node20424;
	wire [4-1:0] node20425;
	wire [4-1:0] node20426;
	wire [4-1:0] node20427;
	wire [4-1:0] node20430;
	wire [4-1:0] node20433;
	wire [4-1:0] node20434;
	wire [4-1:0] node20437;
	wire [4-1:0] node20440;
	wire [4-1:0] node20441;
	wire [4-1:0] node20443;
	wire [4-1:0] node20446;
	wire [4-1:0] node20447;
	wire [4-1:0] node20448;
	wire [4-1:0] node20452;
	wire [4-1:0] node20455;
	wire [4-1:0] node20456;
	wire [4-1:0] node20457;
	wire [4-1:0] node20458;
	wire [4-1:0] node20459;
	wire [4-1:0] node20460;
	wire [4-1:0] node20461;
	wire [4-1:0] node20464;
	wire [4-1:0] node20467;
	wire [4-1:0] node20468;
	wire [4-1:0] node20469;
	wire [4-1:0] node20472;
	wire [4-1:0] node20476;
	wire [4-1:0] node20477;
	wire [4-1:0] node20478;
	wire [4-1:0] node20481;
	wire [4-1:0] node20484;
	wire [4-1:0] node20485;
	wire [4-1:0] node20487;
	wire [4-1:0] node20490;
	wire [4-1:0] node20493;
	wire [4-1:0] node20494;
	wire [4-1:0] node20495;
	wire [4-1:0] node20496;
	wire [4-1:0] node20499;
	wire [4-1:0] node20502;
	wire [4-1:0] node20504;
	wire [4-1:0] node20507;
	wire [4-1:0] node20508;
	wire [4-1:0] node20510;
	wire [4-1:0] node20512;
	wire [4-1:0] node20515;
	wire [4-1:0] node20516;
	wire [4-1:0] node20519;
	wire [4-1:0] node20522;
	wire [4-1:0] node20523;
	wire [4-1:0] node20524;
	wire [4-1:0] node20525;
	wire [4-1:0] node20526;
	wire [4-1:0] node20530;
	wire [4-1:0] node20531;
	wire [4-1:0] node20532;
	wire [4-1:0] node20536;
	wire [4-1:0] node20539;
	wire [4-1:0] node20540;
	wire [4-1:0] node20541;
	wire [4-1:0] node20544;
	wire [4-1:0] node20547;
	wire [4-1:0] node20548;
	wire [4-1:0] node20552;
	wire [4-1:0] node20553;
	wire [4-1:0] node20554;
	wire [4-1:0] node20555;
	wire [4-1:0] node20558;
	wire [4-1:0] node20561;
	wire [4-1:0] node20563;
	wire [4-1:0] node20566;
	wire [4-1:0] node20567;
	wire [4-1:0] node20568;
	wire [4-1:0] node20571;
	wire [4-1:0] node20572;
	wire [4-1:0] node20576;
	wire [4-1:0] node20577;
	wire [4-1:0] node20578;
	wire [4-1:0] node20581;
	wire [4-1:0] node20584;
	wire [4-1:0] node20585;
	wire [4-1:0] node20588;
	wire [4-1:0] node20591;
	wire [4-1:0] node20592;
	wire [4-1:0] node20593;
	wire [4-1:0] node20594;
	wire [4-1:0] node20596;
	wire [4-1:0] node20597;
	wire [4-1:0] node20601;
	wire [4-1:0] node20602;
	wire [4-1:0] node20603;
	wire [4-1:0] node20606;
	wire [4-1:0] node20609;
	wire [4-1:0] node20610;
	wire [4-1:0] node20614;
	wire [4-1:0] node20615;
	wire [4-1:0] node20616;
	wire [4-1:0] node20617;
	wire [4-1:0] node20620;
	wire [4-1:0] node20623;
	wire [4-1:0] node20624;
	wire [4-1:0] node20627;
	wire [4-1:0] node20630;
	wire [4-1:0] node20631;
	wire [4-1:0] node20634;
	wire [4-1:0] node20635;
	wire [4-1:0] node20638;
	wire [4-1:0] node20641;
	wire [4-1:0] node20642;
	wire [4-1:0] node20643;
	wire [4-1:0] node20644;
	wire [4-1:0] node20648;
	wire [4-1:0] node20649;
	wire [4-1:0] node20650;
	wire [4-1:0] node20654;
	wire [4-1:0] node20657;
	wire [4-1:0] node20658;
	wire [4-1:0] node20659;
	wire [4-1:0] node20660;
	wire [4-1:0] node20663;
	wire [4-1:0] node20666;
	wire [4-1:0] node20668;
	wire [4-1:0] node20671;
	wire [4-1:0] node20672;
	wire [4-1:0] node20673;
	wire [4-1:0] node20676;
	wire [4-1:0] node20679;
	wire [4-1:0] node20680;
	wire [4-1:0] node20681;
	wire [4-1:0] node20686;
	wire [4-1:0] node20687;
	wire [4-1:0] node20688;
	wire [4-1:0] node20689;
	wire [4-1:0] node20690;
	wire [4-1:0] node20691;
	wire [4-1:0] node20692;
	wire [4-1:0] node20693;
	wire [4-1:0] node20694;
	wire [4-1:0] node20696;
	wire [4-1:0] node20697;
	wire [4-1:0] node20700;
	wire [4-1:0] node20703;
	wire [4-1:0] node20704;
	wire [4-1:0] node20705;
	wire [4-1:0] node20709;
	wire [4-1:0] node20710;
	wire [4-1:0] node20713;
	wire [4-1:0] node20716;
	wire [4-1:0] node20717;
	wire [4-1:0] node20718;
	wire [4-1:0] node20719;
	wire [4-1:0] node20724;
	wire [4-1:0] node20725;
	wire [4-1:0] node20726;
	wire [4-1:0] node20729;
	wire [4-1:0] node20733;
	wire [4-1:0] node20734;
	wire [4-1:0] node20735;
	wire [4-1:0] node20737;
	wire [4-1:0] node20738;
	wire [4-1:0] node20741;
	wire [4-1:0] node20744;
	wire [4-1:0] node20745;
	wire [4-1:0] node20747;
	wire [4-1:0] node20751;
	wire [4-1:0] node20752;
	wire [4-1:0] node20754;
	wire [4-1:0] node20755;
	wire [4-1:0] node20758;
	wire [4-1:0] node20761;
	wire [4-1:0] node20764;
	wire [4-1:0] node20765;
	wire [4-1:0] node20766;
	wire [4-1:0] node20767;
	wire [4-1:0] node20768;
	wire [4-1:0] node20770;
	wire [4-1:0] node20773;
	wire [4-1:0] node20775;
	wire [4-1:0] node20778;
	wire [4-1:0] node20779;
	wire [4-1:0] node20780;
	wire [4-1:0] node20783;
	wire [4-1:0] node20786;
	wire [4-1:0] node20787;
	wire [4-1:0] node20791;
	wire [4-1:0] node20792;
	wire [4-1:0] node20793;
	wire [4-1:0] node20795;
	wire [4-1:0] node20799;
	wire [4-1:0] node20800;
	wire [4-1:0] node20802;
	wire [4-1:0] node20805;
	wire [4-1:0] node20806;
	wire [4-1:0] node20810;
	wire [4-1:0] node20811;
	wire [4-1:0] node20812;
	wire [4-1:0] node20813;
	wire [4-1:0] node20817;
	wire [4-1:0] node20818;
	wire [4-1:0] node20820;
	wire [4-1:0] node20823;
	wire [4-1:0] node20825;
	wire [4-1:0] node20828;
	wire [4-1:0] node20829;
	wire [4-1:0] node20830;
	wire [4-1:0] node20831;
	wire [4-1:0] node20834;
	wire [4-1:0] node20838;
	wire [4-1:0] node20839;
	wire [4-1:0] node20840;
	wire [4-1:0] node20843;
	wire [4-1:0] node20846;
	wire [4-1:0] node20847;
	wire [4-1:0] node20850;
	wire [4-1:0] node20853;
	wire [4-1:0] node20854;
	wire [4-1:0] node20855;
	wire [4-1:0] node20856;
	wire [4-1:0] node20857;
	wire [4-1:0] node20858;
	wire [4-1:0] node20861;
	wire [4-1:0] node20864;
	wire [4-1:0] node20866;
	wire [4-1:0] node20869;
	wire [4-1:0] node20870;
	wire [4-1:0] node20871;
	wire [4-1:0] node20874;
	wire [4-1:0] node20877;
	wire [4-1:0] node20879;
	wire [4-1:0] node20882;
	wire [4-1:0] node20883;
	wire [4-1:0] node20884;
	wire [4-1:0] node20885;
	wire [4-1:0] node20888;
	wire [4-1:0] node20891;
	wire [4-1:0] node20892;
	wire [4-1:0] node20896;
	wire [4-1:0] node20897;
	wire [4-1:0] node20899;
	wire [4-1:0] node20902;
	wire [4-1:0] node20904;
	wire [4-1:0] node20906;
	wire [4-1:0] node20909;
	wire [4-1:0] node20910;
	wire [4-1:0] node20911;
	wire [4-1:0] node20912;
	wire [4-1:0] node20915;
	wire [4-1:0] node20917;
	wire [4-1:0] node20918;
	wire [4-1:0] node20922;
	wire [4-1:0] node20923;
	wire [4-1:0] node20925;
	wire [4-1:0] node20926;
	wire [4-1:0] node20930;
	wire [4-1:0] node20931;
	wire [4-1:0] node20932;
	wire [4-1:0] node20935;
	wire [4-1:0] node20938;
	wire [4-1:0] node20940;
	wire [4-1:0] node20943;
	wire [4-1:0] node20944;
	wire [4-1:0] node20945;
	wire [4-1:0] node20946;
	wire [4-1:0] node20947;
	wire [4-1:0] node20951;
	wire [4-1:0] node20952;
	wire [4-1:0] node20956;
	wire [4-1:0] node20957;
	wire [4-1:0] node20958;
	wire [4-1:0] node20962;
	wire [4-1:0] node20963;
	wire [4-1:0] node20967;
	wire [4-1:0] node20968;
	wire [4-1:0] node20969;
	wire [4-1:0] node20970;
	wire [4-1:0] node20973;
	wire [4-1:0] node20976;
	wire [4-1:0] node20978;
	wire [4-1:0] node20981;
	wire [4-1:0] node20984;
	wire [4-1:0] node20985;
	wire [4-1:0] node20986;
	wire [4-1:0] node20987;
	wire [4-1:0] node20988;
	wire [4-1:0] node20989;
	wire [4-1:0] node20991;
	wire [4-1:0] node20993;
	wire [4-1:0] node20996;
	wire [4-1:0] node20997;
	wire [4-1:0] node20998;
	wire [4-1:0] node21002;
	wire [4-1:0] node21004;
	wire [4-1:0] node21007;
	wire [4-1:0] node21008;
	wire [4-1:0] node21011;
	wire [4-1:0] node21012;
	wire [4-1:0] node21015;
	wire [4-1:0] node21018;
	wire [4-1:0] node21019;
	wire [4-1:0] node21020;
	wire [4-1:0] node21022;
	wire [4-1:0] node21025;
	wire [4-1:0] node21028;
	wire [4-1:0] node21029;
	wire [4-1:0] node21030;
	wire [4-1:0] node21031;
	wire [4-1:0] node21035;
	wire [4-1:0] node21036;
	wire [4-1:0] node21040;
	wire [4-1:0] node21042;
	wire [4-1:0] node21044;
	wire [4-1:0] node21047;
	wire [4-1:0] node21048;
	wire [4-1:0] node21049;
	wire [4-1:0] node21050;
	wire [4-1:0] node21051;
	wire [4-1:0] node21052;
	wire [4-1:0] node21055;
	wire [4-1:0] node21058;
	wire [4-1:0] node21059;
	wire [4-1:0] node21063;
	wire [4-1:0] node21064;
	wire [4-1:0] node21066;
	wire [4-1:0] node21070;
	wire [4-1:0] node21071;
	wire [4-1:0] node21072;
	wire [4-1:0] node21073;
	wire [4-1:0] node21076;
	wire [4-1:0] node21079;
	wire [4-1:0] node21081;
	wire [4-1:0] node21084;
	wire [4-1:0] node21085;
	wire [4-1:0] node21086;
	wire [4-1:0] node21089;
	wire [4-1:0] node21093;
	wire [4-1:0] node21094;
	wire [4-1:0] node21095;
	wire [4-1:0] node21096;
	wire [4-1:0] node21100;
	wire [4-1:0] node21101;
	wire [4-1:0] node21104;
	wire [4-1:0] node21107;
	wire [4-1:0] node21108;
	wire [4-1:0] node21109;
	wire [4-1:0] node21112;
	wire [4-1:0] node21115;
	wire [4-1:0] node21117;
	wire [4-1:0] node21120;
	wire [4-1:0] node21121;
	wire [4-1:0] node21122;
	wire [4-1:0] node21123;
	wire [4-1:0] node21124;
	wire [4-1:0] node21125;
	wire [4-1:0] node21127;
	wire [4-1:0] node21130;
	wire [4-1:0] node21132;
	wire [4-1:0] node21135;
	wire [4-1:0] node21136;
	wire [4-1:0] node21137;
	wire [4-1:0] node21140;
	wire [4-1:0] node21143;
	wire [4-1:0] node21146;
	wire [4-1:0] node21147;
	wire [4-1:0] node21148;
	wire [4-1:0] node21149;
	wire [4-1:0] node21152;
	wire [4-1:0] node21155;
	wire [4-1:0] node21156;
	wire [4-1:0] node21160;
	wire [4-1:0] node21162;
	wire [4-1:0] node21163;
	wire [4-1:0] node21166;
	wire [4-1:0] node21169;
	wire [4-1:0] node21170;
	wire [4-1:0] node21171;
	wire [4-1:0] node21172;
	wire [4-1:0] node21174;
	wire [4-1:0] node21177;
	wire [4-1:0] node21178;
	wire [4-1:0] node21181;
	wire [4-1:0] node21184;
	wire [4-1:0] node21187;
	wire [4-1:0] node21188;
	wire [4-1:0] node21190;
	wire [4-1:0] node21192;
	wire [4-1:0] node21195;
	wire [4-1:0] node21196;
	wire [4-1:0] node21197;
	wire [4-1:0] node21201;
	wire [4-1:0] node21202;
	wire [4-1:0] node21205;
	wire [4-1:0] node21208;
	wire [4-1:0] node21209;
	wire [4-1:0] node21210;
	wire [4-1:0] node21211;
	wire [4-1:0] node21212;
	wire [4-1:0] node21213;
	wire [4-1:0] node21216;
	wire [4-1:0] node21220;
	wire [4-1:0] node21222;
	wire [4-1:0] node21223;
	wire [4-1:0] node21227;
	wire [4-1:0] node21229;
	wire [4-1:0] node21230;
	wire [4-1:0] node21231;
	wire [4-1:0] node21235;
	wire [4-1:0] node21236;
	wire [4-1:0] node21239;
	wire [4-1:0] node21242;
	wire [4-1:0] node21243;
	wire [4-1:0] node21244;
	wire [4-1:0] node21245;
	wire [4-1:0] node21249;
	wire [4-1:0] node21250;
	wire [4-1:0] node21253;
	wire [4-1:0] node21256;
	wire [4-1:0] node21257;
	wire [4-1:0] node21258;
	wire [4-1:0] node21260;
	wire [4-1:0] node21263;
	wire [4-1:0] node21264;
	wire [4-1:0] node21267;
	wire [4-1:0] node21270;
	wire [4-1:0] node21272;
	wire [4-1:0] node21273;
	wire [4-1:0] node21277;
	wire [4-1:0] node21278;
	wire [4-1:0] node21279;
	wire [4-1:0] node21280;
	wire [4-1:0] node21281;
	wire [4-1:0] node21282;
	wire [4-1:0] node21283;
	wire [4-1:0] node21285;
	wire [4-1:0] node21286;
	wire [4-1:0] node21289;
	wire [4-1:0] node21292;
	wire [4-1:0] node21293;
	wire [4-1:0] node21294;
	wire [4-1:0] node21298;
	wire [4-1:0] node21299;
	wire [4-1:0] node21302;
	wire [4-1:0] node21305;
	wire [4-1:0] node21306;
	wire [4-1:0] node21308;
	wire [4-1:0] node21309;
	wire [4-1:0] node21312;
	wire [4-1:0] node21315;
	wire [4-1:0] node21316;
	wire [4-1:0] node21320;
	wire [4-1:0] node21321;
	wire [4-1:0] node21322;
	wire [4-1:0] node21323;
	wire [4-1:0] node21324;
	wire [4-1:0] node21328;
	wire [4-1:0] node21330;
	wire [4-1:0] node21333;
	wire [4-1:0] node21335;
	wire [4-1:0] node21336;
	wire [4-1:0] node21339;
	wire [4-1:0] node21342;
	wire [4-1:0] node21343;
	wire [4-1:0] node21345;
	wire [4-1:0] node21347;
	wire [4-1:0] node21350;
	wire [4-1:0] node21351;
	wire [4-1:0] node21353;
	wire [4-1:0] node21357;
	wire [4-1:0] node21358;
	wire [4-1:0] node21359;
	wire [4-1:0] node21360;
	wire [4-1:0] node21361;
	wire [4-1:0] node21363;
	wire [4-1:0] node21366;
	wire [4-1:0] node21367;
	wire [4-1:0] node21371;
	wire [4-1:0] node21372;
	wire [4-1:0] node21374;
	wire [4-1:0] node21377;
	wire [4-1:0] node21378;
	wire [4-1:0] node21381;
	wire [4-1:0] node21384;
	wire [4-1:0] node21385;
	wire [4-1:0] node21387;
	wire [4-1:0] node21388;
	wire [4-1:0] node21392;
	wire [4-1:0] node21393;
	wire [4-1:0] node21394;
	wire [4-1:0] node21398;
	wire [4-1:0] node21399;
	wire [4-1:0] node21402;
	wire [4-1:0] node21405;
	wire [4-1:0] node21406;
	wire [4-1:0] node21407;
	wire [4-1:0] node21408;
	wire [4-1:0] node21409;
	wire [4-1:0] node21412;
	wire [4-1:0] node21415;
	wire [4-1:0] node21416;
	wire [4-1:0] node21420;
	wire [4-1:0] node21421;
	wire [4-1:0] node21423;
	wire [4-1:0] node21426;
	wire [4-1:0] node21427;
	wire [4-1:0] node21431;
	wire [4-1:0] node21432;
	wire [4-1:0] node21433;
	wire [4-1:0] node21434;
	wire [4-1:0] node21438;
	wire [4-1:0] node21439;
	wire [4-1:0] node21443;
	wire [4-1:0] node21444;
	wire [4-1:0] node21446;
	wire [4-1:0] node21449;
	wire [4-1:0] node21452;
	wire [4-1:0] node21453;
	wire [4-1:0] node21454;
	wire [4-1:0] node21455;
	wire [4-1:0] node21456;
	wire [4-1:0] node21458;
	wire [4-1:0] node21460;
	wire [4-1:0] node21463;
	wire [4-1:0] node21464;
	wire [4-1:0] node21466;
	wire [4-1:0] node21469;
	wire [4-1:0] node21470;
	wire [4-1:0] node21473;
	wire [4-1:0] node21476;
	wire [4-1:0] node21477;
	wire [4-1:0] node21478;
	wire [4-1:0] node21481;
	wire [4-1:0] node21482;
	wire [4-1:0] node21486;
	wire [4-1:0] node21487;
	wire [4-1:0] node21488;
	wire [4-1:0] node21491;
	wire [4-1:0] node21494;
	wire [4-1:0] node21495;
	wire [4-1:0] node21499;
	wire [4-1:0] node21500;
	wire [4-1:0] node21501;
	wire [4-1:0] node21503;
	wire [4-1:0] node21506;
	wire [4-1:0] node21507;
	wire [4-1:0] node21508;
	wire [4-1:0] node21511;
	wire [4-1:0] node21514;
	wire [4-1:0] node21515;
	wire [4-1:0] node21518;
	wire [4-1:0] node21521;
	wire [4-1:0] node21522;
	wire [4-1:0] node21523;
	wire [4-1:0] node21524;
	wire [4-1:0] node21527;
	wire [4-1:0] node21530;
	wire [4-1:0] node21531;
	wire [4-1:0] node21535;
	wire [4-1:0] node21536;
	wire [4-1:0] node21537;
	wire [4-1:0] node21541;
	wire [4-1:0] node21543;
	wire [4-1:0] node21546;
	wire [4-1:0] node21547;
	wire [4-1:0] node21548;
	wire [4-1:0] node21549;
	wire [4-1:0] node21550;
	wire [4-1:0] node21552;
	wire [4-1:0] node21555;
	wire [4-1:0] node21556;
	wire [4-1:0] node21560;
	wire [4-1:0] node21561;
	wire [4-1:0] node21562;
	wire [4-1:0] node21565;
	wire [4-1:0] node21568;
	wire [4-1:0] node21571;
	wire [4-1:0] node21572;
	wire [4-1:0] node21574;
	wire [4-1:0] node21575;
	wire [4-1:0] node21579;
	wire [4-1:0] node21581;
	wire [4-1:0] node21584;
	wire [4-1:0] node21585;
	wire [4-1:0] node21586;
	wire [4-1:0] node21587;
	wire [4-1:0] node21588;
	wire [4-1:0] node21591;
	wire [4-1:0] node21594;
	wire [4-1:0] node21597;
	wire [4-1:0] node21598;
	wire [4-1:0] node21599;
	wire [4-1:0] node21602;
	wire [4-1:0] node21605;
	wire [4-1:0] node21607;
	wire [4-1:0] node21610;
	wire [4-1:0] node21611;
	wire [4-1:0] node21614;
	wire [4-1:0] node21615;
	wire [4-1:0] node21617;
	wire [4-1:0] node21620;
	wire [4-1:0] node21623;
	wire [4-1:0] node21624;
	wire [4-1:0] node21625;
	wire [4-1:0] node21626;
	wire [4-1:0] node21627;
	wire [4-1:0] node21628;
	wire [4-1:0] node21631;
	wire [4-1:0] node21632;
	wire [4-1:0] node21635;
	wire [4-1:0] node21636;
	wire [4-1:0] node21640;
	wire [4-1:0] node21641;
	wire [4-1:0] node21642;
	wire [4-1:0] node21645;
	wire [4-1:0] node21648;
	wire [4-1:0] node21649;
	wire [4-1:0] node21651;
	wire [4-1:0] node21654;
	wire [4-1:0] node21657;
	wire [4-1:0] node21658;
	wire [4-1:0] node21659;
	wire [4-1:0] node21662;
	wire [4-1:0] node21664;
	wire [4-1:0] node21667;
	wire [4-1:0] node21669;
	wire [4-1:0] node21670;
	wire [4-1:0] node21672;
	wire [4-1:0] node21675;
	wire [4-1:0] node21678;
	wire [4-1:0] node21679;
	wire [4-1:0] node21680;
	wire [4-1:0] node21681;
	wire [4-1:0] node21683;
	wire [4-1:0] node21684;
	wire [4-1:0] node21687;
	wire [4-1:0] node21690;
	wire [4-1:0] node21691;
	wire [4-1:0] node21692;
	wire [4-1:0] node21697;
	wire [4-1:0] node21698;
	wire [4-1:0] node21699;
	wire [4-1:0] node21700;
	wire [4-1:0] node21706;
	wire [4-1:0] node21707;
	wire [4-1:0] node21708;
	wire [4-1:0] node21709;
	wire [4-1:0] node21710;
	wire [4-1:0] node21713;
	wire [4-1:0] node21716;
	wire [4-1:0] node21717;
	wire [4-1:0] node21720;
	wire [4-1:0] node21723;
	wire [4-1:0] node21724;
	wire [4-1:0] node21726;
	wire [4-1:0] node21729;
	wire [4-1:0] node21730;
	wire [4-1:0] node21733;
	wire [4-1:0] node21736;
	wire [4-1:0] node21737;
	wire [4-1:0] node21739;
	wire [4-1:0] node21740;
	wire [4-1:0] node21744;
	wire [4-1:0] node21745;
	wire [4-1:0] node21746;
	wire [4-1:0] node21751;
	wire [4-1:0] node21752;
	wire [4-1:0] node21753;
	wire [4-1:0] node21754;
	wire [4-1:0] node21755;
	wire [4-1:0] node21757;
	wire [4-1:0] node21758;
	wire [4-1:0] node21762;
	wire [4-1:0] node21763;
	wire [4-1:0] node21766;
	wire [4-1:0] node21767;
	wire [4-1:0] node21771;
	wire [4-1:0] node21772;
	wire [4-1:0] node21773;
	wire [4-1:0] node21777;
	wire [4-1:0] node21778;
	wire [4-1:0] node21779;
	wire [4-1:0] node21783;
	wire [4-1:0] node21784;
	wire [4-1:0] node21788;
	wire [4-1:0] node21789;
	wire [4-1:0] node21790;
	wire [4-1:0] node21791;
	wire [4-1:0] node21792;
	wire [4-1:0] node21795;
	wire [4-1:0] node21799;
	wire [4-1:0] node21800;
	wire [4-1:0] node21801;
	wire [4-1:0] node21805;
	wire [4-1:0] node21808;
	wire [4-1:0] node21809;
	wire [4-1:0] node21810;
	wire [4-1:0] node21813;
	wire [4-1:0] node21816;
	wire [4-1:0] node21817;
	wire [4-1:0] node21821;
	wire [4-1:0] node21822;
	wire [4-1:0] node21823;
	wire [4-1:0] node21824;
	wire [4-1:0] node21825;
	wire [4-1:0] node21828;
	wire [4-1:0] node21830;
	wire [4-1:0] node21833;
	wire [4-1:0] node21834;
	wire [4-1:0] node21836;
	wire [4-1:0] node21839;
	wire [4-1:0] node21841;
	wire [4-1:0] node21844;
	wire [4-1:0] node21845;
	wire [4-1:0] node21848;
	wire [4-1:0] node21849;
	wire [4-1:0] node21852;
	wire [4-1:0] node21853;
	wire [4-1:0] node21857;
	wire [4-1:0] node21858;
	wire [4-1:0] node21859;
	wire [4-1:0] node21860;
	wire [4-1:0] node21863;
	wire [4-1:0] node21864;
	wire [4-1:0] node21867;
	wire [4-1:0] node21870;
	wire [4-1:0] node21871;
	wire [4-1:0] node21873;
	wire [4-1:0] node21877;
	wire [4-1:0] node21878;
	wire [4-1:0] node21879;
	wire [4-1:0] node21881;
	wire [4-1:0] node21885;
	wire [4-1:0] node21888;
	wire [4-1:0] node21889;
	wire [4-1:0] node21890;
	wire [4-1:0] node21891;
	wire [4-1:0] node21892;
	wire [4-1:0] node21893;
	wire [4-1:0] node21894;
	wire [4-1:0] node21895;
	wire [4-1:0] node21896;
	wire [4-1:0] node21899;
	wire [4-1:0] node21902;
	wire [4-1:0] node21904;
	wire [4-1:0] node21905;
	wire [4-1:0] node21908;
	wire [4-1:0] node21911;
	wire [4-1:0] node21912;
	wire [4-1:0] node21913;
	wire [4-1:0] node21916;
	wire [4-1:0] node21919;
	wire [4-1:0] node21921;
	wire [4-1:0] node21923;
	wire [4-1:0] node21926;
	wire [4-1:0] node21927;
	wire [4-1:0] node21928;
	wire [4-1:0] node21929;
	wire [4-1:0] node21932;
	wire [4-1:0] node21933;
	wire [4-1:0] node21937;
	wire [4-1:0] node21938;
	wire [4-1:0] node21941;
	wire [4-1:0] node21944;
	wire [4-1:0] node21945;
	wire [4-1:0] node21947;
	wire [4-1:0] node21950;
	wire [4-1:0] node21951;
	wire [4-1:0] node21954;
	wire [4-1:0] node21957;
	wire [4-1:0] node21958;
	wire [4-1:0] node21959;
	wire [4-1:0] node21960;
	wire [4-1:0] node21962;
	wire [4-1:0] node21964;
	wire [4-1:0] node21967;
	wire [4-1:0] node21968;
	wire [4-1:0] node21971;
	wire [4-1:0] node21974;
	wire [4-1:0] node21975;
	wire [4-1:0] node21977;
	wire [4-1:0] node21980;
	wire [4-1:0] node21981;
	wire [4-1:0] node21984;
	wire [4-1:0] node21987;
	wire [4-1:0] node21988;
	wire [4-1:0] node21989;
	wire [4-1:0] node21991;
	wire [4-1:0] node21994;
	wire [4-1:0] node21995;
	wire [4-1:0] node21999;
	wire [4-1:0] node22000;
	wire [4-1:0] node22001;
	wire [4-1:0] node22006;
	wire [4-1:0] node22007;
	wire [4-1:0] node22008;
	wire [4-1:0] node22009;
	wire [4-1:0] node22010;
	wire [4-1:0] node22011;
	wire [4-1:0] node22014;
	wire [4-1:0] node22017;
	wire [4-1:0] node22018;
	wire [4-1:0] node22022;
	wire [4-1:0] node22023;
	wire [4-1:0] node22026;
	wire [4-1:0] node22029;
	wire [4-1:0] node22030;
	wire [4-1:0] node22031;
	wire [4-1:0] node22034;
	wire [4-1:0] node22037;
	wire [4-1:0] node22038;
	wire [4-1:0] node22041;
	wire [4-1:0] node22044;
	wire [4-1:0] node22045;
	wire [4-1:0] node22046;
	wire [4-1:0] node22047;
	wire [4-1:0] node22049;
	wire [4-1:0] node22051;
	wire [4-1:0] node22054;
	wire [4-1:0] node22055;
	wire [4-1:0] node22056;
	wire [4-1:0] node22060;
	wire [4-1:0] node22062;
	wire [4-1:0] node22065;
	wire [4-1:0] node22066;
	wire [4-1:0] node22067;
	wire [4-1:0] node22070;
	wire [4-1:0] node22071;
	wire [4-1:0] node22074;
	wire [4-1:0] node22077;
	wire [4-1:0] node22078;
	wire [4-1:0] node22080;
	wire [4-1:0] node22084;
	wire [4-1:0] node22085;
	wire [4-1:0] node22086;
	wire [4-1:0] node22087;
	wire [4-1:0] node22088;
	wire [4-1:0] node22092;
	wire [4-1:0] node22093;
	wire [4-1:0] node22096;
	wire [4-1:0] node22099;
	wire [4-1:0] node22101;
	wire [4-1:0] node22104;
	wire [4-1:0] node22105;
	wire [4-1:0] node22106;
	wire [4-1:0] node22110;
	wire [4-1:0] node22111;
	wire [4-1:0] node22114;
	wire [4-1:0] node22117;
	wire [4-1:0] node22118;
	wire [4-1:0] node22119;
	wire [4-1:0] node22120;
	wire [4-1:0] node22121;
	wire [4-1:0] node22122;
	wire [4-1:0] node22125;
	wire [4-1:0] node22128;
	wire [4-1:0] node22130;
	wire [4-1:0] node22131;
	wire [4-1:0] node22134;
	wire [4-1:0] node22137;
	wire [4-1:0] node22138;
	wire [4-1:0] node22139;
	wire [4-1:0] node22142;
	wire [4-1:0] node22145;
	wire [4-1:0] node22146;
	wire [4-1:0] node22147;
	wire [4-1:0] node22150;
	wire [4-1:0] node22153;
	wire [4-1:0] node22154;
	wire [4-1:0] node22157;
	wire [4-1:0] node22160;
	wire [4-1:0] node22161;
	wire [4-1:0] node22162;
	wire [4-1:0] node22163;
	wire [4-1:0] node22165;
	wire [4-1:0] node22168;
	wire [4-1:0] node22170;
	wire [4-1:0] node22173;
	wire [4-1:0] node22174;
	wire [4-1:0] node22176;
	wire [4-1:0] node22179;
	wire [4-1:0] node22182;
	wire [4-1:0] node22183;
	wire [4-1:0] node22184;
	wire [4-1:0] node22187;
	wire [4-1:0] node22189;
	wire [4-1:0] node22192;
	wire [4-1:0] node22193;
	wire [4-1:0] node22195;
	wire [4-1:0] node22198;
	wire [4-1:0] node22200;
	wire [4-1:0] node22203;
	wire [4-1:0] node22204;
	wire [4-1:0] node22205;
	wire [4-1:0] node22206;
	wire [4-1:0] node22207;
	wire [4-1:0] node22210;
	wire [4-1:0] node22213;
	wire [4-1:0] node22215;
	wire [4-1:0] node22216;
	wire [4-1:0] node22217;
	wire [4-1:0] node22220;
	wire [4-1:0] node22224;
	wire [4-1:0] node22225;
	wire [4-1:0] node22226;
	wire [4-1:0] node22227;
	wire [4-1:0] node22228;
	wire [4-1:0] node22231;
	wire [4-1:0] node22234;
	wire [4-1:0] node22236;
	wire [4-1:0] node22239;
	wire [4-1:0] node22241;
	wire [4-1:0] node22244;
	wire [4-1:0] node22246;
	wire [4-1:0] node22247;
	wire [4-1:0] node22250;
	wire [4-1:0] node22253;
	wire [4-1:0] node22254;
	wire [4-1:0] node22255;
	wire [4-1:0] node22256;
	wire [4-1:0] node22257;
	wire [4-1:0] node22259;
	wire [4-1:0] node22263;
	wire [4-1:0] node22264;
	wire [4-1:0] node22267;
	wire [4-1:0] node22270;
	wire [4-1:0] node22271;
	wire [4-1:0] node22272;
	wire [4-1:0] node22273;
	wire [4-1:0] node22278;
	wire [4-1:0] node22281;
	wire [4-1:0] node22282;
	wire [4-1:0] node22283;
	wire [4-1:0] node22286;
	wire [4-1:0] node22287;
	wire [4-1:0] node22290;
	wire [4-1:0] node22293;
	wire [4-1:0] node22295;
	wire [4-1:0] node22296;
	wire [4-1:0] node22297;
	wire [4-1:0] node22301;
	wire [4-1:0] node22304;
	wire [4-1:0] node22305;
	wire [4-1:0] node22306;
	wire [4-1:0] node22307;
	wire [4-1:0] node22308;
	wire [4-1:0] node22309;
	wire [4-1:0] node22310;
	wire [4-1:0] node22311;
	wire [4-1:0] node22315;
	wire [4-1:0] node22316;
	wire [4-1:0] node22318;
	wire [4-1:0] node22322;
	wire [4-1:0] node22323;
	wire [4-1:0] node22324;
	wire [4-1:0] node22328;
	wire [4-1:0] node22330;
	wire [4-1:0] node22333;
	wire [4-1:0] node22334;
	wire [4-1:0] node22335;
	wire [4-1:0] node22336;
	wire [4-1:0] node22337;
	wire [4-1:0] node22340;
	wire [4-1:0] node22343;
	wire [4-1:0] node22345;
	wire [4-1:0] node22348;
	wire [4-1:0] node22349;
	wire [4-1:0] node22352;
	wire [4-1:0] node22355;
	wire [4-1:0] node22356;
	wire [4-1:0] node22357;
	wire [4-1:0] node22360;
	wire [4-1:0] node22363;
	wire [4-1:0] node22364;
	wire [4-1:0] node22367;
	wire [4-1:0] node22370;
	wire [4-1:0] node22371;
	wire [4-1:0] node22372;
	wire [4-1:0] node22374;
	wire [4-1:0] node22376;
	wire [4-1:0] node22379;
	wire [4-1:0] node22380;
	wire [4-1:0] node22383;
	wire [4-1:0] node22386;
	wire [4-1:0] node22387;
	wire [4-1:0] node22388;
	wire [4-1:0] node22391;
	wire [4-1:0] node22394;
	wire [4-1:0] node22395;
	wire [4-1:0] node22397;
	wire [4-1:0] node22400;
	wire [4-1:0] node22401;
	wire [4-1:0] node22404;
	wire [4-1:0] node22407;
	wire [4-1:0] node22408;
	wire [4-1:0] node22409;
	wire [4-1:0] node22410;
	wire [4-1:0] node22411;
	wire [4-1:0] node22412;
	wire [4-1:0] node22413;
	wire [4-1:0] node22416;
	wire [4-1:0] node22419;
	wire [4-1:0] node22420;
	wire [4-1:0] node22425;
	wire [4-1:0] node22426;
	wire [4-1:0] node22427;
	wire [4-1:0] node22430;
	wire [4-1:0] node22433;
	wire [4-1:0] node22436;
	wire [4-1:0] node22437;
	wire [4-1:0] node22438;
	wire [4-1:0] node22439;
	wire [4-1:0] node22440;
	wire [4-1:0] node22444;
	wire [4-1:0] node22447;
	wire [4-1:0] node22449;
	wire [4-1:0] node22452;
	wire [4-1:0] node22453;
	wire [4-1:0] node22454;
	wire [4-1:0] node22456;
	wire [4-1:0] node22459;
	wire [4-1:0] node22460;
	wire [4-1:0] node22464;
	wire [4-1:0] node22467;
	wire [4-1:0] node22468;
	wire [4-1:0] node22469;
	wire [4-1:0] node22470;
	wire [4-1:0] node22472;
	wire [4-1:0] node22475;
	wire [4-1:0] node22477;
	wire [4-1:0] node22480;
	wire [4-1:0] node22481;
	wire [4-1:0] node22482;
	wire [4-1:0] node22485;
	wire [4-1:0] node22488;
	wire [4-1:0] node22490;
	wire [4-1:0] node22491;
	wire [4-1:0] node22495;
	wire [4-1:0] node22496;
	wire [4-1:0] node22497;
	wire [4-1:0] node22498;
	wire [4-1:0] node22499;
	wire [4-1:0] node22502;
	wire [4-1:0] node22505;
	wire [4-1:0] node22506;
	wire [4-1:0] node22510;
	wire [4-1:0] node22512;
	wire [4-1:0] node22513;
	wire [4-1:0] node22516;
	wire [4-1:0] node22519;
	wire [4-1:0] node22520;
	wire [4-1:0] node22521;
	wire [4-1:0] node22523;
	wire [4-1:0] node22526;
	wire [4-1:0] node22527;
	wire [4-1:0] node22530;
	wire [4-1:0] node22533;
	wire [4-1:0] node22534;
	wire [4-1:0] node22536;
	wire [4-1:0] node22539;
	wire [4-1:0] node22541;
	wire [4-1:0] node22544;
	wire [4-1:0] node22545;
	wire [4-1:0] node22546;
	wire [4-1:0] node22547;
	wire [4-1:0] node22548;
	wire [4-1:0] node22549;
	wire [4-1:0] node22550;
	wire [4-1:0] node22551;
	wire [4-1:0] node22554;
	wire [4-1:0] node22558;
	wire [4-1:0] node22560;
	wire [4-1:0] node22561;
	wire [4-1:0] node22564;
	wire [4-1:0] node22567;
	wire [4-1:0] node22568;
	wire [4-1:0] node22570;
	wire [4-1:0] node22571;
	wire [4-1:0] node22575;
	wire [4-1:0] node22578;
	wire [4-1:0] node22579;
	wire [4-1:0] node22580;
	wire [4-1:0] node22581;
	wire [4-1:0] node22584;
	wire [4-1:0] node22587;
	wire [4-1:0] node22590;
	wire [4-1:0] node22592;
	wire [4-1:0] node22593;
	wire [4-1:0] node22596;
	wire [4-1:0] node22599;
	wire [4-1:0] node22600;
	wire [4-1:0] node22601;
	wire [4-1:0] node22602;
	wire [4-1:0] node22603;
	wire [4-1:0] node22604;
	wire [4-1:0] node22608;
	wire [4-1:0] node22609;
	wire [4-1:0] node22613;
	wire [4-1:0] node22614;
	wire [4-1:0] node22615;
	wire [4-1:0] node22619;
	wire [4-1:0] node22621;
	wire [4-1:0] node22624;
	wire [4-1:0] node22625;
	wire [4-1:0] node22627;
	wire [4-1:0] node22630;
	wire [4-1:0] node22631;
	wire [4-1:0] node22635;
	wire [4-1:0] node22636;
	wire [4-1:0] node22637;
	wire [4-1:0] node22640;
	wire [4-1:0] node22643;
	wire [4-1:0] node22644;
	wire [4-1:0] node22645;
	wire [4-1:0] node22647;
	wire [4-1:0] node22650;
	wire [4-1:0] node22651;
	wire [4-1:0] node22654;
	wire [4-1:0] node22657;
	wire [4-1:0] node22658;
	wire [4-1:0] node22662;
	wire [4-1:0] node22663;
	wire [4-1:0] node22664;
	wire [4-1:0] node22665;
	wire [4-1:0] node22666;
	wire [4-1:0] node22668;
	wire [4-1:0] node22671;
	wire [4-1:0] node22672;
	wire [4-1:0] node22673;
	wire [4-1:0] node22676;
	wire [4-1:0] node22679;
	wire [4-1:0] node22681;
	wire [4-1:0] node22684;
	wire [4-1:0] node22686;
	wire [4-1:0] node22687;
	wire [4-1:0] node22689;
	wire [4-1:0] node22692;
	wire [4-1:0] node22693;
	wire [4-1:0] node22697;
	wire [4-1:0] node22698;
	wire [4-1:0] node22699;
	wire [4-1:0] node22700;
	wire [4-1:0] node22703;
	wire [4-1:0] node22706;
	wire [4-1:0] node22708;
	wire [4-1:0] node22711;
	wire [4-1:0] node22712;
	wire [4-1:0] node22713;
	wire [4-1:0] node22716;
	wire [4-1:0] node22719;
	wire [4-1:0] node22721;
	wire [4-1:0] node22723;
	wire [4-1:0] node22726;
	wire [4-1:0] node22727;
	wire [4-1:0] node22728;
	wire [4-1:0] node22729;
	wire [4-1:0] node22730;
	wire [4-1:0] node22731;
	wire [4-1:0] node22734;
	wire [4-1:0] node22738;
	wire [4-1:0] node22739;
	wire [4-1:0] node22742;
	wire [4-1:0] node22745;
	wire [4-1:0] node22746;
	wire [4-1:0] node22748;
	wire [4-1:0] node22751;
	wire [4-1:0] node22753;
	wire [4-1:0] node22754;
	wire [4-1:0] node22757;
	wire [4-1:0] node22760;
	wire [4-1:0] node22761;
	wire [4-1:0] node22762;
	wire [4-1:0] node22763;
	wire [4-1:0] node22766;
	wire [4-1:0] node22769;
	wire [4-1:0] node22770;
	wire [4-1:0] node22772;
	wire [4-1:0] node22775;
	wire [4-1:0] node22776;
	wire [4-1:0] node22779;
	wire [4-1:0] node22782;
	wire [4-1:0] node22784;
	wire [4-1:0] node22785;
	wire [4-1:0] node22786;
	wire [4-1:0] node22790;
	wire [4-1:0] node22791;
	wire [4-1:0] node22794;
	wire [4-1:0] node22797;
	wire [4-1:0] node22798;
	wire [4-1:0] node22799;
	wire [4-1:0] node22800;
	wire [4-1:0] node22801;
	wire [4-1:0] node22802;
	wire [4-1:0] node22803;
	wire [4-1:0] node22804;
	wire [4-1:0] node22805;
	wire [4-1:0] node22806;
	wire [4-1:0] node22807;
	wire [4-1:0] node22808;
	wire [4-1:0] node22809;
	wire [4-1:0] node22812;
	wire [4-1:0] node22815;
	wire [4-1:0] node22816;
	wire [4-1:0] node22820;
	wire [4-1:0] node22821;
	wire [4-1:0] node22823;
	wire [4-1:0] node22827;
	wire [4-1:0] node22828;
	wire [4-1:0] node22829;
	wire [4-1:0] node22830;
	wire [4-1:0] node22833;
	wire [4-1:0] node22837;
	wire [4-1:0] node22838;
	wire [4-1:0] node22841;
	wire [4-1:0] node22844;
	wire [4-1:0] node22845;
	wire [4-1:0] node22846;
	wire [4-1:0] node22847;
	wire [4-1:0] node22850;
	wire [4-1:0] node22851;
	wire [4-1:0] node22854;
	wire [4-1:0] node22857;
	wire [4-1:0] node22859;
	wire [4-1:0] node22861;
	wire [4-1:0] node22864;
	wire [4-1:0] node22865;
	wire [4-1:0] node22867;
	wire [4-1:0] node22868;
	wire [4-1:0] node22871;
	wire [4-1:0] node22874;
	wire [4-1:0] node22876;
	wire [4-1:0] node22877;
	wire [4-1:0] node22881;
	wire [4-1:0] node22882;
	wire [4-1:0] node22883;
	wire [4-1:0] node22884;
	wire [4-1:0] node22886;
	wire [4-1:0] node22887;
	wire [4-1:0] node22890;
	wire [4-1:0] node22893;
	wire [4-1:0] node22894;
	wire [4-1:0] node22895;
	wire [4-1:0] node22898;
	wire [4-1:0] node22902;
	wire [4-1:0] node22903;
	wire [4-1:0] node22904;
	wire [4-1:0] node22905;
	wire [4-1:0] node22908;
	wire [4-1:0] node22911;
	wire [4-1:0] node22912;
	wire [4-1:0] node22915;
	wire [4-1:0] node22918;
	wire [4-1:0] node22920;
	wire [4-1:0] node22921;
	wire [4-1:0] node22925;
	wire [4-1:0] node22926;
	wire [4-1:0] node22927;
	wire [4-1:0] node22928;
	wire [4-1:0] node22929;
	wire [4-1:0] node22933;
	wire [4-1:0] node22934;
	wire [4-1:0] node22938;
	wire [4-1:0] node22941;
	wire [4-1:0] node22942;
	wire [4-1:0] node22944;
	wire [4-1:0] node22945;
	wire [4-1:0] node22948;
	wire [4-1:0] node22951;
	wire [4-1:0] node22952;
	wire [4-1:0] node22955;
	wire [4-1:0] node22956;
	wire [4-1:0] node22959;
	wire [4-1:0] node22962;
	wire [4-1:0] node22963;
	wire [4-1:0] node22964;
	wire [4-1:0] node22965;
	wire [4-1:0] node22966;
	wire [4-1:0] node22968;
	wire [4-1:0] node22970;
	wire [4-1:0] node22973;
	wire [4-1:0] node22974;
	wire [4-1:0] node22976;
	wire [4-1:0] node22979;
	wire [4-1:0] node22980;
	wire [4-1:0] node22984;
	wire [4-1:0] node22985;
	wire [4-1:0] node22987;
	wire [4-1:0] node22988;
	wire [4-1:0] node22991;
	wire [4-1:0] node22994;
	wire [4-1:0] node22995;
	wire [4-1:0] node22996;
	wire [4-1:0] node22999;
	wire [4-1:0] node23002;
	wire [4-1:0] node23004;
	wire [4-1:0] node23007;
	wire [4-1:0] node23008;
	wire [4-1:0] node23009;
	wire [4-1:0] node23011;
	wire [4-1:0] node23012;
	wire [4-1:0] node23015;
	wire [4-1:0] node23018;
	wire [4-1:0] node23019;
	wire [4-1:0] node23020;
	wire [4-1:0] node23023;
	wire [4-1:0] node23026;
	wire [4-1:0] node23027;
	wire [4-1:0] node23030;
	wire [4-1:0] node23033;
	wire [4-1:0] node23034;
	wire [4-1:0] node23035;
	wire [4-1:0] node23037;
	wire [4-1:0] node23040;
	wire [4-1:0] node23041;
	wire [4-1:0] node23044;
	wire [4-1:0] node23047;
	wire [4-1:0] node23048;
	wire [4-1:0] node23049;
	wire [4-1:0] node23052;
	wire [4-1:0] node23055;
	wire [4-1:0] node23058;
	wire [4-1:0] node23059;
	wire [4-1:0] node23060;
	wire [4-1:0] node23061;
	wire [4-1:0] node23064;
	wire [4-1:0] node23065;
	wire [4-1:0] node23066;
	wire [4-1:0] node23071;
	wire [4-1:0] node23072;
	wire [4-1:0] node23073;
	wire [4-1:0] node23076;
	wire [4-1:0] node23077;
	wire [4-1:0] node23080;
	wire [4-1:0] node23083;
	wire [4-1:0] node23084;
	wire [4-1:0] node23087;
	wire [4-1:0] node23088;
	wire [4-1:0] node23092;
	wire [4-1:0] node23093;
	wire [4-1:0] node23094;
	wire [4-1:0] node23095;
	wire [4-1:0] node23096;
	wire [4-1:0] node23099;
	wire [4-1:0] node23102;
	wire [4-1:0] node23104;
	wire [4-1:0] node23107;
	wire [4-1:0] node23109;
	wire [4-1:0] node23112;
	wire [4-1:0] node23113;
	wire [4-1:0] node23114;
	wire [4-1:0] node23116;
	wire [4-1:0] node23119;
	wire [4-1:0] node23120;
	wire [4-1:0] node23124;
	wire [4-1:0] node23127;
	wire [4-1:0] node23128;
	wire [4-1:0] node23129;
	wire [4-1:0] node23130;
	wire [4-1:0] node23131;
	wire [4-1:0] node23132;
	wire [4-1:0] node23133;
	wire [4-1:0] node23135;
	wire [4-1:0] node23138;
	wire [4-1:0] node23139;
	wire [4-1:0] node23143;
	wire [4-1:0] node23144;
	wire [4-1:0] node23145;
	wire [4-1:0] node23149;
	wire [4-1:0] node23151;
	wire [4-1:0] node23154;
	wire [4-1:0] node23155;
	wire [4-1:0] node23156;
	wire [4-1:0] node23158;
	wire [4-1:0] node23161;
	wire [4-1:0] node23162;
	wire [4-1:0] node23166;
	wire [4-1:0] node23167;
	wire [4-1:0] node23169;
	wire [4-1:0] node23172;
	wire [4-1:0] node23173;
	wire [4-1:0] node23177;
	wire [4-1:0] node23178;
	wire [4-1:0] node23179;
	wire [4-1:0] node23180;
	wire [4-1:0] node23184;
	wire [4-1:0] node23186;
	wire [4-1:0] node23188;
	wire [4-1:0] node23191;
	wire [4-1:0] node23192;
	wire [4-1:0] node23194;
	wire [4-1:0] node23195;
	wire [4-1:0] node23199;
	wire [4-1:0] node23200;
	wire [4-1:0] node23201;
	wire [4-1:0] node23204;
	wire [4-1:0] node23207;
	wire [4-1:0] node23210;
	wire [4-1:0] node23211;
	wire [4-1:0] node23212;
	wire [4-1:0] node23213;
	wire [4-1:0] node23215;
	wire [4-1:0] node23217;
	wire [4-1:0] node23220;
	wire [4-1:0] node23221;
	wire [4-1:0] node23222;
	wire [4-1:0] node23225;
	wire [4-1:0] node23228;
	wire [4-1:0] node23231;
	wire [4-1:0] node23232;
	wire [4-1:0] node23234;
	wire [4-1:0] node23237;
	wire [4-1:0] node23238;
	wire [4-1:0] node23239;
	wire [4-1:0] node23243;
	wire [4-1:0] node23244;
	wire [4-1:0] node23247;
	wire [4-1:0] node23250;
	wire [4-1:0] node23251;
	wire [4-1:0] node23252;
	wire [4-1:0] node23253;
	wire [4-1:0] node23254;
	wire [4-1:0] node23257;
	wire [4-1:0] node23261;
	wire [4-1:0] node23263;
	wire [4-1:0] node23265;
	wire [4-1:0] node23268;
	wire [4-1:0] node23269;
	wire [4-1:0] node23270;
	wire [4-1:0] node23271;
	wire [4-1:0] node23275;
	wire [4-1:0] node23276;
	wire [4-1:0] node23279;
	wire [4-1:0] node23282;
	wire [4-1:0] node23283;
	wire [4-1:0] node23286;
	wire [4-1:0] node23289;
	wire [4-1:0] node23290;
	wire [4-1:0] node23291;
	wire [4-1:0] node23292;
	wire [4-1:0] node23293;
	wire [4-1:0] node23294;
	wire [4-1:0] node23295;
	wire [4-1:0] node23298;
	wire [4-1:0] node23302;
	wire [4-1:0] node23303;
	wire [4-1:0] node23304;
	wire [4-1:0] node23307;
	wire [4-1:0] node23310;
	wire [4-1:0] node23312;
	wire [4-1:0] node23315;
	wire [4-1:0] node23316;
	wire [4-1:0] node23317;
	wire [4-1:0] node23321;
	wire [4-1:0] node23322;
	wire [4-1:0] node23323;
	wire [4-1:0] node23326;
	wire [4-1:0] node23329;
	wire [4-1:0] node23330;
	wire [4-1:0] node23334;
	wire [4-1:0] node23335;
	wire [4-1:0] node23336;
	wire [4-1:0] node23338;
	wire [4-1:0] node23339;
	wire [4-1:0] node23343;
	wire [4-1:0] node23344;
	wire [4-1:0] node23347;
	wire [4-1:0] node23349;
	wire [4-1:0] node23352;
	wire [4-1:0] node23353;
	wire [4-1:0] node23354;
	wire [4-1:0] node23355;
	wire [4-1:0] node23358;
	wire [4-1:0] node23361;
	wire [4-1:0] node23364;
	wire [4-1:0] node23365;
	wire [4-1:0] node23366;
	wire [4-1:0] node23369;
	wire [4-1:0] node23372;
	wire [4-1:0] node23374;
	wire [4-1:0] node23377;
	wire [4-1:0] node23378;
	wire [4-1:0] node23379;
	wire [4-1:0] node23380;
	wire [4-1:0] node23381;
	wire [4-1:0] node23382;
	wire [4-1:0] node23385;
	wire [4-1:0] node23388;
	wire [4-1:0] node23389;
	wire [4-1:0] node23393;
	wire [4-1:0] node23394;
	wire [4-1:0] node23397;
	wire [4-1:0] node23398;
	wire [4-1:0] node23401;
	wire [4-1:0] node23404;
	wire [4-1:0] node23405;
	wire [4-1:0] node23407;
	wire [4-1:0] node23408;
	wire [4-1:0] node23412;
	wire [4-1:0] node23413;
	wire [4-1:0] node23416;
	wire [4-1:0] node23418;
	wire [4-1:0] node23421;
	wire [4-1:0] node23422;
	wire [4-1:0] node23423;
	wire [4-1:0] node23424;
	wire [4-1:0] node23425;
	wire [4-1:0] node23429;
	wire [4-1:0] node23430;
	wire [4-1:0] node23433;
	wire [4-1:0] node23436;
	wire [4-1:0] node23437;
	wire [4-1:0] node23438;
	wire [4-1:0] node23442;
	wire [4-1:0] node23444;
	wire [4-1:0] node23447;
	wire [4-1:0] node23448;
	wire [4-1:0] node23450;
	wire [4-1:0] node23452;
	wire [4-1:0] node23455;
	wire [4-1:0] node23456;
	wire [4-1:0] node23458;
	wire [4-1:0] node23462;
	wire [4-1:0] node23463;
	wire [4-1:0] node23464;
	wire [4-1:0] node23465;
	wire [4-1:0] node23466;
	wire [4-1:0] node23467;
	wire [4-1:0] node23468;
	wire [4-1:0] node23469;
	wire [4-1:0] node23472;
	wire [4-1:0] node23475;
	wire [4-1:0] node23476;
	wire [4-1:0] node23479;
	wire [4-1:0] node23482;
	wire [4-1:0] node23483;
	wire [4-1:0] node23484;
	wire [4-1:0] node23488;
	wire [4-1:0] node23489;
	wire [4-1:0] node23492;
	wire [4-1:0] node23495;
	wire [4-1:0] node23496;
	wire [4-1:0] node23497;
	wire [4-1:0] node23498;
	wire [4-1:0] node23502;
	wire [4-1:0] node23503;
	wire [4-1:0] node23507;
	wire [4-1:0] node23508;
	wire [4-1:0] node23509;
	wire [4-1:0] node23512;
	wire [4-1:0] node23515;
	wire [4-1:0] node23517;
	wire [4-1:0] node23520;
	wire [4-1:0] node23521;
	wire [4-1:0] node23522;
	wire [4-1:0] node23523;
	wire [4-1:0] node23524;
	wire [4-1:0] node23527;
	wire [4-1:0] node23530;
	wire [4-1:0] node23531;
	wire [4-1:0] node23532;
	wire [4-1:0] node23536;
	wire [4-1:0] node23537;
	wire [4-1:0] node23541;
	wire [4-1:0] node23542;
	wire [4-1:0] node23543;
	wire [4-1:0] node23546;
	wire [4-1:0] node23549;
	wire [4-1:0] node23550;
	wire [4-1:0] node23551;
	wire [4-1:0] node23554;
	wire [4-1:0] node23557;
	wire [4-1:0] node23558;
	wire [4-1:0] node23562;
	wire [4-1:0] node23563;
	wire [4-1:0] node23564;
	wire [4-1:0] node23566;
	wire [4-1:0] node23567;
	wire [4-1:0] node23571;
	wire [4-1:0] node23572;
	wire [4-1:0] node23573;
	wire [4-1:0] node23577;
	wire [4-1:0] node23578;
	wire [4-1:0] node23582;
	wire [4-1:0] node23583;
	wire [4-1:0] node23584;
	wire [4-1:0] node23585;
	wire [4-1:0] node23588;
	wire [4-1:0] node23591;
	wire [4-1:0] node23593;
	wire [4-1:0] node23596;
	wire [4-1:0] node23597;
	wire [4-1:0] node23600;
	wire [4-1:0] node23603;
	wire [4-1:0] node23604;
	wire [4-1:0] node23605;
	wire [4-1:0] node23606;
	wire [4-1:0] node23609;
	wire [4-1:0] node23610;
	wire [4-1:0] node23611;
	wire [4-1:0] node23614;
	wire [4-1:0] node23617;
	wire [4-1:0] node23618;
	wire [4-1:0] node23621;
	wire [4-1:0] node23624;
	wire [4-1:0] node23625;
	wire [4-1:0] node23626;
	wire [4-1:0] node23628;
	wire [4-1:0] node23631;
	wire [4-1:0] node23632;
	wire [4-1:0] node23636;
	wire [4-1:0] node23637;
	wire [4-1:0] node23639;
	wire [4-1:0] node23642;
	wire [4-1:0] node23643;
	wire [4-1:0] node23644;
	wire [4-1:0] node23649;
	wire [4-1:0] node23650;
	wire [4-1:0] node23651;
	wire [4-1:0] node23652;
	wire [4-1:0] node23653;
	wire [4-1:0] node23656;
	wire [4-1:0] node23659;
	wire [4-1:0] node23661;
	wire [4-1:0] node23664;
	wire [4-1:0] node23665;
	wire [4-1:0] node23666;
	wire [4-1:0] node23669;
	wire [4-1:0] node23672;
	wire [4-1:0] node23675;
	wire [4-1:0] node23676;
	wire [4-1:0] node23677;
	wire [4-1:0] node23678;
	wire [4-1:0] node23681;
	wire [4-1:0] node23684;
	wire [4-1:0] node23685;
	wire [4-1:0] node23686;
	wire [4-1:0] node23691;
	wire [4-1:0] node23692;
	wire [4-1:0] node23693;
	wire [4-1:0] node23695;
	wire [4-1:0] node23698;
	wire [4-1:0] node23701;
	wire [4-1:0] node23703;
	wire [4-1:0] node23706;
	wire [4-1:0] node23707;
	wire [4-1:0] node23708;
	wire [4-1:0] node23709;
	wire [4-1:0] node23710;
	wire [4-1:0] node23711;
	wire [4-1:0] node23712;
	wire [4-1:0] node23713;
	wire [4-1:0] node23717;
	wire [4-1:0] node23718;
	wire [4-1:0] node23722;
	wire [4-1:0] node23723;
	wire [4-1:0] node23725;
	wire [4-1:0] node23728;
	wire [4-1:0] node23731;
	wire [4-1:0] node23732;
	wire [4-1:0] node23733;
	wire [4-1:0] node23735;
	wire [4-1:0] node23739;
	wire [4-1:0] node23740;
	wire [4-1:0] node23742;
	wire [4-1:0] node23746;
	wire [4-1:0] node23747;
	wire [4-1:0] node23748;
	wire [4-1:0] node23749;
	wire [4-1:0] node23751;
	wire [4-1:0] node23754;
	wire [4-1:0] node23755;
	wire [4-1:0] node23758;
	wire [4-1:0] node23761;
	wire [4-1:0] node23762;
	wire [4-1:0] node23764;
	wire [4-1:0] node23767;
	wire [4-1:0] node23768;
	wire [4-1:0] node23771;
	wire [4-1:0] node23774;
	wire [4-1:0] node23775;
	wire [4-1:0] node23776;
	wire [4-1:0] node23777;
	wire [4-1:0] node23780;
	wire [4-1:0] node23783;
	wire [4-1:0] node23784;
	wire [4-1:0] node23787;
	wire [4-1:0] node23790;
	wire [4-1:0] node23791;
	wire [4-1:0] node23792;
	wire [4-1:0] node23797;
	wire [4-1:0] node23798;
	wire [4-1:0] node23799;
	wire [4-1:0] node23800;
	wire [4-1:0] node23802;
	wire [4-1:0] node23805;
	wire [4-1:0] node23806;
	wire [4-1:0] node23809;
	wire [4-1:0] node23812;
	wire [4-1:0] node23813;
	wire [4-1:0] node23814;
	wire [4-1:0] node23815;
	wire [4-1:0] node23819;
	wire [4-1:0] node23821;
	wire [4-1:0] node23824;
	wire [4-1:0] node23826;
	wire [4-1:0] node23829;
	wire [4-1:0] node23830;
	wire [4-1:0] node23831;
	wire [4-1:0] node23832;
	wire [4-1:0] node23834;
	wire [4-1:0] node23838;
	wire [4-1:0] node23840;
	wire [4-1:0] node23843;
	wire [4-1:0] node23844;
	wire [4-1:0] node23845;
	wire [4-1:0] node23846;
	wire [4-1:0] node23849;
	wire [4-1:0] node23853;
	wire [4-1:0] node23854;
	wire [4-1:0] node23857;
	wire [4-1:0] node23860;
	wire [4-1:0] node23861;
	wire [4-1:0] node23862;
	wire [4-1:0] node23863;
	wire [4-1:0] node23864;
	wire [4-1:0] node23865;
	wire [4-1:0] node23867;
	wire [4-1:0] node23870;
	wire [4-1:0] node23871;
	wire [4-1:0] node23875;
	wire [4-1:0] node23876;
	wire [4-1:0] node23880;
	wire [4-1:0] node23881;
	wire [4-1:0] node23882;
	wire [4-1:0] node23883;
	wire [4-1:0] node23887;
	wire [4-1:0] node23888;
	wire [4-1:0] node23892;
	wire [4-1:0] node23894;
	wire [4-1:0] node23897;
	wire [4-1:0] node23898;
	wire [4-1:0] node23899;
	wire [4-1:0] node23900;
	wire [4-1:0] node23903;
	wire [4-1:0] node23906;
	wire [4-1:0] node23907;
	wire [4-1:0] node23909;
	wire [4-1:0] node23913;
	wire [4-1:0] node23914;
	wire [4-1:0] node23915;
	wire [4-1:0] node23918;
	wire [4-1:0] node23921;
	wire [4-1:0] node23923;
	wire [4-1:0] node23925;
	wire [4-1:0] node23928;
	wire [4-1:0] node23929;
	wire [4-1:0] node23930;
	wire [4-1:0] node23931;
	wire [4-1:0] node23932;
	wire [4-1:0] node23933;
	wire [4-1:0] node23936;
	wire [4-1:0] node23940;
	wire [4-1:0] node23941;
	wire [4-1:0] node23944;
	wire [4-1:0] node23947;
	wire [4-1:0] node23948;
	wire [4-1:0] node23949;
	wire [4-1:0] node23952;
	wire [4-1:0] node23955;
	wire [4-1:0] node23956;
	wire [4-1:0] node23959;
	wire [4-1:0] node23962;
	wire [4-1:0] node23963;
	wire [4-1:0] node23964;
	wire [4-1:0] node23966;
	wire [4-1:0] node23969;
	wire [4-1:0] node23971;
	wire [4-1:0] node23974;
	wire [4-1:0] node23975;
	wire [4-1:0] node23978;
	wire [4-1:0] node23979;
	wire [4-1:0] node23981;
	wire [4-1:0] node23985;
	wire [4-1:0] node23986;
	wire [4-1:0] node23987;
	wire [4-1:0] node23988;
	wire [4-1:0] node23989;
	wire [4-1:0] node23990;
	wire [4-1:0] node23991;
	wire [4-1:0] node23992;
	wire [4-1:0] node23993;
	wire [4-1:0] node23994;
	wire [4-1:0] node23997;
	wire [4-1:0] node24001;
	wire [4-1:0] node24002;
	wire [4-1:0] node24005;
	wire [4-1:0] node24008;
	wire [4-1:0] node24009;
	wire [4-1:0] node24011;
	wire [4-1:0] node24012;
	wire [4-1:0] node24015;
	wire [4-1:0] node24018;
	wire [4-1:0] node24019;
	wire [4-1:0] node24020;
	wire [4-1:0] node24024;
	wire [4-1:0] node24027;
	wire [4-1:0] node24028;
	wire [4-1:0] node24029;
	wire [4-1:0] node24031;
	wire [4-1:0] node24034;
	wire [4-1:0] node24036;
	wire [4-1:0] node24039;
	wire [4-1:0] node24041;
	wire [4-1:0] node24042;
	wire [4-1:0] node24043;
	wire [4-1:0] node24047;
	wire [4-1:0] node24050;
	wire [4-1:0] node24051;
	wire [4-1:0] node24052;
	wire [4-1:0] node24053;
	wire [4-1:0] node24054;
	wire [4-1:0] node24058;
	wire [4-1:0] node24059;
	wire [4-1:0] node24060;
	wire [4-1:0] node24063;
	wire [4-1:0] node24067;
	wire [4-1:0] node24068;
	wire [4-1:0] node24069;
	wire [4-1:0] node24070;
	wire [4-1:0] node24073;
	wire [4-1:0] node24077;
	wire [4-1:0] node24079;
	wire [4-1:0] node24080;
	wire [4-1:0] node24083;
	wire [4-1:0] node24086;
	wire [4-1:0] node24087;
	wire [4-1:0] node24088;
	wire [4-1:0] node24090;
	wire [4-1:0] node24091;
	wire [4-1:0] node24095;
	wire [4-1:0] node24097;
	wire [4-1:0] node24100;
	wire [4-1:0] node24101;
	wire [4-1:0] node24103;
	wire [4-1:0] node24106;
	wire [4-1:0] node24107;
	wire [4-1:0] node24110;
	wire [4-1:0] node24113;
	wire [4-1:0] node24114;
	wire [4-1:0] node24115;
	wire [4-1:0] node24116;
	wire [4-1:0] node24117;
	wire [4-1:0] node24119;
	wire [4-1:0] node24121;
	wire [4-1:0] node24124;
	wire [4-1:0] node24125;
	wire [4-1:0] node24127;
	wire [4-1:0] node24130;
	wire [4-1:0] node24131;
	wire [4-1:0] node24135;
	wire [4-1:0] node24136;
	wire [4-1:0] node24137;
	wire [4-1:0] node24138;
	wire [4-1:0] node24143;
	wire [4-1:0] node24144;
	wire [4-1:0] node24147;
	wire [4-1:0] node24150;
	wire [4-1:0] node24151;
	wire [4-1:0] node24152;
	wire [4-1:0] node24153;
	wire [4-1:0] node24154;
	wire [4-1:0] node24157;
	wire [4-1:0] node24160;
	wire [4-1:0] node24163;
	wire [4-1:0] node24164;
	wire [4-1:0] node24167;
	wire [4-1:0] node24170;
	wire [4-1:0] node24171;
	wire [4-1:0] node24172;
	wire [4-1:0] node24173;
	wire [4-1:0] node24178;
	wire [4-1:0] node24179;
	wire [4-1:0] node24182;
	wire [4-1:0] node24185;
	wire [4-1:0] node24186;
	wire [4-1:0] node24187;
	wire [4-1:0] node24188;
	wire [4-1:0] node24189;
	wire [4-1:0] node24190;
	wire [4-1:0] node24194;
	wire [4-1:0] node24196;
	wire [4-1:0] node24199;
	wire [4-1:0] node24201;
	wire [4-1:0] node24202;
	wire [4-1:0] node24206;
	wire [4-1:0] node24207;
	wire [4-1:0] node24208;
	wire [4-1:0] node24209;
	wire [4-1:0] node24212;
	wire [4-1:0] node24215;
	wire [4-1:0] node24218;
	wire [4-1:0] node24219;
	wire [4-1:0] node24221;
	wire [4-1:0] node24224;
	wire [4-1:0] node24225;
	wire [4-1:0] node24229;
	wire [4-1:0] node24230;
	wire [4-1:0] node24231;
	wire [4-1:0] node24233;
	wire [4-1:0] node24236;
	wire [4-1:0] node24238;
	wire [4-1:0] node24241;
	wire [4-1:0] node24242;
	wire [4-1:0] node24243;
	wire [4-1:0] node24244;
	wire [4-1:0] node24247;
	wire [4-1:0] node24251;
	wire [4-1:0] node24253;
	wire [4-1:0] node24254;
	wire [4-1:0] node24258;
	wire [4-1:0] node24259;
	wire [4-1:0] node24260;
	wire [4-1:0] node24261;
	wire [4-1:0] node24262;
	wire [4-1:0] node24264;
	wire [4-1:0] node24266;
	wire [4-1:0] node24269;
	wire [4-1:0] node24270;
	wire [4-1:0] node24271;
	wire [4-1:0] node24272;
	wire [4-1:0] node24275;
	wire [4-1:0] node24278;
	wire [4-1:0] node24279;
	wire [4-1:0] node24282;
	wire [4-1:0] node24286;
	wire [4-1:0] node24287;
	wire [4-1:0] node24288;
	wire [4-1:0] node24290;
	wire [4-1:0] node24292;
	wire [4-1:0] node24295;
	wire [4-1:0] node24296;
	wire [4-1:0] node24299;
	wire [4-1:0] node24302;
	wire [4-1:0] node24303;
	wire [4-1:0] node24304;
	wire [4-1:0] node24305;
	wire [4-1:0] node24310;
	wire [4-1:0] node24311;
	wire [4-1:0] node24312;
	wire [4-1:0] node24316;
	wire [4-1:0] node24317;
	wire [4-1:0] node24321;
	wire [4-1:0] node24322;
	wire [4-1:0] node24323;
	wire [4-1:0] node24324;
	wire [4-1:0] node24326;
	wire [4-1:0] node24329;
	wire [4-1:0] node24330;
	wire [4-1:0] node24333;
	wire [4-1:0] node24336;
	wire [4-1:0] node24337;
	wire [4-1:0] node24338;
	wire [4-1:0] node24339;
	wire [4-1:0] node24344;
	wire [4-1:0] node24345;
	wire [4-1:0] node24349;
	wire [4-1:0] node24350;
	wire [4-1:0] node24351;
	wire [4-1:0] node24353;
	wire [4-1:0] node24356;
	wire [4-1:0] node24357;
	wire [4-1:0] node24358;
	wire [4-1:0] node24363;
	wire [4-1:0] node24364;
	wire [4-1:0] node24365;
	wire [4-1:0] node24367;
	wire [4-1:0] node24371;
	wire [4-1:0] node24372;
	wire [4-1:0] node24376;
	wire [4-1:0] node24377;
	wire [4-1:0] node24378;
	wire [4-1:0] node24379;
	wire [4-1:0] node24380;
	wire [4-1:0] node24381;
	wire [4-1:0] node24383;
	wire [4-1:0] node24386;
	wire [4-1:0] node24389;
	wire [4-1:0] node24390;
	wire [4-1:0] node24391;
	wire [4-1:0] node24394;
	wire [4-1:0] node24398;
	wire [4-1:0] node24399;
	wire [4-1:0] node24400;
	wire [4-1:0] node24403;
	wire [4-1:0] node24405;
	wire [4-1:0] node24408;
	wire [4-1:0] node24409;
	wire [4-1:0] node24411;
	wire [4-1:0] node24415;
	wire [4-1:0] node24416;
	wire [4-1:0] node24417;
	wire [4-1:0] node24418;
	wire [4-1:0] node24419;
	wire [4-1:0] node24424;
	wire [4-1:0] node24425;
	wire [4-1:0] node24426;
	wire [4-1:0] node24429;
	wire [4-1:0] node24432;
	wire [4-1:0] node24434;
	wire [4-1:0] node24437;
	wire [4-1:0] node24438;
	wire [4-1:0] node24439;
	wire [4-1:0] node24443;
	wire [4-1:0] node24445;
	wire [4-1:0] node24446;
	wire [4-1:0] node24450;
	wire [4-1:0] node24451;
	wire [4-1:0] node24452;
	wire [4-1:0] node24453;
	wire [4-1:0] node24454;
	wire [4-1:0] node24456;
	wire [4-1:0] node24459;
	wire [4-1:0] node24460;
	wire [4-1:0] node24463;
	wire [4-1:0] node24466;
	wire [4-1:0] node24468;
	wire [4-1:0] node24469;
	wire [4-1:0] node24473;
	wire [4-1:0] node24474;
	wire [4-1:0] node24475;
	wire [4-1:0] node24477;
	wire [4-1:0] node24481;
	wire [4-1:0] node24482;
	wire [4-1:0] node24485;
	wire [4-1:0] node24488;
	wire [4-1:0] node24489;
	wire [4-1:0] node24490;
	wire [4-1:0] node24491;
	wire [4-1:0] node24494;
	wire [4-1:0] node24497;
	wire [4-1:0] node24498;
	wire [4-1:0] node24501;
	wire [4-1:0] node24504;
	wire [4-1:0] node24505;
	wire [4-1:0] node24506;
	wire [4-1:0] node24509;
	wire [4-1:0] node24513;
	wire [4-1:0] node24514;
	wire [4-1:0] node24515;
	wire [4-1:0] node24516;
	wire [4-1:0] node24517;
	wire [4-1:0] node24518;
	wire [4-1:0] node24519;
	wire [4-1:0] node24520;
	wire [4-1:0] node24524;
	wire [4-1:0] node24525;
	wire [4-1:0] node24528;
	wire [4-1:0] node24531;
	wire [4-1:0] node24532;
	wire [4-1:0] node24533;
	wire [4-1:0] node24534;
	wire [4-1:0] node24537;
	wire [4-1:0] node24540;
	wire [4-1:0] node24541;
	wire [4-1:0] node24544;
	wire [4-1:0] node24547;
	wire [4-1:0] node24548;
	wire [4-1:0] node24551;
	wire [4-1:0] node24554;
	wire [4-1:0] node24555;
	wire [4-1:0] node24556;
	wire [4-1:0] node24558;
	wire [4-1:0] node24561;
	wire [4-1:0] node24562;
	wire [4-1:0] node24563;
	wire [4-1:0] node24566;
	wire [4-1:0] node24570;
	wire [4-1:0] node24571;
	wire [4-1:0] node24572;
	wire [4-1:0] node24573;
	wire [4-1:0] node24578;
	wire [4-1:0] node24579;
	wire [4-1:0] node24580;
	wire [4-1:0] node24584;
	wire [4-1:0] node24585;
	wire [4-1:0] node24589;
	wire [4-1:0] node24590;
	wire [4-1:0] node24591;
	wire [4-1:0] node24592;
	wire [4-1:0] node24593;
	wire [4-1:0] node24597;
	wire [4-1:0] node24598;
	wire [4-1:0] node24602;
	wire [4-1:0] node24603;
	wire [4-1:0] node24604;
	wire [4-1:0] node24605;
	wire [4-1:0] node24610;
	wire [4-1:0] node24611;
	wire [4-1:0] node24614;
	wire [4-1:0] node24617;
	wire [4-1:0] node24618;
	wire [4-1:0] node24619;
	wire [4-1:0] node24620;
	wire [4-1:0] node24621;
	wire [4-1:0] node24625;
	wire [4-1:0] node24628;
	wire [4-1:0] node24629;
	wire [4-1:0] node24630;
	wire [4-1:0] node24633;
	wire [4-1:0] node24637;
	wire [4-1:0] node24638;
	wire [4-1:0] node24639;
	wire [4-1:0] node24640;
	wire [4-1:0] node24644;
	wire [4-1:0] node24645;
	wire [4-1:0] node24649;
	wire [4-1:0] node24650;
	wire [4-1:0] node24653;
	wire [4-1:0] node24654;
	wire [4-1:0] node24658;
	wire [4-1:0] node24659;
	wire [4-1:0] node24660;
	wire [4-1:0] node24661;
	wire [4-1:0] node24662;
	wire [4-1:0] node24664;
	wire [4-1:0] node24667;
	wire [4-1:0] node24668;
	wire [4-1:0] node24672;
	wire [4-1:0] node24673;
	wire [4-1:0] node24674;
	wire [4-1:0] node24676;
	wire [4-1:0] node24679;
	wire [4-1:0] node24680;
	wire [4-1:0] node24683;
	wire [4-1:0] node24686;
	wire [4-1:0] node24687;
	wire [4-1:0] node24690;
	wire [4-1:0] node24693;
	wire [4-1:0] node24694;
	wire [4-1:0] node24695;
	wire [4-1:0] node24697;
	wire [4-1:0] node24698;
	wire [4-1:0] node24702;
	wire [4-1:0] node24704;
	wire [4-1:0] node24705;
	wire [4-1:0] node24708;
	wire [4-1:0] node24711;
	wire [4-1:0] node24712;
	wire [4-1:0] node24713;
	wire [4-1:0] node24716;
	wire [4-1:0] node24719;
	wire [4-1:0] node24720;
	wire [4-1:0] node24721;
	wire [4-1:0] node24724;
	wire [4-1:0] node24728;
	wire [4-1:0] node24729;
	wire [4-1:0] node24730;
	wire [4-1:0] node24732;
	wire [4-1:0] node24733;
	wire [4-1:0] node24734;
	wire [4-1:0] node24738;
	wire [4-1:0] node24739;
	wire [4-1:0] node24743;
	wire [4-1:0] node24744;
	wire [4-1:0] node24745;
	wire [4-1:0] node24748;
	wire [4-1:0] node24751;
	wire [4-1:0] node24752;
	wire [4-1:0] node24753;
	wire [4-1:0] node24756;
	wire [4-1:0] node24759;
	wire [4-1:0] node24761;
	wire [4-1:0] node24764;
	wire [4-1:0] node24765;
	wire [4-1:0] node24766;
	wire [4-1:0] node24768;
	wire [4-1:0] node24771;
	wire [4-1:0] node24773;
	wire [4-1:0] node24776;
	wire [4-1:0] node24777;
	wire [4-1:0] node24778;
	wire [4-1:0] node24781;
	wire [4-1:0] node24784;
	wire [4-1:0] node24785;
	wire [4-1:0] node24789;
	wire [4-1:0] node24790;
	wire [4-1:0] node24791;
	wire [4-1:0] node24792;
	wire [4-1:0] node24793;
	wire [4-1:0] node24794;
	wire [4-1:0] node24795;
	wire [4-1:0] node24796;
	wire [4-1:0] node24800;
	wire [4-1:0] node24803;
	wire [4-1:0] node24805;
	wire [4-1:0] node24808;
	wire [4-1:0] node24809;
	wire [4-1:0] node24810;
	wire [4-1:0] node24814;
	wire [4-1:0] node24815;
	wire [4-1:0] node24816;
	wire [4-1:0] node24820;
	wire [4-1:0] node24821;
	wire [4-1:0] node24825;
	wire [4-1:0] node24826;
	wire [4-1:0] node24827;
	wire [4-1:0] node24828;
	wire [4-1:0] node24832;
	wire [4-1:0] node24833;
	wire [4-1:0] node24834;
	wire [4-1:0] node24839;
	wire [4-1:0] node24840;
	wire [4-1:0] node24843;
	wire [4-1:0] node24846;
	wire [4-1:0] node24847;
	wire [4-1:0] node24848;
	wire [4-1:0] node24849;
	wire [4-1:0] node24851;
	wire [4-1:0] node24852;
	wire [4-1:0] node24857;
	wire [4-1:0] node24860;
	wire [4-1:0] node24861;
	wire [4-1:0] node24862;
	wire [4-1:0] node24864;
	wire [4-1:0] node24867;
	wire [4-1:0] node24868;
	wire [4-1:0] node24869;
	wire [4-1:0] node24874;
	wire [4-1:0] node24876;
	wire [4-1:0] node24878;
	wire [4-1:0] node24881;
	wire [4-1:0] node24882;
	wire [4-1:0] node24883;
	wire [4-1:0] node24884;
	wire [4-1:0] node24885;
	wire [4-1:0] node24886;
	wire [4-1:0] node24887;
	wire [4-1:0] node24892;
	wire [4-1:0] node24893;
	wire [4-1:0] node24894;
	wire [4-1:0] node24899;
	wire [4-1:0] node24900;
	wire [4-1:0] node24901;
	wire [4-1:0] node24905;
	wire [4-1:0] node24906;
	wire [4-1:0] node24907;
	wire [4-1:0] node24912;
	wire [4-1:0] node24913;
	wire [4-1:0] node24914;
	wire [4-1:0] node24916;
	wire [4-1:0] node24917;
	wire [4-1:0] node24920;
	wire [4-1:0] node24923;
	wire [4-1:0] node24926;
	wire [4-1:0] node24927;
	wire [4-1:0] node24928;
	wire [4-1:0] node24931;
	wire [4-1:0] node24934;
	wire [4-1:0] node24935;
	wire [4-1:0] node24938;
	wire [4-1:0] node24941;
	wire [4-1:0] node24942;
	wire [4-1:0] node24943;
	wire [4-1:0] node24944;
	wire [4-1:0] node24946;
	wire [4-1:0] node24947;
	wire [4-1:0] node24951;
	wire [4-1:0] node24954;
	wire [4-1:0] node24955;
	wire [4-1:0] node24958;
	wire [4-1:0] node24960;
	wire [4-1:0] node24962;
	wire [4-1:0] node24965;
	wire [4-1:0] node24966;
	wire [4-1:0] node24967;
	wire [4-1:0] node24969;
	wire [4-1:0] node24971;
	wire [4-1:0] node24974;
	wire [4-1:0] node24977;
	wire [4-1:0] node24978;
	wire [4-1:0] node24979;
	wire [4-1:0] node24980;
	wire [4-1:0] node24984;
	wire [4-1:0] node24985;
	wire [4-1:0] node24988;
	wire [4-1:0] node24991;
	wire [4-1:0] node24993;
	wire [4-1:0] node24995;
	wire [4-1:0] node24998;
	wire [4-1:0] node24999;
	wire [4-1:0] node25000;
	wire [4-1:0] node25001;
	wire [4-1:0] node25002;
	wire [4-1:0] node25003;
	wire [4-1:0] node25004;
	wire [4-1:0] node25005;
	wire [4-1:0] node25006;
	wire [4-1:0] node25007;
	wire [4-1:0] node25009;
	wire [4-1:0] node25012;
	wire [4-1:0] node25015;
	wire [4-1:0] node25016;
	wire [4-1:0] node25019;
	wire [4-1:0] node25020;
	wire [4-1:0] node25023;
	wire [4-1:0] node25026;
	wire [4-1:0] node25028;
	wire [4-1:0] node25029;
	wire [4-1:0] node25030;
	wire [4-1:0] node25033;
	wire [4-1:0] node25036;
	wire [4-1:0] node25037;
	wire [4-1:0] node25040;
	wire [4-1:0] node25043;
	wire [4-1:0] node25044;
	wire [4-1:0] node25045;
	wire [4-1:0] node25046;
	wire [4-1:0] node25048;
	wire [4-1:0] node25051;
	wire [4-1:0] node25052;
	wire [4-1:0] node25056;
	wire [4-1:0] node25059;
	wire [4-1:0] node25060;
	wire [4-1:0] node25062;
	wire [4-1:0] node25064;
	wire [4-1:0] node25067;
	wire [4-1:0] node25068;
	wire [4-1:0] node25070;
	wire [4-1:0] node25074;
	wire [4-1:0] node25075;
	wire [4-1:0] node25076;
	wire [4-1:0] node25077;
	wire [4-1:0] node25079;
	wire [4-1:0] node25082;
	wire [4-1:0] node25083;
	wire [4-1:0] node25087;
	wire [4-1:0] node25088;
	wire [4-1:0] node25091;
	wire [4-1:0] node25093;
	wire [4-1:0] node25096;
	wire [4-1:0] node25097;
	wire [4-1:0] node25098;
	wire [4-1:0] node25099;
	wire [4-1:0] node25100;
	wire [4-1:0] node25103;
	wire [4-1:0] node25107;
	wire [4-1:0] node25109;
	wire [4-1:0] node25110;
	wire [4-1:0] node25113;
	wire [4-1:0] node25116;
	wire [4-1:0] node25117;
	wire [4-1:0] node25118;
	wire [4-1:0] node25119;
	wire [4-1:0] node25123;
	wire [4-1:0] node25124;
	wire [4-1:0] node25127;
	wire [4-1:0] node25130;
	wire [4-1:0] node25131;
	wire [4-1:0] node25135;
	wire [4-1:0] node25136;
	wire [4-1:0] node25137;
	wire [4-1:0] node25138;
	wire [4-1:0] node25139;
	wire [4-1:0] node25140;
	wire [4-1:0] node25141;
	wire [4-1:0] node25145;
	wire [4-1:0] node25147;
	wire [4-1:0] node25150;
	wire [4-1:0] node25151;
	wire [4-1:0] node25155;
	wire [4-1:0] node25156;
	wire [4-1:0] node25157;
	wire [4-1:0] node25158;
	wire [4-1:0] node25161;
	wire [4-1:0] node25164;
	wire [4-1:0] node25165;
	wire [4-1:0] node25169;
	wire [4-1:0] node25170;
	wire [4-1:0] node25171;
	wire [4-1:0] node25174;
	wire [4-1:0] node25177;
	wire [4-1:0] node25178;
	wire [4-1:0] node25181;
	wire [4-1:0] node25184;
	wire [4-1:0] node25185;
	wire [4-1:0] node25186;
	wire [4-1:0] node25187;
	wire [4-1:0] node25191;
	wire [4-1:0] node25192;
	wire [4-1:0] node25195;
	wire [4-1:0] node25197;
	wire [4-1:0] node25200;
	wire [4-1:0] node25201;
	wire [4-1:0] node25202;
	wire [4-1:0] node25205;
	wire [4-1:0] node25209;
	wire [4-1:0] node25210;
	wire [4-1:0] node25211;
	wire [4-1:0] node25212;
	wire [4-1:0] node25213;
	wire [4-1:0] node25214;
	wire [4-1:0] node25217;
	wire [4-1:0] node25220;
	wire [4-1:0] node25221;
	wire [4-1:0] node25224;
	wire [4-1:0] node25228;
	wire [4-1:0] node25229;
	wire [4-1:0] node25230;
	wire [4-1:0] node25232;
	wire [4-1:0] node25235;
	wire [4-1:0] node25236;
	wire [4-1:0] node25240;
	wire [4-1:0] node25241;
	wire [4-1:0] node25243;
	wire [4-1:0] node25246;
	wire [4-1:0] node25247;
	wire [4-1:0] node25250;
	wire [4-1:0] node25253;
	wire [4-1:0] node25254;
	wire [4-1:0] node25255;
	wire [4-1:0] node25256;
	wire [4-1:0] node25260;
	wire [4-1:0] node25261;
	wire [4-1:0] node25265;
	wire [4-1:0] node25266;
	wire [4-1:0] node25267;
	wire [4-1:0] node25269;
	wire [4-1:0] node25273;
	wire [4-1:0] node25276;
	wire [4-1:0] node25277;
	wire [4-1:0] node25278;
	wire [4-1:0] node25279;
	wire [4-1:0] node25280;
	wire [4-1:0] node25281;
	wire [4-1:0] node25284;
	wire [4-1:0] node25285;
	wire [4-1:0] node25289;
	wire [4-1:0] node25290;
	wire [4-1:0] node25291;
	wire [4-1:0] node25294;
	wire [4-1:0] node25297;
	wire [4-1:0] node25300;
	wire [4-1:0] node25301;
	wire [4-1:0] node25302;
	wire [4-1:0] node25305;
	wire [4-1:0] node25307;
	wire [4-1:0] node25310;
	wire [4-1:0] node25311;
	wire [4-1:0] node25312;
	wire [4-1:0] node25315;
	wire [4-1:0] node25319;
	wire [4-1:0] node25320;
	wire [4-1:0] node25321;
	wire [4-1:0] node25322;
	wire [4-1:0] node25323;
	wire [4-1:0] node25327;
	wire [4-1:0] node25329;
	wire [4-1:0] node25332;
	wire [4-1:0] node25333;
	wire [4-1:0] node25334;
	wire [4-1:0] node25337;
	wire [4-1:0] node25340;
	wire [4-1:0] node25341;
	wire [4-1:0] node25344;
	wire [4-1:0] node25345;
	wire [4-1:0] node25348;
	wire [4-1:0] node25351;
	wire [4-1:0] node25352;
	wire [4-1:0] node25353;
	wire [4-1:0] node25354;
	wire [4-1:0] node25355;
	wire [4-1:0] node25358;
	wire [4-1:0] node25361;
	wire [4-1:0] node25363;
	wire [4-1:0] node25366;
	wire [4-1:0] node25367;
	wire [4-1:0] node25370;
	wire [4-1:0] node25373;
	wire [4-1:0] node25374;
	wire [4-1:0] node25375;
	wire [4-1:0] node25379;
	wire [4-1:0] node25382;
	wire [4-1:0] node25383;
	wire [4-1:0] node25384;
	wire [4-1:0] node25385;
	wire [4-1:0] node25387;
	wire [4-1:0] node25388;
	wire [4-1:0] node25389;
	wire [4-1:0] node25392;
	wire [4-1:0] node25396;
	wire [4-1:0] node25397;
	wire [4-1:0] node25398;
	wire [4-1:0] node25401;
	wire [4-1:0] node25404;
	wire [4-1:0] node25405;
	wire [4-1:0] node25408;
	wire [4-1:0] node25411;
	wire [4-1:0] node25412;
	wire [4-1:0] node25413;
	wire [4-1:0] node25416;
	wire [4-1:0] node25418;
	wire [4-1:0] node25421;
	wire [4-1:0] node25422;
	wire [4-1:0] node25424;
	wire [4-1:0] node25427;
	wire [4-1:0] node25428;
	wire [4-1:0] node25432;
	wire [4-1:0] node25433;
	wire [4-1:0] node25434;
	wire [4-1:0] node25435;
	wire [4-1:0] node25436;
	wire [4-1:0] node25438;
	wire [4-1:0] node25441;
	wire [4-1:0] node25442;
	wire [4-1:0] node25445;
	wire [4-1:0] node25448;
	wire [4-1:0] node25449;
	wire [4-1:0] node25452;
	wire [4-1:0] node25455;
	wire [4-1:0] node25456;
	wire [4-1:0] node25457;
	wire [4-1:0] node25461;
	wire [4-1:0] node25464;
	wire [4-1:0] node25465;
	wire [4-1:0] node25466;
	wire [4-1:0] node25467;
	wire [4-1:0] node25471;
	wire [4-1:0] node25472;
	wire [4-1:0] node25475;
	wire [4-1:0] node25478;
	wire [4-1:0] node25479;
	wire [4-1:0] node25480;
	wire [4-1:0] node25484;
	wire [4-1:0] node25485;
	wire [4-1:0] node25486;
	wire [4-1:0] node25490;
	wire [4-1:0] node25493;
	wire [4-1:0] node25494;
	wire [4-1:0] node25495;
	wire [4-1:0] node25496;
	wire [4-1:0] node25497;
	wire [4-1:0] node25498;
	wire [4-1:0] node25500;
	wire [4-1:0] node25503;
	wire [4-1:0] node25504;
	wire [4-1:0] node25505;
	wire [4-1:0] node25507;
	wire [4-1:0] node25510;
	wire [4-1:0] node25512;
	wire [4-1:0] node25515;
	wire [4-1:0] node25516;
	wire [4-1:0] node25518;
	wire [4-1:0] node25521;
	wire [4-1:0] node25524;
	wire [4-1:0] node25525;
	wire [4-1:0] node25526;
	wire [4-1:0] node25528;
	wire [4-1:0] node25530;
	wire [4-1:0] node25533;
	wire [4-1:0] node25534;
	wire [4-1:0] node25538;
	wire [4-1:0] node25539;
	wire [4-1:0] node25540;
	wire [4-1:0] node25541;
	wire [4-1:0] node25546;
	wire [4-1:0] node25548;
	wire [4-1:0] node25551;
	wire [4-1:0] node25552;
	wire [4-1:0] node25553;
	wire [4-1:0] node25554;
	wire [4-1:0] node25555;
	wire [4-1:0] node25557;
	wire [4-1:0] node25560;
	wire [4-1:0] node25562;
	wire [4-1:0] node25565;
	wire [4-1:0] node25566;
	wire [4-1:0] node25570;
	wire [4-1:0] node25571;
	wire [4-1:0] node25573;
	wire [4-1:0] node25574;
	wire [4-1:0] node25578;
	wire [4-1:0] node25579;
	wire [4-1:0] node25583;
	wire [4-1:0] node25584;
	wire [4-1:0] node25585;
	wire [4-1:0] node25586;
	wire [4-1:0] node25587;
	wire [4-1:0] node25591;
	wire [4-1:0] node25592;
	wire [4-1:0] node25596;
	wire [4-1:0] node25597;
	wire [4-1:0] node25600;
	wire [4-1:0] node25601;
	wire [4-1:0] node25605;
	wire [4-1:0] node25606;
	wire [4-1:0] node25607;
	wire [4-1:0] node25608;
	wire [4-1:0] node25614;
	wire [4-1:0] node25615;
	wire [4-1:0] node25616;
	wire [4-1:0] node25617;
	wire [4-1:0] node25618;
	wire [4-1:0] node25621;
	wire [4-1:0] node25623;
	wire [4-1:0] node25625;
	wire [4-1:0] node25628;
	wire [4-1:0] node25629;
	wire [4-1:0] node25631;
	wire [4-1:0] node25634;
	wire [4-1:0] node25635;
	wire [4-1:0] node25637;
	wire [4-1:0] node25640;
	wire [4-1:0] node25642;
	wire [4-1:0] node25645;
	wire [4-1:0] node25646;
	wire [4-1:0] node25647;
	wire [4-1:0] node25648;
	wire [4-1:0] node25651;
	wire [4-1:0] node25655;
	wire [4-1:0] node25656;
	wire [4-1:0] node25658;
	wire [4-1:0] node25661;
	wire [4-1:0] node25662;
	wire [4-1:0] node25665;
	wire [4-1:0] node25668;
	wire [4-1:0] node25669;
	wire [4-1:0] node25670;
	wire [4-1:0] node25671;
	wire [4-1:0] node25673;
	wire [4-1:0] node25674;
	wire [4-1:0] node25678;
	wire [4-1:0] node25679;
	wire [4-1:0] node25680;
	wire [4-1:0] node25683;
	wire [4-1:0] node25687;
	wire [4-1:0] node25688;
	wire [4-1:0] node25689;
	wire [4-1:0] node25691;
	wire [4-1:0] node25695;
	wire [4-1:0] node25696;
	wire [4-1:0] node25697;
	wire [4-1:0] node25700;
	wire [4-1:0] node25703;
	wire [4-1:0] node25706;
	wire [4-1:0] node25707;
	wire [4-1:0] node25708;
	wire [4-1:0] node25710;
	wire [4-1:0] node25712;
	wire [4-1:0] node25715;
	wire [4-1:0] node25718;
	wire [4-1:0] node25719;
	wire [4-1:0] node25722;
	wire [4-1:0] node25723;
	wire [4-1:0] node25724;
	wire [4-1:0] node25727;
	wire [4-1:0] node25731;
	wire [4-1:0] node25732;
	wire [4-1:0] node25733;
	wire [4-1:0] node25734;
	wire [4-1:0] node25735;
	wire [4-1:0] node25736;
	wire [4-1:0] node25737;
	wire [4-1:0] node25740;
	wire [4-1:0] node25743;
	wire [4-1:0] node25744;
	wire [4-1:0] node25747;
	wire [4-1:0] node25750;
	wire [4-1:0] node25751;
	wire [4-1:0] node25752;
	wire [4-1:0] node25755;
	wire [4-1:0] node25759;
	wire [4-1:0] node25760;
	wire [4-1:0] node25761;
	wire [4-1:0] node25763;
	wire [4-1:0] node25767;
	wire [4-1:0] node25769;
	wire [4-1:0] node25771;
	wire [4-1:0] node25774;
	wire [4-1:0] node25775;
	wire [4-1:0] node25776;
	wire [4-1:0] node25777;
	wire [4-1:0] node25779;
	wire [4-1:0] node25782;
	wire [4-1:0] node25784;
	wire [4-1:0] node25787;
	wire [4-1:0] node25788;
	wire [4-1:0] node25790;
	wire [4-1:0] node25793;
	wire [4-1:0] node25795;
	wire [4-1:0] node25798;
	wire [4-1:0] node25799;
	wire [4-1:0] node25800;
	wire [4-1:0] node25802;
	wire [4-1:0] node25805;
	wire [4-1:0] node25806;
	wire [4-1:0] node25810;
	wire [4-1:0] node25811;
	wire [4-1:0] node25812;
	wire [4-1:0] node25814;
	wire [4-1:0] node25817;
	wire [4-1:0] node25819;
	wire [4-1:0] node25823;
	wire [4-1:0] node25824;
	wire [4-1:0] node25825;
	wire [4-1:0] node25826;
	wire [4-1:0] node25827;
	wire [4-1:0] node25828;
	wire [4-1:0] node25831;
	wire [4-1:0] node25834;
	wire [4-1:0] node25835;
	wire [4-1:0] node25838;
	wire [4-1:0] node25841;
	wire [4-1:0] node25842;
	wire [4-1:0] node25844;
	wire [4-1:0] node25845;
	wire [4-1:0] node25849;
	wire [4-1:0] node25850;
	wire [4-1:0] node25853;
	wire [4-1:0] node25856;
	wire [4-1:0] node25857;
	wire [4-1:0] node25858;
	wire [4-1:0] node25860;
	wire [4-1:0] node25863;
	wire [4-1:0] node25864;
	wire [4-1:0] node25867;
	wire [4-1:0] node25870;
	wire [4-1:0] node25871;
	wire [4-1:0] node25872;
	wire [4-1:0] node25875;
	wire [4-1:0] node25878;
	wire [4-1:0] node25879;
	wire [4-1:0] node25882;
	wire [4-1:0] node25885;
	wire [4-1:0] node25886;
	wire [4-1:0] node25887;
	wire [4-1:0] node25888;
	wire [4-1:0] node25889;
	wire [4-1:0] node25890;
	wire [4-1:0] node25893;
	wire [4-1:0] node25897;
	wire [4-1:0] node25899;
	wire [4-1:0] node25900;
	wire [4-1:0] node25903;
	wire [4-1:0] node25906;
	wire [4-1:0] node25907;
	wire [4-1:0] node25909;
	wire [4-1:0] node25912;
	wire [4-1:0] node25914;
	wire [4-1:0] node25917;
	wire [4-1:0] node25918;
	wire [4-1:0] node25919;
	wire [4-1:0] node25921;
	wire [4-1:0] node25924;
	wire [4-1:0] node25925;
	wire [4-1:0] node25926;
	wire [4-1:0] node25931;
	wire [4-1:0] node25932;
	wire [4-1:0] node25933;
	wire [4-1:0] node25936;
	wire [4-1:0] node25940;
	wire [4-1:0] node25941;
	wire [4-1:0] node25942;
	wire [4-1:0] node25943;
	wire [4-1:0] node25944;
	wire [4-1:0] node25945;
	wire [4-1:0] node25946;
	wire [4-1:0] node25947;
	wire [4-1:0] node25948;
	wire [4-1:0] node25949;
	wire [4-1:0] node25952;
	wire [4-1:0] node25956;
	wire [4-1:0] node25957;
	wire [4-1:0] node25959;
	wire [4-1:0] node25962;
	wire [4-1:0] node25965;
	wire [4-1:0] node25966;
	wire [4-1:0] node25967;
	wire [4-1:0] node25968;
	wire [4-1:0] node25971;
	wire [4-1:0] node25974;
	wire [4-1:0] node25975;
	wire [4-1:0] node25979;
	wire [4-1:0] node25980;
	wire [4-1:0] node25981;
	wire [4-1:0] node25985;
	wire [4-1:0] node25987;
	wire [4-1:0] node25990;
	wire [4-1:0] node25991;
	wire [4-1:0] node25992;
	wire [4-1:0] node25993;
	wire [4-1:0] node25995;
	wire [4-1:0] node25998;
	wire [4-1:0] node25999;
	wire [4-1:0] node26002;
	wire [4-1:0] node26005;
	wire [4-1:0] node26007;
	wire [4-1:0] node26010;
	wire [4-1:0] node26011;
	wire [4-1:0] node26012;
	wire [4-1:0] node26013;
	wire [4-1:0] node26017;
	wire [4-1:0] node26018;
	wire [4-1:0] node26022;
	wire [4-1:0] node26024;
	wire [4-1:0] node26027;
	wire [4-1:0] node26028;
	wire [4-1:0] node26029;
	wire [4-1:0] node26030;
	wire [4-1:0] node26032;
	wire [4-1:0] node26033;
	wire [4-1:0] node26037;
	wire [4-1:0] node26040;
	wire [4-1:0] node26041;
	wire [4-1:0] node26043;
	wire [4-1:0] node26045;
	wire [4-1:0] node26049;
	wire [4-1:0] node26050;
	wire [4-1:0] node26051;
	wire [4-1:0] node26053;
	wire [4-1:0] node26054;
	wire [4-1:0] node26058;
	wire [4-1:0] node26059;
	wire [4-1:0] node26062;
	wire [4-1:0] node26065;
	wire [4-1:0] node26066;
	wire [4-1:0] node26067;
	wire [4-1:0] node26068;
	wire [4-1:0] node26071;
	wire [4-1:0] node26075;
	wire [4-1:0] node26076;
	wire [4-1:0] node26077;
	wire [4-1:0] node26081;
	wire [4-1:0] node26084;
	wire [4-1:0] node26085;
	wire [4-1:0] node26086;
	wire [4-1:0] node26087;
	wire [4-1:0] node26089;
	wire [4-1:0] node26090;
	wire [4-1:0] node26092;
	wire [4-1:0] node26095;
	wire [4-1:0] node26096;
	wire [4-1:0] node26099;
	wire [4-1:0] node26102;
	wire [4-1:0] node26103;
	wire [4-1:0] node26104;
	wire [4-1:0] node26105;
	wire [4-1:0] node26110;
	wire [4-1:0] node26111;
	wire [4-1:0] node26112;
	wire [4-1:0] node26115;
	wire [4-1:0] node26119;
	wire [4-1:0] node26120;
	wire [4-1:0] node26121;
	wire [4-1:0] node26122;
	wire [4-1:0] node26123;
	wire [4-1:0] node26126;
	wire [4-1:0] node26130;
	wire [4-1:0] node26131;
	wire [4-1:0] node26132;
	wire [4-1:0] node26135;
	wire [4-1:0] node26139;
	wire [4-1:0] node26140;
	wire [4-1:0] node26141;
	wire [4-1:0] node26145;
	wire [4-1:0] node26147;
	wire [4-1:0] node26150;
	wire [4-1:0] node26151;
	wire [4-1:0] node26152;
	wire [4-1:0] node26155;
	wire [4-1:0] node26157;
	wire [4-1:0] node26158;
	wire [4-1:0] node26159;
	wire [4-1:0] node26162;
	wire [4-1:0] node26166;
	wire [4-1:0] node26167;
	wire [4-1:0] node26168;
	wire [4-1:0] node26170;
	wire [4-1:0] node26171;
	wire [4-1:0] node26175;
	wire [4-1:0] node26177;
	wire [4-1:0] node26178;
	wire [4-1:0] node26181;
	wire [4-1:0] node26184;
	wire [4-1:0] node26185;
	wire [4-1:0] node26186;
	wire [4-1:0] node26187;
	wire [4-1:0] node26190;
	wire [4-1:0] node26193;
	wire [4-1:0] node26196;
	wire [4-1:0] node26197;
	wire [4-1:0] node26200;
	wire [4-1:0] node26203;
	wire [4-1:0] node26204;
	wire [4-1:0] node26205;
	wire [4-1:0] node26206;
	wire [4-1:0] node26207;
	wire [4-1:0] node26208;
	wire [4-1:0] node26209;
	wire [4-1:0] node26212;
	wire [4-1:0] node26215;
	wire [4-1:0] node26216;
	wire [4-1:0] node26220;
	wire [4-1:0] node26221;
	wire [4-1:0] node26223;
	wire [4-1:0] node26225;
	wire [4-1:0] node26228;
	wire [4-1:0] node26229;
	wire [4-1:0] node26231;
	wire [4-1:0] node26234;
	wire [4-1:0] node26235;
	wire [4-1:0] node26239;
	wire [4-1:0] node26240;
	wire [4-1:0] node26241;
	wire [4-1:0] node26242;
	wire [4-1:0] node26245;
	wire [4-1:0] node26247;
	wire [4-1:0] node26250;
	wire [4-1:0] node26251;
	wire [4-1:0] node26253;
	wire [4-1:0] node26256;
	wire [4-1:0] node26259;
	wire [4-1:0] node26260;
	wire [4-1:0] node26261;
	wire [4-1:0] node26264;
	wire [4-1:0] node26267;
	wire [4-1:0] node26268;
	wire [4-1:0] node26269;
	wire [4-1:0] node26273;
	wire [4-1:0] node26274;
	wire [4-1:0] node26278;
	wire [4-1:0] node26279;
	wire [4-1:0] node26280;
	wire [4-1:0] node26281;
	wire [4-1:0] node26282;
	wire [4-1:0] node26283;
	wire [4-1:0] node26286;
	wire [4-1:0] node26290;
	wire [4-1:0] node26291;
	wire [4-1:0] node26295;
	wire [4-1:0] node26296;
	wire [4-1:0] node26298;
	wire [4-1:0] node26299;
	wire [4-1:0] node26302;
	wire [4-1:0] node26305;
	wire [4-1:0] node26308;
	wire [4-1:0] node26309;
	wire [4-1:0] node26310;
	wire [4-1:0] node26311;
	wire [4-1:0] node26312;
	wire [4-1:0] node26315;
	wire [4-1:0] node26318;
	wire [4-1:0] node26319;
	wire [4-1:0] node26322;
	wire [4-1:0] node26325;
	wire [4-1:0] node26326;
	wire [4-1:0] node26327;
	wire [4-1:0] node26330;
	wire [4-1:0] node26333;
	wire [4-1:0] node26334;
	wire [4-1:0] node26337;
	wire [4-1:0] node26340;
	wire [4-1:0] node26341;
	wire [4-1:0] node26342;
	wire [4-1:0] node26343;
	wire [4-1:0] node26346;
	wire [4-1:0] node26350;
	wire [4-1:0] node26351;
	wire [4-1:0] node26352;
	wire [4-1:0] node26356;
	wire [4-1:0] node26359;
	wire [4-1:0] node26360;
	wire [4-1:0] node26361;
	wire [4-1:0] node26362;
	wire [4-1:0] node26363;
	wire [4-1:0] node26365;
	wire [4-1:0] node26366;
	wire [4-1:0] node26370;
	wire [4-1:0] node26371;
	wire [4-1:0] node26372;
	wire [4-1:0] node26375;
	wire [4-1:0] node26378;
	wire [4-1:0] node26381;
	wire [4-1:0] node26382;
	wire [4-1:0] node26383;
	wire [4-1:0] node26386;
	wire [4-1:0] node26388;
	wire [4-1:0] node26391;
	wire [4-1:0] node26392;
	wire [4-1:0] node26393;
	wire [4-1:0] node26396;
	wire [4-1:0] node26399;
	wire [4-1:0] node26402;
	wire [4-1:0] node26403;
	wire [4-1:0] node26404;
	wire [4-1:0] node26405;
	wire [4-1:0] node26407;
	wire [4-1:0] node26410;
	wire [4-1:0] node26411;
	wire [4-1:0] node26414;
	wire [4-1:0] node26417;
	wire [4-1:0] node26418;
	wire [4-1:0] node26419;
	wire [4-1:0] node26424;
	wire [4-1:0] node26425;
	wire [4-1:0] node26427;
	wire [4-1:0] node26428;
	wire [4-1:0] node26432;
	wire [4-1:0] node26433;
	wire [4-1:0] node26435;
	wire [4-1:0] node26438;
	wire [4-1:0] node26441;
	wire [4-1:0] node26442;
	wire [4-1:0] node26443;
	wire [4-1:0] node26444;
	wire [4-1:0] node26445;
	wire [4-1:0] node26448;
	wire [4-1:0] node26450;
	wire [4-1:0] node26453;
	wire [4-1:0] node26454;
	wire [4-1:0] node26455;
	wire [4-1:0] node26459;
	wire [4-1:0] node26462;
	wire [4-1:0] node26463;
	wire [4-1:0] node26464;
	wire [4-1:0] node26465;
	wire [4-1:0] node26468;
	wire [4-1:0] node26471;
	wire [4-1:0] node26474;
	wire [4-1:0] node26475;
	wire [4-1:0] node26476;
	wire [4-1:0] node26480;
	wire [4-1:0] node26482;
	wire [4-1:0] node26485;
	wire [4-1:0] node26486;
	wire [4-1:0] node26487;
	wire [4-1:0] node26488;
	wire [4-1:0] node26490;
	wire [4-1:0] node26493;
	wire [4-1:0] node26496;
	wire [4-1:0] node26497;
	wire [4-1:0] node26498;
	wire [4-1:0] node26503;
	wire [4-1:0] node26504;
	wire [4-1:0] node26505;
	wire [4-1:0] node26508;
	wire [4-1:0] node26509;
	wire [4-1:0] node26512;
	wire [4-1:0] node26515;
	wire [4-1:0] node26516;
	wire [4-1:0] node26519;
	wire [4-1:0] node26522;
	wire [4-1:0] node26523;
	wire [4-1:0] node26524;
	wire [4-1:0] node26525;
	wire [4-1:0] node26526;
	wire [4-1:0] node26527;
	wire [4-1:0] node26529;
	wire [4-1:0] node26530;
	wire [4-1:0] node26532;
	wire [4-1:0] node26536;
	wire [4-1:0] node26537;
	wire [4-1:0] node26539;
	wire [4-1:0] node26541;
	wire [4-1:0] node26544;
	wire [4-1:0] node26545;
	wire [4-1:0] node26546;
	wire [4-1:0] node26549;
	wire [4-1:0] node26552;
	wire [4-1:0] node26553;
	wire [4-1:0] node26557;
	wire [4-1:0] node26558;
	wire [4-1:0] node26559;
	wire [4-1:0] node26560;
	wire [4-1:0] node26563;
	wire [4-1:0] node26565;
	wire [4-1:0] node26568;
	wire [4-1:0] node26569;
	wire [4-1:0] node26573;
	wire [4-1:0] node26574;
	wire [4-1:0] node26576;
	wire [4-1:0] node26579;
	wire [4-1:0] node26581;
	wire [4-1:0] node26582;
	wire [4-1:0] node26586;
	wire [4-1:0] node26587;
	wire [4-1:0] node26588;
	wire [4-1:0] node26589;
	wire [4-1:0] node26591;
	wire [4-1:0] node26593;
	wire [4-1:0] node26596;
	wire [4-1:0] node26597;
	wire [4-1:0] node26601;
	wire [4-1:0] node26602;
	wire [4-1:0] node26603;
	wire [4-1:0] node26605;
	wire [4-1:0] node26608;
	wire [4-1:0] node26610;
	wire [4-1:0] node26613;
	wire [4-1:0] node26614;
	wire [4-1:0] node26618;
	wire [4-1:0] node26619;
	wire [4-1:0] node26620;
	wire [4-1:0] node26621;
	wire [4-1:0] node26622;
	wire [4-1:0] node26626;
	wire [4-1:0] node26629;
	wire [4-1:0] node26630;
	wire [4-1:0] node26631;
	wire [4-1:0] node26634;
	wire [4-1:0] node26638;
	wire [4-1:0] node26639;
	wire [4-1:0] node26640;
	wire [4-1:0] node26641;
	wire [4-1:0] node26646;
	wire [4-1:0] node26647;
	wire [4-1:0] node26651;
	wire [4-1:0] node26652;
	wire [4-1:0] node26653;
	wire [4-1:0] node26654;
	wire [4-1:0] node26656;
	wire [4-1:0] node26658;
	wire [4-1:0] node26661;
	wire [4-1:0] node26662;
	wire [4-1:0] node26663;
	wire [4-1:0] node26666;
	wire [4-1:0] node26669;
	wire [4-1:0] node26670;
	wire [4-1:0] node26671;
	wire [4-1:0] node26675;
	wire [4-1:0] node26676;
	wire [4-1:0] node26679;
	wire [4-1:0] node26682;
	wire [4-1:0] node26683;
	wire [4-1:0] node26684;
	wire [4-1:0] node26685;
	wire [4-1:0] node26689;
	wire [4-1:0] node26690;
	wire [4-1:0] node26691;
	wire [4-1:0] node26696;
	wire [4-1:0] node26697;
	wire [4-1:0] node26698;
	wire [4-1:0] node26700;
	wire [4-1:0] node26704;
	wire [4-1:0] node26705;
	wire [4-1:0] node26708;
	wire [4-1:0] node26711;
	wire [4-1:0] node26712;
	wire [4-1:0] node26713;
	wire [4-1:0] node26714;
	wire [4-1:0] node26715;
	wire [4-1:0] node26719;
	wire [4-1:0] node26720;
	wire [4-1:0] node26721;
	wire [4-1:0] node26726;
	wire [4-1:0] node26727;
	wire [4-1:0] node26728;
	wire [4-1:0] node26730;
	wire [4-1:0] node26733;
	wire [4-1:0] node26735;
	wire [4-1:0] node26738;
	wire [4-1:0] node26739;
	wire [4-1:0] node26740;
	wire [4-1:0] node26745;
	wire [4-1:0] node26746;
	wire [4-1:0] node26747;
	wire [4-1:0] node26748;
	wire [4-1:0] node26750;
	wire [4-1:0] node26754;
	wire [4-1:0] node26755;
	wire [4-1:0] node26758;
	wire [4-1:0] node26761;
	wire [4-1:0] node26762;
	wire [4-1:0] node26764;
	wire [4-1:0] node26765;
	wire [4-1:0] node26769;
	wire [4-1:0] node26770;
	wire [4-1:0] node26772;
	wire [4-1:0] node26775;
	wire [4-1:0] node26776;
	wire [4-1:0] node26779;
	wire [4-1:0] node26782;
	wire [4-1:0] node26783;
	wire [4-1:0] node26784;
	wire [4-1:0] node26785;
	wire [4-1:0] node26786;
	wire [4-1:0] node26787;
	wire [4-1:0] node26789;
	wire [4-1:0] node26792;
	wire [4-1:0] node26794;
	wire [4-1:0] node26797;
	wire [4-1:0] node26798;
	wire [4-1:0] node26800;
	wire [4-1:0] node26803;
	wire [4-1:0] node26805;
	wire [4-1:0] node26808;
	wire [4-1:0] node26809;
	wire [4-1:0] node26811;
	wire [4-1:0] node26813;
	wire [4-1:0] node26816;
	wire [4-1:0] node26818;
	wire [4-1:0] node26820;
	wire [4-1:0] node26823;
	wire [4-1:0] node26824;
	wire [4-1:0] node26825;
	wire [4-1:0] node26826;
	wire [4-1:0] node26829;
	wire [4-1:0] node26832;
	wire [4-1:0] node26833;
	wire [4-1:0] node26834;
	wire [4-1:0] node26837;
	wire [4-1:0] node26840;
	wire [4-1:0] node26841;
	wire [4-1:0] node26845;
	wire [4-1:0] node26846;
	wire [4-1:0] node26847;
	wire [4-1:0] node26848;
	wire [4-1:0] node26851;
	wire [4-1:0] node26854;
	wire [4-1:0] node26855;
	wire [4-1:0] node26859;
	wire [4-1:0] node26860;
	wire [4-1:0] node26861;
	wire [4-1:0] node26864;
	wire [4-1:0] node26867;
	wire [4-1:0] node26868;
	wire [4-1:0] node26869;
	wire [4-1:0] node26872;
	wire [4-1:0] node26875;
	wire [4-1:0] node26876;
	wire [4-1:0] node26879;
	wire [4-1:0] node26882;
	wire [4-1:0] node26883;
	wire [4-1:0] node26884;
	wire [4-1:0] node26885;
	wire [4-1:0] node26886;
	wire [4-1:0] node26887;
	wire [4-1:0] node26890;
	wire [4-1:0] node26893;
	wire [4-1:0] node26894;
	wire [4-1:0] node26896;
	wire [4-1:0] node26899;
	wire [4-1:0] node26900;
	wire [4-1:0] node26903;
	wire [4-1:0] node26906;
	wire [4-1:0] node26907;
	wire [4-1:0] node26908;
	wire [4-1:0] node26909;
	wire [4-1:0] node26912;
	wire [4-1:0] node26917;
	wire [4-1:0] node26918;
	wire [4-1:0] node26919;
	wire [4-1:0] node26921;
	wire [4-1:0] node26924;
	wire [4-1:0] node26925;
	wire [4-1:0] node26928;
	wire [4-1:0] node26931;
	wire [4-1:0] node26932;
	wire [4-1:0] node26933;
	wire [4-1:0] node26934;
	wire [4-1:0] node26937;
	wire [4-1:0] node26940;
	wire [4-1:0] node26941;
	wire [4-1:0] node26944;
	wire [4-1:0] node26947;
	wire [4-1:0] node26949;
	wire [4-1:0] node26952;
	wire [4-1:0] node26953;
	wire [4-1:0] node26954;
	wire [4-1:0] node26955;
	wire [4-1:0] node26957;
	wire [4-1:0] node26960;
	wire [4-1:0] node26961;
	wire [4-1:0] node26964;
	wire [4-1:0] node26967;
	wire [4-1:0] node26968;
	wire [4-1:0] node26970;
	wire [4-1:0] node26973;
	wire [4-1:0] node26974;
	wire [4-1:0] node26977;
	wire [4-1:0] node26980;
	wire [4-1:0] node26981;
	wire [4-1:0] node26982;
	wire [4-1:0] node26983;
	wire [4-1:0] node26984;
	wire [4-1:0] node26987;
	wire [4-1:0] node26990;
	wire [4-1:0] node26991;
	wire [4-1:0] node26994;
	wire [4-1:0] node26997;
	wire [4-1:0] node27000;
	wire [4-1:0] node27001;
	wire [4-1:0] node27002;
	wire [4-1:0] node27005;
	wire [4-1:0] node27008;
	wire [4-1:0] node27009;
	wire [4-1:0] node27012;
	wire [4-1:0] node27015;
	wire [4-1:0] node27016;
	wire [4-1:0] node27017;
	wire [4-1:0] node27018;
	wire [4-1:0] node27019;
	wire [4-1:0] node27020;
	wire [4-1:0] node27021;
	wire [4-1:0] node27022;
	wire [4-1:0] node27023;
	wire [4-1:0] node27024;
	wire [4-1:0] node27026;
	wire [4-1:0] node27028;
	wire [4-1:0] node27031;
	wire [4-1:0] node27032;
	wire [4-1:0] node27035;
	wire [4-1:0] node27038;
	wire [4-1:0] node27039;
	wire [4-1:0] node27040;
	wire [4-1:0] node27043;
	wire [4-1:0] node27046;
	wire [4-1:0] node27047;
	wire [4-1:0] node27050;
	wire [4-1:0] node27053;
	wire [4-1:0] node27054;
	wire [4-1:0] node27055;
	wire [4-1:0] node27056;
	wire [4-1:0] node27060;
	wire [4-1:0] node27062;
	wire [4-1:0] node27065;
	wire [4-1:0] node27066;
	wire [4-1:0] node27068;
	wire [4-1:0] node27069;
	wire [4-1:0] node27072;
	wire [4-1:0] node27075;
	wire [4-1:0] node27076;
	wire [4-1:0] node27079;
	wire [4-1:0] node27082;
	wire [4-1:0] node27083;
	wire [4-1:0] node27084;
	wire [4-1:0] node27085;
	wire [4-1:0] node27086;
	wire [4-1:0] node27089;
	wire [4-1:0] node27090;
	wire [4-1:0] node27093;
	wire [4-1:0] node27096;
	wire [4-1:0] node27098;
	wire [4-1:0] node27099;
	wire [4-1:0] node27103;
	wire [4-1:0] node27104;
	wire [4-1:0] node27105;
	wire [4-1:0] node27108;
	wire [4-1:0] node27111;
	wire [4-1:0] node27113;
	wire [4-1:0] node27116;
	wire [4-1:0] node27117;
	wire [4-1:0] node27118;
	wire [4-1:0] node27119;
	wire [4-1:0] node27120;
	wire [4-1:0] node27123;
	wire [4-1:0] node27126;
	wire [4-1:0] node27127;
	wire [4-1:0] node27131;
	wire [4-1:0] node27132;
	wire [4-1:0] node27136;
	wire [4-1:0] node27137;
	wire [4-1:0] node27138;
	wire [4-1:0] node27141;
	wire [4-1:0] node27144;
	wire [4-1:0] node27145;
	wire [4-1:0] node27148;
	wire [4-1:0] node27151;
	wire [4-1:0] node27152;
	wire [4-1:0] node27153;
	wire [4-1:0] node27154;
	wire [4-1:0] node27155;
	wire [4-1:0] node27156;
	wire [4-1:0] node27157;
	wire [4-1:0] node27161;
	wire [4-1:0] node27162;
	wire [4-1:0] node27166;
	wire [4-1:0] node27168;
	wire [4-1:0] node27169;
	wire [4-1:0] node27172;
	wire [4-1:0] node27175;
	wire [4-1:0] node27176;
	wire [4-1:0] node27178;
	wire [4-1:0] node27179;
	wire [4-1:0] node27183;
	wire [4-1:0] node27184;
	wire [4-1:0] node27185;
	wire [4-1:0] node27189;
	wire [4-1:0] node27191;
	wire [4-1:0] node27194;
	wire [4-1:0] node27195;
	wire [4-1:0] node27196;
	wire [4-1:0] node27198;
	wire [4-1:0] node27199;
	wire [4-1:0] node27202;
	wire [4-1:0] node27205;
	wire [4-1:0] node27207;
	wire [4-1:0] node27210;
	wire [4-1:0] node27212;
	wire [4-1:0] node27213;
	wire [4-1:0] node27214;
	wire [4-1:0] node27217;
	wire [4-1:0] node27220;
	wire [4-1:0] node27221;
	wire [4-1:0] node27225;
	wire [4-1:0] node27226;
	wire [4-1:0] node27227;
	wire [4-1:0] node27228;
	wire [4-1:0] node27229;
	wire [4-1:0] node27232;
	wire [4-1:0] node27235;
	wire [4-1:0] node27236;
	wire [4-1:0] node27240;
	wire [4-1:0] node27241;
	wire [4-1:0] node27242;
	wire [4-1:0] node27243;
	wire [4-1:0] node27246;
	wire [4-1:0] node27250;
	wire [4-1:0] node27252;
	wire [4-1:0] node27254;
	wire [4-1:0] node27257;
	wire [4-1:0] node27258;
	wire [4-1:0] node27259;
	wire [4-1:0] node27262;
	wire [4-1:0] node27263;
	wire [4-1:0] node27264;
	wire [4-1:0] node27267;
	wire [4-1:0] node27271;
	wire [4-1:0] node27272;
	wire [4-1:0] node27274;
	wire [4-1:0] node27278;
	wire [4-1:0] node27279;
	wire [4-1:0] node27280;
	wire [4-1:0] node27281;
	wire [4-1:0] node27282;
	wire [4-1:0] node27283;
	wire [4-1:0] node27285;
	wire [4-1:0] node27288;
	wire [4-1:0] node27291;
	wire [4-1:0] node27293;
	wire [4-1:0] node27295;
	wire [4-1:0] node27298;
	wire [4-1:0] node27299;
	wire [4-1:0] node27300;
	wire [4-1:0] node27303;
	wire [4-1:0] node27305;
	wire [4-1:0] node27308;
	wire [4-1:0] node27309;
	wire [4-1:0] node27310;
	wire [4-1:0] node27314;
	wire [4-1:0] node27317;
	wire [4-1:0] node27318;
	wire [4-1:0] node27319;
	wire [4-1:0] node27320;
	wire [4-1:0] node27321;
	wire [4-1:0] node27324;
	wire [4-1:0] node27325;
	wire [4-1:0] node27329;
	wire [4-1:0] node27331;
	wire [4-1:0] node27334;
	wire [4-1:0] node27335;
	wire [4-1:0] node27336;
	wire [4-1:0] node27339;
	wire [4-1:0] node27342;
	wire [4-1:0] node27343;
	wire [4-1:0] node27344;
	wire [4-1:0] node27347;
	wire [4-1:0] node27350;
	wire [4-1:0] node27351;
	wire [4-1:0] node27355;
	wire [4-1:0] node27356;
	wire [4-1:0] node27357;
	wire [4-1:0] node27358;
	wire [4-1:0] node27360;
	wire [4-1:0] node27363;
	wire [4-1:0] node27365;
	wire [4-1:0] node27368;
	wire [4-1:0] node27370;
	wire [4-1:0] node27373;
	wire [4-1:0] node27374;
	wire [4-1:0] node27375;
	wire [4-1:0] node27378;
	wire [4-1:0] node27380;
	wire [4-1:0] node27383;
	wire [4-1:0] node27384;
	wire [4-1:0] node27387;
	wire [4-1:0] node27390;
	wire [4-1:0] node27391;
	wire [4-1:0] node27392;
	wire [4-1:0] node27393;
	wire [4-1:0] node27394;
	wire [4-1:0] node27397;
	wire [4-1:0] node27400;
	wire [4-1:0] node27401;
	wire [4-1:0] node27403;
	wire [4-1:0] node27404;
	wire [4-1:0] node27408;
	wire [4-1:0] node27409;
	wire [4-1:0] node27412;
	wire [4-1:0] node27415;
	wire [4-1:0] node27416;
	wire [4-1:0] node27417;
	wire [4-1:0] node27418;
	wire [4-1:0] node27421;
	wire [4-1:0] node27424;
	wire [4-1:0] node27425;
	wire [4-1:0] node27428;
	wire [4-1:0] node27431;
	wire [4-1:0] node27432;
	wire [4-1:0] node27433;
	wire [4-1:0] node27434;
	wire [4-1:0] node27438;
	wire [4-1:0] node27441;
	wire [4-1:0] node27442;
	wire [4-1:0] node27445;
	wire [4-1:0] node27448;
	wire [4-1:0] node27449;
	wire [4-1:0] node27450;
	wire [4-1:0] node27451;
	wire [4-1:0] node27452;
	wire [4-1:0] node27455;
	wire [4-1:0] node27458;
	wire [4-1:0] node27459;
	wire [4-1:0] node27463;
	wire [4-1:0] node27464;
	wire [4-1:0] node27465;
	wire [4-1:0] node27466;
	wire [4-1:0] node27470;
	wire [4-1:0] node27471;
	wire [4-1:0] node27474;
	wire [4-1:0] node27477;
	wire [4-1:0] node27478;
	wire [4-1:0] node27481;
	wire [4-1:0] node27484;
	wire [4-1:0] node27485;
	wire [4-1:0] node27486;
	wire [4-1:0] node27488;
	wire [4-1:0] node27489;
	wire [4-1:0] node27492;
	wire [4-1:0] node27495;
	wire [4-1:0] node27496;
	wire [4-1:0] node27499;
	wire [4-1:0] node27502;
	wire [4-1:0] node27503;
	wire [4-1:0] node27504;
	wire [4-1:0] node27507;
	wire [4-1:0] node27510;
	wire [4-1:0] node27511;
	wire [4-1:0] node27514;
	wire [4-1:0] node27517;
	wire [4-1:0] node27518;
	wire [4-1:0] node27519;
	wire [4-1:0] node27520;
	wire [4-1:0] node27521;
	wire [4-1:0] node27522;
	wire [4-1:0] node27524;
	wire [4-1:0] node27526;
	wire [4-1:0] node27527;
	wire [4-1:0] node27531;
	wire [4-1:0] node27532;
	wire [4-1:0] node27534;
	wire [4-1:0] node27535;
	wire [4-1:0] node27539;
	wire [4-1:0] node27540;
	wire [4-1:0] node27541;
	wire [4-1:0] node27544;
	wire [4-1:0] node27547;
	wire [4-1:0] node27548;
	wire [4-1:0] node27552;
	wire [4-1:0] node27553;
	wire [4-1:0] node27554;
	wire [4-1:0] node27556;
	wire [4-1:0] node27559;
	wire [4-1:0] node27560;
	wire [4-1:0] node27562;
	wire [4-1:0] node27566;
	wire [4-1:0] node27567;
	wire [4-1:0] node27568;
	wire [4-1:0] node27569;
	wire [4-1:0] node27573;
	wire [4-1:0] node27574;
	wire [4-1:0] node27578;
	wire [4-1:0] node27581;
	wire [4-1:0] node27582;
	wire [4-1:0] node27583;
	wire [4-1:0] node27584;
	wire [4-1:0] node27585;
	wire [4-1:0] node27588;
	wire [4-1:0] node27590;
	wire [4-1:0] node27593;
	wire [4-1:0] node27594;
	wire [4-1:0] node27598;
	wire [4-1:0] node27599;
	wire [4-1:0] node27600;
	wire [4-1:0] node27603;
	wire [4-1:0] node27604;
	wire [4-1:0] node27609;
	wire [4-1:0] node27610;
	wire [4-1:0] node27611;
	wire [4-1:0] node27612;
	wire [4-1:0] node27616;
	wire [4-1:0] node27617;
	wire [4-1:0] node27619;
	wire [4-1:0] node27622;
	wire [4-1:0] node27625;
	wire [4-1:0] node27626;
	wire [4-1:0] node27627;
	wire [4-1:0] node27630;
	wire [4-1:0] node27631;
	wire [4-1:0] node27634;
	wire [4-1:0] node27637;
	wire [4-1:0] node27638;
	wire [4-1:0] node27641;
	wire [4-1:0] node27644;
	wire [4-1:0] node27645;
	wire [4-1:0] node27646;
	wire [4-1:0] node27647;
	wire [4-1:0] node27648;
	wire [4-1:0] node27650;
	wire [4-1:0] node27653;
	wire [4-1:0] node27654;
	wire [4-1:0] node27658;
	wire [4-1:0] node27659;
	wire [4-1:0] node27660;
	wire [4-1:0] node27661;
	wire [4-1:0] node27664;
	wire [4-1:0] node27667;
	wire [4-1:0] node27668;
	wire [4-1:0] node27671;
	wire [4-1:0] node27674;
	wire [4-1:0] node27676;
	wire [4-1:0] node27677;
	wire [4-1:0] node27681;
	wire [4-1:0] node27682;
	wire [4-1:0] node27683;
	wire [4-1:0] node27684;
	wire [4-1:0] node27688;
	wire [4-1:0] node27689;
	wire [4-1:0] node27692;
	wire [4-1:0] node27693;
	wire [4-1:0] node27697;
	wire [4-1:0] node27698;
	wire [4-1:0] node27700;
	wire [4-1:0] node27701;
	wire [4-1:0] node27704;
	wire [4-1:0] node27707;
	wire [4-1:0] node27708;
	wire [4-1:0] node27709;
	wire [4-1:0] node27713;
	wire [4-1:0] node27715;
	wire [4-1:0] node27718;
	wire [4-1:0] node27719;
	wire [4-1:0] node27720;
	wire [4-1:0] node27721;
	wire [4-1:0] node27723;
	wire [4-1:0] node27724;
	wire [4-1:0] node27727;
	wire [4-1:0] node27731;
	wire [4-1:0] node27732;
	wire [4-1:0] node27733;
	wire [4-1:0] node27735;
	wire [4-1:0] node27739;
	wire [4-1:0] node27740;
	wire [4-1:0] node27743;
	wire [4-1:0] node27746;
	wire [4-1:0] node27747;
	wire [4-1:0] node27748;
	wire [4-1:0] node27749;
	wire [4-1:0] node27751;
	wire [4-1:0] node27754;
	wire [4-1:0] node27757;
	wire [4-1:0] node27760;
	wire [4-1:0] node27761;
	wire [4-1:0] node27763;
	wire [4-1:0] node27766;
	wire [4-1:0] node27767;
	wire [4-1:0] node27769;
	wire [4-1:0] node27772;
	wire [4-1:0] node27773;
	wire [4-1:0] node27777;
	wire [4-1:0] node27778;
	wire [4-1:0] node27779;
	wire [4-1:0] node27780;
	wire [4-1:0] node27781;
	wire [4-1:0] node27782;
	wire [4-1:0] node27785;
	wire [4-1:0] node27788;
	wire [4-1:0] node27789;
	wire [4-1:0] node27790;
	wire [4-1:0] node27793;
	wire [4-1:0] node27796;
	wire [4-1:0] node27797;
	wire [4-1:0] node27798;
	wire [4-1:0] node27801;
	wire [4-1:0] node27804;
	wire [4-1:0] node27805;
	wire [4-1:0] node27808;
	wire [4-1:0] node27811;
	wire [4-1:0] node27812;
	wire [4-1:0] node27813;
	wire [4-1:0] node27816;
	wire [4-1:0] node27818;
	wire [4-1:0] node27821;
	wire [4-1:0] node27822;
	wire [4-1:0] node27824;
	wire [4-1:0] node27827;
	wire [4-1:0] node27829;
	wire [4-1:0] node27832;
	wire [4-1:0] node27833;
	wire [4-1:0] node27834;
	wire [4-1:0] node27835;
	wire [4-1:0] node27836;
	wire [4-1:0] node27839;
	wire [4-1:0] node27842;
	wire [4-1:0] node27843;
	wire [4-1:0] node27846;
	wire [4-1:0] node27849;
	wire [4-1:0] node27850;
	wire [4-1:0] node27851;
	wire [4-1:0] node27853;
	wire [4-1:0] node27856;
	wire [4-1:0] node27857;
	wire [4-1:0] node27861;
	wire [4-1:0] node27862;
	wire [4-1:0] node27865;
	wire [4-1:0] node27866;
	wire [4-1:0] node27869;
	wire [4-1:0] node27872;
	wire [4-1:0] node27873;
	wire [4-1:0] node27874;
	wire [4-1:0] node27876;
	wire [4-1:0] node27879;
	wire [4-1:0] node27882;
	wire [4-1:0] node27883;
	wire [4-1:0] node27885;
	wire [4-1:0] node27886;
	wire [4-1:0] node27889;
	wire [4-1:0] node27892;
	wire [4-1:0] node27893;
	wire [4-1:0] node27896;
	wire [4-1:0] node27899;
	wire [4-1:0] node27900;
	wire [4-1:0] node27901;
	wire [4-1:0] node27902;
	wire [4-1:0] node27903;
	wire [4-1:0] node27905;
	wire [4-1:0] node27906;
	wire [4-1:0] node27909;
	wire [4-1:0] node27912;
	wire [4-1:0] node27913;
	wire [4-1:0] node27915;
	wire [4-1:0] node27919;
	wire [4-1:0] node27920;
	wire [4-1:0] node27921;
	wire [4-1:0] node27922;
	wire [4-1:0] node27926;
	wire [4-1:0] node27927;
	wire [4-1:0] node27930;
	wire [4-1:0] node27934;
	wire [4-1:0] node27935;
	wire [4-1:0] node27936;
	wire [4-1:0] node27938;
	wire [4-1:0] node27941;
	wire [4-1:0] node27942;
	wire [4-1:0] node27943;
	wire [4-1:0] node27946;
	wire [4-1:0] node27950;
	wire [4-1:0] node27951;
	wire [4-1:0] node27952;
	wire [4-1:0] node27953;
	wire [4-1:0] node27958;
	wire [4-1:0] node27959;
	wire [4-1:0] node27963;
	wire [4-1:0] node27964;
	wire [4-1:0] node27965;
	wire [4-1:0] node27966;
	wire [4-1:0] node27967;
	wire [4-1:0] node27968;
	wire [4-1:0] node27971;
	wire [4-1:0] node27975;
	wire [4-1:0] node27976;
	wire [4-1:0] node27977;
	wire [4-1:0] node27981;
	wire [4-1:0] node27983;
	wire [4-1:0] node27986;
	wire [4-1:0] node27987;
	wire [4-1:0] node27988;
	wire [4-1:0] node27989;
	wire [4-1:0] node27992;
	wire [4-1:0] node27996;
	wire [4-1:0] node27997;
	wire [4-1:0] node27998;
	wire [4-1:0] node28001;
	wire [4-1:0] node28004;
	wire [4-1:0] node28006;
	wire [4-1:0] node28009;
	wire [4-1:0] node28010;
	wire [4-1:0] node28011;
	wire [4-1:0] node28012;
	wire [4-1:0] node28013;
	wire [4-1:0] node28016;
	wire [4-1:0] node28020;
	wire [4-1:0] node28021;
	wire [4-1:0] node28023;
	wire [4-1:0] node28027;
	wire [4-1:0] node28028;
	wire [4-1:0] node28029;
	wire [4-1:0] node28032;
	wire [4-1:0] node28034;
	wire [4-1:0] node28037;
	wire [4-1:0] node28038;
	wire [4-1:0] node28039;
	wire [4-1:0] node28042;
	wire [4-1:0] node28045;
	wire [4-1:0] node28046;
	wire [4-1:0] node28050;
	wire [4-1:0] node28051;
	wire [4-1:0] node28052;
	wire [4-1:0] node28053;
	wire [4-1:0] node28054;
	wire [4-1:0] node28055;
	wire [4-1:0] node28056;
	wire [4-1:0] node28057;
	wire [4-1:0] node28058;
	wire [4-1:0] node28060;
	wire [4-1:0] node28064;
	wire [4-1:0] node28067;
	wire [4-1:0] node28068;
	wire [4-1:0] node28070;
	wire [4-1:0] node28071;
	wire [4-1:0] node28075;
	wire [4-1:0] node28076;
	wire [4-1:0] node28079;
	wire [4-1:0] node28082;
	wire [4-1:0] node28083;
	wire [4-1:0] node28084;
	wire [4-1:0] node28086;
	wire [4-1:0] node28087;
	wire [4-1:0] node28091;
	wire [4-1:0] node28093;
	wire [4-1:0] node28096;
	wire [4-1:0] node28097;
	wire [4-1:0] node28099;
	wire [4-1:0] node28101;
	wire [4-1:0] node28104;
	wire [4-1:0] node28106;
	wire [4-1:0] node28109;
	wire [4-1:0] node28110;
	wire [4-1:0] node28111;
	wire [4-1:0] node28112;
	wire [4-1:0] node28113;
	wire [4-1:0] node28117;
	wire [4-1:0] node28118;
	wire [4-1:0] node28122;
	wire [4-1:0] node28123;
	wire [4-1:0] node28124;
	wire [4-1:0] node28125;
	wire [4-1:0] node28129;
	wire [4-1:0] node28130;
	wire [4-1:0] node28133;
	wire [4-1:0] node28136;
	wire [4-1:0] node28137;
	wire [4-1:0] node28138;
	wire [4-1:0] node28143;
	wire [4-1:0] node28144;
	wire [4-1:0] node28145;
	wire [4-1:0] node28147;
	wire [4-1:0] node28148;
	wire [4-1:0] node28151;
	wire [4-1:0] node28154;
	wire [4-1:0] node28155;
	wire [4-1:0] node28156;
	wire [4-1:0] node28159;
	wire [4-1:0] node28163;
	wire [4-1:0] node28164;
	wire [4-1:0] node28165;
	wire [4-1:0] node28166;
	wire [4-1:0] node28169;
	wire [4-1:0] node28173;
	wire [4-1:0] node28174;
	wire [4-1:0] node28177;
	wire [4-1:0] node28180;
	wire [4-1:0] node28181;
	wire [4-1:0] node28182;
	wire [4-1:0] node28183;
	wire [4-1:0] node28184;
	wire [4-1:0] node28185;
	wire [4-1:0] node28187;
	wire [4-1:0] node28190;
	wire [4-1:0] node28192;
	wire [4-1:0] node28196;
	wire [4-1:0] node28197;
	wire [4-1:0] node28199;
	wire [4-1:0] node28202;
	wire [4-1:0] node28203;
	wire [4-1:0] node28204;
	wire [4-1:0] node28208;
	wire [4-1:0] node28211;
	wire [4-1:0] node28212;
	wire [4-1:0] node28213;
	wire [4-1:0] node28216;
	wire [4-1:0] node28217;
	wire [4-1:0] node28221;
	wire [4-1:0] node28222;
	wire [4-1:0] node28223;
	wire [4-1:0] node28224;
	wire [4-1:0] node28228;
	wire [4-1:0] node28230;
	wire [4-1:0] node28233;
	wire [4-1:0] node28234;
	wire [4-1:0] node28235;
	wire [4-1:0] node28238;
	wire [4-1:0] node28242;
	wire [4-1:0] node28243;
	wire [4-1:0] node28244;
	wire [4-1:0] node28245;
	wire [4-1:0] node28246;
	wire [4-1:0] node28247;
	wire [4-1:0] node28250;
	wire [4-1:0] node28254;
	wire [4-1:0] node28255;
	wire [4-1:0] node28257;
	wire [4-1:0] node28260;
	wire [4-1:0] node28262;
	wire [4-1:0] node28265;
	wire [4-1:0] node28266;
	wire [4-1:0] node28267;
	wire [4-1:0] node28268;
	wire [4-1:0] node28271;
	wire [4-1:0] node28274;
	wire [4-1:0] node28276;
	wire [4-1:0] node28279;
	wire [4-1:0] node28280;
	wire [4-1:0] node28283;
	wire [4-1:0] node28286;
	wire [4-1:0] node28287;
	wire [4-1:0] node28288;
	wire [4-1:0] node28289;
	wire [4-1:0] node28290;
	wire [4-1:0] node28294;
	wire [4-1:0] node28295;
	wire [4-1:0] node28299;
	wire [4-1:0] node28300;
	wire [4-1:0] node28301;
	wire [4-1:0] node28305;
	wire [4-1:0] node28306;
	wire [4-1:0] node28309;
	wire [4-1:0] node28312;
	wire [4-1:0] node28313;
	wire [4-1:0] node28314;
	wire [4-1:0] node28316;
	wire [4-1:0] node28320;
	wire [4-1:0] node28322;
	wire [4-1:0] node28324;
	wire [4-1:0] node28327;
	wire [4-1:0] node28328;
	wire [4-1:0] node28329;
	wire [4-1:0] node28330;
	wire [4-1:0] node28331;
	wire [4-1:0] node28332;
	wire [4-1:0] node28333;
	wire [4-1:0] node28335;
	wire [4-1:0] node28338;
	wire [4-1:0] node28339;
	wire [4-1:0] node28342;
	wire [4-1:0] node28345;
	wire [4-1:0] node28347;
	wire [4-1:0] node28348;
	wire [4-1:0] node28351;
	wire [4-1:0] node28354;
	wire [4-1:0] node28355;
	wire [4-1:0] node28356;
	wire [4-1:0] node28357;
	wire [4-1:0] node28360;
	wire [4-1:0] node28364;
	wire [4-1:0] node28365;
	wire [4-1:0] node28366;
	wire [4-1:0] node28369;
	wire [4-1:0] node28373;
	wire [4-1:0] node28374;
	wire [4-1:0] node28375;
	wire [4-1:0] node28377;
	wire [4-1:0] node28378;
	wire [4-1:0] node28381;
	wire [4-1:0] node28384;
	wire [4-1:0] node28385;
	wire [4-1:0] node28387;
	wire [4-1:0] node28390;
	wire [4-1:0] node28393;
	wire [4-1:0] node28394;
	wire [4-1:0] node28395;
	wire [4-1:0] node28397;
	wire [4-1:0] node28400;
	wire [4-1:0] node28401;
	wire [4-1:0] node28405;
	wire [4-1:0] node28406;
	wire [4-1:0] node28410;
	wire [4-1:0] node28411;
	wire [4-1:0] node28412;
	wire [4-1:0] node28413;
	wire [4-1:0] node28414;
	wire [4-1:0] node28416;
	wire [4-1:0] node28419;
	wire [4-1:0] node28421;
	wire [4-1:0] node28425;
	wire [4-1:0] node28426;
	wire [4-1:0] node28427;
	wire [4-1:0] node28430;
	wire [4-1:0] node28433;
	wire [4-1:0] node28434;
	wire [4-1:0] node28437;
	wire [4-1:0] node28440;
	wire [4-1:0] node28441;
	wire [4-1:0] node28442;
	wire [4-1:0] node28443;
	wire [4-1:0] node28445;
	wire [4-1:0] node28448;
	wire [4-1:0] node28451;
	wire [4-1:0] node28452;
	wire [4-1:0] node28455;
	wire [4-1:0] node28456;
	wire [4-1:0] node28460;
	wire [4-1:0] node28461;
	wire [4-1:0] node28464;
	wire [4-1:0] node28466;
	wire [4-1:0] node28467;
	wire [4-1:0] node28471;
	wire [4-1:0] node28472;
	wire [4-1:0] node28473;
	wire [4-1:0] node28474;
	wire [4-1:0] node28475;
	wire [4-1:0] node28476;
	wire [4-1:0] node28479;
	wire [4-1:0] node28481;
	wire [4-1:0] node28484;
	wire [4-1:0] node28485;
	wire [4-1:0] node28486;
	wire [4-1:0] node28490;
	wire [4-1:0] node28491;
	wire [4-1:0] node28494;
	wire [4-1:0] node28497;
	wire [4-1:0] node28498;
	wire [4-1:0] node28499;
	wire [4-1:0] node28502;
	wire [4-1:0] node28505;
	wire [4-1:0] node28506;
	wire [4-1:0] node28507;
	wire [4-1:0] node28510;
	wire [4-1:0] node28513;
	wire [4-1:0] node28514;
	wire [4-1:0] node28518;
	wire [4-1:0] node28519;
	wire [4-1:0] node28520;
	wire [4-1:0] node28521;
	wire [4-1:0] node28522;
	wire [4-1:0] node28526;
	wire [4-1:0] node28529;
	wire [4-1:0] node28531;
	wire [4-1:0] node28534;
	wire [4-1:0] node28535;
	wire [4-1:0] node28536;
	wire [4-1:0] node28538;
	wire [4-1:0] node28541;
	wire [4-1:0] node28542;
	wire [4-1:0] node28545;
	wire [4-1:0] node28548;
	wire [4-1:0] node28549;
	wire [4-1:0] node28552;
	wire [4-1:0] node28555;
	wire [4-1:0] node28556;
	wire [4-1:0] node28557;
	wire [4-1:0] node28558;
	wire [4-1:0] node28560;
	wire [4-1:0] node28561;
	wire [4-1:0] node28564;
	wire [4-1:0] node28567;
	wire [4-1:0] node28569;
	wire [4-1:0] node28570;
	wire [4-1:0] node28574;
	wire [4-1:0] node28575;
	wire [4-1:0] node28576;
	wire [4-1:0] node28580;
	wire [4-1:0] node28581;
	wire [4-1:0] node28585;
	wire [4-1:0] node28586;
	wire [4-1:0] node28587;
	wire [4-1:0] node28589;
	wire [4-1:0] node28592;
	wire [4-1:0] node28593;
	wire [4-1:0] node28597;
	wire [4-1:0] node28598;
	wire [4-1:0] node28600;
	wire [4-1:0] node28603;
	wire [4-1:0] node28604;
	wire [4-1:0] node28605;
	wire [4-1:0] node28608;
	wire [4-1:0] node28612;
	wire [4-1:0] node28613;
	wire [4-1:0] node28614;
	wire [4-1:0] node28615;
	wire [4-1:0] node28616;
	wire [4-1:0] node28617;
	wire [4-1:0] node28618;
	wire [4-1:0] node28619;
	wire [4-1:0] node28620;
	wire [4-1:0] node28623;
	wire [4-1:0] node28627;
	wire [4-1:0] node28628;
	wire [4-1:0] node28629;
	wire [4-1:0] node28633;
	wire [4-1:0] node28634;
	wire [4-1:0] node28637;
	wire [4-1:0] node28640;
	wire [4-1:0] node28641;
	wire [4-1:0] node28642;
	wire [4-1:0] node28643;
	wire [4-1:0] node28646;
	wire [4-1:0] node28650;
	wire [4-1:0] node28651;
	wire [4-1:0] node28652;
	wire [4-1:0] node28656;
	wire [4-1:0] node28658;
	wire [4-1:0] node28661;
	wire [4-1:0] node28662;
	wire [4-1:0] node28663;
	wire [4-1:0] node28664;
	wire [4-1:0] node28668;
	wire [4-1:0] node28669;
	wire [4-1:0] node28670;
	wire [4-1:0] node28674;
	wire [4-1:0] node28675;
	wire [4-1:0] node28678;
	wire [4-1:0] node28681;
	wire [4-1:0] node28682;
	wire [4-1:0] node28684;
	wire [4-1:0] node28687;
	wire [4-1:0] node28688;
	wire [4-1:0] node28691;
	wire [4-1:0] node28694;
	wire [4-1:0] node28695;
	wire [4-1:0] node28696;
	wire [4-1:0] node28697;
	wire [4-1:0] node28699;
	wire [4-1:0] node28702;
	wire [4-1:0] node28703;
	wire [4-1:0] node28705;
	wire [4-1:0] node28709;
	wire [4-1:0] node28710;
	wire [4-1:0] node28711;
	wire [4-1:0] node28712;
	wire [4-1:0] node28715;
	wire [4-1:0] node28719;
	wire [4-1:0] node28720;
	wire [4-1:0] node28722;
	wire [4-1:0] node28725;
	wire [4-1:0] node28728;
	wire [4-1:0] node28729;
	wire [4-1:0] node28730;
	wire [4-1:0] node28732;
	wire [4-1:0] node28734;
	wire [4-1:0] node28737;
	wire [4-1:0] node28738;
	wire [4-1:0] node28739;
	wire [4-1:0] node28742;
	wire [4-1:0] node28745;
	wire [4-1:0] node28748;
	wire [4-1:0] node28749;
	wire [4-1:0] node28750;
	wire [4-1:0] node28754;
	wire [4-1:0] node28755;
	wire [4-1:0] node28758;
	wire [4-1:0] node28761;
	wire [4-1:0] node28762;
	wire [4-1:0] node28763;
	wire [4-1:0] node28764;
	wire [4-1:0] node28765;
	wire [4-1:0] node28767;
	wire [4-1:0] node28768;
	wire [4-1:0] node28772;
	wire [4-1:0] node28773;
	wire [4-1:0] node28774;
	wire [4-1:0] node28777;
	wire [4-1:0] node28780;
	wire [4-1:0] node28782;
	wire [4-1:0] node28785;
	wire [4-1:0] node28786;
	wire [4-1:0] node28787;
	wire [4-1:0] node28788;
	wire [4-1:0] node28792;
	wire [4-1:0] node28793;
	wire [4-1:0] node28797;
	wire [4-1:0] node28798;
	wire [4-1:0] node28800;
	wire [4-1:0] node28803;
	wire [4-1:0] node28804;
	wire [4-1:0] node28807;
	wire [4-1:0] node28810;
	wire [4-1:0] node28811;
	wire [4-1:0] node28812;
	wire [4-1:0] node28813;
	wire [4-1:0] node28814;
	wire [4-1:0] node28817;
	wire [4-1:0] node28821;
	wire [4-1:0] node28822;
	wire [4-1:0] node28823;
	wire [4-1:0] node28826;
	wire [4-1:0] node28829;
	wire [4-1:0] node28831;
	wire [4-1:0] node28834;
	wire [4-1:0] node28835;
	wire [4-1:0] node28839;
	wire [4-1:0] node28840;
	wire [4-1:0] node28841;
	wire [4-1:0] node28842;
	wire [4-1:0] node28843;
	wire [4-1:0] node28845;
	wire [4-1:0] node28848;
	wire [4-1:0] node28849;
	wire [4-1:0] node28852;
	wire [4-1:0] node28856;
	wire [4-1:0] node28857;
	wire [4-1:0] node28859;
	wire [4-1:0] node28862;
	wire [4-1:0] node28863;
	wire [4-1:0] node28865;
	wire [4-1:0] node28869;
	wire [4-1:0] node28870;
	wire [4-1:0] node28871;
	wire [4-1:0] node28872;
	wire [4-1:0] node28873;
	wire [4-1:0] node28876;
	wire [4-1:0] node28879;
	wire [4-1:0] node28882;
	wire [4-1:0] node28883;
	wire [4-1:0] node28884;
	wire [4-1:0] node28888;
	wire [4-1:0] node28889;
	wire [4-1:0] node28892;
	wire [4-1:0] node28895;
	wire [4-1:0] node28896;
	wire [4-1:0] node28897;
	wire [4-1:0] node28898;
	wire [4-1:0] node28901;
	wire [4-1:0] node28905;
	wire [4-1:0] node28906;
	wire [4-1:0] node28907;
	wire [4-1:0] node28910;
	wire [4-1:0] node28914;
	wire [4-1:0] node28915;
	wire [4-1:0] node28916;
	wire [4-1:0] node28917;
	wire [4-1:0] node28918;
	wire [4-1:0] node28919;
	wire [4-1:0] node28921;
	wire [4-1:0] node28924;
	wire [4-1:0] node28926;
	wire [4-1:0] node28929;
	wire [4-1:0] node28930;
	wire [4-1:0] node28933;
	wire [4-1:0] node28934;
	wire [4-1:0] node28936;
	wire [4-1:0] node28940;
	wire [4-1:0] node28941;
	wire [4-1:0] node28942;
	wire [4-1:0] node28944;
	wire [4-1:0] node28947;
	wire [4-1:0] node28949;
	wire [4-1:0] node28952;
	wire [4-1:0] node28953;
	wire [4-1:0] node28955;
	wire [4-1:0] node28958;
	wire [4-1:0] node28960;
	wire [4-1:0] node28963;
	wire [4-1:0] node28964;
	wire [4-1:0] node28965;
	wire [4-1:0] node28966;
	wire [4-1:0] node28967;
	wire [4-1:0] node28972;
	wire [4-1:0] node28973;
	wire [4-1:0] node28974;
	wire [4-1:0] node28978;
	wire [4-1:0] node28979;
	wire [4-1:0] node28981;
	wire [4-1:0] node28985;
	wire [4-1:0] node28986;
	wire [4-1:0] node28987;
	wire [4-1:0] node28988;
	wire [4-1:0] node28991;
	wire [4-1:0] node28994;
	wire [4-1:0] node28995;
	wire [4-1:0] node28996;
	wire [4-1:0] node28999;
	wire [4-1:0] node29002;
	wire [4-1:0] node29003;
	wire [4-1:0] node29007;
	wire [4-1:0] node29008;
	wire [4-1:0] node29010;
	wire [4-1:0] node29013;
	wire [4-1:0] node29014;
	wire [4-1:0] node29017;
	wire [4-1:0] node29020;
	wire [4-1:0] node29021;
	wire [4-1:0] node29022;
	wire [4-1:0] node29023;
	wire [4-1:0] node29024;
	wire [4-1:0] node29027;
	wire [4-1:0] node29030;
	wire [4-1:0] node29031;
	wire [4-1:0] node29032;
	wire [4-1:0] node29034;
	wire [4-1:0] node29038;
	wire [4-1:0] node29040;
	wire [4-1:0] node29043;
	wire [4-1:0] node29044;
	wire [4-1:0] node29045;
	wire [4-1:0] node29046;
	wire [4-1:0] node29047;
	wire [4-1:0] node29052;
	wire [4-1:0] node29054;
	wire [4-1:0] node29055;
	wire [4-1:0] node29059;
	wire [4-1:0] node29060;
	wire [4-1:0] node29062;
	wire [4-1:0] node29065;
	wire [4-1:0] node29067;
	wire [4-1:0] node29068;
	wire [4-1:0] node29071;
	wire [4-1:0] node29074;
	wire [4-1:0] node29075;
	wire [4-1:0] node29076;
	wire [4-1:0] node29077;
	wire [4-1:0] node29078;
	wire [4-1:0] node29081;
	wire [4-1:0] node29084;
	wire [4-1:0] node29085;
	wire [4-1:0] node29087;
	wire [4-1:0] node29091;
	wire [4-1:0] node29092;
	wire [4-1:0] node29094;
	wire [4-1:0] node29097;
	wire [4-1:0] node29098;
	wire [4-1:0] node29099;
	wire [4-1:0] node29102;
	wire [4-1:0] node29106;
	wire [4-1:0] node29107;
	wire [4-1:0] node29108;
	wire [4-1:0] node29109;
	wire [4-1:0] node29112;
	wire [4-1:0] node29116;
	wire [4-1:0] node29117;
	wire [4-1:0] node29118;
	wire [4-1:0] node29121;
	wire [4-1:0] node29124;
	wire [4-1:0] node29125;
	wire [4-1:0] node29128;
	wire [4-1:0] node29131;
	wire [4-1:0] node29132;
	wire [4-1:0] node29133;
	wire [4-1:0] node29134;
	wire [4-1:0] node29135;
	wire [4-1:0] node29136;
	wire [4-1:0] node29137;
	wire [4-1:0] node29138;
	wire [4-1:0] node29139;
	wire [4-1:0] node29140;
	wire [4-1:0] node29143;
	wire [4-1:0] node29146;
	wire [4-1:0] node29147;
	wire [4-1:0] node29150;
	wire [4-1:0] node29153;
	wire [4-1:0] node29154;
	wire [4-1:0] node29156;
	wire [4-1:0] node29157;
	wire [4-1:0] node29160;
	wire [4-1:0] node29163;
	wire [4-1:0] node29164;
	wire [4-1:0] node29165;
	wire [4-1:0] node29170;
	wire [4-1:0] node29171;
	wire [4-1:0] node29172;
	wire [4-1:0] node29173;
	wire [4-1:0] node29177;
	wire [4-1:0] node29178;
	wire [4-1:0] node29182;
	wire [4-1:0] node29183;
	wire [4-1:0] node29187;
	wire [4-1:0] node29188;
	wire [4-1:0] node29189;
	wire [4-1:0] node29190;
	wire [4-1:0] node29192;
	wire [4-1:0] node29193;
	wire [4-1:0] node29198;
	wire [4-1:0] node29199;
	wire [4-1:0] node29202;
	wire [4-1:0] node29205;
	wire [4-1:0] node29206;
	wire [4-1:0] node29207;
	wire [4-1:0] node29208;
	wire [4-1:0] node29209;
	wire [4-1:0] node29213;
	wire [4-1:0] node29214;
	wire [4-1:0] node29218;
	wire [4-1:0] node29219;
	wire [4-1:0] node29220;
	wire [4-1:0] node29224;
	wire [4-1:0] node29225;
	wire [4-1:0] node29229;
	wire [4-1:0] node29230;
	wire [4-1:0] node29231;
	wire [4-1:0] node29232;
	wire [4-1:0] node29236;
	wire [4-1:0] node29237;
	wire [4-1:0] node29241;
	wire [4-1:0] node29244;
	wire [4-1:0] node29245;
	wire [4-1:0] node29246;
	wire [4-1:0] node29247;
	wire [4-1:0] node29248;
	wire [4-1:0] node29249;
	wire [4-1:0] node29250;
	wire [4-1:0] node29256;
	wire [4-1:0] node29257;
	wire [4-1:0] node29258;
	wire [4-1:0] node29262;
	wire [4-1:0] node29265;
	wire [4-1:0] node29266;
	wire [4-1:0] node29267;
	wire [4-1:0] node29268;
	wire [4-1:0] node29273;
	wire [4-1:0] node29274;
	wire [4-1:0] node29276;
	wire [4-1:0] node29277;
	wire [4-1:0] node29280;
	wire [4-1:0] node29283;
	wire [4-1:0] node29284;
	wire [4-1:0] node29287;
	wire [4-1:0] node29290;
	wire [4-1:0] node29291;
	wire [4-1:0] node29292;
	wire [4-1:0] node29293;
	wire [4-1:0] node29295;
	wire [4-1:0] node29297;
	wire [4-1:0] node29300;
	wire [4-1:0] node29301;
	wire [4-1:0] node29304;
	wire [4-1:0] node29305;
	wire [4-1:0] node29309;
	wire [4-1:0] node29310;
	wire [4-1:0] node29311;
	wire [4-1:0] node29315;
	wire [4-1:0] node29318;
	wire [4-1:0] node29319;
	wire [4-1:0] node29320;
	wire [4-1:0] node29322;
	wire [4-1:0] node29324;
	wire [4-1:0] node29327;
	wire [4-1:0] node29328;
	wire [4-1:0] node29329;
	wire [4-1:0] node29334;
	wire [4-1:0] node29335;
	wire [4-1:0] node29337;
	wire [4-1:0] node29338;
	wire [4-1:0] node29342;
	wire [4-1:0] node29343;
	wire [4-1:0] node29344;
	wire [4-1:0] node29348;
	wire [4-1:0] node29349;
	wire [4-1:0] node29352;
	wire [4-1:0] node29355;
	wire [4-1:0] node29356;
	wire [4-1:0] node29357;
	wire [4-1:0] node29358;
	wire [4-1:0] node29359;
	wire [4-1:0] node29360;
	wire [4-1:0] node29362;
	wire [4-1:0] node29366;
	wire [4-1:0] node29367;
	wire [4-1:0] node29368;
	wire [4-1:0] node29369;
	wire [4-1:0] node29372;
	wire [4-1:0] node29375;
	wire [4-1:0] node29376;
	wire [4-1:0] node29379;
	wire [4-1:0] node29382;
	wire [4-1:0] node29383;
	wire [4-1:0] node29386;
	wire [4-1:0] node29389;
	wire [4-1:0] node29390;
	wire [4-1:0] node29391;
	wire [4-1:0] node29393;
	wire [4-1:0] node29396;
	wire [4-1:0] node29397;
	wire [4-1:0] node29398;
	wire [4-1:0] node29403;
	wire [4-1:0] node29404;
	wire [4-1:0] node29405;
	wire [4-1:0] node29408;
	wire [4-1:0] node29411;
	wire [4-1:0] node29414;
	wire [4-1:0] node29415;
	wire [4-1:0] node29416;
	wire [4-1:0] node29417;
	wire [4-1:0] node29418;
	wire [4-1:0] node29421;
	wire [4-1:0] node29424;
	wire [4-1:0] node29425;
	wire [4-1:0] node29429;
	wire [4-1:0] node29430;
	wire [4-1:0] node29433;
	wire [4-1:0] node29434;
	wire [4-1:0] node29438;
	wire [4-1:0] node29439;
	wire [4-1:0] node29440;
	wire [4-1:0] node29442;
	wire [4-1:0] node29445;
	wire [4-1:0] node29446;
	wire [4-1:0] node29447;
	wire [4-1:0] node29451;
	wire [4-1:0] node29454;
	wire [4-1:0] node29455;
	wire [4-1:0] node29456;
	wire [4-1:0] node29458;
	wire [4-1:0] node29461;
	wire [4-1:0] node29462;
	wire [4-1:0] node29467;
	wire [4-1:0] node29468;
	wire [4-1:0] node29469;
	wire [4-1:0] node29470;
	wire [4-1:0] node29471;
	wire [4-1:0] node29472;
	wire [4-1:0] node29473;
	wire [4-1:0] node29477;
	wire [4-1:0] node29478;
	wire [4-1:0] node29482;
	wire [4-1:0] node29484;
	wire [4-1:0] node29487;
	wire [4-1:0] node29488;
	wire [4-1:0] node29489;
	wire [4-1:0] node29491;
	wire [4-1:0] node29495;
	wire [4-1:0] node29496;
	wire [4-1:0] node29499;
	wire [4-1:0] node29502;
	wire [4-1:0] node29503;
	wire [4-1:0] node29505;
	wire [4-1:0] node29506;
	wire [4-1:0] node29510;
	wire [4-1:0] node29511;
	wire [4-1:0] node29512;
	wire [4-1:0] node29513;
	wire [4-1:0] node29516;
	wire [4-1:0] node29520;
	wire [4-1:0] node29522;
	wire [4-1:0] node29523;
	wire [4-1:0] node29526;
	wire [4-1:0] node29529;
	wire [4-1:0] node29530;
	wire [4-1:0] node29531;
	wire [4-1:0] node29532;
	wire [4-1:0] node29533;
	wire [4-1:0] node29534;
	wire [4-1:0] node29537;
	wire [4-1:0] node29541;
	wire [4-1:0] node29542;
	wire [4-1:0] node29543;
	wire [4-1:0] node29546;
	wire [4-1:0] node29549;
	wire [4-1:0] node29550;
	wire [4-1:0] node29554;
	wire [4-1:0] node29555;
	wire [4-1:0] node29556;
	wire [4-1:0] node29558;
	wire [4-1:0] node29562;
	wire [4-1:0] node29563;
	wire [4-1:0] node29566;
	wire [4-1:0] node29567;
	wire [4-1:0] node29571;
	wire [4-1:0] node29572;
	wire [4-1:0] node29573;
	wire [4-1:0] node29574;
	wire [4-1:0] node29575;
	wire [4-1:0] node29578;
	wire [4-1:0] node29581;
	wire [4-1:0] node29583;
	wire [4-1:0] node29586;
	wire [4-1:0] node29588;
	wire [4-1:0] node29591;
	wire [4-1:0] node29593;
	wire [4-1:0] node29594;
	wire [4-1:0] node29597;
	wire [4-1:0] node29600;
	wire [4-1:0] node29601;
	wire [4-1:0] node29602;
	wire [4-1:0] node29603;
	wire [4-1:0] node29604;
	wire [4-1:0] node29605;
	wire [4-1:0] node29606;
	wire [4-1:0] node29607;
	wire [4-1:0] node29610;
	wire [4-1:0] node29613;
	wire [4-1:0] node29614;
	wire [4-1:0] node29617;
	wire [4-1:0] node29620;
	wire [4-1:0] node29621;
	wire [4-1:0] node29622;
	wire [4-1:0] node29623;
	wire [4-1:0] node29627;
	wire [4-1:0] node29628;
	wire [4-1:0] node29631;
	wire [4-1:0] node29634;
	wire [4-1:0] node29635;
	wire [4-1:0] node29636;
	wire [4-1:0] node29640;
	wire [4-1:0] node29642;
	wire [4-1:0] node29645;
	wire [4-1:0] node29646;
	wire [4-1:0] node29647;
	wire [4-1:0] node29649;
	wire [4-1:0] node29652;
	wire [4-1:0] node29655;
	wire [4-1:0] node29656;
	wire [4-1:0] node29657;
	wire [4-1:0] node29660;
	wire [4-1:0] node29663;
	wire [4-1:0] node29664;
	wire [4-1:0] node29667;
	wire [4-1:0] node29670;
	wire [4-1:0] node29671;
	wire [4-1:0] node29672;
	wire [4-1:0] node29673;
	wire [4-1:0] node29674;
	wire [4-1:0] node29675;
	wire [4-1:0] node29678;
	wire [4-1:0] node29681;
	wire [4-1:0] node29683;
	wire [4-1:0] node29686;
	wire [4-1:0] node29687;
	wire [4-1:0] node29689;
	wire [4-1:0] node29692;
	wire [4-1:0] node29694;
	wire [4-1:0] node29697;
	wire [4-1:0] node29698;
	wire [4-1:0] node29699;
	wire [4-1:0] node29701;
	wire [4-1:0] node29705;
	wire [4-1:0] node29707;
	wire [4-1:0] node29710;
	wire [4-1:0] node29711;
	wire [4-1:0] node29712;
	wire [4-1:0] node29713;
	wire [4-1:0] node29714;
	wire [4-1:0] node29718;
	wire [4-1:0] node29719;
	wire [4-1:0] node29723;
	wire [4-1:0] node29725;
	wire [4-1:0] node29728;
	wire [4-1:0] node29729;
	wire [4-1:0] node29731;
	wire [4-1:0] node29735;
	wire [4-1:0] node29736;
	wire [4-1:0] node29737;
	wire [4-1:0] node29738;
	wire [4-1:0] node29739;
	wire [4-1:0] node29741;
	wire [4-1:0] node29742;
	wire [4-1:0] node29745;
	wire [4-1:0] node29748;
	wire [4-1:0] node29750;
	wire [4-1:0] node29751;
	wire [4-1:0] node29755;
	wire [4-1:0] node29756;
	wire [4-1:0] node29759;
	wire [4-1:0] node29762;
	wire [4-1:0] node29763;
	wire [4-1:0] node29764;
	wire [4-1:0] node29765;
	wire [4-1:0] node29769;
	wire [4-1:0] node29770;
	wire [4-1:0] node29773;
	wire [4-1:0] node29776;
	wire [4-1:0] node29777;
	wire [4-1:0] node29778;
	wire [4-1:0] node29782;
	wire [4-1:0] node29783;
	wire [4-1:0] node29784;
	wire [4-1:0] node29787;
	wire [4-1:0] node29791;
	wire [4-1:0] node29792;
	wire [4-1:0] node29793;
	wire [4-1:0] node29795;
	wire [4-1:0] node29796;
	wire [4-1:0] node29799;
	wire [4-1:0] node29802;
	wire [4-1:0] node29803;
	wire [4-1:0] node29804;
	wire [4-1:0] node29805;
	wire [4-1:0] node29809;
	wire [4-1:0] node29812;
	wire [4-1:0] node29814;
	wire [4-1:0] node29817;
	wire [4-1:0] node29818;
	wire [4-1:0] node29819;
	wire [4-1:0] node29820;
	wire [4-1:0] node29822;
	wire [4-1:0] node29825;
	wire [4-1:0] node29827;
	wire [4-1:0] node29830;
	wire [4-1:0] node29831;
	wire [4-1:0] node29834;
	wire [4-1:0] node29837;
	wire [4-1:0] node29838;
	wire [4-1:0] node29841;
	wire [4-1:0] node29843;
	wire [4-1:0] node29846;
	wire [4-1:0] node29847;
	wire [4-1:0] node29848;
	wire [4-1:0] node29849;
	wire [4-1:0] node29850;
	wire [4-1:0] node29851;
	wire [4-1:0] node29853;
	wire [4-1:0] node29855;
	wire [4-1:0] node29858;
	wire [4-1:0] node29859;
	wire [4-1:0] node29863;
	wire [4-1:0] node29864;
	wire [4-1:0] node29865;
	wire [4-1:0] node29867;
	wire [4-1:0] node29870;
	wire [4-1:0] node29873;
	wire [4-1:0] node29874;
	wire [4-1:0] node29877;
	wire [4-1:0] node29880;
	wire [4-1:0] node29881;
	wire [4-1:0] node29882;
	wire [4-1:0] node29883;
	wire [4-1:0] node29885;
	wire [4-1:0] node29889;
	wire [4-1:0] node29891;
	wire [4-1:0] node29894;
	wire [4-1:0] node29895;
	wire [4-1:0] node29896;
	wire [4-1:0] node29897;
	wire [4-1:0] node29901;
	wire [4-1:0] node29904;
	wire [4-1:0] node29906;
	wire [4-1:0] node29909;
	wire [4-1:0] node29910;
	wire [4-1:0] node29911;
	wire [4-1:0] node29912;
	wire [4-1:0] node29913;
	wire [4-1:0] node29915;
	wire [4-1:0] node29918;
	wire [4-1:0] node29919;
	wire [4-1:0] node29923;
	wire [4-1:0] node29925;
	wire [4-1:0] node29928;
	wire [4-1:0] node29929;
	wire [4-1:0] node29932;
	wire [4-1:0] node29934;
	wire [4-1:0] node29935;
	wire [4-1:0] node29939;
	wire [4-1:0] node29940;
	wire [4-1:0] node29941;
	wire [4-1:0] node29942;
	wire [4-1:0] node29943;
	wire [4-1:0] node29947;
	wire [4-1:0] node29948;
	wire [4-1:0] node29951;
	wire [4-1:0] node29954;
	wire [4-1:0] node29956;
	wire [4-1:0] node29959;
	wire [4-1:0] node29961;
	wire [4-1:0] node29962;
	wire [4-1:0] node29963;
	wire [4-1:0] node29968;
	wire [4-1:0] node29969;
	wire [4-1:0] node29970;
	wire [4-1:0] node29971;
	wire [4-1:0] node29972;
	wire [4-1:0] node29973;
	wire [4-1:0] node29975;
	wire [4-1:0] node29978;
	wire [4-1:0] node29980;
	wire [4-1:0] node29983;
	wire [4-1:0] node29984;
	wire [4-1:0] node29987;
	wire [4-1:0] node29988;
	wire [4-1:0] node29992;
	wire [4-1:0] node29993;
	wire [4-1:0] node29994;
	wire [4-1:0] node29995;
	wire [4-1:0] node29999;
	wire [4-1:0] node30000;
	wire [4-1:0] node30004;
	wire [4-1:0] node30007;
	wire [4-1:0] node30008;
	wire [4-1:0] node30009;
	wire [4-1:0] node30010;
	wire [4-1:0] node30014;
	wire [4-1:0] node30015;
	wire [4-1:0] node30019;
	wire [4-1:0] node30020;
	wire [4-1:0] node30021;
	wire [4-1:0] node30024;
	wire [4-1:0] node30028;
	wire [4-1:0] node30029;
	wire [4-1:0] node30030;
	wire [4-1:0] node30031;
	wire [4-1:0] node30032;
	wire [4-1:0] node30033;
	wire [4-1:0] node30036;
	wire [4-1:0] node30039;
	wire [4-1:0] node30040;
	wire [4-1:0] node30044;
	wire [4-1:0] node30046;
	wire [4-1:0] node30049;
	wire [4-1:0] node30050;
	wire [4-1:0] node30052;
	wire [4-1:0] node30055;
	wire [4-1:0] node30056;
	wire [4-1:0] node30057;
	wire [4-1:0] node30060;
	wire [4-1:0] node30063;
	wire [4-1:0] node30064;
	wire [4-1:0] node30068;
	wire [4-1:0] node30069;
	wire [4-1:0] node30070;
	wire [4-1:0] node30072;
	wire [4-1:0] node30075;
	wire [4-1:0] node30076;
	wire [4-1:0] node30079;
	wire [4-1:0] node30082;
	wire [4-1:0] node30083;
	wire [4-1:0] node30084;
	wire [4-1:0] node30085;
	wire [4-1:0] node30089;
	wire [4-1:0] node30090;
	wire [4-1:0] node30094;
	wire [4-1:0] node30095;
	wire [4-1:0] node30099;
	wire [4-1:0] node30100;
	wire [4-1:0] node30101;
	wire [4-1:0] node30102;
	wire [4-1:0] node30103;
	wire [4-1:0] node30104;
	wire [4-1:0] node30105;
	wire [4-1:0] node30106;
	wire [4-1:0] node30107;
	wire [4-1:0] node30108;
	wire [4-1:0] node30111;
	wire [4-1:0] node30114;
	wire [4-1:0] node30116;
	wire [4-1:0] node30119;
	wire [4-1:0] node30120;
	wire [4-1:0] node30121;
	wire [4-1:0] node30124;
	wire [4-1:0] node30128;
	wire [4-1:0] node30129;
	wire [4-1:0] node30130;
	wire [4-1:0] node30131;
	wire [4-1:0] node30134;
	wire [4-1:0] node30138;
	wire [4-1:0] node30141;
	wire [4-1:0] node30142;
	wire [4-1:0] node30143;
	wire [4-1:0] node30146;
	wire [4-1:0] node30147;
	wire [4-1:0] node30150;
	wire [4-1:0] node30153;
	wire [4-1:0] node30154;
	wire [4-1:0] node30156;
	wire [4-1:0] node30157;
	wire [4-1:0] node30160;
	wire [4-1:0] node30163;
	wire [4-1:0] node30164;
	wire [4-1:0] node30166;
	wire [4-1:0] node30170;
	wire [4-1:0] node30171;
	wire [4-1:0] node30172;
	wire [4-1:0] node30173;
	wire [4-1:0] node30174;
	wire [4-1:0] node30175;
	wire [4-1:0] node30180;
	wire [4-1:0] node30181;
	wire [4-1:0] node30183;
	wire [4-1:0] node30186;
	wire [4-1:0] node30187;
	wire [4-1:0] node30190;
	wire [4-1:0] node30193;
	wire [4-1:0] node30194;
	wire [4-1:0] node30195;
	wire [4-1:0] node30196;
	wire [4-1:0] node30200;
	wire [4-1:0] node30201;
	wire [4-1:0] node30205;
	wire [4-1:0] node30207;
	wire [4-1:0] node30208;
	wire [4-1:0] node30211;
	wire [4-1:0] node30214;
	wire [4-1:0] node30215;
	wire [4-1:0] node30216;
	wire [4-1:0] node30217;
	wire [4-1:0] node30219;
	wire [4-1:0] node30223;
	wire [4-1:0] node30224;
	wire [4-1:0] node30226;
	wire [4-1:0] node30230;
	wire [4-1:0] node30231;
	wire [4-1:0] node30233;
	wire [4-1:0] node30234;
	wire [4-1:0] node30237;
	wire [4-1:0] node30240;
	wire [4-1:0] node30241;
	wire [4-1:0] node30244;
	wire [4-1:0] node30245;
	wire [4-1:0] node30249;
	wire [4-1:0] node30250;
	wire [4-1:0] node30251;
	wire [4-1:0] node30252;
	wire [4-1:0] node30254;
	wire [4-1:0] node30255;
	wire [4-1:0] node30257;
	wire [4-1:0] node30261;
	wire [4-1:0] node30262;
	wire [4-1:0] node30263;
	wire [4-1:0] node30266;
	wire [4-1:0] node30269;
	wire [4-1:0] node30271;
	wire [4-1:0] node30274;
	wire [4-1:0] node30275;
	wire [4-1:0] node30276;
	wire [4-1:0] node30277;
	wire [4-1:0] node30278;
	wire [4-1:0] node30283;
	wire [4-1:0] node30284;
	wire [4-1:0] node30286;
	wire [4-1:0] node30289;
	wire [4-1:0] node30291;
	wire [4-1:0] node30294;
	wire [4-1:0] node30295;
	wire [4-1:0] node30296;
	wire [4-1:0] node30298;
	wire [4-1:0] node30301;
	wire [4-1:0] node30302;
	wire [4-1:0] node30305;
	wire [4-1:0] node30308;
	wire [4-1:0] node30309;
	wire [4-1:0] node30310;
	wire [4-1:0] node30313;
	wire [4-1:0] node30317;
	wire [4-1:0] node30318;
	wire [4-1:0] node30319;
	wire [4-1:0] node30320;
	wire [4-1:0] node30321;
	wire [4-1:0] node30322;
	wire [4-1:0] node30327;
	wire [4-1:0] node30329;
	wire [4-1:0] node30331;
	wire [4-1:0] node30334;
	wire [4-1:0] node30335;
	wire [4-1:0] node30337;
	wire [4-1:0] node30338;
	wire [4-1:0] node30342;
	wire [4-1:0] node30343;
	wire [4-1:0] node30345;
	wire [4-1:0] node30349;
	wire [4-1:0] node30350;
	wire [4-1:0] node30351;
	wire [4-1:0] node30352;
	wire [4-1:0] node30356;
	wire [4-1:0] node30357;
	wire [4-1:0] node30358;
	wire [4-1:0] node30362;
	wire [4-1:0] node30363;
	wire [4-1:0] node30366;
	wire [4-1:0] node30369;
	wire [4-1:0] node30370;
	wire [4-1:0] node30371;
	wire [4-1:0] node30373;
	wire [4-1:0] node30377;
	wire [4-1:0] node30379;
	wire [4-1:0] node30380;
	wire [4-1:0] node30383;
	wire [4-1:0] node30386;
	wire [4-1:0] node30387;
	wire [4-1:0] node30388;
	wire [4-1:0] node30389;
	wire [4-1:0] node30390;
	wire [4-1:0] node30391;
	wire [4-1:0] node30392;
	wire [4-1:0] node30394;
	wire [4-1:0] node30398;
	wire [4-1:0] node30399;
	wire [4-1:0] node30401;
	wire [4-1:0] node30404;
	wire [4-1:0] node30406;
	wire [4-1:0] node30409;
	wire [4-1:0] node30410;
	wire [4-1:0] node30411;
	wire [4-1:0] node30412;
	wire [4-1:0] node30416;
	wire [4-1:0] node30417;
	wire [4-1:0] node30420;
	wire [4-1:0] node30423;
	wire [4-1:0] node30425;
	wire [4-1:0] node30426;
	wire [4-1:0] node30429;
	wire [4-1:0] node30432;
	wire [4-1:0] node30433;
	wire [4-1:0] node30434;
	wire [4-1:0] node30435;
	wire [4-1:0] node30437;
	wire [4-1:0] node30441;
	wire [4-1:0] node30443;
	wire [4-1:0] node30446;
	wire [4-1:0] node30447;
	wire [4-1:0] node30449;
	wire [4-1:0] node30451;
	wire [4-1:0] node30454;
	wire [4-1:0] node30455;
	wire [4-1:0] node30456;
	wire [4-1:0] node30460;
	wire [4-1:0] node30461;
	wire [4-1:0] node30465;
	wire [4-1:0] node30466;
	wire [4-1:0] node30467;
	wire [4-1:0] node30468;
	wire [4-1:0] node30471;
	wire [4-1:0] node30472;
	wire [4-1:0] node30473;
	wire [4-1:0] node30476;
	wire [4-1:0] node30480;
	wire [4-1:0] node30481;
	wire [4-1:0] node30482;
	wire [4-1:0] node30483;
	wire [4-1:0] node30487;
	wire [4-1:0] node30488;
	wire [4-1:0] node30491;
	wire [4-1:0] node30494;
	wire [4-1:0] node30495;
	wire [4-1:0] node30496;
	wire [4-1:0] node30499;
	wire [4-1:0] node30503;
	wire [4-1:0] node30504;
	wire [4-1:0] node30505;
	wire [4-1:0] node30506;
	wire [4-1:0] node30507;
	wire [4-1:0] node30510;
	wire [4-1:0] node30514;
	wire [4-1:0] node30515;
	wire [4-1:0] node30517;
	wire [4-1:0] node30520;
	wire [4-1:0] node30521;
	wire [4-1:0] node30525;
	wire [4-1:0] node30526;
	wire [4-1:0] node30527;
	wire [4-1:0] node30530;
	wire [4-1:0] node30531;
	wire [4-1:0] node30535;
	wire [4-1:0] node30537;
	wire [4-1:0] node30540;
	wire [4-1:0] node30541;
	wire [4-1:0] node30542;
	wire [4-1:0] node30543;
	wire [4-1:0] node30544;
	wire [4-1:0] node30545;
	wire [4-1:0] node30546;
	wire [4-1:0] node30551;
	wire [4-1:0] node30552;
	wire [4-1:0] node30553;
	wire [4-1:0] node30558;
	wire [4-1:0] node30559;
	wire [4-1:0] node30561;
	wire [4-1:0] node30563;
	wire [4-1:0] node30566;
	wire [4-1:0] node30568;
	wire [4-1:0] node30570;
	wire [4-1:0] node30573;
	wire [4-1:0] node30574;
	wire [4-1:0] node30575;
	wire [4-1:0] node30576;
	wire [4-1:0] node30577;
	wire [4-1:0] node30580;
	wire [4-1:0] node30584;
	wire [4-1:0] node30586;
	wire [4-1:0] node30588;
	wire [4-1:0] node30591;
	wire [4-1:0] node30592;
	wire [4-1:0] node30593;
	wire [4-1:0] node30594;
	wire [4-1:0] node30598;
	wire [4-1:0] node30600;
	wire [4-1:0] node30603;
	wire [4-1:0] node30605;
	wire [4-1:0] node30607;
	wire [4-1:0] node30610;
	wire [4-1:0] node30611;
	wire [4-1:0] node30612;
	wire [4-1:0] node30613;
	wire [4-1:0] node30615;
	wire [4-1:0] node30616;
	wire [4-1:0] node30619;
	wire [4-1:0] node30622;
	wire [4-1:0] node30624;
	wire [4-1:0] node30626;
	wire [4-1:0] node30629;
	wire [4-1:0] node30630;
	wire [4-1:0] node30631;
	wire [4-1:0] node30633;
	wire [4-1:0] node30636;
	wire [4-1:0] node30639;
	wire [4-1:0] node30640;
	wire [4-1:0] node30643;
	wire [4-1:0] node30646;
	wire [4-1:0] node30647;
	wire [4-1:0] node30648;
	wire [4-1:0] node30649;
	wire [4-1:0] node30650;
	wire [4-1:0] node30653;
	wire [4-1:0] node30656;
	wire [4-1:0] node30657;
	wire [4-1:0] node30660;
	wire [4-1:0] node30663;
	wire [4-1:0] node30664;
	wire [4-1:0] node30665;
	wire [4-1:0] node30668;
	wire [4-1:0] node30672;
	wire [4-1:0] node30673;
	wire [4-1:0] node30674;
	wire [4-1:0] node30675;
	wire [4-1:0] node30678;
	wire [4-1:0] node30682;
	wire [4-1:0] node30683;
	wire [4-1:0] node30687;
	wire [4-1:0] node30688;
	wire [4-1:0] node30689;
	wire [4-1:0] node30690;
	wire [4-1:0] node30691;
	wire [4-1:0] node30692;
	wire [4-1:0] node30693;
	wire [4-1:0] node30694;
	wire [4-1:0] node30695;
	wire [4-1:0] node30699;
	wire [4-1:0] node30701;
	wire [4-1:0] node30704;
	wire [4-1:0] node30706;
	wire [4-1:0] node30707;
	wire [4-1:0] node30710;
	wire [4-1:0] node30713;
	wire [4-1:0] node30714;
	wire [4-1:0] node30717;
	wire [4-1:0] node30718;
	wire [4-1:0] node30719;
	wire [4-1:0] node30723;
	wire [4-1:0] node30725;
	wire [4-1:0] node30728;
	wire [4-1:0] node30729;
	wire [4-1:0] node30730;
	wire [4-1:0] node30731;
	wire [4-1:0] node30735;
	wire [4-1:0] node30737;
	wire [4-1:0] node30740;
	wire [4-1:0] node30741;
	wire [4-1:0] node30742;
	wire [4-1:0] node30743;
	wire [4-1:0] node30746;
	wire [4-1:0] node30749;
	wire [4-1:0] node30750;
	wire [4-1:0] node30753;
	wire [4-1:0] node30756;
	wire [4-1:0] node30757;
	wire [4-1:0] node30760;
	wire [4-1:0] node30763;
	wire [4-1:0] node30764;
	wire [4-1:0] node30765;
	wire [4-1:0] node30766;
	wire [4-1:0] node30768;
	wire [4-1:0] node30771;
	wire [4-1:0] node30772;
	wire [4-1:0] node30773;
	wire [4-1:0] node30776;
	wire [4-1:0] node30780;
	wire [4-1:0] node30781;
	wire [4-1:0] node30784;
	wire [4-1:0] node30785;
	wire [4-1:0] node30789;
	wire [4-1:0] node30790;
	wire [4-1:0] node30791;
	wire [4-1:0] node30794;
	wire [4-1:0] node30795;
	wire [4-1:0] node30798;
	wire [4-1:0] node30801;
	wire [4-1:0] node30803;
	wire [4-1:0] node30806;
	wire [4-1:0] node30807;
	wire [4-1:0] node30808;
	wire [4-1:0] node30809;
	wire [4-1:0] node30810;
	wire [4-1:0] node30811;
	wire [4-1:0] node30816;
	wire [4-1:0] node30817;
	wire [4-1:0] node30819;
	wire [4-1:0] node30822;
	wire [4-1:0] node30823;
	wire [4-1:0] node30826;
	wire [4-1:0] node30829;
	wire [4-1:0] node30830;
	wire [4-1:0] node30831;
	wire [4-1:0] node30832;
	wire [4-1:0] node30834;
	wire [4-1:0] node30838;
	wire [4-1:0] node30839;
	wire [4-1:0] node30841;
	wire [4-1:0] node30844;
	wire [4-1:0] node30845;
	wire [4-1:0] node30848;
	wire [4-1:0] node30851;
	wire [4-1:0] node30852;
	wire [4-1:0] node30855;
	wire [4-1:0] node30856;
	wire [4-1:0] node30859;
	wire [4-1:0] node30862;
	wire [4-1:0] node30863;
	wire [4-1:0] node30864;
	wire [4-1:0] node30865;
	wire [4-1:0] node30867;
	wire [4-1:0] node30870;
	wire [4-1:0] node30871;
	wire [4-1:0] node30874;
	wire [4-1:0] node30877;
	wire [4-1:0] node30878;
	wire [4-1:0] node30879;
	wire [4-1:0] node30882;
	wire [4-1:0] node30885;
	wire [4-1:0] node30887;
	wire [4-1:0] node30890;
	wire [4-1:0] node30891;
	wire [4-1:0] node30892;
	wire [4-1:0] node30893;
	wire [4-1:0] node30897;
	wire [4-1:0] node30899;
	wire [4-1:0] node30902;
	wire [4-1:0] node30903;
	wire [4-1:0] node30905;
	wire [4-1:0] node30907;
	wire [4-1:0] node30910;
	wire [4-1:0] node30911;
	wire [4-1:0] node30912;
	wire [4-1:0] node30917;
	wire [4-1:0] node30918;
	wire [4-1:0] node30919;
	wire [4-1:0] node30920;
	wire [4-1:0] node30921;
	wire [4-1:0] node30922;
	wire [4-1:0] node30923;
	wire [4-1:0] node30926;
	wire [4-1:0] node30929;
	wire [4-1:0] node30930;
	wire [4-1:0] node30932;
	wire [4-1:0] node30935;
	wire [4-1:0] node30936;
	wire [4-1:0] node30939;
	wire [4-1:0] node30942;
	wire [4-1:0] node30943;
	wire [4-1:0] node30944;
	wire [4-1:0] node30947;
	wire [4-1:0] node30950;
	wire [4-1:0] node30953;
	wire [4-1:0] node30954;
	wire [4-1:0] node30955;
	wire [4-1:0] node30956;
	wire [4-1:0] node30959;
	wire [4-1:0] node30962;
	wire [4-1:0] node30964;
	wire [4-1:0] node30965;
	wire [4-1:0] node30969;
	wire [4-1:0] node30970;
	wire [4-1:0] node30971;
	wire [4-1:0] node30972;
	wire [4-1:0] node30975;
	wire [4-1:0] node30978;
	wire [4-1:0] node30979;
	wire [4-1:0] node30983;
	wire [4-1:0] node30985;
	wire [4-1:0] node30988;
	wire [4-1:0] node30989;
	wire [4-1:0] node30990;
	wire [4-1:0] node30991;
	wire [4-1:0] node30992;
	wire [4-1:0] node30995;
	wire [4-1:0] node30998;
	wire [4-1:0] node30999;
	wire [4-1:0] node31002;
	wire [4-1:0] node31005;
	wire [4-1:0] node31006;
	wire [4-1:0] node31007;
	wire [4-1:0] node31008;
	wire [4-1:0] node31011;
	wire [4-1:0] node31014;
	wire [4-1:0] node31015;
	wire [4-1:0] node31018;
	wire [4-1:0] node31021;
	wire [4-1:0] node31022;
	wire [4-1:0] node31024;
	wire [4-1:0] node31027;
	wire [4-1:0] node31028;
	wire [4-1:0] node31032;
	wire [4-1:0] node31033;
	wire [4-1:0] node31036;
	wire [4-1:0] node31037;
	wire [4-1:0] node31038;
	wire [4-1:0] node31039;
	wire [4-1:0] node31043;
	wire [4-1:0] node31045;
	wire [4-1:0] node31048;
	wire [4-1:0] node31051;
	wire [4-1:0] node31052;
	wire [4-1:0] node31053;
	wire [4-1:0] node31054;
	wire [4-1:0] node31055;
	wire [4-1:0] node31056;
	wire [4-1:0] node31057;
	wire [4-1:0] node31060;
	wire [4-1:0] node31063;
	wire [4-1:0] node31065;
	wire [4-1:0] node31068;
	wire [4-1:0] node31070;
	wire [4-1:0] node31071;
	wire [4-1:0] node31074;
	wire [4-1:0] node31077;
	wire [4-1:0] node31078;
	wire [4-1:0] node31080;
	wire [4-1:0] node31083;
	wire [4-1:0] node31085;
	wire [4-1:0] node31086;
	wire [4-1:0] node31089;
	wire [4-1:0] node31092;
	wire [4-1:0] node31093;
	wire [4-1:0] node31094;
	wire [4-1:0] node31095;
	wire [4-1:0] node31099;
	wire [4-1:0] node31100;
	wire [4-1:0] node31102;
	wire [4-1:0] node31105;
	wire [4-1:0] node31107;
	wire [4-1:0] node31110;
	wire [4-1:0] node31111;
	wire [4-1:0] node31112;
	wire [4-1:0] node31115;
	wire [4-1:0] node31118;
	wire [4-1:0] node31119;
	wire [4-1:0] node31121;
	wire [4-1:0] node31124;
	wire [4-1:0] node31126;
	wire [4-1:0] node31129;
	wire [4-1:0] node31130;
	wire [4-1:0] node31131;
	wire [4-1:0] node31132;
	wire [4-1:0] node31134;
	wire [4-1:0] node31137;
	wire [4-1:0] node31138;
	wire [4-1:0] node31141;
	wire [4-1:0] node31144;
	wire [4-1:0] node31145;
	wire [4-1:0] node31146;
	wire [4-1:0] node31147;
	wire [4-1:0] node31152;
	wire [4-1:0] node31153;
	wire [4-1:0] node31154;
	wire [4-1:0] node31157;
	wire [4-1:0] node31160;
	wire [4-1:0] node31161;
	wire [4-1:0] node31165;
	wire [4-1:0] node31166;
	wire [4-1:0] node31167;
	wire [4-1:0] node31168;
	wire [4-1:0] node31172;
	wire [4-1:0] node31173;
	wire [4-1:0] node31176;
	wire [4-1:0] node31179;
	wire [4-1:0] node31180;
	wire [4-1:0] node31181;
	wire [4-1:0] node31184;
	wire [4-1:0] node31187;
	wire [4-1:0] node31189;
	wire [4-1:0] node31192;
	wire [4-1:0] node31193;
	wire [4-1:0] node31194;
	wire [4-1:0] node31195;
	wire [4-1:0] node31196;
	wire [4-1:0] node31197;
	wire [4-1:0] node31198;
	wire [4-1:0] node31199;
	wire [4-1:0] node31200;
	wire [4-1:0] node31201;
	wire [4-1:0] node31202;
	wire [4-1:0] node31203;
	wire [4-1:0] node31204;
	wire [4-1:0] node31206;
	wire [4-1:0] node31207;
	wire [4-1:0] node31210;
	wire [4-1:0] node31213;
	wire [4-1:0] node31214;
	wire [4-1:0] node31217;
	wire [4-1:0] node31218;
	wire [4-1:0] node31221;
	wire [4-1:0] node31224;
	wire [4-1:0] node31225;
	wire [4-1:0] node31227;
	wire [4-1:0] node31229;
	wire [4-1:0] node31232;
	wire [4-1:0] node31233;
	wire [4-1:0] node31234;
	wire [4-1:0] node31237;
	wire [4-1:0] node31241;
	wire [4-1:0] node31242;
	wire [4-1:0] node31243;
	wire [4-1:0] node31244;
	wire [4-1:0] node31245;
	wire [4-1:0] node31248;
	wire [4-1:0] node31252;
	wire [4-1:0] node31253;
	wire [4-1:0] node31255;
	wire [4-1:0] node31258;
	wire [4-1:0] node31259;
	wire [4-1:0] node31262;
	wire [4-1:0] node31265;
	wire [4-1:0] node31266;
	wire [4-1:0] node31267;
	wire [4-1:0] node31269;
	wire [4-1:0] node31272;
	wire [4-1:0] node31273;
	wire [4-1:0] node31276;
	wire [4-1:0] node31279;
	wire [4-1:0] node31280;
	wire [4-1:0] node31284;
	wire [4-1:0] node31285;
	wire [4-1:0] node31286;
	wire [4-1:0] node31287;
	wire [4-1:0] node31288;
	wire [4-1:0] node31289;
	wire [4-1:0] node31293;
	wire [4-1:0] node31294;
	wire [4-1:0] node31298;
	wire [4-1:0] node31299;
	wire [4-1:0] node31300;
	wire [4-1:0] node31303;
	wire [4-1:0] node31306;
	wire [4-1:0] node31307;
	wire [4-1:0] node31311;
	wire [4-1:0] node31312;
	wire [4-1:0] node31314;
	wire [4-1:0] node31316;
	wire [4-1:0] node31319;
	wire [4-1:0] node31320;
	wire [4-1:0] node31322;
	wire [4-1:0] node31326;
	wire [4-1:0] node31327;
	wire [4-1:0] node31328;
	wire [4-1:0] node31329;
	wire [4-1:0] node31330;
	wire [4-1:0] node31333;
	wire [4-1:0] node31336;
	wire [4-1:0] node31338;
	wire [4-1:0] node31341;
	wire [4-1:0] node31343;
	wire [4-1:0] node31345;
	wire [4-1:0] node31348;
	wire [4-1:0] node31349;
	wire [4-1:0] node31350;
	wire [4-1:0] node31351;
	wire [4-1:0] node31354;
	wire [4-1:0] node31357;
	wire [4-1:0] node31359;
	wire [4-1:0] node31362;
	wire [4-1:0] node31363;
	wire [4-1:0] node31365;
	wire [4-1:0] node31368;
	wire [4-1:0] node31369;
	wire [4-1:0] node31373;
	wire [4-1:0] node31374;
	wire [4-1:0] node31375;
	wire [4-1:0] node31376;
	wire [4-1:0] node31377;
	wire [4-1:0] node31379;
	wire [4-1:0] node31380;
	wire [4-1:0] node31384;
	wire [4-1:0] node31386;
	wire [4-1:0] node31388;
	wire [4-1:0] node31391;
	wire [4-1:0] node31392;
	wire [4-1:0] node31393;
	wire [4-1:0] node31396;
	wire [4-1:0] node31399;
	wire [4-1:0] node31401;
	wire [4-1:0] node31402;
	wire [4-1:0] node31406;
	wire [4-1:0] node31407;
	wire [4-1:0] node31408;
	wire [4-1:0] node31409;
	wire [4-1:0] node31411;
	wire [4-1:0] node31414;
	wire [4-1:0] node31416;
	wire [4-1:0] node31419;
	wire [4-1:0] node31422;
	wire [4-1:0] node31423;
	wire [4-1:0] node31424;
	wire [4-1:0] node31428;
	wire [4-1:0] node31429;
	wire [4-1:0] node31432;
	wire [4-1:0] node31434;
	wire [4-1:0] node31437;
	wire [4-1:0] node31438;
	wire [4-1:0] node31439;
	wire [4-1:0] node31440;
	wire [4-1:0] node31442;
	wire [4-1:0] node31443;
	wire [4-1:0] node31446;
	wire [4-1:0] node31449;
	wire [4-1:0] node31451;
	wire [4-1:0] node31452;
	wire [4-1:0] node31455;
	wire [4-1:0] node31458;
	wire [4-1:0] node31460;
	wire [4-1:0] node31462;
	wire [4-1:0] node31464;
	wire [4-1:0] node31467;
	wire [4-1:0] node31468;
	wire [4-1:0] node31469;
	wire [4-1:0] node31470;
	wire [4-1:0] node31472;
	wire [4-1:0] node31476;
	wire [4-1:0] node31477;
	wire [4-1:0] node31478;
	wire [4-1:0] node31482;
	wire [4-1:0] node31483;
	wire [4-1:0] node31487;
	wire [4-1:0] node31488;
	wire [4-1:0] node31489;
	wire [4-1:0] node31491;
	wire [4-1:0] node31494;
	wire [4-1:0] node31495;
	wire [4-1:0] node31498;
	wire [4-1:0] node31501;
	wire [4-1:0] node31502;
	wire [4-1:0] node31504;
	wire [4-1:0] node31508;
	wire [4-1:0] node31509;
	wire [4-1:0] node31510;
	wire [4-1:0] node31511;
	wire [4-1:0] node31512;
	wire [4-1:0] node31513;
	wire [4-1:0] node31514;
	wire [4-1:0] node31516;
	wire [4-1:0] node31520;
	wire [4-1:0] node31521;
	wire [4-1:0] node31523;
	wire [4-1:0] node31526;
	wire [4-1:0] node31528;
	wire [4-1:0] node31531;
	wire [4-1:0] node31532;
	wire [4-1:0] node31533;
	wire [4-1:0] node31535;
	wire [4-1:0] node31538;
	wire [4-1:0] node31539;
	wire [4-1:0] node31542;
	wire [4-1:0] node31545;
	wire [4-1:0] node31548;
	wire [4-1:0] node31549;
	wire [4-1:0] node31550;
	wire [4-1:0] node31553;
	wire [4-1:0] node31554;
	wire [4-1:0] node31556;
	wire [4-1:0] node31559;
	wire [4-1:0] node31560;
	wire [4-1:0] node31564;
	wire [4-1:0] node31565;
	wire [4-1:0] node31566;
	wire [4-1:0] node31567;
	wire [4-1:0] node31572;
	wire [4-1:0] node31574;
	wire [4-1:0] node31577;
	wire [4-1:0] node31578;
	wire [4-1:0] node31579;
	wire [4-1:0] node31580;
	wire [4-1:0] node31581;
	wire [4-1:0] node31582;
	wire [4-1:0] node31585;
	wire [4-1:0] node31588;
	wire [4-1:0] node31590;
	wire [4-1:0] node31593;
	wire [4-1:0] node31594;
	wire [4-1:0] node31596;
	wire [4-1:0] node31599;
	wire [4-1:0] node31600;
	wire [4-1:0] node31604;
	wire [4-1:0] node31605;
	wire [4-1:0] node31606;
	wire [4-1:0] node31611;
	wire [4-1:0] node31612;
	wire [4-1:0] node31613;
	wire [4-1:0] node31614;
	wire [4-1:0] node31615;
	wire [4-1:0] node31618;
	wire [4-1:0] node31621;
	wire [4-1:0] node31622;
	wire [4-1:0] node31626;
	wire [4-1:0] node31628;
	wire [4-1:0] node31629;
	wire [4-1:0] node31632;
	wire [4-1:0] node31635;
	wire [4-1:0] node31636;
	wire [4-1:0] node31637;
	wire [4-1:0] node31638;
	wire [4-1:0] node31643;
	wire [4-1:0] node31644;
	wire [4-1:0] node31645;
	wire [4-1:0] node31648;
	wire [4-1:0] node31651;
	wire [4-1:0] node31652;
	wire [4-1:0] node31656;
	wire [4-1:0] node31657;
	wire [4-1:0] node31658;
	wire [4-1:0] node31659;
	wire [4-1:0] node31660;
	wire [4-1:0] node31663;
	wire [4-1:0] node31664;
	wire [4-1:0] node31666;
	wire [4-1:0] node31669;
	wire [4-1:0] node31670;
	wire [4-1:0] node31674;
	wire [4-1:0] node31675;
	wire [4-1:0] node31677;
	wire [4-1:0] node31678;
	wire [4-1:0] node31681;
	wire [4-1:0] node31685;
	wire [4-1:0] node31686;
	wire [4-1:0] node31687;
	wire [4-1:0] node31689;
	wire [4-1:0] node31690;
	wire [4-1:0] node31694;
	wire [4-1:0] node31696;
	wire [4-1:0] node31697;
	wire [4-1:0] node31700;
	wire [4-1:0] node31703;
	wire [4-1:0] node31704;
	wire [4-1:0] node31706;
	wire [4-1:0] node31707;
	wire [4-1:0] node31710;
	wire [4-1:0] node31713;
	wire [4-1:0] node31715;
	wire [4-1:0] node31716;
	wire [4-1:0] node31719;
	wire [4-1:0] node31722;
	wire [4-1:0] node31723;
	wire [4-1:0] node31724;
	wire [4-1:0] node31725;
	wire [4-1:0] node31726;
	wire [4-1:0] node31728;
	wire [4-1:0] node31731;
	wire [4-1:0] node31732;
	wire [4-1:0] node31735;
	wire [4-1:0] node31738;
	wire [4-1:0] node31740;
	wire [4-1:0] node31743;
	wire [4-1:0] node31744;
	wire [4-1:0] node31745;
	wire [4-1:0] node31746;
	wire [4-1:0] node31749;
	wire [4-1:0] node31752;
	wire [4-1:0] node31754;
	wire [4-1:0] node31757;
	wire [4-1:0] node31758;
	wire [4-1:0] node31759;
	wire [4-1:0] node31762;
	wire [4-1:0] node31765;
	wire [4-1:0] node31766;
	wire [4-1:0] node31769;
	wire [4-1:0] node31772;
	wire [4-1:0] node31773;
	wire [4-1:0] node31774;
	wire [4-1:0] node31776;
	wire [4-1:0] node31777;
	wire [4-1:0] node31780;
	wire [4-1:0] node31783;
	wire [4-1:0] node31784;
	wire [4-1:0] node31786;
	wire [4-1:0] node31789;
	wire [4-1:0] node31791;
	wire [4-1:0] node31794;
	wire [4-1:0] node31795;
	wire [4-1:0] node31796;
	wire [4-1:0] node31798;
	wire [4-1:0] node31802;
	wire [4-1:0] node31803;
	wire [4-1:0] node31804;
	wire [4-1:0] node31807;
	wire [4-1:0] node31810;
	wire [4-1:0] node31811;
	wire [4-1:0] node31815;
	wire [4-1:0] node31816;
	wire [4-1:0] node31817;
	wire [4-1:0] node31818;
	wire [4-1:0] node31819;
	wire [4-1:0] node31820;
	wire [4-1:0] node31822;
	wire [4-1:0] node31823;
	wire [4-1:0] node31826;
	wire [4-1:0] node31829;
	wire [4-1:0] node31830;
	wire [4-1:0] node31831;
	wire [4-1:0] node31834;
	wire [4-1:0] node31837;
	wire [4-1:0] node31838;
	wire [4-1:0] node31839;
	wire [4-1:0] node31844;
	wire [4-1:0] node31845;
	wire [4-1:0] node31846;
	wire [4-1:0] node31847;
	wire [4-1:0] node31851;
	wire [4-1:0] node31852;
	wire [4-1:0] node31855;
	wire [4-1:0] node31858;
	wire [4-1:0] node31859;
	wire [4-1:0] node31860;
	wire [4-1:0] node31862;
	wire [4-1:0] node31865;
	wire [4-1:0] node31867;
	wire [4-1:0] node31870;
	wire [4-1:0] node31871;
	wire [4-1:0] node31873;
	wire [4-1:0] node31876;
	wire [4-1:0] node31877;
	wire [4-1:0] node31881;
	wire [4-1:0] node31882;
	wire [4-1:0] node31883;
	wire [4-1:0] node31884;
	wire [4-1:0] node31886;
	wire [4-1:0] node31888;
	wire [4-1:0] node31891;
	wire [4-1:0] node31893;
	wire [4-1:0] node31894;
	wire [4-1:0] node31897;
	wire [4-1:0] node31900;
	wire [4-1:0] node31901;
	wire [4-1:0] node31902;
	wire [4-1:0] node31906;
	wire [4-1:0] node31907;
	wire [4-1:0] node31909;
	wire [4-1:0] node31912;
	wire [4-1:0] node31913;
	wire [4-1:0] node31916;
	wire [4-1:0] node31919;
	wire [4-1:0] node31920;
	wire [4-1:0] node31921;
	wire [4-1:0] node31923;
	wire [4-1:0] node31924;
	wire [4-1:0] node31927;
	wire [4-1:0] node31930;
	wire [4-1:0] node31932;
	wire [4-1:0] node31933;
	wire [4-1:0] node31936;
	wire [4-1:0] node31939;
	wire [4-1:0] node31940;
	wire [4-1:0] node31941;
	wire [4-1:0] node31945;
	wire [4-1:0] node31946;
	wire [4-1:0] node31947;
	wire [4-1:0] node31951;
	wire [4-1:0] node31952;
	wire [4-1:0] node31956;
	wire [4-1:0] node31957;
	wire [4-1:0] node31958;
	wire [4-1:0] node31959;
	wire [4-1:0] node31960;
	wire [4-1:0] node31961;
	wire [4-1:0] node31963;
	wire [4-1:0] node31966;
	wire [4-1:0] node31968;
	wire [4-1:0] node31971;
	wire [4-1:0] node31972;
	wire [4-1:0] node31973;
	wire [4-1:0] node31976;
	wire [4-1:0] node31979;
	wire [4-1:0] node31980;
	wire [4-1:0] node31984;
	wire [4-1:0] node31985;
	wire [4-1:0] node31986;
	wire [4-1:0] node31989;
	wire [4-1:0] node31991;
	wire [4-1:0] node31994;
	wire [4-1:0] node31996;
	wire [4-1:0] node31997;
	wire [4-1:0] node32001;
	wire [4-1:0] node32002;
	wire [4-1:0] node32003;
	wire [4-1:0] node32004;
	wire [4-1:0] node32006;
	wire [4-1:0] node32009;
	wire [4-1:0] node32010;
	wire [4-1:0] node32014;
	wire [4-1:0] node32015;
	wire [4-1:0] node32017;
	wire [4-1:0] node32020;
	wire [4-1:0] node32022;
	wire [4-1:0] node32025;
	wire [4-1:0] node32026;
	wire [4-1:0] node32028;
	wire [4-1:0] node32029;
	wire [4-1:0] node32033;
	wire [4-1:0] node32035;
	wire [4-1:0] node32036;
	wire [4-1:0] node32039;
	wire [4-1:0] node32042;
	wire [4-1:0] node32043;
	wire [4-1:0] node32044;
	wire [4-1:0] node32045;
	wire [4-1:0] node32046;
	wire [4-1:0] node32047;
	wire [4-1:0] node32050;
	wire [4-1:0] node32054;
	wire [4-1:0] node32055;
	wire [4-1:0] node32056;
	wire [4-1:0] node32060;
	wire [4-1:0] node32062;
	wire [4-1:0] node32065;
	wire [4-1:0] node32066;
	wire [4-1:0] node32067;
	wire [4-1:0] node32068;
	wire [4-1:0] node32072;
	wire [4-1:0] node32073;
	wire [4-1:0] node32077;
	wire [4-1:0] node32078;
	wire [4-1:0] node32079;
	wire [4-1:0] node32083;
	wire [4-1:0] node32084;
	wire [4-1:0] node32087;
	wire [4-1:0] node32090;
	wire [4-1:0] node32091;
	wire [4-1:0] node32092;
	wire [4-1:0] node32093;
	wire [4-1:0] node32094;
	wire [4-1:0] node32097;
	wire [4-1:0] node32100;
	wire [4-1:0] node32101;
	wire [4-1:0] node32104;
	wire [4-1:0] node32107;
	wire [4-1:0] node32108;
	wire [4-1:0] node32110;
	wire [4-1:0] node32113;
	wire [4-1:0] node32114;
	wire [4-1:0] node32117;
	wire [4-1:0] node32120;
	wire [4-1:0] node32121;
	wire [4-1:0] node32123;
	wire [4-1:0] node32126;
	wire [4-1:0] node32127;
	wire [4-1:0] node32128;
	wire [4-1:0] node32132;
	wire [4-1:0] node32135;
	wire [4-1:0] node32136;
	wire [4-1:0] node32137;
	wire [4-1:0] node32138;
	wire [4-1:0] node32139;
	wire [4-1:0] node32140;
	wire [4-1:0] node32141;
	wire [4-1:0] node32142;
	wire [4-1:0] node32145;
	wire [4-1:0] node32148;
	wire [4-1:0] node32151;
	wire [4-1:0] node32152;
	wire [4-1:0] node32153;
	wire [4-1:0] node32157;
	wire [4-1:0] node32160;
	wire [4-1:0] node32161;
	wire [4-1:0] node32164;
	wire [4-1:0] node32166;
	wire [4-1:0] node32167;
	wire [4-1:0] node32170;
	wire [4-1:0] node32173;
	wire [4-1:0] node32174;
	wire [4-1:0] node32175;
	wire [4-1:0] node32176;
	wire [4-1:0] node32177;
	wire [4-1:0] node32181;
	wire [4-1:0] node32182;
	wire [4-1:0] node32186;
	wire [4-1:0] node32187;
	wire [4-1:0] node32188;
	wire [4-1:0] node32193;
	wire [4-1:0] node32194;
	wire [4-1:0] node32195;
	wire [4-1:0] node32197;
	wire [4-1:0] node32200;
	wire [4-1:0] node32202;
	wire [4-1:0] node32205;
	wire [4-1:0] node32206;
	wire [4-1:0] node32207;
	wire [4-1:0] node32210;
	wire [4-1:0] node32214;
	wire [4-1:0] node32215;
	wire [4-1:0] node32216;
	wire [4-1:0] node32217;
	wire [4-1:0] node32219;
	wire [4-1:0] node32221;
	wire [4-1:0] node32224;
	wire [4-1:0] node32227;
	wire [4-1:0] node32228;
	wire [4-1:0] node32229;
	wire [4-1:0] node32231;
	wire [4-1:0] node32234;
	wire [4-1:0] node32236;
	wire [4-1:0] node32239;
	wire [4-1:0] node32240;
	wire [4-1:0] node32241;
	wire [4-1:0] node32244;
	wire [4-1:0] node32247;
	wire [4-1:0] node32248;
	wire [4-1:0] node32251;
	wire [4-1:0] node32254;
	wire [4-1:0] node32255;
	wire [4-1:0] node32256;
	wire [4-1:0] node32257;
	wire [4-1:0] node32259;
	wire [4-1:0] node32262;
	wire [4-1:0] node32265;
	wire [4-1:0] node32266;
	wire [4-1:0] node32267;
	wire [4-1:0] node32270;
	wire [4-1:0] node32274;
	wire [4-1:0] node32275;
	wire [4-1:0] node32276;
	wire [4-1:0] node32278;
	wire [4-1:0] node32281;
	wire [4-1:0] node32282;
	wire [4-1:0] node32285;
	wire [4-1:0] node32288;
	wire [4-1:0] node32289;
	wire [4-1:0] node32290;
	wire [4-1:0] node32294;
	wire [4-1:0] node32296;
	wire [4-1:0] node32299;
	wire [4-1:0] node32300;
	wire [4-1:0] node32301;
	wire [4-1:0] node32302;
	wire [4-1:0] node32303;
	wire [4-1:0] node32304;
	wire [4-1:0] node32305;
	wire [4-1:0] node32308;
	wire [4-1:0] node32311;
	wire [4-1:0] node32312;
	wire [4-1:0] node32315;
	wire [4-1:0] node32318;
	wire [4-1:0] node32319;
	wire [4-1:0] node32321;
	wire [4-1:0] node32324;
	wire [4-1:0] node32325;
	wire [4-1:0] node32328;
	wire [4-1:0] node32331;
	wire [4-1:0] node32332;
	wire [4-1:0] node32333;
	wire [4-1:0] node32334;
	wire [4-1:0] node32338;
	wire [4-1:0] node32340;
	wire [4-1:0] node32343;
	wire [4-1:0] node32344;
	wire [4-1:0] node32345;
	wire [4-1:0] node32349;
	wire [4-1:0] node32351;
	wire [4-1:0] node32354;
	wire [4-1:0] node32355;
	wire [4-1:0] node32356;
	wire [4-1:0] node32358;
	wire [4-1:0] node32359;
	wire [4-1:0] node32362;
	wire [4-1:0] node32365;
	wire [4-1:0] node32367;
	wire [4-1:0] node32370;
	wire [4-1:0] node32371;
	wire [4-1:0] node32373;
	wire [4-1:0] node32374;
	wire [4-1:0] node32378;
	wire [4-1:0] node32380;
	wire [4-1:0] node32382;
	wire [4-1:0] node32385;
	wire [4-1:0] node32386;
	wire [4-1:0] node32387;
	wire [4-1:0] node32388;
	wire [4-1:0] node32389;
	wire [4-1:0] node32390;
	wire [4-1:0] node32393;
	wire [4-1:0] node32397;
	wire [4-1:0] node32398;
	wire [4-1:0] node32400;
	wire [4-1:0] node32404;
	wire [4-1:0] node32405;
	wire [4-1:0] node32406;
	wire [4-1:0] node32410;
	wire [4-1:0] node32411;
	wire [4-1:0] node32415;
	wire [4-1:0] node32416;
	wire [4-1:0] node32417;
	wire [4-1:0] node32420;
	wire [4-1:0] node32423;
	wire [4-1:0] node32424;
	wire [4-1:0] node32425;
	wire [4-1:0] node32426;
	wire [4-1:0] node32429;
	wire [4-1:0] node32433;
	wire [4-1:0] node32434;
	wire [4-1:0] node32437;
	wire [4-1:0] node32439;
	wire [4-1:0] node32442;
	wire [4-1:0] node32443;
	wire [4-1:0] node32444;
	wire [4-1:0] node32445;
	wire [4-1:0] node32446;
	wire [4-1:0] node32447;
	wire [4-1:0] node32448;
	wire [4-1:0] node32449;
	wire [4-1:0] node32451;
	wire [4-1:0] node32452;
	wire [4-1:0] node32456;
	wire [4-1:0] node32457;
	wire [4-1:0] node32459;
	wire [4-1:0] node32462;
	wire [4-1:0] node32463;
	wire [4-1:0] node32466;
	wire [4-1:0] node32469;
	wire [4-1:0] node32470;
	wire [4-1:0] node32471;
	wire [4-1:0] node32472;
	wire [4-1:0] node32475;
	wire [4-1:0] node32478;
	wire [4-1:0] node32480;
	wire [4-1:0] node32483;
	wire [4-1:0] node32484;
	wire [4-1:0] node32486;
	wire [4-1:0] node32489;
	wire [4-1:0] node32490;
	wire [4-1:0] node32493;
	wire [4-1:0] node32496;
	wire [4-1:0] node32497;
	wire [4-1:0] node32498;
	wire [4-1:0] node32499;
	wire [4-1:0] node32500;
	wire [4-1:0] node32503;
	wire [4-1:0] node32506;
	wire [4-1:0] node32508;
	wire [4-1:0] node32512;
	wire [4-1:0] node32513;
	wire [4-1:0] node32514;
	wire [4-1:0] node32515;
	wire [4-1:0] node32518;
	wire [4-1:0] node32522;
	wire [4-1:0] node32523;
	wire [4-1:0] node32524;
	wire [4-1:0] node32527;
	wire [4-1:0] node32530;
	wire [4-1:0] node32531;
	wire [4-1:0] node32534;
	wire [4-1:0] node32537;
	wire [4-1:0] node32538;
	wire [4-1:0] node32539;
	wire [4-1:0] node32540;
	wire [4-1:0] node32541;
	wire [4-1:0] node32545;
	wire [4-1:0] node32547;
	wire [4-1:0] node32548;
	wire [4-1:0] node32551;
	wire [4-1:0] node32554;
	wire [4-1:0] node32555;
	wire [4-1:0] node32558;
	wire [4-1:0] node32559;
	wire [4-1:0] node32560;
	wire [4-1:0] node32563;
	wire [4-1:0] node32566;
	wire [4-1:0] node32569;
	wire [4-1:0] node32570;
	wire [4-1:0] node32571;
	wire [4-1:0] node32572;
	wire [4-1:0] node32573;
	wire [4-1:0] node32578;
	wire [4-1:0] node32579;
	wire [4-1:0] node32580;
	wire [4-1:0] node32583;
	wire [4-1:0] node32587;
	wire [4-1:0] node32588;
	wire [4-1:0] node32589;
	wire [4-1:0] node32590;
	wire [4-1:0] node32594;
	wire [4-1:0] node32595;
	wire [4-1:0] node32599;
	wire [4-1:0] node32600;
	wire [4-1:0] node32602;
	wire [4-1:0] node32606;
	wire [4-1:0] node32607;
	wire [4-1:0] node32608;
	wire [4-1:0] node32609;
	wire [4-1:0] node32610;
	wire [4-1:0] node32611;
	wire [4-1:0] node32612;
	wire [4-1:0] node32617;
	wire [4-1:0] node32618;
	wire [4-1:0] node32619;
	wire [4-1:0] node32623;
	wire [4-1:0] node32626;
	wire [4-1:0] node32627;
	wire [4-1:0] node32628;
	wire [4-1:0] node32629;
	wire [4-1:0] node32632;
	wire [4-1:0] node32635;
	wire [4-1:0] node32636;
	wire [4-1:0] node32639;
	wire [4-1:0] node32642;
	wire [4-1:0] node32643;
	wire [4-1:0] node32644;
	wire [4-1:0] node32648;
	wire [4-1:0] node32650;
	wire [4-1:0] node32653;
	wire [4-1:0] node32654;
	wire [4-1:0] node32655;
	wire [4-1:0] node32656;
	wire [4-1:0] node32659;
	wire [4-1:0] node32662;
	wire [4-1:0] node32664;
	wire [4-1:0] node32667;
	wire [4-1:0] node32668;
	wire [4-1:0] node32671;
	wire [4-1:0] node32672;
	wire [4-1:0] node32675;
	wire [4-1:0] node32678;
	wire [4-1:0] node32679;
	wire [4-1:0] node32680;
	wire [4-1:0] node32681;
	wire [4-1:0] node32682;
	wire [4-1:0] node32683;
	wire [4-1:0] node32686;
	wire [4-1:0] node32690;
	wire [4-1:0] node32691;
	wire [4-1:0] node32694;
	wire [4-1:0] node32697;
	wire [4-1:0] node32698;
	wire [4-1:0] node32699;
	wire [4-1:0] node32702;
	wire [4-1:0] node32706;
	wire [4-1:0] node32707;
	wire [4-1:0] node32708;
	wire [4-1:0] node32710;
	wire [4-1:0] node32712;
	wire [4-1:0] node32715;
	wire [4-1:0] node32717;
	wire [4-1:0] node32718;
	wire [4-1:0] node32722;
	wire [4-1:0] node32723;
	wire [4-1:0] node32724;
	wire [4-1:0] node32727;
	wire [4-1:0] node32730;
	wire [4-1:0] node32732;
	wire [4-1:0] node32733;
	wire [4-1:0] node32736;
	wire [4-1:0] node32739;
	wire [4-1:0] node32740;
	wire [4-1:0] node32741;
	wire [4-1:0] node32742;
	wire [4-1:0] node32743;
	wire [4-1:0] node32744;
	wire [4-1:0] node32745;
	wire [4-1:0] node32748;
	wire [4-1:0] node32751;
	wire [4-1:0] node32753;
	wire [4-1:0] node32756;
	wire [4-1:0] node32757;
	wire [4-1:0] node32758;
	wire [4-1:0] node32761;
	wire [4-1:0] node32764;
	wire [4-1:0] node32767;
	wire [4-1:0] node32768;
	wire [4-1:0] node32769;
	wire [4-1:0] node32770;
	wire [4-1:0] node32774;
	wire [4-1:0] node32775;
	wire [4-1:0] node32779;
	wire [4-1:0] node32780;
	wire [4-1:0] node32781;
	wire [4-1:0] node32785;
	wire [4-1:0] node32787;
	wire [4-1:0] node32788;
	wire [4-1:0] node32791;
	wire [4-1:0] node32794;
	wire [4-1:0] node32795;
	wire [4-1:0] node32796;
	wire [4-1:0] node32797;
	wire [4-1:0] node32798;
	wire [4-1:0] node32801;
	wire [4-1:0] node32802;
	wire [4-1:0] node32806;
	wire [4-1:0] node32809;
	wire [4-1:0] node32810;
	wire [4-1:0] node32812;
	wire [4-1:0] node32814;
	wire [4-1:0] node32817;
	wire [4-1:0] node32819;
	wire [4-1:0] node32820;
	wire [4-1:0] node32823;
	wire [4-1:0] node32826;
	wire [4-1:0] node32827;
	wire [4-1:0] node32828;
	wire [4-1:0] node32830;
	wire [4-1:0] node32833;
	wire [4-1:0] node32834;
	wire [4-1:0] node32835;
	wire [4-1:0] node32839;
	wire [4-1:0] node32842;
	wire [4-1:0] node32843;
	wire [4-1:0] node32844;
	wire [4-1:0] node32847;
	wire [4-1:0] node32850;
	wire [4-1:0] node32851;
	wire [4-1:0] node32854;
	wire [4-1:0] node32857;
	wire [4-1:0] node32858;
	wire [4-1:0] node32859;
	wire [4-1:0] node32860;
	wire [4-1:0] node32862;
	wire [4-1:0] node32863;
	wire [4-1:0] node32866;
	wire [4-1:0] node32869;
	wire [4-1:0] node32870;
	wire [4-1:0] node32871;
	wire [4-1:0] node32874;
	wire [4-1:0] node32877;
	wire [4-1:0] node32878;
	wire [4-1:0] node32882;
	wire [4-1:0] node32883;
	wire [4-1:0] node32884;
	wire [4-1:0] node32886;
	wire [4-1:0] node32888;
	wire [4-1:0] node32891;
	wire [4-1:0] node32892;
	wire [4-1:0] node32893;
	wire [4-1:0] node32897;
	wire [4-1:0] node32898;
	wire [4-1:0] node32901;
	wire [4-1:0] node32904;
	wire [4-1:0] node32905;
	wire [4-1:0] node32906;
	wire [4-1:0] node32907;
	wire [4-1:0] node32910;
	wire [4-1:0] node32914;
	wire [4-1:0] node32917;
	wire [4-1:0] node32918;
	wire [4-1:0] node32919;
	wire [4-1:0] node32921;
	wire [4-1:0] node32922;
	wire [4-1:0] node32925;
	wire [4-1:0] node32928;
	wire [4-1:0] node32929;
	wire [4-1:0] node32932;
	wire [4-1:0] node32933;
	wire [4-1:0] node32934;
	wire [4-1:0] node32937;
	wire [4-1:0] node32941;
	wire [4-1:0] node32942;
	wire [4-1:0] node32943;
	wire [4-1:0] node32945;
	wire [4-1:0] node32946;
	wire [4-1:0] node32949;
	wire [4-1:0] node32953;
	wire [4-1:0] node32954;
	wire [4-1:0] node32957;
	wire [4-1:0] node32958;
	wire [4-1:0] node32961;
	wire [4-1:0] node32964;
	wire [4-1:0] node32965;
	wire [4-1:0] node32966;
	wire [4-1:0] node32967;
	wire [4-1:0] node32968;
	wire [4-1:0] node32969;
	wire [4-1:0] node32970;
	wire [4-1:0] node32971;
	wire [4-1:0] node32974;
	wire [4-1:0] node32977;
	wire [4-1:0] node32978;
	wire [4-1:0] node32981;
	wire [4-1:0] node32984;
	wire [4-1:0] node32985;
	wire [4-1:0] node32986;
	wire [4-1:0] node32989;
	wire [4-1:0] node32992;
	wire [4-1:0] node32993;
	wire [4-1:0] node32994;
	wire [4-1:0] node32998;
	wire [4-1:0] node33000;
	wire [4-1:0] node33003;
	wire [4-1:0] node33004;
	wire [4-1:0] node33005;
	wire [4-1:0] node33007;
	wire [4-1:0] node33010;
	wire [4-1:0] node33011;
	wire [4-1:0] node33013;
	wire [4-1:0] node33016;
	wire [4-1:0] node33017;
	wire [4-1:0] node33021;
	wire [4-1:0] node33022;
	wire [4-1:0] node33023;
	wire [4-1:0] node33024;
	wire [4-1:0] node33027;
	wire [4-1:0] node33031;
	wire [4-1:0] node33032;
	wire [4-1:0] node33034;
	wire [4-1:0] node33037;
	wire [4-1:0] node33038;
	wire [4-1:0] node33041;
	wire [4-1:0] node33044;
	wire [4-1:0] node33045;
	wire [4-1:0] node33046;
	wire [4-1:0] node33047;
	wire [4-1:0] node33049;
	wire [4-1:0] node33052;
	wire [4-1:0] node33053;
	wire [4-1:0] node33056;
	wire [4-1:0] node33059;
	wire [4-1:0] node33060;
	wire [4-1:0] node33061;
	wire [4-1:0] node33063;
	wire [4-1:0] node33068;
	wire [4-1:0] node33069;
	wire [4-1:0] node33070;
	wire [4-1:0] node33071;
	wire [4-1:0] node33072;
	wire [4-1:0] node33076;
	wire [4-1:0] node33077;
	wire [4-1:0] node33080;
	wire [4-1:0] node33083;
	wire [4-1:0] node33084;
	wire [4-1:0] node33088;
	wire [4-1:0] node33089;
	wire [4-1:0] node33090;
	wire [4-1:0] node33093;
	wire [4-1:0] node33096;
	wire [4-1:0] node33097;
	wire [4-1:0] node33099;
	wire [4-1:0] node33102;
	wire [4-1:0] node33104;
	wire [4-1:0] node33107;
	wire [4-1:0] node33108;
	wire [4-1:0] node33109;
	wire [4-1:0] node33110;
	wire [4-1:0] node33111;
	wire [4-1:0] node33112;
	wire [4-1:0] node33114;
	wire [4-1:0] node33118;
	wire [4-1:0] node33120;
	wire [4-1:0] node33122;
	wire [4-1:0] node33125;
	wire [4-1:0] node33126;
	wire [4-1:0] node33127;
	wire [4-1:0] node33128;
	wire [4-1:0] node33132;
	wire [4-1:0] node33133;
	wire [4-1:0] node33136;
	wire [4-1:0] node33140;
	wire [4-1:0] node33141;
	wire [4-1:0] node33142;
	wire [4-1:0] node33145;
	wire [4-1:0] node33146;
	wire [4-1:0] node33150;
	wire [4-1:0] node33151;
	wire [4-1:0] node33152;
	wire [4-1:0] node33153;
	wire [4-1:0] node33156;
	wire [4-1:0] node33159;
	wire [4-1:0] node33160;
	wire [4-1:0] node33163;
	wire [4-1:0] node33166;
	wire [4-1:0] node33167;
	wire [4-1:0] node33170;
	wire [4-1:0] node33173;
	wire [4-1:0] node33174;
	wire [4-1:0] node33175;
	wire [4-1:0] node33177;
	wire [4-1:0] node33178;
	wire [4-1:0] node33181;
	wire [4-1:0] node33184;
	wire [4-1:0] node33186;
	wire [4-1:0] node33189;
	wire [4-1:0] node33190;
	wire [4-1:0] node33192;
	wire [4-1:0] node33195;
	wire [4-1:0] node33196;
	wire [4-1:0] node33199;
	wire [4-1:0] node33202;
	wire [4-1:0] node33203;
	wire [4-1:0] node33204;
	wire [4-1:0] node33205;
	wire [4-1:0] node33206;
	wire [4-1:0] node33207;
	wire [4-1:0] node33208;
	wire [4-1:0] node33212;
	wire [4-1:0] node33213;
	wire [4-1:0] node33215;
	wire [4-1:0] node33218;
	wire [4-1:0] node33220;
	wire [4-1:0] node33223;
	wire [4-1:0] node33224;
	wire [4-1:0] node33225;
	wire [4-1:0] node33228;
	wire [4-1:0] node33232;
	wire [4-1:0] node33233;
	wire [4-1:0] node33234;
	wire [4-1:0] node33235;
	wire [4-1:0] node33238;
	wire [4-1:0] node33241;
	wire [4-1:0] node33243;
	wire [4-1:0] node33246;
	wire [4-1:0] node33247;
	wire [4-1:0] node33248;
	wire [4-1:0] node33251;
	wire [4-1:0] node33254;
	wire [4-1:0] node33255;
	wire [4-1:0] node33258;
	wire [4-1:0] node33261;
	wire [4-1:0] node33262;
	wire [4-1:0] node33263;
	wire [4-1:0] node33264;
	wire [4-1:0] node33265;
	wire [4-1:0] node33268;
	wire [4-1:0] node33271;
	wire [4-1:0] node33272;
	wire [4-1:0] node33275;
	wire [4-1:0] node33278;
	wire [4-1:0] node33279;
	wire [4-1:0] node33281;
	wire [4-1:0] node33285;
	wire [4-1:0] node33286;
	wire [4-1:0] node33287;
	wire [4-1:0] node33290;
	wire [4-1:0] node33291;
	wire [4-1:0] node33294;
	wire [4-1:0] node33297;
	wire [4-1:0] node33299;
	wire [4-1:0] node33302;
	wire [4-1:0] node33303;
	wire [4-1:0] node33304;
	wire [4-1:0] node33305;
	wire [4-1:0] node33306;
	wire [4-1:0] node33307;
	wire [4-1:0] node33310;
	wire [4-1:0] node33313;
	wire [4-1:0] node33314;
	wire [4-1:0] node33318;
	wire [4-1:0] node33320;
	wire [4-1:0] node33321;
	wire [4-1:0] node33322;
	wire [4-1:0] node33325;
	wire [4-1:0] node33328;
	wire [4-1:0] node33329;
	wire [4-1:0] node33333;
	wire [4-1:0] node33334;
	wire [4-1:0] node33335;
	wire [4-1:0] node33338;
	wire [4-1:0] node33341;
	wire [4-1:0] node33342;
	wire [4-1:0] node33346;
	wire [4-1:0] node33347;
	wire [4-1:0] node33348;
	wire [4-1:0] node33349;
	wire [4-1:0] node33351;
	wire [4-1:0] node33354;
	wire [4-1:0] node33355;
	wire [4-1:0] node33358;
	wire [4-1:0] node33361;
	wire [4-1:0] node33362;
	wire [4-1:0] node33363;
	wire [4-1:0] node33366;
	wire [4-1:0] node33369;
	wire [4-1:0] node33370;
	wire [4-1:0] node33374;
	wire [4-1:0] node33375;
	wire [4-1:0] node33376;
	wire [4-1:0] node33377;
	wire [4-1:0] node33380;
	wire [4-1:0] node33383;
	wire [4-1:0] node33384;
	wire [4-1:0] node33385;
	wire [4-1:0] node33388;
	wire [4-1:0] node33392;
	wire [4-1:0] node33393;
	wire [4-1:0] node33395;
	wire [4-1:0] node33398;
	wire [4-1:0] node33400;
	wire [4-1:0] node33403;
	wire [4-1:0] node33404;
	wire [4-1:0] node33405;
	wire [4-1:0] node33406;
	wire [4-1:0] node33407;
	wire [4-1:0] node33408;
	wire [4-1:0] node33409;
	wire [4-1:0] node33410;
	wire [4-1:0] node33411;
	wire [4-1:0] node33412;
	wire [4-1:0] node33413;
	wire [4-1:0] node33417;
	wire [4-1:0] node33419;
	wire [4-1:0] node33422;
	wire [4-1:0] node33424;
	wire [4-1:0] node33425;
	wire [4-1:0] node33429;
	wire [4-1:0] node33430;
	wire [4-1:0] node33431;
	wire [4-1:0] node33432;
	wire [4-1:0] node33436;
	wire [4-1:0] node33438;
	wire [4-1:0] node33441;
	wire [4-1:0] node33443;
	wire [4-1:0] node33446;
	wire [4-1:0] node33447;
	wire [4-1:0] node33448;
	wire [4-1:0] node33449;
	wire [4-1:0] node33450;
	wire [4-1:0] node33453;
	wire [4-1:0] node33456;
	wire [4-1:0] node33457;
	wire [4-1:0] node33461;
	wire [4-1:0] node33462;
	wire [4-1:0] node33463;
	wire [4-1:0] node33467;
	wire [4-1:0] node33468;
	wire [4-1:0] node33471;
	wire [4-1:0] node33474;
	wire [4-1:0] node33475;
	wire [4-1:0] node33476;
	wire [4-1:0] node33479;
	wire [4-1:0] node33482;
	wire [4-1:0] node33483;
	wire [4-1:0] node33484;
	wire [4-1:0] node33487;
	wire [4-1:0] node33490;
	wire [4-1:0] node33491;
	wire [4-1:0] node33494;
	wire [4-1:0] node33497;
	wire [4-1:0] node33498;
	wire [4-1:0] node33499;
	wire [4-1:0] node33500;
	wire [4-1:0] node33501;
	wire [4-1:0] node33504;
	wire [4-1:0] node33507;
	wire [4-1:0] node33508;
	wire [4-1:0] node33509;
	wire [4-1:0] node33512;
	wire [4-1:0] node33515;
	wire [4-1:0] node33516;
	wire [4-1:0] node33519;
	wire [4-1:0] node33522;
	wire [4-1:0] node33523;
	wire [4-1:0] node33524;
	wire [4-1:0] node33528;
	wire [4-1:0] node33529;
	wire [4-1:0] node33530;
	wire [4-1:0] node33534;
	wire [4-1:0] node33537;
	wire [4-1:0] node33538;
	wire [4-1:0] node33539;
	wire [4-1:0] node33540;
	wire [4-1:0] node33541;
	wire [4-1:0] node33545;
	wire [4-1:0] node33548;
	wire [4-1:0] node33550;
	wire [4-1:0] node33553;
	wire [4-1:0] node33554;
	wire [4-1:0] node33555;
	wire [4-1:0] node33558;
	wire [4-1:0] node33559;
	wire [4-1:0] node33563;
	wire [4-1:0] node33564;
	wire [4-1:0] node33568;
	wire [4-1:0] node33569;
	wire [4-1:0] node33570;
	wire [4-1:0] node33571;
	wire [4-1:0] node33572;
	wire [4-1:0] node33574;
	wire [4-1:0] node33575;
	wire [4-1:0] node33578;
	wire [4-1:0] node33582;
	wire [4-1:0] node33584;
	wire [4-1:0] node33585;
	wire [4-1:0] node33587;
	wire [4-1:0] node33591;
	wire [4-1:0] node33592;
	wire [4-1:0] node33593;
	wire [4-1:0] node33595;
	wire [4-1:0] node33596;
	wire [4-1:0] node33600;
	wire [4-1:0] node33601;
	wire [4-1:0] node33603;
	wire [4-1:0] node33606;
	wire [4-1:0] node33607;
	wire [4-1:0] node33611;
	wire [4-1:0] node33612;
	wire [4-1:0] node33614;
	wire [4-1:0] node33615;
	wire [4-1:0] node33618;
	wire [4-1:0] node33621;
	wire [4-1:0] node33622;
	wire [4-1:0] node33624;
	wire [4-1:0] node33627;
	wire [4-1:0] node33630;
	wire [4-1:0] node33631;
	wire [4-1:0] node33632;
	wire [4-1:0] node33633;
	wire [4-1:0] node33634;
	wire [4-1:0] node33638;
	wire [4-1:0] node33639;
	wire [4-1:0] node33641;
	wire [4-1:0] node33644;
	wire [4-1:0] node33646;
	wire [4-1:0] node33649;
	wire [4-1:0] node33650;
	wire [4-1:0] node33653;
	wire [4-1:0] node33654;
	wire [4-1:0] node33655;
	wire [4-1:0] node33659;
	wire [4-1:0] node33660;
	wire [4-1:0] node33664;
	wire [4-1:0] node33665;
	wire [4-1:0] node33666;
	wire [4-1:0] node33667;
	wire [4-1:0] node33668;
	wire [4-1:0] node33671;
	wire [4-1:0] node33675;
	wire [4-1:0] node33676;
	wire [4-1:0] node33679;
	wire [4-1:0] node33682;
	wire [4-1:0] node33683;
	wire [4-1:0] node33684;
	wire [4-1:0] node33688;
	wire [4-1:0] node33689;
	wire [4-1:0] node33690;
	wire [4-1:0] node33694;
	wire [4-1:0] node33695;
	wire [4-1:0] node33699;
	wire [4-1:0] node33700;
	wire [4-1:0] node33701;
	wire [4-1:0] node33702;
	wire [4-1:0] node33703;
	wire [4-1:0] node33704;
	wire [4-1:0] node33708;
	wire [4-1:0] node33709;
	wire [4-1:0] node33712;
	wire [4-1:0] node33715;
	wire [4-1:0] node33716;
	wire [4-1:0] node33717;
	wire [4-1:0] node33719;
	wire [4-1:0] node33722;
	wire [4-1:0] node33724;
	wire [4-1:0] node33727;
	wire [4-1:0] node33728;
	wire [4-1:0] node33729;
	wire [4-1:0] node33732;
	wire [4-1:0] node33735;
	wire [4-1:0] node33736;
	wire [4-1:0] node33739;
	wire [4-1:0] node33741;
	wire [4-1:0] node33744;
	wire [4-1:0] node33745;
	wire [4-1:0] node33746;
	wire [4-1:0] node33747;
	wire [4-1:0] node33748;
	wire [4-1:0] node33751;
	wire [4-1:0] node33754;
	wire [4-1:0] node33755;
	wire [4-1:0] node33758;
	wire [4-1:0] node33761;
	wire [4-1:0] node33762;
	wire [4-1:0] node33763;
	wire [4-1:0] node33764;
	wire [4-1:0] node33767;
	wire [4-1:0] node33770;
	wire [4-1:0] node33771;
	wire [4-1:0] node33774;
	wire [4-1:0] node33777;
	wire [4-1:0] node33778;
	wire [4-1:0] node33781;
	wire [4-1:0] node33784;
	wire [4-1:0] node33785;
	wire [4-1:0] node33786;
	wire [4-1:0] node33787;
	wire [4-1:0] node33788;
	wire [4-1:0] node33791;
	wire [4-1:0] node33795;
	wire [4-1:0] node33797;
	wire [4-1:0] node33800;
	wire [4-1:0] node33801;
	wire [4-1:0] node33802;
	wire [4-1:0] node33806;
	wire [4-1:0] node33807;
	wire [4-1:0] node33810;
	wire [4-1:0] node33813;
	wire [4-1:0] node33814;
	wire [4-1:0] node33815;
	wire [4-1:0] node33816;
	wire [4-1:0] node33817;
	wire [4-1:0] node33818;
	wire [4-1:0] node33819;
	wire [4-1:0] node33822;
	wire [4-1:0] node33825;
	wire [4-1:0] node33826;
	wire [4-1:0] node33830;
	wire [4-1:0] node33831;
	wire [4-1:0] node33833;
	wire [4-1:0] node33836;
	wire [4-1:0] node33837;
	wire [4-1:0] node33840;
	wire [4-1:0] node33843;
	wire [4-1:0] node33844;
	wire [4-1:0] node33846;
	wire [4-1:0] node33848;
	wire [4-1:0] node33851;
	wire [4-1:0] node33852;
	wire [4-1:0] node33854;
	wire [4-1:0] node33857;
	wire [4-1:0] node33860;
	wire [4-1:0] node33861;
	wire [4-1:0] node33862;
	wire [4-1:0] node33864;
	wire [4-1:0] node33865;
	wire [4-1:0] node33869;
	wire [4-1:0] node33870;
	wire [4-1:0] node33871;
	wire [4-1:0] node33875;
	wire [4-1:0] node33878;
	wire [4-1:0] node33879;
	wire [4-1:0] node33880;
	wire [4-1:0] node33881;
	wire [4-1:0] node33885;
	wire [4-1:0] node33886;
	wire [4-1:0] node33889;
	wire [4-1:0] node33892;
	wire [4-1:0] node33893;
	wire [4-1:0] node33894;
	wire [4-1:0] node33898;
	wire [4-1:0] node33901;
	wire [4-1:0] node33902;
	wire [4-1:0] node33903;
	wire [4-1:0] node33904;
	wire [4-1:0] node33905;
	wire [4-1:0] node33906;
	wire [4-1:0] node33910;
	wire [4-1:0] node33912;
	wire [4-1:0] node33915;
	wire [4-1:0] node33918;
	wire [4-1:0] node33919;
	wire [4-1:0] node33920;
	wire [4-1:0] node33921;
	wire [4-1:0] node33925;
	wire [4-1:0] node33927;
	wire [4-1:0] node33930;
	wire [4-1:0] node33931;
	wire [4-1:0] node33932;
	wire [4-1:0] node33935;
	wire [4-1:0] node33938;
	wire [4-1:0] node33939;
	wire [4-1:0] node33942;
	wire [4-1:0] node33945;
	wire [4-1:0] node33946;
	wire [4-1:0] node33947;
	wire [4-1:0] node33948;
	wire [4-1:0] node33949;
	wire [4-1:0] node33952;
	wire [4-1:0] node33956;
	wire [4-1:0] node33957;
	wire [4-1:0] node33959;
	wire [4-1:0] node33963;
	wire [4-1:0] node33964;
	wire [4-1:0] node33965;
	wire [4-1:0] node33966;
	wire [4-1:0] node33969;
	wire [4-1:0] node33972;
	wire [4-1:0] node33975;
	wire [4-1:0] node33976;
	wire [4-1:0] node33977;
	wire [4-1:0] node33980;
	wire [4-1:0] node33983;
	wire [4-1:0] node33986;
	wire [4-1:0] node33987;
	wire [4-1:0] node33988;
	wire [4-1:0] node33989;
	wire [4-1:0] node33990;
	wire [4-1:0] node33991;
	wire [4-1:0] node33992;
	wire [4-1:0] node33993;
	wire [4-1:0] node33996;
	wire [4-1:0] node33999;
	wire [4-1:0] node34000;
	wire [4-1:0] node34001;
	wire [4-1:0] node34005;
	wire [4-1:0] node34006;
	wire [4-1:0] node34010;
	wire [4-1:0] node34011;
	wire [4-1:0] node34012;
	wire [4-1:0] node34013;
	wire [4-1:0] node34016;
	wire [4-1:0] node34020;
	wire [4-1:0] node34021;
	wire [4-1:0] node34022;
	wire [4-1:0] node34025;
	wire [4-1:0] node34029;
	wire [4-1:0] node34030;
	wire [4-1:0] node34031;
	wire [4-1:0] node34032;
	wire [4-1:0] node34035;
	wire [4-1:0] node34036;
	wire [4-1:0] node34040;
	wire [4-1:0] node34041;
	wire [4-1:0] node34043;
	wire [4-1:0] node34047;
	wire [4-1:0] node34048;
	wire [4-1:0] node34049;
	wire [4-1:0] node34053;
	wire [4-1:0] node34054;
	wire [4-1:0] node34055;
	wire [4-1:0] node34058;
	wire [4-1:0] node34061;
	wire [4-1:0] node34064;
	wire [4-1:0] node34065;
	wire [4-1:0] node34066;
	wire [4-1:0] node34067;
	wire [4-1:0] node34068;
	wire [4-1:0] node34070;
	wire [4-1:0] node34073;
	wire [4-1:0] node34074;
	wire [4-1:0] node34078;
	wire [4-1:0] node34079;
	wire [4-1:0] node34080;
	wire [4-1:0] node34085;
	wire [4-1:0] node34086;
	wire [4-1:0] node34087;
	wire [4-1:0] node34090;
	wire [4-1:0] node34093;
	wire [4-1:0] node34094;
	wire [4-1:0] node34097;
	wire [4-1:0] node34100;
	wire [4-1:0] node34101;
	wire [4-1:0] node34102;
	wire [4-1:0] node34103;
	wire [4-1:0] node34106;
	wire [4-1:0] node34108;
	wire [4-1:0] node34111;
	wire [4-1:0] node34112;
	wire [4-1:0] node34113;
	wire [4-1:0] node34116;
	wire [4-1:0] node34119;
	wire [4-1:0] node34120;
	wire [4-1:0] node34124;
	wire [4-1:0] node34125;
	wire [4-1:0] node34126;
	wire [4-1:0] node34127;
	wire [4-1:0] node34130;
	wire [4-1:0] node34133;
	wire [4-1:0] node34136;
	wire [4-1:0] node34137;
	wire [4-1:0] node34141;
	wire [4-1:0] node34142;
	wire [4-1:0] node34143;
	wire [4-1:0] node34144;
	wire [4-1:0] node34145;
	wire [4-1:0] node34146;
	wire [4-1:0] node34148;
	wire [4-1:0] node34151;
	wire [4-1:0] node34154;
	wire [4-1:0] node34155;
	wire [4-1:0] node34156;
	wire [4-1:0] node34160;
	wire [4-1:0] node34161;
	wire [4-1:0] node34165;
	wire [4-1:0] node34166;
	wire [4-1:0] node34167;
	wire [4-1:0] node34169;
	wire [4-1:0] node34172;
	wire [4-1:0] node34175;
	wire [4-1:0] node34176;
	wire [4-1:0] node34177;
	wire [4-1:0] node34181;
	wire [4-1:0] node34184;
	wire [4-1:0] node34185;
	wire [4-1:0] node34186;
	wire [4-1:0] node34187;
	wire [4-1:0] node34190;
	wire [4-1:0] node34193;
	wire [4-1:0] node34194;
	wire [4-1:0] node34195;
	wire [4-1:0] node34198;
	wire [4-1:0] node34202;
	wire [4-1:0] node34203;
	wire [4-1:0] node34204;
	wire [4-1:0] node34206;
	wire [4-1:0] node34209;
	wire [4-1:0] node34210;
	wire [4-1:0] node34213;
	wire [4-1:0] node34216;
	wire [4-1:0] node34217;
	wire [4-1:0] node34219;
	wire [4-1:0] node34223;
	wire [4-1:0] node34224;
	wire [4-1:0] node34225;
	wire [4-1:0] node34226;
	wire [4-1:0] node34227;
	wire [4-1:0] node34230;
	wire [4-1:0] node34233;
	wire [4-1:0] node34234;
	wire [4-1:0] node34237;
	wire [4-1:0] node34238;
	wire [4-1:0] node34241;
	wire [4-1:0] node34244;
	wire [4-1:0] node34245;
	wire [4-1:0] node34246;
	wire [4-1:0] node34249;
	wire [4-1:0] node34250;
	wire [4-1:0] node34253;
	wire [4-1:0] node34256;
	wire [4-1:0] node34259;
	wire [4-1:0] node34260;
	wire [4-1:0] node34261;
	wire [4-1:0] node34262;
	wire [4-1:0] node34263;
	wire [4-1:0] node34266;
	wire [4-1:0] node34269;
	wire [4-1:0] node34270;
	wire [4-1:0] node34274;
	wire [4-1:0] node34276;
	wire [4-1:0] node34277;
	wire [4-1:0] node34281;
	wire [4-1:0] node34282;
	wire [4-1:0] node34284;
	wire [4-1:0] node34285;
	wire [4-1:0] node34289;
	wire [4-1:0] node34291;
	wire [4-1:0] node34292;
	wire [4-1:0] node34296;
	wire [4-1:0] node34297;
	wire [4-1:0] node34298;
	wire [4-1:0] node34299;
	wire [4-1:0] node34300;
	wire [4-1:0] node34301;
	wire [4-1:0] node34302;
	wire [4-1:0] node34305;
	wire [4-1:0] node34308;
	wire [4-1:0] node34309;
	wire [4-1:0] node34312;
	wire [4-1:0] node34315;
	wire [4-1:0] node34316;
	wire [4-1:0] node34317;
	wire [4-1:0] node34320;
	wire [4-1:0] node34323;
	wire [4-1:0] node34324;
	wire [4-1:0] node34327;
	wire [4-1:0] node34330;
	wire [4-1:0] node34331;
	wire [4-1:0] node34332;
	wire [4-1:0] node34335;
	wire [4-1:0] node34337;
	wire [4-1:0] node34340;
	wire [4-1:0] node34341;
	wire [4-1:0] node34343;
	wire [4-1:0] node34346;
	wire [4-1:0] node34347;
	wire [4-1:0] node34350;
	wire [4-1:0] node34353;
	wire [4-1:0] node34354;
	wire [4-1:0] node34355;
	wire [4-1:0] node34357;
	wire [4-1:0] node34358;
	wire [4-1:0] node34361;
	wire [4-1:0] node34364;
	wire [4-1:0] node34365;
	wire [4-1:0] node34366;
	wire [4-1:0] node34370;
	wire [4-1:0] node34373;
	wire [4-1:0] node34374;
	wire [4-1:0] node34375;
	wire [4-1:0] node34376;
	wire [4-1:0] node34378;
	wire [4-1:0] node34382;
	wire [4-1:0] node34383;
	wire [4-1:0] node34386;
	wire [4-1:0] node34389;
	wire [4-1:0] node34390;
	wire [4-1:0] node34391;
	wire [4-1:0] node34392;
	wire [4-1:0] node34395;
	wire [4-1:0] node34399;
	wire [4-1:0] node34401;
	wire [4-1:0] node34403;
	wire [4-1:0] node34406;
	wire [4-1:0] node34407;
	wire [4-1:0] node34408;
	wire [4-1:0] node34409;
	wire [4-1:0] node34410;
	wire [4-1:0] node34411;
	wire [4-1:0] node34412;
	wire [4-1:0] node34415;
	wire [4-1:0] node34419;
	wire [4-1:0] node34420;
	wire [4-1:0] node34421;
	wire [4-1:0] node34424;
	wire [4-1:0] node34428;
	wire [4-1:0] node34429;
	wire [4-1:0] node34430;
	wire [4-1:0] node34431;
	wire [4-1:0] node34434;
	wire [4-1:0] node34437;
	wire [4-1:0] node34438;
	wire [4-1:0] node34441;
	wire [4-1:0] node34445;
	wire [4-1:0] node34446;
	wire [4-1:0] node34447;
	wire [4-1:0] node34449;
	wire [4-1:0] node34450;
	wire [4-1:0] node34454;
	wire [4-1:0] node34455;
	wire [4-1:0] node34456;
	wire [4-1:0] node34459;
	wire [4-1:0] node34463;
	wire [4-1:0] node34464;
	wire [4-1:0] node34465;
	wire [4-1:0] node34469;
	wire [4-1:0] node34470;
	wire [4-1:0] node34474;
	wire [4-1:0] node34475;
	wire [4-1:0] node34476;
	wire [4-1:0] node34477;
	wire [4-1:0] node34479;
	wire [4-1:0] node34480;
	wire [4-1:0] node34484;
	wire [4-1:0] node34486;
	wire [4-1:0] node34489;
	wire [4-1:0] node34490;
	wire [4-1:0] node34491;
	wire [4-1:0] node34492;
	wire [4-1:0] node34496;
	wire [4-1:0] node34497;
	wire [4-1:0] node34500;
	wire [4-1:0] node34503;
	wire [4-1:0] node34504;
	wire [4-1:0] node34506;
	wire [4-1:0] node34509;
	wire [4-1:0] node34511;
	wire [4-1:0] node34514;
	wire [4-1:0] node34515;
	wire [4-1:0] node34516;
	wire [4-1:0] node34517;
	wire [4-1:0] node34518;
	wire [4-1:0] node34523;
	wire [4-1:0] node34524;
	wire [4-1:0] node34525;
	wire [4-1:0] node34530;
	wire [4-1:0] node34531;
	wire [4-1:0] node34532;
	wire [4-1:0] node34534;
	wire [4-1:0] node34537;
	wire [4-1:0] node34539;
	wire [4-1:0] node34542;
	wire [4-1:0] node34543;
	wire [4-1:0] node34544;
	wire [4-1:0] node34547;
	wire [4-1:0] node34551;
	wire [4-1:0] node34552;
	wire [4-1:0] node34553;
	wire [4-1:0] node34554;
	wire [4-1:0] node34555;
	wire [4-1:0] node34556;
	wire [4-1:0] node34557;
	wire [4-1:0] node34558;
	wire [4-1:0] node34559;
	wire [4-1:0] node34562;
	wire [4-1:0] node34565;
	wire [4-1:0] node34567;
	wire [4-1:0] node34568;
	wire [4-1:0] node34572;
	wire [4-1:0] node34573;
	wire [4-1:0] node34574;
	wire [4-1:0] node34577;
	wire [4-1:0] node34580;
	wire [4-1:0] node34581;
	wire [4-1:0] node34582;
	wire [4-1:0] node34586;
	wire [4-1:0] node34587;
	wire [4-1:0] node34590;
	wire [4-1:0] node34593;
	wire [4-1:0] node34594;
	wire [4-1:0] node34595;
	wire [4-1:0] node34598;
	wire [4-1:0] node34599;
	wire [4-1:0] node34600;
	wire [4-1:0] node34603;
	wire [4-1:0] node34607;
	wire [4-1:0] node34608;
	wire [4-1:0] node34610;
	wire [4-1:0] node34613;
	wire [4-1:0] node34614;
	wire [4-1:0] node34615;
	wire [4-1:0] node34618;
	wire [4-1:0] node34622;
	wire [4-1:0] node34623;
	wire [4-1:0] node34624;
	wire [4-1:0] node34625;
	wire [4-1:0] node34627;
	wire [4-1:0] node34630;
	wire [4-1:0] node34631;
	wire [4-1:0] node34632;
	wire [4-1:0] node34635;
	wire [4-1:0] node34638;
	wire [4-1:0] node34640;
	wire [4-1:0] node34643;
	wire [4-1:0] node34644;
	wire [4-1:0] node34647;
	wire [4-1:0] node34649;
	wire [4-1:0] node34652;
	wire [4-1:0] node34653;
	wire [4-1:0] node34654;
	wire [4-1:0] node34656;
	wire [4-1:0] node34657;
	wire [4-1:0] node34660;
	wire [4-1:0] node34663;
	wire [4-1:0] node34665;
	wire [4-1:0] node34666;
	wire [4-1:0] node34669;
	wire [4-1:0] node34672;
	wire [4-1:0] node34673;
	wire [4-1:0] node34674;
	wire [4-1:0] node34678;
	wire [4-1:0] node34680;
	wire [4-1:0] node34683;
	wire [4-1:0] node34684;
	wire [4-1:0] node34685;
	wire [4-1:0] node34686;
	wire [4-1:0] node34687;
	wire [4-1:0] node34688;
	wire [4-1:0] node34691;
	wire [4-1:0] node34693;
	wire [4-1:0] node34696;
	wire [4-1:0] node34699;
	wire [4-1:0] node34700;
	wire [4-1:0] node34701;
	wire [4-1:0] node34704;
	wire [4-1:0] node34706;
	wire [4-1:0] node34709;
	wire [4-1:0] node34712;
	wire [4-1:0] node34713;
	wire [4-1:0] node34714;
	wire [4-1:0] node34715;
	wire [4-1:0] node34718;
	wire [4-1:0] node34721;
	wire [4-1:0] node34722;
	wire [4-1:0] node34725;
	wire [4-1:0] node34728;
	wire [4-1:0] node34729;
	wire [4-1:0] node34730;
	wire [4-1:0] node34731;
	wire [4-1:0] node34734;
	wire [4-1:0] node34737;
	wire [4-1:0] node34738;
	wire [4-1:0] node34742;
	wire [4-1:0] node34743;
	wire [4-1:0] node34744;
	wire [4-1:0] node34747;
	wire [4-1:0] node34750;
	wire [4-1:0] node34751;
	wire [4-1:0] node34755;
	wire [4-1:0] node34756;
	wire [4-1:0] node34757;
	wire [4-1:0] node34758;
	wire [4-1:0] node34761;
	wire [4-1:0] node34763;
	wire [4-1:0] node34764;
	wire [4-1:0] node34768;
	wire [4-1:0] node34769;
	wire [4-1:0] node34772;
	wire [4-1:0] node34773;
	wire [4-1:0] node34774;
	wire [4-1:0] node34778;
	wire [4-1:0] node34781;
	wire [4-1:0] node34782;
	wire [4-1:0] node34783;
	wire [4-1:0] node34784;
	wire [4-1:0] node34785;
	wire [4-1:0] node34790;
	wire [4-1:0] node34792;
	wire [4-1:0] node34793;
	wire [4-1:0] node34796;
	wire [4-1:0] node34799;
	wire [4-1:0] node34800;
	wire [4-1:0] node34802;
	wire [4-1:0] node34803;
	wire [4-1:0] node34807;
	wire [4-1:0] node34808;
	wire [4-1:0] node34809;
	wire [4-1:0] node34814;
	wire [4-1:0] node34815;
	wire [4-1:0] node34816;
	wire [4-1:0] node34817;
	wire [4-1:0] node34818;
	wire [4-1:0] node34819;
	wire [4-1:0] node34822;
	wire [4-1:0] node34824;
	wire [4-1:0] node34827;
	wire [4-1:0] node34828;
	wire [4-1:0] node34829;
	wire [4-1:0] node34832;
	wire [4-1:0] node34835;
	wire [4-1:0] node34836;
	wire [4-1:0] node34839;
	wire [4-1:0] node34842;
	wire [4-1:0] node34843;
	wire [4-1:0] node34844;
	wire [4-1:0] node34845;
	wire [4-1:0] node34847;
	wire [4-1:0] node34850;
	wire [4-1:0] node34851;
	wire [4-1:0] node34855;
	wire [4-1:0] node34856;
	wire [4-1:0] node34859;
	wire [4-1:0] node34862;
	wire [4-1:0] node34863;
	wire [4-1:0] node34864;
	wire [4-1:0] node34867;
	wire [4-1:0] node34871;
	wire [4-1:0] node34872;
	wire [4-1:0] node34873;
	wire [4-1:0] node34874;
	wire [4-1:0] node34875;
	wire [4-1:0] node34878;
	wire [4-1:0] node34881;
	wire [4-1:0] node34882;
	wire [4-1:0] node34885;
	wire [4-1:0] node34888;
	wire [4-1:0] node34889;
	wire [4-1:0] node34890;
	wire [4-1:0] node34894;
	wire [4-1:0] node34897;
	wire [4-1:0] node34898;
	wire [4-1:0] node34899;
	wire [4-1:0] node34900;
	wire [4-1:0] node34904;
	wire [4-1:0] node34905;
	wire [4-1:0] node34908;
	wire [4-1:0] node34911;
	wire [4-1:0] node34912;
	wire [4-1:0] node34913;
	wire [4-1:0] node34917;
	wire [4-1:0] node34920;
	wire [4-1:0] node34921;
	wire [4-1:0] node34922;
	wire [4-1:0] node34923;
	wire [4-1:0] node34924;
	wire [4-1:0] node34925;
	wire [4-1:0] node34926;
	wire [4-1:0] node34930;
	wire [4-1:0] node34931;
	wire [4-1:0] node34935;
	wire [4-1:0] node34937;
	wire [4-1:0] node34938;
	wire [4-1:0] node34941;
	wire [4-1:0] node34944;
	wire [4-1:0] node34945;
	wire [4-1:0] node34946;
	wire [4-1:0] node34949;
	wire [4-1:0] node34952;
	wire [4-1:0] node34953;
	wire [4-1:0] node34956;
	wire [4-1:0] node34959;
	wire [4-1:0] node34960;
	wire [4-1:0] node34961;
	wire [4-1:0] node34962;
	wire [4-1:0] node34965;
	wire [4-1:0] node34968;
	wire [4-1:0] node34970;
	wire [4-1:0] node34973;
	wire [4-1:0] node34974;
	wire [4-1:0] node34975;
	wire [4-1:0] node34978;
	wire [4-1:0] node34981;
	wire [4-1:0] node34982;
	wire [4-1:0] node34985;
	wire [4-1:0] node34988;
	wire [4-1:0] node34989;
	wire [4-1:0] node34990;
	wire [4-1:0] node34991;
	wire [4-1:0] node34992;
	wire [4-1:0] node34995;
	wire [4-1:0] node34998;
	wire [4-1:0] node34999;
	wire [4-1:0] node35002;
	wire [4-1:0] node35005;
	wire [4-1:0] node35006;
	wire [4-1:0] node35007;
	wire [4-1:0] node35010;
	wire [4-1:0] node35013;
	wire [4-1:0] node35014;
	wire [4-1:0] node35017;
	wire [4-1:0] node35020;
	wire [4-1:0] node35021;
	wire [4-1:0] node35022;
	wire [4-1:0] node35023;
	wire [4-1:0] node35027;
	wire [4-1:0] node35028;
	wire [4-1:0] node35032;
	wire [4-1:0] node35033;
	wire [4-1:0] node35034;
	wire [4-1:0] node35038;
	wire [4-1:0] node35039;
	wire [4-1:0] node35040;
	wire [4-1:0] node35043;
	wire [4-1:0] node35046;
	wire [4-1:0] node35048;
	wire [4-1:0] node35051;
	wire [4-1:0] node35052;
	wire [4-1:0] node35053;
	wire [4-1:0] node35054;
	wire [4-1:0] node35055;
	wire [4-1:0] node35056;
	wire [4-1:0] node35057;
	wire [4-1:0] node35059;
	wire [4-1:0] node35061;
	wire [4-1:0] node35064;
	wire [4-1:0] node35065;
	wire [4-1:0] node35066;
	wire [4-1:0] node35070;
	wire [4-1:0] node35071;
	wire [4-1:0] node35074;
	wire [4-1:0] node35077;
	wire [4-1:0] node35078;
	wire [4-1:0] node35079;
	wire [4-1:0] node35080;
	wire [4-1:0] node35084;
	wire [4-1:0] node35087;
	wire [4-1:0] node35088;
	wire [4-1:0] node35092;
	wire [4-1:0] node35093;
	wire [4-1:0] node35094;
	wire [4-1:0] node35097;
	wire [4-1:0] node35098;
	wire [4-1:0] node35100;
	wire [4-1:0] node35103;
	wire [4-1:0] node35106;
	wire [4-1:0] node35107;
	wire [4-1:0] node35108;
	wire [4-1:0] node35111;
	wire [4-1:0] node35114;
	wire [4-1:0] node35115;
	wire [4-1:0] node35116;
	wire [4-1:0] node35119;
	wire [4-1:0] node35123;
	wire [4-1:0] node35124;
	wire [4-1:0] node35125;
	wire [4-1:0] node35127;
	wire [4-1:0] node35128;
	wire [4-1:0] node35129;
	wire [4-1:0] node35132;
	wire [4-1:0] node35135;
	wire [4-1:0] node35136;
	wire [4-1:0] node35140;
	wire [4-1:0] node35141;
	wire [4-1:0] node35144;
	wire [4-1:0] node35146;
	wire [4-1:0] node35147;
	wire [4-1:0] node35151;
	wire [4-1:0] node35152;
	wire [4-1:0] node35153;
	wire [4-1:0] node35155;
	wire [4-1:0] node35156;
	wire [4-1:0] node35159;
	wire [4-1:0] node35162;
	wire [4-1:0] node35163;
	wire [4-1:0] node35164;
	wire [4-1:0] node35169;
	wire [4-1:0] node35170;
	wire [4-1:0] node35172;
	wire [4-1:0] node35175;
	wire [4-1:0] node35176;
	wire [4-1:0] node35179;
	wire [4-1:0] node35182;
	wire [4-1:0] node35183;
	wire [4-1:0] node35184;
	wire [4-1:0] node35185;
	wire [4-1:0] node35186;
	wire [4-1:0] node35187;
	wire [4-1:0] node35190;
	wire [4-1:0] node35192;
	wire [4-1:0] node35195;
	wire [4-1:0] node35196;
	wire [4-1:0] node35200;
	wire [4-1:0] node35201;
	wire [4-1:0] node35202;
	wire [4-1:0] node35205;
	wire [4-1:0] node35208;
	wire [4-1:0] node35209;
	wire [4-1:0] node35210;
	wire [4-1:0] node35215;
	wire [4-1:0] node35216;
	wire [4-1:0] node35217;
	wire [4-1:0] node35218;
	wire [4-1:0] node35219;
	wire [4-1:0] node35223;
	wire [4-1:0] node35225;
	wire [4-1:0] node35228;
	wire [4-1:0] node35229;
	wire [4-1:0] node35230;
	wire [4-1:0] node35234;
	wire [4-1:0] node35235;
	wire [4-1:0] node35239;
	wire [4-1:0] node35241;
	wire [4-1:0] node35242;
	wire [4-1:0] node35246;
	wire [4-1:0] node35247;
	wire [4-1:0] node35248;
	wire [4-1:0] node35249;
	wire [4-1:0] node35250;
	wire [4-1:0] node35251;
	wire [4-1:0] node35256;
	wire [4-1:0] node35257;
	wire [4-1:0] node35260;
	wire [4-1:0] node35262;
	wire [4-1:0] node35265;
	wire [4-1:0] node35266;
	wire [4-1:0] node35267;
	wire [4-1:0] node35270;
	wire [4-1:0] node35271;
	wire [4-1:0] node35274;
	wire [4-1:0] node35277;
	wire [4-1:0] node35278;
	wire [4-1:0] node35281;
	wire [4-1:0] node35284;
	wire [4-1:0] node35285;
	wire [4-1:0] node35286;
	wire [4-1:0] node35287;
	wire [4-1:0] node35290;
	wire [4-1:0] node35293;
	wire [4-1:0] node35294;
	wire [4-1:0] node35297;
	wire [4-1:0] node35300;
	wire [4-1:0] node35301;
	wire [4-1:0] node35302;
	wire [4-1:0] node35304;
	wire [4-1:0] node35307;
	wire [4-1:0] node35310;
	wire [4-1:0] node35311;
	wire [4-1:0] node35314;
	wire [4-1:0] node35317;
	wire [4-1:0] node35318;
	wire [4-1:0] node35319;
	wire [4-1:0] node35320;
	wire [4-1:0] node35321;
	wire [4-1:0] node35322;
	wire [4-1:0] node35323;
	wire [4-1:0] node35324;
	wire [4-1:0] node35327;
	wire [4-1:0] node35330;
	wire [4-1:0] node35331;
	wire [4-1:0] node35334;
	wire [4-1:0] node35337;
	wire [4-1:0] node35338;
	wire [4-1:0] node35340;
	wire [4-1:0] node35343;
	wire [4-1:0] node35345;
	wire [4-1:0] node35348;
	wire [4-1:0] node35349;
	wire [4-1:0] node35351;
	wire [4-1:0] node35352;
	wire [4-1:0] node35355;
	wire [4-1:0] node35358;
	wire [4-1:0] node35359;
	wire [4-1:0] node35361;
	wire [4-1:0] node35365;
	wire [4-1:0] node35366;
	wire [4-1:0] node35367;
	wire [4-1:0] node35368;
	wire [4-1:0] node35369;
	wire [4-1:0] node35373;
	wire [4-1:0] node35376;
	wire [4-1:0] node35378;
	wire [4-1:0] node35379;
	wire [4-1:0] node35382;
	wire [4-1:0] node35385;
	wire [4-1:0] node35386;
	wire [4-1:0] node35387;
	wire [4-1:0] node35388;
	wire [4-1:0] node35391;
	wire [4-1:0] node35394;
	wire [4-1:0] node35397;
	wire [4-1:0] node35398;
	wire [4-1:0] node35399;
	wire [4-1:0] node35402;
	wire [4-1:0] node35405;
	wire [4-1:0] node35408;
	wire [4-1:0] node35409;
	wire [4-1:0] node35410;
	wire [4-1:0] node35411;
	wire [4-1:0] node35414;
	wire [4-1:0] node35416;
	wire [4-1:0] node35419;
	wire [4-1:0] node35420;
	wire [4-1:0] node35421;
	wire [4-1:0] node35424;
	wire [4-1:0] node35427;
	wire [4-1:0] node35429;
	wire [4-1:0] node35432;
	wire [4-1:0] node35433;
	wire [4-1:0] node35434;
	wire [4-1:0] node35436;
	wire [4-1:0] node35438;
	wire [4-1:0] node35441;
	wire [4-1:0] node35442;
	wire [4-1:0] node35444;
	wire [4-1:0] node35447;
	wire [4-1:0] node35448;
	wire [4-1:0] node35451;
	wire [4-1:0] node35454;
	wire [4-1:0] node35455;
	wire [4-1:0] node35456;
	wire [4-1:0] node35457;
	wire [4-1:0] node35462;
	wire [4-1:0] node35463;
	wire [4-1:0] node35464;
	wire [4-1:0] node35467;
	wire [4-1:0] node35471;
	wire [4-1:0] node35472;
	wire [4-1:0] node35473;
	wire [4-1:0] node35474;
	wire [4-1:0] node35475;
	wire [4-1:0] node35476;
	wire [4-1:0] node35477;
	wire [4-1:0] node35481;
	wire [4-1:0] node35482;
	wire [4-1:0] node35485;
	wire [4-1:0] node35488;
	wire [4-1:0] node35489;
	wire [4-1:0] node35491;
	wire [4-1:0] node35494;
	wire [4-1:0] node35495;
	wire [4-1:0] node35498;
	wire [4-1:0] node35501;
	wire [4-1:0] node35502;
	wire [4-1:0] node35503;
	wire [4-1:0] node35504;
	wire [4-1:0] node35507;
	wire [4-1:0] node35511;
	wire [4-1:0] node35512;
	wire [4-1:0] node35513;
	wire [4-1:0] node35517;
	wire [4-1:0] node35518;
	wire [4-1:0] node35521;
	wire [4-1:0] node35524;
	wire [4-1:0] node35525;
	wire [4-1:0] node35526;
	wire [4-1:0] node35527;
	wire [4-1:0] node35528;
	wire [4-1:0] node35531;
	wire [4-1:0] node35534;
	wire [4-1:0] node35535;
	wire [4-1:0] node35539;
	wire [4-1:0] node35541;
	wire [4-1:0] node35543;
	wire [4-1:0] node35546;
	wire [4-1:0] node35547;
	wire [4-1:0] node35548;
	wire [4-1:0] node35551;
	wire [4-1:0] node35552;
	wire [4-1:0] node35555;
	wire [4-1:0] node35558;
	wire [4-1:0] node35559;
	wire [4-1:0] node35563;
	wire [4-1:0] node35564;
	wire [4-1:0] node35565;
	wire [4-1:0] node35566;
	wire [4-1:0] node35568;
	wire [4-1:0] node35569;
	wire [4-1:0] node35573;
	wire [4-1:0] node35574;
	wire [4-1:0] node35575;
	wire [4-1:0] node35578;
	wire [4-1:0] node35582;
	wire [4-1:0] node35583;
	wire [4-1:0] node35584;
	wire [4-1:0] node35586;
	wire [4-1:0] node35589;
	wire [4-1:0] node35590;
	wire [4-1:0] node35593;
	wire [4-1:0] node35596;
	wire [4-1:0] node35597;
	wire [4-1:0] node35600;
	wire [4-1:0] node35601;
	wire [4-1:0] node35604;
	wire [4-1:0] node35607;
	wire [4-1:0] node35608;
	wire [4-1:0] node35609;
	wire [4-1:0] node35612;
	wire [4-1:0] node35613;
	wire [4-1:0] node35614;
	wire [4-1:0] node35617;
	wire [4-1:0] node35621;
	wire [4-1:0] node35622;
	wire [4-1:0] node35623;
	wire [4-1:0] node35624;
	wire [4-1:0] node35628;
	wire [4-1:0] node35629;
	wire [4-1:0] node35633;
	wire [4-1:0] node35634;
	wire [4-1:0] node35637;
	wire [4-1:0] node35638;
	wire [4-1:0] node35641;
	wire [4-1:0] node35644;
	wire [4-1:0] node35645;
	wire [4-1:0] node35646;
	wire [4-1:0] node35647;
	wire [4-1:0] node35648;
	wire [4-1:0] node35649;
	wire [4-1:0] node35650;
	wire [4-1:0] node35651;
	wire [4-1:0] node35652;
	wire [4-1:0] node35653;
	wire [4-1:0] node35655;
	wire [4-1:0] node35658;
	wire [4-1:0] node35660;
	wire [4-1:0] node35663;
	wire [4-1:0] node35664;
	wire [4-1:0] node35665;
	wire [4-1:0] node35666;
	wire [4-1:0] node35670;
	wire [4-1:0] node35671;
	wire [4-1:0] node35674;
	wire [4-1:0] node35677;
	wire [4-1:0] node35679;
	wire [4-1:0] node35680;
	wire [4-1:0] node35684;
	wire [4-1:0] node35685;
	wire [4-1:0] node35686;
	wire [4-1:0] node35687;
	wire [4-1:0] node35689;
	wire [4-1:0] node35693;
	wire [4-1:0] node35695;
	wire [4-1:0] node35697;
	wire [4-1:0] node35700;
	wire [4-1:0] node35701;
	wire [4-1:0] node35703;
	wire [4-1:0] node35704;
	wire [4-1:0] node35707;
	wire [4-1:0] node35710;
	wire [4-1:0] node35711;
	wire [4-1:0] node35714;
	wire [4-1:0] node35717;
	wire [4-1:0] node35718;
	wire [4-1:0] node35719;
	wire [4-1:0] node35720;
	wire [4-1:0] node35721;
	wire [4-1:0] node35722;
	wire [4-1:0] node35726;
	wire [4-1:0] node35727;
	wire [4-1:0] node35731;
	wire [4-1:0] node35732;
	wire [4-1:0] node35733;
	wire [4-1:0] node35736;
	wire [4-1:0] node35739;
	wire [4-1:0] node35742;
	wire [4-1:0] node35743;
	wire [4-1:0] node35744;
	wire [4-1:0] node35745;
	wire [4-1:0] node35749;
	wire [4-1:0] node35752;
	wire [4-1:0] node35753;
	wire [4-1:0] node35756;
	wire [4-1:0] node35757;
	wire [4-1:0] node35760;
	wire [4-1:0] node35763;
	wire [4-1:0] node35764;
	wire [4-1:0] node35765;
	wire [4-1:0] node35766;
	wire [4-1:0] node35768;
	wire [4-1:0] node35772;
	wire [4-1:0] node35773;
	wire [4-1:0] node35776;
	wire [4-1:0] node35779;
	wire [4-1:0] node35780;
	wire [4-1:0] node35781;
	wire [4-1:0] node35784;
	wire [4-1:0] node35787;
	wire [4-1:0] node35788;
	wire [4-1:0] node35791;
	wire [4-1:0] node35794;
	wire [4-1:0] node35795;
	wire [4-1:0] node35796;
	wire [4-1:0] node35797;
	wire [4-1:0] node35798;
	wire [4-1:0] node35801;
	wire [4-1:0] node35802;
	wire [4-1:0] node35806;
	wire [4-1:0] node35807;
	wire [4-1:0] node35808;
	wire [4-1:0] node35811;
	wire [4-1:0] node35813;
	wire [4-1:0] node35816;
	wire [4-1:0] node35817;
	wire [4-1:0] node35818;
	wire [4-1:0] node35821;
	wire [4-1:0] node35824;
	wire [4-1:0] node35825;
	wire [4-1:0] node35829;
	wire [4-1:0] node35830;
	wire [4-1:0] node35831;
	wire [4-1:0] node35832;
	wire [4-1:0] node35833;
	wire [4-1:0] node35836;
	wire [4-1:0] node35840;
	wire [4-1:0] node35843;
	wire [4-1:0] node35844;
	wire [4-1:0] node35845;
	wire [4-1:0] node35847;
	wire [4-1:0] node35850;
	wire [4-1:0] node35851;
	wire [4-1:0] node35854;
	wire [4-1:0] node35857;
	wire [4-1:0] node35858;
	wire [4-1:0] node35859;
	wire [4-1:0] node35863;
	wire [4-1:0] node35866;
	wire [4-1:0] node35867;
	wire [4-1:0] node35868;
	wire [4-1:0] node35869;
	wire [4-1:0] node35870;
	wire [4-1:0] node35873;
	wire [4-1:0] node35874;
	wire [4-1:0] node35877;
	wire [4-1:0] node35880;
	wire [4-1:0] node35882;
	wire [4-1:0] node35885;
	wire [4-1:0] node35886;
	wire [4-1:0] node35887;
	wire [4-1:0] node35888;
	wire [4-1:0] node35892;
	wire [4-1:0] node35895;
	wire [4-1:0] node35896;
	wire [4-1:0] node35897;
	wire [4-1:0] node35900;
	wire [4-1:0] node35904;
	wire [4-1:0] node35905;
	wire [4-1:0] node35906;
	wire [4-1:0] node35907;
	wire [4-1:0] node35909;
	wire [4-1:0] node35912;
	wire [4-1:0] node35914;
	wire [4-1:0] node35917;
	wire [4-1:0] node35919;
	wire [4-1:0] node35922;
	wire [4-1:0] node35923;
	wire [4-1:0] node35924;
	wire [4-1:0] node35925;
	wire [4-1:0] node35928;
	wire [4-1:0] node35931;
	wire [4-1:0] node35933;
	wire [4-1:0] node35937;
	wire [4-1:0] node35938;
	wire [4-1:0] node35939;
	wire [4-1:0] node35940;
	wire [4-1:0] node35941;
	wire [4-1:0] node35942;
	wire [4-1:0] node35944;
	wire [4-1:0] node35945;
	wire [4-1:0] node35948;
	wire [4-1:0] node35951;
	wire [4-1:0] node35952;
	wire [4-1:0] node35953;
	wire [4-1:0] node35956;
	wire [4-1:0] node35959;
	wire [4-1:0] node35960;
	wire [4-1:0] node35963;
	wire [4-1:0] node35966;
	wire [4-1:0] node35967;
	wire [4-1:0] node35968;
	wire [4-1:0] node35971;
	wire [4-1:0] node35974;
	wire [4-1:0] node35975;
	wire [4-1:0] node35976;
	wire [4-1:0] node35979;
	wire [4-1:0] node35982;
	wire [4-1:0] node35984;
	wire [4-1:0] node35987;
	wire [4-1:0] node35988;
	wire [4-1:0] node35989;
	wire [4-1:0] node35990;
	wire [4-1:0] node35991;
	wire [4-1:0] node35994;
	wire [4-1:0] node35997;
	wire [4-1:0] node35999;
	wire [4-1:0] node36002;
	wire [4-1:0] node36004;
	wire [4-1:0] node36005;
	wire [4-1:0] node36009;
	wire [4-1:0] node36010;
	wire [4-1:0] node36011;
	wire [4-1:0] node36013;
	wire [4-1:0] node36017;
	wire [4-1:0] node36018;
	wire [4-1:0] node36021;
	wire [4-1:0] node36024;
	wire [4-1:0] node36025;
	wire [4-1:0] node36026;
	wire [4-1:0] node36027;
	wire [4-1:0] node36028;
	wire [4-1:0] node36029;
	wire [4-1:0] node36032;
	wire [4-1:0] node36035;
	wire [4-1:0] node36037;
	wire [4-1:0] node36040;
	wire [4-1:0] node36042;
	wire [4-1:0] node36045;
	wire [4-1:0] node36046;
	wire [4-1:0] node36048;
	wire [4-1:0] node36050;
	wire [4-1:0] node36053;
	wire [4-1:0] node36055;
	wire [4-1:0] node36058;
	wire [4-1:0] node36059;
	wire [4-1:0] node36060;
	wire [4-1:0] node36061;
	wire [4-1:0] node36064;
	wire [4-1:0] node36066;
	wire [4-1:0] node36069;
	wire [4-1:0] node36070;
	wire [4-1:0] node36072;
	wire [4-1:0] node36075;
	wire [4-1:0] node36076;
	wire [4-1:0] node36080;
	wire [4-1:0] node36081;
	wire [4-1:0] node36082;
	wire [4-1:0] node36085;
	wire [4-1:0] node36087;
	wire [4-1:0] node36090;
	wire [4-1:0] node36092;
	wire [4-1:0] node36095;
	wire [4-1:0] node36096;
	wire [4-1:0] node36097;
	wire [4-1:0] node36098;
	wire [4-1:0] node36099;
	wire [4-1:0] node36100;
	wire [4-1:0] node36101;
	wire [4-1:0] node36105;
	wire [4-1:0] node36106;
	wire [4-1:0] node36109;
	wire [4-1:0] node36112;
	wire [4-1:0] node36113;
	wire [4-1:0] node36117;
	wire [4-1:0] node36118;
	wire [4-1:0] node36119;
	wire [4-1:0] node36122;
	wire [4-1:0] node36124;
	wire [4-1:0] node36127;
	wire [4-1:0] node36128;
	wire [4-1:0] node36131;
	wire [4-1:0] node36133;
	wire [4-1:0] node36136;
	wire [4-1:0] node36137;
	wire [4-1:0] node36138;
	wire [4-1:0] node36140;
	wire [4-1:0] node36144;
	wire [4-1:0] node36145;
	wire [4-1:0] node36148;
	wire [4-1:0] node36149;
	wire [4-1:0] node36150;
	wire [4-1:0] node36154;
	wire [4-1:0] node36155;
	wire [4-1:0] node36159;
	wire [4-1:0] node36160;
	wire [4-1:0] node36161;
	wire [4-1:0] node36162;
	wire [4-1:0] node36164;
	wire [4-1:0] node36165;
	wire [4-1:0] node36168;
	wire [4-1:0] node36171;
	wire [4-1:0] node36174;
	wire [4-1:0] node36175;
	wire [4-1:0] node36176;
	wire [4-1:0] node36178;
	wire [4-1:0] node36181;
	wire [4-1:0] node36182;
	wire [4-1:0] node36185;
	wire [4-1:0] node36188;
	wire [4-1:0] node36189;
	wire [4-1:0] node36190;
	wire [4-1:0] node36194;
	wire [4-1:0] node36197;
	wire [4-1:0] node36198;
	wire [4-1:0] node36199;
	wire [4-1:0] node36201;
	wire [4-1:0] node36204;
	wire [4-1:0] node36206;
	wire [4-1:0] node36207;
	wire [4-1:0] node36210;
	wire [4-1:0] node36213;
	wire [4-1:0] node36214;
	wire [4-1:0] node36215;
	wire [4-1:0] node36217;
	wire [4-1:0] node36220;
	wire [4-1:0] node36223;
	wire [4-1:0] node36224;
	wire [4-1:0] node36227;
	wire [4-1:0] node36230;
	wire [4-1:0] node36231;
	wire [4-1:0] node36232;
	wire [4-1:0] node36233;
	wire [4-1:0] node36234;
	wire [4-1:0] node36235;
	wire [4-1:0] node36236;
	wire [4-1:0] node36238;
	wire [4-1:0] node36239;
	wire [4-1:0] node36242;
	wire [4-1:0] node36245;
	wire [4-1:0] node36247;
	wire [4-1:0] node36250;
	wire [4-1:0] node36251;
	wire [4-1:0] node36252;
	wire [4-1:0] node36253;
	wire [4-1:0] node36257;
	wire [4-1:0] node36259;
	wire [4-1:0] node36262;
	wire [4-1:0] node36263;
	wire [4-1:0] node36264;
	wire [4-1:0] node36268;
	wire [4-1:0] node36271;
	wire [4-1:0] node36272;
	wire [4-1:0] node36273;
	wire [4-1:0] node36274;
	wire [4-1:0] node36275;
	wire [4-1:0] node36278;
	wire [4-1:0] node36282;
	wire [4-1:0] node36284;
	wire [4-1:0] node36287;
	wire [4-1:0] node36288;
	wire [4-1:0] node36289;
	wire [4-1:0] node36291;
	wire [4-1:0] node36294;
	wire [4-1:0] node36295;
	wire [4-1:0] node36298;
	wire [4-1:0] node36301;
	wire [4-1:0] node36302;
	wire [4-1:0] node36306;
	wire [4-1:0] node36307;
	wire [4-1:0] node36308;
	wire [4-1:0] node36309;
	wire [4-1:0] node36310;
	wire [4-1:0] node36311;
	wire [4-1:0] node36314;
	wire [4-1:0] node36318;
	wire [4-1:0] node36319;
	wire [4-1:0] node36320;
	wire [4-1:0] node36325;
	wire [4-1:0] node36326;
	wire [4-1:0] node36327;
	wire [4-1:0] node36328;
	wire [4-1:0] node36333;
	wire [4-1:0] node36334;
	wire [4-1:0] node36335;
	wire [4-1:0] node36340;
	wire [4-1:0] node36341;
	wire [4-1:0] node36342;
	wire [4-1:0] node36345;
	wire [4-1:0] node36346;
	wire [4-1:0] node36347;
	wire [4-1:0] node36350;
	wire [4-1:0] node36354;
	wire [4-1:0] node36355;
	wire [4-1:0] node36356;
	wire [4-1:0] node36357;
	wire [4-1:0] node36360;
	wire [4-1:0] node36363;
	wire [4-1:0] node36365;
	wire [4-1:0] node36368;
	wire [4-1:0] node36369;
	wire [4-1:0] node36370;
	wire [4-1:0] node36373;
	wire [4-1:0] node36376;
	wire [4-1:0] node36377;
	wire [4-1:0] node36380;
	wire [4-1:0] node36383;
	wire [4-1:0] node36384;
	wire [4-1:0] node36385;
	wire [4-1:0] node36386;
	wire [4-1:0] node36387;
	wire [4-1:0] node36388;
	wire [4-1:0] node36391;
	wire [4-1:0] node36392;
	wire [4-1:0] node36396;
	wire [4-1:0] node36397;
	wire [4-1:0] node36400;
	wire [4-1:0] node36403;
	wire [4-1:0] node36404;
	wire [4-1:0] node36405;
	wire [4-1:0] node36408;
	wire [4-1:0] node36411;
	wire [4-1:0] node36412;
	wire [4-1:0] node36415;
	wire [4-1:0] node36418;
	wire [4-1:0] node36419;
	wire [4-1:0] node36421;
	wire [4-1:0] node36423;
	wire [4-1:0] node36424;
	wire [4-1:0] node36427;
	wire [4-1:0] node36430;
	wire [4-1:0] node36431;
	wire [4-1:0] node36432;
	wire [4-1:0] node36433;
	wire [4-1:0] node36437;
	wire [4-1:0] node36438;
	wire [4-1:0] node36441;
	wire [4-1:0] node36444;
	wire [4-1:0] node36445;
	wire [4-1:0] node36447;
	wire [4-1:0] node36451;
	wire [4-1:0] node36452;
	wire [4-1:0] node36453;
	wire [4-1:0] node36454;
	wire [4-1:0] node36455;
	wire [4-1:0] node36458;
	wire [4-1:0] node36459;
	wire [4-1:0] node36462;
	wire [4-1:0] node36465;
	wire [4-1:0] node36466;
	wire [4-1:0] node36467;
	wire [4-1:0] node36471;
	wire [4-1:0] node36474;
	wire [4-1:0] node36475;
	wire [4-1:0] node36476;
	wire [4-1:0] node36479;
	wire [4-1:0] node36481;
	wire [4-1:0] node36484;
	wire [4-1:0] node36485;
	wire [4-1:0] node36486;
	wire [4-1:0] node36489;
	wire [4-1:0] node36493;
	wire [4-1:0] node36494;
	wire [4-1:0] node36495;
	wire [4-1:0] node36496;
	wire [4-1:0] node36497;
	wire [4-1:0] node36500;
	wire [4-1:0] node36503;
	wire [4-1:0] node36505;
	wire [4-1:0] node36508;
	wire [4-1:0] node36509;
	wire [4-1:0] node36512;
	wire [4-1:0] node36515;
	wire [4-1:0] node36516;
	wire [4-1:0] node36517;
	wire [4-1:0] node36518;
	wire [4-1:0] node36521;
	wire [4-1:0] node36525;
	wire [4-1:0] node36527;
	wire [4-1:0] node36528;
	wire [4-1:0] node36532;
	wire [4-1:0] node36533;
	wire [4-1:0] node36534;
	wire [4-1:0] node36535;
	wire [4-1:0] node36536;
	wire [4-1:0] node36537;
	wire [4-1:0] node36538;
	wire [4-1:0] node36542;
	wire [4-1:0] node36543;
	wire [4-1:0] node36546;
	wire [4-1:0] node36549;
	wire [4-1:0] node36550;
	wire [4-1:0] node36553;
	wire [4-1:0] node36556;
	wire [4-1:0] node36557;
	wire [4-1:0] node36559;
	wire [4-1:0] node36562;
	wire [4-1:0] node36563;
	wire [4-1:0] node36564;
	wire [4-1:0] node36566;
	wire [4-1:0] node36569;
	wire [4-1:0] node36570;
	wire [4-1:0] node36573;
	wire [4-1:0] node36576;
	wire [4-1:0] node36577;
	wire [4-1:0] node36578;
	wire [4-1:0] node36582;
	wire [4-1:0] node36585;
	wire [4-1:0] node36586;
	wire [4-1:0] node36587;
	wire [4-1:0] node36588;
	wire [4-1:0] node36589;
	wire [4-1:0] node36590;
	wire [4-1:0] node36593;
	wire [4-1:0] node36596;
	wire [4-1:0] node36597;
	wire [4-1:0] node36600;
	wire [4-1:0] node36603;
	wire [4-1:0] node36604;
	wire [4-1:0] node36605;
	wire [4-1:0] node36608;
	wire [4-1:0] node36611;
	wire [4-1:0] node36612;
	wire [4-1:0] node36615;
	wire [4-1:0] node36618;
	wire [4-1:0] node36619;
	wire [4-1:0] node36620;
	wire [4-1:0] node36621;
	wire [4-1:0] node36625;
	wire [4-1:0] node36626;
	wire [4-1:0] node36629;
	wire [4-1:0] node36632;
	wire [4-1:0] node36633;
	wire [4-1:0] node36634;
	wire [4-1:0] node36638;
	wire [4-1:0] node36640;
	wire [4-1:0] node36643;
	wire [4-1:0] node36644;
	wire [4-1:0] node36645;
	wire [4-1:0] node36646;
	wire [4-1:0] node36649;
	wire [4-1:0] node36652;
	wire [4-1:0] node36654;
	wire [4-1:0] node36655;
	wire [4-1:0] node36659;
	wire [4-1:0] node36660;
	wire [4-1:0] node36661;
	wire [4-1:0] node36662;
	wire [4-1:0] node36667;
	wire [4-1:0] node36668;
	wire [4-1:0] node36669;
	wire [4-1:0] node36672;
	wire [4-1:0] node36675;
	wire [4-1:0] node36676;
	wire [4-1:0] node36680;
	wire [4-1:0] node36681;
	wire [4-1:0] node36682;
	wire [4-1:0] node36683;
	wire [4-1:0] node36684;
	wire [4-1:0] node36686;
	wire [4-1:0] node36687;
	wire [4-1:0] node36690;
	wire [4-1:0] node36693;
	wire [4-1:0] node36694;
	wire [4-1:0] node36697;
	wire [4-1:0] node36700;
	wire [4-1:0] node36701;
	wire [4-1:0] node36702;
	wire [4-1:0] node36705;
	wire [4-1:0] node36708;
	wire [4-1:0] node36709;
	wire [4-1:0] node36710;
	wire [4-1:0] node36713;
	wire [4-1:0] node36717;
	wire [4-1:0] node36718;
	wire [4-1:0] node36719;
	wire [4-1:0] node36721;
	wire [4-1:0] node36724;
	wire [4-1:0] node36725;
	wire [4-1:0] node36728;
	wire [4-1:0] node36731;
	wire [4-1:0] node36732;
	wire [4-1:0] node36733;
	wire [4-1:0] node36736;
	wire [4-1:0] node36739;
	wire [4-1:0] node36740;
	wire [4-1:0] node36741;
	wire [4-1:0] node36744;
	wire [4-1:0] node36748;
	wire [4-1:0] node36749;
	wire [4-1:0] node36750;
	wire [4-1:0] node36751;
	wire [4-1:0] node36753;
	wire [4-1:0] node36754;
	wire [4-1:0] node36757;
	wire [4-1:0] node36760;
	wire [4-1:0] node36763;
	wire [4-1:0] node36764;
	wire [4-1:0] node36765;
	wire [4-1:0] node36768;
	wire [4-1:0] node36771;
	wire [4-1:0] node36774;
	wire [4-1:0] node36775;
	wire [4-1:0] node36776;
	wire [4-1:0] node36777;
	wire [4-1:0] node36778;
	wire [4-1:0] node36781;
	wire [4-1:0] node36785;
	wire [4-1:0] node36786;
	wire [4-1:0] node36789;
	wire [4-1:0] node36792;
	wire [4-1:0] node36793;
	wire [4-1:0] node36794;
	wire [4-1:0] node36797;
	wire [4-1:0] node36801;
	wire [4-1:0] node36802;
	wire [4-1:0] node36803;
	wire [4-1:0] node36804;
	wire [4-1:0] node36805;
	wire [4-1:0] node36806;
	wire [4-1:0] node36807;
	wire [4-1:0] node36808;
	wire [4-1:0] node36809;
	wire [4-1:0] node36812;
	wire [4-1:0] node36814;
	wire [4-1:0] node36817;
	wire [4-1:0] node36818;
	wire [4-1:0] node36822;
	wire [4-1:0] node36823;
	wire [4-1:0] node36824;
	wire [4-1:0] node36827;
	wire [4-1:0] node36829;
	wire [4-1:0] node36832;
	wire [4-1:0] node36833;
	wire [4-1:0] node36834;
	wire [4-1:0] node36837;
	wire [4-1:0] node36840;
	wire [4-1:0] node36841;
	wire [4-1:0] node36845;
	wire [4-1:0] node36846;
	wire [4-1:0] node36847;
	wire [4-1:0] node36848;
	wire [4-1:0] node36850;
	wire [4-1:0] node36853;
	wire [4-1:0] node36854;
	wire [4-1:0] node36857;
	wire [4-1:0] node36860;
	wire [4-1:0] node36861;
	wire [4-1:0] node36865;
	wire [4-1:0] node36866;
	wire [4-1:0] node36867;
	wire [4-1:0] node36869;
	wire [4-1:0] node36872;
	wire [4-1:0] node36873;
	wire [4-1:0] node36877;
	wire [4-1:0] node36878;
	wire [4-1:0] node36879;
	wire [4-1:0] node36883;
	wire [4-1:0] node36886;
	wire [4-1:0] node36887;
	wire [4-1:0] node36888;
	wire [4-1:0] node36889;
	wire [4-1:0] node36890;
	wire [4-1:0] node36894;
	wire [4-1:0] node36896;
	wire [4-1:0] node36898;
	wire [4-1:0] node36901;
	wire [4-1:0] node36902;
	wire [4-1:0] node36903;
	wire [4-1:0] node36905;
	wire [4-1:0] node36908;
	wire [4-1:0] node36909;
	wire [4-1:0] node36913;
	wire [4-1:0] node36914;
	wire [4-1:0] node36916;
	wire [4-1:0] node36920;
	wire [4-1:0] node36921;
	wire [4-1:0] node36922;
	wire [4-1:0] node36923;
	wire [4-1:0] node36926;
	wire [4-1:0] node36927;
	wire [4-1:0] node36931;
	wire [4-1:0] node36933;
	wire [4-1:0] node36936;
	wire [4-1:0] node36937;
	wire [4-1:0] node36938;
	wire [4-1:0] node36939;
	wire [4-1:0] node36942;
	wire [4-1:0] node36946;
	wire [4-1:0] node36947;
	wire [4-1:0] node36951;
	wire [4-1:0] node36952;
	wire [4-1:0] node36953;
	wire [4-1:0] node36954;
	wire [4-1:0] node36956;
	wire [4-1:0] node36957;
	wire [4-1:0] node36959;
	wire [4-1:0] node36963;
	wire [4-1:0] node36964;
	wire [4-1:0] node36965;
	wire [4-1:0] node36969;
	wire [4-1:0] node36970;
	wire [4-1:0] node36973;
	wire [4-1:0] node36976;
	wire [4-1:0] node36977;
	wire [4-1:0] node36978;
	wire [4-1:0] node36979;
	wire [4-1:0] node36980;
	wire [4-1:0] node36983;
	wire [4-1:0] node36986;
	wire [4-1:0] node36987;
	wire [4-1:0] node36990;
	wire [4-1:0] node36993;
	wire [4-1:0] node36995;
	wire [4-1:0] node36996;
	wire [4-1:0] node37000;
	wire [4-1:0] node37001;
	wire [4-1:0] node37003;
	wire [4-1:0] node37004;
	wire [4-1:0] node37007;
	wire [4-1:0] node37010;
	wire [4-1:0] node37013;
	wire [4-1:0] node37014;
	wire [4-1:0] node37015;
	wire [4-1:0] node37016;
	wire [4-1:0] node37017;
	wire [4-1:0] node37019;
	wire [4-1:0] node37022;
	wire [4-1:0] node37023;
	wire [4-1:0] node37027;
	wire [4-1:0] node37028;
	wire [4-1:0] node37031;
	wire [4-1:0] node37034;
	wire [4-1:0] node37035;
	wire [4-1:0] node37036;
	wire [4-1:0] node37037;
	wire [4-1:0] node37040;
	wire [4-1:0] node37043;
	wire [4-1:0] node37046;
	wire [4-1:0] node37048;
	wire [4-1:0] node37051;
	wire [4-1:0] node37052;
	wire [4-1:0] node37053;
	wire [4-1:0] node37054;
	wire [4-1:0] node37055;
	wire [4-1:0] node37059;
	wire [4-1:0] node37060;
	wire [4-1:0] node37063;
	wire [4-1:0] node37066;
	wire [4-1:0] node37067;
	wire [4-1:0] node37068;
	wire [4-1:0] node37071;
	wire [4-1:0] node37074;
	wire [4-1:0] node37075;
	wire [4-1:0] node37078;
	wire [4-1:0] node37081;
	wire [4-1:0] node37082;
	wire [4-1:0] node37084;
	wire [4-1:0] node37085;
	wire [4-1:0] node37089;
	wire [4-1:0] node37092;
	wire [4-1:0] node37093;
	wire [4-1:0] node37094;
	wire [4-1:0] node37095;
	wire [4-1:0] node37096;
	wire [4-1:0] node37097;
	wire [4-1:0] node37099;
	wire [4-1:0] node37101;
	wire [4-1:0] node37104;
	wire [4-1:0] node37105;
	wire [4-1:0] node37108;
	wire [4-1:0] node37111;
	wire [4-1:0] node37112;
	wire [4-1:0] node37113;
	wire [4-1:0] node37117;
	wire [4-1:0] node37118;
	wire [4-1:0] node37121;
	wire [4-1:0] node37124;
	wire [4-1:0] node37125;
	wire [4-1:0] node37126;
	wire [4-1:0] node37129;
	wire [4-1:0] node37132;
	wire [4-1:0] node37133;
	wire [4-1:0] node37134;
	wire [4-1:0] node37137;
	wire [4-1:0] node37140;
	wire [4-1:0] node37141;
	wire [4-1:0] node37145;
	wire [4-1:0] node37146;
	wire [4-1:0] node37147;
	wire [4-1:0] node37148;
	wire [4-1:0] node37149;
	wire [4-1:0] node37152;
	wire [4-1:0] node37155;
	wire [4-1:0] node37156;
	wire [4-1:0] node37159;
	wire [4-1:0] node37162;
	wire [4-1:0] node37163;
	wire [4-1:0] node37164;
	wire [4-1:0] node37168;
	wire [4-1:0] node37169;
	wire [4-1:0] node37172;
	wire [4-1:0] node37175;
	wire [4-1:0] node37176;
	wire [4-1:0] node37177;
	wire [4-1:0] node37180;
	wire [4-1:0] node37182;
	wire [4-1:0] node37185;
	wire [4-1:0] node37186;
	wire [4-1:0] node37187;
	wire [4-1:0] node37190;
	wire [4-1:0] node37194;
	wire [4-1:0] node37195;
	wire [4-1:0] node37196;
	wire [4-1:0] node37197;
	wire [4-1:0] node37198;
	wire [4-1:0] node37199;
	wire [4-1:0] node37201;
	wire [4-1:0] node37204;
	wire [4-1:0] node37207;
	wire [4-1:0] node37208;
	wire [4-1:0] node37211;
	wire [4-1:0] node37212;
	wire [4-1:0] node37215;
	wire [4-1:0] node37218;
	wire [4-1:0] node37219;
	wire [4-1:0] node37220;
	wire [4-1:0] node37221;
	wire [4-1:0] node37226;
	wire [4-1:0] node37227;
	wire [4-1:0] node37230;
	wire [4-1:0] node37233;
	wire [4-1:0] node37234;
	wire [4-1:0] node37235;
	wire [4-1:0] node37236;
	wire [4-1:0] node37238;
	wire [4-1:0] node37241;
	wire [4-1:0] node37244;
	wire [4-1:0] node37246;
	wire [4-1:0] node37247;
	wire [4-1:0] node37251;
	wire [4-1:0] node37253;
	wire [4-1:0] node37254;
	wire [4-1:0] node37255;
	wire [4-1:0] node37259;
	wire [4-1:0] node37262;
	wire [4-1:0] node37263;
	wire [4-1:0] node37264;
	wire [4-1:0] node37265;
	wire [4-1:0] node37266;
	wire [4-1:0] node37269;
	wire [4-1:0] node37273;
	wire [4-1:0] node37274;
	wire [4-1:0] node37275;
	wire [4-1:0] node37276;
	wire [4-1:0] node37280;
	wire [4-1:0] node37281;
	wire [4-1:0] node37285;
	wire [4-1:0] node37287;
	wire [4-1:0] node37288;
	wire [4-1:0] node37291;
	wire [4-1:0] node37294;
	wire [4-1:0] node37295;
	wire [4-1:0] node37296;
	wire [4-1:0] node37297;
	wire [4-1:0] node37298;
	wire [4-1:0] node37301;
	wire [4-1:0] node37304;
	wire [4-1:0] node37305;
	wire [4-1:0] node37308;
	wire [4-1:0] node37311;
	wire [4-1:0] node37312;
	wire [4-1:0] node37314;
	wire [4-1:0] node37317;
	wire [4-1:0] node37318;
	wire [4-1:0] node37321;
	wire [4-1:0] node37324;
	wire [4-1:0] node37325;
	wire [4-1:0] node37326;
	wire [4-1:0] node37328;
	wire [4-1:0] node37332;
	wire [4-1:0] node37333;
	wire [4-1:0] node37334;
	wire [4-1:0] node37337;
	wire [4-1:0] node37340;
	wire [4-1:0] node37341;
	wire [4-1:0] node37345;
	wire [4-1:0] node37346;
	wire [4-1:0] node37347;
	wire [4-1:0] node37348;
	wire [4-1:0] node37349;
	wire [4-1:0] node37350;
	wire [4-1:0] node37351;
	wire [4-1:0] node37352;
	wire [4-1:0] node37355;
	wire [4-1:0] node37357;
	wire [4-1:0] node37360;
	wire [4-1:0] node37361;
	wire [4-1:0] node37362;
	wire [4-1:0] node37366;
	wire [4-1:0] node37369;
	wire [4-1:0] node37370;
	wire [4-1:0] node37371;
	wire [4-1:0] node37372;
	wire [4-1:0] node37375;
	wire [4-1:0] node37378;
	wire [4-1:0] node37379;
	wire [4-1:0] node37382;
	wire [4-1:0] node37385;
	wire [4-1:0] node37386;
	wire [4-1:0] node37387;
	wire [4-1:0] node37390;
	wire [4-1:0] node37393;
	wire [4-1:0] node37395;
	wire [4-1:0] node37398;
	wire [4-1:0] node37399;
	wire [4-1:0] node37400;
	wire [4-1:0] node37402;
	wire [4-1:0] node37405;
	wire [4-1:0] node37406;
	wire [4-1:0] node37409;
	wire [4-1:0] node37412;
	wire [4-1:0] node37413;
	wire [4-1:0] node37415;
	wire [4-1:0] node37418;
	wire [4-1:0] node37420;
	wire [4-1:0] node37423;
	wire [4-1:0] node37424;
	wire [4-1:0] node37425;
	wire [4-1:0] node37426;
	wire [4-1:0] node37428;
	wire [4-1:0] node37429;
	wire [4-1:0] node37432;
	wire [4-1:0] node37435;
	wire [4-1:0] node37436;
	wire [4-1:0] node37439;
	wire [4-1:0] node37440;
	wire [4-1:0] node37443;
	wire [4-1:0] node37446;
	wire [4-1:0] node37447;
	wire [4-1:0] node37448;
	wire [4-1:0] node37449;
	wire [4-1:0] node37453;
	wire [4-1:0] node37456;
	wire [4-1:0] node37457;
	wire [4-1:0] node37460;
	wire [4-1:0] node37463;
	wire [4-1:0] node37464;
	wire [4-1:0] node37465;
	wire [4-1:0] node37466;
	wire [4-1:0] node37468;
	wire [4-1:0] node37471;
	wire [4-1:0] node37472;
	wire [4-1:0] node37476;
	wire [4-1:0] node37478;
	wire [4-1:0] node37480;
	wire [4-1:0] node37483;
	wire [4-1:0] node37484;
	wire [4-1:0] node37486;
	wire [4-1:0] node37490;
	wire [4-1:0] node37491;
	wire [4-1:0] node37492;
	wire [4-1:0] node37493;
	wire [4-1:0] node37494;
	wire [4-1:0] node37495;
	wire [4-1:0] node37497;
	wire [4-1:0] node37501;
	wire [4-1:0] node37504;
	wire [4-1:0] node37505;
	wire [4-1:0] node37506;
	wire [4-1:0] node37509;
	wire [4-1:0] node37512;
	wire [4-1:0] node37513;
	wire [4-1:0] node37515;
	wire [4-1:0] node37518;
	wire [4-1:0] node37519;
	wire [4-1:0] node37523;
	wire [4-1:0] node37524;
	wire [4-1:0] node37525;
	wire [4-1:0] node37527;
	wire [4-1:0] node37528;
	wire [4-1:0] node37531;
	wire [4-1:0] node37534;
	wire [4-1:0] node37535;
	wire [4-1:0] node37536;
	wire [4-1:0] node37539;
	wire [4-1:0] node37543;
	wire [4-1:0] node37545;
	wire [4-1:0] node37546;
	wire [4-1:0] node37550;
	wire [4-1:0] node37551;
	wire [4-1:0] node37552;
	wire [4-1:0] node37553;
	wire [4-1:0] node37555;
	wire [4-1:0] node37558;
	wire [4-1:0] node37560;
	wire [4-1:0] node37563;
	wire [4-1:0] node37564;
	wire [4-1:0] node37565;
	wire [4-1:0] node37566;
	wire [4-1:0] node37569;
	wire [4-1:0] node37573;
	wire [4-1:0] node37575;
	wire [4-1:0] node37578;
	wire [4-1:0] node37579;
	wire [4-1:0] node37580;
	wire [4-1:0] node37583;
	wire [4-1:0] node37584;
	wire [4-1:0] node37585;
	wire [4-1:0] node37590;
	wire [4-1:0] node37591;
	wire [4-1:0] node37593;
	wire [4-1:0] node37594;
	wire [4-1:0] node37598;
	wire [4-1:0] node37599;
	wire [4-1:0] node37600;
	wire [4-1:0] node37605;
	wire [4-1:0] node37606;
	wire [4-1:0] node37607;
	wire [4-1:0] node37608;
	wire [4-1:0] node37609;
	wire [4-1:0] node37610;
	wire [4-1:0] node37611;
	wire [4-1:0] node37612;
	wire [4-1:0] node37615;
	wire [4-1:0] node37618;
	wire [4-1:0] node37619;
	wire [4-1:0] node37622;
	wire [4-1:0] node37625;
	wire [4-1:0] node37627;
	wire [4-1:0] node37630;
	wire [4-1:0] node37631;
	wire [4-1:0] node37632;
	wire [4-1:0] node37633;
	wire [4-1:0] node37637;
	wire [4-1:0] node37638;
	wire [4-1:0] node37642;
	wire [4-1:0] node37643;
	wire [4-1:0] node37644;
	wire [4-1:0] node37647;
	wire [4-1:0] node37650;
	wire [4-1:0] node37651;
	wire [4-1:0] node37655;
	wire [4-1:0] node37656;
	wire [4-1:0] node37657;
	wire [4-1:0] node37658;
	wire [4-1:0] node37661;
	wire [4-1:0] node37662;
	wire [4-1:0] node37666;
	wire [4-1:0] node37667;
	wire [4-1:0] node37668;
	wire [4-1:0] node37671;
	wire [4-1:0] node37674;
	wire [4-1:0] node37676;
	wire [4-1:0] node37679;
	wire [4-1:0] node37680;
	wire [4-1:0] node37681;
	wire [4-1:0] node37682;
	wire [4-1:0] node37685;
	wire [4-1:0] node37688;
	wire [4-1:0] node37691;
	wire [4-1:0] node37692;
	wire [4-1:0] node37694;
	wire [4-1:0] node37698;
	wire [4-1:0] node37699;
	wire [4-1:0] node37700;
	wire [4-1:0] node37701;
	wire [4-1:0] node37702;
	wire [4-1:0] node37705;
	wire [4-1:0] node37708;
	wire [4-1:0] node37710;
	wire [4-1:0] node37713;
	wire [4-1:0] node37714;
	wire [4-1:0] node37715;
	wire [4-1:0] node37718;
	wire [4-1:0] node37721;
	wire [4-1:0] node37724;
	wire [4-1:0] node37725;
	wire [4-1:0] node37726;
	wire [4-1:0] node37727;
	wire [4-1:0] node37728;
	wire [4-1:0] node37732;
	wire [4-1:0] node37733;
	wire [4-1:0] node37737;
	wire [4-1:0] node37738;
	wire [4-1:0] node37740;
	wire [4-1:0] node37744;
	wire [4-1:0] node37745;
	wire [4-1:0] node37747;
	wire [4-1:0] node37748;
	wire [4-1:0] node37751;
	wire [4-1:0] node37754;
	wire [4-1:0] node37755;
	wire [4-1:0] node37756;
	wire [4-1:0] node37759;
	wire [4-1:0] node37762;
	wire [4-1:0] node37763;
	wire [4-1:0] node37767;
	wire [4-1:0] node37768;
	wire [4-1:0] node37769;
	wire [4-1:0] node37770;
	wire [4-1:0] node37771;
	wire [4-1:0] node37772;
	wire [4-1:0] node37775;
	wire [4-1:0] node37778;
	wire [4-1:0] node37781;
	wire [4-1:0] node37782;
	wire [4-1:0] node37785;
	wire [4-1:0] node37788;
	wire [4-1:0] node37789;
	wire [4-1:0] node37790;
	wire [4-1:0] node37791;
	wire [4-1:0] node37794;
	wire [4-1:0] node37797;
	wire [4-1:0] node37798;
	wire [4-1:0] node37801;
	wire [4-1:0] node37804;
	wire [4-1:0] node37805;
	wire [4-1:0] node37806;
	wire [4-1:0] node37809;
	wire [4-1:0] node37812;
	wire [4-1:0] node37815;
	wire [4-1:0] node37816;
	wire [4-1:0] node37817;
	wire [4-1:0] node37818;
	wire [4-1:0] node37819;
	wire [4-1:0] node37823;
	wire [4-1:0] node37824;
	wire [4-1:0] node37827;
	wire [4-1:0] node37830;
	wire [4-1:0] node37831;
	wire [4-1:0] node37832;
	wire [4-1:0] node37833;
	wire [4-1:0] node37837;
	wire [4-1:0] node37838;
	wire [4-1:0] node37843;
	wire [4-1:0] node37844;
	wire [4-1:0] node37845;
	wire [4-1:0] node37846;
	wire [4-1:0] node37850;
	wire [4-1:0] node37851;
	wire [4-1:0] node37854;
	wire [4-1:0] node37857;
	wire [4-1:0] node37858;
	wire [4-1:0] node37859;
	wire [4-1:0] node37860;
	wire [4-1:0] node37865;
	wire [4-1:0] node37866;
	wire [4-1:0] node37870;
	wire [4-1:0] node37871;
	wire [4-1:0] node37872;
	wire [4-1:0] node37873;
	wire [4-1:0] node37874;
	wire [4-1:0] node37875;
	wire [4-1:0] node37876;
	wire [4-1:0] node37877;
	wire [4-1:0] node37878;
	wire [4-1:0] node37879;
	wire [4-1:0] node37882;
	wire [4-1:0] node37885;
	wire [4-1:0] node37886;
	wire [4-1:0] node37890;
	wire [4-1:0] node37892;
	wire [4-1:0] node37894;
	wire [4-1:0] node37897;
	wire [4-1:0] node37898;
	wire [4-1:0] node37899;
	wire [4-1:0] node37900;
	wire [4-1:0] node37903;
	wire [4-1:0] node37904;
	wire [4-1:0] node37907;
	wire [4-1:0] node37910;
	wire [4-1:0] node37911;
	wire [4-1:0] node37914;
	wire [4-1:0] node37916;
	wire [4-1:0] node37919;
	wire [4-1:0] node37920;
	wire [4-1:0] node37922;
	wire [4-1:0] node37925;
	wire [4-1:0] node37927;
	wire [4-1:0] node37928;
	wire [4-1:0] node37931;
	wire [4-1:0] node37934;
	wire [4-1:0] node37935;
	wire [4-1:0] node37936;
	wire [4-1:0] node37937;
	wire [4-1:0] node37938;
	wire [4-1:0] node37942;
	wire [4-1:0] node37945;
	wire [4-1:0] node37946;
	wire [4-1:0] node37948;
	wire [4-1:0] node37950;
	wire [4-1:0] node37953;
	wire [4-1:0] node37954;
	wire [4-1:0] node37955;
	wire [4-1:0] node37959;
	wire [4-1:0] node37962;
	wire [4-1:0] node37963;
	wire [4-1:0] node37964;
	wire [4-1:0] node37966;
	wire [4-1:0] node37968;
	wire [4-1:0] node37971;
	wire [4-1:0] node37972;
	wire [4-1:0] node37973;
	wire [4-1:0] node37977;
	wire [4-1:0] node37978;
	wire [4-1:0] node37981;
	wire [4-1:0] node37984;
	wire [4-1:0] node37985;
	wire [4-1:0] node37987;
	wire [4-1:0] node37988;
	wire [4-1:0] node37992;
	wire [4-1:0] node37993;
	wire [4-1:0] node37997;
	wire [4-1:0] node37998;
	wire [4-1:0] node37999;
	wire [4-1:0] node38000;
	wire [4-1:0] node38001;
	wire [4-1:0] node38002;
	wire [4-1:0] node38005;
	wire [4-1:0] node38007;
	wire [4-1:0] node38010;
	wire [4-1:0] node38012;
	wire [4-1:0] node38013;
	wire [4-1:0] node38016;
	wire [4-1:0] node38019;
	wire [4-1:0] node38020;
	wire [4-1:0] node38021;
	wire [4-1:0] node38022;
	wire [4-1:0] node38026;
	wire [4-1:0] node38029;
	wire [4-1:0] node38030;
	wire [4-1:0] node38031;
	wire [4-1:0] node38034;
	wire [4-1:0] node38037;
	wire [4-1:0] node38040;
	wire [4-1:0] node38041;
	wire [4-1:0] node38042;
	wire [4-1:0] node38043;
	wire [4-1:0] node38044;
	wire [4-1:0] node38047;
	wire [4-1:0] node38050;
	wire [4-1:0] node38053;
	wire [4-1:0] node38054;
	wire [4-1:0] node38055;
	wire [4-1:0] node38058;
	wire [4-1:0] node38061;
	wire [4-1:0] node38064;
	wire [4-1:0] node38065;
	wire [4-1:0] node38066;
	wire [4-1:0] node38067;
	wire [4-1:0] node38070;
	wire [4-1:0] node38073;
	wire [4-1:0] node38074;
	wire [4-1:0] node38077;
	wire [4-1:0] node38080;
	wire [4-1:0] node38081;
	wire [4-1:0] node38082;
	wire [4-1:0] node38085;
	wire [4-1:0] node38088;
	wire [4-1:0] node38089;
	wire [4-1:0] node38093;
	wire [4-1:0] node38094;
	wire [4-1:0] node38095;
	wire [4-1:0] node38096;
	wire [4-1:0] node38097;
	wire [4-1:0] node38098;
	wire [4-1:0] node38103;
	wire [4-1:0] node38105;
	wire [4-1:0] node38108;
	wire [4-1:0] node38109;
	wire [4-1:0] node38110;
	wire [4-1:0] node38112;
	wire [4-1:0] node38115;
	wire [4-1:0] node38118;
	wire [4-1:0] node38119;
	wire [4-1:0] node38120;
	wire [4-1:0] node38124;
	wire [4-1:0] node38125;
	wire [4-1:0] node38129;
	wire [4-1:0] node38130;
	wire [4-1:0] node38131;
	wire [4-1:0] node38132;
	wire [4-1:0] node38133;
	wire [4-1:0] node38137;
	wire [4-1:0] node38138;
	wire [4-1:0] node38142;
	wire [4-1:0] node38143;
	wire [4-1:0] node38144;
	wire [4-1:0] node38147;
	wire [4-1:0] node38150;
	wire [4-1:0] node38151;
	wire [4-1:0] node38154;
	wire [4-1:0] node38157;
	wire [4-1:0] node38158;
	wire [4-1:0] node38159;
	wire [4-1:0] node38160;
	wire [4-1:0] node38165;
	wire [4-1:0] node38167;
	wire [4-1:0] node38168;
	wire [4-1:0] node38171;
	wire [4-1:0] node38174;
	wire [4-1:0] node38175;
	wire [4-1:0] node38176;
	wire [4-1:0] node38177;
	wire [4-1:0] node38178;
	wire [4-1:0] node38179;
	wire [4-1:0] node38180;
	wire [4-1:0] node38181;
	wire [4-1:0] node38186;
	wire [4-1:0] node38187;
	wire [4-1:0] node38188;
	wire [4-1:0] node38191;
	wire [4-1:0] node38194;
	wire [4-1:0] node38196;
	wire [4-1:0] node38199;
	wire [4-1:0] node38200;
	wire [4-1:0] node38202;
	wire [4-1:0] node38203;
	wire [4-1:0] node38207;
	wire [4-1:0] node38208;
	wire [4-1:0] node38209;
	wire [4-1:0] node38212;
	wire [4-1:0] node38215;
	wire [4-1:0] node38217;
	wire [4-1:0] node38220;
	wire [4-1:0] node38221;
	wire [4-1:0] node38222;
	wire [4-1:0] node38223;
	wire [4-1:0] node38224;
	wire [4-1:0] node38229;
	wire [4-1:0] node38231;
	wire [4-1:0] node38234;
	wire [4-1:0] node38235;
	wire [4-1:0] node38238;
	wire [4-1:0] node38239;
	wire [4-1:0] node38240;
	wire [4-1:0] node38244;
	wire [4-1:0] node38245;
	wire [4-1:0] node38248;
	wire [4-1:0] node38251;
	wire [4-1:0] node38252;
	wire [4-1:0] node38253;
	wire [4-1:0] node38254;
	wire [4-1:0] node38257;
	wire [4-1:0] node38259;
	wire [4-1:0] node38262;
	wire [4-1:0] node38263;
	wire [4-1:0] node38264;
	wire [4-1:0] node38267;
	wire [4-1:0] node38269;
	wire [4-1:0] node38272;
	wire [4-1:0] node38273;
	wire [4-1:0] node38277;
	wire [4-1:0] node38278;
	wire [4-1:0] node38279;
	wire [4-1:0] node38282;
	wire [4-1:0] node38283;
	wire [4-1:0] node38284;
	wire [4-1:0] node38287;
	wire [4-1:0] node38290;
	wire [4-1:0] node38293;
	wire [4-1:0] node38294;
	wire [4-1:0] node38295;
	wire [4-1:0] node38296;
	wire [4-1:0] node38300;
	wire [4-1:0] node38302;
	wire [4-1:0] node38305;
	wire [4-1:0] node38306;
	wire [4-1:0] node38309;
	wire [4-1:0] node38312;
	wire [4-1:0] node38313;
	wire [4-1:0] node38314;
	wire [4-1:0] node38315;
	wire [4-1:0] node38316;
	wire [4-1:0] node38317;
	wire [4-1:0] node38319;
	wire [4-1:0] node38323;
	wire [4-1:0] node38325;
	wire [4-1:0] node38326;
	wire [4-1:0] node38330;
	wire [4-1:0] node38331;
	wire [4-1:0] node38332;
	wire [4-1:0] node38333;
	wire [4-1:0] node38337;
	wire [4-1:0] node38341;
	wire [4-1:0] node38342;
	wire [4-1:0] node38343;
	wire [4-1:0] node38345;
	wire [4-1:0] node38346;
	wire [4-1:0] node38350;
	wire [4-1:0] node38351;
	wire [4-1:0] node38352;
	wire [4-1:0] node38355;
	wire [4-1:0] node38358;
	wire [4-1:0] node38359;
	wire [4-1:0] node38362;
	wire [4-1:0] node38365;
	wire [4-1:0] node38366;
	wire [4-1:0] node38368;
	wire [4-1:0] node38369;
	wire [4-1:0] node38373;
	wire [4-1:0] node38374;
	wire [4-1:0] node38375;
	wire [4-1:0] node38378;
	wire [4-1:0] node38382;
	wire [4-1:0] node38383;
	wire [4-1:0] node38384;
	wire [4-1:0] node38385;
	wire [4-1:0] node38386;
	wire [4-1:0] node38387;
	wire [4-1:0] node38391;
	wire [4-1:0] node38394;
	wire [4-1:0] node38396;
	wire [4-1:0] node38397;
	wire [4-1:0] node38401;
	wire [4-1:0] node38402;
	wire [4-1:0] node38405;
	wire [4-1:0] node38408;
	wire [4-1:0] node38409;
	wire [4-1:0] node38410;
	wire [4-1:0] node38411;
	wire [4-1:0] node38412;
	wire [4-1:0] node38416;
	wire [4-1:0] node38418;
	wire [4-1:0] node38421;
	wire [4-1:0] node38422;
	wire [4-1:0] node38425;
	wire [4-1:0] node38426;
	wire [4-1:0] node38429;
	wire [4-1:0] node38432;
	wire [4-1:0] node38433;
	wire [4-1:0] node38434;
	wire [4-1:0] node38435;
	wire [4-1:0] node38439;
	wire [4-1:0] node38441;
	wire [4-1:0] node38444;
	wire [4-1:0] node38445;
	wire [4-1:0] node38446;
	wire [4-1:0] node38450;
	wire [4-1:0] node38453;
	wire [4-1:0] node38454;
	wire [4-1:0] node38455;
	wire [4-1:0] node38456;
	wire [4-1:0] node38457;
	wire [4-1:0] node38458;
	wire [4-1:0] node38459;
	wire [4-1:0] node38460;
	wire [4-1:0] node38461;
	wire [4-1:0] node38465;
	wire [4-1:0] node38467;
	wire [4-1:0] node38470;
	wire [4-1:0] node38471;
	wire [4-1:0] node38474;
	wire [4-1:0] node38477;
	wire [4-1:0] node38478;
	wire [4-1:0] node38480;
	wire [4-1:0] node38482;
	wire [4-1:0] node38485;
	wire [4-1:0] node38486;
	wire [4-1:0] node38487;
	wire [4-1:0] node38490;
	wire [4-1:0] node38494;
	wire [4-1:0] node38495;
	wire [4-1:0] node38496;
	wire [4-1:0] node38498;
	wire [4-1:0] node38501;
	wire [4-1:0] node38503;
	wire [4-1:0] node38506;
	wire [4-1:0] node38507;
	wire [4-1:0] node38508;
	wire [4-1:0] node38509;
	wire [4-1:0] node38512;
	wire [4-1:0] node38516;
	wire [4-1:0] node38517;
	wire [4-1:0] node38521;
	wire [4-1:0] node38522;
	wire [4-1:0] node38523;
	wire [4-1:0] node38524;
	wire [4-1:0] node38525;
	wire [4-1:0] node38527;
	wire [4-1:0] node38530;
	wire [4-1:0] node38531;
	wire [4-1:0] node38535;
	wire [4-1:0] node38536;
	wire [4-1:0] node38538;
	wire [4-1:0] node38542;
	wire [4-1:0] node38543;
	wire [4-1:0] node38544;
	wire [4-1:0] node38548;
	wire [4-1:0] node38549;
	wire [4-1:0] node38553;
	wire [4-1:0] node38554;
	wire [4-1:0] node38555;
	wire [4-1:0] node38556;
	wire [4-1:0] node38560;
	wire [4-1:0] node38561;
	wire [4-1:0] node38563;
	wire [4-1:0] node38567;
	wire [4-1:0] node38568;
	wire [4-1:0] node38569;
	wire [4-1:0] node38571;
	wire [4-1:0] node38574;
	wire [4-1:0] node38576;
	wire [4-1:0] node38579;
	wire [4-1:0] node38581;
	wire [4-1:0] node38582;
	wire [4-1:0] node38585;
	wire [4-1:0] node38588;
	wire [4-1:0] node38589;
	wire [4-1:0] node38590;
	wire [4-1:0] node38591;
	wire [4-1:0] node38592;
	wire [4-1:0] node38593;
	wire [4-1:0] node38594;
	wire [4-1:0] node38598;
	wire [4-1:0] node38600;
	wire [4-1:0] node38603;
	wire [4-1:0] node38605;
	wire [4-1:0] node38606;
	wire [4-1:0] node38609;
	wire [4-1:0] node38612;
	wire [4-1:0] node38613;
	wire [4-1:0] node38614;
	wire [4-1:0] node38618;
	wire [4-1:0] node38619;
	wire [4-1:0] node38620;
	wire [4-1:0] node38623;
	wire [4-1:0] node38627;
	wire [4-1:0] node38628;
	wire [4-1:0] node38629;
	wire [4-1:0] node38630;
	wire [4-1:0] node38633;
	wire [4-1:0] node38635;
	wire [4-1:0] node38638;
	wire [4-1:0] node38641;
	wire [4-1:0] node38642;
	wire [4-1:0] node38643;
	wire [4-1:0] node38644;
	wire [4-1:0] node38649;
	wire [4-1:0] node38650;
	wire [4-1:0] node38652;
	wire [4-1:0] node38655;
	wire [4-1:0] node38656;
	wire [4-1:0] node38659;
	wire [4-1:0] node38662;
	wire [4-1:0] node38663;
	wire [4-1:0] node38664;
	wire [4-1:0] node38665;
	wire [4-1:0] node38666;
	wire [4-1:0] node38669;
	wire [4-1:0] node38672;
	wire [4-1:0] node38673;
	wire [4-1:0] node38674;
	wire [4-1:0] node38677;
	wire [4-1:0] node38680;
	wire [4-1:0] node38682;
	wire [4-1:0] node38685;
	wire [4-1:0] node38686;
	wire [4-1:0] node38687;
	wire [4-1:0] node38691;
	wire [4-1:0] node38693;
	wire [4-1:0] node38696;
	wire [4-1:0] node38697;
	wire [4-1:0] node38698;
	wire [4-1:0] node38701;
	wire [4-1:0] node38702;
	wire [4-1:0] node38703;
	wire [4-1:0] node38708;
	wire [4-1:0] node38709;
	wire [4-1:0] node38711;
	wire [4-1:0] node38712;
	wire [4-1:0] node38715;
	wire [4-1:0] node38718;
	wire [4-1:0] node38720;
	wire [4-1:0] node38723;
	wire [4-1:0] node38724;
	wire [4-1:0] node38725;
	wire [4-1:0] node38726;
	wire [4-1:0] node38727;
	wire [4-1:0] node38728;
	wire [4-1:0] node38730;
	wire [4-1:0] node38733;
	wire [4-1:0] node38734;
	wire [4-1:0] node38737;
	wire [4-1:0] node38740;
	wire [4-1:0] node38741;
	wire [4-1:0] node38742;
	wire [4-1:0] node38746;
	wire [4-1:0] node38748;
	wire [4-1:0] node38751;
	wire [4-1:0] node38752;
	wire [4-1:0] node38753;
	wire [4-1:0] node38754;
	wire [4-1:0] node38756;
	wire [4-1:0] node38759;
	wire [4-1:0] node38761;
	wire [4-1:0] node38764;
	wire [4-1:0] node38765;
	wire [4-1:0] node38766;
	wire [4-1:0] node38769;
	wire [4-1:0] node38773;
	wire [4-1:0] node38774;
	wire [4-1:0] node38775;
	wire [4-1:0] node38779;
	wire [4-1:0] node38780;
	wire [4-1:0] node38784;
	wire [4-1:0] node38785;
	wire [4-1:0] node38786;
	wire [4-1:0] node38787;
	wire [4-1:0] node38788;
	wire [4-1:0] node38792;
	wire [4-1:0] node38793;
	wire [4-1:0] node38797;
	wire [4-1:0] node38798;
	wire [4-1:0] node38799;
	wire [4-1:0] node38800;
	wire [4-1:0] node38803;
	wire [4-1:0] node38806;
	wire [4-1:0] node38807;
	wire [4-1:0] node38811;
	wire [4-1:0] node38813;
	wire [4-1:0] node38816;
	wire [4-1:0] node38817;
	wire [4-1:0] node38818;
	wire [4-1:0] node38821;
	wire [4-1:0] node38823;
	wire [4-1:0] node38825;
	wire [4-1:0] node38828;
	wire [4-1:0] node38829;
	wire [4-1:0] node38830;
	wire [4-1:0] node38831;
	wire [4-1:0] node38834;
	wire [4-1:0] node38838;
	wire [4-1:0] node38840;
	wire [4-1:0] node38843;
	wire [4-1:0] node38844;
	wire [4-1:0] node38845;
	wire [4-1:0] node38846;
	wire [4-1:0] node38847;
	wire [4-1:0] node38850;
	wire [4-1:0] node38852;
	wire [4-1:0] node38855;
	wire [4-1:0] node38856;
	wire [4-1:0] node38857;
	wire [4-1:0] node38859;
	wire [4-1:0] node38862;
	wire [4-1:0] node38863;
	wire [4-1:0] node38867;
	wire [4-1:0] node38870;
	wire [4-1:0] node38871;
	wire [4-1:0] node38872;
	wire [4-1:0] node38873;
	wire [4-1:0] node38874;
	wire [4-1:0] node38877;
	wire [4-1:0] node38880;
	wire [4-1:0] node38881;
	wire [4-1:0] node38885;
	wire [4-1:0] node38886;
	wire [4-1:0] node38889;
	wire [4-1:0] node38892;
	wire [4-1:0] node38893;
	wire [4-1:0] node38895;
	wire [4-1:0] node38898;
	wire [4-1:0] node38901;
	wire [4-1:0] node38902;
	wire [4-1:0] node38903;
	wire [4-1:0] node38904;
	wire [4-1:0] node38905;
	wire [4-1:0] node38907;
	wire [4-1:0] node38910;
	wire [4-1:0] node38911;
	wire [4-1:0] node38914;
	wire [4-1:0] node38917;
	wire [4-1:0] node38918;
	wire [4-1:0] node38920;
	wire [4-1:0] node38923;
	wire [4-1:0] node38925;
	wire [4-1:0] node38928;
	wire [4-1:0] node38929;
	wire [4-1:0] node38930;
	wire [4-1:0] node38931;
	wire [4-1:0] node38934;
	wire [4-1:0] node38938;
	wire [4-1:0] node38940;
	wire [4-1:0] node38943;
	wire [4-1:0] node38944;
	wire [4-1:0] node38945;
	wire [4-1:0] node38947;
	wire [4-1:0] node38950;
	wire [4-1:0] node38951;
	wire [4-1:0] node38955;
	wire [4-1:0] node38956;
	wire [4-1:0] node38957;
	wire [4-1:0] node38960;
	wire [4-1:0] node38963;
	wire [4-1:0] node38964;
	wire [4-1:0] node38965;
	wire [4-1:0] node38968;
	wire [4-1:0] node38971;
	wire [4-1:0] node38973;
	wire [4-1:0] node38976;
	wire [4-1:0] node38977;
	wire [4-1:0] node38978;
	wire [4-1:0] node38979;
	wire [4-1:0] node38980;
	wire [4-1:0] node38981;
	wire [4-1:0] node38982;
	wire [4-1:0] node38983;
	wire [4-1:0] node38984;
	wire [4-1:0] node38985;
	wire [4-1:0] node38988;
	wire [4-1:0] node38992;
	wire [4-1:0] node38993;
	wire [4-1:0] node38995;
	wire [4-1:0] node38999;
	wire [4-1:0] node39001;
	wire [4-1:0] node39003;
	wire [4-1:0] node39005;
	wire [4-1:0] node39008;
	wire [4-1:0] node39009;
	wire [4-1:0] node39010;
	wire [4-1:0] node39011;
	wire [4-1:0] node39015;
	wire [4-1:0] node39016;
	wire [4-1:0] node39017;
	wire [4-1:0] node39020;
	wire [4-1:0] node39023;
	wire [4-1:0] node39025;
	wire [4-1:0] node39028;
	wire [4-1:0] node39029;
	wire [4-1:0] node39031;
	wire [4-1:0] node39034;
	wire [4-1:0] node39035;
	wire [4-1:0] node39036;
	wire [4-1:0] node39039;
	wire [4-1:0] node39043;
	wire [4-1:0] node39044;
	wire [4-1:0] node39045;
	wire [4-1:0] node39046;
	wire [4-1:0] node39047;
	wire [4-1:0] node39049;
	wire [4-1:0] node39053;
	wire [4-1:0] node39054;
	wire [4-1:0] node39055;
	wire [4-1:0] node39059;
	wire [4-1:0] node39060;
	wire [4-1:0] node39064;
	wire [4-1:0] node39065;
	wire [4-1:0] node39066;
	wire [4-1:0] node39067;
	wire [4-1:0] node39070;
	wire [4-1:0] node39074;
	wire [4-1:0] node39075;
	wire [4-1:0] node39076;
	wire [4-1:0] node39079;
	wire [4-1:0] node39082;
	wire [4-1:0] node39084;
	wire [4-1:0] node39087;
	wire [4-1:0] node39088;
	wire [4-1:0] node39089;
	wire [4-1:0] node39090;
	wire [4-1:0] node39091;
	wire [4-1:0] node39094;
	wire [4-1:0] node39097;
	wire [4-1:0] node39098;
	wire [4-1:0] node39101;
	wire [4-1:0] node39104;
	wire [4-1:0] node39106;
	wire [4-1:0] node39107;
	wire [4-1:0] node39111;
	wire [4-1:0] node39112;
	wire [4-1:0] node39113;
	wire [4-1:0] node39114;
	wire [4-1:0] node39117;
	wire [4-1:0] node39120;
	wire [4-1:0] node39121;
	wire [4-1:0] node39124;
	wire [4-1:0] node39127;
	wire [4-1:0] node39129;
	wire [4-1:0] node39130;
	wire [4-1:0] node39133;
	wire [4-1:0] node39136;
	wire [4-1:0] node39137;
	wire [4-1:0] node39138;
	wire [4-1:0] node39139;
	wire [4-1:0] node39140;
	wire [4-1:0] node39142;
	wire [4-1:0] node39144;
	wire [4-1:0] node39147;
	wire [4-1:0] node39148;
	wire [4-1:0] node39149;
	wire [4-1:0] node39152;
	wire [4-1:0] node39155;
	wire [4-1:0] node39157;
	wire [4-1:0] node39160;
	wire [4-1:0] node39161;
	wire [4-1:0] node39163;
	wire [4-1:0] node39165;
	wire [4-1:0] node39168;
	wire [4-1:0] node39169;
	wire [4-1:0] node39170;
	wire [4-1:0] node39175;
	wire [4-1:0] node39176;
	wire [4-1:0] node39177;
	wire [4-1:0] node39178;
	wire [4-1:0] node39180;
	wire [4-1:0] node39184;
	wire [4-1:0] node39185;
	wire [4-1:0] node39189;
	wire [4-1:0] node39190;
	wire [4-1:0] node39192;
	wire [4-1:0] node39193;
	wire [4-1:0] node39197;
	wire [4-1:0] node39198;
	wire [4-1:0] node39199;
	wire [4-1:0] node39202;
	wire [4-1:0] node39206;
	wire [4-1:0] node39207;
	wire [4-1:0] node39208;
	wire [4-1:0] node39209;
	wire [4-1:0] node39210;
	wire [4-1:0] node39214;
	wire [4-1:0] node39216;
	wire [4-1:0] node39219;
	wire [4-1:0] node39221;
	wire [4-1:0] node39222;
	wire [4-1:0] node39223;
	wire [4-1:0] node39226;
	wire [4-1:0] node39229;
	wire [4-1:0] node39230;
	wire [4-1:0] node39233;
	wire [4-1:0] node39236;
	wire [4-1:0] node39237;
	wire [4-1:0] node39238;
	wire [4-1:0] node39239;
	wire [4-1:0] node39240;
	wire [4-1:0] node39243;
	wire [4-1:0] node39246;
	wire [4-1:0] node39248;
	wire [4-1:0] node39251;
	wire [4-1:0] node39253;
	wire [4-1:0] node39256;
	wire [4-1:0] node39257;
	wire [4-1:0] node39258;
	wire [4-1:0] node39259;
	wire [4-1:0] node39263;
	wire [4-1:0] node39265;
	wire [4-1:0] node39268;
	wire [4-1:0] node39269;
	wire [4-1:0] node39270;
	wire [4-1:0] node39274;
	wire [4-1:0] node39276;
	wire [4-1:0] node39279;
	wire [4-1:0] node39280;
	wire [4-1:0] node39281;
	wire [4-1:0] node39282;
	wire [4-1:0] node39283;
	wire [4-1:0] node39284;
	wire [4-1:0] node39285;
	wire [4-1:0] node39287;
	wire [4-1:0] node39290;
	wire [4-1:0] node39291;
	wire [4-1:0] node39295;
	wire [4-1:0] node39296;
	wire [4-1:0] node39298;
	wire [4-1:0] node39301;
	wire [4-1:0] node39302;
	wire [4-1:0] node39306;
	wire [4-1:0] node39307;
	wire [4-1:0] node39308;
	wire [4-1:0] node39309;
	wire [4-1:0] node39312;
	wire [4-1:0] node39316;
	wire [4-1:0] node39317;
	wire [4-1:0] node39318;
	wire [4-1:0] node39323;
	wire [4-1:0] node39324;
	wire [4-1:0] node39325;
	wire [4-1:0] node39326;
	wire [4-1:0] node39328;
	wire [4-1:0] node39331;
	wire [4-1:0] node39332;
	wire [4-1:0] node39336;
	wire [4-1:0] node39337;
	wire [4-1:0] node39339;
	wire [4-1:0] node39343;
	wire [4-1:0] node39344;
	wire [4-1:0] node39345;
	wire [4-1:0] node39347;
	wire [4-1:0] node39350;
	wire [4-1:0] node39352;
	wire [4-1:0] node39355;
	wire [4-1:0] node39356;
	wire [4-1:0] node39357;
	wire [4-1:0] node39362;
	wire [4-1:0] node39363;
	wire [4-1:0] node39364;
	wire [4-1:0] node39365;
	wire [4-1:0] node39366;
	wire [4-1:0] node39369;
	wire [4-1:0] node39370;
	wire [4-1:0] node39373;
	wire [4-1:0] node39376;
	wire [4-1:0] node39377;
	wire [4-1:0] node39378;
	wire [4-1:0] node39382;
	wire [4-1:0] node39384;
	wire [4-1:0] node39387;
	wire [4-1:0] node39388;
	wire [4-1:0] node39389;
	wire [4-1:0] node39390;
	wire [4-1:0] node39394;
	wire [4-1:0] node39397;
	wire [4-1:0] node39398;
	wire [4-1:0] node39399;
	wire [4-1:0] node39402;
	wire [4-1:0] node39406;
	wire [4-1:0] node39407;
	wire [4-1:0] node39408;
	wire [4-1:0] node39409;
	wire [4-1:0] node39410;
	wire [4-1:0] node39415;
	wire [4-1:0] node39416;
	wire [4-1:0] node39417;
	wire [4-1:0] node39420;
	wire [4-1:0] node39423;
	wire [4-1:0] node39425;
	wire [4-1:0] node39428;
	wire [4-1:0] node39429;
	wire [4-1:0] node39430;
	wire [4-1:0] node39432;
	wire [4-1:0] node39435;
	wire [4-1:0] node39436;
	wire [4-1:0] node39439;
	wire [4-1:0] node39442;
	wire [4-1:0] node39444;
	wire [4-1:0] node39447;
	wire [4-1:0] node39448;
	wire [4-1:0] node39449;
	wire [4-1:0] node39450;
	wire [4-1:0] node39451;
	wire [4-1:0] node39453;
	wire [4-1:0] node39454;
	wire [4-1:0] node39458;
	wire [4-1:0] node39459;
	wire [4-1:0] node39460;
	wire [4-1:0] node39464;
	wire [4-1:0] node39465;
	wire [4-1:0] node39469;
	wire [4-1:0] node39470;
	wire [4-1:0] node39471;
	wire [4-1:0] node39472;
	wire [4-1:0] node39475;
	wire [4-1:0] node39479;
	wire [4-1:0] node39480;
	wire [4-1:0] node39481;
	wire [4-1:0] node39486;
	wire [4-1:0] node39487;
	wire [4-1:0] node39488;
	wire [4-1:0] node39490;
	wire [4-1:0] node39492;
	wire [4-1:0] node39495;
	wire [4-1:0] node39496;
	wire [4-1:0] node39497;
	wire [4-1:0] node39501;
	wire [4-1:0] node39502;
	wire [4-1:0] node39506;
	wire [4-1:0] node39507;
	wire [4-1:0] node39508;
	wire [4-1:0] node39510;
	wire [4-1:0] node39513;
	wire [4-1:0] node39514;
	wire [4-1:0] node39517;
	wire [4-1:0] node39520;
	wire [4-1:0] node39523;
	wire [4-1:0] node39524;
	wire [4-1:0] node39525;
	wire [4-1:0] node39526;
	wire [4-1:0] node39527;
	wire [4-1:0] node39528;
	wire [4-1:0] node39531;
	wire [4-1:0] node39535;
	wire [4-1:0] node39536;
	wire [4-1:0] node39537;
	wire [4-1:0] node39542;
	wire [4-1:0] node39543;
	wire [4-1:0] node39546;
	wire [4-1:0] node39547;
	wire [4-1:0] node39548;
	wire [4-1:0] node39552;
	wire [4-1:0] node39553;
	wire [4-1:0] node39556;
	wire [4-1:0] node39559;
	wire [4-1:0] node39560;
	wire [4-1:0] node39561;
	wire [4-1:0] node39563;
	wire [4-1:0] node39564;
	wire [4-1:0] node39568;
	wire [4-1:0] node39569;
	wire [4-1:0] node39573;
	wire [4-1:0] node39574;
	wire [4-1:0] node39575;
	wire [4-1:0] node39576;
	wire [4-1:0] node39579;
	wire [4-1:0] node39583;
	wire [4-1:0] node39584;
	wire [4-1:0] node39585;
	wire [4-1:0] node39588;
	wire [4-1:0] node39591;
	wire [4-1:0] node39593;
	wire [4-1:0] node39596;
	wire [4-1:0] node39597;
	wire [4-1:0] node39598;
	wire [4-1:0] node39599;
	wire [4-1:0] node39600;
	wire [4-1:0] node39601;
	wire [4-1:0] node39602;
	wire [4-1:0] node39603;
	wire [4-1:0] node39607;
	wire [4-1:0] node39608;
	wire [4-1:0] node39609;
	wire [4-1:0] node39612;
	wire [4-1:0] node39615;
	wire [4-1:0] node39616;
	wire [4-1:0] node39620;
	wire [4-1:0] node39621;
	wire [4-1:0] node39622;
	wire [4-1:0] node39626;
	wire [4-1:0] node39628;
	wire [4-1:0] node39631;
	wire [4-1:0] node39632;
	wire [4-1:0] node39633;
	wire [4-1:0] node39634;
	wire [4-1:0] node39638;
	wire [4-1:0] node39639;
	wire [4-1:0] node39643;
	wire [4-1:0] node39644;
	wire [4-1:0] node39645;
	wire [4-1:0] node39648;
	wire [4-1:0] node39651;
	wire [4-1:0] node39653;
	wire [4-1:0] node39656;
	wire [4-1:0] node39657;
	wire [4-1:0] node39658;
	wire [4-1:0] node39659;
	wire [4-1:0] node39660;
	wire [4-1:0] node39662;
	wire [4-1:0] node39666;
	wire [4-1:0] node39667;
	wire [4-1:0] node39668;
	wire [4-1:0] node39671;
	wire [4-1:0] node39674;
	wire [4-1:0] node39675;
	wire [4-1:0] node39679;
	wire [4-1:0] node39680;
	wire [4-1:0] node39681;
	wire [4-1:0] node39682;
	wire [4-1:0] node39685;
	wire [4-1:0] node39688;
	wire [4-1:0] node39690;
	wire [4-1:0] node39693;
	wire [4-1:0] node39694;
	wire [4-1:0] node39695;
	wire [4-1:0] node39699;
	wire [4-1:0] node39700;
	wire [4-1:0] node39703;
	wire [4-1:0] node39706;
	wire [4-1:0] node39707;
	wire [4-1:0] node39708;
	wire [4-1:0] node39709;
	wire [4-1:0] node39711;
	wire [4-1:0] node39715;
	wire [4-1:0] node39717;
	wire [4-1:0] node39719;
	wire [4-1:0] node39722;
	wire [4-1:0] node39723;
	wire [4-1:0] node39724;
	wire [4-1:0] node39725;
	wire [4-1:0] node39728;
	wire [4-1:0] node39731;
	wire [4-1:0] node39733;
	wire [4-1:0] node39736;
	wire [4-1:0] node39737;
	wire [4-1:0] node39738;
	wire [4-1:0] node39742;
	wire [4-1:0] node39743;
	wire [4-1:0] node39746;
	wire [4-1:0] node39749;
	wire [4-1:0] node39750;
	wire [4-1:0] node39751;
	wire [4-1:0] node39752;
	wire [4-1:0] node39754;
	wire [4-1:0] node39755;
	wire [4-1:0] node39758;
	wire [4-1:0] node39761;
	wire [4-1:0] node39762;
	wire [4-1:0] node39763;
	wire [4-1:0] node39767;
	wire [4-1:0] node39769;
	wire [4-1:0] node39772;
	wire [4-1:0] node39773;
	wire [4-1:0] node39774;
	wire [4-1:0] node39775;
	wire [4-1:0] node39777;
	wire [4-1:0] node39781;
	wire [4-1:0] node39782;
	wire [4-1:0] node39783;
	wire [4-1:0] node39788;
	wire [4-1:0] node39789;
	wire [4-1:0] node39790;
	wire [4-1:0] node39793;
	wire [4-1:0] node39796;
	wire [4-1:0] node39797;
	wire [4-1:0] node39798;
	wire [4-1:0] node39801;
	wire [4-1:0] node39805;
	wire [4-1:0] node39806;
	wire [4-1:0] node39807;
	wire [4-1:0] node39808;
	wire [4-1:0] node39811;
	wire [4-1:0] node39813;
	wire [4-1:0] node39815;
	wire [4-1:0] node39818;
	wire [4-1:0] node39819;
	wire [4-1:0] node39820;
	wire [4-1:0] node39821;
	wire [4-1:0] node39825;
	wire [4-1:0] node39827;
	wire [4-1:0] node39830;
	wire [4-1:0] node39831;
	wire [4-1:0] node39832;
	wire [4-1:0] node39836;
	wire [4-1:0] node39838;
	wire [4-1:0] node39841;
	wire [4-1:0] node39842;
	wire [4-1:0] node39843;
	wire [4-1:0] node39844;
	wire [4-1:0] node39846;
	wire [4-1:0] node39849;
	wire [4-1:0] node39851;
	wire [4-1:0] node39854;
	wire [4-1:0] node39855;
	wire [4-1:0] node39857;
	wire [4-1:0] node39860;
	wire [4-1:0] node39861;
	wire [4-1:0] node39865;
	wire [4-1:0] node39866;
	wire [4-1:0] node39868;
	wire [4-1:0] node39869;
	wire [4-1:0] node39872;
	wire [4-1:0] node39875;
	wire [4-1:0] node39878;
	wire [4-1:0] node39879;
	wire [4-1:0] node39880;
	wire [4-1:0] node39881;
	wire [4-1:0] node39882;
	wire [4-1:0] node39883;
	wire [4-1:0] node39885;
	wire [4-1:0] node39886;
	wire [4-1:0] node39889;
	wire [4-1:0] node39892;
	wire [4-1:0] node39893;
	wire [4-1:0] node39894;
	wire [4-1:0] node39898;
	wire [4-1:0] node39900;
	wire [4-1:0] node39903;
	wire [4-1:0] node39904;
	wire [4-1:0] node39905;
	wire [4-1:0] node39909;
	wire [4-1:0] node39911;
	wire [4-1:0] node39914;
	wire [4-1:0] node39915;
	wire [4-1:0] node39916;
	wire [4-1:0] node39919;
	wire [4-1:0] node39920;
	wire [4-1:0] node39921;
	wire [4-1:0] node39924;
	wire [4-1:0] node39927;
	wire [4-1:0] node39929;
	wire [4-1:0] node39932;
	wire [4-1:0] node39933;
	wire [4-1:0] node39934;
	wire [4-1:0] node39937;
	wire [4-1:0] node39940;
	wire [4-1:0] node39941;
	wire [4-1:0] node39944;
	wire [4-1:0] node39947;
	wire [4-1:0] node39948;
	wire [4-1:0] node39949;
	wire [4-1:0] node39950;
	wire [4-1:0] node39952;
	wire [4-1:0] node39953;
	wire [4-1:0] node39956;
	wire [4-1:0] node39959;
	wire [4-1:0] node39960;
	wire [4-1:0] node39962;
	wire [4-1:0] node39966;
	wire [4-1:0] node39967;
	wire [4-1:0] node39968;
	wire [4-1:0] node39969;
	wire [4-1:0] node39972;
	wire [4-1:0] node39976;
	wire [4-1:0] node39977;
	wire [4-1:0] node39978;
	wire [4-1:0] node39982;
	wire [4-1:0] node39983;
	wire [4-1:0] node39987;
	wire [4-1:0] node39988;
	wire [4-1:0] node39989;
	wire [4-1:0] node39991;
	wire [4-1:0] node39994;
	wire [4-1:0] node39995;
	wire [4-1:0] node39998;
	wire [4-1:0] node40001;
	wire [4-1:0] node40002;
	wire [4-1:0] node40005;
	wire [4-1:0] node40006;
	wire [4-1:0] node40009;
	wire [4-1:0] node40012;
	wire [4-1:0] node40013;
	wire [4-1:0] node40014;
	wire [4-1:0] node40015;
	wire [4-1:0] node40016;
	wire [4-1:0] node40017;
	wire [4-1:0] node40020;
	wire [4-1:0] node40023;
	wire [4-1:0] node40024;
	wire [4-1:0] node40027;
	wire [4-1:0] node40030;
	wire [4-1:0] node40031;
	wire [4-1:0] node40032;
	wire [4-1:0] node40033;
	wire [4-1:0] node40037;
	wire [4-1:0] node40038;
	wire [4-1:0] node40041;
	wire [4-1:0] node40045;
	wire [4-1:0] node40046;
	wire [4-1:0] node40047;
	wire [4-1:0] node40048;
	wire [4-1:0] node40049;
	wire [4-1:0] node40053;
	wire [4-1:0] node40054;
	wire [4-1:0] node40058;
	wire [4-1:0] node40060;
	wire [4-1:0] node40063;
	wire [4-1:0] node40064;
	wire [4-1:0] node40065;
	wire [4-1:0] node40068;
	wire [4-1:0] node40071;
	wire [4-1:0] node40074;
	wire [4-1:0] node40075;
	wire [4-1:0] node40076;
	wire [4-1:0] node40077;
	wire [4-1:0] node40079;
	wire [4-1:0] node40080;
	wire [4-1:0] node40083;
	wire [4-1:0] node40086;
	wire [4-1:0] node40088;
	wire [4-1:0] node40091;
	wire [4-1:0] node40093;
	wire [4-1:0] node40094;
	wire [4-1:0] node40097;
	wire [4-1:0] node40100;
	wire [4-1:0] node40101;
	wire [4-1:0] node40102;
	wire [4-1:0] node40104;
	wire [4-1:0] node40107;
	wire [4-1:0] node40108;
	wire [4-1:0] node40109;
	wire [4-1:0] node40113;
	wire [4-1:0] node40114;
	wire [4-1:0] node40117;
	wire [4-1:0] node40120;
	wire [4-1:0] node40121;
	wire [4-1:0] node40122;
	wire [4-1:0] node40126;
	wire [4-1:0] node40127;
	wire [4-1:0] node40128;
	wire [4-1:0] node40131;
	wire [4-1:0] node40135;
	wire [4-1:0] node40136;
	wire [4-1:0] node40137;
	wire [4-1:0] node40138;
	wire [4-1:0] node40139;
	wire [4-1:0] node40140;
	wire [4-1:0] node40141;
	wire [4-1:0] node40142;
	wire [4-1:0] node40143;
	wire [4-1:0] node40144;
	wire [4-1:0] node40145;
	wire [4-1:0] node40148;
	wire [4-1:0] node40149;
	wire [4-1:0] node40150;
	wire [4-1:0] node40155;
	wire [4-1:0] node40156;
	wire [4-1:0] node40157;
	wire [4-1:0] node40158;
	wire [4-1:0] node40161;
	wire [4-1:0] node40165;
	wire [4-1:0] node40166;
	wire [4-1:0] node40168;
	wire [4-1:0] node40171;
	wire [4-1:0] node40172;
	wire [4-1:0] node40175;
	wire [4-1:0] node40178;
	wire [4-1:0] node40179;
	wire [4-1:0] node40180;
	wire [4-1:0] node40181;
	wire [4-1:0] node40182;
	wire [4-1:0] node40186;
	wire [4-1:0] node40187;
	wire [4-1:0] node40190;
	wire [4-1:0] node40193;
	wire [4-1:0] node40195;
	wire [4-1:0] node40196;
	wire [4-1:0] node40200;
	wire [4-1:0] node40201;
	wire [4-1:0] node40202;
	wire [4-1:0] node40203;
	wire [4-1:0] node40206;
	wire [4-1:0] node40209;
	wire [4-1:0] node40212;
	wire [4-1:0] node40213;
	wire [4-1:0] node40214;
	wire [4-1:0] node40217;
	wire [4-1:0] node40220;
	wire [4-1:0] node40223;
	wire [4-1:0] node40224;
	wire [4-1:0] node40225;
	wire [4-1:0] node40226;
	wire [4-1:0] node40227;
	wire [4-1:0] node40229;
	wire [4-1:0] node40232;
	wire [4-1:0] node40233;
	wire [4-1:0] node40236;
	wire [4-1:0] node40239;
	wire [4-1:0] node40240;
	wire [4-1:0] node40242;
	wire [4-1:0] node40245;
	wire [4-1:0] node40248;
	wire [4-1:0] node40249;
	wire [4-1:0] node40250;
	wire [4-1:0] node40251;
	wire [4-1:0] node40254;
	wire [4-1:0] node40257;
	wire [4-1:0] node40260;
	wire [4-1:0] node40261;
	wire [4-1:0] node40265;
	wire [4-1:0] node40266;
	wire [4-1:0] node40267;
	wire [4-1:0] node40268;
	wire [4-1:0] node40269;
	wire [4-1:0] node40273;
	wire [4-1:0] node40275;
	wire [4-1:0] node40278;
	wire [4-1:0] node40280;
	wire [4-1:0] node40281;
	wire [4-1:0] node40284;
	wire [4-1:0] node40287;
	wire [4-1:0] node40288;
	wire [4-1:0] node40289;
	wire [4-1:0] node40290;
	wire [4-1:0] node40295;
	wire [4-1:0] node40296;
	wire [4-1:0] node40297;
	wire [4-1:0] node40301;
	wire [4-1:0] node40302;
	wire [4-1:0] node40306;
	wire [4-1:0] node40307;
	wire [4-1:0] node40308;
	wire [4-1:0] node40309;
	wire [4-1:0] node40310;
	wire [4-1:0] node40311;
	wire [4-1:0] node40313;
	wire [4-1:0] node40316;
	wire [4-1:0] node40319;
	wire [4-1:0] node40320;
	wire [4-1:0] node40321;
	wire [4-1:0] node40326;
	wire [4-1:0] node40327;
	wire [4-1:0] node40328;
	wire [4-1:0] node40329;
	wire [4-1:0] node40333;
	wire [4-1:0] node40334;
	wire [4-1:0] node40338;
	wire [4-1:0] node40340;
	wire [4-1:0] node40341;
	wire [4-1:0] node40345;
	wire [4-1:0] node40346;
	wire [4-1:0] node40347;
	wire [4-1:0] node40348;
	wire [4-1:0] node40350;
	wire [4-1:0] node40354;
	wire [4-1:0] node40355;
	wire [4-1:0] node40358;
	wire [4-1:0] node40359;
	wire [4-1:0] node40363;
	wire [4-1:0] node40364;
	wire [4-1:0] node40365;
	wire [4-1:0] node40368;
	wire [4-1:0] node40369;
	wire [4-1:0] node40372;
	wire [4-1:0] node40375;
	wire [4-1:0] node40377;
	wire [4-1:0] node40378;
	wire [4-1:0] node40381;
	wire [4-1:0] node40384;
	wire [4-1:0] node40385;
	wire [4-1:0] node40386;
	wire [4-1:0] node40387;
	wire [4-1:0] node40388;
	wire [4-1:0] node40391;
	wire [4-1:0] node40392;
	wire [4-1:0] node40396;
	wire [4-1:0] node40398;
	wire [4-1:0] node40400;
	wire [4-1:0] node40403;
	wire [4-1:0] node40404;
	wire [4-1:0] node40405;
	wire [4-1:0] node40406;
	wire [4-1:0] node40409;
	wire [4-1:0] node40413;
	wire [4-1:0] node40416;
	wire [4-1:0] node40417;
	wire [4-1:0] node40418;
	wire [4-1:0] node40419;
	wire [4-1:0] node40420;
	wire [4-1:0] node40424;
	wire [4-1:0] node40425;
	wire [4-1:0] node40428;
	wire [4-1:0] node40431;
	wire [4-1:0] node40432;
	wire [4-1:0] node40435;
	wire [4-1:0] node40436;
	wire [4-1:0] node40439;
	wire [4-1:0] node40442;
	wire [4-1:0] node40443;
	wire [4-1:0] node40444;
	wire [4-1:0] node40445;
	wire [4-1:0] node40449;
	wire [4-1:0] node40451;
	wire [4-1:0] node40454;
	wire [4-1:0] node40457;
	wire [4-1:0] node40458;
	wire [4-1:0] node40459;
	wire [4-1:0] node40460;
	wire [4-1:0] node40461;
	wire [4-1:0] node40462;
	wire [4-1:0] node40463;
	wire [4-1:0] node40466;
	wire [4-1:0] node40469;
	wire [4-1:0] node40470;
	wire [4-1:0] node40471;
	wire [4-1:0] node40475;
	wire [4-1:0] node40477;
	wire [4-1:0] node40480;
	wire [4-1:0] node40481;
	wire [4-1:0] node40482;
	wire [4-1:0] node40485;
	wire [4-1:0] node40486;
	wire [4-1:0] node40489;
	wire [4-1:0] node40492;
	wire [4-1:0] node40494;
	wire [4-1:0] node40495;
	wire [4-1:0] node40499;
	wire [4-1:0] node40500;
	wire [4-1:0] node40501;
	wire [4-1:0] node40502;
	wire [4-1:0] node40503;
	wire [4-1:0] node40506;
	wire [4-1:0] node40510;
	wire [4-1:0] node40512;
	wire [4-1:0] node40513;
	wire [4-1:0] node40516;
	wire [4-1:0] node40519;
	wire [4-1:0] node40520;
	wire [4-1:0] node40522;
	wire [4-1:0] node40523;
	wire [4-1:0] node40526;
	wire [4-1:0] node40529;
	wire [4-1:0] node40530;
	wire [4-1:0] node40531;
	wire [4-1:0] node40534;
	wire [4-1:0] node40538;
	wire [4-1:0] node40539;
	wire [4-1:0] node40540;
	wire [4-1:0] node40541;
	wire [4-1:0] node40542;
	wire [4-1:0] node40543;
	wire [4-1:0] node40546;
	wire [4-1:0] node40550;
	wire [4-1:0] node40552;
	wire [4-1:0] node40554;
	wire [4-1:0] node40557;
	wire [4-1:0] node40558;
	wire [4-1:0] node40559;
	wire [4-1:0] node40560;
	wire [4-1:0] node40564;
	wire [4-1:0] node40566;
	wire [4-1:0] node40569;
	wire [4-1:0] node40570;
	wire [4-1:0] node40572;
	wire [4-1:0] node40575;
	wire [4-1:0] node40577;
	wire [4-1:0] node40580;
	wire [4-1:0] node40581;
	wire [4-1:0] node40582;
	wire [4-1:0] node40583;
	wire [4-1:0] node40585;
	wire [4-1:0] node40588;
	wire [4-1:0] node40590;
	wire [4-1:0] node40593;
	wire [4-1:0] node40594;
	wire [4-1:0] node40597;
	wire [4-1:0] node40600;
	wire [4-1:0] node40601;
	wire [4-1:0] node40602;
	wire [4-1:0] node40603;
	wire [4-1:0] node40608;
	wire [4-1:0] node40609;
	wire [4-1:0] node40611;
	wire [4-1:0] node40614;
	wire [4-1:0] node40615;
	wire [4-1:0] node40618;
	wire [4-1:0] node40621;
	wire [4-1:0] node40622;
	wire [4-1:0] node40623;
	wire [4-1:0] node40624;
	wire [4-1:0] node40625;
	wire [4-1:0] node40626;
	wire [4-1:0] node40627;
	wire [4-1:0] node40631;
	wire [4-1:0] node40632;
	wire [4-1:0] node40636;
	wire [4-1:0] node40637;
	wire [4-1:0] node40638;
	wire [4-1:0] node40641;
	wire [4-1:0] node40644;
	wire [4-1:0] node40645;
	wire [4-1:0] node40649;
	wire [4-1:0] node40650;
	wire [4-1:0] node40651;
	wire [4-1:0] node40654;
	wire [4-1:0] node40656;
	wire [4-1:0] node40659;
	wire [4-1:0] node40660;
	wire [4-1:0] node40661;
	wire [4-1:0] node40666;
	wire [4-1:0] node40667;
	wire [4-1:0] node40668;
	wire [4-1:0] node40670;
	wire [4-1:0] node40673;
	wire [4-1:0] node40674;
	wire [4-1:0] node40675;
	wire [4-1:0] node40680;
	wire [4-1:0] node40681;
	wire [4-1:0] node40682;
	wire [4-1:0] node40683;
	wire [4-1:0] node40687;
	wire [4-1:0] node40688;
	wire [4-1:0] node40691;
	wire [4-1:0] node40694;
	wire [4-1:0] node40695;
	wire [4-1:0] node40697;
	wire [4-1:0] node40701;
	wire [4-1:0] node40702;
	wire [4-1:0] node40703;
	wire [4-1:0] node40704;
	wire [4-1:0] node40705;
	wire [4-1:0] node40707;
	wire [4-1:0] node40710;
	wire [4-1:0] node40713;
	wire [4-1:0] node40714;
	wire [4-1:0] node40715;
	wire [4-1:0] node40719;
	wire [4-1:0] node40720;
	wire [4-1:0] node40723;
	wire [4-1:0] node40726;
	wire [4-1:0] node40727;
	wire [4-1:0] node40728;
	wire [4-1:0] node40731;
	wire [4-1:0] node40732;
	wire [4-1:0] node40736;
	wire [4-1:0] node40737;
	wire [4-1:0] node40738;
	wire [4-1:0] node40743;
	wire [4-1:0] node40744;
	wire [4-1:0] node40745;
	wire [4-1:0] node40746;
	wire [4-1:0] node40748;
	wire [4-1:0] node40752;
	wire [4-1:0] node40754;
	wire [4-1:0] node40756;
	wire [4-1:0] node40759;
	wire [4-1:0] node40760;
	wire [4-1:0] node40761;
	wire [4-1:0] node40762;
	wire [4-1:0] node40765;
	wire [4-1:0] node40768;
	wire [4-1:0] node40770;
	wire [4-1:0] node40773;
	wire [4-1:0] node40774;
	wire [4-1:0] node40775;
	wire [4-1:0] node40778;
	wire [4-1:0] node40782;
	wire [4-1:0] node40783;
	wire [4-1:0] node40784;
	wire [4-1:0] node40785;
	wire [4-1:0] node40786;
	wire [4-1:0] node40787;
	wire [4-1:0] node40788;
	wire [4-1:0] node40790;
	wire [4-1:0] node40793;
	wire [4-1:0] node40794;
	wire [4-1:0] node40795;
	wire [4-1:0] node40798;
	wire [4-1:0] node40801;
	wire [4-1:0] node40802;
	wire [4-1:0] node40806;
	wire [4-1:0] node40807;
	wire [4-1:0] node40808;
	wire [4-1:0] node40809;
	wire [4-1:0] node40812;
	wire [4-1:0] node40816;
	wire [4-1:0] node40817;
	wire [4-1:0] node40818;
	wire [4-1:0] node40821;
	wire [4-1:0] node40825;
	wire [4-1:0] node40826;
	wire [4-1:0] node40827;
	wire [4-1:0] node40829;
	wire [4-1:0] node40831;
	wire [4-1:0] node40834;
	wire [4-1:0] node40835;
	wire [4-1:0] node40837;
	wire [4-1:0] node40840;
	wire [4-1:0] node40842;
	wire [4-1:0] node40845;
	wire [4-1:0] node40846;
	wire [4-1:0] node40847;
	wire [4-1:0] node40848;
	wire [4-1:0] node40851;
	wire [4-1:0] node40854;
	wire [4-1:0] node40856;
	wire [4-1:0] node40859;
	wire [4-1:0] node40860;
	wire [4-1:0] node40861;
	wire [4-1:0] node40864;
	wire [4-1:0] node40868;
	wire [4-1:0] node40869;
	wire [4-1:0] node40870;
	wire [4-1:0] node40871;
	wire [4-1:0] node40872;
	wire [4-1:0] node40873;
	wire [4-1:0] node40876;
	wire [4-1:0] node40879;
	wire [4-1:0] node40880;
	wire [4-1:0] node40884;
	wire [4-1:0] node40885;
	wire [4-1:0] node40886;
	wire [4-1:0] node40889;
	wire [4-1:0] node40892;
	wire [4-1:0] node40893;
	wire [4-1:0] node40896;
	wire [4-1:0] node40899;
	wire [4-1:0] node40900;
	wire [4-1:0] node40901;
	wire [4-1:0] node40902;
	wire [4-1:0] node40906;
	wire [4-1:0] node40907;
	wire [4-1:0] node40910;
	wire [4-1:0] node40913;
	wire [4-1:0] node40914;
	wire [4-1:0] node40915;
	wire [4-1:0] node40918;
	wire [4-1:0] node40921;
	wire [4-1:0] node40922;
	wire [4-1:0] node40926;
	wire [4-1:0] node40927;
	wire [4-1:0] node40928;
	wire [4-1:0] node40929;
	wire [4-1:0] node40930;
	wire [4-1:0] node40934;
	wire [4-1:0] node40935;
	wire [4-1:0] node40939;
	wire [4-1:0] node40940;
	wire [4-1:0] node40941;
	wire [4-1:0] node40945;
	wire [4-1:0] node40946;
	wire [4-1:0] node40950;
	wire [4-1:0] node40951;
	wire [4-1:0] node40952;
	wire [4-1:0] node40956;
	wire [4-1:0] node40957;
	wire [4-1:0] node40959;
	wire [4-1:0] node40963;
	wire [4-1:0] node40964;
	wire [4-1:0] node40965;
	wire [4-1:0] node40966;
	wire [4-1:0] node40967;
	wire [4-1:0] node40969;
	wire [4-1:0] node40970;
	wire [4-1:0] node40973;
	wire [4-1:0] node40976;
	wire [4-1:0] node40978;
	wire [4-1:0] node40979;
	wire [4-1:0] node40982;
	wire [4-1:0] node40985;
	wire [4-1:0] node40986;
	wire [4-1:0] node40987;
	wire [4-1:0] node40989;
	wire [4-1:0] node40992;
	wire [4-1:0] node40993;
	wire [4-1:0] node40996;
	wire [4-1:0] node41000;
	wire [4-1:0] node41001;
	wire [4-1:0] node41002;
	wire [4-1:0] node41004;
	wire [4-1:0] node41005;
	wire [4-1:0] node41008;
	wire [4-1:0] node41011;
	wire [4-1:0] node41012;
	wire [4-1:0] node41013;
	wire [4-1:0] node41016;
	wire [4-1:0] node41020;
	wire [4-1:0] node41021;
	wire [4-1:0] node41022;
	wire [4-1:0] node41023;
	wire [4-1:0] node41026;
	wire [4-1:0] node41029;
	wire [4-1:0] node41030;
	wire [4-1:0] node41034;
	wire [4-1:0] node41035;
	wire [4-1:0] node41039;
	wire [4-1:0] node41040;
	wire [4-1:0] node41041;
	wire [4-1:0] node41042;
	wire [4-1:0] node41043;
	wire [4-1:0] node41045;
	wire [4-1:0] node41049;
	wire [4-1:0] node41050;
	wire [4-1:0] node41051;
	wire [4-1:0] node41054;
	wire [4-1:0] node41057;
	wire [4-1:0] node41058;
	wire [4-1:0] node41062;
	wire [4-1:0] node41063;
	wire [4-1:0] node41066;
	wire [4-1:0] node41067;
	wire [4-1:0] node41071;
	wire [4-1:0] node41072;
	wire [4-1:0] node41073;
	wire [4-1:0] node41075;
	wire [4-1:0] node41078;
	wire [4-1:0] node41080;
	wire [4-1:0] node41083;
	wire [4-1:0] node41084;
	wire [4-1:0] node41085;
	wire [4-1:0] node41087;
	wire [4-1:0] node41090;
	wire [4-1:0] node41091;
	wire [4-1:0] node41095;
	wire [4-1:0] node41097;
	wire [4-1:0] node41100;
	wire [4-1:0] node41101;
	wire [4-1:0] node41102;
	wire [4-1:0] node41103;
	wire [4-1:0] node41104;
	wire [4-1:0] node41105;
	wire [4-1:0] node41106;
	wire [4-1:0] node41107;
	wire [4-1:0] node41110;
	wire [4-1:0] node41114;
	wire [4-1:0] node41116;
	wire [4-1:0] node41117;
	wire [4-1:0] node41120;
	wire [4-1:0] node41123;
	wire [4-1:0] node41124;
	wire [4-1:0] node41126;
	wire [4-1:0] node41127;
	wire [4-1:0] node41130;
	wire [4-1:0] node41133;
	wire [4-1:0] node41134;
	wire [4-1:0] node41135;
	wire [4-1:0] node41139;
	wire [4-1:0] node41141;
	wire [4-1:0] node41144;
	wire [4-1:0] node41145;
	wire [4-1:0] node41146;
	wire [4-1:0] node41148;
	wire [4-1:0] node41149;
	wire [4-1:0] node41153;
	wire [4-1:0] node41155;
	wire [4-1:0] node41157;
	wire [4-1:0] node41160;
	wire [4-1:0] node41161;
	wire [4-1:0] node41162;
	wire [4-1:0] node41163;
	wire [4-1:0] node41167;
	wire [4-1:0] node41168;
	wire [4-1:0] node41171;
	wire [4-1:0] node41175;
	wire [4-1:0] node41176;
	wire [4-1:0] node41177;
	wire [4-1:0] node41178;
	wire [4-1:0] node41180;
	wire [4-1:0] node41183;
	wire [4-1:0] node41184;
	wire [4-1:0] node41186;
	wire [4-1:0] node41189;
	wire [4-1:0] node41190;
	wire [4-1:0] node41193;
	wire [4-1:0] node41196;
	wire [4-1:0] node41197;
	wire [4-1:0] node41198;
	wire [4-1:0] node41200;
	wire [4-1:0] node41203;
	wire [4-1:0] node41204;
	wire [4-1:0] node41207;
	wire [4-1:0] node41210;
	wire [4-1:0] node41211;
	wire [4-1:0] node41212;
	wire [4-1:0] node41216;
	wire [4-1:0] node41217;
	wire [4-1:0] node41221;
	wire [4-1:0] node41222;
	wire [4-1:0] node41223;
	wire [4-1:0] node41225;
	wire [4-1:0] node41227;
	wire [4-1:0] node41230;
	wire [4-1:0] node41231;
	wire [4-1:0] node41232;
	wire [4-1:0] node41235;
	wire [4-1:0] node41238;
	wire [4-1:0] node41239;
	wire [4-1:0] node41243;
	wire [4-1:0] node41244;
	wire [4-1:0] node41245;
	wire [4-1:0] node41248;
	wire [4-1:0] node41249;
	wire [4-1:0] node41253;
	wire [4-1:0] node41254;
	wire [4-1:0] node41255;
	wire [4-1:0] node41260;
	wire [4-1:0] node41261;
	wire [4-1:0] node41262;
	wire [4-1:0] node41263;
	wire [4-1:0] node41264;
	wire [4-1:0] node41265;
	wire [4-1:0] node41266;
	wire [4-1:0] node41270;
	wire [4-1:0] node41271;
	wire [4-1:0] node41274;
	wire [4-1:0] node41277;
	wire [4-1:0] node41278;
	wire [4-1:0] node41279;
	wire [4-1:0] node41282;
	wire [4-1:0] node41286;
	wire [4-1:0] node41287;
	wire [4-1:0] node41290;
	wire [4-1:0] node41293;
	wire [4-1:0] node41294;
	wire [4-1:0] node41295;
	wire [4-1:0] node41297;
	wire [4-1:0] node41300;
	wire [4-1:0] node41301;
	wire [4-1:0] node41303;
	wire [4-1:0] node41307;
	wire [4-1:0] node41308;
	wire [4-1:0] node41309;
	wire [4-1:0] node41310;
	wire [4-1:0] node41313;
	wire [4-1:0] node41317;
	wire [4-1:0] node41318;
	wire [4-1:0] node41320;
	wire [4-1:0] node41323;
	wire [4-1:0] node41325;
	wire [4-1:0] node41328;
	wire [4-1:0] node41329;
	wire [4-1:0] node41330;
	wire [4-1:0] node41331;
	wire [4-1:0] node41332;
	wire [4-1:0] node41336;
	wire [4-1:0] node41337;
	wire [4-1:0] node41338;
	wire [4-1:0] node41341;
	wire [4-1:0] node41344;
	wire [4-1:0] node41346;
	wire [4-1:0] node41349;
	wire [4-1:0] node41350;
	wire [4-1:0] node41351;
	wire [4-1:0] node41352;
	wire [4-1:0] node41356;
	wire [4-1:0] node41357;
	wire [4-1:0] node41361;
	wire [4-1:0] node41362;
	wire [4-1:0] node41365;
	wire [4-1:0] node41368;
	wire [4-1:0] node41369;
	wire [4-1:0] node41370;
	wire [4-1:0] node41373;
	wire [4-1:0] node41374;
	wire [4-1:0] node41377;
	wire [4-1:0] node41378;
	wire [4-1:0] node41382;
	wire [4-1:0] node41383;
	wire [4-1:0] node41384;
	wire [4-1:0] node41385;
	wire [4-1:0] node41388;
	wire [4-1:0] node41391;
	wire [4-1:0] node41393;
	wire [4-1:0] node41396;
	wire [4-1:0] node41397;
	wire [4-1:0] node41398;
	wire [4-1:0] node41401;
	wire [4-1:0] node41405;
	wire [4-1:0] node41406;
	wire [4-1:0] node41407;
	wire [4-1:0] node41408;
	wire [4-1:0] node41409;
	wire [4-1:0] node41410;
	wire [4-1:0] node41411;
	wire [4-1:0] node41412;
	wire [4-1:0] node41415;
	wire [4-1:0] node41418;
	wire [4-1:0] node41419;
	wire [4-1:0] node41421;
	wire [4-1:0] node41424;
	wire [4-1:0] node41425;
	wire [4-1:0] node41428;
	wire [4-1:0] node41431;
	wire [4-1:0] node41432;
	wire [4-1:0] node41433;
	wire [4-1:0] node41434;
	wire [4-1:0] node41435;
	wire [4-1:0] node41438;
	wire [4-1:0] node41441;
	wire [4-1:0] node41442;
	wire [4-1:0] node41446;
	wire [4-1:0] node41448;
	wire [4-1:0] node41451;
	wire [4-1:0] node41452;
	wire [4-1:0] node41453;
	wire [4-1:0] node41457;
	wire [4-1:0] node41458;
	wire [4-1:0] node41461;
	wire [4-1:0] node41464;
	wire [4-1:0] node41465;
	wire [4-1:0] node41466;
	wire [4-1:0] node41467;
	wire [4-1:0] node41470;
	wire [4-1:0] node41473;
	wire [4-1:0] node41474;
	wire [4-1:0] node41475;
	wire [4-1:0] node41479;
	wire [4-1:0] node41480;
	wire [4-1:0] node41483;
	wire [4-1:0] node41486;
	wire [4-1:0] node41487;
	wire [4-1:0] node41488;
	wire [4-1:0] node41489;
	wire [4-1:0] node41491;
	wire [4-1:0] node41494;
	wire [4-1:0] node41495;
	wire [4-1:0] node41498;
	wire [4-1:0] node41501;
	wire [4-1:0] node41503;
	wire [4-1:0] node41506;
	wire [4-1:0] node41507;
	wire [4-1:0] node41508;
	wire [4-1:0] node41513;
	wire [4-1:0] node41514;
	wire [4-1:0] node41515;
	wire [4-1:0] node41516;
	wire [4-1:0] node41517;
	wire [4-1:0] node41521;
	wire [4-1:0] node41522;
	wire [4-1:0] node41523;
	wire [4-1:0] node41526;
	wire [4-1:0] node41529;
	wire [4-1:0] node41530;
	wire [4-1:0] node41533;
	wire [4-1:0] node41536;
	wire [4-1:0] node41537;
	wire [4-1:0] node41539;
	wire [4-1:0] node41541;
	wire [4-1:0] node41544;
	wire [4-1:0] node41545;
	wire [4-1:0] node41547;
	wire [4-1:0] node41550;
	wire [4-1:0] node41551;
	wire [4-1:0] node41554;
	wire [4-1:0] node41557;
	wire [4-1:0] node41558;
	wire [4-1:0] node41559;
	wire [4-1:0] node41560;
	wire [4-1:0] node41561;
	wire [4-1:0] node41564;
	wire [4-1:0] node41567;
	wire [4-1:0] node41569;
	wire [4-1:0] node41572;
	wire [4-1:0] node41573;
	wire [4-1:0] node41574;
	wire [4-1:0] node41577;
	wire [4-1:0] node41580;
	wire [4-1:0] node41581;
	wire [4-1:0] node41584;
	wire [4-1:0] node41587;
	wire [4-1:0] node41588;
	wire [4-1:0] node41589;
	wire [4-1:0] node41592;
	wire [4-1:0] node41595;
	wire [4-1:0] node41596;
	wire [4-1:0] node41598;
	wire [4-1:0] node41599;
	wire [4-1:0] node41602;
	wire [4-1:0] node41605;
	wire [4-1:0] node41607;
	wire [4-1:0] node41610;
	wire [4-1:0] node41611;
	wire [4-1:0] node41612;
	wire [4-1:0] node41613;
	wire [4-1:0] node41614;
	wire [4-1:0] node41615;
	wire [4-1:0] node41616;
	wire [4-1:0] node41620;
	wire [4-1:0] node41621;
	wire [4-1:0] node41622;
	wire [4-1:0] node41626;
	wire [4-1:0] node41627;
	wire [4-1:0] node41630;
	wire [4-1:0] node41633;
	wire [4-1:0] node41634;
	wire [4-1:0] node41635;
	wire [4-1:0] node41638;
	wire [4-1:0] node41641;
	wire [4-1:0] node41642;
	wire [4-1:0] node41643;
	wire [4-1:0] node41646;
	wire [4-1:0] node41650;
	wire [4-1:0] node41651;
	wire [4-1:0] node41652;
	wire [4-1:0] node41654;
	wire [4-1:0] node41657;
	wire [4-1:0] node41659;
	wire [4-1:0] node41662;
	wire [4-1:0] node41663;
	wire [4-1:0] node41665;
	wire [4-1:0] node41668;
	wire [4-1:0] node41669;
	wire [4-1:0] node41672;
	wire [4-1:0] node41675;
	wire [4-1:0] node41676;
	wire [4-1:0] node41677;
	wire [4-1:0] node41678;
	wire [4-1:0] node41679;
	wire [4-1:0] node41682;
	wire [4-1:0] node41685;
	wire [4-1:0] node41686;
	wire [4-1:0] node41687;
	wire [4-1:0] node41692;
	wire [4-1:0] node41693;
	wire [4-1:0] node41694;
	wire [4-1:0] node41697;
	wire [4-1:0] node41700;
	wire [4-1:0] node41701;
	wire [4-1:0] node41704;
	wire [4-1:0] node41707;
	wire [4-1:0] node41708;
	wire [4-1:0] node41709;
	wire [4-1:0] node41710;
	wire [4-1:0] node41711;
	wire [4-1:0] node41714;
	wire [4-1:0] node41718;
	wire [4-1:0] node41719;
	wire [4-1:0] node41721;
	wire [4-1:0] node41724;
	wire [4-1:0] node41725;
	wire [4-1:0] node41729;
	wire [4-1:0] node41730;
	wire [4-1:0] node41733;
	wire [4-1:0] node41735;
	wire [4-1:0] node41738;
	wire [4-1:0] node41739;
	wire [4-1:0] node41740;
	wire [4-1:0] node41741;
	wire [4-1:0] node41742;
	wire [4-1:0] node41744;
	wire [4-1:0] node41747;
	wire [4-1:0] node41749;
	wire [4-1:0] node41752;
	wire [4-1:0] node41753;
	wire [4-1:0] node41754;
	wire [4-1:0] node41755;
	wire [4-1:0] node41759;
	wire [4-1:0] node41762;
	wire [4-1:0] node41764;
	wire [4-1:0] node41766;
	wire [4-1:0] node41769;
	wire [4-1:0] node41770;
	wire [4-1:0] node41771;
	wire [4-1:0] node41772;
	wire [4-1:0] node41773;
	wire [4-1:0] node41776;
	wire [4-1:0] node41779;
	wire [4-1:0] node41780;
	wire [4-1:0] node41783;
	wire [4-1:0] node41786;
	wire [4-1:0] node41787;
	wire [4-1:0] node41788;
	wire [4-1:0] node41791;
	wire [4-1:0] node41795;
	wire [4-1:0] node41797;
	wire [4-1:0] node41798;
	wire [4-1:0] node41799;
	wire [4-1:0] node41804;
	wire [4-1:0] node41805;
	wire [4-1:0] node41806;
	wire [4-1:0] node41807;
	wire [4-1:0] node41808;
	wire [4-1:0] node41813;
	wire [4-1:0] node41814;
	wire [4-1:0] node41815;
	wire [4-1:0] node41818;
	wire [4-1:0] node41821;
	wire [4-1:0] node41823;
	wire [4-1:0] node41826;
	wire [4-1:0] node41827;
	wire [4-1:0] node41828;
	wire [4-1:0] node41829;
	wire [4-1:0] node41832;
	wire [4-1:0] node41835;
	wire [4-1:0] node41836;
	wire [4-1:0] node41840;
	wire [4-1:0] node41841;
	wire [4-1:0] node41842;
	wire [4-1:0] node41846;
	wire [4-1:0] node41848;
	wire [4-1:0] node41851;
	wire [4-1:0] node41852;
	wire [4-1:0] node41853;
	wire [4-1:0] node41854;
	wire [4-1:0] node41855;
	wire [4-1:0] node41856;
	wire [4-1:0] node41857;
	wire [4-1:0] node41858;
	wire [4-1:0] node41860;
	wire [4-1:0] node41864;
	wire [4-1:0] node41867;
	wire [4-1:0] node41868;
	wire [4-1:0] node41869;
	wire [4-1:0] node41871;
	wire [4-1:0] node41874;
	wire [4-1:0] node41875;
	wire [4-1:0] node41879;
	wire [4-1:0] node41880;
	wire [4-1:0] node41883;
	wire [4-1:0] node41886;
	wire [4-1:0] node41887;
	wire [4-1:0] node41888;
	wire [4-1:0] node41890;
	wire [4-1:0] node41891;
	wire [4-1:0] node41895;
	wire [4-1:0] node41896;
	wire [4-1:0] node41900;
	wire [4-1:0] node41901;
	wire [4-1:0] node41902;
	wire [4-1:0] node41903;
	wire [4-1:0] node41908;
	wire [4-1:0] node41909;
	wire [4-1:0] node41913;
	wire [4-1:0] node41914;
	wire [4-1:0] node41915;
	wire [4-1:0] node41916;
	wire [4-1:0] node41917;
	wire [4-1:0] node41918;
	wire [4-1:0] node41922;
	wire [4-1:0] node41923;
	wire [4-1:0] node41927;
	wire [4-1:0] node41928;
	wire [4-1:0] node41929;
	wire [4-1:0] node41932;
	wire [4-1:0] node41935;
	wire [4-1:0] node41936;
	wire [4-1:0] node41939;
	wire [4-1:0] node41942;
	wire [4-1:0] node41943;
	wire [4-1:0] node41945;
	wire [4-1:0] node41946;
	wire [4-1:0] node41950;
	wire [4-1:0] node41951;
	wire [4-1:0] node41955;
	wire [4-1:0] node41956;
	wire [4-1:0] node41957;
	wire [4-1:0] node41959;
	wire [4-1:0] node41961;
	wire [4-1:0] node41964;
	wire [4-1:0] node41965;
	wire [4-1:0] node41966;
	wire [4-1:0] node41969;
	wire [4-1:0] node41972;
	wire [4-1:0] node41973;
	wire [4-1:0] node41977;
	wire [4-1:0] node41978;
	wire [4-1:0] node41979;
	wire [4-1:0] node41980;
	wire [4-1:0] node41983;
	wire [4-1:0] node41986;
	wire [4-1:0] node41988;
	wire [4-1:0] node41991;
	wire [4-1:0] node41992;
	wire [4-1:0] node41994;
	wire [4-1:0] node41997;
	wire [4-1:0] node42000;
	wire [4-1:0] node42001;
	wire [4-1:0] node42002;
	wire [4-1:0] node42003;
	wire [4-1:0] node42004;
	wire [4-1:0] node42007;
	wire [4-1:0] node42008;
	wire [4-1:0] node42012;
	wire [4-1:0] node42013;
	wire [4-1:0] node42015;
	wire [4-1:0] node42016;
	wire [4-1:0] node42020;
	wire [4-1:0] node42021;
	wire [4-1:0] node42023;
	wire [4-1:0] node42027;
	wire [4-1:0] node42028;
	wire [4-1:0] node42029;
	wire [4-1:0] node42030;
	wire [4-1:0] node42031;
	wire [4-1:0] node42034;
	wire [4-1:0] node42038;
	wire [4-1:0] node42039;
	wire [4-1:0] node42040;
	wire [4-1:0] node42043;
	wire [4-1:0] node42046;
	wire [4-1:0] node42048;
	wire [4-1:0] node42051;
	wire [4-1:0] node42052;
	wire [4-1:0] node42053;
	wire [4-1:0] node42054;
	wire [4-1:0] node42057;
	wire [4-1:0] node42060;
	wire [4-1:0] node42063;
	wire [4-1:0] node42064;
	wire [4-1:0] node42066;
	wire [4-1:0] node42070;
	wire [4-1:0] node42071;
	wire [4-1:0] node42072;
	wire [4-1:0] node42073;
	wire [4-1:0] node42074;
	wire [4-1:0] node42075;
	wire [4-1:0] node42080;
	wire [4-1:0] node42082;
	wire [4-1:0] node42083;
	wire [4-1:0] node42086;
	wire [4-1:0] node42089;
	wire [4-1:0] node42090;
	wire [4-1:0] node42092;
	wire [4-1:0] node42093;
	wire [4-1:0] node42096;
	wire [4-1:0] node42099;
	wire [4-1:0] node42101;
	wire [4-1:0] node42103;
	wire [4-1:0] node42106;
	wire [4-1:0] node42107;
	wire [4-1:0] node42108;
	wire [4-1:0] node42109;
	wire [4-1:0] node42112;
	wire [4-1:0] node42115;
	wire [4-1:0] node42116;
	wire [4-1:0] node42119;
	wire [4-1:0] node42120;
	wire [4-1:0] node42124;
	wire [4-1:0] node42125;
	wire [4-1:0] node42126;
	wire [4-1:0] node42127;
	wire [4-1:0] node42130;
	wire [4-1:0] node42133;
	wire [4-1:0] node42134;
	wire [4-1:0] node42137;
	wire [4-1:0] node42140;
	wire [4-1:0] node42141;
	wire [4-1:0] node42143;
	wire [4-1:0] node42146;
	wire [4-1:0] node42147;
	wire [4-1:0] node42150;
	wire [4-1:0] node42153;
	wire [4-1:0] node42154;
	wire [4-1:0] node42155;
	wire [4-1:0] node42156;
	wire [4-1:0] node42157;
	wire [4-1:0] node42158;
	wire [4-1:0] node42161;
	wire [4-1:0] node42164;
	wire [4-1:0] node42166;
	wire [4-1:0] node42167;
	wire [4-1:0] node42168;
	wire [4-1:0] node42173;
	wire [4-1:0] node42174;
	wire [4-1:0] node42175;
	wire [4-1:0] node42176;
	wire [4-1:0] node42177;
	wire [4-1:0] node42180;
	wire [4-1:0] node42183;
	wire [4-1:0] node42186;
	wire [4-1:0] node42187;
	wire [4-1:0] node42188;
	wire [4-1:0] node42193;
	wire [4-1:0] node42194;
	wire [4-1:0] node42195;
	wire [4-1:0] node42196;
	wire [4-1:0] node42199;
	wire [4-1:0] node42203;
	wire [4-1:0] node42204;
	wire [4-1:0] node42205;
	wire [4-1:0] node42209;
	wire [4-1:0] node42210;
	wire [4-1:0] node42213;
	wire [4-1:0] node42216;
	wire [4-1:0] node42217;
	wire [4-1:0] node42218;
	wire [4-1:0] node42219;
	wire [4-1:0] node42220;
	wire [4-1:0] node42223;
	wire [4-1:0] node42225;
	wire [4-1:0] node42228;
	wire [4-1:0] node42229;
	wire [4-1:0] node42230;
	wire [4-1:0] node42233;
	wire [4-1:0] node42236;
	wire [4-1:0] node42238;
	wire [4-1:0] node42241;
	wire [4-1:0] node42242;
	wire [4-1:0] node42244;
	wire [4-1:0] node42245;
	wire [4-1:0] node42249;
	wire [4-1:0] node42251;
	wire [4-1:0] node42254;
	wire [4-1:0] node42255;
	wire [4-1:0] node42256;
	wire [4-1:0] node42257;
	wire [4-1:0] node42258;
	wire [4-1:0] node42262;
	wire [4-1:0] node42265;
	wire [4-1:0] node42267;
	wire [4-1:0] node42270;
	wire [4-1:0] node42271;
	wire [4-1:0] node42272;
	wire [4-1:0] node42273;
	wire [4-1:0] node42276;
	wire [4-1:0] node42279;
	wire [4-1:0] node42280;
	wire [4-1:0] node42284;
	wire [4-1:0] node42287;
	wire [4-1:0] node42288;
	wire [4-1:0] node42289;
	wire [4-1:0] node42290;
	wire [4-1:0] node42291;
	wire [4-1:0] node42292;
	wire [4-1:0] node42295;
	wire [4-1:0] node42298;
	wire [4-1:0] node42299;
	wire [4-1:0] node42302;
	wire [4-1:0] node42305;
	wire [4-1:0] node42306;
	wire [4-1:0] node42308;
	wire [4-1:0] node42311;
	wire [4-1:0] node42314;
	wire [4-1:0] node42315;
	wire [4-1:0] node42316;
	wire [4-1:0] node42319;
	wire [4-1:0] node42320;
	wire [4-1:0] node42323;
	wire [4-1:0] node42324;
	wire [4-1:0] node42328;
	wire [4-1:0] node42329;
	wire [4-1:0] node42330;
	wire [4-1:0] node42331;
	wire [4-1:0] node42335;
	wire [4-1:0] node42336;
	wire [4-1:0] node42339;
	wire [4-1:0] node42342;
	wire [4-1:0] node42343;
	wire [4-1:0] node42344;
	wire [4-1:0] node42347;
	wire [4-1:0] node42351;
	wire [4-1:0] node42352;
	wire [4-1:0] node42353;
	wire [4-1:0] node42355;
	wire [4-1:0] node42357;
	wire [4-1:0] node42360;
	wire [4-1:0] node42361;
	wire [4-1:0] node42363;
	wire [4-1:0] node42366;
	wire [4-1:0] node42367;
	wire [4-1:0] node42371;
	wire [4-1:0] node42372;
	wire [4-1:0] node42373;
	wire [4-1:0] node42374;
	wire [4-1:0] node42377;
	wire [4-1:0] node42380;
	wire [4-1:0] node42382;
	wire [4-1:0] node42385;
	wire [4-1:0] node42386;
	wire [4-1:0] node42387;
	wire [4-1:0] node42389;
	wire [4-1:0] node42392;
	wire [4-1:0] node42393;
	wire [4-1:0] node42397;
	wire [4-1:0] node42398;
	wire [4-1:0] node42399;
	wire [4-1:0] node42402;
	wire [4-1:0] node42406;
	wire [4-1:0] node42407;
	wire [4-1:0] node42408;
	wire [4-1:0] node42409;
	wire [4-1:0] node42410;
	wire [4-1:0] node42411;
	wire [4-1:0] node42412;
	wire [4-1:0] node42413;
	wire [4-1:0] node42414;
	wire [4-1:0] node42417;
	wire [4-1:0] node42418;
	wire [4-1:0] node42419;
	wire [4-1:0] node42422;
	wire [4-1:0] node42425;
	wire [4-1:0] node42426;
	wire [4-1:0] node42429;
	wire [4-1:0] node42432;
	wire [4-1:0] node42433;
	wire [4-1:0] node42435;
	wire [4-1:0] node42436;
	wire [4-1:0] node42439;
	wire [4-1:0] node42442;
	wire [4-1:0] node42443;
	wire [4-1:0] node42444;
	wire [4-1:0] node42447;
	wire [4-1:0] node42450;
	wire [4-1:0] node42451;
	wire [4-1:0] node42455;
	wire [4-1:0] node42456;
	wire [4-1:0] node42457;
	wire [4-1:0] node42458;
	wire [4-1:0] node42462;
	wire [4-1:0] node42463;
	wire [4-1:0] node42464;
	wire [4-1:0] node42468;
	wire [4-1:0] node42469;
	wire [4-1:0] node42472;
	wire [4-1:0] node42475;
	wire [4-1:0] node42476;
	wire [4-1:0] node42477;
	wire [4-1:0] node42479;
	wire [4-1:0] node42483;
	wire [4-1:0] node42484;
	wire [4-1:0] node42488;
	wire [4-1:0] node42489;
	wire [4-1:0] node42490;
	wire [4-1:0] node42491;
	wire [4-1:0] node42493;
	wire [4-1:0] node42494;
	wire [4-1:0] node42497;
	wire [4-1:0] node42500;
	wire [4-1:0] node42502;
	wire [4-1:0] node42504;
	wire [4-1:0] node42507;
	wire [4-1:0] node42508;
	wire [4-1:0] node42510;
	wire [4-1:0] node42512;
	wire [4-1:0] node42516;
	wire [4-1:0] node42517;
	wire [4-1:0] node42518;
	wire [4-1:0] node42519;
	wire [4-1:0] node42522;
	wire [4-1:0] node42523;
	wire [4-1:0] node42526;
	wire [4-1:0] node42529;
	wire [4-1:0] node42530;
	wire [4-1:0] node42531;
	wire [4-1:0] node42534;
	wire [4-1:0] node42538;
	wire [4-1:0] node42540;
	wire [4-1:0] node42543;
	wire [4-1:0] node42544;
	wire [4-1:0] node42545;
	wire [4-1:0] node42546;
	wire [4-1:0] node42547;
	wire [4-1:0] node42550;
	wire [4-1:0] node42551;
	wire [4-1:0] node42553;
	wire [4-1:0] node42557;
	wire [4-1:0] node42559;
	wire [4-1:0] node42561;
	wire [4-1:0] node42564;
	wire [4-1:0] node42565;
	wire [4-1:0] node42566;
	wire [4-1:0] node42568;
	wire [4-1:0] node42570;
	wire [4-1:0] node42573;
	wire [4-1:0] node42575;
	wire [4-1:0] node42578;
	wire [4-1:0] node42579;
	wire [4-1:0] node42580;
	wire [4-1:0] node42582;
	wire [4-1:0] node42585;
	wire [4-1:0] node42587;
	wire [4-1:0] node42590;
	wire [4-1:0] node42591;
	wire [4-1:0] node42594;
	wire [4-1:0] node42597;
	wire [4-1:0] node42598;
	wire [4-1:0] node42599;
	wire [4-1:0] node42600;
	wire [4-1:0] node42603;
	wire [4-1:0] node42604;
	wire [4-1:0] node42605;
	wire [4-1:0] node42608;
	wire [4-1:0] node42611;
	wire [4-1:0] node42612;
	wire [4-1:0] node42615;
	wire [4-1:0] node42618;
	wire [4-1:0] node42619;
	wire [4-1:0] node42621;
	wire [4-1:0] node42624;
	wire [4-1:0] node42625;
	wire [4-1:0] node42627;
	wire [4-1:0] node42630;
	wire [4-1:0] node42632;
	wire [4-1:0] node42635;
	wire [4-1:0] node42636;
	wire [4-1:0] node42637;
	wire [4-1:0] node42639;
	wire [4-1:0] node42640;
	wire [4-1:0] node42644;
	wire [4-1:0] node42645;
	wire [4-1:0] node42646;
	wire [4-1:0] node42649;
	wire [4-1:0] node42653;
	wire [4-1:0] node42654;
	wire [4-1:0] node42655;
	wire [4-1:0] node42657;
	wire [4-1:0] node42660;
	wire [4-1:0] node42661;
	wire [4-1:0] node42665;
	wire [4-1:0] node42667;
	wire [4-1:0] node42670;
	wire [4-1:0] node42671;
	wire [4-1:0] node42672;
	wire [4-1:0] node42673;
	wire [4-1:0] node42674;
	wire [4-1:0] node42675;
	wire [4-1:0] node42677;
	wire [4-1:0] node42680;
	wire [4-1:0] node42681;
	wire [4-1:0] node42683;
	wire [4-1:0] node42686;
	wire [4-1:0] node42689;
	wire [4-1:0] node42690;
	wire [4-1:0] node42693;
	wire [4-1:0] node42694;
	wire [4-1:0] node42695;
	wire [4-1:0] node42699;
	wire [4-1:0] node42700;
	wire [4-1:0] node42704;
	wire [4-1:0] node42705;
	wire [4-1:0] node42706;
	wire [4-1:0] node42707;
	wire [4-1:0] node42708;
	wire [4-1:0] node42711;
	wire [4-1:0] node42714;
	wire [4-1:0] node42717;
	wire [4-1:0] node42718;
	wire [4-1:0] node42722;
	wire [4-1:0] node42723;
	wire [4-1:0] node42724;
	wire [4-1:0] node42726;
	wire [4-1:0] node42730;
	wire [4-1:0] node42731;
	wire [4-1:0] node42735;
	wire [4-1:0] node42736;
	wire [4-1:0] node42737;
	wire [4-1:0] node42738;
	wire [4-1:0] node42739;
	wire [4-1:0] node42742;
	wire [4-1:0] node42745;
	wire [4-1:0] node42746;
	wire [4-1:0] node42747;
	wire [4-1:0] node42752;
	wire [4-1:0] node42753;
	wire [4-1:0] node42754;
	wire [4-1:0] node42758;
	wire [4-1:0] node42759;
	wire [4-1:0] node42761;
	wire [4-1:0] node42764;
	wire [4-1:0] node42765;
	wire [4-1:0] node42768;
	wire [4-1:0] node42771;
	wire [4-1:0] node42772;
	wire [4-1:0] node42773;
	wire [4-1:0] node42774;
	wire [4-1:0] node42776;
	wire [4-1:0] node42779;
	wire [4-1:0] node42781;
	wire [4-1:0] node42784;
	wire [4-1:0] node42785;
	wire [4-1:0] node42789;
	wire [4-1:0] node42790;
	wire [4-1:0] node42791;
	wire [4-1:0] node42796;
	wire [4-1:0] node42797;
	wire [4-1:0] node42798;
	wire [4-1:0] node42799;
	wire [4-1:0] node42800;
	wire [4-1:0] node42801;
	wire [4-1:0] node42802;
	wire [4-1:0] node42805;
	wire [4-1:0] node42808;
	wire [4-1:0] node42809;
	wire [4-1:0] node42812;
	wire [4-1:0] node42815;
	wire [4-1:0] node42816;
	wire [4-1:0] node42819;
	wire [4-1:0] node42822;
	wire [4-1:0] node42823;
	wire [4-1:0] node42824;
	wire [4-1:0] node42827;
	wire [4-1:0] node42830;
	wire [4-1:0] node42832;
	wire [4-1:0] node42835;
	wire [4-1:0] node42836;
	wire [4-1:0] node42837;
	wire [4-1:0] node42839;
	wire [4-1:0] node42840;
	wire [4-1:0] node42843;
	wire [4-1:0] node42846;
	wire [4-1:0] node42847;
	wire [4-1:0] node42850;
	wire [4-1:0] node42852;
	wire [4-1:0] node42855;
	wire [4-1:0] node42856;
	wire [4-1:0] node42857;
	wire [4-1:0] node42858;
	wire [4-1:0] node42862;
	wire [4-1:0] node42863;
	wire [4-1:0] node42866;
	wire [4-1:0] node42869;
	wire [4-1:0] node42870;
	wire [4-1:0] node42874;
	wire [4-1:0] node42875;
	wire [4-1:0] node42876;
	wire [4-1:0] node42877;
	wire [4-1:0] node42879;
	wire [4-1:0] node42880;
	wire [4-1:0] node42884;
	wire [4-1:0] node42887;
	wire [4-1:0] node42888;
	wire [4-1:0] node42889;
	wire [4-1:0] node42891;
	wire [4-1:0] node42894;
	wire [4-1:0] node42896;
	wire [4-1:0] node42899;
	wire [4-1:0] node42901;
	wire [4-1:0] node42903;
	wire [4-1:0] node42906;
	wire [4-1:0] node42907;
	wire [4-1:0] node42908;
	wire [4-1:0] node42911;
	wire [4-1:0] node42914;
	wire [4-1:0] node42915;
	wire [4-1:0] node42916;
	wire [4-1:0] node42919;
	wire [4-1:0] node42922;
	wire [4-1:0] node42923;
	wire [4-1:0] node42925;
	wire [4-1:0] node42928;
	wire [4-1:0] node42929;
	wire [4-1:0] node42932;
	wire [4-1:0] node42935;
	wire [4-1:0] node42936;
	wire [4-1:0] node42937;
	wire [4-1:0] node42938;
	wire [4-1:0] node42939;
	wire [4-1:0] node42940;
	wire [4-1:0] node42941;
	wire [4-1:0] node42943;
	wire [4-1:0] node42946;
	wire [4-1:0] node42949;
	wire [4-1:0] node42950;
	wire [4-1:0] node42951;
	wire [4-1:0] node42952;
	wire [4-1:0] node42955;
	wire [4-1:0] node42959;
	wire [4-1:0] node42961;
	wire [4-1:0] node42964;
	wire [4-1:0] node42965;
	wire [4-1:0] node42966;
	wire [4-1:0] node42967;
	wire [4-1:0] node42970;
	wire [4-1:0] node42971;
	wire [4-1:0] node42974;
	wire [4-1:0] node42977;
	wire [4-1:0] node42978;
	wire [4-1:0] node42979;
	wire [4-1:0] node42982;
	wire [4-1:0] node42986;
	wire [4-1:0] node42987;
	wire [4-1:0] node42988;
	wire [4-1:0] node42989;
	wire [4-1:0] node42992;
	wire [4-1:0] node42995;
	wire [4-1:0] node42996;
	wire [4-1:0] node43000;
	wire [4-1:0] node43001;
	wire [4-1:0] node43005;
	wire [4-1:0] node43006;
	wire [4-1:0] node43007;
	wire [4-1:0] node43008;
	wire [4-1:0] node43009;
	wire [4-1:0] node43011;
	wire [4-1:0] node43014;
	wire [4-1:0] node43016;
	wire [4-1:0] node43019;
	wire [4-1:0] node43020;
	wire [4-1:0] node43023;
	wire [4-1:0] node43025;
	wire [4-1:0] node43028;
	wire [4-1:0] node43029;
	wire [4-1:0] node43031;
	wire [4-1:0] node43034;
	wire [4-1:0] node43035;
	wire [4-1:0] node43038;
	wire [4-1:0] node43041;
	wire [4-1:0] node43042;
	wire [4-1:0] node43043;
	wire [4-1:0] node43044;
	wire [4-1:0] node43048;
	wire [4-1:0] node43049;
	wire [4-1:0] node43053;
	wire [4-1:0] node43054;
	wire [4-1:0] node43055;
	wire [4-1:0] node43056;
	wire [4-1:0] node43059;
	wire [4-1:0] node43063;
	wire [4-1:0] node43064;
	wire [4-1:0] node43066;
	wire [4-1:0] node43069;
	wire [4-1:0] node43070;
	wire [4-1:0] node43073;
	wire [4-1:0] node43076;
	wire [4-1:0] node43077;
	wire [4-1:0] node43078;
	wire [4-1:0] node43079;
	wire [4-1:0] node43081;
	wire [4-1:0] node43082;
	wire [4-1:0] node43085;
	wire [4-1:0] node43088;
	wire [4-1:0] node43089;
	wire [4-1:0] node43090;
	wire [4-1:0] node43093;
	wire [4-1:0] node43096;
	wire [4-1:0] node43098;
	wire [4-1:0] node43101;
	wire [4-1:0] node43102;
	wire [4-1:0] node43103;
	wire [4-1:0] node43104;
	wire [4-1:0] node43107;
	wire [4-1:0] node43110;
	wire [4-1:0] node43112;
	wire [4-1:0] node43115;
	wire [4-1:0] node43116;
	wire [4-1:0] node43117;
	wire [4-1:0] node43118;
	wire [4-1:0] node43123;
	wire [4-1:0] node43124;
	wire [4-1:0] node43127;
	wire [4-1:0] node43130;
	wire [4-1:0] node43131;
	wire [4-1:0] node43132;
	wire [4-1:0] node43133;
	wire [4-1:0] node43135;
	wire [4-1:0] node43138;
	wire [4-1:0] node43141;
	wire [4-1:0] node43143;
	wire [4-1:0] node43146;
	wire [4-1:0] node43147;
	wire [4-1:0] node43148;
	wire [4-1:0] node43149;
	wire [4-1:0] node43153;
	wire [4-1:0] node43156;
	wire [4-1:0] node43157;
	wire [4-1:0] node43158;
	wire [4-1:0] node43162;
	wire [4-1:0] node43165;
	wire [4-1:0] node43166;
	wire [4-1:0] node43167;
	wire [4-1:0] node43168;
	wire [4-1:0] node43169;
	wire [4-1:0] node43171;
	wire [4-1:0] node43174;
	wire [4-1:0] node43176;
	wire [4-1:0] node43179;
	wire [4-1:0] node43180;
	wire [4-1:0] node43182;
	wire [4-1:0] node43185;
	wire [4-1:0] node43187;
	wire [4-1:0] node43190;
	wire [4-1:0] node43191;
	wire [4-1:0] node43192;
	wire [4-1:0] node43193;
	wire [4-1:0] node43194;
	wire [4-1:0] node43198;
	wire [4-1:0] node43199;
	wire [4-1:0] node43203;
	wire [4-1:0] node43204;
	wire [4-1:0] node43205;
	wire [4-1:0] node43209;
	wire [4-1:0] node43210;
	wire [4-1:0] node43214;
	wire [4-1:0] node43215;
	wire [4-1:0] node43217;
	wire [4-1:0] node43219;
	wire [4-1:0] node43222;
	wire [4-1:0] node43223;
	wire [4-1:0] node43226;
	wire [4-1:0] node43229;
	wire [4-1:0] node43230;
	wire [4-1:0] node43231;
	wire [4-1:0] node43232;
	wire [4-1:0] node43233;
	wire [4-1:0] node43237;
	wire [4-1:0] node43238;
	wire [4-1:0] node43242;
	wire [4-1:0] node43243;
	wire [4-1:0] node43244;
	wire [4-1:0] node43248;
	wire [4-1:0] node43250;
	wire [4-1:0] node43253;
	wire [4-1:0] node43254;
	wire [4-1:0] node43255;
	wire [4-1:0] node43256;
	wire [4-1:0] node43260;
	wire [4-1:0] node43261;
	wire [4-1:0] node43265;
	wire [4-1:0] node43266;
	wire [4-1:0] node43267;
	wire [4-1:0] node43271;
	wire [4-1:0] node43272;
	wire [4-1:0] node43276;
	wire [4-1:0] node43277;
	wire [4-1:0] node43278;
	wire [4-1:0] node43279;
	wire [4-1:0] node43280;
	wire [4-1:0] node43281;
	wire [4-1:0] node43282;
	wire [4-1:0] node43283;
	wire [4-1:0] node43284;
	wire [4-1:0] node43286;
	wire [4-1:0] node43291;
	wire [4-1:0] node43292;
	wire [4-1:0] node43294;
	wire [4-1:0] node43295;
	wire [4-1:0] node43298;
	wire [4-1:0] node43301;
	wire [4-1:0] node43303;
	wire [4-1:0] node43306;
	wire [4-1:0] node43307;
	wire [4-1:0] node43308;
	wire [4-1:0] node43309;
	wire [4-1:0] node43310;
	wire [4-1:0] node43313;
	wire [4-1:0] node43318;
	wire [4-1:0] node43319;
	wire [4-1:0] node43322;
	wire [4-1:0] node43324;
	wire [4-1:0] node43327;
	wire [4-1:0] node43328;
	wire [4-1:0] node43329;
	wire [4-1:0] node43330;
	wire [4-1:0] node43333;
	wire [4-1:0] node43336;
	wire [4-1:0] node43337;
	wire [4-1:0] node43338;
	wire [4-1:0] node43340;
	wire [4-1:0] node43345;
	wire [4-1:0] node43346;
	wire [4-1:0] node43347;
	wire [4-1:0] node43349;
	wire [4-1:0] node43352;
	wire [4-1:0] node43353;
	wire [4-1:0] node43354;
	wire [4-1:0] node43358;
	wire [4-1:0] node43360;
	wire [4-1:0] node43363;
	wire [4-1:0] node43364;
	wire [4-1:0] node43365;
	wire [4-1:0] node43369;
	wire [4-1:0] node43370;
	wire [4-1:0] node43373;
	wire [4-1:0] node43376;
	wire [4-1:0] node43377;
	wire [4-1:0] node43378;
	wire [4-1:0] node43379;
	wire [4-1:0] node43380;
	wire [4-1:0] node43381;
	wire [4-1:0] node43384;
	wire [4-1:0] node43386;
	wire [4-1:0] node43389;
	wire [4-1:0] node43390;
	wire [4-1:0] node43391;
	wire [4-1:0] node43396;
	wire [4-1:0] node43397;
	wire [4-1:0] node43398;
	wire [4-1:0] node43401;
	wire [4-1:0] node43402;
	wire [4-1:0] node43406;
	wire [4-1:0] node43407;
	wire [4-1:0] node43410;
	wire [4-1:0] node43413;
	wire [4-1:0] node43414;
	wire [4-1:0] node43415;
	wire [4-1:0] node43416;
	wire [4-1:0] node43419;
	wire [4-1:0] node43422;
	wire [4-1:0] node43423;
	wire [4-1:0] node43424;
	wire [4-1:0] node43428;
	wire [4-1:0] node43430;
	wire [4-1:0] node43433;
	wire [4-1:0] node43434;
	wire [4-1:0] node43436;
	wire [4-1:0] node43437;
	wire [4-1:0] node43440;
	wire [4-1:0] node43443;
	wire [4-1:0] node43444;
	wire [4-1:0] node43446;
	wire [4-1:0] node43449;
	wire [4-1:0] node43450;
	wire [4-1:0] node43453;
	wire [4-1:0] node43456;
	wire [4-1:0] node43457;
	wire [4-1:0] node43458;
	wire [4-1:0] node43460;
	wire [4-1:0] node43461;
	wire [4-1:0] node43464;
	wire [4-1:0] node43467;
	wire [4-1:0] node43468;
	wire [4-1:0] node43469;
	wire [4-1:0] node43473;
	wire [4-1:0] node43474;
	wire [4-1:0] node43477;
	wire [4-1:0] node43480;
	wire [4-1:0] node43481;
	wire [4-1:0] node43482;
	wire [4-1:0] node43485;
	wire [4-1:0] node43488;
	wire [4-1:0] node43489;
	wire [4-1:0] node43490;
	wire [4-1:0] node43494;
	wire [4-1:0] node43495;
	wire [4-1:0] node43496;
	wire [4-1:0] node43499;
	wire [4-1:0] node43503;
	wire [4-1:0] node43504;
	wire [4-1:0] node43505;
	wire [4-1:0] node43506;
	wire [4-1:0] node43507;
	wire [4-1:0] node43509;
	wire [4-1:0] node43512;
	wire [4-1:0] node43514;
	wire [4-1:0] node43517;
	wire [4-1:0] node43518;
	wire [4-1:0] node43520;
	wire [4-1:0] node43523;
	wire [4-1:0] node43525;
	wire [4-1:0] node43528;
	wire [4-1:0] node43529;
	wire [4-1:0] node43530;
	wire [4-1:0] node43531;
	wire [4-1:0] node43535;
	wire [4-1:0] node43536;
	wire [4-1:0] node43540;
	wire [4-1:0] node43541;
	wire [4-1:0] node43542;
	wire [4-1:0] node43546;
	wire [4-1:0] node43547;
	wire [4-1:0] node43551;
	wire [4-1:0] node43552;
	wire [4-1:0] node43553;
	wire [4-1:0] node43554;
	wire [4-1:0] node43555;
	wire [4-1:0] node43556;
	wire [4-1:0] node43560;
	wire [4-1:0] node43561;
	wire [4-1:0] node43565;
	wire [4-1:0] node43566;
	wire [4-1:0] node43567;
	wire [4-1:0] node43572;
	wire [4-1:0] node43573;
	wire [4-1:0] node43574;
	wire [4-1:0] node43575;
	wire [4-1:0] node43578;
	wire [4-1:0] node43581;
	wire [4-1:0] node43582;
	wire [4-1:0] node43585;
	wire [4-1:0] node43588;
	wire [4-1:0] node43589;
	wire [4-1:0] node43590;
	wire [4-1:0] node43593;
	wire [4-1:0] node43596;
	wire [4-1:0] node43598;
	wire [4-1:0] node43601;
	wire [4-1:0] node43602;
	wire [4-1:0] node43603;
	wire [4-1:0] node43604;
	wire [4-1:0] node43605;
	wire [4-1:0] node43608;
	wire [4-1:0] node43611;
	wire [4-1:0] node43612;
	wire [4-1:0] node43616;
	wire [4-1:0] node43617;
	wire [4-1:0] node43618;
	wire [4-1:0] node43621;
	wire [4-1:0] node43624;
	wire [4-1:0] node43626;
	wire [4-1:0] node43629;
	wire [4-1:0] node43630;
	wire [4-1:0] node43633;
	wire [4-1:0] node43636;
	wire [4-1:0] node43637;
	wire [4-1:0] node43638;
	wire [4-1:0] node43639;
	wire [4-1:0] node43640;
	wire [4-1:0] node43641;
	wire [4-1:0] node43642;
	wire [4-1:0] node43644;
	wire [4-1:0] node43647;
	wire [4-1:0] node43649;
	wire [4-1:0] node43652;
	wire [4-1:0] node43653;
	wire [4-1:0] node43656;
	wire [4-1:0] node43657;
	wire [4-1:0] node43661;
	wire [4-1:0] node43662;
	wire [4-1:0] node43664;
	wire [4-1:0] node43665;
	wire [4-1:0] node43668;
	wire [4-1:0] node43671;
	wire [4-1:0] node43672;
	wire [4-1:0] node43673;
	wire [4-1:0] node43674;
	wire [4-1:0] node43677;
	wire [4-1:0] node43681;
	wire [4-1:0] node43683;
	wire [4-1:0] node43686;
	wire [4-1:0] node43687;
	wire [4-1:0] node43688;
	wire [4-1:0] node43689;
	wire [4-1:0] node43690;
	wire [4-1:0] node43693;
	wire [4-1:0] node43696;
	wire [4-1:0] node43697;
	wire [4-1:0] node43700;
	wire [4-1:0] node43703;
	wire [4-1:0] node43704;
	wire [4-1:0] node43706;
	wire [4-1:0] node43710;
	wire [4-1:0] node43711;
	wire [4-1:0] node43712;
	wire [4-1:0] node43713;
	wire [4-1:0] node43715;
	wire [4-1:0] node43718;
	wire [4-1:0] node43720;
	wire [4-1:0] node43723;
	wire [4-1:0] node43724;
	wire [4-1:0] node43727;
	wire [4-1:0] node43729;
	wire [4-1:0] node43732;
	wire [4-1:0] node43733;
	wire [4-1:0] node43734;
	wire [4-1:0] node43738;
	wire [4-1:0] node43741;
	wire [4-1:0] node43742;
	wire [4-1:0] node43743;
	wire [4-1:0] node43744;
	wire [4-1:0] node43745;
	wire [4-1:0] node43748;
	wire [4-1:0] node43751;
	wire [4-1:0] node43752;
	wire [4-1:0] node43754;
	wire [4-1:0] node43755;
	wire [4-1:0] node43758;
	wire [4-1:0] node43761;
	wire [4-1:0] node43762;
	wire [4-1:0] node43763;
	wire [4-1:0] node43768;
	wire [4-1:0] node43769;
	wire [4-1:0] node43770;
	wire [4-1:0] node43771;
	wire [4-1:0] node43774;
	wire [4-1:0] node43777;
	wire [4-1:0] node43779;
	wire [4-1:0] node43780;
	wire [4-1:0] node43783;
	wire [4-1:0] node43786;
	wire [4-1:0] node43787;
	wire [4-1:0] node43788;
	wire [4-1:0] node43792;
	wire [4-1:0] node43793;
	wire [4-1:0] node43796;
	wire [4-1:0] node43799;
	wire [4-1:0] node43800;
	wire [4-1:0] node43801;
	wire [4-1:0] node43802;
	wire [4-1:0] node43804;
	wire [4-1:0] node43805;
	wire [4-1:0] node43809;
	wire [4-1:0] node43810;
	wire [4-1:0] node43813;
	wire [4-1:0] node43816;
	wire [4-1:0] node43817;
	wire [4-1:0] node43818;
	wire [4-1:0] node43821;
	wire [4-1:0] node43824;
	wire [4-1:0] node43825;
	wire [4-1:0] node43829;
	wire [4-1:0] node43830;
	wire [4-1:0] node43831;
	wire [4-1:0] node43834;
	wire [4-1:0] node43837;
	wire [4-1:0] node43838;
	wire [4-1:0] node43841;
	wire [4-1:0] node43844;
	wire [4-1:0] node43845;
	wire [4-1:0] node43846;
	wire [4-1:0] node43847;
	wire [4-1:0] node43848;
	wire [4-1:0] node43849;
	wire [4-1:0] node43852;
	wire [4-1:0] node43855;
	wire [4-1:0] node43856;
	wire [4-1:0] node43857;
	wire [4-1:0] node43860;
	wire [4-1:0] node43863;
	wire [4-1:0] node43865;
	wire [4-1:0] node43868;
	wire [4-1:0] node43869;
	wire [4-1:0] node43870;
	wire [4-1:0] node43873;
	wire [4-1:0] node43876;
	wire [4-1:0] node43878;
	wire [4-1:0] node43879;
	wire [4-1:0] node43881;
	wire [4-1:0] node43884;
	wire [4-1:0] node43885;
	wire [4-1:0] node43889;
	wire [4-1:0] node43890;
	wire [4-1:0] node43891;
	wire [4-1:0] node43892;
	wire [4-1:0] node43893;
	wire [4-1:0] node43894;
	wire [4-1:0] node43897;
	wire [4-1:0] node43901;
	wire [4-1:0] node43903;
	wire [4-1:0] node43906;
	wire [4-1:0] node43907;
	wire [4-1:0] node43908;
	wire [4-1:0] node43911;
	wire [4-1:0] node43914;
	wire [4-1:0] node43915;
	wire [4-1:0] node43918;
	wire [4-1:0] node43921;
	wire [4-1:0] node43922;
	wire [4-1:0] node43925;
	wire [4-1:0] node43928;
	wire [4-1:0] node43929;
	wire [4-1:0] node43930;
	wire [4-1:0] node43931;
	wire [4-1:0] node43932;
	wire [4-1:0] node43935;
	wire [4-1:0] node43938;
	wire [4-1:0] node43939;
	wire [4-1:0] node43940;
	wire [4-1:0] node43943;
	wire [4-1:0] node43947;
	wire [4-1:0] node43948;
	wire [4-1:0] node43951;
	wire [4-1:0] node43954;
	wire [4-1:0] node43955;
	wire [4-1:0] node43956;
	wire [4-1:0] node43957;
	wire [4-1:0] node43958;
	wire [4-1:0] node43963;
	wire [4-1:0] node43964;
	wire [4-1:0] node43965;
	wire [4-1:0] node43969;
	wire [4-1:0] node43972;
	wire [4-1:0] node43973;
	wire [4-1:0] node43974;
	wire [4-1:0] node43977;
	wire [4-1:0] node43978;
	wire [4-1:0] node43982;
	wire [4-1:0] node43983;
	wire [4-1:0] node43984;
	wire [4-1:0] node43988;
	wire [4-1:0] node43991;
	wire [4-1:0] node43992;
	wire [4-1:0] node43993;
	wire [4-1:0] node43994;
	wire [4-1:0] node43995;
	wire [4-1:0] node43996;
	wire [4-1:0] node43997;
	wire [4-1:0] node43998;
	wire [4-1:0] node43999;
	wire [4-1:0] node44000;
	wire [4-1:0] node44002;
	wire [4-1:0] node44005;
	wire [4-1:0] node44007;
	wire [4-1:0] node44010;
	wire [4-1:0] node44011;
	wire [4-1:0] node44013;
	wire [4-1:0] node44016;
	wire [4-1:0] node44018;
	wire [4-1:0] node44019;
	wire [4-1:0] node44022;
	wire [4-1:0] node44025;
	wire [4-1:0] node44026;
	wire [4-1:0] node44027;
	wire [4-1:0] node44029;
	wire [4-1:0] node44030;
	wire [4-1:0] node44034;
	wire [4-1:0] node44035;
	wire [4-1:0] node44036;
	wire [4-1:0] node44039;
	wire [4-1:0] node44042;
	wire [4-1:0] node44044;
	wire [4-1:0] node44047;
	wire [4-1:0] node44048;
	wire [4-1:0] node44049;
	wire [4-1:0] node44052;
	wire [4-1:0] node44055;
	wire [4-1:0] node44056;
	wire [4-1:0] node44059;
	wire [4-1:0] node44062;
	wire [4-1:0] node44063;
	wire [4-1:0] node44064;
	wire [4-1:0] node44065;
	wire [4-1:0] node44066;
	wire [4-1:0] node44068;
	wire [4-1:0] node44072;
	wire [4-1:0] node44073;
	wire [4-1:0] node44074;
	wire [4-1:0] node44078;
	wire [4-1:0] node44081;
	wire [4-1:0] node44082;
	wire [4-1:0] node44083;
	wire [4-1:0] node44087;
	wire [4-1:0] node44089;
	wire [4-1:0] node44090;
	wire [4-1:0] node44093;
	wire [4-1:0] node44096;
	wire [4-1:0] node44097;
	wire [4-1:0] node44098;
	wire [4-1:0] node44099;
	wire [4-1:0] node44102;
	wire [4-1:0] node44105;
	wire [4-1:0] node44106;
	wire [4-1:0] node44110;
	wire [4-1:0] node44112;
	wire [4-1:0] node44113;
	wire [4-1:0] node44115;
	wire [4-1:0] node44118;
	wire [4-1:0] node44119;
	wire [4-1:0] node44123;
	wire [4-1:0] node44124;
	wire [4-1:0] node44125;
	wire [4-1:0] node44126;
	wire [4-1:0] node44127;
	wire [4-1:0] node44128;
	wire [4-1:0] node44132;
	wire [4-1:0] node44133;
	wire [4-1:0] node44134;
	wire [4-1:0] node44139;
	wire [4-1:0] node44140;
	wire [4-1:0] node44141;
	wire [4-1:0] node44146;
	wire [4-1:0] node44147;
	wire [4-1:0] node44148;
	wire [4-1:0] node44150;
	wire [4-1:0] node44153;
	wire [4-1:0] node44154;
	wire [4-1:0] node44155;
	wire [4-1:0] node44158;
	wire [4-1:0] node44161;
	wire [4-1:0] node44163;
	wire [4-1:0] node44166;
	wire [4-1:0] node44167;
	wire [4-1:0] node44168;
	wire [4-1:0] node44172;
	wire [4-1:0] node44173;
	wire [4-1:0] node44177;
	wire [4-1:0] node44178;
	wire [4-1:0] node44179;
	wire [4-1:0] node44181;
	wire [4-1:0] node44183;
	wire [4-1:0] node44186;
	wire [4-1:0] node44187;
	wire [4-1:0] node44188;
	wire [4-1:0] node44192;
	wire [4-1:0] node44193;
	wire [4-1:0] node44194;
	wire [4-1:0] node44199;
	wire [4-1:0] node44200;
	wire [4-1:0] node44201;
	wire [4-1:0] node44202;
	wire [4-1:0] node44203;
	wire [4-1:0] node44209;
	wire [4-1:0] node44210;
	wire [4-1:0] node44211;
	wire [4-1:0] node44212;
	wire [4-1:0] node44215;
	wire [4-1:0] node44218;
	wire [4-1:0] node44219;
	wire [4-1:0] node44222;
	wire [4-1:0] node44225;
	wire [4-1:0] node44226;
	wire [4-1:0] node44227;
	wire [4-1:0] node44232;
	wire [4-1:0] node44233;
	wire [4-1:0] node44234;
	wire [4-1:0] node44235;
	wire [4-1:0] node44236;
	wire [4-1:0] node44237;
	wire [4-1:0] node44238;
	wire [4-1:0] node44241;
	wire [4-1:0] node44244;
	wire [4-1:0] node44246;
	wire [4-1:0] node44249;
	wire [4-1:0] node44250;
	wire [4-1:0] node44251;
	wire [4-1:0] node44254;
	wire [4-1:0] node44257;
	wire [4-1:0] node44258;
	wire [4-1:0] node44259;
	wire [4-1:0] node44262;
	wire [4-1:0] node44266;
	wire [4-1:0] node44267;
	wire [4-1:0] node44269;
	wire [4-1:0] node44272;
	wire [4-1:0] node44273;
	wire [4-1:0] node44274;
	wire [4-1:0] node44277;
	wire [4-1:0] node44280;
	wire [4-1:0] node44281;
	wire [4-1:0] node44284;
	wire [4-1:0] node44287;
	wire [4-1:0] node44288;
	wire [4-1:0] node44289;
	wire [4-1:0] node44290;
	wire [4-1:0] node44292;
	wire [4-1:0] node44295;
	wire [4-1:0] node44297;
	wire [4-1:0] node44300;
	wire [4-1:0] node44303;
	wire [4-1:0] node44304;
	wire [4-1:0] node44305;
	wire [4-1:0] node44306;
	wire [4-1:0] node44311;
	wire [4-1:0] node44312;
	wire [4-1:0] node44313;
	wire [4-1:0] node44317;
	wire [4-1:0] node44318;
	wire [4-1:0] node44322;
	wire [4-1:0] node44323;
	wire [4-1:0] node44324;
	wire [4-1:0] node44325;
	wire [4-1:0] node44326;
	wire [4-1:0] node44327;
	wire [4-1:0] node44331;
	wire [4-1:0] node44332;
	wire [4-1:0] node44335;
	wire [4-1:0] node44338;
	wire [4-1:0] node44339;
	wire [4-1:0] node44340;
	wire [4-1:0] node44341;
	wire [4-1:0] node44346;
	wire [4-1:0] node44349;
	wire [4-1:0] node44350;
	wire [4-1:0] node44351;
	wire [4-1:0] node44353;
	wire [4-1:0] node44354;
	wire [4-1:0] node44358;
	wire [4-1:0] node44359;
	wire [4-1:0] node44362;
	wire [4-1:0] node44365;
	wire [4-1:0] node44366;
	wire [4-1:0] node44367;
	wire [4-1:0] node44371;
	wire [4-1:0] node44372;
	wire [4-1:0] node44375;
	wire [4-1:0] node44378;
	wire [4-1:0] node44379;
	wire [4-1:0] node44380;
	wire [4-1:0] node44381;
	wire [4-1:0] node44382;
	wire [4-1:0] node44385;
	wire [4-1:0] node44388;
	wire [4-1:0] node44389;
	wire [4-1:0] node44392;
	wire [4-1:0] node44395;
	wire [4-1:0] node44396;
	wire [4-1:0] node44398;
	wire [4-1:0] node44399;
	wire [4-1:0] node44402;
	wire [4-1:0] node44405;
	wire [4-1:0] node44406;
	wire [4-1:0] node44407;
	wire [4-1:0] node44410;
	wire [4-1:0] node44414;
	wire [4-1:0] node44415;
	wire [4-1:0] node44416;
	wire [4-1:0] node44419;
	wire [4-1:0] node44421;
	wire [4-1:0] node44422;
	wire [4-1:0] node44426;
	wire [4-1:0] node44427;
	wire [4-1:0] node44429;
	wire [4-1:0] node44432;
	wire [4-1:0] node44433;
	wire [4-1:0] node44436;
	wire [4-1:0] node44439;
	wire [4-1:0] node44440;
	wire [4-1:0] node44441;
	wire [4-1:0] node44442;
	wire [4-1:0] node44443;
	wire [4-1:0] node44444;
	wire [4-1:0] node44445;
	wire [4-1:0] node44446;
	wire [4-1:0] node44449;
	wire [4-1:0] node44452;
	wire [4-1:0] node44453;
	wire [4-1:0] node44455;
	wire [4-1:0] node44458;
	wire [4-1:0] node44460;
	wire [4-1:0] node44463;
	wire [4-1:0] node44464;
	wire [4-1:0] node44466;
	wire [4-1:0] node44468;
	wire [4-1:0] node44471;
	wire [4-1:0] node44472;
	wire [4-1:0] node44475;
	wire [4-1:0] node44478;
	wire [4-1:0] node44479;
	wire [4-1:0] node44481;
	wire [4-1:0] node44482;
	wire [4-1:0] node44485;
	wire [4-1:0] node44486;
	wire [4-1:0] node44489;
	wire [4-1:0] node44492;
	wire [4-1:0] node44493;
	wire [4-1:0] node44494;
	wire [4-1:0] node44496;
	wire [4-1:0] node44499;
	wire [4-1:0] node44502;
	wire [4-1:0] node44505;
	wire [4-1:0] node44506;
	wire [4-1:0] node44507;
	wire [4-1:0] node44508;
	wire [4-1:0] node44509;
	wire [4-1:0] node44512;
	wire [4-1:0] node44515;
	wire [4-1:0] node44516;
	wire [4-1:0] node44517;
	wire [4-1:0] node44521;
	wire [4-1:0] node44522;
	wire [4-1:0] node44525;
	wire [4-1:0] node44528;
	wire [4-1:0] node44529;
	wire [4-1:0] node44531;
	wire [4-1:0] node44534;
	wire [4-1:0] node44535;
	wire [4-1:0] node44536;
	wire [4-1:0] node44539;
	wire [4-1:0] node44543;
	wire [4-1:0] node44544;
	wire [4-1:0] node44545;
	wire [4-1:0] node44546;
	wire [4-1:0] node44547;
	wire [4-1:0] node44551;
	wire [4-1:0] node44555;
	wire [4-1:0] node44556;
	wire [4-1:0] node44557;
	wire [4-1:0] node44560;
	wire [4-1:0] node44563;
	wire [4-1:0] node44564;
	wire [4-1:0] node44567;
	wire [4-1:0] node44568;
	wire [4-1:0] node44572;
	wire [4-1:0] node44573;
	wire [4-1:0] node44574;
	wire [4-1:0] node44575;
	wire [4-1:0] node44576;
	wire [4-1:0] node44577;
	wire [4-1:0] node44580;
	wire [4-1:0] node44583;
	wire [4-1:0] node44584;
	wire [4-1:0] node44587;
	wire [4-1:0] node44590;
	wire [4-1:0] node44591;
	wire [4-1:0] node44592;
	wire [4-1:0] node44595;
	wire [4-1:0] node44598;
	wire [4-1:0] node44599;
	wire [4-1:0] node44602;
	wire [4-1:0] node44605;
	wire [4-1:0] node44606;
	wire [4-1:0] node44607;
	wire [4-1:0] node44608;
	wire [4-1:0] node44611;
	wire [4-1:0] node44615;
	wire [4-1:0] node44616;
	wire [4-1:0] node44617;
	wire [4-1:0] node44620;
	wire [4-1:0] node44621;
	wire [4-1:0] node44625;
	wire [4-1:0] node44626;
	wire [4-1:0] node44629;
	wire [4-1:0] node44632;
	wire [4-1:0] node44633;
	wire [4-1:0] node44634;
	wire [4-1:0] node44635;
	wire [4-1:0] node44636;
	wire [4-1:0] node44639;
	wire [4-1:0] node44642;
	wire [4-1:0] node44643;
	wire [4-1:0] node44647;
	wire [4-1:0] node44648;
	wire [4-1:0] node44651;
	wire [4-1:0] node44654;
	wire [4-1:0] node44655;
	wire [4-1:0] node44656;
	wire [4-1:0] node44659;
	wire [4-1:0] node44662;
	wire [4-1:0] node44663;
	wire [4-1:0] node44666;
	wire [4-1:0] node44669;
	wire [4-1:0] node44670;
	wire [4-1:0] node44671;
	wire [4-1:0] node44672;
	wire [4-1:0] node44673;
	wire [4-1:0] node44674;
	wire [4-1:0] node44675;
	wire [4-1:0] node44678;
	wire [4-1:0] node44681;
	wire [4-1:0] node44682;
	wire [4-1:0] node44685;
	wire [4-1:0] node44688;
	wire [4-1:0] node44689;
	wire [4-1:0] node44692;
	wire [4-1:0] node44695;
	wire [4-1:0] node44696;
	wire [4-1:0] node44697;
	wire [4-1:0] node44700;
	wire [4-1:0] node44703;
	wire [4-1:0] node44704;
	wire [4-1:0] node44706;
	wire [4-1:0] node44709;
	wire [4-1:0] node44710;
	wire [4-1:0] node44713;
	wire [4-1:0] node44716;
	wire [4-1:0] node44717;
	wire [4-1:0] node44718;
	wire [4-1:0] node44720;
	wire [4-1:0] node44723;
	wire [4-1:0] node44724;
	wire [4-1:0] node44727;
	wire [4-1:0] node44730;
	wire [4-1:0] node44731;
	wire [4-1:0] node44732;
	wire [4-1:0] node44735;
	wire [4-1:0] node44738;
	wire [4-1:0] node44739;
	wire [4-1:0] node44740;
	wire [4-1:0] node44741;
	wire [4-1:0] node44744;
	wire [4-1:0] node44747;
	wire [4-1:0] node44748;
	wire [4-1:0] node44751;
	wire [4-1:0] node44754;
	wire [4-1:0] node44755;
	wire [4-1:0] node44756;
	wire [4-1:0] node44759;
	wire [4-1:0] node44762;
	wire [4-1:0] node44763;
	wire [4-1:0] node44766;
	wire [4-1:0] node44769;
	wire [4-1:0] node44770;
	wire [4-1:0] node44771;
	wire [4-1:0] node44772;
	wire [4-1:0] node44773;
	wire [4-1:0] node44774;
	wire [4-1:0] node44777;
	wire [4-1:0] node44780;
	wire [4-1:0] node44782;
	wire [4-1:0] node44785;
	wire [4-1:0] node44786;
	wire [4-1:0] node44789;
	wire [4-1:0] node44792;
	wire [4-1:0] node44793;
	wire [4-1:0] node44794;
	wire [4-1:0] node44797;
	wire [4-1:0] node44800;
	wire [4-1:0] node44801;
	wire [4-1:0] node44804;
	wire [4-1:0] node44807;
	wire [4-1:0] node44808;
	wire [4-1:0] node44809;
	wire [4-1:0] node44810;
	wire [4-1:0] node44811;
	wire [4-1:0] node44815;
	wire [4-1:0] node44817;
	wire [4-1:0] node44820;
	wire [4-1:0] node44821;
	wire [4-1:0] node44824;
	wire [4-1:0] node44827;
	wire [4-1:0] node44828;
	wire [4-1:0] node44829;
	wire [4-1:0] node44832;
	wire [4-1:0] node44835;
	wire [4-1:0] node44836;
	wire [4-1:0] node44837;
	wire [4-1:0] node44838;
	wire [4-1:0] node44841;
	wire [4-1:0] node44844;
	wire [4-1:0] node44845;
	wire [4-1:0] node44848;
	wire [4-1:0] node44851;
	wire [4-1:0] node44852;
	wire [4-1:0] node44855;
	wire [4-1:0] node44858;
	wire [4-1:0] node44859;
	wire [4-1:0] node44860;
	wire [4-1:0] node44861;
	wire [4-1:0] node44862;
	wire [4-1:0] node44863;
	wire [4-1:0] node44864;
	wire [4-1:0] node44865;
	wire [4-1:0] node44868;
	wire [4-1:0] node44869;
	wire [4-1:0] node44871;
	wire [4-1:0] node44874;
	wire [4-1:0] node44875;
	wire [4-1:0] node44878;
	wire [4-1:0] node44881;
	wire [4-1:0] node44882;
	wire [4-1:0] node44883;
	wire [4-1:0] node44884;
	wire [4-1:0] node44888;
	wire [4-1:0] node44890;
	wire [4-1:0] node44893;
	wire [4-1:0] node44894;
	wire [4-1:0] node44898;
	wire [4-1:0] node44899;
	wire [4-1:0] node44901;
	wire [4-1:0] node44902;
	wire [4-1:0] node44904;
	wire [4-1:0] node44908;
	wire [4-1:0] node44909;
	wire [4-1:0] node44910;
	wire [4-1:0] node44913;
	wire [4-1:0] node44916;
	wire [4-1:0] node44918;
	wire [4-1:0] node44921;
	wire [4-1:0] node44922;
	wire [4-1:0] node44923;
	wire [4-1:0] node44924;
	wire [4-1:0] node44925;
	wire [4-1:0] node44926;
	wire [4-1:0] node44929;
	wire [4-1:0] node44933;
	wire [4-1:0] node44934;
	wire [4-1:0] node44935;
	wire [4-1:0] node44938;
	wire [4-1:0] node44941;
	wire [4-1:0] node44944;
	wire [4-1:0] node44945;
	wire [4-1:0] node44946;
	wire [4-1:0] node44949;
	wire [4-1:0] node44952;
	wire [4-1:0] node44953;
	wire [4-1:0] node44955;
	wire [4-1:0] node44959;
	wire [4-1:0] node44960;
	wire [4-1:0] node44961;
	wire [4-1:0] node44962;
	wire [4-1:0] node44965;
	wire [4-1:0] node44968;
	wire [4-1:0] node44970;
	wire [4-1:0] node44973;
	wire [4-1:0] node44974;
	wire [4-1:0] node44977;
	wire [4-1:0] node44979;
	wire [4-1:0] node44980;
	wire [4-1:0] node44983;
	wire [4-1:0] node44986;
	wire [4-1:0] node44987;
	wire [4-1:0] node44988;
	wire [4-1:0] node44989;
	wire [4-1:0] node44990;
	wire [4-1:0] node44991;
	wire [4-1:0] node44994;
	wire [4-1:0] node44997;
	wire [4-1:0] node44998;
	wire [4-1:0] node45002;
	wire [4-1:0] node45003;
	wire [4-1:0] node45004;
	wire [4-1:0] node45005;
	wire [4-1:0] node45008;
	wire [4-1:0] node45011;
	wire [4-1:0] node45012;
	wire [4-1:0] node45017;
	wire [4-1:0] node45018;
	wire [4-1:0] node45019;
	wire [4-1:0] node45020;
	wire [4-1:0] node45024;
	wire [4-1:0] node45025;
	wire [4-1:0] node45027;
	wire [4-1:0] node45030;
	wire [4-1:0] node45031;
	wire [4-1:0] node45035;
	wire [4-1:0] node45036;
	wire [4-1:0] node45037;
	wire [4-1:0] node45040;
	wire [4-1:0] node45043;
	wire [4-1:0] node45044;
	wire [4-1:0] node45045;
	wire [4-1:0] node45048;
	wire [4-1:0] node45051;
	wire [4-1:0] node45053;
	wire [4-1:0] node45056;
	wire [4-1:0] node45057;
	wire [4-1:0] node45058;
	wire [4-1:0] node45059;
	wire [4-1:0] node45060;
	wire [4-1:0] node45062;
	wire [4-1:0] node45065;
	wire [4-1:0] node45066;
	wire [4-1:0] node45069;
	wire [4-1:0] node45072;
	wire [4-1:0] node45073;
	wire [4-1:0] node45074;
	wire [4-1:0] node45077;
	wire [4-1:0] node45080;
	wire [4-1:0] node45081;
	wire [4-1:0] node45085;
	wire [4-1:0] node45086;
	wire [4-1:0] node45087;
	wire [4-1:0] node45090;
	wire [4-1:0] node45094;
	wire [4-1:0] node45095;
	wire [4-1:0] node45096;
	wire [4-1:0] node45097;
	wire [4-1:0] node45101;
	wire [4-1:0] node45102;
	wire [4-1:0] node45106;
	wire [4-1:0] node45107;
	wire [4-1:0] node45110;
	wire [4-1:0] node45112;
	wire [4-1:0] node45113;
	wire [4-1:0] node45117;
	wire [4-1:0] node45118;
	wire [4-1:0] node45119;
	wire [4-1:0] node45120;
	wire [4-1:0] node45121;
	wire [4-1:0] node45122;
	wire [4-1:0] node45125;
	wire [4-1:0] node45128;
	wire [4-1:0] node45129;
	wire [4-1:0] node45130;
	wire [4-1:0] node45134;
	wire [4-1:0] node45135;
	wire [4-1:0] node45138;
	wire [4-1:0] node45141;
	wire [4-1:0] node45142;
	wire [4-1:0] node45143;
	wire [4-1:0] node45144;
	wire [4-1:0] node45148;
	wire [4-1:0] node45151;
	wire [4-1:0] node45152;
	wire [4-1:0] node45153;
	wire [4-1:0] node45157;
	wire [4-1:0] node45160;
	wire [4-1:0] node45161;
	wire [4-1:0] node45162;
	wire [4-1:0] node45163;
	wire [4-1:0] node45164;
	wire [4-1:0] node45168;
	wire [4-1:0] node45169;
	wire [4-1:0] node45173;
	wire [4-1:0] node45174;
	wire [4-1:0] node45175;
	wire [4-1:0] node45179;
	wire [4-1:0] node45180;
	wire [4-1:0] node45184;
	wire [4-1:0] node45185;
	wire [4-1:0] node45186;
	wire [4-1:0] node45187;
	wire [4-1:0] node45190;
	wire [4-1:0] node45193;
	wire [4-1:0] node45194;
	wire [4-1:0] node45197;
	wire [4-1:0] node45200;
	wire [4-1:0] node45201;
	wire [4-1:0] node45202;
	wire [4-1:0] node45205;
	wire [4-1:0] node45208;
	wire [4-1:0] node45210;
	wire [4-1:0] node45213;
	wire [4-1:0] node45214;
	wire [4-1:0] node45215;
	wire [4-1:0] node45216;
	wire [4-1:0] node45217;
	wire [4-1:0] node45218;
	wire [4-1:0] node45219;
	wire [4-1:0] node45222;
	wire [4-1:0] node45225;
	wire [4-1:0] node45226;
	wire [4-1:0] node45229;
	wire [4-1:0] node45232;
	wire [4-1:0] node45233;
	wire [4-1:0] node45236;
	wire [4-1:0] node45239;
	wire [4-1:0] node45240;
	wire [4-1:0] node45241;
	wire [4-1:0] node45244;
	wire [4-1:0] node45247;
	wire [4-1:0] node45248;
	wire [4-1:0] node45251;
	wire [4-1:0] node45254;
	wire [4-1:0] node45255;
	wire [4-1:0] node45256;
	wire [4-1:0] node45257;
	wire [4-1:0] node45261;
	wire [4-1:0] node45262;
	wire [4-1:0] node45263;
	wire [4-1:0] node45266;
	wire [4-1:0] node45269;
	wire [4-1:0] node45272;
	wire [4-1:0] node45273;
	wire [4-1:0] node45276;
	wire [4-1:0] node45278;
	wire [4-1:0] node45280;
	wire [4-1:0] node45283;
	wire [4-1:0] node45284;
	wire [4-1:0] node45285;
	wire [4-1:0] node45286;
	wire [4-1:0] node45288;
	wire [4-1:0] node45291;
	wire [4-1:0] node45292;
	wire [4-1:0] node45295;
	wire [4-1:0] node45298;
	wire [4-1:0] node45299;
	wire [4-1:0] node45303;
	wire [4-1:0] node45304;
	wire [4-1:0] node45305;
	wire [4-1:0] node45309;
	wire [4-1:0] node45310;
	wire [4-1:0] node45311;
	wire [4-1:0] node45314;
	wire [4-1:0] node45317;
	wire [4-1:0] node45318;
	wire [4-1:0] node45321;
	wire [4-1:0] node45324;
	wire [4-1:0] node45325;
	wire [4-1:0] node45326;
	wire [4-1:0] node45327;
	wire [4-1:0] node45328;
	wire [4-1:0] node45329;
	wire [4-1:0] node45330;
	wire [4-1:0] node45333;
	wire [4-1:0] node45335;
	wire [4-1:0] node45338;
	wire [4-1:0] node45339;
	wire [4-1:0] node45340;
	wire [4-1:0] node45341;
	wire [4-1:0] node45344;
	wire [4-1:0] node45348;
	wire [4-1:0] node45349;
	wire [4-1:0] node45352;
	wire [4-1:0] node45355;
	wire [4-1:0] node45356;
	wire [4-1:0] node45357;
	wire [4-1:0] node45360;
	wire [4-1:0] node45361;
	wire [4-1:0] node45363;
	wire [4-1:0] node45366;
	wire [4-1:0] node45367;
	wire [4-1:0] node45370;
	wire [4-1:0] node45373;
	wire [4-1:0] node45374;
	wire [4-1:0] node45375;
	wire [4-1:0] node45379;
	wire [4-1:0] node45380;
	wire [4-1:0] node45383;
	wire [4-1:0] node45386;
	wire [4-1:0] node45387;
	wire [4-1:0] node45388;
	wire [4-1:0] node45389;
	wire [4-1:0] node45390;
	wire [4-1:0] node45394;
	wire [4-1:0] node45395;
	wire [4-1:0] node45396;
	wire [4-1:0] node45399;
	wire [4-1:0] node45402;
	wire [4-1:0] node45404;
	wire [4-1:0] node45407;
	wire [4-1:0] node45408;
	wire [4-1:0] node45409;
	wire [4-1:0] node45413;
	wire [4-1:0] node45414;
	wire [4-1:0] node45417;
	wire [4-1:0] node45420;
	wire [4-1:0] node45421;
	wire [4-1:0] node45422;
	wire [4-1:0] node45423;
	wire [4-1:0] node45424;
	wire [4-1:0] node45427;
	wire [4-1:0] node45430;
	wire [4-1:0] node45431;
	wire [4-1:0] node45435;
	wire [4-1:0] node45436;
	wire [4-1:0] node45438;
	wire [4-1:0] node45441;
	wire [4-1:0] node45442;
	wire [4-1:0] node45445;
	wire [4-1:0] node45448;
	wire [4-1:0] node45449;
	wire [4-1:0] node45450;
	wire [4-1:0] node45451;
	wire [4-1:0] node45454;
	wire [4-1:0] node45457;
	wire [4-1:0] node45458;
	wire [4-1:0] node45462;
	wire [4-1:0] node45465;
	wire [4-1:0] node45466;
	wire [4-1:0] node45467;
	wire [4-1:0] node45468;
	wire [4-1:0] node45469;
	wire [4-1:0] node45470;
	wire [4-1:0] node45471;
	wire [4-1:0] node45475;
	wire [4-1:0] node45476;
	wire [4-1:0] node45480;
	wire [4-1:0] node45481;
	wire [4-1:0] node45484;
	wire [4-1:0] node45487;
	wire [4-1:0] node45488;
	wire [4-1:0] node45490;
	wire [4-1:0] node45491;
	wire [4-1:0] node45495;
	wire [4-1:0] node45496;
	wire [4-1:0] node45499;
	wire [4-1:0] node45502;
	wire [4-1:0] node45503;
	wire [4-1:0] node45504;
	wire [4-1:0] node45506;
	wire [4-1:0] node45507;
	wire [4-1:0] node45510;
	wire [4-1:0] node45513;
	wire [4-1:0] node45515;
	wire [4-1:0] node45518;
	wire [4-1:0] node45519;
	wire [4-1:0] node45521;
	wire [4-1:0] node45523;
	wire [4-1:0] node45526;
	wire [4-1:0] node45527;
	wire [4-1:0] node45530;
	wire [4-1:0] node45533;
	wire [4-1:0] node45534;
	wire [4-1:0] node45535;
	wire [4-1:0] node45537;
	wire [4-1:0] node45540;
	wire [4-1:0] node45541;
	wire [4-1:0] node45543;
	wire [4-1:0] node45546;
	wire [4-1:0] node45547;
	wire [4-1:0] node45551;
	wire [4-1:0] node45552;
	wire [4-1:0] node45553;
	wire [4-1:0] node45554;
	wire [4-1:0] node45558;
	wire [4-1:0] node45561;
	wire [4-1:0] node45562;
	wire [4-1:0] node45563;
	wire [4-1:0] node45567;
	wire [4-1:0] node45568;
	wire [4-1:0] node45572;
	wire [4-1:0] node45573;
	wire [4-1:0] node45574;
	wire [4-1:0] node45575;
	wire [4-1:0] node45576;
	wire [4-1:0] node45577;
	wire [4-1:0] node45578;
	wire [4-1:0] node45581;
	wire [4-1:0] node45584;
	wire [4-1:0] node45585;
	wire [4-1:0] node45586;
	wire [4-1:0] node45589;
	wire [4-1:0] node45593;
	wire [4-1:0] node45594;
	wire [4-1:0] node45597;
	wire [4-1:0] node45600;
	wire [4-1:0] node45601;
	wire [4-1:0] node45602;
	wire [4-1:0] node45603;
	wire [4-1:0] node45606;
	wire [4-1:0] node45609;
	wire [4-1:0] node45610;
	wire [4-1:0] node45613;
	wire [4-1:0] node45616;
	wire [4-1:0] node45617;
	wire [4-1:0] node45618;
	wire [4-1:0] node45621;
	wire [4-1:0] node45624;
	wire [4-1:0] node45625;
	wire [4-1:0] node45629;
	wire [4-1:0] node45630;
	wire [4-1:0] node45631;
	wire [4-1:0] node45632;
	wire [4-1:0] node45636;
	wire [4-1:0] node45637;
	wire [4-1:0] node45641;
	wire [4-1:0] node45642;
	wire [4-1:0] node45643;
	wire [4-1:0] node45647;
	wire [4-1:0] node45648;
	wire [4-1:0] node45652;
	wire [4-1:0] node45653;
	wire [4-1:0] node45654;
	wire [4-1:0] node45655;
	wire [4-1:0] node45657;
	wire [4-1:0] node45658;
	wire [4-1:0] node45661;
	wire [4-1:0] node45664;
	wire [4-1:0] node45665;
	wire [4-1:0] node45667;
	wire [4-1:0] node45670;
	wire [4-1:0] node45672;
	wire [4-1:0] node45675;
	wire [4-1:0] node45676;
	wire [4-1:0] node45677;
	wire [4-1:0] node45679;
	wire [4-1:0] node45682;
	wire [4-1:0] node45683;
	wire [4-1:0] node45685;
	wire [4-1:0] node45688;
	wire [4-1:0] node45691;
	wire [4-1:0] node45692;
	wire [4-1:0] node45694;
	wire [4-1:0] node45697;
	wire [4-1:0] node45698;
	wire [4-1:0] node45702;
	wire [4-1:0] node45703;
	wire [4-1:0] node45704;
	wire [4-1:0] node45705;
	wire [4-1:0] node45706;
	wire [4-1:0] node45707;
	wire [4-1:0] node45711;
	wire [4-1:0] node45712;
	wire [4-1:0] node45716;
	wire [4-1:0] node45718;
	wire [4-1:0] node45719;
	wire [4-1:0] node45723;
	wire [4-1:0] node45725;
	wire [4-1:0] node45726;
	wire [4-1:0] node45729;
	wire [4-1:0] node45732;
	wire [4-1:0] node45733;
	wire [4-1:0] node45734;
	wire [4-1:0] node45738;
	wire [4-1:0] node45739;
	wire [4-1:0] node45740;
	wire [4-1:0] node45744;
	wire [4-1:0] node45745;
	wire [4-1:0] node45749;
	wire [4-1:0] node45750;
	wire [4-1:0] node45751;
	wire [4-1:0] node45752;
	wire [4-1:0] node45753;
	wire [4-1:0] node45754;
	wire [4-1:0] node45755;
	wire [4-1:0] node45756;
	wire [4-1:0] node45757;
	wire [4-1:0] node45760;
	wire [4-1:0] node45763;
	wire [4-1:0] node45764;
	wire [4-1:0] node45765;
	wire [4-1:0] node45768;
	wire [4-1:0] node45771;
	wire [4-1:0] node45772;
	wire [4-1:0] node45775;
	wire [4-1:0] node45778;
	wire [4-1:0] node45779;
	wire [4-1:0] node45780;
	wire [4-1:0] node45782;
	wire [4-1:0] node45785;
	wire [4-1:0] node45786;
	wire [4-1:0] node45788;
	wire [4-1:0] node45791;
	wire [4-1:0] node45793;
	wire [4-1:0] node45796;
	wire [4-1:0] node45797;
	wire [4-1:0] node45798;
	wire [4-1:0] node45799;
	wire [4-1:0] node45802;
	wire [4-1:0] node45806;
	wire [4-1:0] node45808;
	wire [4-1:0] node45809;
	wire [4-1:0] node45812;
	wire [4-1:0] node45815;
	wire [4-1:0] node45816;
	wire [4-1:0] node45817;
	wire [4-1:0] node45818;
	wire [4-1:0] node45821;
	wire [4-1:0] node45824;
	wire [4-1:0] node45826;
	wire [4-1:0] node45827;
	wire [4-1:0] node45830;
	wire [4-1:0] node45833;
	wire [4-1:0] node45834;
	wire [4-1:0] node45835;
	wire [4-1:0] node45836;
	wire [4-1:0] node45837;
	wire [4-1:0] node45841;
	wire [4-1:0] node45844;
	wire [4-1:0] node45845;
	wire [4-1:0] node45849;
	wire [4-1:0] node45850;
	wire [4-1:0] node45851;
	wire [4-1:0] node45854;
	wire [4-1:0] node45858;
	wire [4-1:0] node45859;
	wire [4-1:0] node45860;
	wire [4-1:0] node45861;
	wire [4-1:0] node45862;
	wire [4-1:0] node45864;
	wire [4-1:0] node45867;
	wire [4-1:0] node45868;
	wire [4-1:0] node45869;
	wire [4-1:0] node45872;
	wire [4-1:0] node45875;
	wire [4-1:0] node45876;
	wire [4-1:0] node45879;
	wire [4-1:0] node45882;
	wire [4-1:0] node45883;
	wire [4-1:0] node45884;
	wire [4-1:0] node45886;
	wire [4-1:0] node45889;
	wire [4-1:0] node45890;
	wire [4-1:0] node45894;
	wire [4-1:0] node45896;
	wire [4-1:0] node45899;
	wire [4-1:0] node45900;
	wire [4-1:0] node45901;
	wire [4-1:0] node45903;
	wire [4-1:0] node45906;
	wire [4-1:0] node45908;
	wire [4-1:0] node45911;
	wire [4-1:0] node45912;
	wire [4-1:0] node45913;
	wire [4-1:0] node45914;
	wire [4-1:0] node45917;
	wire [4-1:0] node45920;
	wire [4-1:0] node45921;
	wire [4-1:0] node45924;
	wire [4-1:0] node45927;
	wire [4-1:0] node45929;
	wire [4-1:0] node45930;
	wire [4-1:0] node45933;
	wire [4-1:0] node45936;
	wire [4-1:0] node45937;
	wire [4-1:0] node45938;
	wire [4-1:0] node45940;
	wire [4-1:0] node45942;
	wire [4-1:0] node45945;
	wire [4-1:0] node45946;
	wire [4-1:0] node45947;
	wire [4-1:0] node45950;
	wire [4-1:0] node45953;
	wire [4-1:0] node45955;
	wire [4-1:0] node45956;
	wire [4-1:0] node45959;
	wire [4-1:0] node45962;
	wire [4-1:0] node45963;
	wire [4-1:0] node45964;
	wire [4-1:0] node45965;
	wire [4-1:0] node45967;
	wire [4-1:0] node45970;
	wire [4-1:0] node45972;
	wire [4-1:0] node45976;
	wire [4-1:0] node45978;
	wire [4-1:0] node45979;
	wire [4-1:0] node45983;
	wire [4-1:0] node45984;
	wire [4-1:0] node45985;
	wire [4-1:0] node45986;
	wire [4-1:0] node45987;
	wire [4-1:0] node45988;
	wire [4-1:0] node45991;
	wire [4-1:0] node45993;
	wire [4-1:0] node45996;
	wire [4-1:0] node45998;
	wire [4-1:0] node45999;
	wire [4-1:0] node46003;
	wire [4-1:0] node46004;
	wire [4-1:0] node46005;
	wire [4-1:0] node46007;
	wire [4-1:0] node46011;
	wire [4-1:0] node46012;
	wire [4-1:0] node46014;
	wire [4-1:0] node46017;
	wire [4-1:0] node46019;
	wire [4-1:0] node46022;
	wire [4-1:0] node46023;
	wire [4-1:0] node46024;
	wire [4-1:0] node46025;
	wire [4-1:0] node46028;
	wire [4-1:0] node46031;
	wire [4-1:0] node46032;
	wire [4-1:0] node46033;
	wire [4-1:0] node46036;
	wire [4-1:0] node46039;
	wire [4-1:0] node46041;
	wire [4-1:0] node46044;
	wire [4-1:0] node46045;
	wire [4-1:0] node46047;
	wire [4-1:0] node46049;
	wire [4-1:0] node46050;
	wire [4-1:0] node46053;
	wire [4-1:0] node46056;
	wire [4-1:0] node46057;
	wire [4-1:0] node46061;
	wire [4-1:0] node46062;
	wire [4-1:0] node46063;
	wire [4-1:0] node46064;
	wire [4-1:0] node46065;
	wire [4-1:0] node46068;
	wire [4-1:0] node46071;
	wire [4-1:0] node46072;
	wire [4-1:0] node46075;
	wire [4-1:0] node46078;
	wire [4-1:0] node46079;
	wire [4-1:0] node46080;
	wire [4-1:0] node46082;
	wire [4-1:0] node46085;
	wire [4-1:0] node46086;
	wire [4-1:0] node46089;
	wire [4-1:0] node46092;
	wire [4-1:0] node46093;
	wire [4-1:0] node46094;
	wire [4-1:0] node46098;
	wire [4-1:0] node46100;
	wire [4-1:0] node46103;
	wire [4-1:0] node46104;
	wire [4-1:0] node46105;
	wire [4-1:0] node46106;
	wire [4-1:0] node46107;
	wire [4-1:0] node46109;
	wire [4-1:0] node46112;
	wire [4-1:0] node46113;
	wire [4-1:0] node46116;
	wire [4-1:0] node46119;
	wire [4-1:0] node46120;
	wire [4-1:0] node46122;
	wire [4-1:0] node46126;
	wire [4-1:0] node46127;
	wire [4-1:0] node46129;
	wire [4-1:0] node46132;
	wire [4-1:0] node46133;
	wire [4-1:0] node46136;
	wire [4-1:0] node46139;
	wire [4-1:0] node46140;
	wire [4-1:0] node46141;
	wire [4-1:0] node46142;
	wire [4-1:0] node46145;
	wire [4-1:0] node46148;
	wire [4-1:0] node46149;
	wire [4-1:0] node46150;
	wire [4-1:0] node46153;
	wire [4-1:0] node46157;
	wire [4-1:0] node46158;
	wire [4-1:0] node46161;
	wire [4-1:0] node46162;
	wire [4-1:0] node46164;
	wire [4-1:0] node46167;
	wire [4-1:0] node46170;
	wire [4-1:0] node46171;
	wire [4-1:0] node46172;
	wire [4-1:0] node46173;
	wire [4-1:0] node46174;
	wire [4-1:0] node46175;
	wire [4-1:0] node46176;
	wire [4-1:0] node46177;
	wire [4-1:0] node46180;
	wire [4-1:0] node46183;
	wire [4-1:0] node46184;
	wire [4-1:0] node46187;
	wire [4-1:0] node46190;
	wire [4-1:0] node46191;
	wire [4-1:0] node46192;
	wire [4-1:0] node46195;
	wire [4-1:0] node46198;
	wire [4-1:0] node46199;
	wire [4-1:0] node46202;
	wire [4-1:0] node46205;
	wire [4-1:0] node46206;
	wire [4-1:0] node46207;
	wire [4-1:0] node46208;
	wire [4-1:0] node46209;
	wire [4-1:0] node46212;
	wire [4-1:0] node46215;
	wire [4-1:0] node46218;
	wire [4-1:0] node46219;
	wire [4-1:0] node46221;
	wire [4-1:0] node46225;
	wire [4-1:0] node46226;
	wire [4-1:0] node46227;
	wire [4-1:0] node46229;
	wire [4-1:0] node46232;
	wire [4-1:0] node46233;
	wire [4-1:0] node46237;
	wire [4-1:0] node46238;
	wire [4-1:0] node46239;
	wire [4-1:0] node46242;
	wire [4-1:0] node46245;
	wire [4-1:0] node46247;
	wire [4-1:0] node46250;
	wire [4-1:0] node46251;
	wire [4-1:0] node46252;
	wire [4-1:0] node46253;
	wire [4-1:0] node46254;
	wire [4-1:0] node46257;
	wire [4-1:0] node46260;
	wire [4-1:0] node46261;
	wire [4-1:0] node46264;
	wire [4-1:0] node46267;
	wire [4-1:0] node46268;
	wire [4-1:0] node46269;
	wire [4-1:0] node46272;
	wire [4-1:0] node46275;
	wire [4-1:0] node46276;
	wire [4-1:0] node46277;
	wire [4-1:0] node46281;
	wire [4-1:0] node46283;
	wire [4-1:0] node46286;
	wire [4-1:0] node46287;
	wire [4-1:0] node46288;
	wire [4-1:0] node46289;
	wire [4-1:0] node46290;
	wire [4-1:0] node46294;
	wire [4-1:0] node46296;
	wire [4-1:0] node46299;
	wire [4-1:0] node46300;
	wire [4-1:0] node46304;
	wire [4-1:0] node46305;
	wire [4-1:0] node46306;
	wire [4-1:0] node46307;
	wire [4-1:0] node46311;
	wire [4-1:0] node46312;
	wire [4-1:0] node46316;
	wire [4-1:0] node46317;
	wire [4-1:0] node46318;
	wire [4-1:0] node46321;
	wire [4-1:0] node46324;
	wire [4-1:0] node46325;
	wire [4-1:0] node46328;
	wire [4-1:0] node46331;
	wire [4-1:0] node46332;
	wire [4-1:0] node46333;
	wire [4-1:0] node46334;
	wire [4-1:0] node46335;
	wire [4-1:0] node46336;
	wire [4-1:0] node46340;
	wire [4-1:0] node46341;
	wire [4-1:0] node46344;
	wire [4-1:0] node46347;
	wire [4-1:0] node46348;
	wire [4-1:0] node46349;
	wire [4-1:0] node46352;
	wire [4-1:0] node46356;
	wire [4-1:0] node46357;
	wire [4-1:0] node46358;
	wire [4-1:0] node46359;
	wire [4-1:0] node46360;
	wire [4-1:0] node46363;
	wire [4-1:0] node46367;
	wire [4-1:0] node46368;
	wire [4-1:0] node46369;
	wire [4-1:0] node46374;
	wire [4-1:0] node46375;
	wire [4-1:0] node46376;
	wire [4-1:0] node46380;
	wire [4-1:0] node46381;
	wire [4-1:0] node46384;
	wire [4-1:0] node46387;
	wire [4-1:0] node46388;
	wire [4-1:0] node46389;
	wire [4-1:0] node46390;
	wire [4-1:0] node46391;
	wire [4-1:0] node46393;
	wire [4-1:0] node46397;
	wire [4-1:0] node46398;
	wire [4-1:0] node46399;
	wire [4-1:0] node46404;
	wire [4-1:0] node46405;
	wire [4-1:0] node46407;
	wire [4-1:0] node46409;
	wire [4-1:0] node46412;
	wire [4-1:0] node46413;
	wire [4-1:0] node46415;
	wire [4-1:0] node46418;
	wire [4-1:0] node46419;
	wire [4-1:0] node46422;
	wire [4-1:0] node46425;
	wire [4-1:0] node46426;
	wire [4-1:0] node46427;
	wire [4-1:0] node46430;
	wire [4-1:0] node46433;
	wire [4-1:0] node46434;
	wire [4-1:0] node46435;
	wire [4-1:0] node46439;
	wire [4-1:0] node46440;
	wire [4-1:0] node46443;
	wire [4-1:0] node46446;
	wire [4-1:0] node46447;
	wire [4-1:0] node46448;
	wire [4-1:0] node46449;
	wire [4-1:0] node46450;
	wire [4-1:0] node46451;
	wire [4-1:0] node46455;
	wire [4-1:0] node46456;
	wire [4-1:0] node46460;
	wire [4-1:0] node46461;
	wire [4-1:0] node46462;
	wire [4-1:0] node46466;
	wire [4-1:0] node46467;
	wire [4-1:0] node46471;
	wire [4-1:0] node46472;
	wire [4-1:0] node46473;
	wire [4-1:0] node46474;
	wire [4-1:0] node46477;
	wire [4-1:0] node46478;
	wire [4-1:0] node46482;
	wire [4-1:0] node46483;
	wire [4-1:0] node46486;
	wire [4-1:0] node46487;
	wire [4-1:0] node46491;
	wire [4-1:0] node46492;
	wire [4-1:0] node46493;
	wire [4-1:0] node46494;
	wire [4-1:0] node46498;
	wire [4-1:0] node46499;
	wire [4-1:0] node46503;
	wire [4-1:0] node46504;
	wire [4-1:0] node46505;
	wire [4-1:0] node46506;
	wire [4-1:0] node46510;
	wire [4-1:0] node46511;
	wire [4-1:0] node46514;
	wire [4-1:0] node46518;
	wire [4-1:0] node46519;
	wire [4-1:0] node46520;
	wire [4-1:0] node46521;
	wire [4-1:0] node46522;
	wire [4-1:0] node46523;
	wire [4-1:0] node46527;
	wire [4-1:0] node46528;
	wire [4-1:0] node46532;
	wire [4-1:0] node46533;
	wire [4-1:0] node46536;
	wire [4-1:0] node46539;
	wire [4-1:0] node46540;
	wire [4-1:0] node46541;
	wire [4-1:0] node46542;
	wire [4-1:0] node46543;
	wire [4-1:0] node46546;
	wire [4-1:0] node46549;
	wire [4-1:0] node46550;
	wire [4-1:0] node46554;
	wire [4-1:0] node46555;
	wire [4-1:0] node46556;
	wire [4-1:0] node46559;
	wire [4-1:0] node46562;
	wire [4-1:0] node46563;
	wire [4-1:0] node46566;
	wire [4-1:0] node46569;
	wire [4-1:0] node46570;
	wire [4-1:0] node46573;
	wire [4-1:0] node46576;
	wire [4-1:0] node46577;
	wire [4-1:0] node46578;
	wire [4-1:0] node46579;
	wire [4-1:0] node46580;
	wire [4-1:0] node46584;
	wire [4-1:0] node46585;
	wire [4-1:0] node46589;
	wire [4-1:0] node46590;
	wire [4-1:0] node46591;
	wire [4-1:0] node46596;
	wire [4-1:0] node46597;
	wire [4-1:0] node46599;
	wire [4-1:0] node46600;
	wire [4-1:0] node46603;
	wire [4-1:0] node46606;
	wire [4-1:0] node46608;
	wire [4-1:0] node46609;
	wire [4-1:0] node46613;
	wire [4-1:0] node46614;
	wire [4-1:0] node46615;
	wire [4-1:0] node46616;
	wire [4-1:0] node46617;
	wire [4-1:0] node46618;
	wire [4-1:0] node46619;
	wire [4-1:0] node46620;
	wire [4-1:0] node46624;
	wire [4-1:0] node46625;
	wire [4-1:0] node46626;
	wire [4-1:0] node46627;
	wire [4-1:0] node46631;
	wire [4-1:0] node46633;
	wire [4-1:0] node46636;
	wire [4-1:0] node46637;
	wire [4-1:0] node46638;
	wire [4-1:0] node46643;
	wire [4-1:0] node46644;
	wire [4-1:0] node46645;
	wire [4-1:0] node46646;
	wire [4-1:0] node46647;
	wire [4-1:0] node46652;
	wire [4-1:0] node46653;
	wire [4-1:0] node46654;
	wire [4-1:0] node46657;
	wire [4-1:0] node46660;
	wire [4-1:0] node46661;
	wire [4-1:0] node46665;
	wire [4-1:0] node46666;
	wire [4-1:0] node46669;
	wire [4-1:0] node46670;
	wire [4-1:0] node46671;
	wire [4-1:0] node46676;
	wire [4-1:0] node46677;
	wire [4-1:0] node46678;
	wire [4-1:0] node46679;
	wire [4-1:0] node46680;
	wire [4-1:0] node46683;
	wire [4-1:0] node46686;
	wire [4-1:0] node46687;
	wire [4-1:0] node46690;
	wire [4-1:0] node46693;
	wire [4-1:0] node46694;
	wire [4-1:0] node46695;
	wire [4-1:0] node46698;
	wire [4-1:0] node46701;
	wire [4-1:0] node46703;
	wire [4-1:0] node46706;
	wire [4-1:0] node46707;
	wire [4-1:0] node46709;
	wire [4-1:0] node46710;
	wire [4-1:0] node46713;
	wire [4-1:0] node46716;
	wire [4-1:0] node46717;
	wire [4-1:0] node46718;
	wire [4-1:0] node46719;
	wire [4-1:0] node46722;
	wire [4-1:0] node46725;
	wire [4-1:0] node46726;
	wire [4-1:0] node46729;
	wire [4-1:0] node46732;
	wire [4-1:0] node46733;
	wire [4-1:0] node46736;
	wire [4-1:0] node46739;
	wire [4-1:0] node46740;
	wire [4-1:0] node46741;
	wire [4-1:0] node46742;
	wire [4-1:0] node46743;
	wire [4-1:0] node46744;
	wire [4-1:0] node46748;
	wire [4-1:0] node46749;
	wire [4-1:0] node46753;
	wire [4-1:0] node46754;
	wire [4-1:0] node46755;
	wire [4-1:0] node46759;
	wire [4-1:0] node46760;
	wire [4-1:0] node46764;
	wire [4-1:0] node46765;
	wire [4-1:0] node46766;
	wire [4-1:0] node46768;
	wire [4-1:0] node46769;
	wire [4-1:0] node46772;
	wire [4-1:0] node46775;
	wire [4-1:0] node46777;
	wire [4-1:0] node46780;
	wire [4-1:0] node46781;
	wire [4-1:0] node46783;
	wire [4-1:0] node46786;
	wire [4-1:0] node46787;
	wire [4-1:0] node46791;
	wire [4-1:0] node46792;
	wire [4-1:0] node46793;
	wire [4-1:0] node46794;
	wire [4-1:0] node46797;
	wire [4-1:0] node46800;
	wire [4-1:0] node46801;
	wire [4-1:0] node46802;
	wire [4-1:0] node46806;
	wire [4-1:0] node46807;
	wire [4-1:0] node46811;
	wire [4-1:0] node46812;
	wire [4-1:0] node46813;
	wire [4-1:0] node46814;
	wire [4-1:0] node46815;
	wire [4-1:0] node46819;
	wire [4-1:0] node46821;
	wire [4-1:0] node46824;
	wire [4-1:0] node46825;
	wire [4-1:0] node46829;
	wire [4-1:0] node46830;
	wire [4-1:0] node46833;
	wire [4-1:0] node46836;
	wire [4-1:0] node46837;
	wire [4-1:0] node46838;
	wire [4-1:0] node46839;
	wire [4-1:0] node46840;
	wire [4-1:0] node46841;
	wire [4-1:0] node46842;
	wire [4-1:0] node46845;
	wire [4-1:0] node46848;
	wire [4-1:0] node46851;
	wire [4-1:0] node46852;
	wire [4-1:0] node46854;
	wire [4-1:0] node46857;
	wire [4-1:0] node46858;
	wire [4-1:0] node46861;
	wire [4-1:0] node46864;
	wire [4-1:0] node46865;
	wire [4-1:0] node46866;
	wire [4-1:0] node46867;
	wire [4-1:0] node46868;
	wire [4-1:0] node46871;
	wire [4-1:0] node46874;
	wire [4-1:0] node46875;
	wire [4-1:0] node46878;
	wire [4-1:0] node46881;
	wire [4-1:0] node46883;
	wire [4-1:0] node46884;
	wire [4-1:0] node46887;
	wire [4-1:0] node46890;
	wire [4-1:0] node46891;
	wire [4-1:0] node46892;
	wire [4-1:0] node46894;
	wire [4-1:0] node46897;
	wire [4-1:0] node46898;
	wire [4-1:0] node46903;
	wire [4-1:0] node46904;
	wire [4-1:0] node46905;
	wire [4-1:0] node46906;
	wire [4-1:0] node46907;
	wire [4-1:0] node46908;
	wire [4-1:0] node46911;
	wire [4-1:0] node46914;
	wire [4-1:0] node46916;
	wire [4-1:0] node46919;
	wire [4-1:0] node46920;
	wire [4-1:0] node46922;
	wire [4-1:0] node46925;
	wire [4-1:0] node46927;
	wire [4-1:0] node46930;
	wire [4-1:0] node46931;
	wire [4-1:0] node46933;
	wire [4-1:0] node46934;
	wire [4-1:0] node46938;
	wire [4-1:0] node46939;
	wire [4-1:0] node46940;
	wire [4-1:0] node46944;
	wire [4-1:0] node46947;
	wire [4-1:0] node46948;
	wire [4-1:0] node46949;
	wire [4-1:0] node46950;
	wire [4-1:0] node46954;
	wire [4-1:0] node46955;
	wire [4-1:0] node46956;
	wire [4-1:0] node46959;
	wire [4-1:0] node46963;
	wire [4-1:0] node46964;
	wire [4-1:0] node46967;
	wire [4-1:0] node46970;
	wire [4-1:0] node46971;
	wire [4-1:0] node46972;
	wire [4-1:0] node46973;
	wire [4-1:0] node46974;
	wire [4-1:0] node46977;
	wire [4-1:0] node46979;
	wire [4-1:0] node46982;
	wire [4-1:0] node46983;
	wire [4-1:0] node46984;
	wire [4-1:0] node46986;
	wire [4-1:0] node46990;
	wire [4-1:0] node46991;
	wire [4-1:0] node46994;
	wire [4-1:0] node46997;
	wire [4-1:0] node46998;
	wire [4-1:0] node46999;
	wire [4-1:0] node47000;
	wire [4-1:0] node47003;
	wire [4-1:0] node47007;
	wire [4-1:0] node47008;
	wire [4-1:0] node47011;
	wire [4-1:0] node47014;
	wire [4-1:0] node47015;
	wire [4-1:0] node47016;
	wire [4-1:0] node47017;
	wire [4-1:0] node47018;
	wire [4-1:0] node47020;
	wire [4-1:0] node47023;
	wire [4-1:0] node47026;
	wire [4-1:0] node47027;
	wire [4-1:0] node47028;
	wire [4-1:0] node47032;
	wire [4-1:0] node47033;
	wire [4-1:0] node47037;
	wire [4-1:0] node47038;
	wire [4-1:0] node47039;
	wire [4-1:0] node47042;
	wire [4-1:0] node47046;
	wire [4-1:0] node47047;
	wire [4-1:0] node47048;
	wire [4-1:0] node47049;
	wire [4-1:0] node47053;
	wire [4-1:0] node47054;
	wire [4-1:0] node47055;
	wire [4-1:0] node47060;
	wire [4-1:0] node47061;
	wire [4-1:0] node47062;
	wire [4-1:0] node47063;
	wire [4-1:0] node47066;
	wire [4-1:0] node47071;
	wire [4-1:0] node47072;
	wire [4-1:0] node47073;
	wire [4-1:0] node47074;
	wire [4-1:0] node47075;
	wire [4-1:0] node47076;
	wire [4-1:0] node47077;
	wire [4-1:0] node47078;
	wire [4-1:0] node47081;
	wire [4-1:0] node47084;
	wire [4-1:0] node47085;
	wire [4-1:0] node47089;
	wire [4-1:0] node47090;
	wire [4-1:0] node47093;
	wire [4-1:0] node47094;
	wire [4-1:0] node47095;
	wire [4-1:0] node47100;
	wire [4-1:0] node47101;
	wire [4-1:0] node47102;
	wire [4-1:0] node47103;
	wire [4-1:0] node47107;
	wire [4-1:0] node47108;
	wire [4-1:0] node47111;
	wire [4-1:0] node47114;
	wire [4-1:0] node47115;
	wire [4-1:0] node47118;
	wire [4-1:0] node47121;
	wire [4-1:0] node47122;
	wire [4-1:0] node47123;
	wire [4-1:0] node47124;
	wire [4-1:0] node47125;
	wire [4-1:0] node47129;
	wire [4-1:0] node47130;
	wire [4-1:0] node47134;
	wire [4-1:0] node47135;
	wire [4-1:0] node47136;
	wire [4-1:0] node47140;
	wire [4-1:0] node47141;
	wire [4-1:0] node47145;
	wire [4-1:0] node47146;
	wire [4-1:0] node47147;
	wire [4-1:0] node47148;
	wire [4-1:0] node47149;
	wire [4-1:0] node47153;
	wire [4-1:0] node47156;
	wire [4-1:0] node47157;
	wire [4-1:0] node47160;
	wire [4-1:0] node47163;
	wire [4-1:0] node47164;
	wire [4-1:0] node47165;
	wire [4-1:0] node47167;
	wire [4-1:0] node47172;
	wire [4-1:0] node47173;
	wire [4-1:0] node47174;
	wire [4-1:0] node47175;
	wire [4-1:0] node47176;
	wire [4-1:0] node47177;
	wire [4-1:0] node47180;
	wire [4-1:0] node47183;
	wire [4-1:0] node47184;
	wire [4-1:0] node47187;
	wire [4-1:0] node47190;
	wire [4-1:0] node47191;
	wire [4-1:0] node47194;
	wire [4-1:0] node47197;
	wire [4-1:0] node47198;
	wire [4-1:0] node47199;
	wire [4-1:0] node47200;
	wire [4-1:0] node47201;
	wire [4-1:0] node47205;
	wire [4-1:0] node47208;
	wire [4-1:0] node47209;
	wire [4-1:0] node47212;
	wire [4-1:0] node47215;
	wire [4-1:0] node47216;
	wire [4-1:0] node47219;
	wire [4-1:0] node47222;
	wire [4-1:0] node47223;
	wire [4-1:0] node47224;
	wire [4-1:0] node47225;
	wire [4-1:0] node47228;
	wire [4-1:0] node47230;
	wire [4-1:0] node47233;
	wire [4-1:0] node47234;
	wire [4-1:0] node47237;
	wire [4-1:0] node47240;
	wire [4-1:0] node47241;
	wire [4-1:0] node47242;
	wire [4-1:0] node47243;
	wire [4-1:0] node47246;
	wire [4-1:0] node47249;
	wire [4-1:0] node47251;
	wire [4-1:0] node47254;
	wire [4-1:0] node47255;
	wire [4-1:0] node47258;
	wire [4-1:0] node47261;
	wire [4-1:0] node47262;
	wire [4-1:0] node47263;
	wire [4-1:0] node47264;
	wire [4-1:0] node47265;
	wire [4-1:0] node47266;
	wire [4-1:0] node47267;
	wire [4-1:0] node47270;
	wire [4-1:0] node47273;
	wire [4-1:0] node47274;
	wire [4-1:0] node47278;
	wire [4-1:0] node47279;
	wire [4-1:0] node47280;
	wire [4-1:0] node47281;
	wire [4-1:0] node47284;
	wire [4-1:0] node47287;
	wire [4-1:0] node47288;
	wire [4-1:0] node47291;
	wire [4-1:0] node47295;
	wire [4-1:0] node47296;
	wire [4-1:0] node47297;
	wire [4-1:0] node47298;
	wire [4-1:0] node47302;
	wire [4-1:0] node47303;
	wire [4-1:0] node47307;
	wire [4-1:0] node47309;
	wire [4-1:0] node47312;
	wire [4-1:0] node47313;
	wire [4-1:0] node47314;
	wire [4-1:0] node47315;
	wire [4-1:0] node47317;
	wire [4-1:0] node47321;
	wire [4-1:0] node47322;
	wire [4-1:0] node47323;
	wire [4-1:0] node47326;
	wire [4-1:0] node47329;
	wire [4-1:0] node47330;
	wire [4-1:0] node47331;
	wire [4-1:0] node47334;
	wire [4-1:0] node47338;
	wire [4-1:0] node47339;
	wire [4-1:0] node47340;
	wire [4-1:0] node47341;
	wire [4-1:0] node47343;
	wire [4-1:0] node47346;
	wire [4-1:0] node47347;
	wire [4-1:0] node47351;
	wire [4-1:0] node47352;
	wire [4-1:0] node47355;
	wire [4-1:0] node47358;
	wire [4-1:0] node47359;
	wire [4-1:0] node47360;
	wire [4-1:0] node47361;
	wire [4-1:0] node47364;
	wire [4-1:0] node47368;
	wire [4-1:0] node47369;
	wire [4-1:0] node47370;
	wire [4-1:0] node47375;
	wire [4-1:0] node47376;
	wire [4-1:0] node47377;
	wire [4-1:0] node47378;
	wire [4-1:0] node47379;
	wire [4-1:0] node47383;
	wire [4-1:0] node47384;
	wire [4-1:0] node47388;
	wire [4-1:0] node47389;
	wire [4-1:0] node47390;
	wire [4-1:0] node47393;
	wire [4-1:0] node47397;
	wire [4-1:0] node47398;
	wire [4-1:0] node47399;
	wire [4-1:0] node47400;
	wire [4-1:0] node47404;
	wire [4-1:0] node47405;
	wire [4-1:0] node47409;
	wire [4-1:0] node47410;
	wire [4-1:0] node47411;
	wire [4-1:0] node47415;
	wire [4-1:0] node47416;
	wire [4-1:0] node47420;
	wire [4-1:0] node47421;
	wire [4-1:0] node47422;
	wire [4-1:0] node47423;
	wire [4-1:0] node47424;
	wire [4-1:0] node47425;
	wire [4-1:0] node47426;
	wire [4-1:0] node47427;
	wire [4-1:0] node47428;
	wire [4-1:0] node47429;
	wire [4-1:0] node47430;
	wire [4-1:0] node47431;
	wire [4-1:0] node47432;
	wire [4-1:0] node47435;
	wire [4-1:0] node47438;
	wire [4-1:0] node47439;
	wire [4-1:0] node47440;
	wire [4-1:0] node47443;
	wire [4-1:0] node47447;
	wire [4-1:0] node47448;
	wire [4-1:0] node47451;
	wire [4-1:0] node47452;
	wire [4-1:0] node47456;
	wire [4-1:0] node47457;
	wire [4-1:0] node47458;
	wire [4-1:0] node47460;
	wire [4-1:0] node47463;
	wire [4-1:0] node47465;
	wire [4-1:0] node47467;
	wire [4-1:0] node47470;
	wire [4-1:0] node47471;
	wire [4-1:0] node47473;
	wire [4-1:0] node47474;
	wire [4-1:0] node47478;
	wire [4-1:0] node47481;
	wire [4-1:0] node47482;
	wire [4-1:0] node47483;
	wire [4-1:0] node47484;
	wire [4-1:0] node47485;
	wire [4-1:0] node47486;
	wire [4-1:0] node47491;
	wire [4-1:0] node47492;
	wire [4-1:0] node47493;
	wire [4-1:0] node47497;
	wire [4-1:0] node47498;
	wire [4-1:0] node47501;
	wire [4-1:0] node47504;
	wire [4-1:0] node47505;
	wire [4-1:0] node47506;
	wire [4-1:0] node47507;
	wire [4-1:0] node47511;
	wire [4-1:0] node47514;
	wire [4-1:0] node47515;
	wire [4-1:0] node47519;
	wire [4-1:0] node47520;
	wire [4-1:0] node47521;
	wire [4-1:0] node47522;
	wire [4-1:0] node47523;
	wire [4-1:0] node47527;
	wire [4-1:0] node47528;
	wire [4-1:0] node47532;
	wire [4-1:0] node47533;
	wire [4-1:0] node47535;
	wire [4-1:0] node47538;
	wire [4-1:0] node47539;
	wire [4-1:0] node47543;
	wire [4-1:0] node47544;
	wire [4-1:0] node47545;
	wire [4-1:0] node47548;
	wire [4-1:0] node47549;
	wire [4-1:0] node47553;
	wire [4-1:0] node47554;
	wire [4-1:0] node47555;
	wire [4-1:0] node47559;
	wire [4-1:0] node47562;
	wire [4-1:0] node47563;
	wire [4-1:0] node47564;
	wire [4-1:0] node47565;
	wire [4-1:0] node47566;
	wire [4-1:0] node47567;
	wire [4-1:0] node47570;
	wire [4-1:0] node47573;
	wire [4-1:0] node47574;
	wire [4-1:0] node47577;
	wire [4-1:0] node47580;
	wire [4-1:0] node47581;
	wire [4-1:0] node47582;
	wire [4-1:0] node47584;
	wire [4-1:0] node47587;
	wire [4-1:0] node47588;
	wire [4-1:0] node47591;
	wire [4-1:0] node47594;
	wire [4-1:0] node47595;
	wire [4-1:0] node47599;
	wire [4-1:0] node47600;
	wire [4-1:0] node47601;
	wire [4-1:0] node47604;
	wire [4-1:0] node47606;
	wire [4-1:0] node47608;
	wire [4-1:0] node47611;
	wire [4-1:0] node47612;
	wire [4-1:0] node47613;
	wire [4-1:0] node47614;
	wire [4-1:0] node47617;
	wire [4-1:0] node47621;
	wire [4-1:0] node47622;
	wire [4-1:0] node47626;
	wire [4-1:0] node47627;
	wire [4-1:0] node47628;
	wire [4-1:0] node47629;
	wire [4-1:0] node47632;
	wire [4-1:0] node47633;
	wire [4-1:0] node47636;
	wire [4-1:0] node47639;
	wire [4-1:0] node47640;
	wire [4-1:0] node47641;
	wire [4-1:0] node47643;
	wire [4-1:0] node47647;
	wire [4-1:0] node47648;
	wire [4-1:0] node47652;
	wire [4-1:0] node47653;
	wire [4-1:0] node47654;
	wire [4-1:0] node47655;
	wire [4-1:0] node47658;
	wire [4-1:0] node47659;
	wire [4-1:0] node47663;
	wire [4-1:0] node47665;
	wire [4-1:0] node47666;
	wire [4-1:0] node47670;
	wire [4-1:0] node47671;
	wire [4-1:0] node47673;
	wire [4-1:0] node47676;
	wire [4-1:0] node47677;
	wire [4-1:0] node47678;
	wire [4-1:0] node47682;
	wire [4-1:0] node47685;
	wire [4-1:0] node47686;
	wire [4-1:0] node47687;
	wire [4-1:0] node47688;
	wire [4-1:0] node47689;
	wire [4-1:0] node47690;
	wire [4-1:0] node47691;
	wire [4-1:0] node47695;
	wire [4-1:0] node47696;
	wire [4-1:0] node47697;
	wire [4-1:0] node47700;
	wire [4-1:0] node47704;
	wire [4-1:0] node47706;
	wire [4-1:0] node47707;
	wire [4-1:0] node47710;
	wire [4-1:0] node47713;
	wire [4-1:0] node47714;
	wire [4-1:0] node47715;
	wire [4-1:0] node47716;
	wire [4-1:0] node47718;
	wire [4-1:0] node47721;
	wire [4-1:0] node47722;
	wire [4-1:0] node47725;
	wire [4-1:0] node47728;
	wire [4-1:0] node47729;
	wire [4-1:0] node47730;
	wire [4-1:0] node47733;
	wire [4-1:0] node47736;
	wire [4-1:0] node47738;
	wire [4-1:0] node47741;
	wire [4-1:0] node47742;
	wire [4-1:0] node47743;
	wire [4-1:0] node47747;
	wire [4-1:0] node47749;
	wire [4-1:0] node47752;
	wire [4-1:0] node47753;
	wire [4-1:0] node47754;
	wire [4-1:0] node47755;
	wire [4-1:0] node47756;
	wire [4-1:0] node47760;
	wire [4-1:0] node47761;
	wire [4-1:0] node47764;
	wire [4-1:0] node47767;
	wire [4-1:0] node47768;
	wire [4-1:0] node47769;
	wire [4-1:0] node47773;
	wire [4-1:0] node47774;
	wire [4-1:0] node47776;
	wire [4-1:0] node47779;
	wire [4-1:0] node47780;
	wire [4-1:0] node47784;
	wire [4-1:0] node47785;
	wire [4-1:0] node47786;
	wire [4-1:0] node47788;
	wire [4-1:0] node47791;
	wire [4-1:0] node47792;
	wire [4-1:0] node47795;
	wire [4-1:0] node47798;
	wire [4-1:0] node47799;
	wire [4-1:0] node47800;
	wire [4-1:0] node47803;
	wire [4-1:0] node47806;
	wire [4-1:0] node47807;
	wire [4-1:0] node47811;
	wire [4-1:0] node47812;
	wire [4-1:0] node47813;
	wire [4-1:0] node47814;
	wire [4-1:0] node47815;
	wire [4-1:0] node47816;
	wire [4-1:0] node47818;
	wire [4-1:0] node47821;
	wire [4-1:0] node47824;
	wire [4-1:0] node47825;
	wire [4-1:0] node47829;
	wire [4-1:0] node47830;
	wire [4-1:0] node47831;
	wire [4-1:0] node47834;
	wire [4-1:0] node47837;
	wire [4-1:0] node47839;
	wire [4-1:0] node47842;
	wire [4-1:0] node47843;
	wire [4-1:0] node47844;
	wire [4-1:0] node47846;
	wire [4-1:0] node47849;
	wire [4-1:0] node47850;
	wire [4-1:0] node47853;
	wire [4-1:0] node47855;
	wire [4-1:0] node47858;
	wire [4-1:0] node47859;
	wire [4-1:0] node47860;
	wire [4-1:0] node47863;
	wire [4-1:0] node47866;
	wire [4-1:0] node47869;
	wire [4-1:0] node47870;
	wire [4-1:0] node47871;
	wire [4-1:0] node47872;
	wire [4-1:0] node47873;
	wire [4-1:0] node47876;
	wire [4-1:0] node47880;
	wire [4-1:0] node47881;
	wire [4-1:0] node47883;
	wire [4-1:0] node47886;
	wire [4-1:0] node47887;
	wire [4-1:0] node47889;
	wire [4-1:0] node47892;
	wire [4-1:0] node47895;
	wire [4-1:0] node47896;
	wire [4-1:0] node47897;
	wire [4-1:0] node47898;
	wire [4-1:0] node47899;
	wire [4-1:0] node47903;
	wire [4-1:0] node47907;
	wire [4-1:0] node47908;
	wire [4-1:0] node47909;
	wire [4-1:0] node47910;
	wire [4-1:0] node47913;
	wire [4-1:0] node47916;
	wire [4-1:0] node47918;
	wire [4-1:0] node47921;
	wire [4-1:0] node47922;
	wire [4-1:0] node47923;
	wire [4-1:0] node47927;
	wire [4-1:0] node47928;
	wire [4-1:0] node47931;
	wire [4-1:0] node47934;
	wire [4-1:0] node47935;
	wire [4-1:0] node47936;
	wire [4-1:0] node47937;
	wire [4-1:0] node47938;
	wire [4-1:0] node47939;
	wire [4-1:0] node47940;
	wire [4-1:0] node47942;
	wire [4-1:0] node47944;
	wire [4-1:0] node47947;
	wire [4-1:0] node47949;
	wire [4-1:0] node47950;
	wire [4-1:0] node47954;
	wire [4-1:0] node47955;
	wire [4-1:0] node47956;
	wire [4-1:0] node47960;
	wire [4-1:0] node47962;
	wire [4-1:0] node47964;
	wire [4-1:0] node47967;
	wire [4-1:0] node47968;
	wire [4-1:0] node47969;
	wire [4-1:0] node47970;
	wire [4-1:0] node47971;
	wire [4-1:0] node47975;
	wire [4-1:0] node47976;
	wire [4-1:0] node47979;
	wire [4-1:0] node47982;
	wire [4-1:0] node47983;
	wire [4-1:0] node47986;
	wire [4-1:0] node47988;
	wire [4-1:0] node47991;
	wire [4-1:0] node47992;
	wire [4-1:0] node47994;
	wire [4-1:0] node47996;
	wire [4-1:0] node47999;
	wire [4-1:0] node48000;
	wire [4-1:0] node48001;
	wire [4-1:0] node48004;
	wire [4-1:0] node48007;
	wire [4-1:0] node48008;
	wire [4-1:0] node48012;
	wire [4-1:0] node48013;
	wire [4-1:0] node48014;
	wire [4-1:0] node48015;
	wire [4-1:0] node48016;
	wire [4-1:0] node48017;
	wire [4-1:0] node48020;
	wire [4-1:0] node48023;
	wire [4-1:0] node48026;
	wire [4-1:0] node48028;
	wire [4-1:0] node48029;
	wire [4-1:0] node48032;
	wire [4-1:0] node48035;
	wire [4-1:0] node48036;
	wire [4-1:0] node48037;
	wire [4-1:0] node48038;
	wire [4-1:0] node48042;
	wire [4-1:0] node48043;
	wire [4-1:0] node48046;
	wire [4-1:0] node48049;
	wire [4-1:0] node48050;
	wire [4-1:0] node48051;
	wire [4-1:0] node48056;
	wire [4-1:0] node48057;
	wire [4-1:0] node48058;
	wire [4-1:0] node48059;
	wire [4-1:0] node48060;
	wire [4-1:0] node48064;
	wire [4-1:0] node48066;
	wire [4-1:0] node48069;
	wire [4-1:0] node48071;
	wire [4-1:0] node48074;
	wire [4-1:0] node48075;
	wire [4-1:0] node48077;
	wire [4-1:0] node48080;
	wire [4-1:0] node48082;
	wire [4-1:0] node48083;
	wire [4-1:0] node48086;
	wire [4-1:0] node48089;
	wire [4-1:0] node48090;
	wire [4-1:0] node48091;
	wire [4-1:0] node48092;
	wire [4-1:0] node48093;
	wire [4-1:0] node48094;
	wire [4-1:0] node48098;
	wire [4-1:0] node48099;
	wire [4-1:0] node48103;
	wire [4-1:0] node48104;
	wire [4-1:0] node48106;
	wire [4-1:0] node48107;
	wire [4-1:0] node48111;
	wire [4-1:0] node48112;
	wire [4-1:0] node48113;
	wire [4-1:0] node48117;
	wire [4-1:0] node48118;
	wire [4-1:0] node48122;
	wire [4-1:0] node48123;
	wire [4-1:0] node48124;
	wire [4-1:0] node48126;
	wire [4-1:0] node48127;
	wire [4-1:0] node48131;
	wire [4-1:0] node48132;
	wire [4-1:0] node48133;
	wire [4-1:0] node48136;
	wire [4-1:0] node48140;
	wire [4-1:0] node48141;
	wire [4-1:0] node48142;
	wire [4-1:0] node48145;
	wire [4-1:0] node48146;
	wire [4-1:0] node48151;
	wire [4-1:0] node48152;
	wire [4-1:0] node48153;
	wire [4-1:0] node48154;
	wire [4-1:0] node48155;
	wire [4-1:0] node48158;
	wire [4-1:0] node48161;
	wire [4-1:0] node48162;
	wire [4-1:0] node48165;
	wire [4-1:0] node48167;
	wire [4-1:0] node48170;
	wire [4-1:0] node48171;
	wire [4-1:0] node48172;
	wire [4-1:0] node48173;
	wire [4-1:0] node48176;
	wire [4-1:0] node48180;
	wire [4-1:0] node48181;
	wire [4-1:0] node48184;
	wire [4-1:0] node48187;
	wire [4-1:0] node48188;
	wire [4-1:0] node48189;
	wire [4-1:0] node48191;
	wire [4-1:0] node48194;
	wire [4-1:0] node48197;
	wire [4-1:0] node48198;
	wire [4-1:0] node48199;
	wire [4-1:0] node48202;
	wire [4-1:0] node48203;
	wire [4-1:0] node48206;
	wire [4-1:0] node48209;
	wire [4-1:0] node48211;
	wire [4-1:0] node48214;
	wire [4-1:0] node48215;
	wire [4-1:0] node48216;
	wire [4-1:0] node48217;
	wire [4-1:0] node48218;
	wire [4-1:0] node48219;
	wire [4-1:0] node48222;
	wire [4-1:0] node48225;
	wire [4-1:0] node48226;
	wire [4-1:0] node48228;
	wire [4-1:0] node48229;
	wire [4-1:0] node48233;
	wire [4-1:0] node48235;
	wire [4-1:0] node48238;
	wire [4-1:0] node48239;
	wire [4-1:0] node48241;
	wire [4-1:0] node48242;
	wire [4-1:0] node48246;
	wire [4-1:0] node48247;
	wire [4-1:0] node48248;
	wire [4-1:0] node48251;
	wire [4-1:0] node48254;
	wire [4-1:0] node48255;
	wire [4-1:0] node48259;
	wire [4-1:0] node48260;
	wire [4-1:0] node48261;
	wire [4-1:0] node48262;
	wire [4-1:0] node48264;
	wire [4-1:0] node48267;
	wire [4-1:0] node48268;
	wire [4-1:0] node48271;
	wire [4-1:0] node48274;
	wire [4-1:0] node48275;
	wire [4-1:0] node48277;
	wire [4-1:0] node48280;
	wire [4-1:0] node48281;
	wire [4-1:0] node48282;
	wire [4-1:0] node48286;
	wire [4-1:0] node48289;
	wire [4-1:0] node48290;
	wire [4-1:0] node48291;
	wire [4-1:0] node48292;
	wire [4-1:0] node48293;
	wire [4-1:0] node48296;
	wire [4-1:0] node48299;
	wire [4-1:0] node48300;
	wire [4-1:0] node48303;
	wire [4-1:0] node48306;
	wire [4-1:0] node48307;
	wire [4-1:0] node48310;
	wire [4-1:0] node48313;
	wire [4-1:0] node48314;
	wire [4-1:0] node48315;
	wire [4-1:0] node48318;
	wire [4-1:0] node48321;
	wire [4-1:0] node48322;
	wire [4-1:0] node48323;
	wire [4-1:0] node48327;
	wire [4-1:0] node48329;
	wire [4-1:0] node48332;
	wire [4-1:0] node48333;
	wire [4-1:0] node48334;
	wire [4-1:0] node48335;
	wire [4-1:0] node48336;
	wire [4-1:0] node48337;
	wire [4-1:0] node48341;
	wire [4-1:0] node48342;
	wire [4-1:0] node48343;
	wire [4-1:0] node48347;
	wire [4-1:0] node48350;
	wire [4-1:0] node48351;
	wire [4-1:0] node48352;
	wire [4-1:0] node48355;
	wire [4-1:0] node48357;
	wire [4-1:0] node48360;
	wire [4-1:0] node48361;
	wire [4-1:0] node48362;
	wire [4-1:0] node48365;
	wire [4-1:0] node48368;
	wire [4-1:0] node48369;
	wire [4-1:0] node48373;
	wire [4-1:0] node48374;
	wire [4-1:0] node48375;
	wire [4-1:0] node48376;
	wire [4-1:0] node48377;
	wire [4-1:0] node48380;
	wire [4-1:0] node48383;
	wire [4-1:0] node48385;
	wire [4-1:0] node48388;
	wire [4-1:0] node48389;
	wire [4-1:0] node48392;
	wire [4-1:0] node48395;
	wire [4-1:0] node48396;
	wire [4-1:0] node48397;
	wire [4-1:0] node48398;
	wire [4-1:0] node48402;
	wire [4-1:0] node48404;
	wire [4-1:0] node48407;
	wire [4-1:0] node48408;
	wire [4-1:0] node48411;
	wire [4-1:0] node48414;
	wire [4-1:0] node48415;
	wire [4-1:0] node48416;
	wire [4-1:0] node48417;
	wire [4-1:0] node48418;
	wire [4-1:0] node48421;
	wire [4-1:0] node48423;
	wire [4-1:0] node48426;
	wire [4-1:0] node48427;
	wire [4-1:0] node48430;
	wire [4-1:0] node48431;
	wire [4-1:0] node48435;
	wire [4-1:0] node48436;
	wire [4-1:0] node48438;
	wire [4-1:0] node48439;
	wire [4-1:0] node48443;
	wire [4-1:0] node48444;
	wire [4-1:0] node48445;
	wire [4-1:0] node48450;
	wire [4-1:0] node48451;
	wire [4-1:0] node48452;
	wire [4-1:0] node48454;
	wire [4-1:0] node48457;
	wire [4-1:0] node48458;
	wire [4-1:0] node48461;
	wire [4-1:0] node48464;
	wire [4-1:0] node48465;
	wire [4-1:0] node48466;
	wire [4-1:0] node48470;
	wire [4-1:0] node48471;
	wire [4-1:0] node48472;
	wire [4-1:0] node48476;
	wire [4-1:0] node48479;
	wire [4-1:0] node48480;
	wire [4-1:0] node48481;
	wire [4-1:0] node48482;
	wire [4-1:0] node48483;
	wire [4-1:0] node48484;
	wire [4-1:0] node48485;
	wire [4-1:0] node48486;
	wire [4-1:0] node48487;
	wire [4-1:0] node48490;
	wire [4-1:0] node48493;
	wire [4-1:0] node48495;
	wire [4-1:0] node48497;
	wire [4-1:0] node48500;
	wire [4-1:0] node48501;
	wire [4-1:0] node48502;
	wire [4-1:0] node48503;
	wire [4-1:0] node48507;
	wire [4-1:0] node48509;
	wire [4-1:0] node48512;
	wire [4-1:0] node48513;
	wire [4-1:0] node48514;
	wire [4-1:0] node48519;
	wire [4-1:0] node48520;
	wire [4-1:0] node48521;
	wire [4-1:0] node48522;
	wire [4-1:0] node48523;
	wire [4-1:0] node48526;
	wire [4-1:0] node48529;
	wire [4-1:0] node48531;
	wire [4-1:0] node48534;
	wire [4-1:0] node48535;
	wire [4-1:0] node48536;
	wire [4-1:0] node48539;
	wire [4-1:0] node48542;
	wire [4-1:0] node48543;
	wire [4-1:0] node48546;
	wire [4-1:0] node48549;
	wire [4-1:0] node48550;
	wire [4-1:0] node48552;
	wire [4-1:0] node48553;
	wire [4-1:0] node48556;
	wire [4-1:0] node48559;
	wire [4-1:0] node48560;
	wire [4-1:0] node48561;
	wire [4-1:0] node48564;
	wire [4-1:0] node48567;
	wire [4-1:0] node48568;
	wire [4-1:0] node48571;
	wire [4-1:0] node48574;
	wire [4-1:0] node48575;
	wire [4-1:0] node48576;
	wire [4-1:0] node48577;
	wire [4-1:0] node48578;
	wire [4-1:0] node48579;
	wire [4-1:0] node48582;
	wire [4-1:0] node48586;
	wire [4-1:0] node48587;
	wire [4-1:0] node48588;
	wire [4-1:0] node48592;
	wire [4-1:0] node48594;
	wire [4-1:0] node48597;
	wire [4-1:0] node48599;
	wire [4-1:0] node48600;
	wire [4-1:0] node48603;
	wire [4-1:0] node48605;
	wire [4-1:0] node48608;
	wire [4-1:0] node48609;
	wire [4-1:0] node48610;
	wire [4-1:0] node48611;
	wire [4-1:0] node48615;
	wire [4-1:0] node48616;
	wire [4-1:0] node48617;
	wire [4-1:0] node48622;
	wire [4-1:0] node48623;
	wire [4-1:0] node48624;
	wire [4-1:0] node48625;
	wire [4-1:0] node48628;
	wire [4-1:0] node48632;
	wire [4-1:0] node48634;
	wire [4-1:0] node48636;
	wire [4-1:0] node48639;
	wire [4-1:0] node48640;
	wire [4-1:0] node48641;
	wire [4-1:0] node48642;
	wire [4-1:0] node48643;
	wire [4-1:0] node48644;
	wire [4-1:0] node48647;
	wire [4-1:0] node48650;
	wire [4-1:0] node48653;
	wire [4-1:0] node48654;
	wire [4-1:0] node48655;
	wire [4-1:0] node48657;
	wire [4-1:0] node48661;
	wire [4-1:0] node48663;
	wire [4-1:0] node48664;
	wire [4-1:0] node48667;
	wire [4-1:0] node48670;
	wire [4-1:0] node48671;
	wire [4-1:0] node48672;
	wire [4-1:0] node48673;
	wire [4-1:0] node48674;
	wire [4-1:0] node48677;
	wire [4-1:0] node48680;
	wire [4-1:0] node48681;
	wire [4-1:0] node48685;
	wire [4-1:0] node48686;
	wire [4-1:0] node48687;
	wire [4-1:0] node48691;
	wire [4-1:0] node48692;
	wire [4-1:0] node48695;
	wire [4-1:0] node48698;
	wire [4-1:0] node48699;
	wire [4-1:0] node48701;
	wire [4-1:0] node48703;
	wire [4-1:0] node48706;
	wire [4-1:0] node48707;
	wire [4-1:0] node48709;
	wire [4-1:0] node48712;
	wire [4-1:0] node48713;
	wire [4-1:0] node48716;
	wire [4-1:0] node48719;
	wire [4-1:0] node48720;
	wire [4-1:0] node48721;
	wire [4-1:0] node48722;
	wire [4-1:0] node48723;
	wire [4-1:0] node48726;
	wire [4-1:0] node48729;
	wire [4-1:0] node48731;
	wire [4-1:0] node48732;
	wire [4-1:0] node48735;
	wire [4-1:0] node48738;
	wire [4-1:0] node48739;
	wire [4-1:0] node48741;
	wire [4-1:0] node48742;
	wire [4-1:0] node48746;
	wire [4-1:0] node48747;
	wire [4-1:0] node48748;
	wire [4-1:0] node48751;
	wire [4-1:0] node48754;
	wire [4-1:0] node48756;
	wire [4-1:0] node48759;
	wire [4-1:0] node48760;
	wire [4-1:0] node48761;
	wire [4-1:0] node48762;
	wire [4-1:0] node48765;
	wire [4-1:0] node48768;
	wire [4-1:0] node48769;
	wire [4-1:0] node48772;
	wire [4-1:0] node48775;
	wire [4-1:0] node48776;
	wire [4-1:0] node48778;
	wire [4-1:0] node48781;
	wire [4-1:0] node48783;
	wire [4-1:0] node48786;
	wire [4-1:0] node48787;
	wire [4-1:0] node48788;
	wire [4-1:0] node48789;
	wire [4-1:0] node48790;
	wire [4-1:0] node48791;
	wire [4-1:0] node48794;
	wire [4-1:0] node48796;
	wire [4-1:0] node48799;
	wire [4-1:0] node48800;
	wire [4-1:0] node48801;
	wire [4-1:0] node48802;
	wire [4-1:0] node48805;
	wire [4-1:0] node48809;
	wire [4-1:0] node48810;
	wire [4-1:0] node48813;
	wire [4-1:0] node48816;
	wire [4-1:0] node48817;
	wire [4-1:0] node48818;
	wire [4-1:0] node48819;
	wire [4-1:0] node48822;
	wire [4-1:0] node48825;
	wire [4-1:0] node48826;
	wire [4-1:0] node48829;
	wire [4-1:0] node48832;
	wire [4-1:0] node48833;
	wire [4-1:0] node48836;
	wire [4-1:0] node48837;
	wire [4-1:0] node48840;
	wire [4-1:0] node48843;
	wire [4-1:0] node48844;
	wire [4-1:0] node48845;
	wire [4-1:0] node48846;
	wire [4-1:0] node48848;
	wire [4-1:0] node48852;
	wire [4-1:0] node48853;
	wire [4-1:0] node48855;
	wire [4-1:0] node48858;
	wire [4-1:0] node48860;
	wire [4-1:0] node48863;
	wire [4-1:0] node48864;
	wire [4-1:0] node48865;
	wire [4-1:0] node48868;
	wire [4-1:0] node48870;
	wire [4-1:0] node48873;
	wire [4-1:0] node48874;
	wire [4-1:0] node48875;
	wire [4-1:0] node48878;
	wire [4-1:0] node48881;
	wire [4-1:0] node48882;
	wire [4-1:0] node48883;
	wire [4-1:0] node48886;
	wire [4-1:0] node48889;
	wire [4-1:0] node48891;
	wire [4-1:0] node48894;
	wire [4-1:0] node48895;
	wire [4-1:0] node48896;
	wire [4-1:0] node48897;
	wire [4-1:0] node48898;
	wire [4-1:0] node48899;
	wire [4-1:0] node48902;
	wire [4-1:0] node48905;
	wire [4-1:0] node48907;
	wire [4-1:0] node48910;
	wire [4-1:0] node48912;
	wire [4-1:0] node48913;
	wire [4-1:0] node48916;
	wire [4-1:0] node48919;
	wire [4-1:0] node48920;
	wire [4-1:0] node48921;
	wire [4-1:0] node48923;
	wire [4-1:0] node48924;
	wire [4-1:0] node48927;
	wire [4-1:0] node48930;
	wire [4-1:0] node48931;
	wire [4-1:0] node48933;
	wire [4-1:0] node48936;
	wire [4-1:0] node48937;
	wire [4-1:0] node48940;
	wire [4-1:0] node48943;
	wire [4-1:0] node48944;
	wire [4-1:0] node48945;
	wire [4-1:0] node48948;
	wire [4-1:0] node48951;
	wire [4-1:0] node48952;
	wire [4-1:0] node48953;
	wire [4-1:0] node48956;
	wire [4-1:0] node48959;
	wire [4-1:0] node48960;
	wire [4-1:0] node48964;
	wire [4-1:0] node48965;
	wire [4-1:0] node48966;
	wire [4-1:0] node48968;
	wire [4-1:0] node48969;
	wire [4-1:0] node48972;
	wire [4-1:0] node48975;
	wire [4-1:0] node48976;
	wire [4-1:0] node48978;
	wire [4-1:0] node48979;
	wire [4-1:0] node48982;
	wire [4-1:0] node48985;
	wire [4-1:0] node48986;
	wire [4-1:0] node48989;
	wire [4-1:0] node48992;
	wire [4-1:0] node48993;
	wire [4-1:0] node48994;
	wire [4-1:0] node48995;
	wire [4-1:0] node48998;
	wire [4-1:0] node49001;
	wire [4-1:0] node49002;
	wire [4-1:0] node49005;
	wire [4-1:0] node49008;
	wire [4-1:0] node49009;
	wire [4-1:0] node49010;
	wire [4-1:0] node49013;
	wire [4-1:0] node49016;
	wire [4-1:0] node49018;
	wire [4-1:0] node49021;
	wire [4-1:0] node49022;
	wire [4-1:0] node49023;
	wire [4-1:0] node49024;
	wire [4-1:0] node49025;
	wire [4-1:0] node49026;
	wire [4-1:0] node49027;
	wire [4-1:0] node49030;
	wire [4-1:0] node49031;
	wire [4-1:0] node49034;
	wire [4-1:0] node49036;
	wire [4-1:0] node49039;
	wire [4-1:0] node49040;
	wire [4-1:0] node49041;
	wire [4-1:0] node49042;
	wire [4-1:0] node49047;
	wire [4-1:0] node49049;
	wire [4-1:0] node49050;
	wire [4-1:0] node49054;
	wire [4-1:0] node49055;
	wire [4-1:0] node49056;
	wire [4-1:0] node49057;
	wire [4-1:0] node49058;
	wire [4-1:0] node49061;
	wire [4-1:0] node49064;
	wire [4-1:0] node49065;
	wire [4-1:0] node49068;
	wire [4-1:0] node49071;
	wire [4-1:0] node49072;
	wire [4-1:0] node49073;
	wire [4-1:0] node49076;
	wire [4-1:0] node49079;
	wire [4-1:0] node49080;
	wire [4-1:0] node49083;
	wire [4-1:0] node49086;
	wire [4-1:0] node49087;
	wire [4-1:0] node49088;
	wire [4-1:0] node49092;
	wire [4-1:0] node49094;
	wire [4-1:0] node49097;
	wire [4-1:0] node49098;
	wire [4-1:0] node49099;
	wire [4-1:0] node49100;
	wire [4-1:0] node49101;
	wire [4-1:0] node49104;
	wire [4-1:0] node49106;
	wire [4-1:0] node49109;
	wire [4-1:0] node49110;
	wire [4-1:0] node49113;
	wire [4-1:0] node49115;
	wire [4-1:0] node49118;
	wire [4-1:0] node49119;
	wire [4-1:0] node49122;
	wire [4-1:0] node49124;
	wire [4-1:0] node49127;
	wire [4-1:0] node49128;
	wire [4-1:0] node49129;
	wire [4-1:0] node49130;
	wire [4-1:0] node49131;
	wire [4-1:0] node49135;
	wire [4-1:0] node49136;
	wire [4-1:0] node49139;
	wire [4-1:0] node49142;
	wire [4-1:0] node49143;
	wire [4-1:0] node49144;
	wire [4-1:0] node49147;
	wire [4-1:0] node49150;
	wire [4-1:0] node49152;
	wire [4-1:0] node49155;
	wire [4-1:0] node49156;
	wire [4-1:0] node49157;
	wire [4-1:0] node49159;
	wire [4-1:0] node49163;
	wire [4-1:0] node49165;
	wire [4-1:0] node49166;
	wire [4-1:0] node49169;
	wire [4-1:0] node49172;
	wire [4-1:0] node49173;
	wire [4-1:0] node49174;
	wire [4-1:0] node49175;
	wire [4-1:0] node49176;
	wire [4-1:0] node49178;
	wire [4-1:0] node49181;
	wire [4-1:0] node49182;
	wire [4-1:0] node49185;
	wire [4-1:0] node49188;
	wire [4-1:0] node49189;
	wire [4-1:0] node49190;
	wire [4-1:0] node49192;
	wire [4-1:0] node49195;
	wire [4-1:0] node49196;
	wire [4-1:0] node49199;
	wire [4-1:0] node49202;
	wire [4-1:0] node49203;
	wire [4-1:0] node49204;
	wire [4-1:0] node49207;
	wire [4-1:0] node49210;
	wire [4-1:0] node49211;
	wire [4-1:0] node49214;
	wire [4-1:0] node49217;
	wire [4-1:0] node49218;
	wire [4-1:0] node49219;
	wire [4-1:0] node49220;
	wire [4-1:0] node49221;
	wire [4-1:0] node49224;
	wire [4-1:0] node49227;
	wire [4-1:0] node49229;
	wire [4-1:0] node49232;
	wire [4-1:0] node49233;
	wire [4-1:0] node49237;
	wire [4-1:0] node49238;
	wire [4-1:0] node49240;
	wire [4-1:0] node49241;
	wire [4-1:0] node49244;
	wire [4-1:0] node49247;
	wire [4-1:0] node49248;
	wire [4-1:0] node49251;
	wire [4-1:0] node49254;
	wire [4-1:0] node49255;
	wire [4-1:0] node49256;
	wire [4-1:0] node49257;
	wire [4-1:0] node49258;
	wire [4-1:0] node49263;
	wire [4-1:0] node49265;
	wire [4-1:0] node49266;
	wire [4-1:0] node49269;
	wire [4-1:0] node49272;
	wire [4-1:0] node49273;
	wire [4-1:0] node49274;
	wire [4-1:0] node49275;
	wire [4-1:0] node49276;
	wire [4-1:0] node49280;
	wire [4-1:0] node49282;
	wire [4-1:0] node49285;
	wire [4-1:0] node49286;
	wire [4-1:0] node49290;
	wire [4-1:0] node49291;
	wire [4-1:0] node49292;
	wire [4-1:0] node49296;
	wire [4-1:0] node49297;
	wire [4-1:0] node49301;
	wire [4-1:0] node49302;
	wire [4-1:0] node49303;
	wire [4-1:0] node49304;
	wire [4-1:0] node49305;
	wire [4-1:0] node49306;
	wire [4-1:0] node49307;
	wire [4-1:0] node49309;
	wire [4-1:0] node49312;
	wire [4-1:0] node49313;
	wire [4-1:0] node49317;
	wire [4-1:0] node49318;
	wire [4-1:0] node49319;
	wire [4-1:0] node49323;
	wire [4-1:0] node49324;
	wire [4-1:0] node49328;
	wire [4-1:0] node49329;
	wire [4-1:0] node49330;
	wire [4-1:0] node49331;
	wire [4-1:0] node49335;
	wire [4-1:0] node49336;
	wire [4-1:0] node49339;
	wire [4-1:0] node49342;
	wire [4-1:0] node49343;
	wire [4-1:0] node49344;
	wire [4-1:0] node49348;
	wire [4-1:0] node49349;
	wire [4-1:0] node49353;
	wire [4-1:0] node49354;
	wire [4-1:0] node49355;
	wire [4-1:0] node49356;
	wire [4-1:0] node49359;
	wire [4-1:0] node49361;
	wire [4-1:0] node49364;
	wire [4-1:0] node49366;
	wire [4-1:0] node49368;
	wire [4-1:0] node49371;
	wire [4-1:0] node49372;
	wire [4-1:0] node49373;
	wire [4-1:0] node49377;
	wire [4-1:0] node49378;
	wire [4-1:0] node49380;
	wire [4-1:0] node49383;
	wire [4-1:0] node49386;
	wire [4-1:0] node49387;
	wire [4-1:0] node49388;
	wire [4-1:0] node49389;
	wire [4-1:0] node49390;
	wire [4-1:0] node49392;
	wire [4-1:0] node49395;
	wire [4-1:0] node49396;
	wire [4-1:0] node49400;
	wire [4-1:0] node49401;
	wire [4-1:0] node49404;
	wire [4-1:0] node49407;
	wire [4-1:0] node49408;
	wire [4-1:0] node49409;
	wire [4-1:0] node49413;
	wire [4-1:0] node49416;
	wire [4-1:0] node49417;
	wire [4-1:0] node49418;
	wire [4-1:0] node49419;
	wire [4-1:0] node49422;
	wire [4-1:0] node49423;
	wire [4-1:0] node49427;
	wire [4-1:0] node49428;
	wire [4-1:0] node49431;
	wire [4-1:0] node49434;
	wire [4-1:0] node49435;
	wire [4-1:0] node49436;
	wire [4-1:0] node49439;
	wire [4-1:0] node49443;
	wire [4-1:0] node49444;
	wire [4-1:0] node49445;
	wire [4-1:0] node49446;
	wire [4-1:0] node49447;
	wire [4-1:0] node49449;
	wire [4-1:0] node49452;
	wire [4-1:0] node49454;
	wire [4-1:0] node49457;
	wire [4-1:0] node49458;
	wire [4-1:0] node49460;
	wire [4-1:0] node49463;
	wire [4-1:0] node49465;
	wire [4-1:0] node49468;
	wire [4-1:0] node49469;
	wire [4-1:0] node49470;
	wire [4-1:0] node49471;
	wire [4-1:0] node49472;
	wire [4-1:0] node49475;
	wire [4-1:0] node49479;
	wire [4-1:0] node49480;
	wire [4-1:0] node49484;
	wire [4-1:0] node49487;
	wire [4-1:0] node49488;
	wire [4-1:0] node49489;
	wire [4-1:0] node49490;
	wire [4-1:0] node49492;
	wire [4-1:0] node49493;
	wire [4-1:0] node49496;
	wire [4-1:0] node49499;
	wire [4-1:0] node49500;
	wire [4-1:0] node49502;
	wire [4-1:0] node49505;
	wire [4-1:0] node49506;
	wire [4-1:0] node49509;
	wire [4-1:0] node49512;
	wire [4-1:0] node49513;
	wire [4-1:0] node49516;
	wire [4-1:0] node49519;
	wire [4-1:0] node49520;
	wire [4-1:0] node49521;
	wire [4-1:0] node49522;
	wire [4-1:0] node49526;
	wire [4-1:0] node49527;
	wire [4-1:0] node49531;
	wire [4-1:0] node49532;
	wire [4-1:0] node49534;
	wire [4-1:0] node49537;
	wire [4-1:0] node49538;
	wire [4-1:0] node49542;
	wire [4-1:0] node49543;
	wire [4-1:0] node49544;
	wire [4-1:0] node49545;
	wire [4-1:0] node49546;
	wire [4-1:0] node49547;
	wire [4-1:0] node49548;
	wire [4-1:0] node49549;
	wire [4-1:0] node49550;
	wire [4-1:0] node49551;
	wire [4-1:0] node49552;
	wire [4-1:0] node49555;
	wire [4-1:0] node49559;
	wire [4-1:0] node49561;
	wire [4-1:0] node49564;
	wire [4-1:0] node49565;
	wire [4-1:0] node49566;
	wire [4-1:0] node49567;
	wire [4-1:0] node49570;
	wire [4-1:0] node49574;
	wire [4-1:0] node49575;
	wire [4-1:0] node49576;
	wire [4-1:0] node49580;
	wire [4-1:0] node49581;
	wire [4-1:0] node49584;
	wire [4-1:0] node49587;
	wire [4-1:0] node49588;
	wire [4-1:0] node49589;
	wire [4-1:0] node49590;
	wire [4-1:0] node49592;
	wire [4-1:0] node49595;
	wire [4-1:0] node49597;
	wire [4-1:0] node49600;
	wire [4-1:0] node49602;
	wire [4-1:0] node49605;
	wire [4-1:0] node49606;
	wire [4-1:0] node49608;
	wire [4-1:0] node49609;
	wire [4-1:0] node49612;
	wire [4-1:0] node49615;
	wire [4-1:0] node49616;
	wire [4-1:0] node49619;
	wire [4-1:0] node49622;
	wire [4-1:0] node49623;
	wire [4-1:0] node49624;
	wire [4-1:0] node49625;
	wire [4-1:0] node49626;
	wire [4-1:0] node49629;
	wire [4-1:0] node49632;
	wire [4-1:0] node49633;
	wire [4-1:0] node49634;
	wire [4-1:0] node49637;
	wire [4-1:0] node49640;
	wire [4-1:0] node49641;
	wire [4-1:0] node49644;
	wire [4-1:0] node49647;
	wire [4-1:0] node49648;
	wire [4-1:0] node49651;
	wire [4-1:0] node49652;
	wire [4-1:0] node49653;
	wire [4-1:0] node49656;
	wire [4-1:0] node49659;
	wire [4-1:0] node49660;
	wire [4-1:0] node49663;
	wire [4-1:0] node49666;
	wire [4-1:0] node49667;
	wire [4-1:0] node49668;
	wire [4-1:0] node49670;
	wire [4-1:0] node49673;
	wire [4-1:0] node49674;
	wire [4-1:0] node49676;
	wire [4-1:0] node49679;
	wire [4-1:0] node49680;
	wire [4-1:0] node49684;
	wire [4-1:0] node49685;
	wire [4-1:0] node49686;
	wire [4-1:0] node49687;
	wire [4-1:0] node49690;
	wire [4-1:0] node49693;
	wire [4-1:0] node49694;
	wire [4-1:0] node49697;
	wire [4-1:0] node49700;
	wire [4-1:0] node49701;
	wire [4-1:0] node49702;
	wire [4-1:0] node49707;
	wire [4-1:0] node49708;
	wire [4-1:0] node49709;
	wire [4-1:0] node49710;
	wire [4-1:0] node49711;
	wire [4-1:0] node49713;
	wire [4-1:0] node49714;
	wire [4-1:0] node49718;
	wire [4-1:0] node49719;
	wire [4-1:0] node49723;
	wire [4-1:0] node49724;
	wire [4-1:0] node49725;
	wire [4-1:0] node49726;
	wire [4-1:0] node49729;
	wire [4-1:0] node49733;
	wire [4-1:0] node49735;
	wire [4-1:0] node49738;
	wire [4-1:0] node49739;
	wire [4-1:0] node49740;
	wire [4-1:0] node49741;
	wire [4-1:0] node49742;
	wire [4-1:0] node49745;
	wire [4-1:0] node49748;
	wire [4-1:0] node49749;
	wire [4-1:0] node49752;
	wire [4-1:0] node49755;
	wire [4-1:0] node49756;
	wire [4-1:0] node49757;
	wire [4-1:0] node49760;
	wire [4-1:0] node49763;
	wire [4-1:0] node49765;
	wire [4-1:0] node49768;
	wire [4-1:0] node49769;
	wire [4-1:0] node49771;
	wire [4-1:0] node49774;
	wire [4-1:0] node49775;
	wire [4-1:0] node49778;
	wire [4-1:0] node49780;
	wire [4-1:0] node49783;
	wire [4-1:0] node49784;
	wire [4-1:0] node49785;
	wire [4-1:0] node49786;
	wire [4-1:0] node49788;
	wire [4-1:0] node49790;
	wire [4-1:0] node49793;
	wire [4-1:0] node49795;
	wire [4-1:0] node49796;
	wire [4-1:0] node49799;
	wire [4-1:0] node49802;
	wire [4-1:0] node49803;
	wire [4-1:0] node49805;
	wire [4-1:0] node49807;
	wire [4-1:0] node49810;
	wire [4-1:0] node49811;
	wire [4-1:0] node49814;
	wire [4-1:0] node49817;
	wire [4-1:0] node49818;
	wire [4-1:0] node49819;
	wire [4-1:0] node49820;
	wire [4-1:0] node49821;
	wire [4-1:0] node49825;
	wire [4-1:0] node49828;
	wire [4-1:0] node49829;
	wire [4-1:0] node49830;
	wire [4-1:0] node49834;
	wire [4-1:0] node49835;
	wire [4-1:0] node49838;
	wire [4-1:0] node49841;
	wire [4-1:0] node49842;
	wire [4-1:0] node49843;
	wire [4-1:0] node49846;
	wire [4-1:0] node49849;
	wire [4-1:0] node49851;
	wire [4-1:0] node49854;
	wire [4-1:0] node49855;
	wire [4-1:0] node49856;
	wire [4-1:0] node49857;
	wire [4-1:0] node49858;
	wire [4-1:0] node49859;
	wire [4-1:0] node49861;
	wire [4-1:0] node49864;
	wire [4-1:0] node49865;
	wire [4-1:0] node49868;
	wire [4-1:0] node49871;
	wire [4-1:0] node49872;
	wire [4-1:0] node49874;
	wire [4-1:0] node49877;
	wire [4-1:0] node49878;
	wire [4-1:0] node49881;
	wire [4-1:0] node49884;
	wire [4-1:0] node49885;
	wire [4-1:0] node49886;
	wire [4-1:0] node49887;
	wire [4-1:0] node49888;
	wire [4-1:0] node49893;
	wire [4-1:0] node49894;
	wire [4-1:0] node49897;
	wire [4-1:0] node49899;
	wire [4-1:0] node49902;
	wire [4-1:0] node49903;
	wire [4-1:0] node49904;
	wire [4-1:0] node49907;
	wire [4-1:0] node49910;
	wire [4-1:0] node49911;
	wire [4-1:0] node49912;
	wire [4-1:0] node49916;
	wire [4-1:0] node49918;
	wire [4-1:0] node49921;
	wire [4-1:0] node49922;
	wire [4-1:0] node49923;
	wire [4-1:0] node49924;
	wire [4-1:0] node49927;
	wire [4-1:0] node49929;
	wire [4-1:0] node49932;
	wire [4-1:0] node49933;
	wire [4-1:0] node49934;
	wire [4-1:0] node49936;
	wire [4-1:0] node49939;
	wire [4-1:0] node49942;
	wire [4-1:0] node49943;
	wire [4-1:0] node49946;
	wire [4-1:0] node49949;
	wire [4-1:0] node49950;
	wire [4-1:0] node49951;
	wire [4-1:0] node49952;
	wire [4-1:0] node49957;
	wire [4-1:0] node49958;
	wire [4-1:0] node49959;
	wire [4-1:0] node49962;
	wire [4-1:0] node49965;
	wire [4-1:0] node49966;
	wire [4-1:0] node49968;
	wire [4-1:0] node49971;
	wire [4-1:0] node49972;
	wire [4-1:0] node49976;
	wire [4-1:0] node49977;
	wire [4-1:0] node49978;
	wire [4-1:0] node49979;
	wire [4-1:0] node49980;
	wire [4-1:0] node49981;
	wire [4-1:0] node49984;
	wire [4-1:0] node49987;
	wire [4-1:0] node49988;
	wire [4-1:0] node49991;
	wire [4-1:0] node49994;
	wire [4-1:0] node49995;
	wire [4-1:0] node49998;
	wire [4-1:0] node50001;
	wire [4-1:0] node50002;
	wire [4-1:0] node50003;
	wire [4-1:0] node50004;
	wire [4-1:0] node50005;
	wire [4-1:0] node50008;
	wire [4-1:0] node50011;
	wire [4-1:0] node50012;
	wire [4-1:0] node50016;
	wire [4-1:0] node50018;
	wire [4-1:0] node50021;
	wire [4-1:0] node50022;
	wire [4-1:0] node50023;
	wire [4-1:0] node50027;
	wire [4-1:0] node50030;
	wire [4-1:0] node50031;
	wire [4-1:0] node50032;
	wire [4-1:0] node50033;
	wire [4-1:0] node50034;
	wire [4-1:0] node50037;
	wire [4-1:0] node50040;
	wire [4-1:0] node50041;
	wire [4-1:0] node50043;
	wire [4-1:0] node50046;
	wire [4-1:0] node50049;
	wire [4-1:0] node50050;
	wire [4-1:0] node50053;
	wire [4-1:0] node50056;
	wire [4-1:0] node50057;
	wire [4-1:0] node50058;
	wire [4-1:0] node50059;
	wire [4-1:0] node50060;
	wire [4-1:0] node50063;
	wire [4-1:0] node50067;
	wire [4-1:0] node50068;
	wire [4-1:0] node50071;
	wire [4-1:0] node50074;
	wire [4-1:0] node50075;
	wire [4-1:0] node50076;
	wire [4-1:0] node50080;
	wire [4-1:0] node50083;
	wire [4-1:0] node50084;
	wire [4-1:0] node50085;
	wire [4-1:0] node50086;
	wire [4-1:0] node50087;
	wire [4-1:0] node50088;
	wire [4-1:0] node50089;
	wire [4-1:0] node50091;
	wire [4-1:0] node50092;
	wire [4-1:0] node50095;
	wire [4-1:0] node50098;
	wire [4-1:0] node50099;
	wire [4-1:0] node50100;
	wire [4-1:0] node50103;
	wire [4-1:0] node50106;
	wire [4-1:0] node50107;
	wire [4-1:0] node50111;
	wire [4-1:0] node50112;
	wire [4-1:0] node50113;
	wire [4-1:0] node50114;
	wire [4-1:0] node50118;
	wire [4-1:0] node50119;
	wire [4-1:0] node50123;
	wire [4-1:0] node50124;
	wire [4-1:0] node50125;
	wire [4-1:0] node50128;
	wire [4-1:0] node50131;
	wire [4-1:0] node50133;
	wire [4-1:0] node50136;
	wire [4-1:0] node50137;
	wire [4-1:0] node50138;
	wire [4-1:0] node50139;
	wire [4-1:0] node50140;
	wire [4-1:0] node50143;
	wire [4-1:0] node50146;
	wire [4-1:0] node50147;
	wire [4-1:0] node50151;
	wire [4-1:0] node50154;
	wire [4-1:0] node50155;
	wire [4-1:0] node50157;
	wire [4-1:0] node50160;
	wire [4-1:0] node50161;
	wire [4-1:0] node50162;
	wire [4-1:0] node50166;
	wire [4-1:0] node50167;
	wire [4-1:0] node50171;
	wire [4-1:0] node50172;
	wire [4-1:0] node50173;
	wire [4-1:0] node50174;
	wire [4-1:0] node50175;
	wire [4-1:0] node50176;
	wire [4-1:0] node50179;
	wire [4-1:0] node50183;
	wire [4-1:0] node50185;
	wire [4-1:0] node50186;
	wire [4-1:0] node50190;
	wire [4-1:0] node50191;
	wire [4-1:0] node50193;
	wire [4-1:0] node50195;
	wire [4-1:0] node50198;
	wire [4-1:0] node50199;
	wire [4-1:0] node50200;
	wire [4-1:0] node50203;
	wire [4-1:0] node50207;
	wire [4-1:0] node50208;
	wire [4-1:0] node50209;
	wire [4-1:0] node50210;
	wire [4-1:0] node50211;
	wire [4-1:0] node50215;
	wire [4-1:0] node50218;
	wire [4-1:0] node50220;
	wire [4-1:0] node50221;
	wire [4-1:0] node50224;
	wire [4-1:0] node50227;
	wire [4-1:0] node50228;
	wire [4-1:0] node50230;
	wire [4-1:0] node50232;
	wire [4-1:0] node50235;
	wire [4-1:0] node50236;
	wire [4-1:0] node50238;
	wire [4-1:0] node50242;
	wire [4-1:0] node50243;
	wire [4-1:0] node50244;
	wire [4-1:0] node50245;
	wire [4-1:0] node50247;
	wire [4-1:0] node50248;
	wire [4-1:0] node50251;
	wire [4-1:0] node50254;
	wire [4-1:0] node50255;
	wire [4-1:0] node50256;
	wire [4-1:0] node50259;
	wire [4-1:0] node50262;
	wire [4-1:0] node50263;
	wire [4-1:0] node50265;
	wire [4-1:0] node50269;
	wire [4-1:0] node50270;
	wire [4-1:0] node50271;
	wire [4-1:0] node50272;
	wire [4-1:0] node50275;
	wire [4-1:0] node50278;
	wire [4-1:0] node50279;
	wire [4-1:0] node50282;
	wire [4-1:0] node50285;
	wire [4-1:0] node50286;
	wire [4-1:0] node50287;
	wire [4-1:0] node50288;
	wire [4-1:0] node50291;
	wire [4-1:0] node50294;
	wire [4-1:0] node50295;
	wire [4-1:0] node50298;
	wire [4-1:0] node50301;
	wire [4-1:0] node50302;
	wire [4-1:0] node50306;
	wire [4-1:0] node50307;
	wire [4-1:0] node50308;
	wire [4-1:0] node50309;
	wire [4-1:0] node50310;
	wire [4-1:0] node50311;
	wire [4-1:0] node50314;
	wire [4-1:0] node50317;
	wire [4-1:0] node50320;
	wire [4-1:0] node50321;
	wire [4-1:0] node50324;
	wire [4-1:0] node50326;
	wire [4-1:0] node50329;
	wire [4-1:0] node50330;
	wire [4-1:0] node50333;
	wire [4-1:0] node50334;
	wire [4-1:0] node50335;
	wire [4-1:0] node50338;
	wire [4-1:0] node50341;
	wire [4-1:0] node50344;
	wire [4-1:0] node50345;
	wire [4-1:0] node50346;
	wire [4-1:0] node50349;
	wire [4-1:0] node50351;
	wire [4-1:0] node50352;
	wire [4-1:0] node50355;
	wire [4-1:0] node50358;
	wire [4-1:0] node50359;
	wire [4-1:0] node50360;
	wire [4-1:0] node50364;
	wire [4-1:0] node50366;
	wire [4-1:0] node50367;
	wire [4-1:0] node50370;
	wire [4-1:0] node50373;
	wire [4-1:0] node50374;
	wire [4-1:0] node50375;
	wire [4-1:0] node50376;
	wire [4-1:0] node50377;
	wire [4-1:0] node50378;
	wire [4-1:0] node50379;
	wire [4-1:0] node50380;
	wire [4-1:0] node50384;
	wire [4-1:0] node50385;
	wire [4-1:0] node50389;
	wire [4-1:0] node50391;
	wire [4-1:0] node50394;
	wire [4-1:0] node50395;
	wire [4-1:0] node50397;
	wire [4-1:0] node50400;
	wire [4-1:0] node50401;
	wire [4-1:0] node50404;
	wire [4-1:0] node50407;
	wire [4-1:0] node50408;
	wire [4-1:0] node50409;
	wire [4-1:0] node50410;
	wire [4-1:0] node50413;
	wire [4-1:0] node50416;
	wire [4-1:0] node50417;
	wire [4-1:0] node50418;
	wire [4-1:0] node50423;
	wire [4-1:0] node50424;
	wire [4-1:0] node50426;
	wire [4-1:0] node50429;
	wire [4-1:0] node50431;
	wire [4-1:0] node50432;
	wire [4-1:0] node50435;
	wire [4-1:0] node50438;
	wire [4-1:0] node50439;
	wire [4-1:0] node50440;
	wire [4-1:0] node50441;
	wire [4-1:0] node50444;
	wire [4-1:0] node50445;
	wire [4-1:0] node50448;
	wire [4-1:0] node50451;
	wire [4-1:0] node50452;
	wire [4-1:0] node50453;
	wire [4-1:0] node50457;
	wire [4-1:0] node50460;
	wire [4-1:0] node50461;
	wire [4-1:0] node50462;
	wire [4-1:0] node50463;
	wire [4-1:0] node50465;
	wire [4-1:0] node50468;
	wire [4-1:0] node50471;
	wire [4-1:0] node50472;
	wire [4-1:0] node50475;
	wire [4-1:0] node50478;
	wire [4-1:0] node50479;
	wire [4-1:0] node50480;
	wire [4-1:0] node50484;
	wire [4-1:0] node50487;
	wire [4-1:0] node50488;
	wire [4-1:0] node50489;
	wire [4-1:0] node50490;
	wire [4-1:0] node50491;
	wire [4-1:0] node50492;
	wire [4-1:0] node50496;
	wire [4-1:0] node50497;
	wire [4-1:0] node50499;
	wire [4-1:0] node50502;
	wire [4-1:0] node50505;
	wire [4-1:0] node50506;
	wire [4-1:0] node50507;
	wire [4-1:0] node50510;
	wire [4-1:0] node50513;
	wire [4-1:0] node50515;
	wire [4-1:0] node50516;
	wire [4-1:0] node50520;
	wire [4-1:0] node50521;
	wire [4-1:0] node50522;
	wire [4-1:0] node50523;
	wire [4-1:0] node50524;
	wire [4-1:0] node50527;
	wire [4-1:0] node50530;
	wire [4-1:0] node50531;
	wire [4-1:0] node50534;
	wire [4-1:0] node50537;
	wire [4-1:0] node50538;
	wire [4-1:0] node50542;
	wire [4-1:0] node50545;
	wire [4-1:0] node50546;
	wire [4-1:0] node50547;
	wire [4-1:0] node50548;
	wire [4-1:0] node50549;
	wire [4-1:0] node50554;
	wire [4-1:0] node50556;
	wire [4-1:0] node50557;
	wire [4-1:0] node50561;
	wire [4-1:0] node50562;
	wire [4-1:0] node50563;
	wire [4-1:0] node50564;
	wire [4-1:0] node50565;
	wire [4-1:0] node50570;
	wire [4-1:0] node50571;
	wire [4-1:0] node50573;
	wire [4-1:0] node50576;
	wire [4-1:0] node50578;
	wire [4-1:0] node50581;
	wire [4-1:0] node50582;
	wire [4-1:0] node50584;
	wire [4-1:0] node50588;
	wire [4-1:0] node50589;
	wire [4-1:0] node50590;
	wire [4-1:0] node50591;
	wire [4-1:0] node50592;
	wire [4-1:0] node50593;
	wire [4-1:0] node50594;
	wire [4-1:0] node50595;
	wire [4-1:0] node50596;
	wire [4-1:0] node50597;
	wire [4-1:0] node50600;
	wire [4-1:0] node50603;
	wire [4-1:0] node50604;
	wire [4-1:0] node50607;
	wire [4-1:0] node50610;
	wire [4-1:0] node50611;
	wire [4-1:0] node50612;
	wire [4-1:0] node50615;
	wire [4-1:0] node50619;
	wire [4-1:0] node50620;
	wire [4-1:0] node50621;
	wire [4-1:0] node50623;
	wire [4-1:0] node50626;
	wire [4-1:0] node50627;
	wire [4-1:0] node50631;
	wire [4-1:0] node50632;
	wire [4-1:0] node50633;
	wire [4-1:0] node50637;
	wire [4-1:0] node50639;
	wire [4-1:0] node50642;
	wire [4-1:0] node50643;
	wire [4-1:0] node50645;
	wire [4-1:0] node50646;
	wire [4-1:0] node50649;
	wire [4-1:0] node50652;
	wire [4-1:0] node50653;
	wire [4-1:0] node50654;
	wire [4-1:0] node50655;
	wire [4-1:0] node50659;
	wire [4-1:0] node50662;
	wire [4-1:0] node50663;
	wire [4-1:0] node50664;
	wire [4-1:0] node50667;
	wire [4-1:0] node50670;
	wire [4-1:0] node50671;
	wire [4-1:0] node50674;
	wire [4-1:0] node50677;
	wire [4-1:0] node50678;
	wire [4-1:0] node50679;
	wire [4-1:0] node50680;
	wire [4-1:0] node50683;
	wire [4-1:0] node50684;
	wire [4-1:0] node50685;
	wire [4-1:0] node50688;
	wire [4-1:0] node50691;
	wire [4-1:0] node50692;
	wire [4-1:0] node50695;
	wire [4-1:0] node50698;
	wire [4-1:0] node50699;
	wire [4-1:0] node50700;
	wire [4-1:0] node50701;
	wire [4-1:0] node50706;
	wire [4-1:0] node50707;
	wire [4-1:0] node50709;
	wire [4-1:0] node50712;
	wire [4-1:0] node50714;
	wire [4-1:0] node50717;
	wire [4-1:0] node50718;
	wire [4-1:0] node50719;
	wire [4-1:0] node50722;
	wire [4-1:0] node50725;
	wire [4-1:0] node50726;
	wire [4-1:0] node50727;
	wire [4-1:0] node50732;
	wire [4-1:0] node50733;
	wire [4-1:0] node50734;
	wire [4-1:0] node50735;
	wire [4-1:0] node50736;
	wire [4-1:0] node50737;
	wire [4-1:0] node50740;
	wire [4-1:0] node50743;
	wire [4-1:0] node50744;
	wire [4-1:0] node50746;
	wire [4-1:0] node50749;
	wire [4-1:0] node50750;
	wire [4-1:0] node50754;
	wire [4-1:0] node50755;
	wire [4-1:0] node50757;
	wire [4-1:0] node50759;
	wire [4-1:0] node50762;
	wire [4-1:0] node50763;
	wire [4-1:0] node50767;
	wire [4-1:0] node50768;
	wire [4-1:0] node50769;
	wire [4-1:0] node50770;
	wire [4-1:0] node50771;
	wire [4-1:0] node50774;
	wire [4-1:0] node50777;
	wire [4-1:0] node50778;
	wire [4-1:0] node50782;
	wire [4-1:0] node50783;
	wire [4-1:0] node50786;
	wire [4-1:0] node50789;
	wire [4-1:0] node50790;
	wire [4-1:0] node50793;
	wire [4-1:0] node50796;
	wire [4-1:0] node50797;
	wire [4-1:0] node50798;
	wire [4-1:0] node50799;
	wire [4-1:0] node50801;
	wire [4-1:0] node50802;
	wire [4-1:0] node50806;
	wire [4-1:0] node50808;
	wire [4-1:0] node50811;
	wire [4-1:0] node50812;
	wire [4-1:0] node50816;
	wire [4-1:0] node50817;
	wire [4-1:0] node50819;
	wire [4-1:0] node50822;
	wire [4-1:0] node50823;
	wire [4-1:0] node50825;
	wire [4-1:0] node50826;
	wire [4-1:0] node50831;
	wire [4-1:0] node50832;
	wire [4-1:0] node50833;
	wire [4-1:0] node50834;
	wire [4-1:0] node50835;
	wire [4-1:0] node50838;
	wire [4-1:0] node50841;
	wire [4-1:0] node50842;
	wire [4-1:0] node50843;
	wire [4-1:0] node50844;
	wire [4-1:0] node50846;
	wire [4-1:0] node50850;
	wire [4-1:0] node50852;
	wire [4-1:0] node50854;
	wire [4-1:0] node50857;
	wire [4-1:0] node50858;
	wire [4-1:0] node50861;
	wire [4-1:0] node50864;
	wire [4-1:0] node50865;
	wire [4-1:0] node50866;
	wire [4-1:0] node50867;
	wire [4-1:0] node50868;
	wire [4-1:0] node50869;
	wire [4-1:0] node50872;
	wire [4-1:0] node50876;
	wire [4-1:0] node50877;
	wire [4-1:0] node50880;
	wire [4-1:0] node50883;
	wire [4-1:0] node50884;
	wire [4-1:0] node50885;
	wire [4-1:0] node50888;
	wire [4-1:0] node50891;
	wire [4-1:0] node50892;
	wire [4-1:0] node50895;
	wire [4-1:0] node50898;
	wire [4-1:0] node50899;
	wire [4-1:0] node50900;
	wire [4-1:0] node50902;
	wire [4-1:0] node50905;
	wire [4-1:0] node50907;
	wire [4-1:0] node50909;
	wire [4-1:0] node50912;
	wire [4-1:0] node50913;
	wire [4-1:0] node50914;
	wire [4-1:0] node50916;
	wire [4-1:0] node50919;
	wire [4-1:0] node50920;
	wire [4-1:0] node50924;
	wire [4-1:0] node50925;
	wire [4-1:0] node50927;
	wire [4-1:0] node50931;
	wire [4-1:0] node50932;
	wire [4-1:0] node50933;
	wire [4-1:0] node50934;
	wire [4-1:0] node50935;
	wire [4-1:0] node50936;
	wire [4-1:0] node50937;
	wire [4-1:0] node50941;
	wire [4-1:0] node50942;
	wire [4-1:0] node50945;
	wire [4-1:0] node50948;
	wire [4-1:0] node50949;
	wire [4-1:0] node50950;
	wire [4-1:0] node50954;
	wire [4-1:0] node50955;
	wire [4-1:0] node50958;
	wire [4-1:0] node50961;
	wire [4-1:0] node50963;
	wire [4-1:0] node50965;
	wire [4-1:0] node50966;
	wire [4-1:0] node50969;
	wire [4-1:0] node50972;
	wire [4-1:0] node50973;
	wire [4-1:0] node50976;
	wire [4-1:0] node50979;
	wire [4-1:0] node50980;
	wire [4-1:0] node50981;
	wire [4-1:0] node50983;
	wire [4-1:0] node50984;
	wire [4-1:0] node50987;
	wire [4-1:0] node50990;
	wire [4-1:0] node50991;
	wire [4-1:0] node50993;
	wire [4-1:0] node50997;
	wire [4-1:0] node50998;
	wire [4-1:0] node50999;
	wire [4-1:0] node51000;
	wire [4-1:0] node51003;
	wire [4-1:0] node51006;
	wire [4-1:0] node51009;
	wire [4-1:0] node51011;
	wire [4-1:0] node51012;
	wire [4-1:0] node51015;
	wire [4-1:0] node51018;
	wire [4-1:0] node51019;
	wire [4-1:0] node51020;
	wire [4-1:0] node51021;
	wire [4-1:0] node51022;
	wire [4-1:0] node51023;
	wire [4-1:0] node51024;
	wire [4-1:0] node51025;
	wire [4-1:0] node51028;
	wire [4-1:0] node51031;
	wire [4-1:0] node51032;
	wire [4-1:0] node51034;
	wire [4-1:0] node51037;
	wire [4-1:0] node51038;
	wire [4-1:0] node51042;
	wire [4-1:0] node51043;
	wire [4-1:0] node51044;
	wire [4-1:0] node51046;
	wire [4-1:0] node51049;
	wire [4-1:0] node51050;
	wire [4-1:0] node51055;
	wire [4-1:0] node51056;
	wire [4-1:0] node51057;
	wire [4-1:0] node51059;
	wire [4-1:0] node51062;
	wire [4-1:0] node51063;
	wire [4-1:0] node51064;
	wire [4-1:0] node51067;
	wire [4-1:0] node51070;
	wire [4-1:0] node51071;
	wire [4-1:0] node51074;
	wire [4-1:0] node51077;
	wire [4-1:0] node51078;
	wire [4-1:0] node51079;
	wire [4-1:0] node51080;
	wire [4-1:0] node51084;
	wire [4-1:0] node51087;
	wire [4-1:0] node51088;
	wire [4-1:0] node51091;
	wire [4-1:0] node51094;
	wire [4-1:0] node51095;
	wire [4-1:0] node51096;
	wire [4-1:0] node51097;
	wire [4-1:0] node51098;
	wire [4-1:0] node51101;
	wire [4-1:0] node51105;
	wire [4-1:0] node51106;
	wire [4-1:0] node51107;
	wire [4-1:0] node51108;
	wire [4-1:0] node51113;
	wire [4-1:0] node51114;
	wire [4-1:0] node51115;
	wire [4-1:0] node51119;
	wire [4-1:0] node51120;
	wire [4-1:0] node51123;
	wire [4-1:0] node51126;
	wire [4-1:0] node51127;
	wire [4-1:0] node51128;
	wire [4-1:0] node51129;
	wire [4-1:0] node51132;
	wire [4-1:0] node51135;
	wire [4-1:0] node51136;
	wire [4-1:0] node51137;
	wire [4-1:0] node51140;
	wire [4-1:0] node51143;
	wire [4-1:0] node51144;
	wire [4-1:0] node51147;
	wire [4-1:0] node51150;
	wire [4-1:0] node51151;
	wire [4-1:0] node51152;
	wire [4-1:0] node51153;
	wire [4-1:0] node51158;
	wire [4-1:0] node51159;
	wire [4-1:0] node51161;
	wire [4-1:0] node51164;
	wire [4-1:0] node51166;
	wire [4-1:0] node51169;
	wire [4-1:0] node51170;
	wire [4-1:0] node51171;
	wire [4-1:0] node51172;
	wire [4-1:0] node51173;
	wire [4-1:0] node51177;
	wire [4-1:0] node51179;
	wire [4-1:0] node51181;
	wire [4-1:0] node51184;
	wire [4-1:0] node51185;
	wire [4-1:0] node51186;
	wire [4-1:0] node51188;
	wire [4-1:0] node51189;
	wire [4-1:0] node51193;
	wire [4-1:0] node51194;
	wire [4-1:0] node51195;
	wire [4-1:0] node51199;
	wire [4-1:0] node51200;
	wire [4-1:0] node51204;
	wire [4-1:0] node51205;
	wire [4-1:0] node51206;
	wire [4-1:0] node51207;
	wire [4-1:0] node51211;
	wire [4-1:0] node51212;
	wire [4-1:0] node51217;
	wire [4-1:0] node51218;
	wire [4-1:0] node51219;
	wire [4-1:0] node51220;
	wire [4-1:0] node51221;
	wire [4-1:0] node51226;
	wire [4-1:0] node51227;
	wire [4-1:0] node51228;
	wire [4-1:0] node51231;
	wire [4-1:0] node51234;
	wire [4-1:0] node51236;
	wire [4-1:0] node51239;
	wire [4-1:0] node51240;
	wire [4-1:0] node51241;
	wire [4-1:0] node51243;
	wire [4-1:0] node51246;
	wire [4-1:0] node51247;
	wire [4-1:0] node51250;
	wire [4-1:0] node51253;
	wire [4-1:0] node51254;
	wire [4-1:0] node51255;
	wire [4-1:0] node51256;
	wire [4-1:0] node51260;
	wire [4-1:0] node51263;
	wire [4-1:0] node51264;
	wire [4-1:0] node51267;
	wire [4-1:0] node51270;
	wire [4-1:0] node51271;
	wire [4-1:0] node51272;
	wire [4-1:0] node51273;
	wire [4-1:0] node51274;
	wire [4-1:0] node51276;
	wire [4-1:0] node51279;
	wire [4-1:0] node51281;
	wire [4-1:0] node51284;
	wire [4-1:0] node51285;
	wire [4-1:0] node51287;
	wire [4-1:0] node51290;
	wire [4-1:0] node51292;
	wire [4-1:0] node51295;
	wire [4-1:0] node51296;
	wire [4-1:0] node51297;
	wire [4-1:0] node51298;
	wire [4-1:0] node51299;
	wire [4-1:0] node51303;
	wire [4-1:0] node51304;
	wire [4-1:0] node51308;
	wire [4-1:0] node51309;
	wire [4-1:0] node51310;
	wire [4-1:0] node51315;
	wire [4-1:0] node51316;
	wire [4-1:0] node51319;
	wire [4-1:0] node51320;
	wire [4-1:0] node51321;
	wire [4-1:0] node51325;
	wire [4-1:0] node51326;
	wire [4-1:0] node51330;
	wire [4-1:0] node51331;
	wire [4-1:0] node51332;
	wire [4-1:0] node51333;
	wire [4-1:0] node51334;
	wire [4-1:0] node51335;
	wire [4-1:0] node51337;
	wire [4-1:0] node51340;
	wire [4-1:0] node51342;
	wire [4-1:0] node51345;
	wire [4-1:0] node51347;
	wire [4-1:0] node51348;
	wire [4-1:0] node51351;
	wire [4-1:0] node51354;
	wire [4-1:0] node51355;
	wire [4-1:0] node51357;
	wire [4-1:0] node51358;
	wire [4-1:0] node51362;
	wire [4-1:0] node51363;
	wire [4-1:0] node51366;
	wire [4-1:0] node51369;
	wire [4-1:0] node51370;
	wire [4-1:0] node51371;
	wire [4-1:0] node51373;
	wire [4-1:0] node51374;
	wire [4-1:0] node51377;
	wire [4-1:0] node51380;
	wire [4-1:0] node51381;
	wire [4-1:0] node51382;
	wire [4-1:0] node51386;
	wire [4-1:0] node51387;
	wire [4-1:0] node51391;
	wire [4-1:0] node51393;
	wire [4-1:0] node51396;
	wire [4-1:0] node51397;
	wire [4-1:0] node51398;
	wire [4-1:0] node51399;
	wire [4-1:0] node51403;
	wire [4-1:0] node51404;
	wire [4-1:0] node51408;
	wire [4-1:0] node51410;
	wire [4-1:0] node51411;
	wire [4-1:0] node51415;
	wire [4-1:0] node51416;
	wire [4-1:0] node51417;
	wire [4-1:0] node51418;
	wire [4-1:0] node51419;
	wire [4-1:0] node51420;
	wire [4-1:0] node51421;
	wire [4-1:0] node51422;
	wire [4-1:0] node51423;
	wire [4-1:0] node51424;
	wire [4-1:0] node51425;
	wire [4-1:0] node51427;
	wire [4-1:0] node51431;
	wire [4-1:0] node51432;
	wire [4-1:0] node51433;
	wire [4-1:0] node51437;
	wire [4-1:0] node51439;
	wire [4-1:0] node51442;
	wire [4-1:0] node51443;
	wire [4-1:0] node51444;
	wire [4-1:0] node51445;
	wire [4-1:0] node51449;
	wire [4-1:0] node51451;
	wire [4-1:0] node51454;
	wire [4-1:0] node51455;
	wire [4-1:0] node51459;
	wire [4-1:0] node51460;
	wire [4-1:0] node51461;
	wire [4-1:0] node51462;
	wire [4-1:0] node51465;
	wire [4-1:0] node51466;
	wire [4-1:0] node51471;
	wire [4-1:0] node51472;
	wire [4-1:0] node51475;
	wire [4-1:0] node51477;
	wire [4-1:0] node51480;
	wire [4-1:0] node51481;
	wire [4-1:0] node51482;
	wire [4-1:0] node51483;
	wire [4-1:0] node51484;
	wire [4-1:0] node51487;
	wire [4-1:0] node51490;
	wire [4-1:0] node51492;
	wire [4-1:0] node51493;
	wire [4-1:0] node51496;
	wire [4-1:0] node51499;
	wire [4-1:0] node51500;
	wire [4-1:0] node51502;
	wire [4-1:0] node51503;
	wire [4-1:0] node51507;
	wire [4-1:0] node51508;
	wire [4-1:0] node51510;
	wire [4-1:0] node51513;
	wire [4-1:0] node51515;
	wire [4-1:0] node51518;
	wire [4-1:0] node51519;
	wire [4-1:0] node51520;
	wire [4-1:0] node51521;
	wire [4-1:0] node51522;
	wire [4-1:0] node51525;
	wire [4-1:0] node51528;
	wire [4-1:0] node51530;
	wire [4-1:0] node51533;
	wire [4-1:0] node51534;
	wire [4-1:0] node51535;
	wire [4-1:0] node51538;
	wire [4-1:0] node51541;
	wire [4-1:0] node51543;
	wire [4-1:0] node51546;
	wire [4-1:0] node51547;
	wire [4-1:0] node51548;
	wire [4-1:0] node51549;
	wire [4-1:0] node51553;
	wire [4-1:0] node51555;
	wire [4-1:0] node51558;
	wire [4-1:0] node51560;
	wire [4-1:0] node51563;
	wire [4-1:0] node51564;
	wire [4-1:0] node51565;
	wire [4-1:0] node51566;
	wire [4-1:0] node51567;
	wire [4-1:0] node51568;
	wire [4-1:0] node51570;
	wire [4-1:0] node51573;
	wire [4-1:0] node51574;
	wire [4-1:0] node51577;
	wire [4-1:0] node51580;
	wire [4-1:0] node51581;
	wire [4-1:0] node51582;
	wire [4-1:0] node51585;
	wire [4-1:0] node51589;
	wire [4-1:0] node51590;
	wire [4-1:0] node51592;
	wire [4-1:0] node51593;
	wire [4-1:0] node51596;
	wire [4-1:0] node51599;
	wire [4-1:0] node51600;
	wire [4-1:0] node51601;
	wire [4-1:0] node51604;
	wire [4-1:0] node51608;
	wire [4-1:0] node51609;
	wire [4-1:0] node51610;
	wire [4-1:0] node51611;
	wire [4-1:0] node51614;
	wire [4-1:0] node51615;
	wire [4-1:0] node51619;
	wire [4-1:0] node51620;
	wire [4-1:0] node51622;
	wire [4-1:0] node51625;
	wire [4-1:0] node51628;
	wire [4-1:0] node51629;
	wire [4-1:0] node51630;
	wire [4-1:0] node51631;
	wire [4-1:0] node51634;
	wire [4-1:0] node51638;
	wire [4-1:0] node51639;
	wire [4-1:0] node51643;
	wire [4-1:0] node51644;
	wire [4-1:0] node51645;
	wire [4-1:0] node51646;
	wire [4-1:0] node51647;
	wire [4-1:0] node51650;
	wire [4-1:0] node51653;
	wire [4-1:0] node51654;
	wire [4-1:0] node51655;
	wire [4-1:0] node51658;
	wire [4-1:0] node51661;
	wire [4-1:0] node51662;
	wire [4-1:0] node51665;
	wire [4-1:0] node51668;
	wire [4-1:0] node51669;
	wire [4-1:0] node51670;
	wire [4-1:0] node51672;
	wire [4-1:0] node51676;
	wire [4-1:0] node51678;
	wire [4-1:0] node51679;
	wire [4-1:0] node51682;
	wire [4-1:0] node51685;
	wire [4-1:0] node51686;
	wire [4-1:0] node51687;
	wire [4-1:0] node51688;
	wire [4-1:0] node51692;
	wire [4-1:0] node51693;
	wire [4-1:0] node51695;
	wire [4-1:0] node51698;
	wire [4-1:0] node51701;
	wire [4-1:0] node51702;
	wire [4-1:0] node51703;
	wire [4-1:0] node51706;
	wire [4-1:0] node51709;
	wire [4-1:0] node51710;
	wire [4-1:0] node51713;
	wire [4-1:0] node51716;
	wire [4-1:0] node51717;
	wire [4-1:0] node51718;
	wire [4-1:0] node51719;
	wire [4-1:0] node51720;
	wire [4-1:0] node51721;
	wire [4-1:0] node51723;
	wire [4-1:0] node51726;
	wire [4-1:0] node51727;
	wire [4-1:0] node51731;
	wire [4-1:0] node51732;
	wire [4-1:0] node51735;
	wire [4-1:0] node51736;
	wire [4-1:0] node51739;
	wire [4-1:0] node51742;
	wire [4-1:0] node51743;
	wire [4-1:0] node51745;
	wire [4-1:0] node51746;
	wire [4-1:0] node51747;
	wire [4-1:0] node51750;
	wire [4-1:0] node51753;
	wire [4-1:0] node51754;
	wire [4-1:0] node51757;
	wire [4-1:0] node51760;
	wire [4-1:0] node51761;
	wire [4-1:0] node51762;
	wire [4-1:0] node51765;
	wire [4-1:0] node51768;
	wire [4-1:0] node51769;
	wire [4-1:0] node51772;
	wire [4-1:0] node51775;
	wire [4-1:0] node51776;
	wire [4-1:0] node51777;
	wire [4-1:0] node51778;
	wire [4-1:0] node51779;
	wire [4-1:0] node51780;
	wire [4-1:0] node51783;
	wire [4-1:0] node51786;
	wire [4-1:0] node51787;
	wire [4-1:0] node51791;
	wire [4-1:0] node51793;
	wire [4-1:0] node51796;
	wire [4-1:0] node51797;
	wire [4-1:0] node51798;
	wire [4-1:0] node51802;
	wire [4-1:0] node51804;
	wire [4-1:0] node51805;
	wire [4-1:0] node51808;
	wire [4-1:0] node51811;
	wire [4-1:0] node51812;
	wire [4-1:0] node51813;
	wire [4-1:0] node51814;
	wire [4-1:0] node51815;
	wire [4-1:0] node51818;
	wire [4-1:0] node51822;
	wire [4-1:0] node51823;
	wire [4-1:0] node51824;
	wire [4-1:0] node51829;
	wire [4-1:0] node51830;
	wire [4-1:0] node51831;
	wire [4-1:0] node51834;
	wire [4-1:0] node51838;
	wire [4-1:0] node51839;
	wire [4-1:0] node51840;
	wire [4-1:0] node51841;
	wire [4-1:0] node51842;
	wire [4-1:0] node51843;
	wire [4-1:0] node51846;
	wire [4-1:0] node51849;
	wire [4-1:0] node51851;
	wire [4-1:0] node51854;
	wire [4-1:0] node51855;
	wire [4-1:0] node51856;
	wire [4-1:0] node51857;
	wire [4-1:0] node51860;
	wire [4-1:0] node51863;
	wire [4-1:0] node51864;
	wire [4-1:0] node51868;
	wire [4-1:0] node51870;
	wire [4-1:0] node51873;
	wire [4-1:0] node51874;
	wire [4-1:0] node51876;
	wire [4-1:0] node51877;
	wire [4-1:0] node51880;
	wire [4-1:0] node51883;
	wire [4-1:0] node51884;
	wire [4-1:0] node51885;
	wire [4-1:0] node51888;
	wire [4-1:0] node51891;
	wire [4-1:0] node51892;
	wire [4-1:0] node51896;
	wire [4-1:0] node51897;
	wire [4-1:0] node51898;
	wire [4-1:0] node51899;
	wire [4-1:0] node51900;
	wire [4-1:0] node51904;
	wire [4-1:0] node51907;
	wire [4-1:0] node51908;
	wire [4-1:0] node51909;
	wire [4-1:0] node51913;
	wire [4-1:0] node51916;
	wire [4-1:0] node51917;
	wire [4-1:0] node51919;
	wire [4-1:0] node51920;
	wire [4-1:0] node51923;
	wire [4-1:0] node51926;
	wire [4-1:0] node51927;
	wire [4-1:0] node51928;
	wire [4-1:0] node51932;
	wire [4-1:0] node51935;
	wire [4-1:0] node51936;
	wire [4-1:0] node51937;
	wire [4-1:0] node51938;
	wire [4-1:0] node51939;
	wire [4-1:0] node51940;
	wire [4-1:0] node51941;
	wire [4-1:0] node51942;
	wire [4-1:0] node51943;
	wire [4-1:0] node51948;
	wire [4-1:0] node51950;
	wire [4-1:0] node51951;
	wire [4-1:0] node51954;
	wire [4-1:0] node51957;
	wire [4-1:0] node51959;
	wire [4-1:0] node51960;
	wire [4-1:0] node51961;
	wire [4-1:0] node51964;
	wire [4-1:0] node51967;
	wire [4-1:0] node51968;
	wire [4-1:0] node51971;
	wire [4-1:0] node51974;
	wire [4-1:0] node51975;
	wire [4-1:0] node51976;
	wire [4-1:0] node51977;
	wire [4-1:0] node51978;
	wire [4-1:0] node51981;
	wire [4-1:0] node51985;
	wire [4-1:0] node51986;
	wire [4-1:0] node51987;
	wire [4-1:0] node51990;
	wire [4-1:0] node51993;
	wire [4-1:0] node51996;
	wire [4-1:0] node51997;
	wire [4-1:0] node51998;
	wire [4-1:0] node51999;
	wire [4-1:0] node52002;
	wire [4-1:0] node52006;
	wire [4-1:0] node52008;
	wire [4-1:0] node52011;
	wire [4-1:0] node52012;
	wire [4-1:0] node52013;
	wire [4-1:0] node52014;
	wire [4-1:0] node52015;
	wire [4-1:0] node52016;
	wire [4-1:0] node52019;
	wire [4-1:0] node52022;
	wire [4-1:0] node52024;
	wire [4-1:0] node52027;
	wire [4-1:0] node52030;
	wire [4-1:0] node52031;
	wire [4-1:0] node52032;
	wire [4-1:0] node52035;
	wire [4-1:0] node52036;
	wire [4-1:0] node52040;
	wire [4-1:0] node52043;
	wire [4-1:0] node52044;
	wire [4-1:0] node52045;
	wire [4-1:0] node52046;
	wire [4-1:0] node52048;
	wire [4-1:0] node52051;
	wire [4-1:0] node52053;
	wire [4-1:0] node52056;
	wire [4-1:0] node52057;
	wire [4-1:0] node52059;
	wire [4-1:0] node52062;
	wire [4-1:0] node52064;
	wire [4-1:0] node52067;
	wire [4-1:0] node52068;
	wire [4-1:0] node52070;
	wire [4-1:0] node52072;
	wire [4-1:0] node52075;
	wire [4-1:0] node52076;
	wire [4-1:0] node52077;
	wire [4-1:0] node52080;
	wire [4-1:0] node52084;
	wire [4-1:0] node52085;
	wire [4-1:0] node52086;
	wire [4-1:0] node52087;
	wire [4-1:0] node52088;
	wire [4-1:0] node52090;
	wire [4-1:0] node52093;
	wire [4-1:0] node52095;
	wire [4-1:0] node52098;
	wire [4-1:0] node52100;
	wire [4-1:0] node52103;
	wire [4-1:0] node52104;
	wire [4-1:0] node52105;
	wire [4-1:0] node52106;
	wire [4-1:0] node52110;
	wire [4-1:0] node52113;
	wire [4-1:0] node52115;
	wire [4-1:0] node52118;
	wire [4-1:0] node52119;
	wire [4-1:0] node52120;
	wire [4-1:0] node52121;
	wire [4-1:0] node52122;
	wire [4-1:0] node52126;
	wire [4-1:0] node52127;
	wire [4-1:0] node52129;
	wire [4-1:0] node52132;
	wire [4-1:0] node52134;
	wire [4-1:0] node52137;
	wire [4-1:0] node52138;
	wire [4-1:0] node52139;
	wire [4-1:0] node52143;
	wire [4-1:0] node52146;
	wire [4-1:0] node52147;
	wire [4-1:0] node52148;
	wire [4-1:0] node52151;
	wire [4-1:0] node52154;
	wire [4-1:0] node52155;
	wire [4-1:0] node52157;
	wire [4-1:0] node52160;
	wire [4-1:0] node52161;
	wire [4-1:0] node52164;
	wire [4-1:0] node52166;
	wire [4-1:0] node52169;
	wire [4-1:0] node52170;
	wire [4-1:0] node52171;
	wire [4-1:0] node52172;
	wire [4-1:0] node52173;
	wire [4-1:0] node52174;
	wire [4-1:0] node52175;
	wire [4-1:0] node52178;
	wire [4-1:0] node52181;
	wire [4-1:0] node52183;
	wire [4-1:0] node52186;
	wire [4-1:0] node52187;
	wire [4-1:0] node52190;
	wire [4-1:0] node52193;
	wire [4-1:0] node52194;
	wire [4-1:0] node52195;
	wire [4-1:0] node52198;
	wire [4-1:0] node52201;
	wire [4-1:0] node52202;
	wire [4-1:0] node52204;
	wire [4-1:0] node52207;
	wire [4-1:0] node52208;
	wire [4-1:0] node52211;
	wire [4-1:0] node52214;
	wire [4-1:0] node52215;
	wire [4-1:0] node52216;
	wire [4-1:0] node52217;
	wire [4-1:0] node52219;
	wire [4-1:0] node52222;
	wire [4-1:0] node52223;
	wire [4-1:0] node52227;
	wire [4-1:0] node52228;
	wire [4-1:0] node52231;
	wire [4-1:0] node52234;
	wire [4-1:0] node52235;
	wire [4-1:0] node52236;
	wire [4-1:0] node52239;
	wire [4-1:0] node52242;
	wire [4-1:0] node52243;
	wire [4-1:0] node52246;
	wire [4-1:0] node52249;
	wire [4-1:0] node52250;
	wire [4-1:0] node52251;
	wire [4-1:0] node52252;
	wire [4-1:0] node52253;
	wire [4-1:0] node52254;
	wire [4-1:0] node52257;
	wire [4-1:0] node52260;
	wire [4-1:0] node52261;
	wire [4-1:0] node52264;
	wire [4-1:0] node52267;
	wire [4-1:0] node52268;
	wire [4-1:0] node52271;
	wire [4-1:0] node52274;
	wire [4-1:0] node52275;
	wire [4-1:0] node52276;
	wire [4-1:0] node52279;
	wire [4-1:0] node52282;
	wire [4-1:0] node52283;
	wire [4-1:0] node52286;
	wire [4-1:0] node52289;
	wire [4-1:0] node52290;
	wire [4-1:0] node52291;
	wire [4-1:0] node52292;
	wire [4-1:0] node52293;
	wire [4-1:0] node52297;
	wire [4-1:0] node52300;
	wire [4-1:0] node52301;
	wire [4-1:0] node52302;
	wire [4-1:0] node52306;
	wire [4-1:0] node52309;
	wire [4-1:0] node52310;
	wire [4-1:0] node52311;
	wire [4-1:0] node52312;
	wire [4-1:0] node52316;
	wire [4-1:0] node52319;
	wire [4-1:0] node52320;
	wire [4-1:0] node52321;
	wire [4-1:0] node52325;
	wire [4-1:0] node52328;
	wire [4-1:0] node52329;
	wire [4-1:0] node52330;
	wire [4-1:0] node52331;
	wire [4-1:0] node52332;
	wire [4-1:0] node52333;
	wire [4-1:0] node52334;
	wire [4-1:0] node52335;
	wire [4-1:0] node52337;
	wire [4-1:0] node52339;
	wire [4-1:0] node52342;
	wire [4-1:0] node52343;
	wire [4-1:0] node52347;
	wire [4-1:0] node52348;
	wire [4-1:0] node52351;
	wire [4-1:0] node52354;
	wire [4-1:0] node52355;
	wire [4-1:0] node52356;
	wire [4-1:0] node52357;
	wire [4-1:0] node52358;
	wire [4-1:0] node52362;
	wire [4-1:0] node52363;
	wire [4-1:0] node52367;
	wire [4-1:0] node52369;
	wire [4-1:0] node52370;
	wire [4-1:0] node52373;
	wire [4-1:0] node52376;
	wire [4-1:0] node52377;
	wire [4-1:0] node52379;
	wire [4-1:0] node52382;
	wire [4-1:0] node52383;
	wire [4-1:0] node52384;
	wire [4-1:0] node52387;
	wire [4-1:0] node52390;
	wire [4-1:0] node52392;
	wire [4-1:0] node52395;
	wire [4-1:0] node52396;
	wire [4-1:0] node52397;
	wire [4-1:0] node52398;
	wire [4-1:0] node52399;
	wire [4-1:0] node52403;
	wire [4-1:0] node52405;
	wire [4-1:0] node52408;
	wire [4-1:0] node52409;
	wire [4-1:0] node52411;
	wire [4-1:0] node52412;
	wire [4-1:0] node52415;
	wire [4-1:0] node52418;
	wire [4-1:0] node52419;
	wire [4-1:0] node52422;
	wire [4-1:0] node52425;
	wire [4-1:0] node52426;
	wire [4-1:0] node52428;
	wire [4-1:0] node52429;
	wire [4-1:0] node52431;
	wire [4-1:0] node52435;
	wire [4-1:0] node52436;
	wire [4-1:0] node52439;
	wire [4-1:0] node52440;
	wire [4-1:0] node52441;
	wire [4-1:0] node52444;
	wire [4-1:0] node52448;
	wire [4-1:0] node52449;
	wire [4-1:0] node52450;
	wire [4-1:0] node52451;
	wire [4-1:0] node52452;
	wire [4-1:0] node52455;
	wire [4-1:0] node52456;
	wire [4-1:0] node52459;
	wire [4-1:0] node52462;
	wire [4-1:0] node52463;
	wire [4-1:0] node52464;
	wire [4-1:0] node52468;
	wire [4-1:0] node52471;
	wire [4-1:0] node52472;
	wire [4-1:0] node52473;
	wire [4-1:0] node52475;
	wire [4-1:0] node52476;
	wire [4-1:0] node52480;
	wire [4-1:0] node52482;
	wire [4-1:0] node52485;
	wire [4-1:0] node52486;
	wire [4-1:0] node52487;
	wire [4-1:0] node52490;
	wire [4-1:0] node52493;
	wire [4-1:0] node52494;
	wire [4-1:0] node52497;
	wire [4-1:0] node52500;
	wire [4-1:0] node52501;
	wire [4-1:0] node52502;
	wire [4-1:0] node52503;
	wire [4-1:0] node52504;
	wire [4-1:0] node52505;
	wire [4-1:0] node52509;
	wire [4-1:0] node52512;
	wire [4-1:0] node52513;
	wire [4-1:0] node52517;
	wire [4-1:0] node52518;
	wire [4-1:0] node52519;
	wire [4-1:0] node52523;
	wire [4-1:0] node52526;
	wire [4-1:0] node52527;
	wire [4-1:0] node52528;
	wire [4-1:0] node52529;
	wire [4-1:0] node52532;
	wire [4-1:0] node52535;
	wire [4-1:0] node52536;
	wire [4-1:0] node52539;
	wire [4-1:0] node52540;
	wire [4-1:0] node52544;
	wire [4-1:0] node52545;
	wire [4-1:0] node52548;
	wire [4-1:0] node52550;
	wire [4-1:0] node52553;
	wire [4-1:0] node52554;
	wire [4-1:0] node52555;
	wire [4-1:0] node52556;
	wire [4-1:0] node52557;
	wire [4-1:0] node52560;
	wire [4-1:0] node52563;
	wire [4-1:0] node52564;
	wire [4-1:0] node52566;
	wire [4-1:0] node52567;
	wire [4-1:0] node52571;
	wire [4-1:0] node52572;
	wire [4-1:0] node52575;
	wire [4-1:0] node52578;
	wire [4-1:0] node52579;
	wire [4-1:0] node52580;
	wire [4-1:0] node52582;
	wire [4-1:0] node52584;
	wire [4-1:0] node52587;
	wire [4-1:0] node52588;
	wire [4-1:0] node52589;
	wire [4-1:0] node52590;
	wire [4-1:0] node52595;
	wire [4-1:0] node52596;
	wire [4-1:0] node52600;
	wire [4-1:0] node52601;
	wire [4-1:0] node52602;
	wire [4-1:0] node52603;
	wire [4-1:0] node52604;
	wire [4-1:0] node52607;
	wire [4-1:0] node52610;
	wire [4-1:0] node52612;
	wire [4-1:0] node52615;
	wire [4-1:0] node52616;
	wire [4-1:0] node52620;
	wire [4-1:0] node52621;
	wire [4-1:0] node52622;
	wire [4-1:0] node52626;
	wire [4-1:0] node52627;
	wire [4-1:0] node52630;
	wire [4-1:0] node52633;
	wire [4-1:0] node52634;
	wire [4-1:0] node52635;
	wire [4-1:0] node52636;
	wire [4-1:0] node52637;
	wire [4-1:0] node52641;
	wire [4-1:0] node52642;
	wire [4-1:0] node52646;
	wire [4-1:0] node52647;
	wire [4-1:0] node52648;
	wire [4-1:0] node52652;
	wire [4-1:0] node52653;
	wire [4-1:0] node52657;
	wire [4-1:0] node52658;
	wire [4-1:0] node52659;
	wire [4-1:0] node52660;
	wire [4-1:0] node52661;
	wire [4-1:0] node52665;
	wire [4-1:0] node52666;
	wire [4-1:0] node52669;
	wire [4-1:0] node52672;
	wire [4-1:0] node52673;
	wire [4-1:0] node52675;
	wire [4-1:0] node52678;
	wire [4-1:0] node52679;
	wire [4-1:0] node52680;
	wire [4-1:0] node52683;
	wire [4-1:0] node52687;
	wire [4-1:0] node52688;
	wire [4-1:0] node52689;
	wire [4-1:0] node52690;
	wire [4-1:0] node52691;
	wire [4-1:0] node52694;
	wire [4-1:0] node52698;
	wire [4-1:0] node52700;
	wire [4-1:0] node52701;
	wire [4-1:0] node52704;
	wire [4-1:0] node52707;
	wire [4-1:0] node52708;
	wire [4-1:0] node52709;
	wire [4-1:0] node52712;
	wire [4-1:0] node52714;
	wire [4-1:0] node52717;
	wire [4-1:0] node52718;
	wire [4-1:0] node52721;
	wire [4-1:0] node52724;
	wire [4-1:0] node52725;
	wire [4-1:0] node52726;
	wire [4-1:0] node52727;
	wire [4-1:0] node52728;
	wire [4-1:0] node52729;
	wire [4-1:0] node52730;
	wire [4-1:0] node52732;
	wire [4-1:0] node52735;
	wire [4-1:0] node52737;
	wire [4-1:0] node52740;
	wire [4-1:0] node52741;
	wire [4-1:0] node52743;
	wire [4-1:0] node52745;
	wire [4-1:0] node52749;
	wire [4-1:0] node52750;
	wire [4-1:0] node52751;
	wire [4-1:0] node52753;
	wire [4-1:0] node52756;
	wire [4-1:0] node52758;
	wire [4-1:0] node52761;
	wire [4-1:0] node52762;
	wire [4-1:0] node52763;
	wire [4-1:0] node52765;
	wire [4-1:0] node52769;
	wire [4-1:0] node52770;
	wire [4-1:0] node52772;
	wire [4-1:0] node52775;
	wire [4-1:0] node52776;
	wire [4-1:0] node52780;
	wire [4-1:0] node52781;
	wire [4-1:0] node52782;
	wire [4-1:0] node52783;
	wire [4-1:0] node52785;
	wire [4-1:0] node52786;
	wire [4-1:0] node52789;
	wire [4-1:0] node52792;
	wire [4-1:0] node52795;
	wire [4-1:0] node52796;
	wire [4-1:0] node52797;
	wire [4-1:0] node52798;
	wire [4-1:0] node52802;
	wire [4-1:0] node52803;
	wire [4-1:0] node52807;
	wire [4-1:0] node52808;
	wire [4-1:0] node52809;
	wire [4-1:0] node52812;
	wire [4-1:0] node52816;
	wire [4-1:0] node52817;
	wire [4-1:0] node52818;
	wire [4-1:0] node52819;
	wire [4-1:0] node52820;
	wire [4-1:0] node52825;
	wire [4-1:0] node52826;
	wire [4-1:0] node52827;
	wire [4-1:0] node52830;
	wire [4-1:0] node52834;
	wire [4-1:0] node52835;
	wire [4-1:0] node52836;
	wire [4-1:0] node52839;
	wire [4-1:0] node52842;
	wire [4-1:0] node52845;
	wire [4-1:0] node52846;
	wire [4-1:0] node52847;
	wire [4-1:0] node52848;
	wire [4-1:0] node52849;
	wire [4-1:0] node52850;
	wire [4-1:0] node52854;
	wire [4-1:0] node52855;
	wire [4-1:0] node52858;
	wire [4-1:0] node52861;
	wire [4-1:0] node52862;
	wire [4-1:0] node52863;
	wire [4-1:0] node52867;
	wire [4-1:0] node52868;
	wire [4-1:0] node52871;
	wire [4-1:0] node52872;
	wire [4-1:0] node52876;
	wire [4-1:0] node52877;
	wire [4-1:0] node52878;
	wire [4-1:0] node52879;
	wire [4-1:0] node52880;
	wire [4-1:0] node52883;
	wire [4-1:0] node52887;
	wire [4-1:0] node52888;
	wire [4-1:0] node52889;
	wire [4-1:0] node52893;
	wire [4-1:0] node52896;
	wire [4-1:0] node52897;
	wire [4-1:0] node52898;
	wire [4-1:0] node52900;
	wire [4-1:0] node52904;
	wire [4-1:0] node52905;
	wire [4-1:0] node52909;
	wire [4-1:0] node52910;
	wire [4-1:0] node52911;
	wire [4-1:0] node52912;
	wire [4-1:0] node52913;
	wire [4-1:0] node52917;
	wire [4-1:0] node52918;
	wire [4-1:0] node52919;
	wire [4-1:0] node52924;
	wire [4-1:0] node52925;
	wire [4-1:0] node52928;
	wire [4-1:0] node52929;
	wire [4-1:0] node52930;
	wire [4-1:0] node52934;
	wire [4-1:0] node52937;
	wire [4-1:0] node52938;
	wire [4-1:0] node52939;
	wire [4-1:0] node52940;
	wire [4-1:0] node52943;
	wire [4-1:0] node52946;
	wire [4-1:0] node52947;
	wire [4-1:0] node52950;
	wire [4-1:0] node52953;
	wire [4-1:0] node52954;
	wire [4-1:0] node52955;
	wire [4-1:0] node52957;
	wire [4-1:0] node52960;
	wire [4-1:0] node52962;
	wire [4-1:0] node52965;
	wire [4-1:0] node52966;
	wire [4-1:0] node52967;
	wire [4-1:0] node52971;
	wire [4-1:0] node52974;
	wire [4-1:0] node52975;
	wire [4-1:0] node52976;
	wire [4-1:0] node52977;
	wire [4-1:0] node52978;
	wire [4-1:0] node52979;
	wire [4-1:0] node52982;
	wire [4-1:0] node52984;
	wire [4-1:0] node52987;
	wire [4-1:0] node52988;
	wire [4-1:0] node52991;
	wire [4-1:0] node52993;
	wire [4-1:0] node52996;
	wire [4-1:0] node52997;
	wire [4-1:0] node52999;
	wire [4-1:0] node53001;
	wire [4-1:0] node53004;
	wire [4-1:0] node53005;
	wire [4-1:0] node53007;
	wire [4-1:0] node53010;
	wire [4-1:0] node53013;
	wire [4-1:0] node53014;
	wire [4-1:0] node53015;
	wire [4-1:0] node53016;
	wire [4-1:0] node53017;
	wire [4-1:0] node53021;
	wire [4-1:0] node53022;
	wire [4-1:0] node53023;
	wire [4-1:0] node53026;
	wire [4-1:0] node53029;
	wire [4-1:0] node53031;
	wire [4-1:0] node53034;
	wire [4-1:0] node53035;
	wire [4-1:0] node53037;
	wire [4-1:0] node53038;
	wire [4-1:0] node53041;
	wire [4-1:0] node53044;
	wire [4-1:0] node53045;
	wire [4-1:0] node53047;
	wire [4-1:0] node53051;
	wire [4-1:0] node53052;
	wire [4-1:0] node53053;
	wire [4-1:0] node53054;
	wire [4-1:0] node53055;
	wire [4-1:0] node53060;
	wire [4-1:0] node53061;
	wire [4-1:0] node53065;
	wire [4-1:0] node53066;
	wire [4-1:0] node53067;
	wire [4-1:0] node53070;
	wire [4-1:0] node53073;
	wire [4-1:0] node53074;
	wire [4-1:0] node53077;
	wire [4-1:0] node53080;
	wire [4-1:0] node53081;
	wire [4-1:0] node53082;
	wire [4-1:0] node53083;
	wire [4-1:0] node53084;
	wire [4-1:0] node53086;
	wire [4-1:0] node53089;
	wire [4-1:0] node53090;
	wire [4-1:0] node53094;
	wire [4-1:0] node53095;
	wire [4-1:0] node53096;
	wire [4-1:0] node53099;
	wire [4-1:0] node53102;
	wire [4-1:0] node53103;
	wire [4-1:0] node53106;
	wire [4-1:0] node53109;
	wire [4-1:0] node53110;
	wire [4-1:0] node53111;
	wire [4-1:0] node53115;
	wire [4-1:0] node53117;
	wire [4-1:0] node53120;
	wire [4-1:0] node53121;
	wire [4-1:0] node53122;
	wire [4-1:0] node53123;
	wire [4-1:0] node53124;
	wire [4-1:0] node53127;
	wire [4-1:0] node53130;
	wire [4-1:0] node53131;
	wire [4-1:0] node53132;
	wire [4-1:0] node53135;
	wire [4-1:0] node53138;
	wire [4-1:0] node53139;
	wire [4-1:0] node53142;
	wire [4-1:0] node53145;
	wire [4-1:0] node53146;
	wire [4-1:0] node53149;
	wire [4-1:0] node53152;
	wire [4-1:0] node53153;
	wire [4-1:0] node53154;
	wire [4-1:0] node53156;
	wire [4-1:0] node53157;
	wire [4-1:0] node53160;
	wire [4-1:0] node53163;
	wire [4-1:0] node53164;
	wire [4-1:0] node53165;
	wire [4-1:0] node53168;
	wire [4-1:0] node53172;
	wire [4-1:0] node53173;
	wire [4-1:0] node53176;
	wire [4-1:0] node53179;
	wire [4-1:0] node53180;
	wire [4-1:0] node53181;
	wire [4-1:0] node53182;
	wire [4-1:0] node53183;
	wire [4-1:0] node53184;
	wire [4-1:0] node53185;
	wire [4-1:0] node53186;
	wire [4-1:0] node53187;
	wire [4-1:0] node53190;
	wire [4-1:0] node53191;
	wire [4-1:0] node53195;
	wire [4-1:0] node53196;
	wire [4-1:0] node53200;
	wire [4-1:0] node53201;
	wire [4-1:0] node53203;
	wire [4-1:0] node53204;
	wire [4-1:0] node53207;
	wire [4-1:0] node53210;
	wire [4-1:0] node53211;
	wire [4-1:0] node53214;
	wire [4-1:0] node53217;
	wire [4-1:0] node53218;
	wire [4-1:0] node53219;
	wire [4-1:0] node53220;
	wire [4-1:0] node53221;
	wire [4-1:0] node53222;
	wire [4-1:0] node53226;
	wire [4-1:0] node53230;
	wire [4-1:0] node53231;
	wire [4-1:0] node53232;
	wire [4-1:0] node53236;
	wire [4-1:0] node53239;
	wire [4-1:0] node53240;
	wire [4-1:0] node53241;
	wire [4-1:0] node53242;
	wire [4-1:0] node53246;
	wire [4-1:0] node53247;
	wire [4-1:0] node53248;
	wire [4-1:0] node53251;
	wire [4-1:0] node53254;
	wire [4-1:0] node53255;
	wire [4-1:0] node53258;
	wire [4-1:0] node53261;
	wire [4-1:0] node53262;
	wire [4-1:0] node53263;
	wire [4-1:0] node53266;
	wire [4-1:0] node53269;
	wire [4-1:0] node53270;
	wire [4-1:0] node53273;
	wire [4-1:0] node53276;
	wire [4-1:0] node53277;
	wire [4-1:0] node53278;
	wire [4-1:0] node53279;
	wire [4-1:0] node53280;
	wire [4-1:0] node53281;
	wire [4-1:0] node53282;
	wire [4-1:0] node53285;
	wire [4-1:0] node53288;
	wire [4-1:0] node53289;
	wire [4-1:0] node53292;
	wire [4-1:0] node53295;
	wire [4-1:0] node53296;
	wire [4-1:0] node53298;
	wire [4-1:0] node53301;
	wire [4-1:0] node53304;
	wire [4-1:0] node53305;
	wire [4-1:0] node53306;
	wire [4-1:0] node53309;
	wire [4-1:0] node53312;
	wire [4-1:0] node53313;
	wire [4-1:0] node53317;
	wire [4-1:0] node53318;
	wire [4-1:0] node53319;
	wire [4-1:0] node53320;
	wire [4-1:0] node53323;
	wire [4-1:0] node53326;
	wire [4-1:0] node53329;
	wire [4-1:0] node53330;
	wire [4-1:0] node53332;
	wire [4-1:0] node53333;
	wire [4-1:0] node53336;
	wire [4-1:0] node53339;
	wire [4-1:0] node53341;
	wire [4-1:0] node53344;
	wire [4-1:0] node53345;
	wire [4-1:0] node53346;
	wire [4-1:0] node53347;
	wire [4-1:0] node53348;
	wire [4-1:0] node53350;
	wire [4-1:0] node53354;
	wire [4-1:0] node53355;
	wire [4-1:0] node53356;
	wire [4-1:0] node53360;
	wire [4-1:0] node53361;
	wire [4-1:0] node53364;
	wire [4-1:0] node53367;
	wire [4-1:0] node53368;
	wire [4-1:0] node53369;
	wire [4-1:0] node53373;
	wire [4-1:0] node53375;
	wire [4-1:0] node53378;
	wire [4-1:0] node53379;
	wire [4-1:0] node53380;
	wire [4-1:0] node53381;
	wire [4-1:0] node53382;
	wire [4-1:0] node53386;
	wire [4-1:0] node53388;
	wire [4-1:0] node53391;
	wire [4-1:0] node53392;
	wire [4-1:0] node53395;
	wire [4-1:0] node53398;
	wire [4-1:0] node53399;
	wire [4-1:0] node53400;
	wire [4-1:0] node53403;
	wire [4-1:0] node53406;
	wire [4-1:0] node53409;
	wire [4-1:0] node53410;
	wire [4-1:0] node53411;
	wire [4-1:0] node53412;
	wire [4-1:0] node53413;
	wire [4-1:0] node53414;
	wire [4-1:0] node53415;
	wire [4-1:0] node53416;
	wire [4-1:0] node53420;
	wire [4-1:0] node53421;
	wire [4-1:0] node53424;
	wire [4-1:0] node53427;
	wire [4-1:0] node53428;
	wire [4-1:0] node53432;
	wire [4-1:0] node53433;
	wire [4-1:0] node53435;
	wire [4-1:0] node53438;
	wire [4-1:0] node53440;
	wire [4-1:0] node53443;
	wire [4-1:0] node53444;
	wire [4-1:0] node53445;
	wire [4-1:0] node53446;
	wire [4-1:0] node53447;
	wire [4-1:0] node53450;
	wire [4-1:0] node53453;
	wire [4-1:0] node53454;
	wire [4-1:0] node53458;
	wire [4-1:0] node53460;
	wire [4-1:0] node53461;
	wire [4-1:0] node53464;
	wire [4-1:0] node53467;
	wire [4-1:0] node53468;
	wire [4-1:0] node53470;
	wire [4-1:0] node53473;
	wire [4-1:0] node53474;
	wire [4-1:0] node53478;
	wire [4-1:0] node53479;
	wire [4-1:0] node53480;
	wire [4-1:0] node53481;
	wire [4-1:0] node53483;
	wire [4-1:0] node53486;
	wire [4-1:0] node53487;
	wire [4-1:0] node53488;
	wire [4-1:0] node53493;
	wire [4-1:0] node53494;
	wire [4-1:0] node53495;
	wire [4-1:0] node53496;
	wire [4-1:0] node53499;
	wire [4-1:0] node53502;
	wire [4-1:0] node53504;
	wire [4-1:0] node53507;
	wire [4-1:0] node53509;
	wire [4-1:0] node53512;
	wire [4-1:0] node53513;
	wire [4-1:0] node53514;
	wire [4-1:0] node53517;
	wire [4-1:0] node53518;
	wire [4-1:0] node53521;
	wire [4-1:0] node53524;
	wire [4-1:0] node53526;
	wire [4-1:0] node53528;
	wire [4-1:0] node53531;
	wire [4-1:0] node53532;
	wire [4-1:0] node53533;
	wire [4-1:0] node53534;
	wire [4-1:0] node53536;
	wire [4-1:0] node53537;
	wire [4-1:0] node53540;
	wire [4-1:0] node53543;
	wire [4-1:0] node53544;
	wire [4-1:0] node53545;
	wire [4-1:0] node53549;
	wire [4-1:0] node53550;
	wire [4-1:0] node53553;
	wire [4-1:0] node53555;
	wire [4-1:0] node53558;
	wire [4-1:0] node53559;
	wire [4-1:0] node53560;
	wire [4-1:0] node53561;
	wire [4-1:0] node53564;
	wire [4-1:0] node53567;
	wire [4-1:0] node53568;
	wire [4-1:0] node53569;
	wire [4-1:0] node53572;
	wire [4-1:0] node53575;
	wire [4-1:0] node53576;
	wire [4-1:0] node53580;
	wire [4-1:0] node53582;
	wire [4-1:0] node53585;
	wire [4-1:0] node53586;
	wire [4-1:0] node53587;
	wire [4-1:0] node53588;
	wire [4-1:0] node53590;
	wire [4-1:0] node53592;
	wire [4-1:0] node53595;
	wire [4-1:0] node53596;
	wire [4-1:0] node53599;
	wire [4-1:0] node53602;
	wire [4-1:0] node53603;
	wire [4-1:0] node53604;
	wire [4-1:0] node53607;
	wire [4-1:0] node53610;
	wire [4-1:0] node53611;
	wire [4-1:0] node53613;
	wire [4-1:0] node53617;
	wire [4-1:0] node53618;
	wire [4-1:0] node53620;
	wire [4-1:0] node53621;
	wire [4-1:0] node53622;
	wire [4-1:0] node53625;
	wire [4-1:0] node53629;
	wire [4-1:0] node53630;
	wire [4-1:0] node53633;
	wire [4-1:0] node53634;
	wire [4-1:0] node53637;
	wire [4-1:0] node53640;
	wire [4-1:0] node53641;
	wire [4-1:0] node53642;
	wire [4-1:0] node53643;
	wire [4-1:0] node53644;
	wire [4-1:0] node53645;
	wire [4-1:0] node53646;
	wire [4-1:0] node53647;
	wire [4-1:0] node53651;
	wire [4-1:0] node53652;
	wire [4-1:0] node53656;
	wire [4-1:0] node53657;
	wire [4-1:0] node53658;
	wire [4-1:0] node53662;
	wire [4-1:0] node53663;
	wire [4-1:0] node53667;
	wire [4-1:0] node53668;
	wire [4-1:0] node53669;
	wire [4-1:0] node53670;
	wire [4-1:0] node53671;
	wire [4-1:0] node53676;
	wire [4-1:0] node53678;
	wire [4-1:0] node53681;
	wire [4-1:0] node53682;
	wire [4-1:0] node53685;
	wire [4-1:0] node53688;
	wire [4-1:0] node53689;
	wire [4-1:0] node53690;
	wire [4-1:0] node53691;
	wire [4-1:0] node53693;
	wire [4-1:0] node53696;
	wire [4-1:0] node53698;
	wire [4-1:0] node53701;
	wire [4-1:0] node53702;
	wire [4-1:0] node53705;
	wire [4-1:0] node53708;
	wire [4-1:0] node53709;
	wire [4-1:0] node53712;
	wire [4-1:0] node53715;
	wire [4-1:0] node53716;
	wire [4-1:0] node53717;
	wire [4-1:0] node53718;
	wire [4-1:0] node53719;
	wire [4-1:0] node53722;
	wire [4-1:0] node53723;
	wire [4-1:0] node53727;
	wire [4-1:0] node53728;
	wire [4-1:0] node53729;
	wire [4-1:0] node53733;
	wire [4-1:0] node53734;
	wire [4-1:0] node53738;
	wire [4-1:0] node53739;
	wire [4-1:0] node53740;
	wire [4-1:0] node53741;
	wire [4-1:0] node53742;
	wire [4-1:0] node53745;
	wire [4-1:0] node53749;
	wire [4-1:0] node53750;
	wire [4-1:0] node53754;
	wire [4-1:0] node53755;
	wire [4-1:0] node53758;
	wire [4-1:0] node53761;
	wire [4-1:0] node53762;
	wire [4-1:0] node53763;
	wire [4-1:0] node53764;
	wire [4-1:0] node53768;
	wire [4-1:0] node53769;
	wire [4-1:0] node53773;
	wire [4-1:0] node53774;
	wire [4-1:0] node53775;
	wire [4-1:0] node53779;
	wire [4-1:0] node53780;
	wire [4-1:0] node53784;
	wire [4-1:0] node53785;
	wire [4-1:0] node53786;
	wire [4-1:0] node53787;
	wire [4-1:0] node53788;
	wire [4-1:0] node53789;
	wire [4-1:0] node53791;
	wire [4-1:0] node53794;
	wire [4-1:0] node53795;
	wire [4-1:0] node53796;
	wire [4-1:0] node53800;
	wire [4-1:0] node53801;
	wire [4-1:0] node53805;
	wire [4-1:0] node53806;
	wire [4-1:0] node53807;
	wire [4-1:0] node53808;
	wire [4-1:0] node53811;
	wire [4-1:0] node53814;
	wire [4-1:0] node53816;
	wire [4-1:0] node53819;
	wire [4-1:0] node53821;
	wire [4-1:0] node53824;
	wire [4-1:0] node53825;
	wire [4-1:0] node53826;
	wire [4-1:0] node53827;
	wire [4-1:0] node53831;
	wire [4-1:0] node53832;
	wire [4-1:0] node53833;
	wire [4-1:0] node53838;
	wire [4-1:0] node53839;
	wire [4-1:0] node53840;
	wire [4-1:0] node53841;
	wire [4-1:0] node53844;
	wire [4-1:0] node53847;
	wire [4-1:0] node53848;
	wire [4-1:0] node53851;
	wire [4-1:0] node53854;
	wire [4-1:0] node53855;
	wire [4-1:0] node53859;
	wire [4-1:0] node53860;
	wire [4-1:0] node53861;
	wire [4-1:0] node53862;
	wire [4-1:0] node53865;
	wire [4-1:0] node53868;
	wire [4-1:0] node53869;
	wire [4-1:0] node53870;
	wire [4-1:0] node53874;
	wire [4-1:0] node53875;
	wire [4-1:0] node53879;
	wire [4-1:0] node53880;
	wire [4-1:0] node53883;
	wire [4-1:0] node53886;
	wire [4-1:0] node53887;
	wire [4-1:0] node53888;
	wire [4-1:0] node53889;
	wire [4-1:0] node53890;
	wire [4-1:0] node53893;
	wire [4-1:0] node53894;
	wire [4-1:0] node53895;
	wire [4-1:0] node53898;
	wire [4-1:0] node53901;
	wire [4-1:0] node53902;
	wire [4-1:0] node53906;
	wire [4-1:0] node53907;
	wire [4-1:0] node53908;
	wire [4-1:0] node53912;
	wire [4-1:0] node53913;
	wire [4-1:0] node53916;
	wire [4-1:0] node53919;
	wire [4-1:0] node53920;
	wire [4-1:0] node53921;
	wire [4-1:0] node53922;
	wire [4-1:0] node53926;
	wire [4-1:0] node53927;
	wire [4-1:0] node53930;
	wire [4-1:0] node53933;
	wire [4-1:0] node53934;
	wire [4-1:0] node53937;
	wire [4-1:0] node53940;
	wire [4-1:0] node53941;
	wire [4-1:0] node53942;
	wire [4-1:0] node53943;
	wire [4-1:0] node53944;
	wire [4-1:0] node53945;
	wire [4-1:0] node53949;
	wire [4-1:0] node53950;
	wire [4-1:0] node53953;
	wire [4-1:0] node53957;
	wire [4-1:0] node53958;
	wire [4-1:0] node53960;
	wire [4-1:0] node53963;
	wire [4-1:0] node53964;
	wire [4-1:0] node53967;
	wire [4-1:0] node53970;
	wire [4-1:0] node53971;
	wire [4-1:0] node53974;
	wire [4-1:0] node53977;
	wire [4-1:0] node53978;
	wire [4-1:0] node53979;
	wire [4-1:0] node53980;
	wire [4-1:0] node53981;
	wire [4-1:0] node53982;
	wire [4-1:0] node53983;
	wire [4-1:0] node53984;
	wire [4-1:0] node53985;
	wire [4-1:0] node53986;
	wire [4-1:0] node53990;
	wire [4-1:0] node53991;
	wire [4-1:0] node53994;
	wire [4-1:0] node53997;
	wire [4-1:0] node53998;
	wire [4-1:0] node54000;
	wire [4-1:0] node54003;
	wire [4-1:0] node54004;
	wire [4-1:0] node54008;
	wire [4-1:0] node54010;
	wire [4-1:0] node54011;
	wire [4-1:0] node54015;
	wire [4-1:0] node54016;
	wire [4-1:0] node54018;
	wire [4-1:0] node54019;
	wire [4-1:0] node54020;
	wire [4-1:0] node54024;
	wire [4-1:0] node54027;
	wire [4-1:0] node54029;
	wire [4-1:0] node54030;
	wire [4-1:0] node54031;
	wire [4-1:0] node54036;
	wire [4-1:0] node54037;
	wire [4-1:0] node54038;
	wire [4-1:0] node54039;
	wire [4-1:0] node54041;
	wire [4-1:0] node54042;
	wire [4-1:0] node54045;
	wire [4-1:0] node54048;
	wire [4-1:0] node54050;
	wire [4-1:0] node54053;
	wire [4-1:0] node54054;
	wire [4-1:0] node54055;
	wire [4-1:0] node54056;
	wire [4-1:0] node54059;
	wire [4-1:0] node54062;
	wire [4-1:0] node54063;
	wire [4-1:0] node54066;
	wire [4-1:0] node54069;
	wire [4-1:0] node54070;
	wire [4-1:0] node54073;
	wire [4-1:0] node54076;
	wire [4-1:0] node54077;
	wire [4-1:0] node54078;
	wire [4-1:0] node54079;
	wire [4-1:0] node54084;
	wire [4-1:0] node54085;
	wire [4-1:0] node54086;
	wire [4-1:0] node54091;
	wire [4-1:0] node54092;
	wire [4-1:0] node54093;
	wire [4-1:0] node54094;
	wire [4-1:0] node54095;
	wire [4-1:0] node54096;
	wire [4-1:0] node54100;
	wire [4-1:0] node54101;
	wire [4-1:0] node54102;
	wire [4-1:0] node54107;
	wire [4-1:0] node54108;
	wire [4-1:0] node54109;
	wire [4-1:0] node54110;
	wire [4-1:0] node54113;
	wire [4-1:0] node54116;
	wire [4-1:0] node54117;
	wire [4-1:0] node54121;
	wire [4-1:0] node54123;
	wire [4-1:0] node54126;
	wire [4-1:0] node54127;
	wire [4-1:0] node54128;
	wire [4-1:0] node54129;
	wire [4-1:0] node54130;
	wire [4-1:0] node54133;
	wire [4-1:0] node54136;
	wire [4-1:0] node54138;
	wire [4-1:0] node54141;
	wire [4-1:0] node54142;
	wire [4-1:0] node54146;
	wire [4-1:0] node54147;
	wire [4-1:0] node54148;
	wire [4-1:0] node54150;
	wire [4-1:0] node54153;
	wire [4-1:0] node54154;
	wire [4-1:0] node54157;
	wire [4-1:0] node54160;
	wire [4-1:0] node54161;
	wire [4-1:0] node54164;
	wire [4-1:0] node54167;
	wire [4-1:0] node54168;
	wire [4-1:0] node54169;
	wire [4-1:0] node54170;
	wire [4-1:0] node54171;
	wire [4-1:0] node54172;
	wire [4-1:0] node54178;
	wire [4-1:0] node54180;
	wire [4-1:0] node54182;
	wire [4-1:0] node54183;
	wire [4-1:0] node54186;
	wire [4-1:0] node54189;
	wire [4-1:0] node54190;
	wire [4-1:0] node54191;
	wire [4-1:0] node54192;
	wire [4-1:0] node54195;
	wire [4-1:0] node54198;
	wire [4-1:0] node54199;
	wire [4-1:0] node54203;
	wire [4-1:0] node54204;
	wire [4-1:0] node54207;
	wire [4-1:0] node54210;
	wire [4-1:0] node54211;
	wire [4-1:0] node54212;
	wire [4-1:0] node54213;
	wire [4-1:0] node54214;
	wire [4-1:0] node54215;
	wire [4-1:0] node54216;
	wire [4-1:0] node54217;
	wire [4-1:0] node54220;
	wire [4-1:0] node54225;
	wire [4-1:0] node54226;
	wire [4-1:0] node54227;
	wire [4-1:0] node54228;
	wire [4-1:0] node54233;
	wire [4-1:0] node54234;
	wire [4-1:0] node54235;
	wire [4-1:0] node54238;
	wire [4-1:0] node54242;
	wire [4-1:0] node54243;
	wire [4-1:0] node54245;
	wire [4-1:0] node54248;
	wire [4-1:0] node54249;
	wire [4-1:0] node54250;
	wire [4-1:0] node54252;
	wire [4-1:0] node54255;
	wire [4-1:0] node54257;
	wire [4-1:0] node54260;
	wire [4-1:0] node54262;
	wire [4-1:0] node54263;
	wire [4-1:0] node54266;
	wire [4-1:0] node54269;
	wire [4-1:0] node54270;
	wire [4-1:0] node54271;
	wire [4-1:0] node54272;
	wire [4-1:0] node54275;
	wire [4-1:0] node54276;
	wire [4-1:0] node54279;
	wire [4-1:0] node54282;
	wire [4-1:0] node54284;
	wire [4-1:0] node54285;
	wire [4-1:0] node54286;
	wire [4-1:0] node54290;
	wire [4-1:0] node54291;
	wire [4-1:0] node54295;
	wire [4-1:0] node54296;
	wire [4-1:0] node54297;
	wire [4-1:0] node54300;
	wire [4-1:0] node54303;
	wire [4-1:0] node54304;
	wire [4-1:0] node54306;
	wire [4-1:0] node54309;
	wire [4-1:0] node54310;
	wire [4-1:0] node54313;
	wire [4-1:0] node54316;
	wire [4-1:0] node54317;
	wire [4-1:0] node54318;
	wire [4-1:0] node54319;
	wire [4-1:0] node54320;
	wire [4-1:0] node54321;
	wire [4-1:0] node54325;
	wire [4-1:0] node54326;
	wire [4-1:0] node54330;
	wire [4-1:0] node54331;
	wire [4-1:0] node54335;
	wire [4-1:0] node54336;
	wire [4-1:0] node54337;
	wire [4-1:0] node54338;
	wire [4-1:0] node54339;
	wire [4-1:0] node54343;
	wire [4-1:0] node54346;
	wire [4-1:0] node54349;
	wire [4-1:0] node54350;
	wire [4-1:0] node54351;
	wire [4-1:0] node54353;
	wire [4-1:0] node54357;
	wire [4-1:0] node54358;
	wire [4-1:0] node54360;
	wire [4-1:0] node54363;
	wire [4-1:0] node54364;
	wire [4-1:0] node54367;
	wire [4-1:0] node54370;
	wire [4-1:0] node54371;
	wire [4-1:0] node54372;
	wire [4-1:0] node54373;
	wire [4-1:0] node54374;
	wire [4-1:0] node54379;
	wire [4-1:0] node54380;
	wire [4-1:0] node54381;
	wire [4-1:0] node54385;
	wire [4-1:0] node54386;
	wire [4-1:0] node54390;
	wire [4-1:0] node54391;
	wire [4-1:0] node54392;
	wire [4-1:0] node54393;
	wire [4-1:0] node54395;
	wire [4-1:0] node54398;
	wire [4-1:0] node54400;
	wire [4-1:0] node54403;
	wire [4-1:0] node54404;
	wire [4-1:0] node54408;
	wire [4-1:0] node54409;
	wire [4-1:0] node54412;
	wire [4-1:0] node54415;
	wire [4-1:0] node54416;
	wire [4-1:0] node54417;
	wire [4-1:0] node54418;
	wire [4-1:0] node54419;
	wire [4-1:0] node54420;
	wire [4-1:0] node54421;
	wire [4-1:0] node54422;
	wire [4-1:0] node54426;
	wire [4-1:0] node54427;
	wire [4-1:0] node54431;
	wire [4-1:0] node54432;
	wire [4-1:0] node54433;
	wire [4-1:0] node54437;
	wire [4-1:0] node54438;
	wire [4-1:0] node54442;
	wire [4-1:0] node54443;
	wire [4-1:0] node54444;
	wire [4-1:0] node54445;
	wire [4-1:0] node54448;
	wire [4-1:0] node54449;
	wire [4-1:0] node54453;
	wire [4-1:0] node54456;
	wire [4-1:0] node54457;
	wire [4-1:0] node54458;
	wire [4-1:0] node54459;
	wire [4-1:0] node54464;
	wire [4-1:0] node54465;
	wire [4-1:0] node54466;
	wire [4-1:0] node54470;
	wire [4-1:0] node54471;
	wire [4-1:0] node54475;
	wire [4-1:0] node54476;
	wire [4-1:0] node54477;
	wire [4-1:0] node54478;
	wire [4-1:0] node54479;
	wire [4-1:0] node54482;
	wire [4-1:0] node54486;
	wire [4-1:0] node54487;
	wire [4-1:0] node54490;
	wire [4-1:0] node54493;
	wire [4-1:0] node54494;
	wire [4-1:0] node54495;
	wire [4-1:0] node54498;
	wire [4-1:0] node54501;
	wire [4-1:0] node54502;
	wire [4-1:0] node54505;
	wire [4-1:0] node54508;
	wire [4-1:0] node54509;
	wire [4-1:0] node54510;
	wire [4-1:0] node54511;
	wire [4-1:0] node54512;
	wire [4-1:0] node54513;
	wire [4-1:0] node54514;
	wire [4-1:0] node54517;
	wire [4-1:0] node54520;
	wire [4-1:0] node54522;
	wire [4-1:0] node54525;
	wire [4-1:0] node54527;
	wire [4-1:0] node54529;
	wire [4-1:0] node54532;
	wire [4-1:0] node54533;
	wire [4-1:0] node54534;
	wire [4-1:0] node54537;
	wire [4-1:0] node54540;
	wire [4-1:0] node54542;
	wire [4-1:0] node54543;
	wire [4-1:0] node54546;
	wire [4-1:0] node54549;
	wire [4-1:0] node54550;
	wire [4-1:0] node54551;
	wire [4-1:0] node54553;
	wire [4-1:0] node54554;
	wire [4-1:0] node54559;
	wire [4-1:0] node54560;
	wire [4-1:0] node54563;
	wire [4-1:0] node54566;
	wire [4-1:0] node54567;
	wire [4-1:0] node54568;
	wire [4-1:0] node54569;
	wire [4-1:0] node54573;
	wire [4-1:0] node54574;
	wire [4-1:0] node54578;
	wire [4-1:0] node54579;
	wire [4-1:0] node54580;
	wire [4-1:0] node54584;
	wire [4-1:0] node54585;
	wire [4-1:0] node54589;
	wire [4-1:0] node54590;
	wire [4-1:0] node54591;
	wire [4-1:0] node54592;
	wire [4-1:0] node54593;
	wire [4-1:0] node54594;
	wire [4-1:0] node54595;
	wire [4-1:0] node54597;
	wire [4-1:0] node54600;
	wire [4-1:0] node54601;
	wire [4-1:0] node54604;
	wire [4-1:0] node54607;
	wire [4-1:0] node54609;
	wire [4-1:0] node54612;
	wire [4-1:0] node54613;
	wire [4-1:0] node54614;
	wire [4-1:0] node54615;
	wire [4-1:0] node54620;
	wire [4-1:0] node54621;
	wire [4-1:0] node54624;
	wire [4-1:0] node54627;
	wire [4-1:0] node54628;
	wire [4-1:0] node54629;
	wire [4-1:0] node54630;
	wire [4-1:0] node54632;
	wire [4-1:0] node54635;
	wire [4-1:0] node54638;
	wire [4-1:0] node54639;
	wire [4-1:0] node54642;
	wire [4-1:0] node54645;
	wire [4-1:0] node54646;
	wire [4-1:0] node54647;
	wire [4-1:0] node54650;
	wire [4-1:0] node54651;
	wire [4-1:0] node54656;
	wire [4-1:0] node54657;
	wire [4-1:0] node54658;
	wire [4-1:0] node54660;
	wire [4-1:0] node54661;
	wire [4-1:0] node54662;
	wire [4-1:0] node54665;
	wire [4-1:0] node54668;
	wire [4-1:0] node54670;
	wire [4-1:0] node54673;
	wire [4-1:0] node54674;
	wire [4-1:0] node54675;
	wire [4-1:0] node54678;
	wire [4-1:0] node54681;
	wire [4-1:0] node54682;
	wire [4-1:0] node54685;
	wire [4-1:0] node54688;
	wire [4-1:0] node54689;
	wire [4-1:0] node54692;
	wire [4-1:0] node54695;
	wire [4-1:0] node54696;
	wire [4-1:0] node54697;
	wire [4-1:0] node54698;
	wire [4-1:0] node54699;
	wire [4-1:0] node54701;
	wire [4-1:0] node54702;
	wire [4-1:0] node54705;
	wire [4-1:0] node54708;
	wire [4-1:0] node54709;
	wire [4-1:0] node54713;
	wire [4-1:0] node54714;
	wire [4-1:0] node54715;
	wire [4-1:0] node54716;
	wire [4-1:0] node54719;
	wire [4-1:0] node54722;
	wire [4-1:0] node54724;
	wire [4-1:0] node54727;
	wire [4-1:0] node54728;
	wire [4-1:0] node54731;
	wire [4-1:0] node54734;
	wire [4-1:0] node54735;
	wire [4-1:0] node54736;
	wire [4-1:0] node54738;
	wire [4-1:0] node54739;
	wire [4-1:0] node54743;
	wire [4-1:0] node54744;
	wire [4-1:0] node54747;
	wire [4-1:0] node54750;
	wire [4-1:0] node54751;
	wire [4-1:0] node54752;
	wire [4-1:0] node54753;
	wire [4-1:0] node54756;
	wire [4-1:0] node54761;
	wire [4-1:0] node54762;
	wire [4-1:0] node54763;
	wire [4-1:0] node54764;
	wire [4-1:0] node54768;
	wire [4-1:0] node54769;
	wire [4-1:0] node54773;
	wire [4-1:0] node54774;
	wire [4-1:0] node54775;
	wire [4-1:0] node54779;
	wire [4-1:0] node54780;
	wire [4-1:0] node54784;
	wire [4-1:0] node54785;
	wire [4-1:0] node54786;
	wire [4-1:0] node54787;
	wire [4-1:0] node54788;
	wire [4-1:0] node54789;
	wire [4-1:0] node54790;
	wire [4-1:0] node54791;
	wire [4-1:0] node54792;
	wire [4-1:0] node54793;
	wire [4-1:0] node54794;
	wire [4-1:0] node54798;
	wire [4-1:0] node54799;
	wire [4-1:0] node54803;
	wire [4-1:0] node54804;
	wire [4-1:0] node54805;
	wire [4-1:0] node54809;
	wire [4-1:0] node54810;
	wire [4-1:0] node54814;
	wire [4-1:0] node54815;
	wire [4-1:0] node54816;
	wire [4-1:0] node54817;
	wire [4-1:0] node54818;
	wire [4-1:0] node54821;
	wire [4-1:0] node54824;
	wire [4-1:0] node54825;
	wire [4-1:0] node54827;
	wire [4-1:0] node54831;
	wire [4-1:0] node54832;
	wire [4-1:0] node54835;
	wire [4-1:0] node54838;
	wire [4-1:0] node54839;
	wire [4-1:0] node54840;
	wire [4-1:0] node54841;
	wire [4-1:0] node54842;
	wire [4-1:0] node54847;
	wire [4-1:0] node54848;
	wire [4-1:0] node54850;
	wire [4-1:0] node54854;
	wire [4-1:0] node54855;
	wire [4-1:0] node54856;
	wire [4-1:0] node54857;
	wire [4-1:0] node54860;
	wire [4-1:0] node54863;
	wire [4-1:0] node54865;
	wire [4-1:0] node54869;
	wire [4-1:0] node54870;
	wire [4-1:0] node54871;
	wire [4-1:0] node54872;
	wire [4-1:0] node54873;
	wire [4-1:0] node54877;
	wire [4-1:0] node54878;
	wire [4-1:0] node54882;
	wire [4-1:0] node54883;
	wire [4-1:0] node54884;
	wire [4-1:0] node54888;
	wire [4-1:0] node54889;
	wire [4-1:0] node54893;
	wire [4-1:0] node54894;
	wire [4-1:0] node54895;
	wire [4-1:0] node54896;
	wire [4-1:0] node54897;
	wire [4-1:0] node54901;
	wire [4-1:0] node54902;
	wire [4-1:0] node54905;
	wire [4-1:0] node54908;
	wire [4-1:0] node54909;
	wire [4-1:0] node54910;
	wire [4-1:0] node54913;
	wire [4-1:0] node54916;
	wire [4-1:0] node54917;
	wire [4-1:0] node54920;
	wire [4-1:0] node54923;
	wire [4-1:0] node54924;
	wire [4-1:0] node54926;
	wire [4-1:0] node54927;
	wire [4-1:0] node54928;
	wire [4-1:0] node54931;
	wire [4-1:0] node54935;
	wire [4-1:0] node54936;
	wire [4-1:0] node54937;
	wire [4-1:0] node54938;
	wire [4-1:0] node54941;
	wire [4-1:0] node54944;
	wire [4-1:0] node54945;
	wire [4-1:0] node54949;
	wire [4-1:0] node54950;
	wire [4-1:0] node54954;
	wire [4-1:0] node54955;
	wire [4-1:0] node54956;
	wire [4-1:0] node54957;
	wire [4-1:0] node54958;
	wire [4-1:0] node54959;
	wire [4-1:0] node54960;
	wire [4-1:0] node54963;
	wire [4-1:0] node54966;
	wire [4-1:0] node54968;
	wire [4-1:0] node54969;
	wire [4-1:0] node54972;
	wire [4-1:0] node54975;
	wire [4-1:0] node54977;
	wire [4-1:0] node54980;
	wire [4-1:0] node54981;
	wire [4-1:0] node54984;
	wire [4-1:0] node54987;
	wire [4-1:0] node54988;
	wire [4-1:0] node54989;
	wire [4-1:0] node54990;
	wire [4-1:0] node54991;
	wire [4-1:0] node54994;
	wire [4-1:0] node54998;
	wire [4-1:0] node54999;
	wire [4-1:0] node55001;
	wire [4-1:0] node55002;
	wire [4-1:0] node55005;
	wire [4-1:0] node55008;
	wire [4-1:0] node55009;
	wire [4-1:0] node55012;
	wire [4-1:0] node55015;
	wire [4-1:0] node55016;
	wire [4-1:0] node55017;
	wire [4-1:0] node55018;
	wire [4-1:0] node55022;
	wire [4-1:0] node55023;
	wire [4-1:0] node55024;
	wire [4-1:0] node55027;
	wire [4-1:0] node55030;
	wire [4-1:0] node55032;
	wire [4-1:0] node55035;
	wire [4-1:0] node55036;
	wire [4-1:0] node55037;
	wire [4-1:0] node55038;
	wire [4-1:0] node55043;
	wire [4-1:0] node55044;
	wire [4-1:0] node55047;
	wire [4-1:0] node55050;
	wire [4-1:0] node55051;
	wire [4-1:0] node55052;
	wire [4-1:0] node55053;
	wire [4-1:0] node55054;
	wire [4-1:0] node55058;
	wire [4-1:0] node55059;
	wire [4-1:0] node55063;
	wire [4-1:0] node55064;
	wire [4-1:0] node55065;
	wire [4-1:0] node55069;
	wire [4-1:0] node55070;
	wire [4-1:0] node55074;
	wire [4-1:0] node55075;
	wire [4-1:0] node55076;
	wire [4-1:0] node55077;
	wire [4-1:0] node55078;
	wire [4-1:0] node55082;
	wire [4-1:0] node55083;
	wire [4-1:0] node55087;
	wire [4-1:0] node55088;
	wire [4-1:0] node55089;
	wire [4-1:0] node55093;
	wire [4-1:0] node55096;
	wire [4-1:0] node55097;
	wire [4-1:0] node55099;
	wire [4-1:0] node55100;
	wire [4-1:0] node55103;
	wire [4-1:0] node55106;
	wire [4-1:0] node55107;
	wire [4-1:0] node55108;
	wire [4-1:0] node55109;
	wire [4-1:0] node55112;
	wire [4-1:0] node55116;
	wire [4-1:0] node55118;
	wire [4-1:0] node55121;
	wire [4-1:0] node55122;
	wire [4-1:0] node55123;
	wire [4-1:0] node55124;
	wire [4-1:0] node55125;
	wire [4-1:0] node55126;
	wire [4-1:0] node55127;
	wire [4-1:0] node55128;
	wire [4-1:0] node55132;
	wire [4-1:0] node55133;
	wire [4-1:0] node55137;
	wire [4-1:0] node55138;
	wire [4-1:0] node55139;
	wire [4-1:0] node55144;
	wire [4-1:0] node55145;
	wire [4-1:0] node55146;
	wire [4-1:0] node55147;
	wire [4-1:0] node55151;
	wire [4-1:0] node55152;
	wire [4-1:0] node55153;
	wire [4-1:0] node55157;
	wire [4-1:0] node55160;
	wire [4-1:0] node55161;
	wire [4-1:0] node55164;
	wire [4-1:0] node55167;
	wire [4-1:0] node55168;
	wire [4-1:0] node55169;
	wire [4-1:0] node55170;
	wire [4-1:0] node55172;
	wire [4-1:0] node55175;
	wire [4-1:0] node55176;
	wire [4-1:0] node55180;
	wire [4-1:0] node55181;
	wire [4-1:0] node55182;
	wire [4-1:0] node55185;
	wire [4-1:0] node55188;
	wire [4-1:0] node55189;
	wire [4-1:0] node55192;
	wire [4-1:0] node55195;
	wire [4-1:0] node55196;
	wire [4-1:0] node55197;
	wire [4-1:0] node55198;
	wire [4-1:0] node55199;
	wire [4-1:0] node55203;
	wire [4-1:0] node55205;
	wire [4-1:0] node55208;
	wire [4-1:0] node55209;
	wire [4-1:0] node55212;
	wire [4-1:0] node55215;
	wire [4-1:0] node55216;
	wire [4-1:0] node55219;
	wire [4-1:0] node55222;
	wire [4-1:0] node55223;
	wire [4-1:0] node55224;
	wire [4-1:0] node55225;
	wire [4-1:0] node55226;
	wire [4-1:0] node55227;
	wire [4-1:0] node55230;
	wire [4-1:0] node55233;
	wire [4-1:0] node55235;
	wire [4-1:0] node55238;
	wire [4-1:0] node55239;
	wire [4-1:0] node55240;
	wire [4-1:0] node55244;
	wire [4-1:0] node55246;
	wire [4-1:0] node55249;
	wire [4-1:0] node55250;
	wire [4-1:0] node55251;
	wire [4-1:0] node55252;
	wire [4-1:0] node55256;
	wire [4-1:0] node55257;
	wire [4-1:0] node55259;
	wire [4-1:0] node55262;
	wire [4-1:0] node55265;
	wire [4-1:0] node55266;
	wire [4-1:0] node55267;
	wire [4-1:0] node55270;
	wire [4-1:0] node55271;
	wire [4-1:0] node55275;
	wire [4-1:0] node55277;
	wire [4-1:0] node55280;
	wire [4-1:0] node55281;
	wire [4-1:0] node55282;
	wire [4-1:0] node55283;
	wire [4-1:0] node55287;
	wire [4-1:0] node55288;
	wire [4-1:0] node55292;
	wire [4-1:0] node55293;
	wire [4-1:0] node55294;
	wire [4-1:0] node55298;
	wire [4-1:0] node55299;
	wire [4-1:0] node55303;
	wire [4-1:0] node55304;
	wire [4-1:0] node55305;
	wire [4-1:0] node55306;
	wire [4-1:0] node55307;
	wire [4-1:0] node55308;
	wire [4-1:0] node55309;
	wire [4-1:0] node55310;
	wire [4-1:0] node55313;
	wire [4-1:0] node55317;
	wire [4-1:0] node55319;
	wire [4-1:0] node55320;
	wire [4-1:0] node55323;
	wire [4-1:0] node55326;
	wire [4-1:0] node55327;
	wire [4-1:0] node55330;
	wire [4-1:0] node55333;
	wire [4-1:0] node55334;
	wire [4-1:0] node55335;
	wire [4-1:0] node55336;
	wire [4-1:0] node55337;
	wire [4-1:0] node55340;
	wire [4-1:0] node55344;
	wire [4-1:0] node55345;
	wire [4-1:0] node55346;
	wire [4-1:0] node55349;
	wire [4-1:0] node55352;
	wire [4-1:0] node55353;
	wire [4-1:0] node55357;
	wire [4-1:0] node55358;
	wire [4-1:0] node55361;
	wire [4-1:0] node55364;
	wire [4-1:0] node55365;
	wire [4-1:0] node55366;
	wire [4-1:0] node55367;
	wire [4-1:0] node55371;
	wire [4-1:0] node55372;
	wire [4-1:0] node55376;
	wire [4-1:0] node55377;
	wire [4-1:0] node55378;
	wire [4-1:0] node55382;
	wire [4-1:0] node55383;
	wire [4-1:0] node55387;
	wire [4-1:0] node55388;
	wire [4-1:0] node55389;
	wire [4-1:0] node55390;
	wire [4-1:0] node55391;
	wire [4-1:0] node55392;
	wire [4-1:0] node55393;
	wire [4-1:0] node55397;
	wire [4-1:0] node55399;
	wire [4-1:0] node55402;
	wire [4-1:0] node55403;
	wire [4-1:0] node55407;
	wire [4-1:0] node55408;
	wire [4-1:0] node55409;
	wire [4-1:0] node55410;
	wire [4-1:0] node55413;
	wire [4-1:0] node55417;
	wire [4-1:0] node55418;
	wire [4-1:0] node55419;
	wire [4-1:0] node55423;
	wire [4-1:0] node55426;
	wire [4-1:0] node55427;
	wire [4-1:0] node55428;
	wire [4-1:0] node55429;
	wire [4-1:0] node55432;
	wire [4-1:0] node55435;
	wire [4-1:0] node55436;
	wire [4-1:0] node55439;
	wire [4-1:0] node55442;
	wire [4-1:0] node55444;
	wire [4-1:0] node55445;
	wire [4-1:0] node55446;
	wire [4-1:0] node55449;
	wire [4-1:0] node55453;
	wire [4-1:0] node55454;
	wire [4-1:0] node55455;
	wire [4-1:0] node55456;
	wire [4-1:0] node55457;
	wire [4-1:0] node55460;
	wire [4-1:0] node55464;
	wire [4-1:0] node55465;
	wire [4-1:0] node55466;
	wire [4-1:0] node55468;
	wire [4-1:0] node55471;
	wire [4-1:0] node55473;
	wire [4-1:0] node55476;
	wire [4-1:0] node55477;
	wire [4-1:0] node55480;
	wire [4-1:0] node55483;
	wire [4-1:0] node55484;
	wire [4-1:0] node55485;
	wire [4-1:0] node55486;
	wire [4-1:0] node55490;
	wire [4-1:0] node55491;
	wire [4-1:0] node55495;
	wire [4-1:0] node55496;
	wire [4-1:0] node55497;
	wire [4-1:0] node55500;
	wire [4-1:0] node55503;
	wire [4-1:0] node55504;
	wire [4-1:0] node55506;
	wire [4-1:0] node55509;
	wire [4-1:0] node55510;
	wire [4-1:0] node55514;
	wire [4-1:0] node55515;
	wire [4-1:0] node55516;
	wire [4-1:0] node55517;
	wire [4-1:0] node55518;
	wire [4-1:0] node55519;
	wire [4-1:0] node55520;
	wire [4-1:0] node55521;
	wire [4-1:0] node55522;
	wire [4-1:0] node55524;
	wire [4-1:0] node55528;
	wire [4-1:0] node55530;
	wire [4-1:0] node55531;
	wire [4-1:0] node55535;
	wire [4-1:0] node55536;
	wire [4-1:0] node55538;
	wire [4-1:0] node55540;
	wire [4-1:0] node55543;
	wire [4-1:0] node55544;
	wire [4-1:0] node55546;
	wire [4-1:0] node55549;
	wire [4-1:0] node55552;
	wire [4-1:0] node55553;
	wire [4-1:0] node55554;
	wire [4-1:0] node55555;
	wire [4-1:0] node55557;
	wire [4-1:0] node55561;
	wire [4-1:0] node55563;
	wire [4-1:0] node55565;
	wire [4-1:0] node55568;
	wire [4-1:0] node55569;
	wire [4-1:0] node55570;
	wire [4-1:0] node55574;
	wire [4-1:0] node55575;
	wire [4-1:0] node55576;
	wire [4-1:0] node55580;
	wire [4-1:0] node55581;
	wire [4-1:0] node55584;
	wire [4-1:0] node55587;
	wire [4-1:0] node55588;
	wire [4-1:0] node55589;
	wire [4-1:0] node55590;
	wire [4-1:0] node55592;
	wire [4-1:0] node55595;
	wire [4-1:0] node55596;
	wire [4-1:0] node55597;
	wire [4-1:0] node55600;
	wire [4-1:0] node55603;
	wire [4-1:0] node55604;
	wire [4-1:0] node55608;
	wire [4-1:0] node55609;
	wire [4-1:0] node55610;
	wire [4-1:0] node55613;
	wire [4-1:0] node55616;
	wire [4-1:0] node55619;
	wire [4-1:0] node55620;
	wire [4-1:0] node55622;
	wire [4-1:0] node55623;
	wire [4-1:0] node55624;
	wire [4-1:0] node55628;
	wire [4-1:0] node55629;
	wire [4-1:0] node55633;
	wire [4-1:0] node55634;
	wire [4-1:0] node55635;
	wire [4-1:0] node55638;
	wire [4-1:0] node55641;
	wire [4-1:0] node55643;
	wire [4-1:0] node55644;
	wire [4-1:0] node55647;
	wire [4-1:0] node55650;
	wire [4-1:0] node55651;
	wire [4-1:0] node55652;
	wire [4-1:0] node55653;
	wire [4-1:0] node55654;
	wire [4-1:0] node55655;
	wire [4-1:0] node55658;
	wire [4-1:0] node55660;
	wire [4-1:0] node55663;
	wire [4-1:0] node55664;
	wire [4-1:0] node55665;
	wire [4-1:0] node55668;
	wire [4-1:0] node55672;
	wire [4-1:0] node55673;
	wire [4-1:0] node55675;
	wire [4-1:0] node55676;
	wire [4-1:0] node55679;
	wire [4-1:0] node55682;
	wire [4-1:0] node55683;
	wire [4-1:0] node55684;
	wire [4-1:0] node55687;
	wire [4-1:0] node55690;
	wire [4-1:0] node55691;
	wire [4-1:0] node55694;
	wire [4-1:0] node55697;
	wire [4-1:0] node55698;
	wire [4-1:0] node55699;
	wire [4-1:0] node55701;
	wire [4-1:0] node55704;
	wire [4-1:0] node55705;
	wire [4-1:0] node55708;
	wire [4-1:0] node55711;
	wire [4-1:0] node55712;
	wire [4-1:0] node55713;
	wire [4-1:0] node55716;
	wire [4-1:0] node55719;
	wire [4-1:0] node55720;
	wire [4-1:0] node55724;
	wire [4-1:0] node55725;
	wire [4-1:0] node55726;
	wire [4-1:0] node55727;
	wire [4-1:0] node55728;
	wire [4-1:0] node55729;
	wire [4-1:0] node55733;
	wire [4-1:0] node55736;
	wire [4-1:0] node55737;
	wire [4-1:0] node55740;
	wire [4-1:0] node55743;
	wire [4-1:0] node55744;
	wire [4-1:0] node55745;
	wire [4-1:0] node55746;
	wire [4-1:0] node55749;
	wire [4-1:0] node55752;
	wire [4-1:0] node55753;
	wire [4-1:0] node55757;
	wire [4-1:0] node55758;
	wire [4-1:0] node55759;
	wire [4-1:0] node55762;
	wire [4-1:0] node55765;
	wire [4-1:0] node55766;
	wire [4-1:0] node55769;
	wire [4-1:0] node55772;
	wire [4-1:0] node55773;
	wire [4-1:0] node55774;
	wire [4-1:0] node55775;
	wire [4-1:0] node55780;
	wire [4-1:0] node55781;
	wire [4-1:0] node55782;
	wire [4-1:0] node55784;
	wire [4-1:0] node55787;
	wire [4-1:0] node55790;
	wire [4-1:0] node55791;
	wire [4-1:0] node55792;
	wire [4-1:0] node55796;
	wire [4-1:0] node55798;
	wire [4-1:0] node55801;
	wire [4-1:0] node55802;
	wire [4-1:0] node55803;
	wire [4-1:0] node55804;
	wire [4-1:0] node55805;
	wire [4-1:0] node55806;
	wire [4-1:0] node55807;
	wire [4-1:0] node55810;
	wire [4-1:0] node55811;
	wire [4-1:0] node55815;
	wire [4-1:0] node55816;
	wire [4-1:0] node55819;
	wire [4-1:0] node55822;
	wire [4-1:0] node55823;
	wire [4-1:0] node55825;
	wire [4-1:0] node55828;
	wire [4-1:0] node55829;
	wire [4-1:0] node55832;
	wire [4-1:0] node55835;
	wire [4-1:0] node55836;
	wire [4-1:0] node55837;
	wire [4-1:0] node55838;
	wire [4-1:0] node55842;
	wire [4-1:0] node55843;
	wire [4-1:0] node55846;
	wire [4-1:0] node55849;
	wire [4-1:0] node55850;
	wire [4-1:0] node55851;
	wire [4-1:0] node55854;
	wire [4-1:0] node55857;
	wire [4-1:0] node55858;
	wire [4-1:0] node55860;
	wire [4-1:0] node55864;
	wire [4-1:0] node55865;
	wire [4-1:0] node55866;
	wire [4-1:0] node55867;
	wire [4-1:0] node55870;
	wire [4-1:0] node55871;
	wire [4-1:0] node55875;
	wire [4-1:0] node55876;
	wire [4-1:0] node55878;
	wire [4-1:0] node55881;
	wire [4-1:0] node55882;
	wire [4-1:0] node55885;
	wire [4-1:0] node55888;
	wire [4-1:0] node55889;
	wire [4-1:0] node55890;
	wire [4-1:0] node55892;
	wire [4-1:0] node55895;
	wire [4-1:0] node55896;
	wire [4-1:0] node55898;
	wire [4-1:0] node55901;
	wire [4-1:0] node55902;
	wire [4-1:0] node55905;
	wire [4-1:0] node55908;
	wire [4-1:0] node55909;
	wire [4-1:0] node55910;
	wire [4-1:0] node55913;
	wire [4-1:0] node55916;
	wire [4-1:0] node55918;
	wire [4-1:0] node55921;
	wire [4-1:0] node55922;
	wire [4-1:0] node55923;
	wire [4-1:0] node55924;
	wire [4-1:0] node55925;
	wire [4-1:0] node55928;
	wire [4-1:0] node55931;
	wire [4-1:0] node55932;
	wire [4-1:0] node55935;
	wire [4-1:0] node55938;
	wire [4-1:0] node55939;
	wire [4-1:0] node55940;
	wire [4-1:0] node55943;
	wire [4-1:0] node55946;
	wire [4-1:0] node55947;
	wire [4-1:0] node55951;
	wire [4-1:0] node55952;
	wire [4-1:0] node55953;
	wire [4-1:0] node55954;
	wire [4-1:0] node55957;
	wire [4-1:0] node55960;
	wire [4-1:0] node55961;
	wire [4-1:0] node55964;
	wire [4-1:0] node55967;
	wire [4-1:0] node55968;
	wire [4-1:0] node55969;
	wire [4-1:0] node55970;
	wire [4-1:0] node55971;
	wire [4-1:0] node55974;
	wire [4-1:0] node55977;
	wire [4-1:0] node55978;
	wire [4-1:0] node55981;
	wire [4-1:0] node55984;
	wire [4-1:0] node55985;
	wire [4-1:0] node55988;
	wire [4-1:0] node55991;
	wire [4-1:0] node55992;
	wire [4-1:0] node55995;
	wire [4-1:0] node55998;
	wire [4-1:0] node55999;
	wire [4-1:0] node56000;
	wire [4-1:0] node56001;
	wire [4-1:0] node56002;
	wire [4-1:0] node56003;
	wire [4-1:0] node56004;
	wire [4-1:0] node56005;
	wire [4-1:0] node56007;
	wire [4-1:0] node56010;
	wire [4-1:0] node56011;
	wire [4-1:0] node56015;
	wire [4-1:0] node56018;
	wire [4-1:0] node56019;
	wire [4-1:0] node56020;
	wire [4-1:0] node56021;
	wire [4-1:0] node56025;
	wire [4-1:0] node56026;
	wire [4-1:0] node56030;
	wire [4-1:0] node56031;
	wire [4-1:0] node56032;
	wire [4-1:0] node56035;
	wire [4-1:0] node56038;
	wire [4-1:0] node56039;
	wire [4-1:0] node56042;
	wire [4-1:0] node56045;
	wire [4-1:0] node56046;
	wire [4-1:0] node56047;
	wire [4-1:0] node56049;
	wire [4-1:0] node56050;
	wire [4-1:0] node56054;
	wire [4-1:0] node56055;
	wire [4-1:0] node56058;
	wire [4-1:0] node56059;
	wire [4-1:0] node56063;
	wire [4-1:0] node56064;
	wire [4-1:0] node56065;
	wire [4-1:0] node56069;
	wire [4-1:0] node56070;
	wire [4-1:0] node56071;
	wire [4-1:0] node56075;
	wire [4-1:0] node56077;
	wire [4-1:0] node56080;
	wire [4-1:0] node56081;
	wire [4-1:0] node56082;
	wire [4-1:0] node56083;
	wire [4-1:0] node56085;
	wire [4-1:0] node56088;
	wire [4-1:0] node56089;
	wire [4-1:0] node56093;
	wire [4-1:0] node56094;
	wire [4-1:0] node56095;
	wire [4-1:0] node56098;
	wire [4-1:0] node56101;
	wire [4-1:0] node56102;
	wire [4-1:0] node56105;
	wire [4-1:0] node56108;
	wire [4-1:0] node56109;
	wire [4-1:0] node56110;
	wire [4-1:0] node56111;
	wire [4-1:0] node56114;
	wire [4-1:0] node56117;
	wire [4-1:0] node56120;
	wire [4-1:0] node56121;
	wire [4-1:0] node56123;
	wire [4-1:0] node56124;
	wire [4-1:0] node56127;
	wire [4-1:0] node56130;
	wire [4-1:0] node56133;
	wire [4-1:0] node56134;
	wire [4-1:0] node56135;
	wire [4-1:0] node56136;
	wire [4-1:0] node56137;
	wire [4-1:0] node56139;
	wire [4-1:0] node56140;
	wire [4-1:0] node56143;
	wire [4-1:0] node56146;
	wire [4-1:0] node56147;
	wire [4-1:0] node56148;
	wire [4-1:0] node56152;
	wire [4-1:0] node56154;
	wire [4-1:0] node56157;
	wire [4-1:0] node56158;
	wire [4-1:0] node56159;
	wire [4-1:0] node56160;
	wire [4-1:0] node56163;
	wire [4-1:0] node56167;
	wire [4-1:0] node56168;
	wire [4-1:0] node56169;
	wire [4-1:0] node56172;
	wire [4-1:0] node56175;
	wire [4-1:0] node56176;
	wire [4-1:0] node56180;
	wire [4-1:0] node56181;
	wire [4-1:0] node56182;
	wire [4-1:0] node56183;
	wire [4-1:0] node56185;
	wire [4-1:0] node56189;
	wire [4-1:0] node56190;
	wire [4-1:0] node56191;
	wire [4-1:0] node56195;
	wire [4-1:0] node56198;
	wire [4-1:0] node56199;
	wire [4-1:0] node56200;
	wire [4-1:0] node56202;
	wire [4-1:0] node56205;
	wire [4-1:0] node56207;
	wire [4-1:0] node56210;
	wire [4-1:0] node56211;
	wire [4-1:0] node56212;
	wire [4-1:0] node56215;
	wire [4-1:0] node56218;
	wire [4-1:0] node56219;
	wire [4-1:0] node56222;
	wire [4-1:0] node56225;
	wire [4-1:0] node56226;
	wire [4-1:0] node56227;
	wire [4-1:0] node56228;
	wire [4-1:0] node56231;
	wire [4-1:0] node56232;
	wire [4-1:0] node56234;
	wire [4-1:0] node56237;
	wire [4-1:0] node56238;
	wire [4-1:0] node56241;
	wire [4-1:0] node56244;
	wire [4-1:0] node56245;
	wire [4-1:0] node56246;
	wire [4-1:0] node56247;
	wire [4-1:0] node56250;
	wire [4-1:0] node56253;
	wire [4-1:0] node56255;
	wire [4-1:0] node56259;
	wire [4-1:0] node56260;
	wire [4-1:0] node56261;
	wire [4-1:0] node56262;
	wire [4-1:0] node56265;
	wire [4-1:0] node56268;
	wire [4-1:0] node56269;
	wire [4-1:0] node56270;
	wire [4-1:0] node56273;
	wire [4-1:0] node56276;
	wire [4-1:0] node56277;
	wire [4-1:0] node56281;
	wire [4-1:0] node56282;
	wire [4-1:0] node56284;
	wire [4-1:0] node56285;
	wire [4-1:0] node56288;
	wire [4-1:0] node56291;
	wire [4-1:0] node56292;
	wire [4-1:0] node56295;
	wire [4-1:0] node56298;
	wire [4-1:0] node56299;
	wire [4-1:0] node56300;
	wire [4-1:0] node56301;
	wire [4-1:0] node56302;
	wire [4-1:0] node56303;
	wire [4-1:0] node56307;
	wire [4-1:0] node56308;
	wire [4-1:0] node56312;
	wire [4-1:0] node56313;
	wire [4-1:0] node56314;
	wire [4-1:0] node56318;
	wire [4-1:0] node56319;
	wire [4-1:0] node56323;
	wire [4-1:0] node56324;
	wire [4-1:0] node56325;
	wire [4-1:0] node56326;
	wire [4-1:0] node56327;
	wire [4-1:0] node56330;
	wire [4-1:0] node56333;
	wire [4-1:0] node56335;
	wire [4-1:0] node56338;
	wire [4-1:0] node56339;
	wire [4-1:0] node56340;
	wire [4-1:0] node56343;
	wire [4-1:0] node56346;
	wire [4-1:0] node56347;
	wire [4-1:0] node56348;
	wire [4-1:0] node56351;
	wire [4-1:0] node56354;
	wire [4-1:0] node56355;
	wire [4-1:0] node56358;
	wire [4-1:0] node56361;
	wire [4-1:0] node56362;
	wire [4-1:0] node56363;
	wire [4-1:0] node56364;
	wire [4-1:0] node56367;
	wire [4-1:0] node56370;
	wire [4-1:0] node56371;
	wire [4-1:0] node56374;
	wire [4-1:0] node56377;
	wire [4-1:0] node56378;
	wire [4-1:0] node56381;
	wire [4-1:0] node56384;
	wire [4-1:0] node56385;
	wire [4-1:0] node56386;
	wire [4-1:0] node56387;
	wire [4-1:0] node56388;
	wire [4-1:0] node56389;
	wire [4-1:0] node56393;
	wire [4-1:0] node56394;
	wire [4-1:0] node56398;
	wire [4-1:0] node56399;
	wire [4-1:0] node56400;
	wire [4-1:0] node56401;
	wire [4-1:0] node56406;
	wire [4-1:0] node56409;
	wire [4-1:0] node56410;
	wire [4-1:0] node56411;
	wire [4-1:0] node56413;
	wire [4-1:0] node56416;
	wire [4-1:0] node56419;
	wire [4-1:0] node56420;
	wire [4-1:0] node56424;
	wire [4-1:0] node56425;
	wire [4-1:0] node56426;
	wire [4-1:0] node56427;
	wire [4-1:0] node56431;
	wire [4-1:0] node56432;
	wire [4-1:0] node56436;
	wire [4-1:0] node56437;
	wire [4-1:0] node56438;
	wire [4-1:0] node56442;
	wire [4-1:0] node56443;
	wire [4-1:0] node56447;
	wire [4-1:0] node56448;
	wire [4-1:0] node56449;
	wire [4-1:0] node56450;
	wire [4-1:0] node56451;
	wire [4-1:0] node56452;
	wire [4-1:0] node56453;
	wire [4-1:0] node56454;
	wire [4-1:0] node56455;
	wire [4-1:0] node56457;
	wire [4-1:0] node56460;
	wire [4-1:0] node56462;
	wire [4-1:0] node56465;
	wire [4-1:0] node56466;
	wire [4-1:0] node56468;
	wire [4-1:0] node56471;
	wire [4-1:0] node56474;
	wire [4-1:0] node56475;
	wire [4-1:0] node56476;
	wire [4-1:0] node56477;
	wire [4-1:0] node56478;
	wire [4-1:0] node56482;
	wire [4-1:0] node56485;
	wire [4-1:0] node56486;
	wire [4-1:0] node56489;
	wire [4-1:0] node56491;
	wire [4-1:0] node56494;
	wire [4-1:0] node56495;
	wire [4-1:0] node56498;
	wire [4-1:0] node56501;
	wire [4-1:0] node56502;
	wire [4-1:0] node56503;
	wire [4-1:0] node56505;
	wire [4-1:0] node56507;
	wire [4-1:0] node56510;
	wire [4-1:0] node56512;
	wire [4-1:0] node56513;
	wire [4-1:0] node56516;
	wire [4-1:0] node56519;
	wire [4-1:0] node56520;
	wire [4-1:0] node56521;
	wire [4-1:0] node56522;
	wire [4-1:0] node56526;
	wire [4-1:0] node56529;
	wire [4-1:0] node56531;
	wire [4-1:0] node56532;
	wire [4-1:0] node56533;
	wire [4-1:0] node56538;
	wire [4-1:0] node56539;
	wire [4-1:0] node56540;
	wire [4-1:0] node56541;
	wire [4-1:0] node56542;
	wire [4-1:0] node56543;
	wire [4-1:0] node56546;
	wire [4-1:0] node56549;
	wire [4-1:0] node56550;
	wire [4-1:0] node56554;
	wire [4-1:0] node56555;
	wire [4-1:0] node56558;
	wire [4-1:0] node56561;
	wire [4-1:0] node56562;
	wire [4-1:0] node56563;
	wire [4-1:0] node56565;
	wire [4-1:0] node56568;
	wire [4-1:0] node56570;
	wire [4-1:0] node56572;
	wire [4-1:0] node56575;
	wire [4-1:0] node56576;
	wire [4-1:0] node56578;
	wire [4-1:0] node56581;
	wire [4-1:0] node56582;
	wire [4-1:0] node56586;
	wire [4-1:0] node56587;
	wire [4-1:0] node56588;
	wire [4-1:0] node56589;
	wire [4-1:0] node56591;
	wire [4-1:0] node56592;
	wire [4-1:0] node56596;
	wire [4-1:0] node56597;
	wire [4-1:0] node56600;
	wire [4-1:0] node56603;
	wire [4-1:0] node56605;
	wire [4-1:0] node56606;
	wire [4-1:0] node56607;
	wire [4-1:0] node56610;
	wire [4-1:0] node56614;
	wire [4-1:0] node56615;
	wire [4-1:0] node56616;
	wire [4-1:0] node56617;
	wire [4-1:0] node56621;
	wire [4-1:0] node56622;
	wire [4-1:0] node56625;
	wire [4-1:0] node56628;
	wire [4-1:0] node56629;
	wire [4-1:0] node56632;
	wire [4-1:0] node56635;
	wire [4-1:0] node56636;
	wire [4-1:0] node56637;
	wire [4-1:0] node56638;
	wire [4-1:0] node56639;
	wire [4-1:0] node56640;
	wire [4-1:0] node56641;
	wire [4-1:0] node56644;
	wire [4-1:0] node56647;
	wire [4-1:0] node56648;
	wire [4-1:0] node56651;
	wire [4-1:0] node56654;
	wire [4-1:0] node56655;
	wire [4-1:0] node56656;
	wire [4-1:0] node56660;
	wire [4-1:0] node56663;
	wire [4-1:0] node56664;
	wire [4-1:0] node56665;
	wire [4-1:0] node56666;
	wire [4-1:0] node56669;
	wire [4-1:0] node56672;
	wire [4-1:0] node56674;
	wire [4-1:0] node56677;
	wire [4-1:0] node56678;
	wire [4-1:0] node56679;
	wire [4-1:0] node56682;
	wire [4-1:0] node56685;
	wire [4-1:0] node56686;
	wire [4-1:0] node56689;
	wire [4-1:0] node56692;
	wire [4-1:0] node56693;
	wire [4-1:0] node56694;
	wire [4-1:0] node56695;
	wire [4-1:0] node56698;
	wire [4-1:0] node56699;
	wire [4-1:0] node56703;
	wire [4-1:0] node56704;
	wire [4-1:0] node56706;
	wire [4-1:0] node56709;
	wire [4-1:0] node56710;
	wire [4-1:0] node56713;
	wire [4-1:0] node56716;
	wire [4-1:0] node56717;
	wire [4-1:0] node56718;
	wire [4-1:0] node56719;
	wire [4-1:0] node56723;
	wire [4-1:0] node56726;
	wire [4-1:0] node56727;
	wire [4-1:0] node56728;
	wire [4-1:0] node56731;
	wire [4-1:0] node56734;
	wire [4-1:0] node56735;
	wire [4-1:0] node56739;
	wire [4-1:0] node56740;
	wire [4-1:0] node56741;
	wire [4-1:0] node56742;
	wire [4-1:0] node56744;
	wire [4-1:0] node56747;
	wire [4-1:0] node56748;
	wire [4-1:0] node56749;
	wire [4-1:0] node56752;
	wire [4-1:0] node56755;
	wire [4-1:0] node56756;
	wire [4-1:0] node56760;
	wire [4-1:0] node56761;
	wire [4-1:0] node56762;
	wire [4-1:0] node56763;
	wire [4-1:0] node56764;
	wire [4-1:0] node56767;
	wire [4-1:0] node56772;
	wire [4-1:0] node56773;
	wire [4-1:0] node56774;
	wire [4-1:0] node56775;
	wire [4-1:0] node56778;
	wire [4-1:0] node56782;
	wire [4-1:0] node56784;
	wire [4-1:0] node56785;
	wire [4-1:0] node56788;
	wire [4-1:0] node56791;
	wire [4-1:0] node56792;
	wire [4-1:0] node56793;
	wire [4-1:0] node56794;
	wire [4-1:0] node56797;
	wire [4-1:0] node56800;
	wire [4-1:0] node56801;
	wire [4-1:0] node56803;
	wire [4-1:0] node56804;
	wire [4-1:0] node56808;
	wire [4-1:0] node56810;
	wire [4-1:0] node56811;
	wire [4-1:0] node56815;
	wire [4-1:0] node56816;
	wire [4-1:0] node56817;
	wire [4-1:0] node56820;
	wire [4-1:0] node56823;
	wire [4-1:0] node56824;
	wire [4-1:0] node56828;
	wire [4-1:0] node56829;
	wire [4-1:0] node56830;
	wire [4-1:0] node56831;
	wire [4-1:0] node56832;
	wire [4-1:0] node56833;
	wire [4-1:0] node56834;
	wire [4-1:0] node56835;
	wire [4-1:0] node56836;
	wire [4-1:0] node56839;
	wire [4-1:0] node56842;
	wire [4-1:0] node56843;
	wire [4-1:0] node56846;
	wire [4-1:0] node56849;
	wire [4-1:0] node56850;
	wire [4-1:0] node56853;
	wire [4-1:0] node56856;
	wire [4-1:0] node56858;
	wire [4-1:0] node56860;
	wire [4-1:0] node56863;
	wire [4-1:0] node56864;
	wire [4-1:0] node56865;
	wire [4-1:0] node56866;
	wire [4-1:0] node56869;
	wire [4-1:0] node56872;
	wire [4-1:0] node56873;
	wire [4-1:0] node56876;
	wire [4-1:0] node56879;
	wire [4-1:0] node56880;
	wire [4-1:0] node56881;
	wire [4-1:0] node56884;
	wire [4-1:0] node56887;
	wire [4-1:0] node56888;
	wire [4-1:0] node56892;
	wire [4-1:0] node56893;
	wire [4-1:0] node56894;
	wire [4-1:0] node56895;
	wire [4-1:0] node56897;
	wire [4-1:0] node56900;
	wire [4-1:0] node56901;
	wire [4-1:0] node56905;
	wire [4-1:0] node56907;
	wire [4-1:0] node56908;
	wire [4-1:0] node56909;
	wire [4-1:0] node56914;
	wire [4-1:0] node56915;
	wire [4-1:0] node56916;
	wire [4-1:0] node56917;
	wire [4-1:0] node56920;
	wire [4-1:0] node56923;
	wire [4-1:0] node56925;
	wire [4-1:0] node56927;
	wire [4-1:0] node56930;
	wire [4-1:0] node56931;
	wire [4-1:0] node56932;
	wire [4-1:0] node56935;
	wire [4-1:0] node56938;
	wire [4-1:0] node56939;
	wire [4-1:0] node56943;
	wire [4-1:0] node56944;
	wire [4-1:0] node56945;
	wire [4-1:0] node56946;
	wire [4-1:0] node56947;
	wire [4-1:0] node56950;
	wire [4-1:0] node56953;
	wire [4-1:0] node56954;
	wire [4-1:0] node56956;
	wire [4-1:0] node56957;
	wire [4-1:0] node56960;
	wire [4-1:0] node56963;
	wire [4-1:0] node56964;
	wire [4-1:0] node56967;
	wire [4-1:0] node56970;
	wire [4-1:0] node56971;
	wire [4-1:0] node56972;
	wire [4-1:0] node56973;
	wire [4-1:0] node56975;
	wire [4-1:0] node56980;
	wire [4-1:0] node56981;
	wire [4-1:0] node56983;
	wire [4-1:0] node56984;
	wire [4-1:0] node56988;
	wire [4-1:0] node56989;
	wire [4-1:0] node56990;
	wire [4-1:0] node56993;
	wire [4-1:0] node56996;
	wire [4-1:0] node56998;
	wire [4-1:0] node57001;
	wire [4-1:0] node57002;
	wire [4-1:0] node57003;
	wire [4-1:0] node57004;
	wire [4-1:0] node57005;
	wire [4-1:0] node57008;
	wire [4-1:0] node57011;
	wire [4-1:0] node57013;
	wire [4-1:0] node57016;
	wire [4-1:0] node57017;
	wire [4-1:0] node57020;
	wire [4-1:0] node57023;
	wire [4-1:0] node57024;
	wire [4-1:0] node57025;
	wire [4-1:0] node57027;
	wire [4-1:0] node57030;
	wire [4-1:0] node57033;
	wire [4-1:0] node57034;
	wire [4-1:0] node57035;
	wire [4-1:0] node57038;
	wire [4-1:0] node57041;
	wire [4-1:0] node57042;
	wire [4-1:0] node57043;
	wire [4-1:0] node57046;
	wire [4-1:0] node57049;
	wire [4-1:0] node57050;
	wire [4-1:0] node57053;
	wire [4-1:0] node57056;
	wire [4-1:0] node57057;
	wire [4-1:0] node57058;
	wire [4-1:0] node57059;
	wire [4-1:0] node57060;
	wire [4-1:0] node57061;
	wire [4-1:0] node57062;
	wire [4-1:0] node57066;
	wire [4-1:0] node57067;
	wire [4-1:0] node57069;
	wire [4-1:0] node57073;
	wire [4-1:0] node57074;
	wire [4-1:0] node57077;
	wire [4-1:0] node57079;
	wire [4-1:0] node57080;
	wire [4-1:0] node57083;
	wire [4-1:0] node57086;
	wire [4-1:0] node57087;
	wire [4-1:0] node57088;
	wire [4-1:0] node57089;
	wire [4-1:0] node57090;
	wire [4-1:0] node57093;
	wire [4-1:0] node57097;
	wire [4-1:0] node57098;
	wire [4-1:0] node57101;
	wire [4-1:0] node57104;
	wire [4-1:0] node57105;
	wire [4-1:0] node57106;
	wire [4-1:0] node57109;
	wire [4-1:0] node57112;
	wire [4-1:0] node57115;
	wire [4-1:0] node57116;
	wire [4-1:0] node57117;
	wire [4-1:0] node57118;
	wire [4-1:0] node57119;
	wire [4-1:0] node57122;
	wire [4-1:0] node57125;
	wire [4-1:0] node57126;
	wire [4-1:0] node57127;
	wire [4-1:0] node57130;
	wire [4-1:0] node57133;
	wire [4-1:0] node57134;
	wire [4-1:0] node57138;
	wire [4-1:0] node57139;
	wire [4-1:0] node57140;
	wire [4-1:0] node57141;
	wire [4-1:0] node57145;
	wire [4-1:0] node57146;
	wire [4-1:0] node57151;
	wire [4-1:0] node57152;
	wire [4-1:0] node57153;
	wire [4-1:0] node57157;
	wire [4-1:0] node57158;
	wire [4-1:0] node57159;
	wire [4-1:0] node57164;
	wire [4-1:0] node57165;
	wire [4-1:0] node57166;
	wire [4-1:0] node57167;
	wire [4-1:0] node57168;
	wire [4-1:0] node57170;
	wire [4-1:0] node57174;
	wire [4-1:0] node57175;
	wire [4-1:0] node57176;
	wire [4-1:0] node57180;
	wire [4-1:0] node57183;
	wire [4-1:0] node57184;
	wire [4-1:0] node57185;
	wire [4-1:0] node57186;
	wire [4-1:0] node57187;
	wire [4-1:0] node57190;
	wire [4-1:0] node57194;
	wire [4-1:0] node57195;
	wire [4-1:0] node57198;
	wire [4-1:0] node57201;
	wire [4-1:0] node57202;
	wire [4-1:0] node57203;
	wire [4-1:0] node57207;
	wire [4-1:0] node57210;
	wire [4-1:0] node57211;
	wire [4-1:0] node57212;
	wire [4-1:0] node57213;
	wire [4-1:0] node57215;
	wire [4-1:0] node57217;
	wire [4-1:0] node57220;
	wire [4-1:0] node57221;
	wire [4-1:0] node57224;
	wire [4-1:0] node57227;
	wire [4-1:0] node57228;
	wire [4-1:0] node57229;
	wire [4-1:0] node57233;
	wire [4-1:0] node57236;
	wire [4-1:0] node57237;
	wire [4-1:0] node57238;
	wire [4-1:0] node57240;
	wire [4-1:0] node57243;
	wire [4-1:0] node57246;
	wire [4-1:0] node57249;
	wire [4-1:0] node57250;
	wire [4-1:0] node57251;
	wire [4-1:0] node57252;
	wire [4-1:0] node57253;
	wire [4-1:0] node57254;
	wire [4-1:0] node57255;
	wire [4-1:0] node57257;
	wire [4-1:0] node57258;
	wire [4-1:0] node57261;
	wire [4-1:0] node57264;
	wire [4-1:0] node57265;
	wire [4-1:0] node57266;
	wire [4-1:0] node57268;
	wire [4-1:0] node57272;
	wire [4-1:0] node57273;
	wire [4-1:0] node57276;
	wire [4-1:0] node57279;
	wire [4-1:0] node57280;
	wire [4-1:0] node57281;
	wire [4-1:0] node57282;
	wire [4-1:0] node57285;
	wire [4-1:0] node57288;
	wire [4-1:0] node57289;
	wire [4-1:0] node57291;
	wire [4-1:0] node57294;
	wire [4-1:0] node57295;
	wire [4-1:0] node57298;
	wire [4-1:0] node57301;
	wire [4-1:0] node57302;
	wire [4-1:0] node57303;
	wire [4-1:0] node57307;
	wire [4-1:0] node57308;
	wire [4-1:0] node57312;
	wire [4-1:0] node57313;
	wire [4-1:0] node57314;
	wire [4-1:0] node57315;
	wire [4-1:0] node57317;
	wire [4-1:0] node57320;
	wire [4-1:0] node57321;
	wire [4-1:0] node57324;
	wire [4-1:0] node57327;
	wire [4-1:0] node57328;
	wire [4-1:0] node57331;
	wire [4-1:0] node57334;
	wire [4-1:0] node57335;
	wire [4-1:0] node57336;
	wire [4-1:0] node57337;
	wire [4-1:0] node57340;
	wire [4-1:0] node57343;
	wire [4-1:0] node57345;
	wire [4-1:0] node57346;
	wire [4-1:0] node57349;
	wire [4-1:0] node57352;
	wire [4-1:0] node57353;
	wire [4-1:0] node57354;
	wire [4-1:0] node57356;
	wire [4-1:0] node57359;
	wire [4-1:0] node57361;
	wire [4-1:0] node57365;
	wire [4-1:0] node57366;
	wire [4-1:0] node57367;
	wire [4-1:0] node57368;
	wire [4-1:0] node57369;
	wire [4-1:0] node57371;
	wire [4-1:0] node57374;
	wire [4-1:0] node57375;
	wire [4-1:0] node57379;
	wire [4-1:0] node57380;
	wire [4-1:0] node57381;
	wire [4-1:0] node57384;
	wire [4-1:0] node57387;
	wire [4-1:0] node57389;
	wire [4-1:0] node57392;
	wire [4-1:0] node57393;
	wire [4-1:0] node57394;
	wire [4-1:0] node57396;
	wire [4-1:0] node57399;
	wire [4-1:0] node57400;
	wire [4-1:0] node57404;
	wire [4-1:0] node57405;
	wire [4-1:0] node57406;
	wire [4-1:0] node57409;
	wire [4-1:0] node57412;
	wire [4-1:0] node57413;
	wire [4-1:0] node57416;
	wire [4-1:0] node57419;
	wire [4-1:0] node57420;
	wire [4-1:0] node57421;
	wire [4-1:0] node57423;
	wire [4-1:0] node57424;
	wire [4-1:0] node57427;
	wire [4-1:0] node57429;
	wire [4-1:0] node57432;
	wire [4-1:0] node57433;
	wire [4-1:0] node57434;
	wire [4-1:0] node57438;
	wire [4-1:0] node57441;
	wire [4-1:0] node57442;
	wire [4-1:0] node57443;
	wire [4-1:0] node57444;
	wire [4-1:0] node57447;
	wire [4-1:0] node57450;
	wire [4-1:0] node57451;
	wire [4-1:0] node57453;
	wire [4-1:0] node57456;
	wire [4-1:0] node57458;
	wire [4-1:0] node57461;
	wire [4-1:0] node57462;
	wire [4-1:0] node57465;
	wire [4-1:0] node57468;
	wire [4-1:0] node57469;
	wire [4-1:0] node57470;
	wire [4-1:0] node57471;
	wire [4-1:0] node57472;
	wire [4-1:0] node57473;
	wire [4-1:0] node57474;
	wire [4-1:0] node57475;
	wire [4-1:0] node57478;
	wire [4-1:0] node57481;
	wire [4-1:0] node57482;
	wire [4-1:0] node57485;
	wire [4-1:0] node57488;
	wire [4-1:0] node57489;
	wire [4-1:0] node57493;
	wire [4-1:0] node57494;
	wire [4-1:0] node57497;
	wire [4-1:0] node57500;
	wire [4-1:0] node57501;
	wire [4-1:0] node57503;
	wire [4-1:0] node57504;
	wire [4-1:0] node57507;
	wire [4-1:0] node57510;
	wire [4-1:0] node57511;
	wire [4-1:0] node57512;
	wire [4-1:0] node57516;
	wire [4-1:0] node57517;
	wire [4-1:0] node57518;
	wire [4-1:0] node57522;
	wire [4-1:0] node57523;
	wire [4-1:0] node57526;
	wire [4-1:0] node57529;
	wire [4-1:0] node57530;
	wire [4-1:0] node57531;
	wire [4-1:0] node57532;
	wire [4-1:0] node57535;
	wire [4-1:0] node57538;
	wire [4-1:0] node57539;
	wire [4-1:0] node57542;
	wire [4-1:0] node57545;
	wire [4-1:0] node57546;
	wire [4-1:0] node57547;
	wire [4-1:0] node57551;
	wire [4-1:0] node57554;
	wire [4-1:0] node57555;
	wire [4-1:0] node57556;
	wire [4-1:0] node57557;
	wire [4-1:0] node57558;
	wire [4-1:0] node57561;
	wire [4-1:0] node57564;
	wire [4-1:0] node57565;
	wire [4-1:0] node57568;
	wire [4-1:0] node57571;
	wire [4-1:0] node57572;
	wire [4-1:0] node57573;
	wire [4-1:0] node57576;
	wire [4-1:0] node57579;
	wire [4-1:0] node57580;
	wire [4-1:0] node57581;
	wire [4-1:0] node57584;
	wire [4-1:0] node57587;
	wire [4-1:0] node57588;
	wire [4-1:0] node57591;
	wire [4-1:0] node57594;
	wire [4-1:0] node57595;
	wire [4-1:0] node57596;
	wire [4-1:0] node57597;
	wire [4-1:0] node57598;
	wire [4-1:0] node57601;
	wire [4-1:0] node57605;
	wire [4-1:0] node57606;
	wire [4-1:0] node57609;
	wire [4-1:0] node57612;
	wire [4-1:0] node57613;
	wire [4-1:0] node57614;
	wire [4-1:0] node57617;
	wire [4-1:0] node57620;
	wire [4-1:0] node57621;
	wire [4-1:0] node57624;
	wire [4-1:0] node57627;
	wire [4-1:0] node57628;
	wire [4-1:0] node57629;
	wire [4-1:0] node57630;
	wire [4-1:0] node57631;
	wire [4-1:0] node57632;
	wire [4-1:0] node57633;
	wire [4-1:0] node57635;
	wire [4-1:0] node57637;
	wire [4-1:0] node57640;
	wire [4-1:0] node57642;
	wire [4-1:0] node57645;
	wire [4-1:0] node57646;
	wire [4-1:0] node57647;
	wire [4-1:0] node57651;
	wire [4-1:0] node57654;
	wire [4-1:0] node57655;
	wire [4-1:0] node57656;
	wire [4-1:0] node57657;
	wire [4-1:0] node57658;
	wire [4-1:0] node57661;
	wire [4-1:0] node57664;
	wire [4-1:0] node57666;
	wire [4-1:0] node57669;
	wire [4-1:0] node57670;
	wire [4-1:0] node57673;
	wire [4-1:0] node57676;
	wire [4-1:0] node57677;
	wire [4-1:0] node57678;
	wire [4-1:0] node57682;
	wire [4-1:0] node57685;
	wire [4-1:0] node57686;
	wire [4-1:0] node57687;
	wire [4-1:0] node57688;
	wire [4-1:0] node57690;
	wire [4-1:0] node57693;
	wire [4-1:0] node57694;
	wire [4-1:0] node57698;
	wire [4-1:0] node57700;
	wire [4-1:0] node57703;
	wire [4-1:0] node57704;
	wire [4-1:0] node57705;
	wire [4-1:0] node57708;
	wire [4-1:0] node57710;
	wire [4-1:0] node57713;
	wire [4-1:0] node57714;
	wire [4-1:0] node57717;
	wire [4-1:0] node57720;
	wire [4-1:0] node57721;
	wire [4-1:0] node57722;
	wire [4-1:0] node57723;
	wire [4-1:0] node57724;
	wire [4-1:0] node57725;
	wire [4-1:0] node57729;
	wire [4-1:0] node57730;
	wire [4-1:0] node57732;
	wire [4-1:0] node57735;
	wire [4-1:0] node57736;
	wire [4-1:0] node57739;
	wire [4-1:0] node57742;
	wire [4-1:0] node57743;
	wire [4-1:0] node57744;
	wire [4-1:0] node57745;
	wire [4-1:0] node57748;
	wire [4-1:0] node57751;
	wire [4-1:0] node57754;
	wire [4-1:0] node57755;
	wire [4-1:0] node57758;
	wire [4-1:0] node57761;
	wire [4-1:0] node57762;
	wire [4-1:0] node57763;
	wire [4-1:0] node57764;
	wire [4-1:0] node57765;
	wire [4-1:0] node57768;
	wire [4-1:0] node57772;
	wire [4-1:0] node57774;
	wire [4-1:0] node57777;
	wire [4-1:0] node57778;
	wire [4-1:0] node57779;
	wire [4-1:0] node57780;
	wire [4-1:0] node57783;
	wire [4-1:0] node57787;
	wire [4-1:0] node57788;
	wire [4-1:0] node57789;
	wire [4-1:0] node57794;
	wire [4-1:0] node57795;
	wire [4-1:0] node57796;
	wire [4-1:0] node57797;
	wire [4-1:0] node57799;
	wire [4-1:0] node57802;
	wire [4-1:0] node57803;
	wire [4-1:0] node57806;
	wire [4-1:0] node57809;
	wire [4-1:0] node57810;
	wire [4-1:0] node57811;
	wire [4-1:0] node57815;
	wire [4-1:0] node57818;
	wire [4-1:0] node57819;
	wire [4-1:0] node57821;
	wire [4-1:0] node57822;
	wire [4-1:0] node57823;
	wire [4-1:0] node57827;
	wire [4-1:0] node57828;
	wire [4-1:0] node57831;
	wire [4-1:0] node57834;
	wire [4-1:0] node57835;
	wire [4-1:0] node57836;
	wire [4-1:0] node57840;
	wire [4-1:0] node57843;
	wire [4-1:0] node57844;
	wire [4-1:0] node57845;
	wire [4-1:0] node57846;
	wire [4-1:0] node57847;
	wire [4-1:0] node57848;
	wire [4-1:0] node57850;
	wire [4-1:0] node57853;
	wire [4-1:0] node57856;
	wire [4-1:0] node57857;
	wire [4-1:0] node57860;
	wire [4-1:0] node57862;
	wire [4-1:0] node57865;
	wire [4-1:0] node57866;
	wire [4-1:0] node57867;
	wire [4-1:0] node57868;
	wire [4-1:0] node57870;
	wire [4-1:0] node57873;
	wire [4-1:0] node57875;
	wire [4-1:0] node57878;
	wire [4-1:0] node57879;
	wire [4-1:0] node57881;
	wire [4-1:0] node57884;
	wire [4-1:0] node57886;
	wire [4-1:0] node57889;
	wire [4-1:0] node57890;
	wire [4-1:0] node57892;
	wire [4-1:0] node57895;
	wire [4-1:0] node57896;
	wire [4-1:0] node57897;
	wire [4-1:0] node57900;
	wire [4-1:0] node57903;
	wire [4-1:0] node57905;
	wire [4-1:0] node57908;
	wire [4-1:0] node57909;
	wire [4-1:0] node57910;
	wire [4-1:0] node57911;
	wire [4-1:0] node57913;
	wire [4-1:0] node57914;
	wire [4-1:0] node57918;
	wire [4-1:0] node57919;
	wire [4-1:0] node57921;
	wire [4-1:0] node57924;
	wire [4-1:0] node57926;
	wire [4-1:0] node57929;
	wire [4-1:0] node57930;
	wire [4-1:0] node57931;
	wire [4-1:0] node57934;
	wire [4-1:0] node57937;
	wire [4-1:0] node57938;
	wire [4-1:0] node57941;
	wire [4-1:0] node57944;
	wire [4-1:0] node57945;
	wire [4-1:0] node57946;
	wire [4-1:0] node57949;
	wire [4-1:0] node57952;
	wire [4-1:0] node57953;
	wire [4-1:0] node57956;
	wire [4-1:0] node57959;
	wire [4-1:0] node57960;
	wire [4-1:0] node57961;
	wire [4-1:0] node57962;
	wire [4-1:0] node57963;
	wire [4-1:0] node57965;
	wire [4-1:0] node57967;
	wire [4-1:0] node57970;
	wire [4-1:0] node57971;
	wire [4-1:0] node57974;
	wire [4-1:0] node57977;
	wire [4-1:0] node57978;
	wire [4-1:0] node57979;
	wire [4-1:0] node57981;
	wire [4-1:0] node57984;
	wire [4-1:0] node57987;
	wire [4-1:0] node57988;
	wire [4-1:0] node57989;
	wire [4-1:0] node57992;
	wire [4-1:0] node57995;
	wire [4-1:0] node57997;
	wire [4-1:0] node58000;
	wire [4-1:0] node58001;
	wire [4-1:0] node58002;
	wire [4-1:0] node58003;
	wire [4-1:0] node58007;
	wire [4-1:0] node58008;
	wire [4-1:0] node58012;
	wire [4-1:0] node58013;
	wire [4-1:0] node58014;
	wire [4-1:0] node58018;
	wire [4-1:0] node58019;
	wire [4-1:0] node58023;
	wire [4-1:0] node58024;
	wire [4-1:0] node58025;
	wire [4-1:0] node58028;
	wire [4-1:0] node58029;
	wire [4-1:0] node58033;
	wire [4-1:0] node58034;
	wire [4-1:0] node58035;
	wire [4-1:0] node58039;
	wire [4-1:0] node58040;
	wire [4-1:0] node58044;
	wire [4-1:0] node58045;
	wire [4-1:0] node58046;
	wire [4-1:0] node58047;
	wire [4-1:0] node58048;
	wire [4-1:0] node58049;
	wire [4-1:0] node58050;
	wire [4-1:0] node58051;
	wire [4-1:0] node58052;
	wire [4-1:0] node58053;
	wire [4-1:0] node58056;
	wire [4-1:0] node58059;
	wire [4-1:0] node58060;
	wire [4-1:0] node58061;
	wire [4-1:0] node58064;
	wire [4-1:0] node58067;
	wire [4-1:0] node58069;
	wire [4-1:0] node58072;
	wire [4-1:0] node58073;
	wire [4-1:0] node58074;
	wire [4-1:0] node58076;
	wire [4-1:0] node58079;
	wire [4-1:0] node58080;
	wire [4-1:0] node58083;
	wire [4-1:0] node58086;
	wire [4-1:0] node58087;
	wire [4-1:0] node58089;
	wire [4-1:0] node58092;
	wire [4-1:0] node58093;
	wire [4-1:0] node58097;
	wire [4-1:0] node58098;
	wire [4-1:0] node58099;
	wire [4-1:0] node58100;
	wire [4-1:0] node58101;
	wire [4-1:0] node58104;
	wire [4-1:0] node58108;
	wire [4-1:0] node58109;
	wire [4-1:0] node58111;
	wire [4-1:0] node58114;
	wire [4-1:0] node58115;
	wire [4-1:0] node58118;
	wire [4-1:0] node58121;
	wire [4-1:0] node58122;
	wire [4-1:0] node58123;
	wire [4-1:0] node58126;
	wire [4-1:0] node58129;
	wire [4-1:0] node58130;
	wire [4-1:0] node58133;
	wire [4-1:0] node58136;
	wire [4-1:0] node58137;
	wire [4-1:0] node58138;
	wire [4-1:0] node58139;
	wire [4-1:0] node58140;
	wire [4-1:0] node58141;
	wire [4-1:0] node58145;
	wire [4-1:0] node58146;
	wire [4-1:0] node58149;
	wire [4-1:0] node58152;
	wire [4-1:0] node58153;
	wire [4-1:0] node58154;
	wire [4-1:0] node58158;
	wire [4-1:0] node58160;
	wire [4-1:0] node58163;
	wire [4-1:0] node58164;
	wire [4-1:0] node58165;
	wire [4-1:0] node58168;
	wire [4-1:0] node58171;
	wire [4-1:0] node58172;
	wire [4-1:0] node58173;
	wire [4-1:0] node58177;
	wire [4-1:0] node58180;
	wire [4-1:0] node58181;
	wire [4-1:0] node58182;
	wire [4-1:0] node58183;
	wire [4-1:0] node58186;
	wire [4-1:0] node58187;
	wire [4-1:0] node58191;
	wire [4-1:0] node58193;
	wire [4-1:0] node58194;
	wire [4-1:0] node58198;
	wire [4-1:0] node58199;
	wire [4-1:0] node58200;
	wire [4-1:0] node58203;
	wire [4-1:0] node58204;
	wire [4-1:0] node58207;
	wire [4-1:0] node58210;
	wire [4-1:0] node58211;
	wire [4-1:0] node58212;
	wire [4-1:0] node58215;
	wire [4-1:0] node58218;
	wire [4-1:0] node58219;
	wire [4-1:0] node58222;
	wire [4-1:0] node58225;
	wire [4-1:0] node58226;
	wire [4-1:0] node58227;
	wire [4-1:0] node58228;
	wire [4-1:0] node58229;
	wire [4-1:0] node58231;
	wire [4-1:0] node58232;
	wire [4-1:0] node58233;
	wire [4-1:0] node58237;
	wire [4-1:0] node58238;
	wire [4-1:0] node58242;
	wire [4-1:0] node58243;
	wire [4-1:0] node58244;
	wire [4-1:0] node58245;
	wire [4-1:0] node58248;
	wire [4-1:0] node58252;
	wire [4-1:0] node58253;
	wire [4-1:0] node58254;
	wire [4-1:0] node58257;
	wire [4-1:0] node58261;
	wire [4-1:0] node58262;
	wire [4-1:0] node58263;
	wire [4-1:0] node58265;
	wire [4-1:0] node58268;
	wire [4-1:0] node58270;
	wire [4-1:0] node58271;
	wire [4-1:0] node58274;
	wire [4-1:0] node58277;
	wire [4-1:0] node58278;
	wire [4-1:0] node58279;
	wire [4-1:0] node58280;
	wire [4-1:0] node58283;
	wire [4-1:0] node58287;
	wire [4-1:0] node58290;
	wire [4-1:0] node58291;
	wire [4-1:0] node58292;
	wire [4-1:0] node58293;
	wire [4-1:0] node58294;
	wire [4-1:0] node58298;
	wire [4-1:0] node58299;
	wire [4-1:0] node58303;
	wire [4-1:0] node58304;
	wire [4-1:0] node58306;
	wire [4-1:0] node58309;
	wire [4-1:0] node58311;
	wire [4-1:0] node58314;
	wire [4-1:0] node58315;
	wire [4-1:0] node58316;
	wire [4-1:0] node58317;
	wire [4-1:0] node58320;
	wire [4-1:0] node58323;
	wire [4-1:0] node58324;
	wire [4-1:0] node58328;
	wire [4-1:0] node58329;
	wire [4-1:0] node58331;
	wire [4-1:0] node58334;
	wire [4-1:0] node58336;
	wire [4-1:0] node58339;
	wire [4-1:0] node58340;
	wire [4-1:0] node58341;
	wire [4-1:0] node58342;
	wire [4-1:0] node58343;
	wire [4-1:0] node58344;
	wire [4-1:0] node58345;
	wire [4-1:0] node58349;
	wire [4-1:0] node58351;
	wire [4-1:0] node58354;
	wire [4-1:0] node58355;
	wire [4-1:0] node58358;
	wire [4-1:0] node58361;
	wire [4-1:0] node58362;
	wire [4-1:0] node58363;
	wire [4-1:0] node58367;
	wire [4-1:0] node58368;
	wire [4-1:0] node58371;
	wire [4-1:0] node58374;
	wire [4-1:0] node58375;
	wire [4-1:0] node58376;
	wire [4-1:0] node58377;
	wire [4-1:0] node58380;
	wire [4-1:0] node58383;
	wire [4-1:0] node58384;
	wire [4-1:0] node58385;
	wire [4-1:0] node58389;
	wire [4-1:0] node58392;
	wire [4-1:0] node58393;
	wire [4-1:0] node58394;
	wire [4-1:0] node58395;
	wire [4-1:0] node58398;
	wire [4-1:0] node58401;
	wire [4-1:0] node58402;
	wire [4-1:0] node58405;
	wire [4-1:0] node58408;
	wire [4-1:0] node58411;
	wire [4-1:0] node58412;
	wire [4-1:0] node58413;
	wire [4-1:0] node58414;
	wire [4-1:0] node58416;
	wire [4-1:0] node58419;
	wire [4-1:0] node58421;
	wire [4-1:0] node58424;
	wire [4-1:0] node58425;
	wire [4-1:0] node58426;
	wire [4-1:0] node58429;
	wire [4-1:0] node58432;
	wire [4-1:0] node58433;
	wire [4-1:0] node58436;
	wire [4-1:0] node58439;
	wire [4-1:0] node58440;
	wire [4-1:0] node58441;
	wire [4-1:0] node58442;
	wire [4-1:0] node58446;
	wire [4-1:0] node58447;
	wire [4-1:0] node58450;
	wire [4-1:0] node58453;
	wire [4-1:0] node58454;
	wire [4-1:0] node58456;
	wire [4-1:0] node58459;
	wire [4-1:0] node58461;
	wire [4-1:0] node58463;
	wire [4-1:0] node58466;
	wire [4-1:0] node58467;
	wire [4-1:0] node58468;
	wire [4-1:0] node58469;
	wire [4-1:0] node58470;
	wire [4-1:0] node58471;
	wire [4-1:0] node58472;
	wire [4-1:0] node58473;
	wire [4-1:0] node58475;
	wire [4-1:0] node58478;
	wire [4-1:0] node58479;
	wire [4-1:0] node58483;
	wire [4-1:0] node58485;
	wire [4-1:0] node58488;
	wire [4-1:0] node58489;
	wire [4-1:0] node58490;
	wire [4-1:0] node58491;
	wire [4-1:0] node58494;
	wire [4-1:0] node58499;
	wire [4-1:0] node58500;
	wire [4-1:0] node58501;
	wire [4-1:0] node58502;
	wire [4-1:0] node58505;
	wire [4-1:0] node58508;
	wire [4-1:0] node58509;
	wire [4-1:0] node58512;
	wire [4-1:0] node58515;
	wire [4-1:0] node58516;
	wire [4-1:0] node58517;
	wire [4-1:0] node58521;
	wire [4-1:0] node58524;
	wire [4-1:0] node58525;
	wire [4-1:0] node58526;
	wire [4-1:0] node58527;
	wire [4-1:0] node58528;
	wire [4-1:0] node58531;
	wire [4-1:0] node58534;
	wire [4-1:0] node58535;
	wire [4-1:0] node58538;
	wire [4-1:0] node58541;
	wire [4-1:0] node58542;
	wire [4-1:0] node58543;
	wire [4-1:0] node58547;
	wire [4-1:0] node58550;
	wire [4-1:0] node58551;
	wire [4-1:0] node58552;
	wire [4-1:0] node58554;
	wire [4-1:0] node58557;
	wire [4-1:0] node58559;
	wire [4-1:0] node58562;
	wire [4-1:0] node58564;
	wire [4-1:0] node58567;
	wire [4-1:0] node58568;
	wire [4-1:0] node58569;
	wire [4-1:0] node58570;
	wire [4-1:0] node58571;
	wire [4-1:0] node58573;
	wire [4-1:0] node58575;
	wire [4-1:0] node58578;
	wire [4-1:0] node58579;
	wire [4-1:0] node58580;
	wire [4-1:0] node58583;
	wire [4-1:0] node58586;
	wire [4-1:0] node58589;
	wire [4-1:0] node58590;
	wire [4-1:0] node58592;
	wire [4-1:0] node58593;
	wire [4-1:0] node58597;
	wire [4-1:0] node58598;
	wire [4-1:0] node58599;
	wire [4-1:0] node58602;
	wire [4-1:0] node58606;
	wire [4-1:0] node58607;
	wire [4-1:0] node58608;
	wire [4-1:0] node58609;
	wire [4-1:0] node58611;
	wire [4-1:0] node58616;
	wire [4-1:0] node58617;
	wire [4-1:0] node58618;
	wire [4-1:0] node58619;
	wire [4-1:0] node58624;
	wire [4-1:0] node58625;
	wire [4-1:0] node58626;
	wire [4-1:0] node58629;
	wire [4-1:0] node58632;
	wire [4-1:0] node58634;
	wire [4-1:0] node58637;
	wire [4-1:0] node58638;
	wire [4-1:0] node58639;
	wire [4-1:0] node58640;
	wire [4-1:0] node58643;
	wire [4-1:0] node58644;
	wire [4-1:0] node58647;
	wire [4-1:0] node58650;
	wire [4-1:0] node58651;
	wire [4-1:0] node58652;
	wire [4-1:0] node58654;
	wire [4-1:0] node58658;
	wire [4-1:0] node58659;
	wire [4-1:0] node58661;
	wire [4-1:0] node58664;
	wire [4-1:0] node58665;
	wire [4-1:0] node58668;
	wire [4-1:0] node58671;
	wire [4-1:0] node58672;
	wire [4-1:0] node58673;
	wire [4-1:0] node58675;
	wire [4-1:0] node58678;
	wire [4-1:0] node58680;
	wire [4-1:0] node58681;
	wire [4-1:0] node58684;
	wire [4-1:0] node58687;
	wire [4-1:0] node58688;
	wire [4-1:0] node58689;
	wire [4-1:0] node58692;
	wire [4-1:0] node58695;
	wire [4-1:0] node58696;
	wire [4-1:0] node58699;
	wire [4-1:0] node58702;
	wire [4-1:0] node58703;
	wire [4-1:0] node58704;
	wire [4-1:0] node58705;
	wire [4-1:0] node58706;
	wire [4-1:0] node58707;
	wire [4-1:0] node58708;
	wire [4-1:0] node58711;
	wire [4-1:0] node58714;
	wire [4-1:0] node58715;
	wire [4-1:0] node58718;
	wire [4-1:0] node58721;
	wire [4-1:0] node58722;
	wire [4-1:0] node58725;
	wire [4-1:0] node58728;
	wire [4-1:0] node58729;
	wire [4-1:0] node58730;
	wire [4-1:0] node58734;
	wire [4-1:0] node58737;
	wire [4-1:0] node58738;
	wire [4-1:0] node58739;
	wire [4-1:0] node58740;
	wire [4-1:0] node58742;
	wire [4-1:0] node58745;
	wire [4-1:0] node58747;
	wire [4-1:0] node58749;
	wire [4-1:0] node58752;
	wire [4-1:0] node58753;
	wire [4-1:0] node58756;
	wire [4-1:0] node58759;
	wire [4-1:0] node58760;
	wire [4-1:0] node58761;
	wire [4-1:0] node58765;
	wire [4-1:0] node58768;
	wire [4-1:0] node58769;
	wire [4-1:0] node58770;
	wire [4-1:0] node58771;
	wire [4-1:0] node58772;
	wire [4-1:0] node58775;
	wire [4-1:0] node58778;
	wire [4-1:0] node58779;
	wire [4-1:0] node58782;
	wire [4-1:0] node58785;
	wire [4-1:0] node58786;
	wire [4-1:0] node58787;
	wire [4-1:0] node58791;
	wire [4-1:0] node58794;
	wire [4-1:0] node58795;
	wire [4-1:0] node58796;
	wire [4-1:0] node58798;
	wire [4-1:0] node58801;
	wire [4-1:0] node58804;
	wire [4-1:0] node58805;
	wire [4-1:0] node58806;
	wire [4-1:0] node58809;
	wire [4-1:0] node58812;
	wire [4-1:0] node58813;
	wire [4-1:0] node58814;
	wire [4-1:0] node58817;
	wire [4-1:0] node58820;
	wire [4-1:0] node58821;
	wire [4-1:0] node58824;
	wire [4-1:0] node58827;
	wire [4-1:0] node58828;
	wire [4-1:0] node58829;
	wire [4-1:0] node58830;
	wire [4-1:0] node58831;
	wire [4-1:0] node58832;
	wire [4-1:0] node58833;
	wire [4-1:0] node58834;
	wire [4-1:0] node58835;
	wire [4-1:0] node58836;
	wire [4-1:0] node58840;
	wire [4-1:0] node58842;
	wire [4-1:0] node58845;
	wire [4-1:0] node58846;
	wire [4-1:0] node58849;
	wire [4-1:0] node58852;
	wire [4-1:0] node58853;
	wire [4-1:0] node58854;
	wire [4-1:0] node58857;
	wire [4-1:0] node58860;
	wire [4-1:0] node58861;
	wire [4-1:0] node58864;
	wire [4-1:0] node58866;
	wire [4-1:0] node58869;
	wire [4-1:0] node58870;
	wire [4-1:0] node58871;
	wire [4-1:0] node58872;
	wire [4-1:0] node58875;
	wire [4-1:0] node58878;
	wire [4-1:0] node58879;
	wire [4-1:0] node58883;
	wire [4-1:0] node58884;
	wire [4-1:0] node58886;
	wire [4-1:0] node58889;
	wire [4-1:0] node58891;
	wire [4-1:0] node58894;
	wire [4-1:0] node58895;
	wire [4-1:0] node58896;
	wire [4-1:0] node58897;
	wire [4-1:0] node58898;
	wire [4-1:0] node58903;
	wire [4-1:0] node58904;
	wire [4-1:0] node58907;
	wire [4-1:0] node58910;
	wire [4-1:0] node58911;
	wire [4-1:0] node58912;
	wire [4-1:0] node58915;
	wire [4-1:0] node58918;
	wire [4-1:0] node58919;
	wire [4-1:0] node58922;
	wire [4-1:0] node58925;
	wire [4-1:0] node58926;
	wire [4-1:0] node58927;
	wire [4-1:0] node58928;
	wire [4-1:0] node58929;
	wire [4-1:0] node58932;
	wire [4-1:0] node58934;
	wire [4-1:0] node58937;
	wire [4-1:0] node58938;
	wire [4-1:0] node58939;
	wire [4-1:0] node58940;
	wire [4-1:0] node58943;
	wire [4-1:0] node58946;
	wire [4-1:0] node58947;
	wire [4-1:0] node58950;
	wire [4-1:0] node58954;
	wire [4-1:0] node58955;
	wire [4-1:0] node58956;
	wire [4-1:0] node58957;
	wire [4-1:0] node58961;
	wire [4-1:0] node58963;
	wire [4-1:0] node58966;
	wire [4-1:0] node58967;
	wire [4-1:0] node58968;
	wire [4-1:0] node58970;
	wire [4-1:0] node58973;
	wire [4-1:0] node58974;
	wire [4-1:0] node58977;
	wire [4-1:0] node58980;
	wire [4-1:0] node58981;
	wire [4-1:0] node58984;
	wire [4-1:0] node58987;
	wire [4-1:0] node58988;
	wire [4-1:0] node58989;
	wire [4-1:0] node58990;
	wire [4-1:0] node58991;
	wire [4-1:0] node58994;
	wire [4-1:0] node58997;
	wire [4-1:0] node58999;
	wire [4-1:0] node59000;
	wire [4-1:0] node59004;
	wire [4-1:0] node59005;
	wire [4-1:0] node59006;
	wire [4-1:0] node59007;
	wire [4-1:0] node59010;
	wire [4-1:0] node59013;
	wire [4-1:0] node59014;
	wire [4-1:0] node59017;
	wire [4-1:0] node59020;
	wire [4-1:0] node59021;
	wire [4-1:0] node59025;
	wire [4-1:0] node59026;
	wire [4-1:0] node59027;
	wire [4-1:0] node59028;
	wire [4-1:0] node59030;
	wire [4-1:0] node59033;
	wire [4-1:0] node59034;
	wire [4-1:0] node59038;
	wire [4-1:0] node59040;
	wire [4-1:0] node59042;
	wire [4-1:0] node59045;
	wire [4-1:0] node59046;
	wire [4-1:0] node59047;
	wire [4-1:0] node59048;
	wire [4-1:0] node59051;
	wire [4-1:0] node59054;
	wire [4-1:0] node59056;
	wire [4-1:0] node59059;
	wire [4-1:0] node59061;
	wire [4-1:0] node59062;
	wire [4-1:0] node59065;
	wire [4-1:0] node59068;
	wire [4-1:0] node59069;
	wire [4-1:0] node59070;
	wire [4-1:0] node59071;
	wire [4-1:0] node59072;
	wire [4-1:0] node59073;
	wire [4-1:0] node59076;
	wire [4-1:0] node59079;
	wire [4-1:0] node59080;
	wire [4-1:0] node59083;
	wire [4-1:0] node59086;
	wire [4-1:0] node59087;
	wire [4-1:0] node59088;
	wire [4-1:0] node59091;
	wire [4-1:0] node59094;
	wire [4-1:0] node59095;
	wire [4-1:0] node59098;
	wire [4-1:0] node59101;
	wire [4-1:0] node59102;
	wire [4-1:0] node59103;
	wire [4-1:0] node59104;
	wire [4-1:0] node59107;
	wire [4-1:0] node59110;
	wire [4-1:0] node59111;
	wire [4-1:0] node59114;
	wire [4-1:0] node59117;
	wire [4-1:0] node59118;
	wire [4-1:0] node59119;
	wire [4-1:0] node59123;
	wire [4-1:0] node59126;
	wire [4-1:0] node59127;
	wire [4-1:0] node59128;
	wire [4-1:0] node59129;
	wire [4-1:0] node59130;
	wire [4-1:0] node59131;
	wire [4-1:0] node59134;
	wire [4-1:0] node59137;
	wire [4-1:0] node59138;
	wire [4-1:0] node59139;
	wire [4-1:0] node59143;
	wire [4-1:0] node59146;
	wire [4-1:0] node59147;
	wire [4-1:0] node59150;
	wire [4-1:0] node59153;
	wire [4-1:0] node59154;
	wire [4-1:0] node59155;
	wire [4-1:0] node59158;
	wire [4-1:0] node59161;
	wire [4-1:0] node59162;
	wire [4-1:0] node59163;
	wire [4-1:0] node59167;
	wire [4-1:0] node59170;
	wire [4-1:0] node59171;
	wire [4-1:0] node59172;
	wire [4-1:0] node59173;
	wire [4-1:0] node59174;
	wire [4-1:0] node59175;
	wire [4-1:0] node59178;
	wire [4-1:0] node59181;
	wire [4-1:0] node59182;
	wire [4-1:0] node59185;
	wire [4-1:0] node59188;
	wire [4-1:0] node59190;
	wire [4-1:0] node59191;
	wire [4-1:0] node59195;
	wire [4-1:0] node59196;
	wire [4-1:0] node59199;
	wire [4-1:0] node59202;
	wire [4-1:0] node59203;
	wire [4-1:0] node59204;
	wire [4-1:0] node59208;
	wire [4-1:0] node59211;
	wire [4-1:0] node59212;
	wire [4-1:0] node59213;
	wire [4-1:0] node59214;
	wire [4-1:0] node59215;
	wire [4-1:0] node59216;
	wire [4-1:0] node59217;
	wire [4-1:0] node59220;
	wire [4-1:0] node59223;
	wire [4-1:0] node59224;
	wire [4-1:0] node59225;
	wire [4-1:0] node59228;
	wire [4-1:0] node59232;
	wire [4-1:0] node59233;
	wire [4-1:0] node59234;
	wire [4-1:0] node59236;
	wire [4-1:0] node59239;
	wire [4-1:0] node59240;
	wire [4-1:0] node59243;
	wire [4-1:0] node59246;
	wire [4-1:0] node59247;
	wire [4-1:0] node59248;
	wire [4-1:0] node59252;
	wire [4-1:0] node59253;
	wire [4-1:0] node59254;
	wire [4-1:0] node59257;
	wire [4-1:0] node59260;
	wire [4-1:0] node59261;
	wire [4-1:0] node59264;
	wire [4-1:0] node59267;
	wire [4-1:0] node59268;
	wire [4-1:0] node59269;
	wire [4-1:0] node59270;
	wire [4-1:0] node59271;
	wire [4-1:0] node59274;
	wire [4-1:0] node59277;
	wire [4-1:0] node59278;
	wire [4-1:0] node59279;
	wire [4-1:0] node59282;
	wire [4-1:0] node59285;
	wire [4-1:0] node59287;
	wire [4-1:0] node59290;
	wire [4-1:0] node59291;
	wire [4-1:0] node59292;
	wire [4-1:0] node59295;
	wire [4-1:0] node59298;
	wire [4-1:0] node59299;
	wire [4-1:0] node59302;
	wire [4-1:0] node59305;
	wire [4-1:0] node59306;
	wire [4-1:0] node59307;
	wire [4-1:0] node59308;
	wire [4-1:0] node59309;
	wire [4-1:0] node59312;
	wire [4-1:0] node59315;
	wire [4-1:0] node59316;
	wire [4-1:0] node59319;
	wire [4-1:0] node59322;
	wire [4-1:0] node59323;
	wire [4-1:0] node59327;
	wire [4-1:0] node59328;
	wire [4-1:0] node59331;
	wire [4-1:0] node59334;
	wire [4-1:0] node59335;
	wire [4-1:0] node59336;
	wire [4-1:0] node59337;
	wire [4-1:0] node59338;
	wire [4-1:0] node59341;
	wire [4-1:0] node59343;
	wire [4-1:0] node59344;
	wire [4-1:0] node59347;
	wire [4-1:0] node59350;
	wire [4-1:0] node59351;
	wire [4-1:0] node59352;
	wire [4-1:0] node59353;
	wire [4-1:0] node59356;
	wire [4-1:0] node59361;
	wire [4-1:0] node59362;
	wire [4-1:0] node59363;
	wire [4-1:0] node59365;
	wire [4-1:0] node59367;
	wire [4-1:0] node59370;
	wire [4-1:0] node59371;
	wire [4-1:0] node59372;
	wire [4-1:0] node59375;
	wire [4-1:0] node59378;
	wire [4-1:0] node59379;
	wire [4-1:0] node59382;
	wire [4-1:0] node59385;
	wire [4-1:0] node59386;
	wire [4-1:0] node59387;
	wire [4-1:0] node59390;
	wire [4-1:0] node59392;
	wire [4-1:0] node59395;
	wire [4-1:0] node59396;
	wire [4-1:0] node59397;
	wire [4-1:0] node59400;
	wire [4-1:0] node59403;
	wire [4-1:0] node59406;
	wire [4-1:0] node59407;
	wire [4-1:0] node59408;
	wire [4-1:0] node59409;
	wire [4-1:0] node59411;
	wire [4-1:0] node59412;
	wire [4-1:0] node59415;
	wire [4-1:0] node59418;
	wire [4-1:0] node59419;
	wire [4-1:0] node59423;
	wire [4-1:0] node59424;
	wire [4-1:0] node59426;
	wire [4-1:0] node59429;
	wire [4-1:0] node59430;
	wire [4-1:0] node59431;
	wire [4-1:0] node59434;
	wire [4-1:0] node59437;
	wire [4-1:0] node59438;
	wire [4-1:0] node59442;
	wire [4-1:0] node59443;
	wire [4-1:0] node59444;
	wire [4-1:0] node59445;
	wire [4-1:0] node59447;
	wire [4-1:0] node59451;
	wire [4-1:0] node59453;
	wire [4-1:0] node59456;
	wire [4-1:0] node59457;
	wire [4-1:0] node59458;
	wire [4-1:0] node59459;
	wire [4-1:0] node59464;
	wire [4-1:0] node59467;
	wire [4-1:0] node59468;
	wire [4-1:0] node59469;
	wire [4-1:0] node59470;
	wire [4-1:0] node59471;
	wire [4-1:0] node59472;
	wire [4-1:0] node59474;
	wire [4-1:0] node59477;
	wire [4-1:0] node59480;
	wire [4-1:0] node59481;
	wire [4-1:0] node59485;
	wire [4-1:0] node59486;
	wire [4-1:0] node59487;
	wire [4-1:0] node59488;
	wire [4-1:0] node59489;
	wire [4-1:0] node59492;
	wire [4-1:0] node59496;
	wire [4-1:0] node59498;
	wire [4-1:0] node59499;
	wire [4-1:0] node59502;
	wire [4-1:0] node59505;
	wire [4-1:0] node59506;
	wire [4-1:0] node59510;
	wire [4-1:0] node59511;
	wire [4-1:0] node59512;
	wire [4-1:0] node59513;
	wire [4-1:0] node59516;
	wire [4-1:0] node59517;
	wire [4-1:0] node59521;
	wire [4-1:0] node59522;
	wire [4-1:0] node59523;
	wire [4-1:0] node59528;
	wire [4-1:0] node59529;
	wire [4-1:0] node59530;
	wire [4-1:0] node59531;
	wire [4-1:0] node59536;
	wire [4-1:0] node59537;
	wire [4-1:0] node59538;
	wire [4-1:0] node59542;
	wire [4-1:0] node59545;
	wire [4-1:0] node59546;
	wire [4-1:0] node59547;
	wire [4-1:0] node59548;
	wire [4-1:0] node59549;
	wire [4-1:0] node59550;
	wire [4-1:0] node59552;
	wire [4-1:0] node59555;
	wire [4-1:0] node59557;
	wire [4-1:0] node59560;
	wire [4-1:0] node59562;
	wire [4-1:0] node59564;
	wire [4-1:0] node59567;
	wire [4-1:0] node59568;
	wire [4-1:0] node59569;
	wire [4-1:0] node59570;
	wire [4-1:0] node59573;
	wire [4-1:0] node59577;
	wire [4-1:0] node59578;
	wire [4-1:0] node59581;
	wire [4-1:0] node59584;
	wire [4-1:0] node59585;
	wire [4-1:0] node59586;
	wire [4-1:0] node59588;
	wire [4-1:0] node59591;
	wire [4-1:0] node59592;
	wire [4-1:0] node59596;
	wire [4-1:0] node59597;
	wire [4-1:0] node59598;
	wire [4-1:0] node59599;
	wire [4-1:0] node59602;
	wire [4-1:0] node59606;
	wire [4-1:0] node59607;
	wire [4-1:0] node59610;
	wire [4-1:0] node59611;
	wire [4-1:0] node59615;
	wire [4-1:0] node59616;
	wire [4-1:0] node59617;
	wire [4-1:0] node59618;
	wire [4-1:0] node59619;
	wire [4-1:0] node59622;
	wire [4-1:0] node59625;
	wire [4-1:0] node59626;
	wire [4-1:0] node59628;
	wire [4-1:0] node59631;
	wire [4-1:0] node59633;
	wire [4-1:0] node59636;
	wire [4-1:0] node59637;
	wire [4-1:0] node59638;
	wire [4-1:0] node59639;
	wire [4-1:0] node59642;
	wire [4-1:0] node59646;
	wire [4-1:0] node59647;
	wire [4-1:0] node59648;
	wire [4-1:0] node59651;
	wire [4-1:0] node59655;
	wire [4-1:0] node59656;
	wire [4-1:0] node59657;
	wire [4-1:0] node59658;
	wire [4-1:0] node59659;
	wire [4-1:0] node59663;
	wire [4-1:0] node59666;
	wire [4-1:0] node59667;
	wire [4-1:0] node59670;
	wire [4-1:0] node59673;
	wire [4-1:0] node59674;
	wire [4-1:0] node59676;
	wire [4-1:0] node59677;
	wire [4-1:0] node59680;
	wire [4-1:0] node59683;
	wire [4-1:0] node59684;
	wire [4-1:0] node59688;
	wire [4-1:0] node59689;
	wire [4-1:0] node59690;
	wire [4-1:0] node59691;
	wire [4-1:0] node59692;
	wire [4-1:0] node59693;
	wire [4-1:0] node59694;
	wire [4-1:0] node59695;
	wire [4-1:0] node59697;
	wire [4-1:0] node59699;
	wire [4-1:0] node59701;
	wire [4-1:0] node59704;
	wire [4-1:0] node59705;
	wire [4-1:0] node59706;
	wire [4-1:0] node59708;
	wire [4-1:0] node59712;
	wire [4-1:0] node59713;
	wire [4-1:0] node59715;
	wire [4-1:0] node59719;
	wire [4-1:0] node59720;
	wire [4-1:0] node59721;
	wire [4-1:0] node59724;
	wire [4-1:0] node59727;
	wire [4-1:0] node59729;
	wire [4-1:0] node59730;
	wire [4-1:0] node59732;
	wire [4-1:0] node59736;
	wire [4-1:0] node59737;
	wire [4-1:0] node59738;
	wire [4-1:0] node59739;
	wire [4-1:0] node59741;
	wire [4-1:0] node59743;
	wire [4-1:0] node59746;
	wire [4-1:0] node59747;
	wire [4-1:0] node59750;
	wire [4-1:0] node59753;
	wire [4-1:0] node59754;
	wire [4-1:0] node59755;
	wire [4-1:0] node59756;
	wire [4-1:0] node59759;
	wire [4-1:0] node59763;
	wire [4-1:0] node59765;
	wire [4-1:0] node59767;
	wire [4-1:0] node59770;
	wire [4-1:0] node59771;
	wire [4-1:0] node59772;
	wire [4-1:0] node59773;
	wire [4-1:0] node59775;
	wire [4-1:0] node59778;
	wire [4-1:0] node59781;
	wire [4-1:0] node59782;
	wire [4-1:0] node59785;
	wire [4-1:0] node59788;
	wire [4-1:0] node59790;
	wire [4-1:0] node59792;
	wire [4-1:0] node59793;
	wire [4-1:0] node59797;
	wire [4-1:0] node59798;
	wire [4-1:0] node59799;
	wire [4-1:0] node59800;
	wire [4-1:0] node59801;
	wire [4-1:0] node59804;
	wire [4-1:0] node59805;
	wire [4-1:0] node59809;
	wire [4-1:0] node59810;
	wire [4-1:0] node59811;
	wire [4-1:0] node59813;
	wire [4-1:0] node59816;
	wire [4-1:0] node59818;
	wire [4-1:0] node59821;
	wire [4-1:0] node59822;
	wire [4-1:0] node59824;
	wire [4-1:0] node59827;
	wire [4-1:0] node59830;
	wire [4-1:0] node59831;
	wire [4-1:0] node59832;
	wire [4-1:0] node59834;
	wire [4-1:0] node59837;
	wire [4-1:0] node59839;
	wire [4-1:0] node59842;
	wire [4-1:0] node59843;
	wire [4-1:0] node59845;
	wire [4-1:0] node59848;
	wire [4-1:0] node59850;
	wire [4-1:0] node59853;
	wire [4-1:0] node59854;
	wire [4-1:0] node59855;
	wire [4-1:0] node59856;
	wire [4-1:0] node59859;
	wire [4-1:0] node59861;
	wire [4-1:0] node59864;
	wire [4-1:0] node59865;
	wire [4-1:0] node59867;
	wire [4-1:0] node59870;
	wire [4-1:0] node59872;
	wire [4-1:0] node59875;
	wire [4-1:0] node59876;
	wire [4-1:0] node59877;
	wire [4-1:0] node59878;
	wire [4-1:0] node59881;
	wire [4-1:0] node59884;
	wire [4-1:0] node59885;
	wire [4-1:0] node59886;
	wire [4-1:0] node59889;
	wire [4-1:0] node59893;
	wire [4-1:0] node59894;
	wire [4-1:0] node59895;
	wire [4-1:0] node59898;
	wire [4-1:0] node59901;
	wire [4-1:0] node59903;
	wire [4-1:0] node59906;
	wire [4-1:0] node59907;
	wire [4-1:0] node59908;
	wire [4-1:0] node59909;
	wire [4-1:0] node59910;
	wire [4-1:0] node59911;
	wire [4-1:0] node59914;
	wire [4-1:0] node59917;
	wire [4-1:0] node59918;
	wire [4-1:0] node59919;
	wire [4-1:0] node59921;
	wire [4-1:0] node59924;
	wire [4-1:0] node59927;
	wire [4-1:0] node59928;
	wire [4-1:0] node59931;
	wire [4-1:0] node59934;
	wire [4-1:0] node59935;
	wire [4-1:0] node59936;
	wire [4-1:0] node59938;
	wire [4-1:0] node59941;
	wire [4-1:0] node59944;
	wire [4-1:0] node59945;
	wire [4-1:0] node59949;
	wire [4-1:0] node59950;
	wire [4-1:0] node59951;
	wire [4-1:0] node59953;
	wire [4-1:0] node59956;
	wire [4-1:0] node59958;
	wire [4-1:0] node59961;
	wire [4-1:0] node59962;
	wire [4-1:0] node59964;
	wire [4-1:0] node59967;
	wire [4-1:0] node59969;
	wire [4-1:0] node59972;
	wire [4-1:0] node59973;
	wire [4-1:0] node59974;
	wire [4-1:0] node59975;
	wire [4-1:0] node59976;
	wire [4-1:0] node59979;
	wire [4-1:0] node59982;
	wire [4-1:0] node59983;
	wire [4-1:0] node59984;
	wire [4-1:0] node59987;
	wire [4-1:0] node59990;
	wire [4-1:0] node59991;
	wire [4-1:0] node59992;
	wire [4-1:0] node59995;
	wire [4-1:0] node59999;
	wire [4-1:0] node60000;
	wire [4-1:0] node60001;
	wire [4-1:0] node60003;
	wire [4-1:0] node60004;
	wire [4-1:0] node60007;
	wire [4-1:0] node60010;
	wire [4-1:0] node60012;
	wire [4-1:0] node60015;
	wire [4-1:0] node60016;
	wire [4-1:0] node60017;
	wire [4-1:0] node60020;
	wire [4-1:0] node60023;
	wire [4-1:0] node60024;
	wire [4-1:0] node60026;
	wire [4-1:0] node60030;
	wire [4-1:0] node60031;
	wire [4-1:0] node60032;
	wire [4-1:0] node60034;
	wire [4-1:0] node60037;
	wire [4-1:0] node60039;
	wire [4-1:0] node60042;
	wire [4-1:0] node60043;
	wire [4-1:0] node60045;
	wire [4-1:0] node60048;
	wire [4-1:0] node60050;
	wire [4-1:0] node60053;
	wire [4-1:0] node60054;
	wire [4-1:0] node60055;
	wire [4-1:0] node60056;
	wire [4-1:0] node60057;
	wire [4-1:0] node60058;
	wire [4-1:0] node60059;
	wire [4-1:0] node60060;
	wire [4-1:0] node60061;
	wire [4-1:0] node60065;
	wire [4-1:0] node60068;
	wire [4-1:0] node60069;
	wire [4-1:0] node60072;
	wire [4-1:0] node60075;
	wire [4-1:0] node60076;
	wire [4-1:0] node60077;
	wire [4-1:0] node60078;
	wire [4-1:0] node60082;
	wire [4-1:0] node60084;
	wire [4-1:0] node60087;
	wire [4-1:0] node60088;
	wire [4-1:0] node60091;
	wire [4-1:0] node60094;
	wire [4-1:0] node60095;
	wire [4-1:0] node60096;
	wire [4-1:0] node60097;
	wire [4-1:0] node60098;
	wire [4-1:0] node60102;
	wire [4-1:0] node60105;
	wire [4-1:0] node60107;
	wire [4-1:0] node60110;
	wire [4-1:0] node60111;
	wire [4-1:0] node60112;
	wire [4-1:0] node60113;
	wire [4-1:0] node60117;
	wire [4-1:0] node60118;
	wire [4-1:0] node60121;
	wire [4-1:0] node60124;
	wire [4-1:0] node60125;
	wire [4-1:0] node60128;
	wire [4-1:0] node60131;
	wire [4-1:0] node60132;
	wire [4-1:0] node60133;
	wire [4-1:0] node60134;
	wire [4-1:0] node60135;
	wire [4-1:0] node60137;
	wire [4-1:0] node60140;
	wire [4-1:0] node60143;
	wire [4-1:0] node60144;
	wire [4-1:0] node60145;
	wire [4-1:0] node60150;
	wire [4-1:0] node60151;
	wire [4-1:0] node60152;
	wire [4-1:0] node60153;
	wire [4-1:0] node60156;
	wire [4-1:0] node60159;
	wire [4-1:0] node60161;
	wire [4-1:0] node60164;
	wire [4-1:0] node60166;
	wire [4-1:0] node60168;
	wire [4-1:0] node60171;
	wire [4-1:0] node60172;
	wire [4-1:0] node60173;
	wire [4-1:0] node60174;
	wire [4-1:0] node60178;
	wire [4-1:0] node60179;
	wire [4-1:0] node60182;
	wire [4-1:0] node60185;
	wire [4-1:0] node60186;
	wire [4-1:0] node60187;
	wire [4-1:0] node60188;
	wire [4-1:0] node60191;
	wire [4-1:0] node60195;
	wire [4-1:0] node60197;
	wire [4-1:0] node60200;
	wire [4-1:0] node60201;
	wire [4-1:0] node60202;
	wire [4-1:0] node60203;
	wire [4-1:0] node60204;
	wire [4-1:0] node60206;
	wire [4-1:0] node60207;
	wire [4-1:0] node60210;
	wire [4-1:0] node60214;
	wire [4-1:0] node60215;
	wire [4-1:0] node60216;
	wire [4-1:0] node60217;
	wire [4-1:0] node60220;
	wire [4-1:0] node60223;
	wire [4-1:0] node60225;
	wire [4-1:0] node60228;
	wire [4-1:0] node60229;
	wire [4-1:0] node60233;
	wire [4-1:0] node60234;
	wire [4-1:0] node60235;
	wire [4-1:0] node60236;
	wire [4-1:0] node60237;
	wire [4-1:0] node60242;
	wire [4-1:0] node60243;
	wire [4-1:0] node60244;
	wire [4-1:0] node60248;
	wire [4-1:0] node60249;
	wire [4-1:0] node60253;
	wire [4-1:0] node60254;
	wire [4-1:0] node60258;
	wire [4-1:0] node60259;
	wire [4-1:0] node60260;
	wire [4-1:0] node60261;
	wire [4-1:0] node60262;
	wire [4-1:0] node60264;
	wire [4-1:0] node60267;
	wire [4-1:0] node60269;
	wire [4-1:0] node60272;
	wire [4-1:0] node60275;
	wire [4-1:0] node60276;
	wire [4-1:0] node60279;
	wire [4-1:0] node60280;
	wire [4-1:0] node60281;
	wire [4-1:0] node60286;
	wire [4-1:0] node60287;
	wire [4-1:0] node60288;
	wire [4-1:0] node60289;
	wire [4-1:0] node60290;
	wire [4-1:0] node60293;
	wire [4-1:0] node60297;
	wire [4-1:0] node60298;
	wire [4-1:0] node60301;
	wire [4-1:0] node60302;
	wire [4-1:0] node60305;
	wire [4-1:0] node60308;
	wire [4-1:0] node60309;
	wire [4-1:0] node60310;
	wire [4-1:0] node60312;
	wire [4-1:0] node60315;
	wire [4-1:0] node60316;
	wire [4-1:0] node60319;
	wire [4-1:0] node60322;
	wire [4-1:0] node60323;
	wire [4-1:0] node60324;
	wire [4-1:0] node60327;
	wire [4-1:0] node60331;
	wire [4-1:0] node60332;
	wire [4-1:0] node60333;
	wire [4-1:0] node60334;
	wire [4-1:0] node60335;
	wire [4-1:0] node60336;
	wire [4-1:0] node60337;
	wire [4-1:0] node60340;
	wire [4-1:0] node60343;
	wire [4-1:0] node60344;
	wire [4-1:0] node60345;
	wire [4-1:0] node60348;
	wire [4-1:0] node60352;
	wire [4-1:0] node60353;
	wire [4-1:0] node60355;
	wire [4-1:0] node60357;
	wire [4-1:0] node60360;
	wire [4-1:0] node60361;
	wire [4-1:0] node60363;
	wire [4-1:0] node60366;
	wire [4-1:0] node60367;
	wire [4-1:0] node60370;
	wire [4-1:0] node60373;
	wire [4-1:0] node60374;
	wire [4-1:0] node60375;
	wire [4-1:0] node60376;
	wire [4-1:0] node60378;
	wire [4-1:0] node60381;
	wire [4-1:0] node60382;
	wire [4-1:0] node60385;
	wire [4-1:0] node60388;
	wire [4-1:0] node60389;
	wire [4-1:0] node60391;
	wire [4-1:0] node60395;
	wire [4-1:0] node60396;
	wire [4-1:0] node60398;
	wire [4-1:0] node60399;
	wire [4-1:0] node60404;
	wire [4-1:0] node60405;
	wire [4-1:0] node60406;
	wire [4-1:0] node60407;
	wire [4-1:0] node60408;
	wire [4-1:0] node60409;
	wire [4-1:0] node60413;
	wire [4-1:0] node60414;
	wire [4-1:0] node60418;
	wire [4-1:0] node60421;
	wire [4-1:0] node60422;
	wire [4-1:0] node60423;
	wire [4-1:0] node60426;
	wire [4-1:0] node60429;
	wire [4-1:0] node60430;
	wire [4-1:0] node60431;
	wire [4-1:0] node60434;
	wire [4-1:0] node60437;
	wire [4-1:0] node60440;
	wire [4-1:0] node60441;
	wire [4-1:0] node60442;
	wire [4-1:0] node60444;
	wire [4-1:0] node60446;
	wire [4-1:0] node60449;
	wire [4-1:0] node60450;
	wire [4-1:0] node60453;
	wire [4-1:0] node60455;
	wire [4-1:0] node60458;
	wire [4-1:0] node60459;
	wire [4-1:0] node60460;
	wire [4-1:0] node60462;
	wire [4-1:0] node60465;
	wire [4-1:0] node60467;
	wire [4-1:0] node60470;
	wire [4-1:0] node60472;
	wire [4-1:0] node60473;
	wire [4-1:0] node60476;
	wire [4-1:0] node60479;
	wire [4-1:0] node60480;
	wire [4-1:0] node60481;
	wire [4-1:0] node60482;
	wire [4-1:0] node60485;
	wire [4-1:0] node60488;
	wire [4-1:0] node60489;
	wire [4-1:0] node60490;
	wire [4-1:0] node60491;
	wire [4-1:0] node60492;
	wire [4-1:0] node60496;
	wire [4-1:0] node60498;
	wire [4-1:0] node60501;
	wire [4-1:0] node60502;
	wire [4-1:0] node60503;
	wire [4-1:0] node60506;
	wire [4-1:0] node60509;
	wire [4-1:0] node60511;
	wire [4-1:0] node60514;
	wire [4-1:0] node60515;
	wire [4-1:0] node60518;
	wire [4-1:0] node60521;
	wire [4-1:0] node60522;
	wire [4-1:0] node60523;
	wire [4-1:0] node60524;
	wire [4-1:0] node60527;
	wire [4-1:0] node60530;
	wire [4-1:0] node60531;
	wire [4-1:0] node60533;
	wire [4-1:0] node60534;
	wire [4-1:0] node60537;
	wire [4-1:0] node60540;
	wire [4-1:0] node60542;
	wire [4-1:0] node60544;
	wire [4-1:0] node60547;
	wire [4-1:0] node60548;
	wire [4-1:0] node60551;
	wire [4-1:0] node60554;
	wire [4-1:0] node60555;
	wire [4-1:0] node60556;
	wire [4-1:0] node60557;
	wire [4-1:0] node60558;
	wire [4-1:0] node60559;
	wire [4-1:0] node60560;
	wire [4-1:0] node60561;
	wire [4-1:0] node60562;
	wire [4-1:0] node60566;
	wire [4-1:0] node60567;
	wire [4-1:0] node60571;
	wire [4-1:0] node60572;
	wire [4-1:0] node60573;
	wire [4-1:0] node60574;
	wire [4-1:0] node60578;
	wire [4-1:0] node60580;
	wire [4-1:0] node60584;
	wire [4-1:0] node60585;
	wire [4-1:0] node60586;
	wire [4-1:0] node60589;
	wire [4-1:0] node60590;
	wire [4-1:0] node60594;
	wire [4-1:0] node60595;
	wire [4-1:0] node60596;
	wire [4-1:0] node60597;
	wire [4-1:0] node60601;
	wire [4-1:0] node60602;
	wire [4-1:0] node60605;
	wire [4-1:0] node60609;
	wire [4-1:0] node60610;
	wire [4-1:0] node60611;
	wire [4-1:0] node60612;
	wire [4-1:0] node60613;
	wire [4-1:0] node60614;
	wire [4-1:0] node60617;
	wire [4-1:0] node60620;
	wire [4-1:0] node60622;
	wire [4-1:0] node60625;
	wire [4-1:0] node60626;
	wire [4-1:0] node60630;
	wire [4-1:0] node60631;
	wire [4-1:0] node60632;
	wire [4-1:0] node60633;
	wire [4-1:0] node60637;
	wire [4-1:0] node60638;
	wire [4-1:0] node60641;
	wire [4-1:0] node60644;
	wire [4-1:0] node60645;
	wire [4-1:0] node60647;
	wire [4-1:0] node60651;
	wire [4-1:0] node60652;
	wire [4-1:0] node60653;
	wire [4-1:0] node60656;
	wire [4-1:0] node60659;
	wire [4-1:0] node60661;
	wire [4-1:0] node60662;
	wire [4-1:0] node60665;
	wire [4-1:0] node60668;
	wire [4-1:0] node60669;
	wire [4-1:0] node60670;
	wire [4-1:0] node60671;
	wire [4-1:0] node60673;
	wire [4-1:0] node60674;
	wire [4-1:0] node60678;
	wire [4-1:0] node60680;
	wire [4-1:0] node60681;
	wire [4-1:0] node60682;
	wire [4-1:0] node60687;
	wire [4-1:0] node60688;
	wire [4-1:0] node60689;
	wire [4-1:0] node60690;
	wire [4-1:0] node60694;
	wire [4-1:0] node60695;
	wire [4-1:0] node60699;
	wire [4-1:0] node60700;
	wire [4-1:0] node60701;
	wire [4-1:0] node60706;
	wire [4-1:0] node60707;
	wire [4-1:0] node60708;
	wire [4-1:0] node60709;
	wire [4-1:0] node60710;
	wire [4-1:0] node60712;
	wire [4-1:0] node60715;
	wire [4-1:0] node60716;
	wire [4-1:0] node60720;
	wire [4-1:0] node60721;
	wire [4-1:0] node60722;
	wire [4-1:0] node60725;
	wire [4-1:0] node60728;
	wire [4-1:0] node60730;
	wire [4-1:0] node60733;
	wire [4-1:0] node60734;
	wire [4-1:0] node60737;
	wire [4-1:0] node60740;
	wire [4-1:0] node60741;
	wire [4-1:0] node60742;
	wire [4-1:0] node60745;
	wire [4-1:0] node60748;
	wire [4-1:0] node60749;
	wire [4-1:0] node60750;
	wire [4-1:0] node60754;
	wire [4-1:0] node60755;
	wire [4-1:0] node60758;
	wire [4-1:0] node60761;
	wire [4-1:0] node60762;
	wire [4-1:0] node60763;
	wire [4-1:0] node60764;
	wire [4-1:0] node60765;
	wire [4-1:0] node60766;
	wire [4-1:0] node60767;
	wire [4-1:0] node60768;
	wire [4-1:0] node60771;
	wire [4-1:0] node60774;
	wire [4-1:0] node60776;
	wire [4-1:0] node60780;
	wire [4-1:0] node60782;
	wire [4-1:0] node60783;
	wire [4-1:0] node60784;
	wire [4-1:0] node60788;
	wire [4-1:0] node60789;
	wire [4-1:0] node60793;
	wire [4-1:0] node60794;
	wire [4-1:0] node60795;
	wire [4-1:0] node60796;
	wire [4-1:0] node60799;
	wire [4-1:0] node60802;
	wire [4-1:0] node60803;
	wire [4-1:0] node60807;
	wire [4-1:0] node60808;
	wire [4-1:0] node60811;
	wire [4-1:0] node60814;
	wire [4-1:0] node60815;
	wire [4-1:0] node60816;
	wire [4-1:0] node60817;
	wire [4-1:0] node60821;
	wire [4-1:0] node60822;
	wire [4-1:0] node60826;
	wire [4-1:0] node60827;
	wire [4-1:0] node60828;
	wire [4-1:0] node60832;
	wire [4-1:0] node60833;
	wire [4-1:0] node60837;
	wire [4-1:0] node60838;
	wire [4-1:0] node60839;
	wire [4-1:0] node60840;
	wire [4-1:0] node60841;
	wire [4-1:0] node60842;
	wire [4-1:0] node60846;
	wire [4-1:0] node60847;
	wire [4-1:0] node60851;
	wire [4-1:0] node60853;
	wire [4-1:0] node60854;
	wire [4-1:0] node60858;
	wire [4-1:0] node60859;
	wire [4-1:0] node60860;
	wire [4-1:0] node60862;
	wire [4-1:0] node60863;
	wire [4-1:0] node60866;
	wire [4-1:0] node60869;
	wire [4-1:0] node60870;
	wire [4-1:0] node60871;
	wire [4-1:0] node60875;
	wire [4-1:0] node60876;
	wire [4-1:0] node60880;
	wire [4-1:0] node60881;
	wire [4-1:0] node60882;
	wire [4-1:0] node60883;
	wire [4-1:0] node60886;
	wire [4-1:0] node60890;
	wire [4-1:0] node60891;
	wire [4-1:0] node60892;
	wire [4-1:0] node60897;
	wire [4-1:0] node60898;
	wire [4-1:0] node60899;
	wire [4-1:0] node60900;
	wire [4-1:0] node60901;
	wire [4-1:0] node60905;
	wire [4-1:0] node60906;
	wire [4-1:0] node60910;
	wire [4-1:0] node60911;
	wire [4-1:0] node60914;
	wire [4-1:0] node60915;
	wire [4-1:0] node60919;
	wire [4-1:0] node60920;
	wire [4-1:0] node60921;
	wire [4-1:0] node60923;
	wire [4-1:0] node60924;
	wire [4-1:0] node60928;
	wire [4-1:0] node60930;
	wire [4-1:0] node60931;
	wire [4-1:0] node60935;
	wire [4-1:0] node60936;
	wire [4-1:0] node60937;
	wire [4-1:0] node60938;
	wire [4-1:0] node60942;
	wire [4-1:0] node60943;
	wire [4-1:0] node60947;
	wire [4-1:0] node60949;
	wire [4-1:0] node60952;
	wire [4-1:0] node60953;
	wire [4-1:0] node60954;
	wire [4-1:0] node60955;
	wire [4-1:0] node60956;
	wire [4-1:0] node60957;
	wire [4-1:0] node60958;
	wire [4-1:0] node60959;
	wire [4-1:0] node60961;
	wire [4-1:0] node60964;
	wire [4-1:0] node60966;
	wire [4-1:0] node60969;
	wire [4-1:0] node60971;
	wire [4-1:0] node60973;
	wire [4-1:0] node60976;
	wire [4-1:0] node60977;
	wire [4-1:0] node60979;
	wire [4-1:0] node60980;
	wire [4-1:0] node60983;
	wire [4-1:0] node60986;
	wire [4-1:0] node60987;
	wire [4-1:0] node60990;
	wire [4-1:0] node60993;
	wire [4-1:0] node60994;
	wire [4-1:0] node60995;
	wire [4-1:0] node60996;
	wire [4-1:0] node60999;
	wire [4-1:0] node61000;
	wire [4-1:0] node61004;
	wire [4-1:0] node61006;
	wire [4-1:0] node61009;
	wire [4-1:0] node61010;
	wire [4-1:0] node61011;
	wire [4-1:0] node61014;
	wire [4-1:0] node61017;
	wire [4-1:0] node61019;
	wire [4-1:0] node61022;
	wire [4-1:0] node61023;
	wire [4-1:0] node61024;
	wire [4-1:0] node61025;
	wire [4-1:0] node61026;
	wire [4-1:0] node61030;
	wire [4-1:0] node61031;
	wire [4-1:0] node61032;
	wire [4-1:0] node61037;
	wire [4-1:0] node61038;
	wire [4-1:0] node61039;
	wire [4-1:0] node61043;
	wire [4-1:0] node61044;
	wire [4-1:0] node61045;
	wire [4-1:0] node61048;
	wire [4-1:0] node61052;
	wire [4-1:0] node61053;
	wire [4-1:0] node61054;
	wire [4-1:0] node61056;
	wire [4-1:0] node61059;
	wire [4-1:0] node61060;
	wire [4-1:0] node61063;
	wire [4-1:0] node61065;
	wire [4-1:0] node61068;
	wire [4-1:0] node61069;
	wire [4-1:0] node61071;
	wire [4-1:0] node61072;
	wire [4-1:0] node61077;
	wire [4-1:0] node61078;
	wire [4-1:0] node61079;
	wire [4-1:0] node61080;
	wire [4-1:0] node61081;
	wire [4-1:0] node61082;
	wire [4-1:0] node61085;
	wire [4-1:0] node61088;
	wire [4-1:0] node61089;
	wire [4-1:0] node61092;
	wire [4-1:0] node61095;
	wire [4-1:0] node61096;
	wire [4-1:0] node61097;
	wire [4-1:0] node61098;
	wire [4-1:0] node61101;
	wire [4-1:0] node61104;
	wire [4-1:0] node61105;
	wire [4-1:0] node61109;
	wire [4-1:0] node61110;
	wire [4-1:0] node61114;
	wire [4-1:0] node61115;
	wire [4-1:0] node61116;
	wire [4-1:0] node61117;
	wire [4-1:0] node61118;
	wire [4-1:0] node61121;
	wire [4-1:0] node61125;
	wire [4-1:0] node61126;
	wire [4-1:0] node61128;
	wire [4-1:0] node61131;
	wire [4-1:0] node61133;
	wire [4-1:0] node61136;
	wire [4-1:0] node61137;
	wire [4-1:0] node61138;
	wire [4-1:0] node61142;
	wire [4-1:0] node61143;
	wire [4-1:0] node61146;
	wire [4-1:0] node61149;
	wire [4-1:0] node61150;
	wire [4-1:0] node61151;
	wire [4-1:0] node61152;
	wire [4-1:0] node61153;
	wire [4-1:0] node61156;
	wire [4-1:0] node61159;
	wire [4-1:0] node61160;
	wire [4-1:0] node61164;
	wire [4-1:0] node61166;
	wire [4-1:0] node61168;
	wire [4-1:0] node61169;
	wire [4-1:0] node61172;
	wire [4-1:0] node61175;
	wire [4-1:0] node61176;
	wire [4-1:0] node61177;
	wire [4-1:0] node61180;
	wire [4-1:0] node61183;
	wire [4-1:0] node61184;
	wire [4-1:0] node61186;
	wire [4-1:0] node61187;
	wire [4-1:0] node61190;
	wire [4-1:0] node61193;
	wire [4-1:0] node61194;
	wire [4-1:0] node61195;
	wire [4-1:0] node61198;
	wire [4-1:0] node61202;
	wire [4-1:0] node61203;
	wire [4-1:0] node61204;
	wire [4-1:0] node61205;
	wire [4-1:0] node61206;
	wire [4-1:0] node61207;
	wire [4-1:0] node61208;
	wire [4-1:0] node61209;
	wire [4-1:0] node61212;
	wire [4-1:0] node61215;
	wire [4-1:0] node61218;
	wire [4-1:0] node61219;
	wire [4-1:0] node61221;
	wire [4-1:0] node61225;
	wire [4-1:0] node61226;
	wire [4-1:0] node61227;
	wire [4-1:0] node61229;
	wire [4-1:0] node61232;
	wire [4-1:0] node61234;
	wire [4-1:0] node61237;
	wire [4-1:0] node61238;
	wire [4-1:0] node61241;
	wire [4-1:0] node61244;
	wire [4-1:0] node61245;
	wire [4-1:0] node61246;
	wire [4-1:0] node61247;
	wire [4-1:0] node61248;
	wire [4-1:0] node61251;
	wire [4-1:0] node61254;
	wire [4-1:0] node61255;
	wire [4-1:0] node61259;
	wire [4-1:0] node61260;
	wire [4-1:0] node61264;
	wire [4-1:0] node61265;
	wire [4-1:0] node61267;
	wire [4-1:0] node61268;
	wire [4-1:0] node61271;
	wire [4-1:0] node61274;
	wire [4-1:0] node61275;
	wire [4-1:0] node61278;
	wire [4-1:0] node61281;
	wire [4-1:0] node61282;
	wire [4-1:0] node61283;
	wire [4-1:0] node61284;
	wire [4-1:0] node61285;
	wire [4-1:0] node61286;
	wire [4-1:0] node61290;
	wire [4-1:0] node61291;
	wire [4-1:0] node61295;
	wire [4-1:0] node61296;
	wire [4-1:0] node61297;
	wire [4-1:0] node61302;
	wire [4-1:0] node61303;
	wire [4-1:0] node61304;
	wire [4-1:0] node61306;
	wire [4-1:0] node61309;
	wire [4-1:0] node61310;
	wire [4-1:0] node61314;
	wire [4-1:0] node61315;
	wire [4-1:0] node61318;
	wire [4-1:0] node61321;
	wire [4-1:0] node61322;
	wire [4-1:0] node61323;
	wire [4-1:0] node61325;
	wire [4-1:0] node61328;
	wire [4-1:0] node61329;
	wire [4-1:0] node61332;
	wire [4-1:0] node61335;
	wire [4-1:0] node61336;
	wire [4-1:0] node61337;
	wire [4-1:0] node61338;
	wire [4-1:0] node61342;
	wire [4-1:0] node61345;
	wire [4-1:0] node61347;
	wire [4-1:0] node61350;
	wire [4-1:0] node61351;
	wire [4-1:0] node61352;
	wire [4-1:0] node61353;
	wire [4-1:0] node61354;
	wire [4-1:0] node61355;
	wire [4-1:0] node61358;
	wire [4-1:0] node61361;
	wire [4-1:0] node61363;
	wire [4-1:0] node61364;
	wire [4-1:0] node61368;
	wire [4-1:0] node61369;
	wire [4-1:0] node61373;
	wire [4-1:0] node61374;
	wire [4-1:0] node61375;
	wire [4-1:0] node61377;
	wire [4-1:0] node61380;
	wire [4-1:0] node61383;
	wire [4-1:0] node61384;
	wire [4-1:0] node61387;
	wire [4-1:0] node61390;
	wire [4-1:0] node61391;
	wire [4-1:0] node61392;
	wire [4-1:0] node61393;
	wire [4-1:0] node61395;
	wire [4-1:0] node61398;
	wire [4-1:0] node61400;
	wire [4-1:0] node61403;
	wire [4-1:0] node61404;
	wire [4-1:0] node61405;
	wire [4-1:0] node61408;
	wire [4-1:0] node61411;
	wire [4-1:0] node61412;
	wire [4-1:0] node61413;
	wire [4-1:0] node61417;
	wire [4-1:0] node61418;
	wire [4-1:0] node61421;
	wire [4-1:0] node61424;
	wire [4-1:0] node61425;
	wire [4-1:0] node61426;
	wire [4-1:0] node61427;
	wire [4-1:0] node61428;
	wire [4-1:0] node61431;
	wire [4-1:0] node61436;
	wire [4-1:0] node61437;
	wire [4-1:0] node61440;

	assign outp = (inp[10]) ? node31192 : node1;
		assign node1 = (inp[6]) ? node14923 : node2;
			assign node2 = (inp[11]) ? node6792 : node3;
				assign node3 = (inp[1]) ? node3427 : node4;
					assign node4 = (inp[13]) ? node1948 : node5;
						assign node5 = (inp[2]) ? node975 : node6;
							assign node6 = (inp[14]) ? node522 : node7;
								assign node7 = (inp[3]) ? node275 : node8;
									assign node8 = (inp[8]) ? node150 : node9;
										assign node9 = (inp[7]) ? node71 : node10;
											assign node10 = (inp[5]) ? node36 : node11;
												assign node11 = (inp[0]) ? node23 : node12;
													assign node12 = (inp[15]) ? node20 : node13;
														assign node13 = (inp[9]) ? node17 : node14;
															assign node14 = (inp[4]) ? 4'b1011 : 4'b1111;
															assign node17 = (inp[4]) ? 4'b1111 : 4'b1011;
														assign node20 = (inp[9]) ? 4'b1101 : 4'b1001;
													assign node23 = (inp[15]) ? 4'b1011 : node24;
														assign node24 = (inp[12]) ? node30 : node25;
															assign node25 = (inp[4]) ? 4'b1001 : node26;
																assign node26 = (inp[9]) ? 4'b1001 : 4'b1101;
															assign node30 = (inp[4]) ? 4'b1101 : node31;
																assign node31 = (inp[9]) ? 4'b1001 : 4'b1101;
												assign node36 = (inp[4]) ? node52 : node37;
													assign node37 = (inp[9]) ? node47 : node38;
														assign node38 = (inp[12]) ? node44 : node39;
															assign node39 = (inp[0]) ? node41 : 4'b1111;
																assign node41 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node44 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node47 = (inp[15]) ? node49 : 4'b1001;
															assign node49 = (inp[0]) ? 4'b1011 : 4'b1001;
													assign node52 = (inp[9]) ? node58 : node53;
														assign node53 = (inp[15]) ? node55 : 4'b1011;
															assign node55 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node58 = (inp[12]) ? node66 : node59;
															assign node59 = (inp[0]) ? node63 : node60;
																assign node60 = (inp[15]) ? 4'b1111 : 4'b1101;
																assign node63 = (inp[15]) ? 4'b1101 : 4'b1111;
															assign node66 = (inp[15]) ? 4'b1111 : node67;
																assign node67 = (inp[0]) ? 4'b1111 : 4'b1101;
											assign node71 = (inp[12]) ? node105 : node72;
												assign node72 = (inp[15]) ? node88 : node73;
													assign node73 = (inp[0]) ? node85 : node74;
														assign node74 = (inp[5]) ? node80 : node75;
															assign node75 = (inp[9]) ? 4'b1110 : node76;
																assign node76 = (inp[4]) ? 4'b1010 : 4'b1110;
															assign node80 = (inp[4]) ? 4'b1100 : node81;
																assign node81 = (inp[9]) ? 4'b1010 : 4'b1110;
														assign node85 = (inp[4]) ? 4'b1000 : 4'b1100;
													assign node88 = (inp[0]) ? node98 : node89;
														assign node89 = (inp[9]) ? node93 : node90;
															assign node90 = (inp[4]) ? 4'b1000 : 4'b1100;
															assign node93 = (inp[4]) ? node95 : 4'b1000;
																assign node95 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node98 = (inp[5]) ? node100 : 4'b1010;
															assign node100 = (inp[9]) ? 4'b1100 : node101;
																assign node101 = (inp[4]) ? 4'b1010 : 4'b1110;
												assign node105 = (inp[5]) ? node125 : node106;
													assign node106 = (inp[15]) ? node116 : node107;
														assign node107 = (inp[0]) ? 4'b1000 : node108;
															assign node108 = (inp[9]) ? node112 : node109;
																assign node109 = (inp[4]) ? 4'b1010 : 4'b1110;
																assign node112 = (inp[4]) ? 4'b1110 : 4'b1010;
														assign node116 = (inp[0]) ? node122 : node117;
															assign node117 = (inp[9]) ? node119 : 4'b1000;
																assign node119 = (inp[4]) ? 4'b1100 : 4'b1000;
															assign node122 = (inp[9]) ? 4'b1010 : 4'b1110;
													assign node125 = (inp[4]) ? node137 : node126;
														assign node126 = (inp[9]) ? node132 : node127;
															assign node127 = (inp[0]) ? node129 : 4'b1100;
																assign node129 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node132 = (inp[15]) ? node134 : 4'b1000;
																assign node134 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node137 = (inp[9]) ? node143 : node138;
															assign node138 = (inp[15]) ? node140 : 4'b1010;
																assign node140 = (inp[0]) ? 4'b1010 : 4'b1000;
															assign node143 = (inp[15]) ? node147 : node144;
																assign node144 = (inp[0]) ? 4'b1110 : 4'b1100;
																assign node147 = (inp[0]) ? 4'b1100 : 4'b1110;
										assign node150 = (inp[7]) ? node218 : node151;
											assign node151 = (inp[12]) ? node185 : node152;
												assign node152 = (inp[0]) ? node162 : node153;
													assign node153 = (inp[15]) ? 4'b1110 : node154;
														assign node154 = (inp[9]) ? node158 : node155;
															assign node155 = (inp[4]) ? 4'b1010 : 4'b1110;
															assign node158 = (inp[4]) ? 4'b1110 : 4'b1010;
													assign node162 = (inp[15]) ? node172 : node163;
														assign node163 = (inp[5]) ? node169 : node164;
															assign node164 = (inp[9]) ? node166 : 4'b1100;
																assign node166 = (inp[4]) ? 4'b1100 : 4'b1000;
															assign node169 = (inp[9]) ? 4'b1110 : 4'b1000;
														assign node172 = (inp[5]) ? node180 : node173;
															assign node173 = (inp[4]) ? node177 : node174;
																assign node174 = (inp[9]) ? 4'b1010 : 4'b1110;
																assign node177 = (inp[9]) ? 4'b1110 : 4'b1010;
															assign node180 = (inp[4]) ? 4'b1100 : node181;
																assign node181 = (inp[9]) ? 4'b1010 : 4'b1110;
												assign node185 = (inp[4]) ? node203 : node186;
													assign node186 = (inp[9]) ? node200 : node187;
														assign node187 = (inp[5]) ? node193 : node188;
															assign node188 = (inp[15]) ? node190 : 4'b1100;
																assign node190 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node193 = (inp[0]) ? node197 : node194;
																assign node194 = (inp[15]) ? 4'b1100 : 4'b1110;
																assign node197 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node200 = (inp[5]) ? 4'b1010 : 4'b1000;
													assign node203 = (inp[9]) ? node211 : node204;
														assign node204 = (inp[0]) ? node208 : node205;
															assign node205 = (inp[15]) ? 4'b1000 : 4'b1010;
															assign node208 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node211 = (inp[15]) ? node213 : 4'b1110;
															assign node213 = (inp[0]) ? 4'b1100 : node214;
																assign node214 = (inp[5]) ? 4'b1110 : 4'b1100;
											assign node218 = (inp[4]) ? node242 : node219;
												assign node219 = (inp[9]) ? node235 : node220;
													assign node220 = (inp[5]) ? node228 : node221;
														assign node221 = (inp[0]) ? node225 : node222;
															assign node222 = (inp[15]) ? 4'b1101 : 4'b1111;
															assign node225 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node228 = (inp[0]) ? node232 : node229;
															assign node229 = (inp[15]) ? 4'b1101 : 4'b1111;
															assign node232 = (inp[15]) ? 4'b1111 : 4'b1101;
													assign node235 = (inp[15]) ? node239 : node236;
														assign node236 = (inp[0]) ? 4'b1001 : 4'b1011;
														assign node239 = (inp[0]) ? 4'b1011 : 4'b1001;
												assign node242 = (inp[9]) ? node250 : node243;
													assign node243 = (inp[0]) ? node247 : node244;
														assign node244 = (inp[15]) ? 4'b1001 : 4'b1011;
														assign node247 = (inp[15]) ? 4'b1011 : 4'b1001;
													assign node250 = (inp[15]) ? node266 : node251;
														assign node251 = (inp[12]) ? node259 : node252;
															assign node252 = (inp[0]) ? node256 : node253;
																assign node253 = (inp[5]) ? 4'b1101 : 4'b1111;
																assign node256 = (inp[5]) ? 4'b1111 : 4'b1101;
															assign node259 = (inp[0]) ? node263 : node260;
																assign node260 = (inp[5]) ? 4'b1101 : 4'b1111;
																assign node263 = (inp[5]) ? 4'b1111 : 4'b1101;
														assign node266 = (inp[12]) ? node272 : node267;
															assign node267 = (inp[0]) ? 4'b1111 : node268;
																assign node268 = (inp[5]) ? 4'b1111 : 4'b1101;
															assign node272 = (inp[0]) ? 4'b1101 : 4'b1111;
									assign node275 = (inp[9]) ? node397 : node276;
										assign node276 = (inp[4]) ? node332 : node277;
											assign node277 = (inp[15]) ? node305 : node278;
												assign node278 = (inp[5]) ? node290 : node279;
													assign node279 = (inp[0]) ? node285 : node280;
														assign node280 = (inp[12]) ? node282 : 4'b1110;
															assign node282 = (inp[8]) ? 4'b1111 : 4'b1110;
														assign node285 = (inp[7]) ? 4'b1100 : node286;
															assign node286 = (inp[8]) ? 4'b1100 : 4'b1101;
													assign node290 = (inp[0]) ? node292 : 4'b1100;
														assign node292 = (inp[12]) ? node300 : node293;
															assign node293 = (inp[7]) ? node297 : node294;
																assign node294 = (inp[8]) ? 4'b1110 : 4'b1111;
																assign node297 = (inp[8]) ? 4'b1111 : 4'b1110;
															assign node300 = (inp[8]) ? 4'b1111 : node301;
																assign node301 = (inp[7]) ? 4'b1110 : 4'b1111;
												assign node305 = (inp[0]) ? node319 : node306;
													assign node306 = (inp[5]) ? node314 : node307;
														assign node307 = (inp[12]) ? node311 : node308;
															assign node308 = (inp[8]) ? 4'b1100 : 4'b1101;
															assign node311 = (inp[8]) ? 4'b1101 : 4'b1100;
														assign node314 = (inp[8]) ? 4'b1111 : node315;
															assign node315 = (inp[7]) ? 4'b1110 : 4'b1111;
													assign node319 = (inp[5]) ? node325 : node320;
														assign node320 = (inp[8]) ? 4'b1110 : node321;
															assign node321 = (inp[7]) ? 4'b1110 : 4'b1111;
														assign node325 = (inp[8]) ? node329 : node326;
															assign node326 = (inp[7]) ? 4'b1100 : 4'b1101;
															assign node329 = (inp[7]) ? 4'b1101 : 4'b1100;
											assign node332 = (inp[0]) ? node366 : node333;
												assign node333 = (inp[15]) ? node351 : node334;
													assign node334 = (inp[5]) ? node344 : node335;
														assign node335 = (inp[12]) ? 4'b1010 : node336;
															assign node336 = (inp[8]) ? node340 : node337;
																assign node337 = (inp[7]) ? 4'b1010 : 4'b1011;
																assign node340 = (inp[7]) ? 4'b1011 : 4'b1010;
														assign node344 = (inp[7]) ? node348 : node345;
															assign node345 = (inp[8]) ? 4'b1000 : 4'b1001;
															assign node348 = (inp[8]) ? 4'b1001 : 4'b1000;
													assign node351 = (inp[5]) ? node359 : node352;
														assign node352 = (inp[7]) ? node356 : node353;
															assign node353 = (inp[8]) ? 4'b1000 : 4'b1001;
															assign node356 = (inp[8]) ? 4'b1001 : 4'b1000;
														assign node359 = (inp[7]) ? node363 : node360;
															assign node360 = (inp[8]) ? 4'b1010 : 4'b1011;
															assign node363 = (inp[8]) ? 4'b1011 : 4'b1010;
												assign node366 = (inp[8]) ? node378 : node367;
													assign node367 = (inp[7]) ? node373 : node368;
														assign node368 = (inp[5]) ? node370 : 4'b1011;
															assign node370 = (inp[15]) ? 4'b1001 : 4'b1011;
														assign node373 = (inp[15]) ? node375 : 4'b1010;
															assign node375 = (inp[5]) ? 4'b1000 : 4'b1010;
													assign node378 = (inp[7]) ? node386 : node379;
														assign node379 = (inp[15]) ? node383 : node380;
															assign node380 = (inp[5]) ? 4'b1010 : 4'b1000;
															assign node383 = (inp[5]) ? 4'b1000 : 4'b1010;
														assign node386 = (inp[12]) ? node392 : node387;
															assign node387 = (inp[15]) ? 4'b1011 : node388;
																assign node388 = (inp[5]) ? 4'b1011 : 4'b1001;
															assign node392 = (inp[15]) ? node394 : 4'b1011;
																assign node394 = (inp[5]) ? 4'b1001 : 4'b1011;
										assign node397 = (inp[4]) ? node473 : node398;
											assign node398 = (inp[0]) ? node432 : node399;
												assign node399 = (inp[8]) ? node419 : node400;
													assign node400 = (inp[7]) ? node414 : node401;
														assign node401 = (inp[12]) ? node407 : node402;
															assign node402 = (inp[5]) ? node404 : 4'b1001;
																assign node404 = (inp[15]) ? 4'b1011 : 4'b1001;
															assign node407 = (inp[5]) ? node411 : node408;
																assign node408 = (inp[15]) ? 4'b1001 : 4'b1011;
																assign node411 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node414 = (inp[12]) ? 4'b1010 : node415;
															assign node415 = (inp[5]) ? 4'b1000 : 4'b1010;
													assign node419 = (inp[7]) ? node425 : node420;
														assign node420 = (inp[15]) ? node422 : 4'b1000;
															assign node422 = (inp[12]) ? 4'b1000 : 4'b1010;
														assign node425 = (inp[5]) ? node429 : node426;
															assign node426 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node429 = (inp[15]) ? 4'b1011 : 4'b1001;
												assign node432 = (inp[12]) ? node454 : node433;
													assign node433 = (inp[5]) ? node441 : node434;
														assign node434 = (inp[15]) ? node436 : 4'b1000;
															assign node436 = (inp[8]) ? node438 : 4'b1010;
																assign node438 = (inp[7]) ? 4'b1011 : 4'b1010;
														assign node441 = (inp[15]) ? node447 : node442;
															assign node442 = (inp[8]) ? node444 : 4'b1011;
																assign node444 = (inp[7]) ? 4'b1011 : 4'b1010;
															assign node447 = (inp[8]) ? node451 : node448;
																assign node448 = (inp[7]) ? 4'b1000 : 4'b1001;
																assign node451 = (inp[7]) ? 4'b1001 : 4'b1000;
													assign node454 = (inp[7]) ? node462 : node455;
														assign node455 = (inp[5]) ? node459 : node456;
															assign node456 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node459 = (inp[15]) ? 4'b1000 : 4'b1010;
														assign node462 = (inp[8]) ? node470 : node463;
															assign node463 = (inp[15]) ? node467 : node464;
																assign node464 = (inp[5]) ? 4'b1010 : 4'b1000;
																assign node467 = (inp[5]) ? 4'b1000 : 4'b1010;
															assign node470 = (inp[15]) ? 4'b1011 : 4'b1001;
											assign node473 = (inp[7]) ? node499 : node474;
												assign node474 = (inp[8]) ? node484 : node475;
													assign node475 = (inp[5]) ? 4'b1111 : node476;
														assign node476 = (inp[0]) ? node480 : node477;
															assign node477 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node480 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node484 = (inp[12]) ? node492 : node485;
														assign node485 = (inp[15]) ? node489 : node486;
															assign node486 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node489 = (inp[0]) ? 4'b1100 : 4'b1110;
														assign node492 = (inp[0]) ? node496 : node493;
															assign node493 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node496 = (inp[15]) ? 4'b1100 : 4'b1110;
												assign node499 = (inp[8]) ? node507 : node500;
													assign node500 = (inp[0]) ? node504 : node501;
														assign node501 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node504 = (inp[15]) ? 4'b1100 : 4'b1110;
													assign node507 = (inp[12]) ? node515 : node508;
														assign node508 = (inp[15]) ? node512 : node509;
															assign node509 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node512 = (inp[0]) ? 4'b1101 : 4'b1111;
														assign node515 = (inp[5]) ? node517 : 4'b1111;
															assign node517 = (inp[0]) ? node519 : 4'b1101;
																assign node519 = (inp[15]) ? 4'b1101 : 4'b1111;
								assign node522 = (inp[7]) ? node760 : node523;
									assign node523 = (inp[8]) ? node605 : node524;
										assign node524 = (inp[4]) ? node564 : node525;
											assign node525 = (inp[9]) ? node545 : node526;
												assign node526 = (inp[0]) ? node534 : node527;
													assign node527 = (inp[15]) ? 4'b1100 : node528;
														assign node528 = (inp[3]) ? node530 : 4'b1110;
															assign node530 = (inp[5]) ? 4'b1100 : 4'b1110;
													assign node534 = (inp[15]) ? node540 : node535;
														assign node535 = (inp[3]) ? node537 : 4'b1100;
															assign node537 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node540 = (inp[5]) ? node542 : 4'b1110;
															assign node542 = (inp[3]) ? 4'b1100 : 4'b1110;
												assign node545 = (inp[3]) ? node553 : node546;
													assign node546 = (inp[0]) ? node550 : node547;
														assign node547 = (inp[15]) ? 4'b1000 : 4'b1010;
														assign node550 = (inp[15]) ? 4'b1010 : 4'b1000;
													assign node553 = (inp[12]) ? node555 : 4'b1010;
														assign node555 = (inp[0]) ? 4'b1010 : node556;
															assign node556 = (inp[5]) ? node560 : node557;
																assign node557 = (inp[15]) ? 4'b1000 : 4'b1010;
																assign node560 = (inp[15]) ? 4'b1010 : 4'b1000;
											assign node564 = (inp[9]) ? node588 : node565;
												assign node565 = (inp[0]) ? node577 : node566;
													assign node566 = (inp[15]) ? node572 : node567;
														assign node567 = (inp[5]) ? node569 : 4'b1010;
															assign node569 = (inp[3]) ? 4'b1000 : 4'b1010;
														assign node572 = (inp[3]) ? node574 : 4'b1000;
															assign node574 = (inp[5]) ? 4'b1010 : 4'b1000;
													assign node577 = (inp[15]) ? node583 : node578;
														assign node578 = (inp[5]) ? node580 : 4'b1000;
															assign node580 = (inp[3]) ? 4'b1010 : 4'b1000;
														assign node583 = (inp[3]) ? node585 : 4'b1010;
															assign node585 = (inp[5]) ? 4'b1000 : 4'b1010;
												assign node588 = (inp[0]) ? node598 : node589;
													assign node589 = (inp[15]) ? node595 : node590;
														assign node590 = (inp[5]) ? 4'b1100 : node591;
															assign node591 = (inp[3]) ? 4'b1100 : 4'b1110;
														assign node595 = (inp[5]) ? 4'b1110 : 4'b1100;
													assign node598 = (inp[15]) ? node602 : node599;
														assign node599 = (inp[3]) ? 4'b1110 : 4'b1100;
														assign node602 = (inp[3]) ? 4'b1100 : 4'b1110;
										assign node605 = (inp[12]) ? node683 : node606;
											assign node606 = (inp[0]) ? node648 : node607;
												assign node607 = (inp[15]) ? node625 : node608;
													assign node608 = (inp[5]) ? node616 : node609;
														assign node609 = (inp[9]) ? node613 : node610;
															assign node610 = (inp[4]) ? 4'b1011 : 4'b1111;
															assign node613 = (inp[4]) ? 4'b1111 : 4'b1011;
														assign node616 = (inp[3]) ? 4'b1101 : node617;
															assign node617 = (inp[4]) ? node621 : node618;
																assign node618 = (inp[9]) ? 4'b1011 : 4'b1111;
																assign node621 = (inp[9]) ? 4'b1101 : 4'b1011;
													assign node625 = (inp[3]) ? node633 : node626;
														assign node626 = (inp[4]) ? node630 : node627;
															assign node627 = (inp[9]) ? 4'b1001 : 4'b1101;
															assign node630 = (inp[9]) ? 4'b1101 : 4'b1001;
														assign node633 = (inp[5]) ? node641 : node634;
															assign node634 = (inp[9]) ? node638 : node635;
																assign node635 = (inp[4]) ? 4'b1001 : 4'b1101;
																assign node638 = (inp[4]) ? 4'b1111 : 4'b1001;
															assign node641 = (inp[4]) ? node645 : node642;
																assign node642 = (inp[9]) ? 4'b1011 : 4'b1111;
																assign node645 = (inp[9]) ? 4'b1111 : 4'b1011;
												assign node648 = (inp[15]) ? node662 : node649;
													assign node649 = (inp[3]) ? node657 : node650;
														assign node650 = (inp[4]) ? node654 : node651;
															assign node651 = (inp[9]) ? 4'b1001 : 4'b1101;
															assign node654 = (inp[9]) ? 4'b1101 : 4'b1001;
														assign node657 = (inp[9]) ? node659 : 4'b1111;
															assign node659 = (inp[5]) ? 4'b1011 : 4'b1001;
													assign node662 = (inp[3]) ? node672 : node663;
														assign node663 = (inp[4]) ? node667 : node664;
															assign node664 = (inp[9]) ? 4'b1011 : 4'b1111;
															assign node667 = (inp[9]) ? node669 : 4'b1011;
																assign node669 = (inp[5]) ? 4'b1101 : 4'b1111;
														assign node672 = (inp[5]) ? node678 : node673;
															assign node673 = (inp[4]) ? node675 : 4'b1011;
																assign node675 = (inp[9]) ? 4'b1101 : 4'b1011;
															assign node678 = (inp[9]) ? 4'b1001 : node679;
																assign node679 = (inp[4]) ? 4'b1001 : 4'b1101;
											assign node683 = (inp[15]) ? node723 : node684;
												assign node684 = (inp[0]) ? node702 : node685;
													assign node685 = (inp[5]) ? node693 : node686;
														assign node686 = (inp[9]) ? node690 : node687;
															assign node687 = (inp[4]) ? 4'b1011 : 4'b1111;
															assign node690 = (inp[4]) ? 4'b1101 : 4'b1011;
														assign node693 = (inp[3]) ? node697 : node694;
															assign node694 = (inp[4]) ? 4'b1101 : 4'b1011;
															assign node697 = (inp[9]) ? 4'b1001 : node698;
																assign node698 = (inp[4]) ? 4'b1001 : 4'b1101;
													assign node702 = (inp[5]) ? node714 : node703;
														assign node703 = (inp[3]) ? node709 : node704;
															assign node704 = (inp[4]) ? node706 : 4'b1101;
																assign node706 = (inp[9]) ? 4'b1101 : 4'b1001;
															assign node709 = (inp[4]) ? 4'b1001 : node710;
																assign node710 = (inp[9]) ? 4'b1001 : 4'b1101;
														assign node714 = (inp[3]) ? node720 : node715;
															assign node715 = (inp[9]) ? node717 : 4'b1001;
																assign node717 = (inp[4]) ? 4'b1111 : 4'b1001;
															assign node720 = (inp[4]) ? 4'b1011 : 4'b1111;
												assign node723 = (inp[0]) ? node741 : node724;
													assign node724 = (inp[5]) ? node732 : node725;
														assign node725 = (inp[9]) ? node729 : node726;
															assign node726 = (inp[4]) ? 4'b1001 : 4'b1101;
															assign node729 = (inp[4]) ? 4'b1111 : 4'b1001;
														assign node732 = (inp[3]) ? 4'b1111 : node733;
															assign node733 = (inp[9]) ? node737 : node734;
																assign node734 = (inp[4]) ? 4'b1001 : 4'b1101;
																assign node737 = (inp[4]) ? 4'b1111 : 4'b1001;
													assign node741 = (inp[3]) ? node749 : node742;
														assign node742 = (inp[5]) ? node744 : 4'b1111;
															assign node744 = (inp[9]) ? 4'b1011 : node745;
																assign node745 = (inp[4]) ? 4'b1011 : 4'b1111;
														assign node749 = (inp[5]) ? node755 : node750;
															assign node750 = (inp[9]) ? node752 : 4'b1011;
																assign node752 = (inp[4]) ? 4'b1101 : 4'b1011;
															assign node755 = (inp[4]) ? node757 : 4'b1001;
																assign node757 = (inp[9]) ? 4'b1101 : 4'b1001;
									assign node760 = (inp[8]) ? node870 : node761;
										assign node761 = (inp[15]) ? node825 : node762;
											assign node762 = (inp[5]) ? node788 : node763;
												assign node763 = (inp[0]) ? node771 : node764;
													assign node764 = (inp[4]) ? node768 : node765;
														assign node765 = (inp[9]) ? 4'b1011 : 4'b1111;
														assign node768 = (inp[9]) ? 4'b1101 : 4'b1011;
													assign node771 = (inp[3]) ? node781 : node772;
														assign node772 = (inp[12]) ? node774 : 4'b1101;
															assign node774 = (inp[4]) ? node778 : node775;
																assign node775 = (inp[9]) ? 4'b1001 : 4'b1101;
																assign node778 = (inp[9]) ? 4'b1101 : 4'b1001;
														assign node781 = (inp[4]) ? node785 : node782;
															assign node782 = (inp[9]) ? 4'b1001 : 4'b1101;
															assign node785 = (inp[9]) ? 4'b1111 : 4'b1001;
												assign node788 = (inp[0]) ? node804 : node789;
													assign node789 = (inp[3]) ? node797 : node790;
														assign node790 = (inp[4]) ? node794 : node791;
															assign node791 = (inp[9]) ? 4'b1011 : 4'b1111;
															assign node794 = (inp[9]) ? 4'b1101 : 4'b1011;
														assign node797 = (inp[4]) ? node801 : node798;
															assign node798 = (inp[9]) ? 4'b1001 : 4'b1101;
															assign node801 = (inp[9]) ? 4'b1101 : 4'b1001;
													assign node804 = (inp[3]) ? node812 : node805;
														assign node805 = (inp[9]) ? node809 : node806;
															assign node806 = (inp[4]) ? 4'b1001 : 4'b1101;
															assign node809 = (inp[4]) ? 4'b1111 : 4'b1001;
														assign node812 = (inp[12]) ? node820 : node813;
															assign node813 = (inp[4]) ? node817 : node814;
																assign node814 = (inp[9]) ? 4'b1011 : 4'b1111;
																assign node817 = (inp[9]) ? 4'b1111 : 4'b1011;
															assign node820 = (inp[9]) ? 4'b1011 : node821;
																assign node821 = (inp[4]) ? 4'b1011 : 4'b1111;
											assign node825 = (inp[0]) ? node855 : node826;
												assign node826 = (inp[3]) ? node836 : node827;
													assign node827 = (inp[4]) ? node831 : node828;
														assign node828 = (inp[9]) ? 4'b1001 : 4'b1101;
														assign node831 = (inp[9]) ? node833 : 4'b1001;
															assign node833 = (inp[5]) ? 4'b1111 : 4'b1101;
													assign node836 = (inp[5]) ? node846 : node837;
														assign node837 = (inp[12]) ? node843 : node838;
															assign node838 = (inp[9]) ? node840 : 4'b1001;
																assign node840 = (inp[4]) ? 4'b1111 : 4'b1001;
															assign node843 = (inp[9]) ? 4'b1111 : 4'b1101;
														assign node846 = (inp[12]) ? node848 : 4'b1011;
															assign node848 = (inp[9]) ? node852 : node849;
																assign node849 = (inp[4]) ? 4'b1011 : 4'b1111;
																assign node852 = (inp[4]) ? 4'b1111 : 4'b1011;
												assign node855 = (inp[4]) ? node863 : node856;
													assign node856 = (inp[9]) ? 4'b1011 : node857;
														assign node857 = (inp[5]) ? node859 : 4'b1111;
															assign node859 = (inp[3]) ? 4'b1101 : 4'b1111;
													assign node863 = (inp[9]) ? 4'b1101 : node864;
														assign node864 = (inp[5]) ? node866 : 4'b1011;
															assign node866 = (inp[3]) ? 4'b1001 : 4'b1011;
										assign node870 = (inp[4]) ? node922 : node871;
											assign node871 = (inp[9]) ? node899 : node872;
												assign node872 = (inp[3]) ? node886 : node873;
													assign node873 = (inp[5]) ? node879 : node874;
														assign node874 = (inp[12]) ? node876 : 4'b1110;
															assign node876 = (inp[15]) ? 4'b1100 : 4'b1110;
														assign node879 = (inp[15]) ? node883 : node880;
															assign node880 = (inp[0]) ? 4'b1100 : 4'b1110;
															assign node883 = (inp[0]) ? 4'b1110 : 4'b1100;
													assign node886 = (inp[12]) ? node894 : node887;
														assign node887 = (inp[5]) ? node889 : 4'b1100;
															assign node889 = (inp[15]) ? 4'b1110 : node890;
																assign node890 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node894 = (inp[5]) ? 4'b1100 : node895;
															assign node895 = (inp[15]) ? 4'b1100 : 4'b1110;
												assign node899 = (inp[15]) ? node911 : node900;
													assign node900 = (inp[0]) ? node906 : node901;
														assign node901 = (inp[3]) ? node903 : 4'b1010;
															assign node903 = (inp[5]) ? 4'b1000 : 4'b1010;
														assign node906 = (inp[3]) ? node908 : 4'b1000;
															assign node908 = (inp[5]) ? 4'b1010 : 4'b1000;
													assign node911 = (inp[0]) ? node917 : node912;
														assign node912 = (inp[3]) ? node914 : 4'b1000;
															assign node914 = (inp[5]) ? 4'b1010 : 4'b1000;
														assign node917 = (inp[5]) ? node919 : 4'b1010;
															assign node919 = (inp[3]) ? 4'b1000 : 4'b1010;
											assign node922 = (inp[9]) ? node954 : node923;
												assign node923 = (inp[5]) ? node939 : node924;
													assign node924 = (inp[12]) ? node932 : node925;
														assign node925 = (inp[0]) ? node929 : node926;
															assign node926 = (inp[15]) ? 4'b1000 : 4'b1010;
															assign node929 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node932 = (inp[0]) ? node936 : node933;
															assign node933 = (inp[15]) ? 4'b1000 : 4'b1010;
															assign node936 = (inp[15]) ? 4'b1010 : 4'b1000;
													assign node939 = (inp[0]) ? node949 : node940;
														assign node940 = (inp[12]) ? node946 : node941;
															assign node941 = (inp[15]) ? node943 : 4'b1010;
																assign node943 = (inp[3]) ? 4'b1010 : 4'b1000;
															assign node946 = (inp[3]) ? 4'b1000 : 4'b1010;
														assign node949 = (inp[15]) ? 4'b1000 : node950;
															assign node950 = (inp[3]) ? 4'b1010 : 4'b1000;
												assign node954 = (inp[0]) ? node964 : node955;
													assign node955 = (inp[15]) ? node959 : node956;
														assign node956 = (inp[3]) ? 4'b1100 : 4'b1110;
														assign node959 = (inp[5]) ? 4'b1110 : node960;
															assign node960 = (inp[12]) ? 4'b1110 : 4'b1100;
													assign node964 = (inp[15]) ? node970 : node965;
														assign node965 = (inp[3]) ? 4'b1110 : node966;
															assign node966 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node970 = (inp[3]) ? 4'b1100 : node971;
															assign node971 = (inp[5]) ? 4'b1100 : 4'b1110;
							assign node975 = (inp[3]) ? node1417 : node976;
								assign node976 = (inp[4]) ? node1186 : node977;
									assign node977 = (inp[9]) ? node1059 : node978;
										assign node978 = (inp[15]) ? node1002 : node979;
											assign node979 = (inp[0]) ? node987 : node980;
												assign node980 = (inp[8]) ? node984 : node981;
													assign node981 = (inp[7]) ? 4'b1111 : 4'b1110;
													assign node984 = (inp[7]) ? 4'b1110 : 4'b1111;
												assign node987 = (inp[14]) ? node995 : node988;
													assign node988 = (inp[8]) ? node992 : node989;
														assign node989 = (inp[7]) ? 4'b1101 : 4'b1100;
														assign node992 = (inp[7]) ? 4'b1100 : 4'b1101;
													assign node995 = (inp[7]) ? node999 : node996;
														assign node996 = (inp[8]) ? 4'b1101 : 4'b1100;
														assign node999 = (inp[8]) ? 4'b1100 : 4'b1101;
											assign node1002 = (inp[0]) ? node1036 : node1003;
												assign node1003 = (inp[5]) ? node1019 : node1004;
													assign node1004 = (inp[14]) ? node1012 : node1005;
														assign node1005 = (inp[7]) ? node1009 : node1006;
															assign node1006 = (inp[8]) ? 4'b1101 : 4'b1100;
															assign node1009 = (inp[8]) ? 4'b1100 : 4'b1101;
														assign node1012 = (inp[7]) ? node1016 : node1013;
															assign node1013 = (inp[8]) ? 4'b1101 : 4'b1100;
															assign node1016 = (inp[8]) ? 4'b1100 : 4'b1101;
													assign node1019 = (inp[14]) ? node1027 : node1020;
														assign node1020 = (inp[12]) ? 4'b1100 : node1021;
															assign node1021 = (inp[7]) ? node1023 : 4'b1100;
																assign node1023 = (inp[8]) ? 4'b1100 : 4'b1101;
														assign node1027 = (inp[12]) ? 4'b1101 : node1028;
															assign node1028 = (inp[7]) ? node1032 : node1029;
																assign node1029 = (inp[8]) ? 4'b1101 : 4'b1100;
																assign node1032 = (inp[8]) ? 4'b1100 : 4'b1101;
												assign node1036 = (inp[12]) ? node1052 : node1037;
													assign node1037 = (inp[14]) ? node1039 : 4'b1111;
														assign node1039 = (inp[5]) ? node1045 : node1040;
															assign node1040 = (inp[7]) ? node1042 : 4'b1110;
																assign node1042 = (inp[8]) ? 4'b1110 : 4'b1111;
															assign node1045 = (inp[8]) ? node1049 : node1046;
																assign node1046 = (inp[7]) ? 4'b1111 : 4'b1110;
																assign node1049 = (inp[7]) ? 4'b1110 : 4'b1111;
													assign node1052 = (inp[14]) ? node1054 : 4'b1110;
														assign node1054 = (inp[8]) ? node1056 : 4'b1111;
															assign node1056 = (inp[7]) ? 4'b1110 : 4'b1111;
										assign node1059 = (inp[5]) ? node1121 : node1060;
											assign node1060 = (inp[15]) ? node1084 : node1061;
												assign node1061 = (inp[0]) ? node1069 : node1062;
													assign node1062 = (inp[7]) ? node1066 : node1063;
														assign node1063 = (inp[8]) ? 4'b1011 : 4'b1010;
														assign node1066 = (inp[8]) ? 4'b1010 : 4'b1011;
													assign node1069 = (inp[14]) ? node1077 : node1070;
														assign node1070 = (inp[7]) ? node1074 : node1071;
															assign node1071 = (inp[8]) ? 4'b1001 : 4'b1000;
															assign node1074 = (inp[8]) ? 4'b1000 : 4'b1001;
														assign node1077 = (inp[8]) ? node1081 : node1078;
															assign node1078 = (inp[7]) ? 4'b1001 : 4'b1000;
															assign node1081 = (inp[7]) ? 4'b1000 : 4'b1001;
												assign node1084 = (inp[0]) ? node1102 : node1085;
													assign node1085 = (inp[12]) ? node1091 : node1086;
														assign node1086 = (inp[8]) ? node1088 : 4'b1001;
															assign node1088 = (inp[7]) ? 4'b1000 : 4'b1001;
														assign node1091 = (inp[14]) ? node1097 : node1092;
															assign node1092 = (inp[7]) ? 4'b1000 : node1093;
																assign node1093 = (inp[8]) ? 4'b1001 : 4'b1000;
															assign node1097 = (inp[8]) ? 4'b1001 : node1098;
																assign node1098 = (inp[7]) ? 4'b1001 : 4'b1000;
													assign node1102 = (inp[12]) ? node1114 : node1103;
														assign node1103 = (inp[14]) ? node1109 : node1104;
															assign node1104 = (inp[8]) ? 4'b1011 : node1105;
																assign node1105 = (inp[7]) ? 4'b1011 : 4'b1010;
															assign node1109 = (inp[7]) ? node1111 : 4'b1010;
																assign node1111 = (inp[8]) ? 4'b1010 : 4'b1011;
														assign node1114 = (inp[14]) ? 4'b1011 : node1115;
															assign node1115 = (inp[7]) ? node1117 : 4'b1011;
																assign node1117 = (inp[8]) ? 4'b1010 : 4'b1011;
											assign node1121 = (inp[14]) ? node1153 : node1122;
												assign node1122 = (inp[15]) ? node1144 : node1123;
													assign node1123 = (inp[0]) ? node1131 : node1124;
														assign node1124 = (inp[12]) ? 4'b1011 : node1125;
															assign node1125 = (inp[7]) ? node1127 : 4'b1011;
																assign node1127 = (inp[8]) ? 4'b1010 : 4'b1011;
														assign node1131 = (inp[12]) ? node1137 : node1132;
															assign node1132 = (inp[7]) ? 4'b1001 : node1133;
																assign node1133 = (inp[8]) ? 4'b1001 : 4'b1000;
															assign node1137 = (inp[7]) ? node1141 : node1138;
																assign node1138 = (inp[8]) ? 4'b1001 : 4'b1000;
																assign node1141 = (inp[8]) ? 4'b1000 : 4'b1001;
													assign node1144 = (inp[0]) ? 4'b1010 : node1145;
														assign node1145 = (inp[8]) ? node1149 : node1146;
															assign node1146 = (inp[7]) ? 4'b1001 : 4'b1000;
															assign node1149 = (inp[7]) ? 4'b1000 : 4'b1001;
												assign node1153 = (inp[0]) ? node1171 : node1154;
													assign node1154 = (inp[15]) ? node1166 : node1155;
														assign node1155 = (inp[12]) ? node1161 : node1156;
															assign node1156 = (inp[8]) ? 4'b1010 : node1157;
																assign node1157 = (inp[7]) ? 4'b1011 : 4'b1010;
															assign node1161 = (inp[7]) ? node1163 : 4'b1011;
																assign node1163 = (inp[8]) ? 4'b1010 : 4'b1011;
														assign node1166 = (inp[12]) ? 4'b1000 : node1167;
															assign node1167 = (inp[7]) ? 4'b1001 : 4'b1000;
													assign node1171 = (inp[15]) ? node1179 : node1172;
														assign node1172 = (inp[8]) ? node1176 : node1173;
															assign node1173 = (inp[7]) ? 4'b1001 : 4'b1000;
															assign node1176 = (inp[7]) ? 4'b1000 : 4'b1001;
														assign node1179 = (inp[8]) ? node1183 : node1180;
															assign node1180 = (inp[7]) ? 4'b1011 : 4'b1010;
															assign node1183 = (inp[7]) ? 4'b1010 : 4'b1011;
									assign node1186 = (inp[9]) ? node1314 : node1187;
										assign node1187 = (inp[12]) ? node1261 : node1188;
											assign node1188 = (inp[14]) ? node1230 : node1189;
												assign node1189 = (inp[5]) ? node1217 : node1190;
													assign node1190 = (inp[7]) ? node1204 : node1191;
														assign node1191 = (inp[8]) ? node1199 : node1192;
															assign node1192 = (inp[15]) ? node1196 : node1193;
																assign node1193 = (inp[0]) ? 4'b1000 : 4'b1010;
																assign node1196 = (inp[0]) ? 4'b1010 : 4'b1000;
															assign node1199 = (inp[0]) ? 4'b1011 : node1200;
																assign node1200 = (inp[15]) ? 4'b1001 : 4'b1011;
														assign node1204 = (inp[8]) ? node1210 : node1205;
															assign node1205 = (inp[15]) ? 4'b1011 : node1206;
																assign node1206 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node1210 = (inp[0]) ? node1214 : node1211;
																assign node1211 = (inp[15]) ? 4'b1000 : 4'b1010;
																assign node1214 = (inp[15]) ? 4'b1010 : 4'b1000;
													assign node1217 = (inp[8]) ? node1223 : node1218;
														assign node1218 = (inp[15]) ? node1220 : 4'b1010;
															assign node1220 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node1223 = (inp[7]) ? node1225 : 4'b1001;
															assign node1225 = (inp[15]) ? 4'b1000 : node1226;
																assign node1226 = (inp[0]) ? 4'b1000 : 4'b1010;
												assign node1230 = (inp[15]) ? node1248 : node1231;
													assign node1231 = (inp[0]) ? node1241 : node1232;
														assign node1232 = (inp[5]) ? node1234 : 4'b1011;
															assign node1234 = (inp[7]) ? node1238 : node1235;
																assign node1235 = (inp[8]) ? 4'b1011 : 4'b1010;
																assign node1238 = (inp[8]) ? 4'b1010 : 4'b1011;
														assign node1241 = (inp[8]) ? node1245 : node1242;
															assign node1242 = (inp[7]) ? 4'b1001 : 4'b1000;
															assign node1245 = (inp[7]) ? 4'b1000 : 4'b1001;
													assign node1248 = (inp[0]) ? node1256 : node1249;
														assign node1249 = (inp[7]) ? node1253 : node1250;
															assign node1250 = (inp[8]) ? 4'b1001 : 4'b1000;
															assign node1253 = (inp[8]) ? 4'b1000 : 4'b1001;
														assign node1256 = (inp[5]) ? node1258 : 4'b1010;
															assign node1258 = (inp[7]) ? 4'b1010 : 4'b1011;
											assign node1261 = (inp[5]) ? node1285 : node1262;
												assign node1262 = (inp[8]) ? node1276 : node1263;
													assign node1263 = (inp[7]) ? node1271 : node1264;
														assign node1264 = (inp[15]) ? node1268 : node1265;
															assign node1265 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node1268 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node1271 = (inp[0]) ? node1273 : 4'b1011;
															assign node1273 = (inp[15]) ? 4'b1011 : 4'b1001;
													assign node1276 = (inp[7]) ? node1278 : 4'b1001;
														assign node1278 = (inp[15]) ? node1282 : node1279;
															assign node1279 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node1282 = (inp[0]) ? 4'b1010 : 4'b1000;
												assign node1285 = (inp[14]) ? node1305 : node1286;
													assign node1286 = (inp[8]) ? node1296 : node1287;
														assign node1287 = (inp[7]) ? node1289 : 4'b1010;
															assign node1289 = (inp[0]) ? node1293 : node1290;
																assign node1290 = (inp[15]) ? 4'b1001 : 4'b1011;
																assign node1293 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node1296 = (inp[7]) ? node1298 : 4'b1011;
															assign node1298 = (inp[15]) ? node1302 : node1299;
																assign node1299 = (inp[0]) ? 4'b1000 : 4'b1010;
																assign node1302 = (inp[0]) ? 4'b1010 : 4'b1000;
													assign node1305 = (inp[15]) ? 4'b1011 : node1306;
														assign node1306 = (inp[0]) ? node1308 : 4'b1011;
															assign node1308 = (inp[8]) ? 4'b1001 : node1309;
																assign node1309 = (inp[7]) ? 4'b1001 : 4'b1000;
										assign node1314 = (inp[0]) ? node1368 : node1315;
											assign node1315 = (inp[14]) ? node1345 : node1316;
												assign node1316 = (inp[8]) ? node1330 : node1317;
													assign node1317 = (inp[7]) ? node1327 : node1318;
														assign node1318 = (inp[12]) ? node1324 : node1319;
															assign node1319 = (inp[5]) ? node1321 : 4'b1100;
																assign node1321 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node1324 = (inp[5]) ? 4'b1100 : 4'b1110;
														assign node1327 = (inp[12]) ? 4'b1111 : 4'b1101;
													assign node1330 = (inp[7]) ? node1338 : node1331;
														assign node1331 = (inp[15]) ? node1335 : node1332;
															assign node1332 = (inp[5]) ? 4'b1101 : 4'b1111;
															assign node1335 = (inp[5]) ? 4'b1111 : 4'b1101;
														assign node1338 = (inp[5]) ? node1342 : node1339;
															assign node1339 = (inp[15]) ? 4'b1100 : 4'b1110;
															assign node1342 = (inp[15]) ? 4'b1110 : 4'b1100;
												assign node1345 = (inp[8]) ? node1361 : node1346;
													assign node1346 = (inp[7]) ? node1354 : node1347;
														assign node1347 = (inp[15]) ? node1351 : node1348;
															assign node1348 = (inp[5]) ? 4'b1100 : 4'b1110;
															assign node1351 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node1354 = (inp[5]) ? node1358 : node1355;
															assign node1355 = (inp[15]) ? 4'b1101 : 4'b1111;
															assign node1358 = (inp[15]) ? 4'b1111 : 4'b1101;
													assign node1361 = (inp[7]) ? node1363 : 4'b1101;
														assign node1363 = (inp[15]) ? node1365 : 4'b1100;
															assign node1365 = (inp[5]) ? 4'b1110 : 4'b1100;
											assign node1368 = (inp[8]) ? node1392 : node1369;
												assign node1369 = (inp[7]) ? node1385 : node1370;
													assign node1370 = (inp[12]) ? node1378 : node1371;
														assign node1371 = (inp[14]) ? node1373 : 4'b1110;
															assign node1373 = (inp[5]) ? node1375 : 4'b1110;
																assign node1375 = (inp[15]) ? 4'b1100 : 4'b1110;
														assign node1378 = (inp[15]) ? node1382 : node1379;
															assign node1379 = (inp[5]) ? 4'b1110 : 4'b1100;
															assign node1382 = (inp[5]) ? 4'b1100 : 4'b1110;
													assign node1385 = (inp[15]) ? node1389 : node1386;
														assign node1386 = (inp[5]) ? 4'b1111 : 4'b1101;
														assign node1389 = (inp[5]) ? 4'b1101 : 4'b1111;
												assign node1392 = (inp[7]) ? node1402 : node1393;
													assign node1393 = (inp[12]) ? node1395 : 4'b1101;
														assign node1395 = (inp[5]) ? node1399 : node1396;
															assign node1396 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node1399 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node1402 = (inp[12]) ? node1410 : node1403;
														assign node1403 = (inp[5]) ? node1407 : node1404;
															assign node1404 = (inp[14]) ? 4'b1100 : 4'b1110;
															assign node1407 = (inp[15]) ? 4'b1100 : 4'b1110;
														assign node1410 = (inp[5]) ? node1414 : node1411;
															assign node1411 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node1414 = (inp[15]) ? 4'b1100 : 4'b1110;
								assign node1417 = (inp[9]) ? node1715 : node1418;
									assign node1418 = (inp[4]) ? node1586 : node1419;
										assign node1419 = (inp[12]) ? node1511 : node1420;
											assign node1420 = (inp[14]) ? node1472 : node1421;
												assign node1421 = (inp[0]) ? node1445 : node1422;
													assign node1422 = (inp[7]) ? node1436 : node1423;
														assign node1423 = (inp[8]) ? node1431 : node1424;
															assign node1424 = (inp[15]) ? node1428 : node1425;
																assign node1425 = (inp[5]) ? 4'b1100 : 4'b1110;
																assign node1428 = (inp[5]) ? 4'b1110 : 4'b1100;
															assign node1431 = (inp[15]) ? 4'b1101 : node1432;
																assign node1432 = (inp[5]) ? 4'b1101 : 4'b1111;
														assign node1436 = (inp[8]) ? node1438 : 4'b1101;
															assign node1438 = (inp[15]) ? node1442 : node1439;
																assign node1439 = (inp[5]) ? 4'b1100 : 4'b1110;
																assign node1442 = (inp[5]) ? 4'b1110 : 4'b1100;
													assign node1445 = (inp[7]) ? node1459 : node1446;
														assign node1446 = (inp[8]) ? node1452 : node1447;
															assign node1447 = (inp[15]) ? 4'b1100 : node1448;
																assign node1448 = (inp[5]) ? 4'b1110 : 4'b1100;
															assign node1452 = (inp[5]) ? node1456 : node1453;
																assign node1453 = (inp[15]) ? 4'b1111 : 4'b1101;
																assign node1456 = (inp[15]) ? 4'b1101 : 4'b1111;
														assign node1459 = (inp[8]) ? node1465 : node1460;
															assign node1460 = (inp[15]) ? node1462 : 4'b1111;
																assign node1462 = (inp[5]) ? 4'b1101 : 4'b1111;
															assign node1465 = (inp[15]) ? node1469 : node1466;
																assign node1466 = (inp[5]) ? 4'b1110 : 4'b1100;
																assign node1469 = (inp[5]) ? 4'b1100 : 4'b1110;
												assign node1472 = (inp[5]) ? node1492 : node1473;
													assign node1473 = (inp[7]) ? node1485 : node1474;
														assign node1474 = (inp[8]) ? node1478 : node1475;
															assign node1475 = (inp[15]) ? 4'b1100 : 4'b1110;
															assign node1478 = (inp[15]) ? node1482 : node1479;
																assign node1479 = (inp[0]) ? 4'b1101 : 4'b1111;
																assign node1482 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node1485 = (inp[8]) ? 4'b1100 : node1486;
															assign node1486 = (inp[15]) ? node1488 : 4'b1101;
																assign node1488 = (inp[0]) ? 4'b1111 : 4'b1101;
													assign node1492 = (inp[8]) ? node1502 : node1493;
														assign node1493 = (inp[7]) ? node1499 : node1494;
															assign node1494 = (inp[15]) ? node1496 : 4'b1100;
																assign node1496 = (inp[0]) ? 4'b1100 : 4'b1110;
															assign node1499 = (inp[0]) ? 4'b1101 : 4'b1111;
														assign node1502 = (inp[7]) ? node1508 : node1503;
															assign node1503 = (inp[0]) ? node1505 : 4'b1101;
																assign node1505 = (inp[15]) ? 4'b1101 : 4'b1111;
															assign node1508 = (inp[15]) ? 4'b1100 : 4'b1110;
											assign node1511 = (inp[5]) ? node1555 : node1512;
												assign node1512 = (inp[7]) ? node1526 : node1513;
													assign node1513 = (inp[8]) ? node1521 : node1514;
														assign node1514 = (inp[0]) ? node1518 : node1515;
															assign node1515 = (inp[15]) ? 4'b1100 : 4'b1110;
															assign node1518 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node1521 = (inp[14]) ? 4'b1101 : node1522;
															assign node1522 = (inp[15]) ? 4'b1111 : 4'b1101;
													assign node1526 = (inp[8]) ? node1542 : node1527;
														assign node1527 = (inp[14]) ? node1535 : node1528;
															assign node1528 = (inp[0]) ? node1532 : node1529;
																assign node1529 = (inp[15]) ? 4'b1101 : 4'b1111;
																assign node1532 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node1535 = (inp[0]) ? node1539 : node1536;
																assign node1536 = (inp[15]) ? 4'b1101 : 4'b1111;
																assign node1539 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node1542 = (inp[14]) ? node1550 : node1543;
															assign node1543 = (inp[15]) ? node1547 : node1544;
																assign node1544 = (inp[0]) ? 4'b1100 : 4'b1110;
																assign node1547 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node1550 = (inp[15]) ? node1552 : 4'b1100;
																assign node1552 = (inp[0]) ? 4'b1110 : 4'b1100;
												assign node1555 = (inp[14]) ? node1575 : node1556;
													assign node1556 = (inp[0]) ? node1566 : node1557;
														assign node1557 = (inp[15]) ? node1561 : node1558;
															assign node1558 = (inp[7]) ? 4'b1101 : 4'b1100;
															assign node1561 = (inp[8]) ? node1563 : 4'b1111;
																assign node1563 = (inp[7]) ? 4'b1110 : 4'b1111;
														assign node1566 = (inp[15]) ? node1568 : 4'b1111;
															assign node1568 = (inp[8]) ? node1572 : node1569;
																assign node1569 = (inp[7]) ? 4'b1101 : 4'b1100;
																assign node1572 = (inp[7]) ? 4'b1100 : 4'b1101;
													assign node1575 = (inp[7]) ? node1579 : node1576;
														assign node1576 = (inp[8]) ? 4'b1111 : 4'b1110;
														assign node1579 = (inp[8]) ? node1581 : 4'b1111;
															assign node1581 = (inp[0]) ? node1583 : 4'b1100;
																assign node1583 = (inp[15]) ? 4'b1100 : 4'b1110;
										assign node1586 = (inp[14]) ? node1658 : node1587;
											assign node1587 = (inp[8]) ? node1625 : node1588;
												assign node1588 = (inp[7]) ? node1604 : node1589;
													assign node1589 = (inp[5]) ? 4'b1000 : node1590;
														assign node1590 = (inp[12]) ? node1596 : node1591;
															assign node1591 = (inp[15]) ? node1593 : 4'b1000;
																assign node1593 = (inp[0]) ? 4'b1010 : 4'b1000;
															assign node1596 = (inp[15]) ? node1600 : node1597;
																assign node1597 = (inp[0]) ? 4'b1000 : 4'b1010;
																assign node1600 = (inp[0]) ? 4'b1010 : 4'b1000;
													assign node1604 = (inp[12]) ? node1618 : node1605;
														assign node1605 = (inp[15]) ? node1613 : node1606;
															assign node1606 = (inp[5]) ? node1610 : node1607;
																assign node1607 = (inp[0]) ? 4'b1001 : 4'b1011;
																assign node1610 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node1613 = (inp[5]) ? 4'b1001 : node1614;
																assign node1614 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node1618 = (inp[5]) ? 4'b1001 : node1619;
															assign node1619 = (inp[15]) ? 4'b1001 : node1620;
																assign node1620 = (inp[0]) ? 4'b1001 : 4'b1011;
												assign node1625 = (inp[7]) ? node1643 : node1626;
													assign node1626 = (inp[15]) ? node1634 : node1627;
														assign node1627 = (inp[5]) ? node1631 : node1628;
															assign node1628 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node1631 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node1634 = (inp[12]) ? node1636 : 4'b1011;
															assign node1636 = (inp[0]) ? node1640 : node1637;
																assign node1637 = (inp[5]) ? 4'b1011 : 4'b1001;
																assign node1640 = (inp[5]) ? 4'b1001 : 4'b1011;
													assign node1643 = (inp[15]) ? node1649 : node1644;
														assign node1644 = (inp[5]) ? node1646 : 4'b1010;
															assign node1646 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node1649 = (inp[12]) ? 4'b1000 : node1650;
															assign node1650 = (inp[5]) ? node1654 : node1651;
																assign node1651 = (inp[0]) ? 4'b1010 : 4'b1000;
																assign node1654 = (inp[0]) ? 4'b1000 : 4'b1010;
											assign node1658 = (inp[0]) ? node1686 : node1659;
												assign node1659 = (inp[7]) ? node1667 : node1660;
													assign node1660 = (inp[8]) ? 4'b1011 : node1661;
														assign node1661 = (inp[15]) ? node1663 : 4'b1010;
															assign node1663 = (inp[5]) ? 4'b1010 : 4'b1000;
													assign node1667 = (inp[8]) ? node1677 : node1668;
														assign node1668 = (inp[12]) ? node1670 : 4'b1001;
															assign node1670 = (inp[5]) ? node1674 : node1671;
																assign node1671 = (inp[15]) ? 4'b1001 : 4'b1011;
																assign node1674 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node1677 = (inp[12]) ? node1679 : 4'b1000;
															assign node1679 = (inp[15]) ? node1683 : node1680;
																assign node1680 = (inp[5]) ? 4'b1000 : 4'b1010;
																assign node1683 = (inp[5]) ? 4'b1010 : 4'b1000;
												assign node1686 = (inp[7]) ? node1700 : node1687;
													assign node1687 = (inp[8]) ? node1693 : node1688;
														assign node1688 = (inp[5]) ? node1690 : 4'b1000;
															assign node1690 = (inp[15]) ? 4'b1000 : 4'b1010;
														assign node1693 = (inp[5]) ? node1697 : node1694;
															assign node1694 = (inp[15]) ? 4'b1011 : 4'b1001;
															assign node1697 = (inp[15]) ? 4'b1001 : 4'b1011;
													assign node1700 = (inp[8]) ? node1706 : node1701;
														assign node1701 = (inp[5]) ? 4'b1011 : node1702;
															assign node1702 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node1706 = (inp[12]) ? 4'b1000 : node1707;
															assign node1707 = (inp[5]) ? node1711 : node1708;
																assign node1708 = (inp[15]) ? 4'b1010 : 4'b1000;
																assign node1711 = (inp[15]) ? 4'b1000 : 4'b1010;
									assign node1715 = (inp[4]) ? node1843 : node1716;
										assign node1716 = (inp[12]) ? node1790 : node1717;
											assign node1717 = (inp[14]) ? node1755 : node1718;
												assign node1718 = (inp[5]) ? node1740 : node1719;
													assign node1719 = (inp[7]) ? node1727 : node1720;
														assign node1720 = (inp[8]) ? 4'b1011 : node1721;
															assign node1721 = (inp[0]) ? node1723 : 4'b1010;
																assign node1723 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node1727 = (inp[8]) ? node1733 : node1728;
															assign node1728 = (inp[15]) ? node1730 : 4'b1001;
																assign node1730 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node1733 = (inp[15]) ? node1737 : node1734;
																assign node1734 = (inp[0]) ? 4'b1000 : 4'b1010;
																assign node1737 = (inp[0]) ? 4'b1010 : 4'b1000;
													assign node1740 = (inp[8]) ? node1746 : node1741;
														assign node1741 = (inp[15]) ? node1743 : 4'b1000;
															assign node1743 = (inp[0]) ? 4'b1000 : 4'b1010;
														assign node1746 = (inp[7]) ? node1748 : 4'b1011;
															assign node1748 = (inp[15]) ? node1752 : node1749;
																assign node1749 = (inp[0]) ? 4'b1010 : 4'b1000;
																assign node1752 = (inp[0]) ? 4'b1000 : 4'b1010;
												assign node1755 = (inp[15]) ? node1769 : node1756;
													assign node1756 = (inp[0]) ? node1762 : node1757;
														assign node1757 = (inp[5]) ? 4'b1001 : node1758;
															assign node1758 = (inp[7]) ? 4'b1011 : 4'b1010;
														assign node1762 = (inp[5]) ? node1764 : 4'b1000;
															assign node1764 = (inp[8]) ? node1766 : 4'b1010;
																assign node1766 = (inp[7]) ? 4'b1010 : 4'b1011;
													assign node1769 = (inp[7]) ? node1779 : node1770;
														assign node1770 = (inp[8]) ? node1772 : 4'b1010;
															assign node1772 = (inp[5]) ? node1776 : node1773;
																assign node1773 = (inp[0]) ? 4'b1011 : 4'b1001;
																assign node1776 = (inp[0]) ? 4'b1001 : 4'b1011;
														assign node1779 = (inp[8]) ? node1785 : node1780;
															assign node1780 = (inp[0]) ? node1782 : 4'b1011;
																assign node1782 = (inp[5]) ? 4'b1001 : 4'b1011;
															assign node1785 = (inp[5]) ? 4'b1010 : node1786;
																assign node1786 = (inp[0]) ? 4'b1010 : 4'b1000;
											assign node1790 = (inp[0]) ? node1810 : node1791;
												assign node1791 = (inp[8]) ? node1797 : node1792;
													assign node1792 = (inp[7]) ? 4'b1001 : node1793;
														assign node1793 = (inp[5]) ? 4'b1010 : 4'b1000;
													assign node1797 = (inp[7]) ? node1805 : node1798;
														assign node1798 = (inp[5]) ? node1802 : node1799;
															assign node1799 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node1802 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node1805 = (inp[5]) ? node1807 : 4'b1010;
															assign node1807 = (inp[15]) ? 4'b1010 : 4'b1000;
												assign node1810 = (inp[15]) ? node1828 : node1811;
													assign node1811 = (inp[5]) ? node1819 : node1812;
														assign node1812 = (inp[8]) ? node1816 : node1813;
															assign node1813 = (inp[7]) ? 4'b1001 : 4'b1000;
															assign node1816 = (inp[7]) ? 4'b1000 : 4'b1001;
														assign node1819 = (inp[14]) ? node1823 : node1820;
															assign node1820 = (inp[8]) ? 4'b1010 : 4'b1011;
															assign node1823 = (inp[7]) ? 4'b1011 : node1824;
																assign node1824 = (inp[8]) ? 4'b1011 : 4'b1010;
													assign node1828 = (inp[5]) ? node1836 : node1829;
														assign node1829 = (inp[8]) ? node1833 : node1830;
															assign node1830 = (inp[7]) ? 4'b1011 : 4'b1010;
															assign node1833 = (inp[7]) ? 4'b1010 : 4'b1011;
														assign node1836 = (inp[8]) ? node1840 : node1837;
															assign node1837 = (inp[7]) ? 4'b1001 : 4'b1000;
															assign node1840 = (inp[7]) ? 4'b1000 : 4'b1001;
										assign node1843 = (inp[5]) ? node1905 : node1844;
											assign node1844 = (inp[12]) ? node1878 : node1845;
												assign node1845 = (inp[8]) ? node1857 : node1846;
													assign node1846 = (inp[7]) ? node1852 : node1847;
														assign node1847 = (inp[15]) ? node1849 : 4'b1110;
															assign node1849 = (inp[0]) ? 4'b1100 : 4'b1110;
														assign node1852 = (inp[0]) ? 4'b1111 : node1853;
															assign node1853 = (inp[15]) ? 4'b1111 : 4'b1101;
													assign node1857 = (inp[7]) ? node1873 : node1858;
														assign node1858 = (inp[14]) ? node1866 : node1859;
															assign node1859 = (inp[0]) ? node1863 : node1860;
																assign node1860 = (inp[15]) ? 4'b1111 : 4'b1101;
																assign node1863 = (inp[15]) ? 4'b1101 : 4'b1111;
															assign node1866 = (inp[0]) ? node1870 : node1867;
																assign node1867 = (inp[15]) ? 4'b1111 : 4'b1101;
																assign node1870 = (inp[15]) ? 4'b1101 : 4'b1111;
														assign node1873 = (inp[0]) ? node1875 : 4'b1110;
															assign node1875 = (inp[14]) ? 4'b1110 : 4'b1100;
												assign node1878 = (inp[0]) ? node1892 : node1879;
													assign node1879 = (inp[15]) ? node1885 : node1880;
														assign node1880 = (inp[8]) ? 4'b1100 : node1881;
															assign node1881 = (inp[7]) ? 4'b1101 : 4'b1100;
														assign node1885 = (inp[7]) ? node1889 : node1886;
															assign node1886 = (inp[8]) ? 4'b1111 : 4'b1110;
															assign node1889 = (inp[8]) ? 4'b1110 : 4'b1111;
													assign node1892 = (inp[15]) ? node1900 : node1893;
														assign node1893 = (inp[8]) ? node1897 : node1894;
															assign node1894 = (inp[7]) ? 4'b1111 : 4'b1110;
															assign node1897 = (inp[7]) ? 4'b1110 : 4'b1111;
														assign node1900 = (inp[8]) ? 4'b1101 : node1901;
															assign node1901 = (inp[7]) ? 4'b1101 : 4'b1100;
											assign node1905 = (inp[14]) ? node1925 : node1906;
												assign node1906 = (inp[15]) ? node1918 : node1907;
													assign node1907 = (inp[0]) ? node1913 : node1908;
														assign node1908 = (inp[7]) ? node1910 : 4'b1101;
															assign node1910 = (inp[8]) ? 4'b1100 : 4'b1101;
														assign node1913 = (inp[7]) ? node1915 : 4'b1111;
															assign node1915 = (inp[8]) ? 4'b1110 : 4'b1111;
													assign node1918 = (inp[0]) ? 4'b1101 : node1919;
														assign node1919 = (inp[8]) ? 4'b1111 : node1920;
															assign node1920 = (inp[7]) ? 4'b1111 : 4'b1110;
												assign node1925 = (inp[15]) ? node1939 : node1926;
													assign node1926 = (inp[0]) ? node1932 : node1927;
														assign node1927 = (inp[7]) ? 4'b1101 : node1928;
															assign node1928 = (inp[8]) ? 4'b1101 : 4'b1100;
														assign node1932 = (inp[8]) ? node1936 : node1933;
															assign node1933 = (inp[7]) ? 4'b1111 : 4'b1110;
															assign node1936 = (inp[7]) ? 4'b1110 : 4'b1111;
													assign node1939 = (inp[0]) ? node1943 : node1940;
														assign node1940 = (inp[12]) ? 4'b1111 : 4'b1110;
														assign node1943 = (inp[8]) ? node1945 : 4'b1101;
															assign node1945 = (inp[7]) ? 4'b1100 : 4'b1101;
						assign node1948 = (inp[7]) ? node2740 : node1949;
							assign node1949 = (inp[8]) ? node2335 : node1950;
								assign node1950 = (inp[14]) ? node2212 : node1951;
									assign node1951 = (inp[2]) ? node2079 : node1952;
										assign node1952 = (inp[4]) ? node2010 : node1953;
											assign node1953 = (inp[9]) ? node1975 : node1954;
												assign node1954 = (inp[0]) ? node1966 : node1955;
													assign node1955 = (inp[15]) ? node1961 : node1956;
														assign node1956 = (inp[3]) ? node1958 : 4'b1111;
															assign node1958 = (inp[5]) ? 4'b1101 : 4'b1111;
														assign node1961 = (inp[3]) ? node1963 : 4'b1101;
															assign node1963 = (inp[5]) ? 4'b1111 : 4'b1101;
													assign node1966 = (inp[15]) ? node1968 : 4'b1101;
														assign node1968 = (inp[12]) ? node1970 : 4'b1101;
															assign node1970 = (inp[5]) ? node1972 : 4'b1111;
																assign node1972 = (inp[3]) ? 4'b1101 : 4'b1111;
												assign node1975 = (inp[5]) ? node1989 : node1976;
													assign node1976 = (inp[12]) ? node1984 : node1977;
														assign node1977 = (inp[0]) ? node1981 : node1978;
															assign node1978 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node1981 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node1984 = (inp[0]) ? node1986 : 4'b1011;
															assign node1986 = (inp[15]) ? 4'b1011 : 4'b1001;
													assign node1989 = (inp[0]) ? node1997 : node1990;
														assign node1990 = (inp[12]) ? node1992 : 4'b1001;
															assign node1992 = (inp[15]) ? node1994 : 4'b1001;
																assign node1994 = (inp[3]) ? 4'b1011 : 4'b1001;
														assign node1997 = (inp[12]) ? node2005 : node1998;
															assign node1998 = (inp[15]) ? node2002 : node1999;
																assign node1999 = (inp[3]) ? 4'b1011 : 4'b1001;
																assign node2002 = (inp[3]) ? 4'b1001 : 4'b1011;
															assign node2005 = (inp[3]) ? node2007 : 4'b1001;
																assign node2007 = (inp[15]) ? 4'b1001 : 4'b1011;
											assign node2010 = (inp[9]) ? node2040 : node2011;
												assign node2011 = (inp[3]) ? node2031 : node2012;
													assign node2012 = (inp[12]) ? node2020 : node2013;
														assign node2013 = (inp[5]) ? 4'b1001 : node2014;
															assign node2014 = (inp[15]) ? 4'b1011 : node2015;
																assign node2015 = (inp[0]) ? 4'b1001 : 4'b1011;
														assign node2020 = (inp[5]) ? node2026 : node2021;
															assign node2021 = (inp[15]) ? node2023 : 4'b1011;
																assign node2023 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node2026 = (inp[0]) ? node2028 : 4'b1011;
																assign node2028 = (inp[15]) ? 4'b1011 : 4'b1001;
													assign node2031 = (inp[5]) ? node2033 : 4'b1001;
														assign node2033 = (inp[15]) ? node2037 : node2034;
															assign node2034 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node2037 = (inp[0]) ? 4'b1001 : 4'b1011;
												assign node2040 = (inp[5]) ? node2054 : node2041;
													assign node2041 = (inp[3]) ? node2047 : node2042;
														assign node2042 = (inp[15]) ? 4'b1111 : node2043;
															assign node2043 = (inp[0]) ? 4'b1101 : 4'b1111;
														assign node2047 = (inp[15]) ? node2051 : node2048;
															assign node2048 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node2051 = (inp[0]) ? 4'b1101 : 4'b1111;
													assign node2054 = (inp[3]) ? node2064 : node2055;
														assign node2055 = (inp[12]) ? node2061 : node2056;
															assign node2056 = (inp[0]) ? node2058 : 4'b1101;
																assign node2058 = (inp[15]) ? 4'b1101 : 4'b1111;
															assign node2061 = (inp[0]) ? 4'b1101 : 4'b1111;
														assign node2064 = (inp[12]) ? node2072 : node2065;
															assign node2065 = (inp[15]) ? node2069 : node2066;
																assign node2066 = (inp[0]) ? 4'b1111 : 4'b1101;
																assign node2069 = (inp[0]) ? 4'b1101 : 4'b1111;
															assign node2072 = (inp[0]) ? node2076 : node2073;
																assign node2073 = (inp[15]) ? 4'b1111 : 4'b1101;
																assign node2076 = (inp[15]) ? 4'b1101 : 4'b1111;
										assign node2079 = (inp[5]) ? node2133 : node2080;
											assign node2080 = (inp[0]) ? node2100 : node2081;
												assign node2081 = (inp[15]) ? node2091 : node2082;
													assign node2082 = (inp[4]) ? node2086 : node2083;
														assign node2083 = (inp[9]) ? 4'b1010 : 4'b1110;
														assign node2086 = (inp[9]) ? node2088 : 4'b1010;
															assign node2088 = (inp[3]) ? 4'b1100 : 4'b1110;
													assign node2091 = (inp[3]) ? 4'b1000 : node2092;
														assign node2092 = (inp[9]) ? node2096 : node2093;
															assign node2093 = (inp[4]) ? 4'b1000 : 4'b1100;
															assign node2096 = (inp[4]) ? 4'b1100 : 4'b1000;
												assign node2100 = (inp[15]) ? node2114 : node2101;
													assign node2101 = (inp[3]) ? node2109 : node2102;
														assign node2102 = (inp[9]) ? node2106 : node2103;
															assign node2103 = (inp[4]) ? 4'b1000 : 4'b1100;
															assign node2106 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node2109 = (inp[9]) ? node2111 : 4'b1000;
															assign node2111 = (inp[4]) ? 4'b1110 : 4'b1000;
													assign node2114 = (inp[12]) ? node2120 : node2115;
														assign node2115 = (inp[4]) ? node2117 : 4'b1110;
															assign node2117 = (inp[3]) ? 4'b1010 : 4'b1110;
														assign node2120 = (inp[3]) ? node2128 : node2121;
															assign node2121 = (inp[9]) ? node2125 : node2122;
																assign node2122 = (inp[4]) ? 4'b1010 : 4'b1110;
																assign node2125 = (inp[4]) ? 4'b1110 : 4'b1010;
															assign node2128 = (inp[4]) ? node2130 : 4'b1010;
																assign node2130 = (inp[9]) ? 4'b1100 : 4'b1010;
											assign node2133 = (inp[12]) ? node2169 : node2134;
												assign node2134 = (inp[9]) ? node2152 : node2135;
													assign node2135 = (inp[4]) ? node2149 : node2136;
														assign node2136 = (inp[15]) ? node2142 : node2137;
															assign node2137 = (inp[3]) ? node2139 : 4'b1100;
																assign node2139 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node2142 = (inp[0]) ? node2146 : node2143;
																assign node2143 = (inp[3]) ? 4'b1110 : 4'b1100;
																assign node2146 = (inp[3]) ? 4'b1100 : 4'b1110;
														assign node2149 = (inp[3]) ? 4'b1000 : 4'b1010;
													assign node2152 = (inp[4]) ? node2164 : node2153;
														assign node2153 = (inp[3]) ? node2159 : node2154;
															assign node2154 = (inp[0]) ? node2156 : 4'b1000;
																assign node2156 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node2159 = (inp[0]) ? node2161 : 4'b1010;
																assign node2161 = (inp[15]) ? 4'b1000 : 4'b1010;
														assign node2164 = (inp[15]) ? node2166 : 4'b1100;
															assign node2166 = (inp[0]) ? 4'b1100 : 4'b1110;
												assign node2169 = (inp[4]) ? node2191 : node2170;
													assign node2170 = (inp[9]) ? node2186 : node2171;
														assign node2171 = (inp[3]) ? node2179 : node2172;
															assign node2172 = (inp[15]) ? node2176 : node2173;
																assign node2173 = (inp[0]) ? 4'b1100 : 4'b1110;
																assign node2176 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node2179 = (inp[15]) ? node2183 : node2180;
																assign node2180 = (inp[0]) ? 4'b1110 : 4'b1100;
																assign node2183 = (inp[0]) ? 4'b1100 : 4'b1110;
														assign node2186 = (inp[15]) ? node2188 : 4'b1010;
															assign node2188 = (inp[3]) ? 4'b1010 : 4'b1000;
													assign node2191 = (inp[9]) ? node2205 : node2192;
														assign node2192 = (inp[0]) ? node2198 : node2193;
															assign node2193 = (inp[3]) ? node2195 : 4'b1010;
																assign node2195 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node2198 = (inp[3]) ? node2202 : node2199;
																assign node2199 = (inp[15]) ? 4'b1010 : 4'b1000;
																assign node2202 = (inp[15]) ? 4'b1000 : 4'b1010;
														assign node2205 = (inp[15]) ? node2209 : node2206;
															assign node2206 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node2209 = (inp[0]) ? 4'b1100 : 4'b1110;
									assign node2212 = (inp[15]) ? node2278 : node2213;
										assign node2213 = (inp[0]) ? node2247 : node2214;
											assign node2214 = (inp[5]) ? node2224 : node2215;
												assign node2215 = (inp[9]) ? node2219 : node2216;
													assign node2216 = (inp[4]) ? 4'b1010 : 4'b1110;
													assign node2219 = (inp[4]) ? node2221 : 4'b1010;
														assign node2221 = (inp[3]) ? 4'b1100 : 4'b1110;
												assign node2224 = (inp[3]) ? node2232 : node2225;
													assign node2225 = (inp[9]) ? node2229 : node2226;
														assign node2226 = (inp[4]) ? 4'b1010 : 4'b1110;
														assign node2229 = (inp[4]) ? 4'b1100 : 4'b1010;
													assign node2232 = (inp[12]) ? node2240 : node2233;
														assign node2233 = (inp[9]) ? node2237 : node2234;
															assign node2234 = (inp[4]) ? 4'b1000 : 4'b1100;
															assign node2237 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node2240 = (inp[9]) ? node2244 : node2241;
															assign node2241 = (inp[4]) ? 4'b1000 : 4'b1100;
															assign node2244 = (inp[4]) ? 4'b1100 : 4'b1000;
											assign node2247 = (inp[3]) ? node2257 : node2248;
												assign node2248 = (inp[9]) ? node2252 : node2249;
													assign node2249 = (inp[4]) ? 4'b1000 : 4'b1100;
													assign node2252 = (inp[4]) ? node2254 : 4'b1000;
														assign node2254 = (inp[2]) ? 4'b1100 : 4'b1110;
												assign node2257 = (inp[5]) ? node2265 : node2258;
													assign node2258 = (inp[4]) ? node2262 : node2259;
														assign node2259 = (inp[9]) ? 4'b1000 : 4'b1100;
														assign node2262 = (inp[9]) ? 4'b1110 : 4'b1000;
													assign node2265 = (inp[2]) ? node2273 : node2266;
														assign node2266 = (inp[4]) ? node2270 : node2267;
															assign node2267 = (inp[12]) ? 4'b1110 : 4'b1010;
															assign node2270 = (inp[12]) ? 4'b1010 : 4'b1110;
														assign node2273 = (inp[9]) ? 4'b1110 : node2274;
															assign node2274 = (inp[4]) ? 4'b1010 : 4'b1110;
										assign node2278 = (inp[0]) ? node2304 : node2279;
											assign node2279 = (inp[3]) ? node2289 : node2280;
												assign node2280 = (inp[9]) ? node2284 : node2281;
													assign node2281 = (inp[4]) ? 4'b1000 : 4'b1100;
													assign node2284 = (inp[4]) ? node2286 : 4'b1000;
														assign node2286 = (inp[5]) ? 4'b1110 : 4'b1100;
												assign node2289 = (inp[5]) ? node2297 : node2290;
													assign node2290 = (inp[4]) ? node2294 : node2291;
														assign node2291 = (inp[9]) ? 4'b1000 : 4'b1100;
														assign node2294 = (inp[9]) ? 4'b1110 : 4'b1000;
													assign node2297 = (inp[4]) ? node2301 : node2298;
														assign node2298 = (inp[9]) ? 4'b1010 : 4'b1110;
														assign node2301 = (inp[9]) ? 4'b1110 : 4'b1010;
											assign node2304 = (inp[3]) ? node2314 : node2305;
												assign node2305 = (inp[9]) ? node2309 : node2306;
													assign node2306 = (inp[4]) ? 4'b1010 : 4'b1110;
													assign node2309 = (inp[4]) ? node2311 : 4'b1010;
														assign node2311 = (inp[5]) ? 4'b1100 : 4'b1110;
												assign node2314 = (inp[5]) ? node2322 : node2315;
													assign node2315 = (inp[4]) ? node2319 : node2316;
														assign node2316 = (inp[9]) ? 4'b1010 : 4'b1110;
														assign node2319 = (inp[9]) ? 4'b1100 : 4'b1010;
													assign node2322 = (inp[12]) ? node2328 : node2323;
														assign node2323 = (inp[4]) ? node2325 : 4'b1100;
															assign node2325 = (inp[9]) ? 4'b1100 : 4'b1000;
														assign node2328 = (inp[4]) ? node2332 : node2329;
															assign node2329 = (inp[9]) ? 4'b1000 : 4'b1100;
															assign node2332 = (inp[9]) ? 4'b1100 : 4'b1000;
								assign node2335 = (inp[14]) ? node2559 : node2336;
									assign node2336 = (inp[2]) ? node2440 : node2337;
										assign node2337 = (inp[15]) ? node2401 : node2338;
											assign node2338 = (inp[12]) ? node2368 : node2339;
												assign node2339 = (inp[0]) ? node2355 : node2340;
													assign node2340 = (inp[5]) ? node2348 : node2341;
														assign node2341 = (inp[3]) ? 4'b1010 : node2342;
															assign node2342 = (inp[4]) ? node2344 : 4'b1110;
																assign node2344 = (inp[9]) ? 4'b1110 : 4'b1010;
														assign node2348 = (inp[4]) ? node2352 : node2349;
															assign node2349 = (inp[3]) ? 4'b1100 : 4'b1010;
															assign node2352 = (inp[9]) ? 4'b1100 : 4'b1000;
													assign node2355 = (inp[5]) ? node2361 : node2356;
														assign node2356 = (inp[9]) ? 4'b1000 : node2357;
															assign node2357 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node2361 = (inp[4]) ? 4'b1110 : node2362;
															assign node2362 = (inp[9]) ? node2364 : 4'b1110;
																assign node2364 = (inp[3]) ? 4'b1010 : 4'b1000;
												assign node2368 = (inp[0]) ? node2382 : node2369;
													assign node2369 = (inp[5]) ? node2375 : node2370;
														assign node2370 = (inp[9]) ? 4'b1010 : node2371;
															assign node2371 = (inp[4]) ? 4'b1010 : 4'b1110;
														assign node2375 = (inp[3]) ? 4'b1000 : node2376;
															assign node2376 = (inp[4]) ? node2378 : 4'b1010;
																assign node2378 = (inp[9]) ? 4'b1100 : 4'b1010;
													assign node2382 = (inp[5]) ? node2392 : node2383;
														assign node2383 = (inp[3]) ? node2385 : 4'b1000;
															assign node2385 = (inp[4]) ? node2389 : node2386;
																assign node2386 = (inp[9]) ? 4'b1000 : 4'b1100;
																assign node2389 = (inp[9]) ? 4'b1110 : 4'b1000;
														assign node2392 = (inp[3]) ? node2396 : node2393;
															assign node2393 = (inp[4]) ? 4'b1110 : 4'b1000;
															assign node2396 = (inp[4]) ? 4'b1010 : node2397;
																assign node2397 = (inp[9]) ? 4'b1010 : 4'b1110;
											assign node2401 = (inp[9]) ? node2423 : node2402;
												assign node2402 = (inp[4]) ? node2412 : node2403;
													assign node2403 = (inp[5]) ? node2407 : node2404;
														assign node2404 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node2407 = (inp[12]) ? 4'b1110 : node2408;
															assign node2408 = (inp[0]) ? 4'b1100 : 4'b1110;
													assign node2412 = (inp[0]) ? node2418 : node2413;
														assign node2413 = (inp[3]) ? node2415 : 4'b1000;
															assign node2415 = (inp[5]) ? 4'b1010 : 4'b1000;
														assign node2418 = (inp[12]) ? 4'b1010 : node2419;
															assign node2419 = (inp[5]) ? 4'b1000 : 4'b1010;
												assign node2423 = (inp[4]) ? node2433 : node2424;
													assign node2424 = (inp[5]) ? node2428 : node2425;
														assign node2425 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node2428 = (inp[3]) ? node2430 : 4'b1000;
															assign node2430 = (inp[0]) ? 4'b1000 : 4'b1010;
													assign node2433 = (inp[0]) ? 4'b1100 : node2434;
														assign node2434 = (inp[3]) ? 4'b1110 : node2435;
															assign node2435 = (inp[5]) ? 4'b1110 : 4'b1100;
										assign node2440 = (inp[12]) ? node2490 : node2441;
											assign node2441 = (inp[9]) ? node2469 : node2442;
												assign node2442 = (inp[4]) ? node2460 : node2443;
													assign node2443 = (inp[15]) ? node2455 : node2444;
														assign node2444 = (inp[0]) ? node2450 : node2445;
															assign node2445 = (inp[3]) ? node2447 : 4'b0111;
																assign node2447 = (inp[5]) ? 4'b0101 : 4'b0111;
															assign node2450 = (inp[5]) ? node2452 : 4'b0101;
																assign node2452 = (inp[3]) ? 4'b0111 : 4'b0101;
														assign node2455 = (inp[0]) ? 4'b0111 : node2456;
															assign node2456 = (inp[3]) ? 4'b0111 : 4'b0101;
													assign node2460 = (inp[5]) ? node2462 : 4'b0011;
														assign node2462 = (inp[15]) ? 4'b0001 : node2463;
															assign node2463 = (inp[3]) ? 4'b0011 : node2464;
																assign node2464 = (inp[0]) ? 4'b0001 : 4'b0011;
												assign node2469 = (inp[4]) ? node2475 : node2470;
													assign node2470 = (inp[5]) ? node2472 : 4'b0001;
														assign node2472 = (inp[15]) ? 4'b0011 : 4'b0001;
													assign node2475 = (inp[5]) ? node2485 : node2476;
														assign node2476 = (inp[15]) ? node2478 : 4'b0111;
															assign node2478 = (inp[0]) ? node2482 : node2479;
																assign node2479 = (inp[3]) ? 4'b0111 : 4'b0101;
																assign node2482 = (inp[3]) ? 4'b0101 : 4'b0111;
														assign node2485 = (inp[0]) ? 4'b0101 : node2486;
															assign node2486 = (inp[15]) ? 4'b0111 : 4'b0101;
											assign node2490 = (inp[15]) ? node2520 : node2491;
												assign node2491 = (inp[3]) ? node2509 : node2492;
													assign node2492 = (inp[0]) ? node2500 : node2493;
														assign node2493 = (inp[9]) ? node2497 : node2494;
															assign node2494 = (inp[4]) ? 4'b0011 : 4'b0111;
															assign node2497 = (inp[5]) ? 4'b0101 : 4'b0111;
														assign node2500 = (inp[5]) ? node2506 : node2501;
															assign node2501 = (inp[9]) ? 4'b0001 : node2502;
																assign node2502 = (inp[4]) ? 4'b0001 : 4'b0101;
															assign node2506 = (inp[9]) ? 4'b0111 : 4'b0001;
													assign node2509 = (inp[5]) ? node2515 : node2510;
														assign node2510 = (inp[0]) ? 4'b0111 : node2511;
															assign node2511 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node2515 = (inp[0]) ? node2517 : 4'b0001;
															assign node2517 = (inp[4]) ? 4'b0111 : 4'b0011;
												assign node2520 = (inp[0]) ? node2536 : node2521;
													assign node2521 = (inp[5]) ? node2529 : node2522;
														assign node2522 = (inp[3]) ? 4'b0001 : node2523;
															assign node2523 = (inp[9]) ? 4'b0001 : node2524;
																assign node2524 = (inp[4]) ? 4'b0001 : 4'b0101;
														assign node2529 = (inp[3]) ? node2533 : node2530;
															assign node2530 = (inp[9]) ? 4'b0001 : 4'b0101;
															assign node2533 = (inp[4]) ? 4'b0011 : 4'b0111;
													assign node2536 = (inp[5]) ? node2546 : node2537;
														assign node2537 = (inp[3]) ? 4'b0011 : node2538;
															assign node2538 = (inp[4]) ? node2542 : node2539;
																assign node2539 = (inp[9]) ? 4'b0011 : 4'b0111;
																assign node2542 = (inp[9]) ? 4'b0111 : 4'b0011;
														assign node2546 = (inp[3]) ? node2552 : node2547;
															assign node2547 = (inp[4]) ? 4'b0101 : node2548;
																assign node2548 = (inp[9]) ? 4'b0011 : 4'b0111;
															assign node2552 = (inp[4]) ? node2556 : node2553;
																assign node2553 = (inp[9]) ? 4'b0001 : 4'b0101;
																assign node2556 = (inp[9]) ? 4'b0101 : 4'b0001;
									assign node2559 = (inp[4]) ? node2677 : node2560;
										assign node2560 = (inp[9]) ? node2600 : node2561;
											assign node2561 = (inp[2]) ? node2581 : node2562;
												assign node2562 = (inp[5]) ? node2570 : node2563;
													assign node2563 = (inp[15]) ? node2567 : node2564;
														assign node2564 = (inp[0]) ? 4'b0101 : 4'b0111;
														assign node2567 = (inp[0]) ? 4'b0111 : 4'b0101;
													assign node2570 = (inp[12]) ? node2572 : 4'b0111;
														assign node2572 = (inp[15]) ? node2574 : 4'b0111;
															assign node2574 = (inp[3]) ? node2578 : node2575;
																assign node2575 = (inp[0]) ? 4'b0111 : 4'b0101;
																assign node2578 = (inp[0]) ? 4'b0101 : 4'b0111;
												assign node2581 = (inp[3]) ? node2587 : node2582;
													assign node2582 = (inp[15]) ? node2584 : 4'b0101;
														assign node2584 = (inp[0]) ? 4'b0111 : 4'b0101;
													assign node2587 = (inp[5]) ? node2595 : node2588;
														assign node2588 = (inp[15]) ? node2592 : node2589;
															assign node2589 = (inp[0]) ? 4'b0101 : 4'b0111;
															assign node2592 = (inp[0]) ? 4'b0111 : 4'b0101;
														assign node2595 = (inp[15]) ? 4'b0111 : node2596;
															assign node2596 = (inp[0]) ? 4'b0111 : 4'b0101;
											assign node2600 = (inp[12]) ? node2644 : node2601;
												assign node2601 = (inp[5]) ? node2627 : node2602;
													assign node2602 = (inp[3]) ? node2612 : node2603;
														assign node2603 = (inp[2]) ? node2605 : 4'b0011;
															assign node2605 = (inp[15]) ? node2609 : node2606;
																assign node2606 = (inp[0]) ? 4'b0001 : 4'b0011;
																assign node2609 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node2612 = (inp[2]) ? node2620 : node2613;
															assign node2613 = (inp[0]) ? node2617 : node2614;
																assign node2614 = (inp[15]) ? 4'b0001 : 4'b0011;
																assign node2617 = (inp[15]) ? 4'b0011 : 4'b0001;
															assign node2620 = (inp[0]) ? node2624 : node2621;
																assign node2621 = (inp[15]) ? 4'b0001 : 4'b0011;
																assign node2624 = (inp[15]) ? 4'b0011 : 4'b0001;
													assign node2627 = (inp[3]) ? node2635 : node2628;
														assign node2628 = (inp[0]) ? node2632 : node2629;
															assign node2629 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node2632 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node2635 = (inp[2]) ? 4'b0011 : node2636;
															assign node2636 = (inp[15]) ? node2640 : node2637;
																assign node2637 = (inp[0]) ? 4'b0011 : 4'b0001;
																assign node2640 = (inp[0]) ? 4'b0001 : 4'b0011;
												assign node2644 = (inp[3]) ? node2662 : node2645;
													assign node2645 = (inp[5]) ? node2655 : node2646;
														assign node2646 = (inp[2]) ? node2652 : node2647;
															assign node2647 = (inp[15]) ? node2649 : 4'b0011;
																assign node2649 = (inp[0]) ? 4'b0011 : 4'b0001;
															assign node2652 = (inp[0]) ? 4'b0001 : 4'b0011;
														assign node2655 = (inp[15]) ? node2659 : node2656;
															assign node2656 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node2659 = (inp[0]) ? 4'b0011 : 4'b0001;
													assign node2662 = (inp[5]) ? node2670 : node2663;
														assign node2663 = (inp[0]) ? node2667 : node2664;
															assign node2664 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node2667 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node2670 = (inp[0]) ? node2674 : node2671;
															assign node2671 = (inp[15]) ? 4'b0011 : 4'b0001;
															assign node2674 = (inp[15]) ? 4'b0001 : 4'b0011;
										assign node2677 = (inp[9]) ? node2717 : node2678;
											assign node2678 = (inp[12]) ? node2704 : node2679;
												assign node2679 = (inp[3]) ? node2695 : node2680;
													assign node2680 = (inp[2]) ? node2688 : node2681;
														assign node2681 = (inp[15]) ? node2685 : node2682;
															assign node2682 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node2685 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node2688 = (inp[15]) ? node2692 : node2689;
															assign node2689 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node2692 = (inp[0]) ? 4'b0011 : 4'b0001;
													assign node2695 = (inp[0]) ? 4'b0001 : node2696;
														assign node2696 = (inp[5]) ? node2700 : node2697;
															assign node2697 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node2700 = (inp[15]) ? 4'b0011 : 4'b0001;
												assign node2704 = (inp[0]) ? node2712 : node2705;
													assign node2705 = (inp[15]) ? node2707 : 4'b0011;
														assign node2707 = (inp[5]) ? node2709 : 4'b0001;
															assign node2709 = (inp[3]) ? 4'b0011 : 4'b0001;
													assign node2712 = (inp[15]) ? 4'b0011 : node2713;
														assign node2713 = (inp[3]) ? 4'b0011 : 4'b0001;
											assign node2717 = (inp[0]) ? node2729 : node2718;
												assign node2718 = (inp[15]) ? node2724 : node2719;
													assign node2719 = (inp[5]) ? 4'b0101 : node2720;
														assign node2720 = (inp[3]) ? 4'b0101 : 4'b0111;
													assign node2724 = (inp[3]) ? 4'b0111 : node2725;
														assign node2725 = (inp[5]) ? 4'b0111 : 4'b0101;
												assign node2729 = (inp[15]) ? node2735 : node2730;
													assign node2730 = (inp[5]) ? 4'b0111 : node2731;
														assign node2731 = (inp[3]) ? 4'b0111 : 4'b0101;
													assign node2735 = (inp[3]) ? 4'b0101 : node2736;
														assign node2736 = (inp[5]) ? 4'b0101 : 4'b0111;
							assign node2740 = (inp[8]) ? node3076 : node2741;
								assign node2741 = (inp[2]) ? node2929 : node2742;
									assign node2742 = (inp[14]) ? node2836 : node2743;
										assign node2743 = (inp[9]) ? node2797 : node2744;
											assign node2744 = (inp[4]) ? node2776 : node2745;
												assign node2745 = (inp[3]) ? node2753 : node2746;
													assign node2746 = (inp[15]) ? node2750 : node2747;
														assign node2747 = (inp[0]) ? 4'b1100 : 4'b1110;
														assign node2750 = (inp[0]) ? 4'b1110 : 4'b1100;
													assign node2753 = (inp[12]) ? node2767 : node2754;
														assign node2754 = (inp[15]) ? node2762 : node2755;
															assign node2755 = (inp[5]) ? node2759 : node2756;
																assign node2756 = (inp[0]) ? 4'b1100 : 4'b1110;
																assign node2759 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node2762 = (inp[5]) ? 4'b1110 : node2763;
																assign node2763 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node2767 = (inp[5]) ? 4'b1100 : node2768;
															assign node2768 = (inp[0]) ? node2772 : node2769;
																assign node2769 = (inp[15]) ? 4'b1100 : 4'b1110;
																assign node2772 = (inp[15]) ? 4'b1110 : 4'b1100;
												assign node2776 = (inp[0]) ? node2788 : node2777;
													assign node2777 = (inp[15]) ? node2783 : node2778;
														assign node2778 = (inp[3]) ? node2780 : 4'b1010;
															assign node2780 = (inp[5]) ? 4'b1000 : 4'b1010;
														assign node2783 = (inp[5]) ? node2785 : 4'b1000;
															assign node2785 = (inp[3]) ? 4'b1010 : 4'b1000;
													assign node2788 = (inp[15]) ? node2792 : node2789;
														assign node2789 = (inp[3]) ? 4'b1010 : 4'b1000;
														assign node2792 = (inp[3]) ? node2794 : 4'b1010;
															assign node2794 = (inp[12]) ? 4'b1010 : 4'b1000;
											assign node2797 = (inp[4]) ? node2815 : node2798;
												assign node2798 = (inp[15]) ? node2808 : node2799;
													assign node2799 = (inp[0]) ? node2805 : node2800;
														assign node2800 = (inp[5]) ? node2802 : 4'b1010;
															assign node2802 = (inp[3]) ? 4'b1000 : 4'b1010;
														assign node2805 = (inp[3]) ? 4'b1010 : 4'b1000;
													assign node2808 = (inp[0]) ? node2810 : 4'b1000;
														assign node2810 = (inp[5]) ? node2812 : 4'b1010;
															assign node2812 = (inp[3]) ? 4'b1000 : 4'b1010;
												assign node2815 = (inp[0]) ? node2825 : node2816;
													assign node2816 = (inp[3]) ? 4'b1100 : node2817;
														assign node2817 = (inp[12]) ? node2819 : 4'b1100;
															assign node2819 = (inp[5]) ? 4'b1110 : node2820;
																assign node2820 = (inp[15]) ? 4'b1100 : 4'b1110;
													assign node2825 = (inp[15]) ? node2831 : node2826;
														assign node2826 = (inp[5]) ? 4'b1110 : node2827;
															assign node2827 = (inp[3]) ? 4'b1110 : 4'b1100;
														assign node2831 = (inp[5]) ? 4'b1100 : node2832;
															assign node2832 = (inp[3]) ? 4'b1100 : 4'b1110;
										assign node2836 = (inp[3]) ? node2880 : node2837;
											assign node2837 = (inp[4]) ? node2859 : node2838;
												assign node2838 = (inp[9]) ? node2846 : node2839;
													assign node2839 = (inp[0]) ? node2843 : node2840;
														assign node2840 = (inp[15]) ? 4'b0101 : 4'b0111;
														assign node2843 = (inp[15]) ? 4'b0111 : 4'b0101;
													assign node2846 = (inp[12]) ? node2852 : node2847;
														assign node2847 = (inp[5]) ? 4'b0001 : node2848;
															assign node2848 = (inp[15]) ? 4'b0001 : 4'b0011;
														assign node2852 = (inp[15]) ? node2856 : node2853;
															assign node2853 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node2856 = (inp[0]) ? 4'b0011 : 4'b0001;
												assign node2859 = (inp[9]) ? node2873 : node2860;
													assign node2860 = (inp[5]) ? node2868 : node2861;
														assign node2861 = (inp[15]) ? node2865 : node2862;
															assign node2862 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node2865 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node2868 = (inp[0]) ? node2870 : 4'b0011;
															assign node2870 = (inp[15]) ? 4'b0011 : 4'b0001;
													assign node2873 = (inp[0]) ? node2875 : 4'b0111;
														assign node2875 = (inp[5]) ? node2877 : 4'b0101;
															assign node2877 = (inp[15]) ? 4'b0101 : 4'b0111;
											assign node2880 = (inp[4]) ? node2912 : node2881;
												assign node2881 = (inp[9]) ? node2899 : node2882;
													assign node2882 = (inp[15]) ? node2892 : node2883;
														assign node2883 = (inp[12]) ? 4'b0101 : node2884;
															assign node2884 = (inp[0]) ? node2888 : node2885;
																assign node2885 = (inp[5]) ? 4'b0101 : 4'b0111;
																assign node2888 = (inp[5]) ? 4'b0111 : 4'b0101;
														assign node2892 = (inp[5]) ? node2896 : node2893;
															assign node2893 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node2896 = (inp[0]) ? 4'b0101 : 4'b0111;
													assign node2899 = (inp[15]) ? node2907 : node2900;
														assign node2900 = (inp[12]) ? node2902 : 4'b0011;
															assign node2902 = (inp[0]) ? node2904 : 4'b0011;
																assign node2904 = (inp[5]) ? 4'b0011 : 4'b0001;
														assign node2907 = (inp[5]) ? 4'b0001 : node2908;
															assign node2908 = (inp[0]) ? 4'b0011 : 4'b0001;
												assign node2912 = (inp[9]) ? node2924 : node2913;
													assign node2913 = (inp[5]) ? node2919 : node2914;
														assign node2914 = (inp[0]) ? node2916 : 4'b0011;
															assign node2916 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node2919 = (inp[0]) ? node2921 : 4'b0001;
															assign node2921 = (inp[15]) ? 4'b0001 : 4'b0011;
													assign node2924 = (inp[0]) ? node2926 : 4'b0101;
														assign node2926 = (inp[15]) ? 4'b0101 : 4'b0111;
									assign node2929 = (inp[5]) ? node2997 : node2930;
										assign node2930 = (inp[15]) ? node2970 : node2931;
											assign node2931 = (inp[0]) ? node2941 : node2932;
												assign node2932 = (inp[4]) ? node2936 : node2933;
													assign node2933 = (inp[9]) ? 4'b0011 : 4'b0111;
													assign node2936 = (inp[3]) ? 4'b0101 : node2937;
														assign node2937 = (inp[9]) ? 4'b0111 : 4'b0011;
												assign node2941 = (inp[3]) ? node2963 : node2942;
													assign node2942 = (inp[14]) ? node2956 : node2943;
														assign node2943 = (inp[12]) ? node2949 : node2944;
															assign node2944 = (inp[4]) ? 4'b0001 : node2945;
																assign node2945 = (inp[9]) ? 4'b0001 : 4'b0101;
															assign node2949 = (inp[9]) ? node2953 : node2950;
																assign node2950 = (inp[4]) ? 4'b0001 : 4'b0101;
																assign node2953 = (inp[4]) ? 4'b0101 : 4'b0001;
														assign node2956 = (inp[9]) ? node2960 : node2957;
															assign node2957 = (inp[4]) ? 4'b0001 : 4'b0101;
															assign node2960 = (inp[4]) ? 4'b0101 : 4'b0001;
													assign node2963 = (inp[9]) ? node2967 : node2964;
														assign node2964 = (inp[4]) ? 4'b0001 : 4'b0101;
														assign node2967 = (inp[4]) ? 4'b0111 : 4'b0001;
											assign node2970 = (inp[0]) ? node2990 : node2971;
												assign node2971 = (inp[14]) ? node2985 : node2972;
													assign node2972 = (inp[3]) ? node2980 : node2973;
														assign node2973 = (inp[4]) ? node2977 : node2974;
															assign node2974 = (inp[9]) ? 4'b0001 : 4'b0101;
															assign node2977 = (inp[9]) ? 4'b0101 : 4'b0001;
														assign node2980 = (inp[9]) ? 4'b0001 : node2981;
															assign node2981 = (inp[4]) ? 4'b0001 : 4'b0101;
													assign node2985 = (inp[4]) ? node2987 : 4'b0001;
														assign node2987 = (inp[9]) ? 4'b0111 : 4'b0001;
												assign node2990 = (inp[9]) ? node2994 : node2991;
													assign node2991 = (inp[4]) ? 4'b0011 : 4'b0111;
													assign node2994 = (inp[3]) ? 4'b0101 : 4'b0111;
										assign node2997 = (inp[3]) ? node3031 : node2998;
											assign node2998 = (inp[0]) ? node3014 : node2999;
												assign node2999 = (inp[15]) ? node3007 : node3000;
													assign node3000 = (inp[9]) ? node3004 : node3001;
														assign node3001 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node3004 = (inp[4]) ? 4'b0101 : 4'b0011;
													assign node3007 = (inp[9]) ? node3011 : node3008;
														assign node3008 = (inp[4]) ? 4'b0001 : 4'b0101;
														assign node3011 = (inp[4]) ? 4'b0111 : 4'b0001;
												assign node3014 = (inp[15]) ? node3024 : node3015;
													assign node3015 = (inp[12]) ? node3017 : 4'b0001;
														assign node3017 = (inp[9]) ? node3021 : node3018;
															assign node3018 = (inp[4]) ? 4'b0001 : 4'b0101;
															assign node3021 = (inp[4]) ? 4'b0111 : 4'b0001;
													assign node3024 = (inp[9]) ? node3028 : node3025;
														assign node3025 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node3028 = (inp[4]) ? 4'b0101 : 4'b0011;
											assign node3031 = (inp[0]) ? node3047 : node3032;
												assign node3032 = (inp[15]) ? node3040 : node3033;
													assign node3033 = (inp[9]) ? node3037 : node3034;
														assign node3034 = (inp[4]) ? 4'b0001 : 4'b0101;
														assign node3037 = (inp[4]) ? 4'b0101 : 4'b0001;
													assign node3040 = (inp[9]) ? node3044 : node3041;
														assign node3041 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node3044 = (inp[4]) ? 4'b0111 : 4'b0011;
												assign node3047 = (inp[15]) ? node3069 : node3048;
													assign node3048 = (inp[12]) ? node3062 : node3049;
														assign node3049 = (inp[14]) ? node3057 : node3050;
															assign node3050 = (inp[9]) ? node3054 : node3051;
																assign node3051 = (inp[4]) ? 4'b0011 : 4'b0111;
																assign node3054 = (inp[4]) ? 4'b0111 : 4'b0011;
															assign node3057 = (inp[9]) ? 4'b0111 : node3058;
																assign node3058 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node3062 = (inp[4]) ? node3066 : node3063;
															assign node3063 = (inp[9]) ? 4'b0011 : 4'b0111;
															assign node3066 = (inp[9]) ? 4'b0111 : 4'b0011;
													assign node3069 = (inp[4]) ? node3073 : node3070;
														assign node3070 = (inp[9]) ? 4'b0001 : 4'b0101;
														assign node3073 = (inp[9]) ? 4'b0101 : 4'b0001;
								assign node3076 = (inp[2]) ? node3264 : node3077;
									assign node3077 = (inp[14]) ? node3175 : node3078;
										assign node3078 = (inp[4]) ? node3118 : node3079;
											assign node3079 = (inp[9]) ? node3103 : node3080;
												assign node3080 = (inp[15]) ? node3092 : node3081;
													assign node3081 = (inp[0]) ? node3087 : node3082;
														assign node3082 = (inp[5]) ? node3084 : 4'b0111;
															assign node3084 = (inp[3]) ? 4'b0101 : 4'b0111;
														assign node3087 = (inp[3]) ? node3089 : 4'b0101;
															assign node3089 = (inp[5]) ? 4'b0111 : 4'b0101;
													assign node3092 = (inp[0]) ? node3096 : node3093;
														assign node3093 = (inp[12]) ? 4'b0101 : 4'b0111;
														assign node3096 = (inp[12]) ? 4'b0111 : node3097;
															assign node3097 = (inp[5]) ? node3099 : 4'b0111;
																assign node3099 = (inp[3]) ? 4'b0101 : 4'b0111;
												assign node3103 = (inp[15]) ? node3107 : node3104;
													assign node3104 = (inp[0]) ? 4'b0001 : 4'b0011;
													assign node3107 = (inp[0]) ? node3113 : node3108;
														assign node3108 = (inp[3]) ? node3110 : 4'b0001;
															assign node3110 = (inp[5]) ? 4'b0011 : 4'b0001;
														assign node3113 = (inp[3]) ? node3115 : 4'b0011;
															assign node3115 = (inp[5]) ? 4'b0001 : 4'b0011;
											assign node3118 = (inp[9]) ? node3138 : node3119;
												assign node3119 = (inp[5]) ? node3127 : node3120;
													assign node3120 = (inp[0]) ? node3124 : node3121;
														assign node3121 = (inp[15]) ? 4'b0001 : 4'b0011;
														assign node3124 = (inp[15]) ? 4'b0011 : 4'b0001;
													assign node3127 = (inp[15]) ? 4'b0001 : node3128;
														assign node3128 = (inp[12]) ? node3132 : node3129;
															assign node3129 = (inp[3]) ? 4'b0011 : 4'b0001;
															assign node3132 = (inp[3]) ? 4'b0001 : node3133;
																assign node3133 = (inp[0]) ? 4'b0001 : 4'b0011;
												assign node3138 = (inp[12]) ? node3152 : node3139;
													assign node3139 = (inp[15]) ? node3147 : node3140;
														assign node3140 = (inp[0]) ? node3142 : 4'b0101;
															assign node3142 = (inp[5]) ? 4'b0111 : node3143;
																assign node3143 = (inp[3]) ? 4'b0111 : 4'b0101;
														assign node3147 = (inp[0]) ? 4'b0101 : node3148;
															assign node3148 = (inp[3]) ? 4'b0111 : 4'b0101;
													assign node3152 = (inp[5]) ? node3166 : node3153;
														assign node3153 = (inp[15]) ? node3161 : node3154;
															assign node3154 = (inp[3]) ? node3158 : node3155;
																assign node3155 = (inp[0]) ? 4'b0101 : 4'b0111;
																assign node3158 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node3161 = (inp[0]) ? 4'b0101 : node3162;
																assign node3162 = (inp[3]) ? 4'b0111 : 4'b0101;
														assign node3166 = (inp[3]) ? 4'b0111 : node3167;
															assign node3167 = (inp[0]) ? node3171 : node3168;
																assign node3168 = (inp[15]) ? 4'b0111 : 4'b0101;
																assign node3171 = (inp[15]) ? 4'b0101 : 4'b0111;
										assign node3175 = (inp[0]) ? node3221 : node3176;
											assign node3176 = (inp[9]) ? node3198 : node3177;
												assign node3177 = (inp[4]) ? node3189 : node3178;
													assign node3178 = (inp[15]) ? node3184 : node3179;
														assign node3179 = (inp[5]) ? node3181 : 4'b0110;
															assign node3181 = (inp[3]) ? 4'b0100 : 4'b0110;
														assign node3184 = (inp[5]) ? node3186 : 4'b0100;
															assign node3186 = (inp[3]) ? 4'b0110 : 4'b0100;
													assign node3189 = (inp[15]) ? node3193 : node3190;
														assign node3190 = (inp[3]) ? 4'b0000 : 4'b0010;
														assign node3193 = (inp[5]) ? node3195 : 4'b0000;
															assign node3195 = (inp[3]) ? 4'b0010 : 4'b0000;
												assign node3198 = (inp[4]) ? node3210 : node3199;
													assign node3199 = (inp[12]) ? node3205 : node3200;
														assign node3200 = (inp[5]) ? node3202 : 4'b0010;
															assign node3202 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node3205 = (inp[5]) ? 4'b0010 : node3206;
															assign node3206 = (inp[15]) ? 4'b0000 : 4'b0010;
													assign node3210 = (inp[15]) ? node3216 : node3211;
														assign node3211 = (inp[3]) ? 4'b0100 : node3212;
															assign node3212 = (inp[5]) ? 4'b0100 : 4'b0110;
														assign node3216 = (inp[5]) ? 4'b0110 : node3217;
															assign node3217 = (inp[3]) ? 4'b0110 : 4'b0100;
											assign node3221 = (inp[5]) ? node3237 : node3222;
												assign node3222 = (inp[15]) ? node3228 : node3223;
													assign node3223 = (inp[4]) ? 4'b0000 : node3224;
														assign node3224 = (inp[9]) ? 4'b0000 : 4'b0100;
													assign node3228 = (inp[3]) ? node3230 : 4'b0010;
														assign node3230 = (inp[9]) ? node3234 : node3231;
															assign node3231 = (inp[4]) ? 4'b0010 : 4'b0110;
															assign node3234 = (inp[4]) ? 4'b0100 : 4'b0010;
												assign node3237 = (inp[15]) ? node3251 : node3238;
													assign node3238 = (inp[3]) ? node3244 : node3239;
														assign node3239 = (inp[9]) ? node3241 : 4'b0000;
															assign node3241 = (inp[4]) ? 4'b0110 : 4'b0000;
														assign node3244 = (inp[4]) ? node3248 : node3245;
															assign node3245 = (inp[9]) ? 4'b0010 : 4'b0110;
															assign node3248 = (inp[9]) ? 4'b0110 : 4'b0010;
													assign node3251 = (inp[3]) ? node3259 : node3252;
														assign node3252 = (inp[4]) ? node3256 : node3253;
															assign node3253 = (inp[9]) ? 4'b0010 : 4'b0110;
															assign node3256 = (inp[9]) ? 4'b0100 : 4'b0010;
														assign node3259 = (inp[9]) ? 4'b0000 : node3260;
															assign node3260 = (inp[4]) ? 4'b0000 : 4'b0100;
									assign node3264 = (inp[3]) ? node3308 : node3265;
										assign node3265 = (inp[0]) ? node3285 : node3266;
											assign node3266 = (inp[15]) ? node3276 : node3267;
												assign node3267 = (inp[9]) ? node3271 : node3268;
													assign node3268 = (inp[4]) ? 4'b0010 : 4'b0110;
													assign node3271 = (inp[4]) ? node3273 : 4'b0010;
														assign node3273 = (inp[5]) ? 4'b0100 : 4'b0110;
												assign node3276 = (inp[4]) ? node3280 : node3277;
													assign node3277 = (inp[9]) ? 4'b0000 : 4'b0100;
													assign node3280 = (inp[9]) ? node3282 : 4'b0000;
														assign node3282 = (inp[5]) ? 4'b0110 : 4'b0100;
											assign node3285 = (inp[15]) ? node3299 : node3286;
												assign node3286 = (inp[5]) ? node3294 : node3287;
													assign node3287 = (inp[4]) ? node3291 : node3288;
														assign node3288 = (inp[9]) ? 4'b0000 : 4'b0100;
														assign node3291 = (inp[9]) ? 4'b0100 : 4'b0000;
													assign node3294 = (inp[4]) ? node3296 : 4'b0000;
														assign node3296 = (inp[9]) ? 4'b0110 : 4'b0000;
												assign node3299 = (inp[4]) ? node3303 : node3300;
													assign node3300 = (inp[9]) ? 4'b0010 : 4'b0110;
													assign node3303 = (inp[9]) ? node3305 : 4'b0010;
														assign node3305 = (inp[5]) ? 4'b0100 : 4'b0110;
										assign node3308 = (inp[12]) ? node3358 : node3309;
											assign node3309 = (inp[4]) ? node3337 : node3310;
												assign node3310 = (inp[9]) ? node3320 : node3311;
													assign node3311 = (inp[5]) ? node3313 : 4'b0110;
														assign node3313 = (inp[0]) ? node3317 : node3314;
															assign node3314 = (inp[15]) ? 4'b0110 : 4'b0100;
															assign node3317 = (inp[15]) ? 4'b0100 : 4'b0110;
													assign node3320 = (inp[5]) ? node3328 : node3321;
														assign node3321 = (inp[14]) ? node3323 : 4'b0010;
															assign node3323 = (inp[0]) ? 4'b0010 : node3324;
																assign node3324 = (inp[15]) ? 4'b0000 : 4'b0010;
														assign node3328 = (inp[14]) ? 4'b0010 : node3329;
															assign node3329 = (inp[15]) ? node3333 : node3330;
																assign node3330 = (inp[0]) ? 4'b0010 : 4'b0000;
																assign node3333 = (inp[0]) ? 4'b0000 : 4'b0010;
												assign node3337 = (inp[9]) ? node3351 : node3338;
													assign node3338 = (inp[0]) ? node3344 : node3339;
														assign node3339 = (inp[15]) ? 4'b0000 : node3340;
															assign node3340 = (inp[5]) ? 4'b0000 : 4'b0010;
														assign node3344 = (inp[14]) ? node3346 : 4'b0010;
															assign node3346 = (inp[15]) ? node3348 : 4'b0000;
																assign node3348 = (inp[5]) ? 4'b0000 : 4'b0010;
													assign node3351 = (inp[0]) ? node3355 : node3352;
														assign node3352 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node3355 = (inp[15]) ? 4'b0100 : 4'b0110;
											assign node3358 = (inp[4]) ? node3400 : node3359;
												assign node3359 = (inp[9]) ? node3389 : node3360;
													assign node3360 = (inp[15]) ? node3374 : node3361;
														assign node3361 = (inp[14]) ? node3369 : node3362;
															assign node3362 = (inp[5]) ? node3366 : node3363;
																assign node3363 = (inp[0]) ? 4'b0100 : 4'b0110;
																assign node3366 = (inp[0]) ? 4'b0110 : 4'b0100;
															assign node3369 = (inp[5]) ? node3371 : 4'b0100;
																assign node3371 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node3374 = (inp[14]) ? node3382 : node3375;
															assign node3375 = (inp[5]) ? node3379 : node3376;
																assign node3376 = (inp[0]) ? 4'b0110 : 4'b0100;
																assign node3379 = (inp[0]) ? 4'b0100 : 4'b0110;
															assign node3382 = (inp[0]) ? node3386 : node3383;
																assign node3383 = (inp[5]) ? 4'b0110 : 4'b0100;
																assign node3386 = (inp[5]) ? 4'b0100 : 4'b0110;
													assign node3389 = (inp[5]) ? node3395 : node3390;
														assign node3390 = (inp[0]) ? node3392 : 4'b0000;
															assign node3392 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node3395 = (inp[15]) ? node3397 : 4'b0010;
															assign node3397 = (inp[0]) ? 4'b0000 : 4'b0010;
												assign node3400 = (inp[9]) ? node3420 : node3401;
													assign node3401 = (inp[14]) ? node3409 : node3402;
														assign node3402 = (inp[15]) ? 4'b0000 : node3403;
															assign node3403 = (inp[5]) ? node3405 : 4'b0000;
																assign node3405 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node3409 = (inp[15]) ? node3415 : node3410;
															assign node3410 = (inp[5]) ? node3412 : 4'b0010;
																assign node3412 = (inp[0]) ? 4'b0010 : 4'b0000;
															assign node3415 = (inp[0]) ? 4'b0000 : node3416;
																assign node3416 = (inp[5]) ? 4'b0010 : 4'b0000;
													assign node3420 = (inp[15]) ? node3424 : node3421;
														assign node3421 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node3424 = (inp[0]) ? 4'b0100 : 4'b0110;
					assign node3427 = (inp[13]) ? node5115 : node3428;
						assign node3428 = (inp[8]) ? node4204 : node3429;
							assign node3429 = (inp[7]) ? node3873 : node3430;
								assign node3430 = (inp[14]) ? node3670 : node3431;
									assign node3431 = (inp[2]) ? node3533 : node3432;
										assign node3432 = (inp[5]) ? node3474 : node3433;
											assign node3433 = (inp[4]) ? node3459 : node3434;
												assign node3434 = (inp[9]) ? node3442 : node3435;
													assign node3435 = (inp[15]) ? node3439 : node3436;
														assign node3436 = (inp[0]) ? 4'b1101 : 4'b1111;
														assign node3439 = (inp[0]) ? 4'b1111 : 4'b1101;
													assign node3442 = (inp[12]) ? node3452 : node3443;
														assign node3443 = (inp[3]) ? 4'b1001 : node3444;
															assign node3444 = (inp[15]) ? node3448 : node3445;
																assign node3445 = (inp[0]) ? 4'b1001 : 4'b1011;
																assign node3448 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node3452 = (inp[0]) ? node3456 : node3453;
															assign node3453 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node3456 = (inp[15]) ? 4'b1011 : 4'b1001;
												assign node3459 = (inp[9]) ? node3465 : node3460;
													assign node3460 = (inp[0]) ? node3462 : 4'b1001;
														assign node3462 = (inp[15]) ? 4'b1011 : 4'b1001;
													assign node3465 = (inp[3]) ? node3467 : 4'b1101;
														assign node3467 = (inp[15]) ? node3471 : node3468;
															assign node3468 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node3471 = (inp[0]) ? 4'b1101 : 4'b1111;
											assign node3474 = (inp[0]) ? node3500 : node3475;
												assign node3475 = (inp[15]) ? node3489 : node3476;
													assign node3476 = (inp[3]) ? node3482 : node3477;
														assign node3477 = (inp[9]) ? node3479 : 4'b1011;
															assign node3479 = (inp[4]) ? 4'b1101 : 4'b1011;
														assign node3482 = (inp[12]) ? node3484 : 4'b1101;
															assign node3484 = (inp[9]) ? 4'b1001 : node3485;
																assign node3485 = (inp[4]) ? 4'b1001 : 4'b1101;
													assign node3489 = (inp[3]) ? node3495 : node3490;
														assign node3490 = (inp[4]) ? 4'b1111 : node3491;
															assign node3491 = (inp[9]) ? 4'b1001 : 4'b1101;
														assign node3495 = (inp[9]) ? 4'b1011 : node3496;
															assign node3496 = (inp[4]) ? 4'b1011 : 4'b1111;
												assign node3500 = (inp[15]) ? node3516 : node3501;
													assign node3501 = (inp[3]) ? node3509 : node3502;
														assign node3502 = (inp[9]) ? node3506 : node3503;
															assign node3503 = (inp[4]) ? 4'b1001 : 4'b1101;
															assign node3506 = (inp[4]) ? 4'b1111 : 4'b1001;
														assign node3509 = (inp[4]) ? node3513 : node3510;
															assign node3510 = (inp[9]) ? 4'b1011 : 4'b1111;
															assign node3513 = (inp[9]) ? 4'b1111 : 4'b1011;
													assign node3516 = (inp[3]) ? node3522 : node3517;
														assign node3517 = (inp[9]) ? 4'b1101 : node3518;
															assign node3518 = (inp[4]) ? 4'b1011 : 4'b1111;
														assign node3522 = (inp[12]) ? node3528 : node3523;
															assign node3523 = (inp[4]) ? 4'b1001 : node3524;
																assign node3524 = (inp[9]) ? 4'b1001 : 4'b1101;
															assign node3528 = (inp[4]) ? 4'b1101 : node3529;
																assign node3529 = (inp[9]) ? 4'b1001 : 4'b1101;
										assign node3533 = (inp[12]) ? node3609 : node3534;
											assign node3534 = (inp[0]) ? node3576 : node3535;
												assign node3535 = (inp[5]) ? node3557 : node3536;
													assign node3536 = (inp[15]) ? node3550 : node3537;
														assign node3537 = (inp[3]) ? node3543 : node3538;
															assign node3538 = (inp[4]) ? node3540 : 4'b1010;
																assign node3540 = (inp[9]) ? 4'b1110 : 4'b1010;
															assign node3543 = (inp[9]) ? node3547 : node3544;
																assign node3544 = (inp[4]) ? 4'b1010 : 4'b1110;
																assign node3547 = (inp[4]) ? 4'b1100 : 4'b1010;
														assign node3550 = (inp[9]) ? node3554 : node3551;
															assign node3551 = (inp[4]) ? 4'b1000 : 4'b1100;
															assign node3554 = (inp[4]) ? 4'b1110 : 4'b1000;
													assign node3557 = (inp[15]) ? node3567 : node3558;
														assign node3558 = (inp[3]) ? node3562 : node3559;
															assign node3559 = (inp[4]) ? 4'b1100 : 4'b1110;
															assign node3562 = (inp[9]) ? node3564 : 4'b1100;
																assign node3564 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node3567 = (inp[3]) ? node3571 : node3568;
															assign node3568 = (inp[4]) ? 4'b1000 : 4'b1100;
															assign node3571 = (inp[4]) ? node3573 : 4'b1110;
																assign node3573 = (inp[9]) ? 4'b1110 : 4'b1010;
												assign node3576 = (inp[15]) ? node3594 : node3577;
													assign node3577 = (inp[5]) ? node3583 : node3578;
														assign node3578 = (inp[4]) ? 4'b1000 : node3579;
															assign node3579 = (inp[9]) ? 4'b1000 : 4'b1100;
														assign node3583 = (inp[3]) ? node3591 : node3584;
															assign node3584 = (inp[9]) ? node3588 : node3585;
																assign node3585 = (inp[4]) ? 4'b1000 : 4'b1100;
																assign node3588 = (inp[4]) ? 4'b1110 : 4'b1000;
															assign node3591 = (inp[9]) ? 4'b1010 : 4'b1110;
													assign node3594 = (inp[3]) ? node3600 : node3595;
														assign node3595 = (inp[9]) ? node3597 : 4'b1010;
															assign node3597 = (inp[4]) ? 4'b1100 : 4'b1010;
														assign node3600 = (inp[4]) ? node3606 : node3601;
															assign node3601 = (inp[5]) ? 4'b1000 : node3602;
																assign node3602 = (inp[9]) ? 4'b1010 : 4'b1110;
															assign node3606 = (inp[9]) ? 4'b1100 : 4'b1000;
											assign node3609 = (inp[4]) ? node3641 : node3610;
												assign node3610 = (inp[9]) ? node3626 : node3611;
													assign node3611 = (inp[0]) ? node3619 : node3612;
														assign node3612 = (inp[15]) ? 4'b1100 : node3613;
															assign node3613 = (inp[5]) ? node3615 : 4'b1110;
																assign node3615 = (inp[3]) ? 4'b1100 : 4'b1110;
														assign node3619 = (inp[15]) ? 4'b1110 : node3620;
															assign node3620 = (inp[3]) ? node3622 : 4'b1100;
																assign node3622 = (inp[5]) ? 4'b1110 : 4'b1100;
													assign node3626 = (inp[5]) ? node3636 : node3627;
														assign node3627 = (inp[3]) ? 4'b1010 : node3628;
															assign node3628 = (inp[15]) ? node3632 : node3629;
																assign node3629 = (inp[0]) ? 4'b1000 : 4'b1010;
																assign node3632 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node3636 = (inp[3]) ? 4'b1000 : node3637;
															assign node3637 = (inp[0]) ? 4'b1000 : 4'b1010;
												assign node3641 = (inp[9]) ? node3655 : node3642;
													assign node3642 = (inp[15]) ? node3648 : node3643;
														assign node3643 = (inp[0]) ? node3645 : 4'b1010;
															assign node3645 = (inp[3]) ? 4'b1010 : 4'b1000;
														assign node3648 = (inp[3]) ? node3650 : 4'b1010;
															assign node3650 = (inp[0]) ? node3652 : 4'b1000;
																assign node3652 = (inp[5]) ? 4'b1000 : 4'b1010;
													assign node3655 = (inp[15]) ? node3661 : node3656;
														assign node3656 = (inp[0]) ? 4'b1110 : node3657;
															assign node3657 = (inp[3]) ? 4'b1100 : 4'b1110;
														assign node3661 = (inp[3]) ? node3667 : node3662;
															assign node3662 = (inp[5]) ? 4'b1100 : node3663;
																assign node3663 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node3667 = (inp[0]) ? 4'b1100 : 4'b1110;
									assign node3670 = (inp[2]) ? node3778 : node3671;
										assign node3671 = (inp[4]) ? node3715 : node3672;
											assign node3672 = (inp[9]) ? node3690 : node3673;
												assign node3673 = (inp[0]) ? node3681 : node3674;
													assign node3674 = (inp[15]) ? 4'b1100 : node3675;
														assign node3675 = (inp[3]) ? node3677 : 4'b1110;
															assign node3677 = (inp[5]) ? 4'b1100 : 4'b1110;
													assign node3681 = (inp[15]) ? node3687 : node3682;
														assign node3682 = (inp[3]) ? node3684 : 4'b1100;
															assign node3684 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node3687 = (inp[3]) ? 4'b1100 : 4'b1110;
												assign node3690 = (inp[3]) ? node3698 : node3691;
													assign node3691 = (inp[15]) ? node3695 : node3692;
														assign node3692 = (inp[0]) ? 4'b1000 : 4'b1010;
														assign node3695 = (inp[0]) ? 4'b1010 : 4'b1000;
													assign node3698 = (inp[0]) ? node3708 : node3699;
														assign node3699 = (inp[12]) ? node3701 : 4'b1010;
															assign node3701 = (inp[15]) ? node3705 : node3702;
																assign node3702 = (inp[5]) ? 4'b1000 : 4'b1010;
																assign node3705 = (inp[5]) ? 4'b1010 : 4'b1000;
														assign node3708 = (inp[5]) ? node3712 : node3709;
															assign node3709 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node3712 = (inp[15]) ? 4'b1000 : 4'b1010;
											assign node3715 = (inp[9]) ? node3747 : node3716;
												assign node3716 = (inp[12]) ? node3734 : node3717;
													assign node3717 = (inp[15]) ? node3727 : node3718;
														assign node3718 = (inp[0]) ? node3724 : node3719;
															assign node3719 = (inp[5]) ? node3721 : 4'b1010;
																assign node3721 = (inp[3]) ? 4'b1000 : 4'b1010;
															assign node3724 = (inp[5]) ? 4'b1010 : 4'b1000;
														assign node3727 = (inp[0]) ? node3729 : 4'b1000;
															assign node3729 = (inp[3]) ? node3731 : 4'b1010;
																assign node3731 = (inp[5]) ? 4'b1000 : 4'b1010;
													assign node3734 = (inp[0]) ? node3744 : node3735;
														assign node3735 = (inp[5]) ? node3739 : node3736;
															assign node3736 = (inp[15]) ? 4'b1000 : 4'b1010;
															assign node3739 = (inp[15]) ? 4'b1010 : node3740;
																assign node3740 = (inp[3]) ? 4'b1000 : 4'b1010;
														assign node3744 = (inp[15]) ? 4'b1010 : 4'b1000;
												assign node3747 = (inp[5]) ? node3763 : node3748;
													assign node3748 = (inp[15]) ? node3756 : node3749;
														assign node3749 = (inp[3]) ? node3753 : node3750;
															assign node3750 = (inp[0]) ? 4'b1100 : 4'b1110;
															assign node3753 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node3756 = (inp[0]) ? node3760 : node3757;
															assign node3757 = (inp[3]) ? 4'b1110 : 4'b1100;
															assign node3760 = (inp[3]) ? 4'b1100 : 4'b1110;
													assign node3763 = (inp[3]) ? node3771 : node3764;
														assign node3764 = (inp[15]) ? node3768 : node3765;
															assign node3765 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node3768 = (inp[0]) ? 4'b1100 : 4'b1110;
														assign node3771 = (inp[15]) ? node3775 : node3772;
															assign node3772 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node3775 = (inp[0]) ? 4'b1100 : 4'b1110;
										assign node3778 = (inp[5]) ? node3816 : node3779;
											assign node3779 = (inp[0]) ? node3797 : node3780;
												assign node3780 = (inp[15]) ? node3788 : node3781;
													assign node3781 = (inp[4]) ? node3785 : node3782;
														assign node3782 = (inp[9]) ? 4'b1010 : 4'b1110;
														assign node3785 = (inp[9]) ? 4'b1100 : 4'b1010;
													assign node3788 = (inp[3]) ? node3790 : 4'b1000;
														assign node3790 = (inp[9]) ? node3794 : node3791;
															assign node3791 = (inp[4]) ? 4'b1000 : 4'b1100;
															assign node3794 = (inp[4]) ? 4'b1110 : 4'b1000;
												assign node3797 = (inp[15]) ? node3807 : node3798;
													assign node3798 = (inp[9]) ? node3802 : node3799;
														assign node3799 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node3802 = (inp[4]) ? node3804 : 4'b1000;
															assign node3804 = (inp[3]) ? 4'b1110 : 4'b1100;
													assign node3807 = (inp[9]) ? node3811 : node3808;
														assign node3808 = (inp[4]) ? 4'b1010 : 4'b1110;
														assign node3811 = (inp[4]) ? node3813 : 4'b1010;
															assign node3813 = (inp[3]) ? 4'b1100 : 4'b1110;
											assign node3816 = (inp[0]) ? node3844 : node3817;
												assign node3817 = (inp[15]) ? node3829 : node3818;
													assign node3818 = (inp[3]) ? node3824 : node3819;
														assign node3819 = (inp[9]) ? 4'b1010 : node3820;
															assign node3820 = (inp[4]) ? 4'b1010 : 4'b1110;
														assign node3824 = (inp[9]) ? node3826 : 4'b1000;
															assign node3826 = (inp[4]) ? 4'b1100 : 4'b1000;
													assign node3829 = (inp[3]) ? node3835 : node3830;
														assign node3830 = (inp[9]) ? 4'b1110 : node3831;
															assign node3831 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node3835 = (inp[12]) ? node3837 : 4'b1110;
															assign node3837 = (inp[4]) ? node3841 : node3838;
																assign node3838 = (inp[9]) ? 4'b1010 : 4'b1110;
																assign node3841 = (inp[9]) ? 4'b1110 : 4'b1010;
												assign node3844 = (inp[12]) ? node3856 : node3845;
													assign node3845 = (inp[4]) ? node3853 : node3846;
														assign node3846 = (inp[9]) ? node3848 : 4'b1110;
															assign node3848 = (inp[15]) ? 4'b1010 : node3849;
																assign node3849 = (inp[3]) ? 4'b1010 : 4'b1000;
														assign node3853 = (inp[9]) ? 4'b1110 : 4'b1010;
													assign node3856 = (inp[3]) ? node3864 : node3857;
														assign node3857 = (inp[15]) ? node3859 : 4'b1000;
															assign node3859 = (inp[9]) ? 4'b1010 : node3860;
																assign node3860 = (inp[4]) ? 4'b1010 : 4'b1110;
														assign node3864 = (inp[15]) ? node3870 : node3865;
															assign node3865 = (inp[9]) ? node3867 : 4'b1110;
																assign node3867 = (inp[4]) ? 4'b1110 : 4'b1010;
															assign node3870 = (inp[4]) ? 4'b1000 : 4'b1100;
								assign node3873 = (inp[2]) ? node4103 : node3874;
									assign node3874 = (inp[14]) ? node3980 : node3875;
										assign node3875 = (inp[0]) ? node3921 : node3876;
											assign node3876 = (inp[15]) ? node3898 : node3877;
												assign node3877 = (inp[5]) ? node3887 : node3878;
													assign node3878 = (inp[4]) ? node3882 : node3879;
														assign node3879 = (inp[9]) ? 4'b1010 : 4'b1110;
														assign node3882 = (inp[9]) ? node3884 : 4'b1010;
															assign node3884 = (inp[3]) ? 4'b1100 : 4'b1110;
													assign node3887 = (inp[3]) ? node3893 : node3888;
														assign node3888 = (inp[9]) ? node3890 : 4'b1010;
															assign node3890 = (inp[4]) ? 4'b1100 : 4'b1010;
														assign node3893 = (inp[4]) ? node3895 : 4'b1000;
															assign node3895 = (inp[9]) ? 4'b1100 : 4'b1000;
												assign node3898 = (inp[5]) ? node3906 : node3899;
													assign node3899 = (inp[4]) ? node3903 : node3900;
														assign node3900 = (inp[9]) ? 4'b1000 : 4'b1100;
														assign node3903 = (inp[9]) ? 4'b1110 : 4'b1000;
													assign node3906 = (inp[3]) ? node3914 : node3907;
														assign node3907 = (inp[4]) ? node3911 : node3908;
															assign node3908 = (inp[9]) ? 4'b1000 : 4'b1100;
															assign node3911 = (inp[9]) ? 4'b1110 : 4'b1000;
														assign node3914 = (inp[4]) ? node3918 : node3915;
															assign node3915 = (inp[9]) ? 4'b1010 : 4'b1110;
															assign node3918 = (inp[9]) ? 4'b1110 : 4'b1010;
											assign node3921 = (inp[15]) ? node3957 : node3922;
												assign node3922 = (inp[3]) ? node3944 : node3923;
													assign node3923 = (inp[5]) ? node3937 : node3924;
														assign node3924 = (inp[12]) ? node3932 : node3925;
															assign node3925 = (inp[4]) ? node3929 : node3926;
																assign node3926 = (inp[9]) ? 4'b1000 : 4'b1100;
																assign node3929 = (inp[9]) ? 4'b1100 : 4'b1000;
															assign node3932 = (inp[9]) ? 4'b1100 : node3933;
																assign node3933 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node3937 = (inp[4]) ? node3941 : node3938;
															assign node3938 = (inp[9]) ? 4'b1000 : 4'b1100;
															assign node3941 = (inp[12]) ? 4'b1000 : 4'b1110;
													assign node3944 = (inp[5]) ? node3952 : node3945;
														assign node3945 = (inp[9]) ? node3949 : node3946;
															assign node3946 = (inp[4]) ? 4'b1000 : 4'b1100;
															assign node3949 = (inp[4]) ? 4'b1110 : 4'b1000;
														assign node3952 = (inp[9]) ? 4'b1010 : node3953;
															assign node3953 = (inp[4]) ? 4'b1010 : 4'b1110;
												assign node3957 = (inp[3]) ? node3967 : node3958;
													assign node3958 = (inp[4]) ? node3962 : node3959;
														assign node3959 = (inp[9]) ? 4'b1010 : 4'b1110;
														assign node3962 = (inp[9]) ? node3964 : 4'b1010;
															assign node3964 = (inp[5]) ? 4'b1100 : 4'b1110;
													assign node3967 = (inp[5]) ? node3973 : node3968;
														assign node3968 = (inp[4]) ? node3970 : 4'b1010;
															assign node3970 = (inp[9]) ? 4'b1100 : 4'b1010;
														assign node3973 = (inp[9]) ? node3977 : node3974;
															assign node3974 = (inp[4]) ? 4'b1000 : 4'b1100;
															assign node3977 = (inp[4]) ? 4'b1100 : 4'b1000;
										assign node3980 = (inp[12]) ? node4040 : node3981;
											assign node3981 = (inp[15]) ? node4011 : node3982;
												assign node3982 = (inp[0]) ? node3994 : node3983;
													assign node3983 = (inp[3]) ? node3987 : node3984;
														assign node3984 = (inp[9]) ? 4'b0011 : 4'b0111;
														assign node3987 = (inp[5]) ? node3989 : 4'b0011;
															assign node3989 = (inp[4]) ? node3991 : 4'b0001;
																assign node3991 = (inp[9]) ? 4'b0101 : 4'b0001;
													assign node3994 = (inp[3]) ? node4004 : node3995;
														assign node3995 = (inp[5]) ? node4001 : node3996;
															assign node3996 = (inp[9]) ? 4'b0101 : node3997;
																assign node3997 = (inp[4]) ? 4'b0001 : 4'b0101;
															assign node4001 = (inp[9]) ? 4'b0001 : 4'b0101;
														assign node4004 = (inp[5]) ? node4006 : 4'b0001;
															assign node4006 = (inp[4]) ? 4'b0111 : node4007;
																assign node4007 = (inp[9]) ? 4'b0011 : 4'b0111;
												assign node4011 = (inp[5]) ? node4025 : node4012;
													assign node4012 = (inp[0]) ? node4018 : node4013;
														assign node4013 = (inp[4]) ? node4015 : 4'b0101;
															assign node4015 = (inp[3]) ? 4'b0111 : 4'b0101;
														assign node4018 = (inp[9]) ? node4022 : node4019;
															assign node4019 = (inp[4]) ? 4'b0011 : 4'b0111;
															assign node4022 = (inp[4]) ? 4'b0101 : 4'b0011;
													assign node4025 = (inp[9]) ? node4035 : node4026;
														assign node4026 = (inp[4]) ? node4028 : 4'b0111;
															assign node4028 = (inp[0]) ? node4032 : node4029;
																assign node4029 = (inp[3]) ? 4'b0011 : 4'b0001;
																assign node4032 = (inp[3]) ? 4'b0001 : 4'b0011;
														assign node4035 = (inp[0]) ? 4'b0101 : node4036;
															assign node4036 = (inp[4]) ? 4'b0111 : 4'b0011;
											assign node4040 = (inp[9]) ? node4066 : node4041;
												assign node4041 = (inp[4]) ? node4055 : node4042;
													assign node4042 = (inp[15]) ? node4048 : node4043;
														assign node4043 = (inp[0]) ? 4'b0101 : node4044;
															assign node4044 = (inp[3]) ? 4'b0101 : 4'b0111;
														assign node4048 = (inp[5]) ? node4052 : node4049;
															assign node4049 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node4052 = (inp[0]) ? 4'b0101 : 4'b0111;
													assign node4055 = (inp[15]) ? node4057 : 4'b0001;
														assign node4057 = (inp[0]) ? node4063 : node4058;
															assign node4058 = (inp[3]) ? node4060 : 4'b0001;
																assign node4060 = (inp[5]) ? 4'b0011 : 4'b0001;
															assign node4063 = (inp[5]) ? 4'b0001 : 4'b0011;
												assign node4066 = (inp[4]) ? node4086 : node4067;
													assign node4067 = (inp[15]) ? node4079 : node4068;
														assign node4068 = (inp[0]) ? node4074 : node4069;
															assign node4069 = (inp[3]) ? node4071 : 4'b0011;
																assign node4071 = (inp[5]) ? 4'b0001 : 4'b0011;
															assign node4074 = (inp[3]) ? node4076 : 4'b0001;
																assign node4076 = (inp[5]) ? 4'b0011 : 4'b0001;
														assign node4079 = (inp[0]) ? node4081 : 4'b0001;
															assign node4081 = (inp[5]) ? node4083 : 4'b0011;
																assign node4083 = (inp[3]) ? 4'b0001 : 4'b0011;
													assign node4086 = (inp[3]) ? node4096 : node4087;
														assign node4087 = (inp[15]) ? node4089 : 4'b0111;
															assign node4089 = (inp[5]) ? node4093 : node4090;
																assign node4090 = (inp[0]) ? 4'b0111 : 4'b0101;
																assign node4093 = (inp[0]) ? 4'b0101 : 4'b0111;
														assign node4096 = (inp[15]) ? node4100 : node4097;
															assign node4097 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node4100 = (inp[0]) ? 4'b0101 : 4'b0111;
									assign node4103 = (inp[4]) ? node4157 : node4104;
										assign node4104 = (inp[9]) ? node4128 : node4105;
											assign node4105 = (inp[15]) ? node4117 : node4106;
												assign node4106 = (inp[0]) ? node4112 : node4107;
													assign node4107 = (inp[5]) ? node4109 : 4'b0111;
														assign node4109 = (inp[3]) ? 4'b0101 : 4'b0111;
													assign node4112 = (inp[3]) ? node4114 : 4'b0101;
														assign node4114 = (inp[5]) ? 4'b0111 : 4'b0101;
												assign node4117 = (inp[0]) ? node4123 : node4118;
													assign node4118 = (inp[5]) ? node4120 : 4'b0101;
														assign node4120 = (inp[3]) ? 4'b0111 : 4'b0101;
													assign node4123 = (inp[3]) ? node4125 : 4'b0111;
														assign node4125 = (inp[12]) ? 4'b0111 : 4'b0101;
											assign node4128 = (inp[12]) ? node4140 : node4129;
												assign node4129 = (inp[0]) ? node4131 : 4'b0011;
													assign node4131 = (inp[15]) ? node4135 : node4132;
														assign node4132 = (inp[3]) ? 4'b0011 : 4'b0001;
														assign node4135 = (inp[5]) ? node4137 : 4'b0011;
															assign node4137 = (inp[3]) ? 4'b0001 : 4'b0011;
												assign node4140 = (inp[15]) ? node4148 : node4141;
													assign node4141 = (inp[0]) ? node4143 : 4'b0011;
														assign node4143 = (inp[3]) ? node4145 : 4'b0001;
															assign node4145 = (inp[5]) ? 4'b0011 : 4'b0001;
													assign node4148 = (inp[0]) ? node4152 : node4149;
														assign node4149 = (inp[5]) ? 4'b0011 : 4'b0001;
														assign node4152 = (inp[5]) ? node4154 : 4'b0011;
															assign node4154 = (inp[3]) ? 4'b0001 : 4'b0011;
										assign node4157 = (inp[9]) ? node4181 : node4158;
											assign node4158 = (inp[15]) ? node4170 : node4159;
												assign node4159 = (inp[0]) ? node4165 : node4160;
													assign node4160 = (inp[5]) ? node4162 : 4'b0011;
														assign node4162 = (inp[3]) ? 4'b0001 : 4'b0011;
													assign node4165 = (inp[3]) ? node4167 : 4'b0001;
														assign node4167 = (inp[5]) ? 4'b0011 : 4'b0001;
												assign node4170 = (inp[0]) ? node4176 : node4171;
													assign node4171 = (inp[5]) ? node4173 : 4'b0001;
														assign node4173 = (inp[3]) ? 4'b0011 : 4'b0001;
													assign node4176 = (inp[5]) ? node4178 : 4'b0011;
														assign node4178 = (inp[3]) ? 4'b0001 : 4'b0011;
											assign node4181 = (inp[15]) ? node4193 : node4182;
												assign node4182 = (inp[0]) ? node4188 : node4183;
													assign node4183 = (inp[5]) ? 4'b0101 : node4184;
														assign node4184 = (inp[3]) ? 4'b0101 : 4'b0111;
													assign node4188 = (inp[3]) ? 4'b0111 : node4189;
														assign node4189 = (inp[5]) ? 4'b0111 : 4'b0101;
												assign node4193 = (inp[0]) ? node4199 : node4194;
													assign node4194 = (inp[5]) ? 4'b0111 : node4195;
														assign node4195 = (inp[3]) ? 4'b0111 : 4'b0101;
													assign node4199 = (inp[5]) ? 4'b0101 : node4200;
														assign node4200 = (inp[3]) ? 4'b0101 : 4'b0111;
							assign node4204 = (inp[7]) ? node4750 : node4205;
								assign node4205 = (inp[14]) ? node4473 : node4206;
									assign node4206 = (inp[2]) ? node4348 : node4207;
										assign node4207 = (inp[5]) ? node4275 : node4208;
											assign node4208 = (inp[12]) ? node4242 : node4209;
												assign node4209 = (inp[4]) ? node4223 : node4210;
													assign node4210 = (inp[9]) ? node4216 : node4211;
														assign node4211 = (inp[0]) ? 4'b1110 : node4212;
															assign node4212 = (inp[15]) ? 4'b1100 : 4'b1110;
														assign node4216 = (inp[0]) ? node4220 : node4217;
															assign node4217 = (inp[15]) ? 4'b1000 : 4'b1010;
															assign node4220 = (inp[15]) ? 4'b1010 : 4'b1000;
													assign node4223 = (inp[9]) ? node4231 : node4224;
														assign node4224 = (inp[3]) ? 4'b1010 : node4225;
															assign node4225 = (inp[0]) ? 4'b1000 : node4226;
																assign node4226 = (inp[15]) ? 4'b1000 : 4'b1010;
														assign node4231 = (inp[3]) ? node4237 : node4232;
															assign node4232 = (inp[0]) ? node4234 : 4'b1110;
																assign node4234 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node4237 = (inp[0]) ? node4239 : 4'b1100;
																assign node4239 = (inp[15]) ? 4'b1100 : 4'b1110;
												assign node4242 = (inp[9]) ? node4254 : node4243;
													assign node4243 = (inp[4]) ? node4249 : node4244;
														assign node4244 = (inp[0]) ? node4246 : 4'b1100;
															assign node4246 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node4249 = (inp[0]) ? node4251 : 4'b1010;
															assign node4251 = (inp[15]) ? 4'b1010 : 4'b1000;
													assign node4254 = (inp[4]) ? node4260 : node4255;
														assign node4255 = (inp[15]) ? node4257 : 4'b1010;
															assign node4257 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node4260 = (inp[15]) ? node4268 : node4261;
															assign node4261 = (inp[3]) ? node4265 : node4262;
																assign node4262 = (inp[0]) ? 4'b1100 : 4'b1110;
																assign node4265 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node4268 = (inp[0]) ? node4272 : node4269;
																assign node4269 = (inp[3]) ? 4'b1110 : 4'b1100;
																assign node4272 = (inp[3]) ? 4'b1100 : 4'b1110;
											assign node4275 = (inp[12]) ? node4315 : node4276;
												assign node4276 = (inp[9]) ? node4300 : node4277;
													assign node4277 = (inp[4]) ? node4285 : node4278;
														assign node4278 = (inp[15]) ? 4'b1100 : node4279;
															assign node4279 = (inp[3]) ? 4'b1110 : node4280;
																assign node4280 = (inp[0]) ? 4'b1100 : 4'b1110;
														assign node4285 = (inp[15]) ? node4293 : node4286;
															assign node4286 = (inp[3]) ? node4290 : node4287;
																assign node4287 = (inp[0]) ? 4'b1000 : 4'b1010;
																assign node4290 = (inp[0]) ? 4'b1010 : 4'b1000;
															assign node4293 = (inp[0]) ? node4297 : node4294;
																assign node4294 = (inp[3]) ? 4'b1010 : 4'b1000;
																assign node4297 = (inp[3]) ? 4'b1000 : 4'b1010;
													assign node4300 = (inp[4]) ? node4310 : node4301;
														assign node4301 = (inp[3]) ? 4'b1000 : node4302;
															assign node4302 = (inp[0]) ? node4306 : node4303;
																assign node4303 = (inp[15]) ? 4'b1000 : 4'b1010;
																assign node4306 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node4310 = (inp[15]) ? node4312 : 4'b1110;
															assign node4312 = (inp[0]) ? 4'b1100 : 4'b1110;
												assign node4315 = (inp[3]) ? node4335 : node4316;
													assign node4316 = (inp[9]) ? node4320 : node4317;
														assign node4317 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node4320 = (inp[4]) ? node4328 : node4321;
															assign node4321 = (inp[0]) ? node4325 : node4322;
																assign node4322 = (inp[15]) ? 4'b1000 : 4'b1010;
																assign node4325 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node4328 = (inp[15]) ? node4332 : node4329;
																assign node4329 = (inp[0]) ? 4'b1110 : 4'b1100;
																assign node4332 = (inp[0]) ? 4'b1100 : 4'b1110;
													assign node4335 = (inp[15]) ? node4339 : node4336;
														assign node4336 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node4339 = (inp[0]) ? node4343 : node4340;
															assign node4340 = (inp[9]) ? 4'b1010 : 4'b1110;
															assign node4343 = (inp[4]) ? node4345 : 4'b1000;
																assign node4345 = (inp[9]) ? 4'b1100 : 4'b1000;
										assign node4348 = (inp[5]) ? node4404 : node4349;
											assign node4349 = (inp[9]) ? node4379 : node4350;
												assign node4350 = (inp[4]) ? node4366 : node4351;
													assign node4351 = (inp[3]) ? node4359 : node4352;
														assign node4352 = (inp[15]) ? node4356 : node4353;
															assign node4353 = (inp[0]) ? 4'b0101 : 4'b0111;
															assign node4356 = (inp[0]) ? 4'b0111 : 4'b0101;
														assign node4359 = (inp[0]) ? node4363 : node4360;
															assign node4360 = (inp[15]) ? 4'b0101 : 4'b0111;
															assign node4363 = (inp[15]) ? 4'b0111 : 4'b0101;
													assign node4366 = (inp[12]) ? node4372 : node4367;
														assign node4367 = (inp[3]) ? 4'b0011 : node4368;
															assign node4368 = (inp[0]) ? 4'b0001 : 4'b0011;
														assign node4372 = (inp[0]) ? node4376 : node4373;
															assign node4373 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node4376 = (inp[15]) ? 4'b0011 : 4'b0001;
												assign node4379 = (inp[4]) ? node4395 : node4380;
													assign node4380 = (inp[12]) ? node4388 : node4381;
														assign node4381 = (inp[3]) ? node4383 : 4'b0001;
															assign node4383 = (inp[15]) ? 4'b0001 : node4384;
																assign node4384 = (inp[0]) ? 4'b0001 : 4'b0011;
														assign node4388 = (inp[15]) ? node4392 : node4389;
															assign node4389 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node4392 = (inp[0]) ? 4'b0011 : 4'b0001;
													assign node4395 = (inp[3]) ? node4397 : 4'b0101;
														assign node4397 = (inp[12]) ? 4'b0111 : node4398;
															assign node4398 = (inp[15]) ? 4'b0101 : node4399;
																assign node4399 = (inp[0]) ? 4'b0111 : 4'b0101;
											assign node4404 = (inp[3]) ? node4428 : node4405;
												assign node4405 = (inp[0]) ? node4419 : node4406;
													assign node4406 = (inp[15]) ? node4414 : node4407;
														assign node4407 = (inp[9]) ? node4411 : node4408;
															assign node4408 = (inp[4]) ? 4'b0011 : 4'b0111;
															assign node4411 = (inp[4]) ? 4'b0101 : 4'b0011;
														assign node4414 = (inp[9]) ? 4'b0111 : node4415;
															assign node4415 = (inp[4]) ? 4'b0001 : 4'b0101;
													assign node4419 = (inp[15]) ? node4423 : node4420;
														assign node4420 = (inp[4]) ? 4'b0111 : 4'b0001;
														assign node4423 = (inp[9]) ? 4'b0011 : node4424;
															assign node4424 = (inp[4]) ? 4'b0011 : 4'b0111;
												assign node4428 = (inp[12]) ? node4454 : node4429;
													assign node4429 = (inp[9]) ? node4441 : node4430;
														assign node4430 = (inp[4]) ? node4436 : node4431;
															assign node4431 = (inp[15]) ? 4'b0101 : node4432;
																assign node4432 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node4436 = (inp[15]) ? node4438 : 4'b0001;
																assign node4438 = (inp[0]) ? 4'b0001 : 4'b0011;
														assign node4441 = (inp[4]) ? node4449 : node4442;
															assign node4442 = (inp[0]) ? node4446 : node4443;
																assign node4443 = (inp[15]) ? 4'b0011 : 4'b0001;
																assign node4446 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node4449 = (inp[0]) ? 4'b0101 : node4450;
																assign node4450 = (inp[15]) ? 4'b0111 : 4'b0101;
													assign node4454 = (inp[9]) ? node4464 : node4455;
														assign node4455 = (inp[4]) ? node4459 : node4456;
															assign node4456 = (inp[15]) ? 4'b0111 : 4'b0101;
															assign node4459 = (inp[15]) ? 4'b0011 : node4460;
																assign node4460 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node4464 = (inp[4]) ? node4468 : node4465;
															assign node4465 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node4468 = (inp[0]) ? node4470 : 4'b0111;
																assign node4470 = (inp[15]) ? 4'b0101 : 4'b0111;
									assign node4473 = (inp[12]) ? node4603 : node4474;
										assign node4474 = (inp[4]) ? node4550 : node4475;
											assign node4475 = (inp[9]) ? node4501 : node4476;
												assign node4476 = (inp[5]) ? node4492 : node4477;
													assign node4477 = (inp[2]) ? node4485 : node4478;
														assign node4478 = (inp[0]) ? node4482 : node4479;
															assign node4479 = (inp[15]) ? 4'b0101 : 4'b0111;
															assign node4482 = (inp[15]) ? 4'b0111 : 4'b0101;
														assign node4485 = (inp[0]) ? node4489 : node4486;
															assign node4486 = (inp[15]) ? 4'b0101 : 4'b0111;
															assign node4489 = (inp[15]) ? 4'b0111 : 4'b0101;
													assign node4492 = (inp[0]) ? 4'b0101 : node4493;
														assign node4493 = (inp[15]) ? node4497 : node4494;
															assign node4494 = (inp[3]) ? 4'b0101 : 4'b0111;
															assign node4497 = (inp[3]) ? 4'b0111 : 4'b0101;
												assign node4501 = (inp[3]) ? node4521 : node4502;
													assign node4502 = (inp[2]) ? node4514 : node4503;
														assign node4503 = (inp[5]) ? node4509 : node4504;
															assign node4504 = (inp[0]) ? 4'b0001 : node4505;
																assign node4505 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node4509 = (inp[0]) ? node4511 : 4'b0001;
																assign node4511 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node4514 = (inp[15]) ? node4518 : node4515;
															assign node4515 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node4518 = (inp[0]) ? 4'b0011 : 4'b0001;
													assign node4521 = (inp[2]) ? node4535 : node4522;
														assign node4522 = (inp[5]) ? node4528 : node4523;
															assign node4523 = (inp[0]) ? 4'b0011 : node4524;
																assign node4524 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node4528 = (inp[0]) ? node4532 : node4529;
																assign node4529 = (inp[15]) ? 4'b0011 : 4'b0001;
																assign node4532 = (inp[15]) ? 4'b0001 : 4'b0011;
														assign node4535 = (inp[15]) ? node4543 : node4536;
															assign node4536 = (inp[5]) ? node4540 : node4537;
																assign node4537 = (inp[0]) ? 4'b0001 : 4'b0011;
																assign node4540 = (inp[0]) ? 4'b0011 : 4'b0001;
															assign node4543 = (inp[5]) ? node4547 : node4544;
																assign node4544 = (inp[0]) ? 4'b0011 : 4'b0001;
																assign node4547 = (inp[0]) ? 4'b0001 : 4'b0011;
											assign node4550 = (inp[9]) ? node4584 : node4551;
												assign node4551 = (inp[2]) ? node4571 : node4552;
													assign node4552 = (inp[15]) ? node4560 : node4553;
														assign node4553 = (inp[0]) ? 4'b0001 : node4554;
															assign node4554 = (inp[3]) ? node4556 : 4'b0011;
																assign node4556 = (inp[5]) ? 4'b0001 : 4'b0011;
														assign node4560 = (inp[0]) ? node4566 : node4561;
															assign node4561 = (inp[3]) ? node4563 : 4'b0001;
																assign node4563 = (inp[5]) ? 4'b0011 : 4'b0001;
															assign node4566 = (inp[5]) ? node4568 : 4'b0011;
																assign node4568 = (inp[3]) ? 4'b0001 : 4'b0011;
													assign node4571 = (inp[5]) ? node4577 : node4572;
														assign node4572 = (inp[3]) ? 4'b0001 : node4573;
															assign node4573 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node4577 = (inp[0]) ? 4'b0011 : node4578;
															assign node4578 = (inp[15]) ? node4580 : 4'b0011;
																assign node4580 = (inp[3]) ? 4'b0011 : 4'b0001;
												assign node4584 = (inp[15]) ? node4592 : node4585;
													assign node4585 = (inp[0]) ? 4'b0111 : node4586;
														assign node4586 = (inp[5]) ? 4'b0101 : node4587;
															assign node4587 = (inp[3]) ? 4'b0101 : 4'b0111;
													assign node4592 = (inp[0]) ? node4598 : node4593;
														assign node4593 = (inp[3]) ? 4'b0111 : node4594;
															assign node4594 = (inp[5]) ? 4'b0111 : 4'b0101;
														assign node4598 = (inp[3]) ? 4'b0101 : node4599;
															assign node4599 = (inp[5]) ? 4'b0101 : 4'b0111;
										assign node4603 = (inp[2]) ? node4687 : node4604;
											assign node4604 = (inp[3]) ? node4646 : node4605;
												assign node4605 = (inp[4]) ? node4627 : node4606;
													assign node4606 = (inp[9]) ? node4620 : node4607;
														assign node4607 = (inp[5]) ? node4613 : node4608;
															assign node4608 = (inp[15]) ? node4610 : 4'b0101;
																assign node4610 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node4613 = (inp[15]) ? node4617 : node4614;
																assign node4614 = (inp[0]) ? 4'b0101 : 4'b0111;
																assign node4617 = (inp[0]) ? 4'b0111 : 4'b0101;
														assign node4620 = (inp[15]) ? node4624 : node4621;
															assign node4621 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node4624 = (inp[0]) ? 4'b0011 : 4'b0001;
													assign node4627 = (inp[9]) ? node4637 : node4628;
														assign node4628 = (inp[5]) ? node4630 : 4'b0011;
															assign node4630 = (inp[15]) ? node4634 : node4631;
																assign node4631 = (inp[0]) ? 4'b0001 : 4'b0011;
																assign node4634 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node4637 = (inp[5]) ? 4'b0111 : node4638;
															assign node4638 = (inp[0]) ? node4642 : node4639;
																assign node4639 = (inp[15]) ? 4'b0101 : 4'b0111;
																assign node4642 = (inp[15]) ? 4'b0111 : 4'b0101;
												assign node4646 = (inp[5]) ? node4670 : node4647;
													assign node4647 = (inp[4]) ? node4657 : node4648;
														assign node4648 = (inp[9]) ? 4'b0011 : node4649;
															assign node4649 = (inp[0]) ? node4653 : node4650;
																assign node4650 = (inp[15]) ? 4'b0101 : 4'b0111;
																assign node4653 = (inp[15]) ? 4'b0111 : 4'b0101;
														assign node4657 = (inp[9]) ? node4663 : node4658;
															assign node4658 = (inp[0]) ? 4'b0011 : node4659;
																assign node4659 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node4663 = (inp[15]) ? node4667 : node4664;
																assign node4664 = (inp[0]) ? 4'b0111 : 4'b0101;
																assign node4667 = (inp[0]) ? 4'b0101 : 4'b0111;
													assign node4670 = (inp[15]) ? node4678 : node4671;
														assign node4671 = (inp[0]) ? node4673 : 4'b0101;
															assign node4673 = (inp[9]) ? node4675 : 4'b0011;
																assign node4675 = (inp[4]) ? 4'b0111 : 4'b0011;
														assign node4678 = (inp[0]) ? 4'b0101 : node4679;
															assign node4679 = (inp[9]) ? node4683 : node4680;
																assign node4680 = (inp[4]) ? 4'b0011 : 4'b0111;
																assign node4683 = (inp[4]) ? 4'b0111 : 4'b0011;
											assign node4687 = (inp[15]) ? node4719 : node4688;
												assign node4688 = (inp[0]) ? node4702 : node4689;
													assign node4689 = (inp[3]) ? node4693 : node4690;
														assign node4690 = (inp[5]) ? 4'b0011 : 4'b0111;
														assign node4693 = (inp[5]) ? node4695 : 4'b0011;
															assign node4695 = (inp[4]) ? node4699 : node4696;
																assign node4696 = (inp[9]) ? 4'b0001 : 4'b0101;
																assign node4699 = (inp[9]) ? 4'b0101 : 4'b0001;
													assign node4702 = (inp[5]) ? node4712 : node4703;
														assign node4703 = (inp[4]) ? node4707 : node4704;
															assign node4704 = (inp[9]) ? 4'b0001 : 4'b0101;
															assign node4707 = (inp[9]) ? node4709 : 4'b0001;
																assign node4709 = (inp[3]) ? 4'b0111 : 4'b0101;
														assign node4712 = (inp[3]) ? 4'b0111 : node4713;
															assign node4713 = (inp[4]) ? node4715 : 4'b0001;
																assign node4715 = (inp[9]) ? 4'b0111 : 4'b0001;
												assign node4719 = (inp[0]) ? node4737 : node4720;
													assign node4720 = (inp[3]) ? node4726 : node4721;
														assign node4721 = (inp[4]) ? node4723 : 4'b0101;
															assign node4723 = (inp[5]) ? 4'b0001 : 4'b0101;
														assign node4726 = (inp[5]) ? node4730 : node4727;
															assign node4727 = (inp[9]) ? 4'b0001 : 4'b0101;
															assign node4730 = (inp[9]) ? node4734 : node4731;
																assign node4731 = (inp[4]) ? 4'b0011 : 4'b0111;
																assign node4734 = (inp[4]) ? 4'b0111 : 4'b0011;
													assign node4737 = (inp[5]) ? node4745 : node4738;
														assign node4738 = (inp[9]) ? node4742 : node4739;
															assign node4739 = (inp[4]) ? 4'b0011 : 4'b0111;
															assign node4742 = (inp[4]) ? 4'b0111 : 4'b0011;
														assign node4745 = (inp[4]) ? 4'b0101 : node4746;
															assign node4746 = (inp[9]) ? 4'b0011 : 4'b0111;
								assign node4750 = (inp[14]) ? node4966 : node4751;
									assign node4751 = (inp[2]) ? node4889 : node4752;
										assign node4752 = (inp[9]) ? node4820 : node4753;
											assign node4753 = (inp[4]) ? node4789 : node4754;
												assign node4754 = (inp[3]) ? node4770 : node4755;
													assign node4755 = (inp[5]) ? node4763 : node4756;
														assign node4756 = (inp[12]) ? 4'b0101 : node4757;
															assign node4757 = (inp[15]) ? node4759 : 4'b0101;
																assign node4759 = (inp[0]) ? 4'b0111 : 4'b0101;
														assign node4763 = (inp[0]) ? node4767 : node4764;
															assign node4764 = (inp[15]) ? 4'b0101 : 4'b0111;
															assign node4767 = (inp[15]) ? 4'b0111 : 4'b0101;
													assign node4770 = (inp[12]) ? node4780 : node4771;
														assign node4771 = (inp[0]) ? node4773 : 4'b0111;
															assign node4773 = (inp[5]) ? node4777 : node4774;
																assign node4774 = (inp[15]) ? 4'b0111 : 4'b0101;
																assign node4777 = (inp[15]) ? 4'b0101 : 4'b0111;
														assign node4780 = (inp[0]) ? node4782 : 4'b0101;
															assign node4782 = (inp[15]) ? node4786 : node4783;
																assign node4783 = (inp[5]) ? 4'b0111 : 4'b0101;
																assign node4786 = (inp[5]) ? 4'b0101 : 4'b0111;
												assign node4789 = (inp[5]) ? node4797 : node4790;
													assign node4790 = (inp[0]) ? node4794 : node4791;
														assign node4791 = (inp[15]) ? 4'b0001 : 4'b0011;
														assign node4794 = (inp[15]) ? 4'b0011 : 4'b0001;
													assign node4797 = (inp[12]) ? node4807 : node4798;
														assign node4798 = (inp[3]) ? node4800 : 4'b0001;
															assign node4800 = (inp[0]) ? node4804 : node4801;
																assign node4801 = (inp[15]) ? 4'b0011 : 4'b0001;
																assign node4804 = (inp[15]) ? 4'b0001 : 4'b0011;
														assign node4807 = (inp[15]) ? node4815 : node4808;
															assign node4808 = (inp[0]) ? node4812 : node4809;
																assign node4809 = (inp[3]) ? 4'b0001 : 4'b0011;
																assign node4812 = (inp[3]) ? 4'b0011 : 4'b0001;
															assign node4815 = (inp[3]) ? 4'b0001 : node4816;
																assign node4816 = (inp[0]) ? 4'b0011 : 4'b0001;
											assign node4820 = (inp[4]) ? node4868 : node4821;
												assign node4821 = (inp[3]) ? node4849 : node4822;
													assign node4822 = (inp[12]) ? node4838 : node4823;
														assign node4823 = (inp[5]) ? node4831 : node4824;
															assign node4824 = (inp[0]) ? node4828 : node4825;
																assign node4825 = (inp[15]) ? 4'b0001 : 4'b0011;
																assign node4828 = (inp[15]) ? 4'b0011 : 4'b0001;
															assign node4831 = (inp[15]) ? node4835 : node4832;
																assign node4832 = (inp[0]) ? 4'b0001 : 4'b0011;
																assign node4835 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node4838 = (inp[5]) ? node4844 : node4839;
															assign node4839 = (inp[15]) ? node4841 : 4'b0001;
																assign node4841 = (inp[0]) ? 4'b0011 : 4'b0001;
															assign node4844 = (inp[15]) ? 4'b0001 : node4845;
																assign node4845 = (inp[0]) ? 4'b0001 : 4'b0011;
													assign node4849 = (inp[0]) ? node4857 : node4850;
														assign node4850 = (inp[15]) ? node4854 : node4851;
															assign node4851 = (inp[5]) ? 4'b0001 : 4'b0011;
															assign node4854 = (inp[5]) ? 4'b0011 : 4'b0001;
														assign node4857 = (inp[12]) ? node4863 : node4858;
															assign node4858 = (inp[5]) ? 4'b0001 : node4859;
																assign node4859 = (inp[15]) ? 4'b0011 : 4'b0001;
															assign node4863 = (inp[15]) ? 4'b0011 : node4864;
																assign node4864 = (inp[5]) ? 4'b0011 : 4'b0001;
												assign node4868 = (inp[3]) ? node4882 : node4869;
													assign node4869 = (inp[15]) ? node4875 : node4870;
														assign node4870 = (inp[12]) ? 4'b0111 : node4871;
															assign node4871 = (inp[0]) ? 4'b0111 : 4'b0101;
														assign node4875 = (inp[0]) ? node4879 : node4876;
															assign node4876 = (inp[5]) ? 4'b0111 : 4'b0101;
															assign node4879 = (inp[5]) ? 4'b0101 : 4'b0111;
													assign node4882 = (inp[0]) ? node4886 : node4883;
														assign node4883 = (inp[15]) ? 4'b0111 : 4'b0101;
														assign node4886 = (inp[15]) ? 4'b0101 : 4'b0111;
										assign node4889 = (inp[9]) ? node4923 : node4890;
											assign node4890 = (inp[4]) ? node4912 : node4891;
												assign node4891 = (inp[15]) ? node4903 : node4892;
													assign node4892 = (inp[0]) ? node4898 : node4893;
														assign node4893 = (inp[3]) ? node4895 : 4'b0110;
															assign node4895 = (inp[5]) ? 4'b0100 : 4'b0110;
														assign node4898 = (inp[5]) ? node4900 : 4'b0100;
															assign node4900 = (inp[3]) ? 4'b0110 : 4'b0100;
													assign node4903 = (inp[0]) ? node4907 : node4904;
														assign node4904 = (inp[3]) ? 4'b0110 : 4'b0100;
														assign node4907 = (inp[3]) ? node4909 : 4'b0110;
															assign node4909 = (inp[5]) ? 4'b0100 : 4'b0110;
												assign node4912 = (inp[0]) ? node4918 : node4913;
													assign node4913 = (inp[15]) ? 4'b0000 : node4914;
														assign node4914 = (inp[5]) ? 4'b0000 : 4'b0010;
													assign node4918 = (inp[15]) ? 4'b0010 : node4919;
														assign node4919 = (inp[3]) ? 4'b0010 : 4'b0000;
											assign node4923 = (inp[4]) ? node4947 : node4924;
												assign node4924 = (inp[15]) ? node4936 : node4925;
													assign node4925 = (inp[0]) ? node4931 : node4926;
														assign node4926 = (inp[3]) ? node4928 : 4'b0010;
															assign node4928 = (inp[5]) ? 4'b0000 : 4'b0010;
														assign node4931 = (inp[3]) ? node4933 : 4'b0000;
															assign node4933 = (inp[12]) ? 4'b0010 : 4'b0000;
													assign node4936 = (inp[0]) ? node4942 : node4937;
														assign node4937 = (inp[3]) ? node4939 : 4'b0000;
															assign node4939 = (inp[5]) ? 4'b0010 : 4'b0000;
														assign node4942 = (inp[3]) ? node4944 : 4'b0010;
															assign node4944 = (inp[5]) ? 4'b0000 : 4'b0010;
												assign node4947 = (inp[0]) ? node4961 : node4948;
													assign node4948 = (inp[12]) ? node4950 : 4'b0110;
														assign node4950 = (inp[15]) ? node4956 : node4951;
															assign node4951 = (inp[5]) ? 4'b0100 : node4952;
																assign node4952 = (inp[3]) ? 4'b0100 : 4'b0110;
															assign node4956 = (inp[3]) ? 4'b0110 : node4957;
																assign node4957 = (inp[5]) ? 4'b0110 : 4'b0100;
													assign node4961 = (inp[15]) ? 4'b0100 : node4962;
														assign node4962 = (inp[5]) ? 4'b0110 : 4'b0100;
									assign node4966 = (inp[3]) ? node5032 : node4967;
										assign node4967 = (inp[15]) ? node4999 : node4968;
											assign node4968 = (inp[0]) ? node4978 : node4969;
												assign node4969 = (inp[4]) ? node4973 : node4970;
													assign node4970 = (inp[9]) ? 4'b0010 : 4'b0110;
													assign node4973 = (inp[9]) ? node4975 : 4'b0010;
														assign node4975 = (inp[5]) ? 4'b0100 : 4'b0110;
												assign node4978 = (inp[5]) ? node4992 : node4979;
													assign node4979 = (inp[12]) ? node4987 : node4980;
														assign node4980 = (inp[4]) ? node4984 : node4981;
															assign node4981 = (inp[9]) ? 4'b0000 : 4'b0100;
															assign node4984 = (inp[9]) ? 4'b0100 : 4'b0000;
														assign node4987 = (inp[4]) ? node4989 : 4'b0100;
															assign node4989 = (inp[9]) ? 4'b0100 : 4'b0000;
													assign node4992 = (inp[9]) ? node4996 : node4993;
														assign node4993 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node4996 = (inp[4]) ? 4'b0110 : 4'b0000;
											assign node4999 = (inp[0]) ? node5023 : node5000;
												assign node5000 = (inp[5]) ? node5016 : node5001;
													assign node5001 = (inp[12]) ? node5009 : node5002;
														assign node5002 = (inp[9]) ? node5006 : node5003;
															assign node5003 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node5006 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node5009 = (inp[4]) ? node5013 : node5010;
															assign node5010 = (inp[9]) ? 4'b0000 : 4'b0100;
															assign node5013 = (inp[9]) ? 4'b0100 : 4'b0000;
													assign node5016 = (inp[9]) ? node5020 : node5017;
														assign node5017 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node5020 = (inp[4]) ? 4'b0110 : 4'b0000;
												assign node5023 = (inp[9]) ? node5027 : node5024;
													assign node5024 = (inp[4]) ? 4'b0010 : 4'b0110;
													assign node5027 = (inp[4]) ? node5029 : 4'b0010;
														assign node5029 = (inp[5]) ? 4'b0100 : 4'b0110;
										assign node5032 = (inp[0]) ? node5082 : node5033;
											assign node5033 = (inp[15]) ? node5063 : node5034;
												assign node5034 = (inp[5]) ? node5040 : node5035;
													assign node5035 = (inp[4]) ? node5037 : 4'b0010;
														assign node5037 = (inp[9]) ? 4'b0100 : 4'b0010;
													assign node5040 = (inp[12]) ? node5056 : node5041;
														assign node5041 = (inp[2]) ? node5049 : node5042;
															assign node5042 = (inp[9]) ? node5046 : node5043;
																assign node5043 = (inp[4]) ? 4'b0000 : 4'b0100;
																assign node5046 = (inp[4]) ? 4'b0100 : 4'b0000;
															assign node5049 = (inp[4]) ? node5053 : node5050;
																assign node5050 = (inp[9]) ? 4'b0000 : 4'b0100;
																assign node5053 = (inp[9]) ? 4'b0100 : 4'b0000;
														assign node5056 = (inp[4]) ? node5060 : node5057;
															assign node5057 = (inp[9]) ? 4'b0000 : 4'b0100;
															assign node5060 = (inp[9]) ? 4'b0100 : 4'b0000;
												assign node5063 = (inp[5]) ? node5071 : node5064;
													assign node5064 = (inp[9]) ? node5068 : node5065;
														assign node5065 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node5068 = (inp[4]) ? 4'b0110 : 4'b0000;
													assign node5071 = (inp[2]) ? node5077 : node5072;
														assign node5072 = (inp[4]) ? node5074 : 4'b0010;
															assign node5074 = (inp[9]) ? 4'b0110 : 4'b0010;
														assign node5077 = (inp[4]) ? 4'b0010 : node5078;
															assign node5078 = (inp[9]) ? 4'b0010 : 4'b0110;
											assign node5082 = (inp[15]) ? node5098 : node5083;
												assign node5083 = (inp[5]) ? node5091 : node5084;
													assign node5084 = (inp[4]) ? node5088 : node5085;
														assign node5085 = (inp[9]) ? 4'b0000 : 4'b0100;
														assign node5088 = (inp[9]) ? 4'b0110 : 4'b0000;
													assign node5091 = (inp[4]) ? node5095 : node5092;
														assign node5092 = (inp[9]) ? 4'b0010 : 4'b0110;
														assign node5095 = (inp[9]) ? 4'b0110 : 4'b0010;
												assign node5098 = (inp[5]) ? node5106 : node5099;
													assign node5099 = (inp[4]) ? node5103 : node5100;
														assign node5100 = (inp[9]) ? 4'b0010 : 4'b0110;
														assign node5103 = (inp[9]) ? 4'b0100 : 4'b0010;
													assign node5106 = (inp[12]) ? 4'b0100 : node5107;
														assign node5107 = (inp[4]) ? node5111 : node5108;
															assign node5108 = (inp[9]) ? 4'b0000 : 4'b0100;
															assign node5111 = (inp[9]) ? 4'b0100 : 4'b0000;
						assign node5115 = (inp[15]) ? node5963 : node5116;
							assign node5116 = (inp[0]) ? node5580 : node5117;
								assign node5117 = (inp[3]) ? node5369 : node5118;
									assign node5118 = (inp[5]) ? node5252 : node5119;
										assign node5119 = (inp[7]) ? node5195 : node5120;
											assign node5120 = (inp[8]) ? node5150 : node5121;
												assign node5121 = (inp[14]) ? node5133 : node5122;
													assign node5122 = (inp[2]) ? node5128 : node5123;
														assign node5123 = (inp[4]) ? 4'b0111 : node5124;
															assign node5124 = (inp[9]) ? 4'b0011 : 4'b0111;
														assign node5128 = (inp[4]) ? 4'b0110 : node5129;
															assign node5129 = (inp[9]) ? 4'b0010 : 4'b0110;
													assign node5133 = (inp[2]) ? node5141 : node5134;
														assign node5134 = (inp[9]) ? node5138 : node5135;
															assign node5135 = (inp[4]) ? 4'b0010 : 4'b0110;
															assign node5138 = (inp[4]) ? 4'b0110 : 4'b0010;
														assign node5141 = (inp[12]) ? node5145 : node5142;
															assign node5142 = (inp[9]) ? 4'b0110 : 4'b0010;
															assign node5145 = (inp[4]) ? 4'b0010 : node5146;
																assign node5146 = (inp[9]) ? 4'b0010 : 4'b0110;
												assign node5150 = (inp[14]) ? node5174 : node5151;
													assign node5151 = (inp[2]) ? node5167 : node5152;
														assign node5152 = (inp[12]) ? node5160 : node5153;
															assign node5153 = (inp[4]) ? node5157 : node5154;
																assign node5154 = (inp[9]) ? 4'b0010 : 4'b0110;
																assign node5157 = (inp[9]) ? 4'b0110 : 4'b0010;
															assign node5160 = (inp[4]) ? node5164 : node5161;
																assign node5161 = (inp[9]) ? 4'b0010 : 4'b0110;
																assign node5164 = (inp[9]) ? 4'b0110 : 4'b0010;
														assign node5167 = (inp[9]) ? node5171 : node5168;
															assign node5168 = (inp[4]) ? 4'b0011 : 4'b0111;
															assign node5171 = (inp[4]) ? 4'b0111 : 4'b0011;
													assign node5174 = (inp[12]) ? node5184 : node5175;
														assign node5175 = (inp[2]) ? 4'b0111 : node5176;
															assign node5176 = (inp[4]) ? node5180 : node5177;
																assign node5177 = (inp[9]) ? 4'b0011 : 4'b0111;
																assign node5180 = (inp[9]) ? 4'b0111 : 4'b0011;
														assign node5184 = (inp[2]) ? node5190 : node5185;
															assign node5185 = (inp[9]) ? node5187 : 4'b0111;
																assign node5187 = (inp[4]) ? 4'b0111 : 4'b0011;
															assign node5190 = (inp[9]) ? 4'b0011 : node5191;
																assign node5191 = (inp[4]) ? 4'b0011 : 4'b0111;
											assign node5195 = (inp[8]) ? node5233 : node5196;
												assign node5196 = (inp[2]) ? node5216 : node5197;
													assign node5197 = (inp[14]) ? node5205 : node5198;
														assign node5198 = (inp[4]) ? node5202 : node5199;
															assign node5199 = (inp[9]) ? 4'b0010 : 4'b0110;
															assign node5202 = (inp[9]) ? 4'b0110 : 4'b0010;
														assign node5205 = (inp[12]) ? node5211 : node5206;
															assign node5206 = (inp[9]) ? 4'b0011 : node5207;
																assign node5207 = (inp[4]) ? 4'b0011 : 4'b0111;
															assign node5211 = (inp[4]) ? node5213 : 4'b0011;
																assign node5213 = (inp[9]) ? 4'b0111 : 4'b0011;
													assign node5216 = (inp[12]) ? node5226 : node5217;
														assign node5217 = (inp[14]) ? node5219 : 4'b0011;
															assign node5219 = (inp[4]) ? node5223 : node5220;
																assign node5220 = (inp[9]) ? 4'b0011 : 4'b0111;
																assign node5223 = (inp[9]) ? 4'b0111 : 4'b0011;
														assign node5226 = (inp[9]) ? node5230 : node5227;
															assign node5227 = (inp[4]) ? 4'b0011 : 4'b0111;
															assign node5230 = (inp[4]) ? 4'b0111 : 4'b0011;
												assign node5233 = (inp[2]) ? node5245 : node5234;
													assign node5234 = (inp[14]) ? node5240 : node5235;
														assign node5235 = (inp[9]) ? node5237 : 4'b0111;
															assign node5237 = (inp[4]) ? 4'b0111 : 4'b0011;
														assign node5240 = (inp[9]) ? 4'b0110 : node5241;
															assign node5241 = (inp[4]) ? 4'b0010 : 4'b0110;
													assign node5245 = (inp[4]) ? node5249 : node5246;
														assign node5246 = (inp[9]) ? 4'b0010 : 4'b0110;
														assign node5249 = (inp[9]) ? 4'b0110 : 4'b0010;
										assign node5252 = (inp[4]) ? node5320 : node5253;
											assign node5253 = (inp[9]) ? node5283 : node5254;
												assign node5254 = (inp[8]) ? node5266 : node5255;
													assign node5255 = (inp[7]) ? node5261 : node5256;
														assign node5256 = (inp[14]) ? 4'b0110 : node5257;
															assign node5257 = (inp[2]) ? 4'b0110 : 4'b0111;
														assign node5261 = (inp[2]) ? 4'b0111 : node5262;
															assign node5262 = (inp[14]) ? 4'b0111 : 4'b0110;
													assign node5266 = (inp[12]) ? node5276 : node5267;
														assign node5267 = (inp[14]) ? 4'b0110 : node5268;
															assign node5268 = (inp[7]) ? node5272 : node5269;
																assign node5269 = (inp[2]) ? 4'b0111 : 4'b0110;
																assign node5272 = (inp[2]) ? 4'b0110 : 4'b0111;
														assign node5276 = (inp[7]) ? node5280 : node5277;
															assign node5277 = (inp[14]) ? 4'b0111 : 4'b0110;
															assign node5280 = (inp[2]) ? 4'b0110 : 4'b0111;
												assign node5283 = (inp[12]) ? node5301 : node5284;
													assign node5284 = (inp[8]) ? node5292 : node5285;
														assign node5285 = (inp[7]) ? node5289 : node5286;
															assign node5286 = (inp[2]) ? 4'b0010 : 4'b0011;
															assign node5289 = (inp[2]) ? 4'b0011 : 4'b0010;
														assign node5292 = (inp[2]) ? 4'b0010 : node5293;
															assign node5293 = (inp[14]) ? node5297 : node5294;
																assign node5294 = (inp[7]) ? 4'b0011 : 4'b0010;
																assign node5297 = (inp[7]) ? 4'b0010 : 4'b0011;
													assign node5301 = (inp[14]) ? node5315 : node5302;
														assign node5302 = (inp[8]) ? node5310 : node5303;
															assign node5303 = (inp[2]) ? node5307 : node5304;
																assign node5304 = (inp[7]) ? 4'b0010 : 4'b0011;
																assign node5307 = (inp[7]) ? 4'b0011 : 4'b0010;
															assign node5310 = (inp[7]) ? 4'b0011 : node5311;
																assign node5311 = (inp[2]) ? 4'b0011 : 4'b0010;
														assign node5315 = (inp[2]) ? node5317 : 4'b0011;
															assign node5317 = (inp[7]) ? 4'b0010 : 4'b0011;
											assign node5320 = (inp[9]) ? node5342 : node5321;
												assign node5321 = (inp[2]) ? node5335 : node5322;
													assign node5322 = (inp[7]) ? node5330 : node5323;
														assign node5323 = (inp[8]) ? node5327 : node5324;
															assign node5324 = (inp[14]) ? 4'b0010 : 4'b0011;
															assign node5327 = (inp[14]) ? 4'b0011 : 4'b0010;
														assign node5330 = (inp[8]) ? 4'b0011 : node5331;
															assign node5331 = (inp[14]) ? 4'b0011 : 4'b0010;
													assign node5335 = (inp[8]) ? node5339 : node5336;
														assign node5336 = (inp[7]) ? 4'b0011 : 4'b0010;
														assign node5339 = (inp[7]) ? 4'b0010 : 4'b0011;
												assign node5342 = (inp[14]) ? node5356 : node5343;
													assign node5343 = (inp[7]) ? 4'b0101 : node5344;
														assign node5344 = (inp[12]) ? node5350 : node5345;
															assign node5345 = (inp[2]) ? 4'b0100 : node5346;
																assign node5346 = (inp[8]) ? 4'b0100 : 4'b0101;
															assign node5350 = (inp[8]) ? 4'b0101 : node5351;
																assign node5351 = (inp[2]) ? 4'b0100 : 4'b0101;
													assign node5356 = (inp[2]) ? node5362 : node5357;
														assign node5357 = (inp[8]) ? node5359 : 4'b0100;
															assign node5359 = (inp[12]) ? 4'b0100 : 4'b0101;
														assign node5362 = (inp[8]) ? node5366 : node5363;
															assign node5363 = (inp[7]) ? 4'b0101 : 4'b0100;
															assign node5366 = (inp[7]) ? 4'b0100 : 4'b0101;
									assign node5369 = (inp[5]) ? node5475 : node5370;
										assign node5370 = (inp[9]) ? node5424 : node5371;
											assign node5371 = (inp[4]) ? node5393 : node5372;
												assign node5372 = (inp[2]) ? node5388 : node5373;
													assign node5373 = (inp[8]) ? node5381 : node5374;
														assign node5374 = (inp[7]) ? node5378 : node5375;
															assign node5375 = (inp[14]) ? 4'b0110 : 4'b0111;
															assign node5378 = (inp[14]) ? 4'b0111 : 4'b0110;
														assign node5381 = (inp[12]) ? 4'b0111 : node5382;
															assign node5382 = (inp[14]) ? node5384 : 4'b0111;
																assign node5384 = (inp[7]) ? 4'b0110 : 4'b0111;
													assign node5388 = (inp[8]) ? node5390 : 4'b0110;
														assign node5390 = (inp[7]) ? 4'b0110 : 4'b0111;
												assign node5393 = (inp[12]) ? node5405 : node5394;
													assign node5394 = (inp[7]) ? node5398 : node5395;
														assign node5395 = (inp[8]) ? 4'b0011 : 4'b0010;
														assign node5398 = (inp[8]) ? 4'b0010 : node5399;
															assign node5399 = (inp[2]) ? 4'b0011 : node5400;
																assign node5400 = (inp[14]) ? 4'b0011 : 4'b0010;
													assign node5405 = (inp[2]) ? node5417 : node5406;
														assign node5406 = (inp[14]) ? node5412 : node5407;
															assign node5407 = (inp[8]) ? node5409 : 4'b0011;
																assign node5409 = (inp[7]) ? 4'b0011 : 4'b0010;
															assign node5412 = (inp[8]) ? node5414 : 4'b0010;
																assign node5414 = (inp[7]) ? 4'b0010 : 4'b0011;
														assign node5417 = (inp[14]) ? node5419 : 4'b0010;
															assign node5419 = (inp[7]) ? node5421 : 4'b0010;
																assign node5421 = (inp[8]) ? 4'b0010 : 4'b0011;
											assign node5424 = (inp[4]) ? node5444 : node5425;
												assign node5425 = (inp[8]) ? node5435 : node5426;
													assign node5426 = (inp[7]) ? node5430 : node5427;
														assign node5427 = (inp[14]) ? 4'b0010 : 4'b0011;
														assign node5430 = (inp[14]) ? 4'b0011 : node5431;
															assign node5431 = (inp[2]) ? 4'b0011 : 4'b0010;
													assign node5435 = (inp[2]) ? node5441 : node5436;
														assign node5436 = (inp[7]) ? node5438 : 4'b0010;
															assign node5438 = (inp[14]) ? 4'b0010 : 4'b0011;
														assign node5441 = (inp[7]) ? 4'b0010 : 4'b0011;
												assign node5444 = (inp[12]) ? node5460 : node5445;
													assign node5445 = (inp[8]) ? node5451 : node5446;
														assign node5446 = (inp[7]) ? node5448 : 4'b0100;
															assign node5448 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node5451 = (inp[7]) ? node5457 : node5452;
															assign node5452 = (inp[2]) ? 4'b0101 : node5453;
																assign node5453 = (inp[14]) ? 4'b0101 : 4'b0100;
															assign node5457 = (inp[2]) ? 4'b0100 : 4'b0101;
													assign node5460 = (inp[7]) ? node5466 : node5461;
														assign node5461 = (inp[8]) ? 4'b0101 : node5462;
															assign node5462 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node5466 = (inp[8]) ? node5472 : node5467;
															assign node5467 = (inp[14]) ? 4'b0101 : node5468;
																assign node5468 = (inp[2]) ? 4'b0101 : 4'b0100;
															assign node5472 = (inp[14]) ? 4'b0100 : 4'b0101;
										assign node5475 = (inp[4]) ? node5523 : node5476;
											assign node5476 = (inp[9]) ? node5500 : node5477;
												assign node5477 = (inp[14]) ? node5493 : node5478;
													assign node5478 = (inp[8]) ? node5486 : node5479;
														assign node5479 = (inp[2]) ? node5483 : node5480;
															assign node5480 = (inp[7]) ? 4'b0100 : 4'b0101;
															assign node5483 = (inp[7]) ? 4'b0101 : 4'b0100;
														assign node5486 = (inp[2]) ? node5490 : node5487;
															assign node5487 = (inp[12]) ? 4'b0100 : 4'b0101;
															assign node5490 = (inp[7]) ? 4'b0100 : 4'b0101;
													assign node5493 = (inp[8]) ? node5497 : node5494;
														assign node5494 = (inp[7]) ? 4'b0101 : 4'b0100;
														assign node5497 = (inp[7]) ? 4'b0100 : 4'b0101;
												assign node5500 = (inp[7]) ? node5512 : node5501;
													assign node5501 = (inp[8]) ? node5507 : node5502;
														assign node5502 = (inp[2]) ? 4'b0000 : node5503;
															assign node5503 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node5507 = (inp[14]) ? 4'b0001 : node5508;
															assign node5508 = (inp[2]) ? 4'b0001 : 4'b0000;
													assign node5512 = (inp[8]) ? node5518 : node5513;
														assign node5513 = (inp[2]) ? 4'b0001 : node5514;
															assign node5514 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node5518 = (inp[14]) ? 4'b0000 : node5519;
															assign node5519 = (inp[2]) ? 4'b0000 : 4'b0001;
											assign node5523 = (inp[9]) ? node5557 : node5524;
												assign node5524 = (inp[12]) ? node5540 : node5525;
													assign node5525 = (inp[14]) ? 4'b0000 : node5526;
														assign node5526 = (inp[2]) ? node5534 : node5527;
															assign node5527 = (inp[8]) ? node5531 : node5528;
																assign node5528 = (inp[7]) ? 4'b0000 : 4'b0001;
																assign node5531 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node5534 = (inp[7]) ? 4'b0000 : node5535;
																assign node5535 = (inp[8]) ? 4'b0001 : 4'b0000;
													assign node5540 = (inp[14]) ? node5550 : node5541;
														assign node5541 = (inp[8]) ? 4'b0000 : node5542;
															assign node5542 = (inp[2]) ? node5546 : node5543;
																assign node5543 = (inp[7]) ? 4'b0000 : 4'b0001;
																assign node5546 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node5550 = (inp[8]) ? node5554 : node5551;
															assign node5551 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node5554 = (inp[7]) ? 4'b0000 : 4'b0001;
												assign node5557 = (inp[7]) ? node5569 : node5558;
													assign node5558 = (inp[8]) ? node5564 : node5559;
														assign node5559 = (inp[14]) ? 4'b0100 : node5560;
															assign node5560 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node5564 = (inp[14]) ? 4'b0101 : node5565;
															assign node5565 = (inp[2]) ? 4'b0101 : 4'b0100;
													assign node5569 = (inp[8]) ? node5575 : node5570;
														assign node5570 = (inp[2]) ? 4'b0101 : node5571;
															assign node5571 = (inp[14]) ? 4'b0101 : 4'b0100;
														assign node5575 = (inp[12]) ? node5577 : 4'b0100;
															assign node5577 = (inp[2]) ? 4'b0100 : 4'b0101;
								assign node5580 = (inp[3]) ? node5728 : node5581;
									assign node5581 = (inp[9]) ? node5645 : node5582;
										assign node5582 = (inp[4]) ? node5626 : node5583;
											assign node5583 = (inp[12]) ? node5603 : node5584;
												assign node5584 = (inp[7]) ? node5592 : node5585;
													assign node5585 = (inp[8]) ? 4'b0101 : node5586;
														assign node5586 = (inp[14]) ? 4'b0100 : node5587;
															assign node5587 = (inp[2]) ? 4'b0100 : 4'b0101;
													assign node5592 = (inp[8]) ? node5598 : node5593;
														assign node5593 = (inp[14]) ? 4'b0101 : node5594;
															assign node5594 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node5598 = (inp[14]) ? 4'b0100 : node5599;
															assign node5599 = (inp[2]) ? 4'b0100 : 4'b0101;
												assign node5603 = (inp[8]) ? node5615 : node5604;
													assign node5604 = (inp[7]) ? node5610 : node5605;
														assign node5605 = (inp[14]) ? 4'b0100 : node5606;
															assign node5606 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node5610 = (inp[14]) ? 4'b0101 : node5611;
															assign node5611 = (inp[2]) ? 4'b0101 : 4'b0100;
													assign node5615 = (inp[7]) ? node5621 : node5616;
														assign node5616 = (inp[14]) ? 4'b0101 : node5617;
															assign node5617 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node5621 = (inp[2]) ? 4'b0100 : node5622;
															assign node5622 = (inp[14]) ? 4'b0100 : 4'b0101;
											assign node5626 = (inp[8]) ? node5634 : node5627;
												assign node5627 = (inp[7]) ? node5629 : 4'b0000;
													assign node5629 = (inp[14]) ? 4'b0001 : node5630;
														assign node5630 = (inp[2]) ? 4'b0001 : 4'b0000;
												assign node5634 = (inp[7]) ? node5640 : node5635;
													assign node5635 = (inp[14]) ? 4'b0001 : node5636;
														assign node5636 = (inp[2]) ? 4'b0001 : 4'b0000;
													assign node5640 = (inp[14]) ? 4'b0000 : node5641;
														assign node5641 = (inp[2]) ? 4'b0000 : 4'b0001;
										assign node5645 = (inp[4]) ? node5669 : node5646;
											assign node5646 = (inp[7]) ? node5658 : node5647;
												assign node5647 = (inp[8]) ? node5653 : node5648;
													assign node5648 = (inp[14]) ? 4'b0000 : node5649;
														assign node5649 = (inp[2]) ? 4'b0000 : 4'b0001;
													assign node5653 = (inp[2]) ? 4'b0001 : node5654;
														assign node5654 = (inp[14]) ? 4'b0001 : 4'b0000;
												assign node5658 = (inp[8]) ? node5664 : node5659;
													assign node5659 = (inp[14]) ? 4'b0001 : node5660;
														assign node5660 = (inp[2]) ? 4'b0001 : 4'b0000;
													assign node5664 = (inp[2]) ? 4'b0000 : node5665;
														assign node5665 = (inp[14]) ? 4'b0000 : 4'b0001;
											assign node5669 = (inp[5]) ? node5703 : node5670;
												assign node5670 = (inp[2]) ? node5690 : node5671;
													assign node5671 = (inp[14]) ? node5685 : node5672;
														assign node5672 = (inp[12]) ? node5680 : node5673;
															assign node5673 = (inp[8]) ? node5677 : node5674;
																assign node5674 = (inp[7]) ? 4'b0100 : 4'b0101;
																assign node5677 = (inp[7]) ? 4'b0101 : 4'b0100;
															assign node5680 = (inp[7]) ? 4'b0101 : node5681;
																assign node5681 = (inp[8]) ? 4'b0100 : 4'b0101;
														assign node5685 = (inp[7]) ? node5687 : 4'b0101;
															assign node5687 = (inp[8]) ? 4'b0100 : 4'b0101;
													assign node5690 = (inp[12]) ? node5698 : node5691;
														assign node5691 = (inp[8]) ? node5695 : node5692;
															assign node5692 = (inp[7]) ? 4'b0101 : 4'b0100;
															assign node5695 = (inp[7]) ? 4'b0100 : 4'b0101;
														assign node5698 = (inp[8]) ? node5700 : 4'b0100;
															assign node5700 = (inp[7]) ? 4'b0100 : 4'b0101;
												assign node5703 = (inp[12]) ? node5719 : node5704;
													assign node5704 = (inp[2]) ? node5714 : node5705;
														assign node5705 = (inp[8]) ? node5707 : 4'b0110;
															assign node5707 = (inp[7]) ? node5711 : node5708;
																assign node5708 = (inp[14]) ? 4'b0111 : 4'b0110;
																assign node5711 = (inp[14]) ? 4'b0110 : 4'b0111;
														assign node5714 = (inp[7]) ? node5716 : 4'b0110;
															assign node5716 = (inp[8]) ? 4'b0110 : 4'b0111;
													assign node5719 = (inp[14]) ? node5721 : 4'b0111;
														assign node5721 = (inp[8]) ? node5725 : node5722;
															assign node5722 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node5725 = (inp[7]) ? 4'b0110 : 4'b0111;
									assign node5728 = (inp[5]) ? node5824 : node5729;
										assign node5729 = (inp[9]) ? node5779 : node5730;
											assign node5730 = (inp[4]) ? node5752 : node5731;
												assign node5731 = (inp[7]) ? node5743 : node5732;
													assign node5732 = (inp[8]) ? node5738 : node5733;
														assign node5733 = (inp[14]) ? 4'b0100 : node5734;
															assign node5734 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node5738 = (inp[14]) ? 4'b0101 : node5739;
															assign node5739 = (inp[2]) ? 4'b0101 : 4'b0100;
													assign node5743 = (inp[8]) ? node5747 : node5744;
														assign node5744 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node5747 = (inp[2]) ? 4'b0100 : node5748;
															assign node5748 = (inp[14]) ? 4'b0100 : 4'b0101;
												assign node5752 = (inp[12]) ? node5770 : node5753;
													assign node5753 = (inp[8]) ? node5761 : node5754;
														assign node5754 = (inp[7]) ? node5756 : 4'b0000;
															assign node5756 = (inp[14]) ? 4'b0001 : node5757;
																assign node5757 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node5761 = (inp[7]) ? node5767 : node5762;
															assign node5762 = (inp[14]) ? 4'b0001 : node5763;
																assign node5763 = (inp[2]) ? 4'b0001 : 4'b0000;
															assign node5767 = (inp[2]) ? 4'b0000 : 4'b0001;
													assign node5770 = (inp[7]) ? node5774 : node5771;
														assign node5771 = (inp[8]) ? 4'b0001 : 4'b0000;
														assign node5774 = (inp[8]) ? 4'b0000 : node5775;
															assign node5775 = (inp[2]) ? 4'b0001 : 4'b0000;
											assign node5779 = (inp[4]) ? node5797 : node5780;
												assign node5780 = (inp[8]) ? node5788 : node5781;
													assign node5781 = (inp[7]) ? node5783 : 4'b0000;
														assign node5783 = (inp[14]) ? 4'b0001 : node5784;
															assign node5784 = (inp[2]) ? 4'b0001 : 4'b0000;
													assign node5788 = (inp[2]) ? node5794 : node5789;
														assign node5789 = (inp[7]) ? 4'b0001 : node5790;
															assign node5790 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node5794 = (inp[7]) ? 4'b0000 : 4'b0001;
												assign node5797 = (inp[14]) ? node5817 : node5798;
													assign node5798 = (inp[8]) ? node5812 : node5799;
														assign node5799 = (inp[12]) ? node5805 : node5800;
															assign node5800 = (inp[7]) ? 4'b0110 : node5801;
																assign node5801 = (inp[2]) ? 4'b0110 : 4'b0111;
															assign node5805 = (inp[7]) ? node5809 : node5806;
																assign node5806 = (inp[2]) ? 4'b0110 : 4'b0111;
																assign node5809 = (inp[2]) ? 4'b0111 : 4'b0110;
														assign node5812 = (inp[7]) ? 4'b0111 : node5813;
															assign node5813 = (inp[2]) ? 4'b0111 : 4'b0110;
													assign node5817 = (inp[8]) ? node5821 : node5818;
														assign node5818 = (inp[7]) ? 4'b0111 : 4'b0110;
														assign node5821 = (inp[7]) ? 4'b0110 : 4'b0111;
										assign node5824 = (inp[12]) ? node5898 : node5825;
											assign node5825 = (inp[2]) ? node5875 : node5826;
												assign node5826 = (inp[14]) ? node5852 : node5827;
													assign node5827 = (inp[9]) ? node5841 : node5828;
														assign node5828 = (inp[4]) ? node5836 : node5829;
															assign node5829 = (inp[7]) ? node5833 : node5830;
																assign node5830 = (inp[8]) ? 4'b0110 : 4'b0111;
																assign node5833 = (inp[8]) ? 4'b0111 : 4'b0110;
															assign node5836 = (inp[7]) ? 4'b0010 : node5837;
																assign node5837 = (inp[8]) ? 4'b0010 : 4'b0011;
														assign node5841 = (inp[4]) ? node5845 : node5842;
															assign node5842 = (inp[7]) ? 4'b0011 : 4'b0010;
															assign node5845 = (inp[7]) ? node5849 : node5846;
																assign node5846 = (inp[8]) ? 4'b0110 : 4'b0111;
																assign node5849 = (inp[8]) ? 4'b0111 : 4'b0110;
													assign node5852 = (inp[8]) ? node5862 : node5853;
														assign node5853 = (inp[7]) ? node5859 : node5854;
															assign node5854 = (inp[9]) ? 4'b0010 : node5855;
																assign node5855 = (inp[4]) ? 4'b0010 : 4'b0110;
															assign node5859 = (inp[9]) ? 4'b0111 : 4'b0011;
														assign node5862 = (inp[7]) ? node5868 : node5863;
															assign node5863 = (inp[4]) ? 4'b0111 : node5864;
																assign node5864 = (inp[9]) ? 4'b0011 : 4'b0111;
															assign node5868 = (inp[4]) ? node5872 : node5869;
																assign node5869 = (inp[9]) ? 4'b0010 : 4'b0110;
																assign node5872 = (inp[9]) ? 4'b0110 : 4'b0010;
												assign node5875 = (inp[8]) ? node5887 : node5876;
													assign node5876 = (inp[7]) ? node5882 : node5877;
														assign node5877 = (inp[9]) ? node5879 : 4'b0110;
															assign node5879 = (inp[4]) ? 4'b0110 : 4'b0010;
														assign node5882 = (inp[9]) ? node5884 : 4'b0111;
															assign node5884 = (inp[4]) ? 4'b0111 : 4'b0011;
													assign node5887 = (inp[7]) ? node5895 : node5888;
														assign node5888 = (inp[4]) ? node5892 : node5889;
															assign node5889 = (inp[9]) ? 4'b0011 : 4'b0111;
															assign node5892 = (inp[9]) ? 4'b0111 : 4'b0011;
														assign node5895 = (inp[9]) ? 4'b0110 : 4'b0010;
											assign node5898 = (inp[8]) ? node5922 : node5899;
												assign node5899 = (inp[7]) ? node5909 : node5900;
													assign node5900 = (inp[2]) ? node5902 : 4'b0011;
														assign node5902 = (inp[9]) ? node5906 : node5903;
															assign node5903 = (inp[4]) ? 4'b0010 : 4'b0110;
															assign node5906 = (inp[4]) ? 4'b0110 : 4'b0010;
													assign node5909 = (inp[2]) ? node5919 : node5910;
														assign node5910 = (inp[14]) ? 4'b0111 : node5911;
															assign node5911 = (inp[9]) ? node5915 : node5912;
																assign node5912 = (inp[4]) ? 4'b0010 : 4'b0110;
																assign node5915 = (inp[4]) ? 4'b0110 : 4'b0010;
														assign node5919 = (inp[9]) ? 4'b0011 : 4'b0111;
												assign node5922 = (inp[7]) ? node5942 : node5923;
													assign node5923 = (inp[14]) ? node5933 : node5924;
														assign node5924 = (inp[2]) ? node5930 : node5925;
															assign node5925 = (inp[4]) ? node5927 : 4'b0010;
																assign node5927 = (inp[9]) ? 4'b0110 : 4'b0010;
															assign node5930 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node5933 = (inp[2]) ? 4'b0111 : node5934;
															assign node5934 = (inp[4]) ? node5938 : node5935;
																assign node5935 = (inp[9]) ? 4'b0011 : 4'b0111;
																assign node5938 = (inp[9]) ? 4'b0111 : 4'b0011;
													assign node5942 = (inp[14]) ? node5950 : node5943;
														assign node5943 = (inp[2]) ? 4'b0010 : node5944;
															assign node5944 = (inp[9]) ? node5946 : 4'b0111;
																assign node5946 = (inp[4]) ? 4'b0111 : 4'b0011;
														assign node5950 = (inp[2]) ? node5956 : node5951;
															assign node5951 = (inp[9]) ? 4'b0010 : node5952;
																assign node5952 = (inp[4]) ? 4'b0010 : 4'b0110;
															assign node5956 = (inp[4]) ? node5960 : node5957;
																assign node5957 = (inp[9]) ? 4'b0010 : 4'b0110;
																assign node5960 = (inp[9]) ? 4'b0110 : 4'b0010;
							assign node5963 = (inp[0]) ? node6417 : node5964;
								assign node5964 = (inp[5]) ? node6160 : node5965;
									assign node5965 = (inp[4]) ? node6075 : node5966;
										assign node5966 = (inp[9]) ? node6018 : node5967;
											assign node5967 = (inp[14]) ? node6003 : node5968;
												assign node5968 = (inp[12]) ? node5984 : node5969;
													assign node5969 = (inp[7]) ? node5977 : node5970;
														assign node5970 = (inp[2]) ? node5974 : node5971;
															assign node5971 = (inp[8]) ? 4'b0100 : 4'b0101;
															assign node5974 = (inp[8]) ? 4'b0101 : 4'b0100;
														assign node5977 = (inp[8]) ? node5981 : node5978;
															assign node5978 = (inp[3]) ? 4'b0101 : 4'b0100;
															assign node5981 = (inp[3]) ? 4'b0100 : 4'b0101;
													assign node5984 = (inp[7]) ? node5992 : node5985;
														assign node5985 = (inp[8]) ? node5989 : node5986;
															assign node5986 = (inp[2]) ? 4'b0100 : 4'b0101;
															assign node5989 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node5992 = (inp[3]) ? node5998 : node5993;
															assign node5993 = (inp[8]) ? 4'b0101 : node5994;
																assign node5994 = (inp[2]) ? 4'b0101 : 4'b0100;
															assign node5998 = (inp[8]) ? node6000 : 4'b0101;
																assign node6000 = (inp[2]) ? 4'b0100 : 4'b0101;
												assign node6003 = (inp[2]) ? node6011 : node6004;
													assign node6004 = (inp[7]) ? node6008 : node6005;
														assign node6005 = (inp[8]) ? 4'b0101 : 4'b0100;
														assign node6008 = (inp[8]) ? 4'b0100 : 4'b0101;
													assign node6011 = (inp[8]) ? node6015 : node6012;
														assign node6012 = (inp[7]) ? 4'b0101 : 4'b0100;
														assign node6015 = (inp[7]) ? 4'b0100 : 4'b0101;
											assign node6018 = (inp[14]) ? node6040 : node6019;
												assign node6019 = (inp[7]) ? node6027 : node6020;
													assign node6020 = (inp[2]) ? node6024 : node6021;
														assign node6021 = (inp[8]) ? 4'b0000 : 4'b0001;
														assign node6024 = (inp[8]) ? 4'b0001 : 4'b0000;
													assign node6027 = (inp[3]) ? node6033 : node6028;
														assign node6028 = (inp[2]) ? node6030 : 4'b0000;
															assign node6030 = (inp[8]) ? 4'b0000 : 4'b0001;
														assign node6033 = (inp[2]) ? node6037 : node6034;
															assign node6034 = (inp[8]) ? 4'b0001 : 4'b0000;
															assign node6037 = (inp[8]) ? 4'b0000 : 4'b0001;
												assign node6040 = (inp[2]) ? node6058 : node6041;
													assign node6041 = (inp[3]) ? node6049 : node6042;
														assign node6042 = (inp[8]) ? node6046 : node6043;
															assign node6043 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node6046 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node6049 = (inp[12]) ? node6051 : 4'b0000;
															assign node6051 = (inp[8]) ? node6055 : node6052;
																assign node6052 = (inp[7]) ? 4'b0001 : 4'b0000;
																assign node6055 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node6058 = (inp[12]) ? node6068 : node6059;
														assign node6059 = (inp[3]) ? node6065 : node6060;
															assign node6060 = (inp[7]) ? 4'b0001 : node6061;
																assign node6061 = (inp[8]) ? 4'b0001 : 4'b0000;
															assign node6065 = (inp[8]) ? 4'b0000 : 4'b0001;
														assign node6068 = (inp[8]) ? node6072 : node6069;
															assign node6069 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node6072 = (inp[7]) ? 4'b0000 : 4'b0001;
										assign node6075 = (inp[9]) ? node6121 : node6076;
											assign node6076 = (inp[2]) ? node6100 : node6077;
												assign node6077 = (inp[14]) ? node6087 : node6078;
													assign node6078 = (inp[12]) ? node6080 : 4'b0000;
														assign node6080 = (inp[8]) ? node6084 : node6081;
															assign node6081 = (inp[7]) ? 4'b0000 : 4'b0001;
															assign node6084 = (inp[7]) ? 4'b0001 : 4'b0000;
													assign node6087 = (inp[3]) ? node6093 : node6088;
														assign node6088 = (inp[12]) ? node6090 : 4'b0001;
															assign node6090 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node6093 = (inp[7]) ? node6097 : node6094;
															assign node6094 = (inp[8]) ? 4'b0001 : 4'b0000;
															assign node6097 = (inp[8]) ? 4'b0000 : 4'b0001;
												assign node6100 = (inp[14]) ? node6108 : node6101;
													assign node6101 = (inp[8]) ? node6105 : node6102;
														assign node6102 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node6105 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node6108 = (inp[3]) ? node6114 : node6109;
														assign node6109 = (inp[7]) ? 4'b0001 : node6110;
															assign node6110 = (inp[8]) ? 4'b0001 : 4'b0000;
														assign node6114 = (inp[7]) ? node6118 : node6115;
															assign node6115 = (inp[8]) ? 4'b0001 : 4'b0000;
															assign node6118 = (inp[8]) ? 4'b0000 : 4'b0001;
											assign node6121 = (inp[3]) ? node6143 : node6122;
												assign node6122 = (inp[2]) ? node6136 : node6123;
													assign node6123 = (inp[12]) ? node6131 : node6124;
														assign node6124 = (inp[8]) ? 4'b0101 : node6125;
															assign node6125 = (inp[14]) ? node6127 : 4'b0100;
																assign node6127 = (inp[7]) ? 4'b0101 : 4'b0100;
														assign node6131 = (inp[7]) ? node6133 : 4'b0101;
															assign node6133 = (inp[8]) ? 4'b0100 : 4'b0101;
													assign node6136 = (inp[8]) ? node6140 : node6137;
														assign node6137 = (inp[7]) ? 4'b0101 : 4'b0100;
														assign node6140 = (inp[7]) ? 4'b0100 : 4'b0101;
												assign node6143 = (inp[7]) ? node6155 : node6144;
													assign node6144 = (inp[8]) ? node6150 : node6145;
														assign node6145 = (inp[14]) ? 4'b0110 : node6146;
															assign node6146 = (inp[2]) ? 4'b0110 : 4'b0111;
														assign node6150 = (inp[2]) ? 4'b0111 : node6151;
															assign node6151 = (inp[14]) ? 4'b0111 : 4'b0110;
													assign node6155 = (inp[8]) ? node6157 : 4'b0111;
														assign node6157 = (inp[14]) ? 4'b0110 : 4'b0111;
									assign node6160 = (inp[3]) ? node6286 : node6161;
										assign node6161 = (inp[9]) ? node6221 : node6162;
											assign node6162 = (inp[4]) ? node6198 : node6163;
												assign node6163 = (inp[14]) ? node6183 : node6164;
													assign node6164 = (inp[12]) ? node6174 : node6165;
														assign node6165 = (inp[8]) ? 4'b0100 : node6166;
															assign node6166 = (inp[2]) ? node6170 : node6167;
																assign node6167 = (inp[7]) ? 4'b0100 : 4'b0101;
																assign node6170 = (inp[7]) ? 4'b0101 : 4'b0100;
														assign node6174 = (inp[8]) ? node6176 : 4'b0100;
															assign node6176 = (inp[2]) ? node6180 : node6177;
																assign node6177 = (inp[7]) ? 4'b0101 : 4'b0100;
																assign node6180 = (inp[7]) ? 4'b0100 : 4'b0101;
													assign node6183 = (inp[2]) ? node6191 : node6184;
														assign node6184 = (inp[12]) ? node6186 : 4'b0101;
															assign node6186 = (inp[7]) ? 4'b0101 : node6187;
																assign node6187 = (inp[8]) ? 4'b0101 : 4'b0100;
														assign node6191 = (inp[8]) ? node6195 : node6192;
															assign node6192 = (inp[7]) ? 4'b0101 : 4'b0100;
															assign node6195 = (inp[7]) ? 4'b0100 : 4'b0101;
												assign node6198 = (inp[8]) ? node6210 : node6199;
													assign node6199 = (inp[7]) ? node6205 : node6200;
														assign node6200 = (inp[2]) ? 4'b0000 : node6201;
															assign node6201 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node6205 = (inp[2]) ? 4'b0001 : node6206;
															assign node6206 = (inp[14]) ? 4'b0001 : 4'b0000;
													assign node6210 = (inp[2]) ? node6218 : node6211;
														assign node6211 = (inp[14]) ? node6215 : node6212;
															assign node6212 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node6215 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node6218 = (inp[7]) ? 4'b0000 : 4'b0001;
											assign node6221 = (inp[4]) ? node6255 : node6222;
												assign node6222 = (inp[14]) ? node6236 : node6223;
													assign node6223 = (inp[7]) ? node6231 : node6224;
														assign node6224 = (inp[8]) ? node6228 : node6225;
															assign node6225 = (inp[2]) ? 4'b0000 : 4'b0001;
															assign node6228 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node6231 = (inp[2]) ? node6233 : 4'b0001;
															assign node6233 = (inp[8]) ? 4'b0000 : 4'b0001;
													assign node6236 = (inp[12]) ? node6248 : node6237;
														assign node6237 = (inp[2]) ? node6243 : node6238;
															assign node6238 = (inp[7]) ? 4'b0001 : node6239;
																assign node6239 = (inp[8]) ? 4'b0001 : 4'b0000;
															assign node6243 = (inp[8]) ? node6245 : 4'b0000;
																assign node6245 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node6248 = (inp[2]) ? 4'b0000 : node6249;
															assign node6249 = (inp[8]) ? 4'b0000 : node6250;
																assign node6250 = (inp[7]) ? 4'b0001 : 4'b0000;
												assign node6255 = (inp[12]) ? node6269 : node6256;
													assign node6256 = (inp[14]) ? node6262 : node6257;
														assign node6257 = (inp[7]) ? node6259 : 4'b0111;
															assign node6259 = (inp[8]) ? 4'b0110 : 4'b0111;
														assign node6262 = (inp[8]) ? node6266 : node6263;
															assign node6263 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node6266 = (inp[7]) ? 4'b0110 : 4'b0111;
													assign node6269 = (inp[8]) ? node6275 : node6270;
														assign node6270 = (inp[14]) ? node6272 : 4'b0110;
															assign node6272 = (inp[7]) ? 4'b0111 : 4'b0110;
														assign node6275 = (inp[7]) ? node6281 : node6276;
															assign node6276 = (inp[2]) ? 4'b0111 : node6277;
																assign node6277 = (inp[14]) ? 4'b0111 : 4'b0110;
															assign node6281 = (inp[2]) ? 4'b0110 : node6282;
																assign node6282 = (inp[14]) ? 4'b0110 : 4'b0111;
										assign node6286 = (inp[14]) ? node6350 : node6287;
											assign node6287 = (inp[8]) ? node6329 : node6288;
												assign node6288 = (inp[7]) ? node6314 : node6289;
													assign node6289 = (inp[2]) ? node6301 : node6290;
														assign node6290 = (inp[12]) ? node6296 : node6291;
															assign node6291 = (inp[4]) ? node6293 : 4'b0011;
																assign node6293 = (inp[9]) ? 4'b0111 : 4'b0011;
															assign node6296 = (inp[9]) ? 4'b0011 : node6297;
																assign node6297 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node6301 = (inp[12]) ? node6309 : node6302;
															assign node6302 = (inp[4]) ? node6306 : node6303;
																assign node6303 = (inp[9]) ? 4'b0010 : 4'b0110;
																assign node6306 = (inp[9]) ? 4'b0110 : 4'b0010;
															assign node6309 = (inp[4]) ? node6311 : 4'b0010;
																assign node6311 = (inp[9]) ? 4'b0110 : 4'b0010;
													assign node6314 = (inp[2]) ? node6322 : node6315;
														assign node6315 = (inp[12]) ? 4'b0010 : node6316;
															assign node6316 = (inp[4]) ? 4'b0110 : node6317;
																assign node6317 = (inp[9]) ? 4'b0010 : 4'b0110;
														assign node6322 = (inp[4]) ? node6326 : node6323;
															assign node6323 = (inp[9]) ? 4'b0011 : 4'b0111;
															assign node6326 = (inp[9]) ? 4'b0111 : 4'b0011;
												assign node6329 = (inp[7]) ? node6347 : node6330;
													assign node6330 = (inp[2]) ? node6338 : node6331;
														assign node6331 = (inp[4]) ? node6335 : node6332;
															assign node6332 = (inp[9]) ? 4'b0010 : 4'b0110;
															assign node6335 = (inp[9]) ? 4'b0110 : 4'b0010;
														assign node6338 = (inp[12]) ? 4'b0011 : node6339;
															assign node6339 = (inp[9]) ? node6343 : node6340;
																assign node6340 = (inp[4]) ? 4'b0011 : 4'b0111;
																assign node6343 = (inp[4]) ? 4'b0111 : 4'b0011;
													assign node6347 = (inp[2]) ? 4'b0010 : 4'b0011;
											assign node6350 = (inp[2]) ? node6382 : node6351;
												assign node6351 = (inp[8]) ? node6367 : node6352;
													assign node6352 = (inp[7]) ? node6360 : node6353;
														assign node6353 = (inp[4]) ? node6357 : node6354;
															assign node6354 = (inp[9]) ? 4'b0010 : 4'b0110;
															assign node6357 = (inp[9]) ? 4'b0110 : 4'b0010;
														assign node6360 = (inp[12]) ? node6362 : 4'b0111;
															assign node6362 = (inp[9]) ? 4'b0011 : node6363;
																assign node6363 = (inp[4]) ? 4'b0011 : 4'b0111;
													assign node6367 = (inp[7]) ? node6373 : node6368;
														assign node6368 = (inp[9]) ? 4'b0111 : node6369;
															assign node6369 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node6373 = (inp[12]) ? node6375 : 4'b0110;
															assign node6375 = (inp[9]) ? node6379 : node6376;
																assign node6376 = (inp[4]) ? 4'b0010 : 4'b0110;
																assign node6379 = (inp[4]) ? 4'b0110 : 4'b0010;
												assign node6382 = (inp[7]) ? node6398 : node6383;
													assign node6383 = (inp[8]) ? node6391 : node6384;
														assign node6384 = (inp[12]) ? node6386 : 4'b0010;
															assign node6386 = (inp[9]) ? node6388 : 4'b0010;
																assign node6388 = (inp[4]) ? 4'b0110 : 4'b0010;
														assign node6391 = (inp[12]) ? 4'b0011 : node6392;
															assign node6392 = (inp[4]) ? 4'b0011 : node6393;
																assign node6393 = (inp[9]) ? 4'b0011 : 4'b0111;
													assign node6398 = (inp[8]) ? node6412 : node6399;
														assign node6399 = (inp[12]) ? node6407 : node6400;
															assign node6400 = (inp[4]) ? node6404 : node6401;
																assign node6401 = (inp[9]) ? 4'b0011 : 4'b0111;
																assign node6404 = (inp[9]) ? 4'b0111 : 4'b0011;
															assign node6407 = (inp[4]) ? node6409 : 4'b0011;
																assign node6409 = (inp[9]) ? 4'b0111 : 4'b0011;
														assign node6412 = (inp[9]) ? node6414 : 4'b0110;
															assign node6414 = (inp[4]) ? 4'b0110 : 4'b0010;
								assign node6417 = (inp[3]) ? node6559 : node6418;
									assign node6418 = (inp[9]) ? node6498 : node6419;
										assign node6419 = (inp[4]) ? node6465 : node6420;
											assign node6420 = (inp[14]) ? node6446 : node6421;
												assign node6421 = (inp[12]) ? node6431 : node6422;
													assign node6422 = (inp[2]) ? 4'b0111 : node6423;
														assign node6423 = (inp[8]) ? node6427 : node6424;
															assign node6424 = (inp[7]) ? 4'b0110 : 4'b0111;
															assign node6427 = (inp[7]) ? 4'b0111 : 4'b0110;
													assign node6431 = (inp[2]) ? node6441 : node6432;
														assign node6432 = (inp[5]) ? 4'b0110 : node6433;
															assign node6433 = (inp[7]) ? node6437 : node6434;
																assign node6434 = (inp[8]) ? 4'b0110 : 4'b0111;
																assign node6437 = (inp[8]) ? 4'b0111 : 4'b0110;
														assign node6441 = (inp[7]) ? 4'b0110 : node6442;
															assign node6442 = (inp[5]) ? 4'b0111 : 4'b0110;
												assign node6446 = (inp[12]) ? node6452 : node6447;
													assign node6447 = (inp[8]) ? node6449 : 4'b0110;
														assign node6449 = (inp[7]) ? 4'b0110 : 4'b0111;
													assign node6452 = (inp[2]) ? node6460 : node6453;
														assign node6453 = (inp[7]) ? node6457 : node6454;
															assign node6454 = (inp[8]) ? 4'b0111 : 4'b0110;
															assign node6457 = (inp[8]) ? 4'b0110 : 4'b0111;
														assign node6460 = (inp[7]) ? node6462 : 4'b0111;
															assign node6462 = (inp[8]) ? 4'b0110 : 4'b0111;
											assign node6465 = (inp[2]) ? node6491 : node6466;
												assign node6466 = (inp[7]) ? node6486 : node6467;
													assign node6467 = (inp[12]) ? node6475 : node6468;
														assign node6468 = (inp[14]) ? node6472 : node6469;
															assign node6469 = (inp[8]) ? 4'b0010 : 4'b0011;
															assign node6472 = (inp[8]) ? 4'b0011 : 4'b0010;
														assign node6475 = (inp[5]) ? node6481 : node6476;
															assign node6476 = (inp[14]) ? 4'b0010 : node6477;
																assign node6477 = (inp[8]) ? 4'b0010 : 4'b0011;
															assign node6481 = (inp[8]) ? node6483 : 4'b0010;
																assign node6483 = (inp[14]) ? 4'b0011 : 4'b0010;
													assign node6486 = (inp[14]) ? 4'b0011 : node6487;
														assign node6487 = (inp[8]) ? 4'b0011 : 4'b0010;
												assign node6491 = (inp[8]) ? node6495 : node6492;
													assign node6492 = (inp[7]) ? 4'b0011 : 4'b0010;
													assign node6495 = (inp[7]) ? 4'b0010 : 4'b0011;
										assign node6498 = (inp[4]) ? node6522 : node6499;
											assign node6499 = (inp[7]) ? node6511 : node6500;
												assign node6500 = (inp[8]) ? node6506 : node6501;
													assign node6501 = (inp[2]) ? 4'b0010 : node6502;
														assign node6502 = (inp[14]) ? 4'b0010 : 4'b0011;
													assign node6506 = (inp[2]) ? 4'b0011 : node6507;
														assign node6507 = (inp[14]) ? 4'b0011 : 4'b0010;
												assign node6511 = (inp[8]) ? node6517 : node6512;
													assign node6512 = (inp[2]) ? 4'b0011 : node6513;
														assign node6513 = (inp[14]) ? 4'b0011 : 4'b0010;
													assign node6517 = (inp[2]) ? 4'b0010 : node6518;
														assign node6518 = (inp[14]) ? 4'b0010 : 4'b0011;
											assign node6522 = (inp[5]) ? node6540 : node6523;
												assign node6523 = (inp[14]) ? node6533 : node6524;
													assign node6524 = (inp[8]) ? 4'b0111 : node6525;
														assign node6525 = (inp[2]) ? node6529 : node6526;
															assign node6526 = (inp[7]) ? 4'b0110 : 4'b0111;
															assign node6529 = (inp[7]) ? 4'b0111 : 4'b0110;
													assign node6533 = (inp[12]) ? 4'b0110 : node6534;
														assign node6534 = (inp[7]) ? node6536 : 4'b0111;
															assign node6536 = (inp[8]) ? 4'b0110 : 4'b0111;
												assign node6540 = (inp[8]) ? node6548 : node6541;
													assign node6541 = (inp[7]) ? 4'b0101 : node6542;
														assign node6542 = (inp[2]) ? 4'b0100 : node6543;
															assign node6543 = (inp[14]) ? 4'b0100 : 4'b0101;
													assign node6548 = (inp[7]) ? node6554 : node6549;
														assign node6549 = (inp[14]) ? 4'b0101 : node6550;
															assign node6550 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node6554 = (inp[14]) ? 4'b0100 : node6555;
															assign node6555 = (inp[2]) ? 4'b0100 : 4'b0101;
									assign node6559 = (inp[5]) ? node6683 : node6560;
										assign node6560 = (inp[9]) ? node6616 : node6561;
											assign node6561 = (inp[4]) ? node6595 : node6562;
												assign node6562 = (inp[2]) ? node6580 : node6563;
													assign node6563 = (inp[8]) ? node6573 : node6564;
														assign node6564 = (inp[12]) ? node6566 : 4'b0111;
															assign node6566 = (inp[14]) ? node6570 : node6567;
																assign node6567 = (inp[7]) ? 4'b0110 : 4'b0111;
																assign node6570 = (inp[7]) ? 4'b0111 : 4'b0110;
														assign node6573 = (inp[7]) ? node6577 : node6574;
															assign node6574 = (inp[14]) ? 4'b0111 : 4'b0110;
															assign node6577 = (inp[14]) ? 4'b0110 : 4'b0111;
													assign node6580 = (inp[14]) ? node6592 : node6581;
														assign node6581 = (inp[12]) ? node6587 : node6582;
															assign node6582 = (inp[7]) ? 4'b0111 : node6583;
																assign node6583 = (inp[8]) ? 4'b0111 : 4'b0110;
															assign node6587 = (inp[8]) ? node6589 : 4'b0110;
																assign node6589 = (inp[7]) ? 4'b0110 : 4'b0111;
														assign node6592 = (inp[12]) ? 4'b0111 : 4'b0110;
												assign node6595 = (inp[7]) ? node6605 : node6596;
													assign node6596 = (inp[8]) ? node6600 : node6597;
														assign node6597 = (inp[2]) ? 4'b0010 : 4'b0011;
														assign node6600 = (inp[14]) ? 4'b0011 : node6601;
															assign node6601 = (inp[2]) ? 4'b0011 : 4'b0010;
													assign node6605 = (inp[8]) ? node6611 : node6606;
														assign node6606 = (inp[2]) ? 4'b0011 : node6607;
															assign node6607 = (inp[14]) ? 4'b0011 : 4'b0010;
														assign node6611 = (inp[2]) ? 4'b0010 : node6612;
															assign node6612 = (inp[12]) ? 4'b0011 : 4'b0010;
											assign node6616 = (inp[4]) ? node6640 : node6617;
												assign node6617 = (inp[12]) ? node6625 : node6618;
													assign node6618 = (inp[8]) ? node6620 : 4'b0010;
														assign node6620 = (inp[7]) ? 4'b0010 : node6621;
															assign node6621 = (inp[2]) ? 4'b0011 : 4'b0010;
													assign node6625 = (inp[7]) ? node6633 : node6626;
														assign node6626 = (inp[8]) ? 4'b0011 : node6627;
															assign node6627 = (inp[2]) ? 4'b0010 : node6628;
																assign node6628 = (inp[14]) ? 4'b0010 : 4'b0011;
														assign node6633 = (inp[8]) ? 4'b0010 : node6634;
															assign node6634 = (inp[14]) ? 4'b0011 : node6635;
																assign node6635 = (inp[2]) ? 4'b0011 : 4'b0010;
												assign node6640 = (inp[12]) ? node6658 : node6641;
													assign node6641 = (inp[14]) ? node6651 : node6642;
														assign node6642 = (inp[8]) ? node6644 : 4'b0101;
															assign node6644 = (inp[7]) ? node6648 : node6645;
																assign node6645 = (inp[2]) ? 4'b0101 : 4'b0100;
																assign node6648 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node6651 = (inp[8]) ? node6655 : node6652;
															assign node6652 = (inp[7]) ? 4'b0101 : 4'b0100;
															assign node6655 = (inp[7]) ? 4'b0100 : 4'b0101;
													assign node6658 = (inp[2]) ? node6674 : node6659;
														assign node6659 = (inp[14]) ? node6667 : node6660;
															assign node6660 = (inp[7]) ? node6664 : node6661;
																assign node6661 = (inp[8]) ? 4'b0100 : 4'b0101;
																assign node6664 = (inp[8]) ? 4'b0101 : 4'b0100;
															assign node6667 = (inp[8]) ? node6671 : node6668;
																assign node6668 = (inp[7]) ? 4'b0101 : 4'b0100;
																assign node6671 = (inp[7]) ? 4'b0100 : 4'b0101;
														assign node6674 = (inp[14]) ? node6676 : 4'b0100;
															assign node6676 = (inp[7]) ? node6680 : node6677;
																assign node6677 = (inp[8]) ? 4'b0101 : 4'b0100;
																assign node6680 = (inp[8]) ? 4'b0100 : 4'b0101;
										assign node6683 = (inp[7]) ? node6741 : node6684;
											assign node6684 = (inp[8]) ? node6712 : node6685;
												assign node6685 = (inp[2]) ? node6703 : node6686;
													assign node6686 = (inp[14]) ? node6700 : node6687;
														assign node6687 = (inp[12]) ? node6695 : node6688;
															assign node6688 = (inp[4]) ? node6692 : node6689;
																assign node6689 = (inp[9]) ? 4'b0001 : 4'b0101;
																assign node6692 = (inp[9]) ? 4'b0101 : 4'b0001;
															assign node6695 = (inp[4]) ? node6697 : 4'b0001;
																assign node6697 = (inp[9]) ? 4'b0101 : 4'b0001;
														assign node6700 = (inp[4]) ? 4'b0100 : 4'b0000;
													assign node6703 = (inp[14]) ? 4'b0100 : node6704;
														assign node6704 = (inp[4]) ? node6708 : node6705;
															assign node6705 = (inp[9]) ? 4'b0000 : 4'b0100;
															assign node6708 = (inp[9]) ? 4'b0100 : 4'b0000;
												assign node6712 = (inp[2]) ? node6728 : node6713;
													assign node6713 = (inp[14]) ? node6721 : node6714;
														assign node6714 = (inp[12]) ? 4'b0100 : node6715;
															assign node6715 = (inp[9]) ? node6717 : 4'b0000;
																assign node6717 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node6721 = (inp[9]) ? node6725 : node6722;
															assign node6722 = (inp[4]) ? 4'b0001 : 4'b0101;
															assign node6725 = (inp[4]) ? 4'b0101 : 4'b0001;
													assign node6728 = (inp[12]) ? node6734 : node6729;
														assign node6729 = (inp[9]) ? node6731 : 4'b0101;
															assign node6731 = (inp[4]) ? 4'b0101 : 4'b0001;
														assign node6734 = (inp[4]) ? node6738 : node6735;
															assign node6735 = (inp[9]) ? 4'b0001 : 4'b0101;
															assign node6738 = (inp[9]) ? 4'b0101 : 4'b0001;
											assign node6741 = (inp[8]) ? node6771 : node6742;
												assign node6742 = (inp[2]) ? node6758 : node6743;
													assign node6743 = (inp[14]) ? node6751 : node6744;
														assign node6744 = (inp[4]) ? node6748 : node6745;
															assign node6745 = (inp[9]) ? 4'b0000 : 4'b0100;
															assign node6748 = (inp[9]) ? 4'b0100 : 4'b0000;
														assign node6751 = (inp[4]) ? node6755 : node6752;
															assign node6752 = (inp[9]) ? 4'b0001 : 4'b0101;
															assign node6755 = (inp[9]) ? 4'b0101 : 4'b0001;
													assign node6758 = (inp[14]) ? node6766 : node6759;
														assign node6759 = (inp[4]) ? node6763 : node6760;
															assign node6760 = (inp[9]) ? 4'b0001 : 4'b0101;
															assign node6763 = (inp[9]) ? 4'b0101 : 4'b0001;
														assign node6766 = (inp[12]) ? 4'b0101 : node6767;
															assign node6767 = (inp[9]) ? 4'b0101 : 4'b0001;
												assign node6771 = (inp[2]) ? node6785 : node6772;
													assign node6772 = (inp[14]) ? node6780 : node6773;
														assign node6773 = (inp[9]) ? node6777 : node6774;
															assign node6774 = (inp[4]) ? 4'b0001 : 4'b0101;
															assign node6777 = (inp[4]) ? 4'b0101 : 4'b0001;
														assign node6780 = (inp[9]) ? node6782 : 4'b0000;
															assign node6782 = (inp[4]) ? 4'b0100 : 4'b0000;
													assign node6785 = (inp[4]) ? node6789 : node6786;
														assign node6786 = (inp[9]) ? 4'b0000 : 4'b0100;
														assign node6789 = (inp[9]) ? 4'b0100 : 4'b0000;
				assign node6792 = (inp[13]) ? node10714 : node6793;
					assign node6793 = (inp[1]) ? node8725 : node6794;
						assign node6794 = (inp[3]) ? node7622 : node6795;
							assign node6795 = (inp[14]) ? node7263 : node6796;
								assign node6796 = (inp[15]) ? node7032 : node6797;
									assign node6797 = (inp[0]) ? node6917 : node6798;
										assign node6798 = (inp[4]) ? node6860 : node6799;
											assign node6799 = (inp[9]) ? node6831 : node6800;
												assign node6800 = (inp[5]) ? node6816 : node6801;
													assign node6801 = (inp[8]) ? node6809 : node6802;
														assign node6802 = (inp[7]) ? node6806 : node6803;
															assign node6803 = (inp[2]) ? 4'b0110 : 4'b0111;
															assign node6806 = (inp[2]) ? 4'b0111 : 4'b0110;
														assign node6809 = (inp[7]) ? node6813 : node6810;
															assign node6810 = (inp[2]) ? 4'b0111 : 4'b0110;
															assign node6813 = (inp[2]) ? 4'b0110 : 4'b0111;
													assign node6816 = (inp[2]) ? node6824 : node6817;
														assign node6817 = (inp[12]) ? 4'b0110 : node6818;
															assign node6818 = (inp[8]) ? 4'b0110 : node6819;
																assign node6819 = (inp[7]) ? 4'b0110 : 4'b0111;
														assign node6824 = (inp[8]) ? node6828 : node6825;
															assign node6825 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node6828 = (inp[7]) ? 4'b0110 : 4'b0111;
												assign node6831 = (inp[8]) ? node6847 : node6832;
													assign node6832 = (inp[12]) ? node6840 : node6833;
														assign node6833 = (inp[7]) ? node6837 : node6834;
															assign node6834 = (inp[2]) ? 4'b0010 : 4'b0011;
															assign node6837 = (inp[2]) ? 4'b0011 : 4'b0010;
														assign node6840 = (inp[2]) ? node6844 : node6841;
															assign node6841 = (inp[7]) ? 4'b0010 : 4'b0011;
															assign node6844 = (inp[7]) ? 4'b0011 : 4'b0010;
													assign node6847 = (inp[12]) ? node6853 : node6848;
														assign node6848 = (inp[2]) ? node6850 : 4'b0011;
															assign node6850 = (inp[7]) ? 4'b0010 : 4'b0011;
														assign node6853 = (inp[7]) ? node6857 : node6854;
															assign node6854 = (inp[2]) ? 4'b0011 : 4'b0010;
															assign node6857 = (inp[2]) ? 4'b0010 : 4'b0011;
											assign node6860 = (inp[9]) ? node6882 : node6861;
												assign node6861 = (inp[12]) ? node6869 : node6862;
													assign node6862 = (inp[2]) ? node6864 : 4'b0011;
														assign node6864 = (inp[8]) ? 4'b0010 : node6865;
															assign node6865 = (inp[7]) ? 4'b0011 : 4'b0010;
													assign node6869 = (inp[2]) ? node6875 : node6870;
														assign node6870 = (inp[8]) ? node6872 : 4'b0010;
															assign node6872 = (inp[7]) ? 4'b0011 : 4'b0010;
														assign node6875 = (inp[7]) ? node6879 : node6876;
															assign node6876 = (inp[8]) ? 4'b0011 : 4'b0010;
															assign node6879 = (inp[8]) ? 4'b0010 : 4'b0011;
												assign node6882 = (inp[5]) ? node6902 : node6883;
													assign node6883 = (inp[7]) ? node6895 : node6884;
														assign node6884 = (inp[12]) ? node6890 : node6885;
															assign node6885 = (inp[2]) ? 4'b0111 : node6886;
																assign node6886 = (inp[8]) ? 4'b0110 : 4'b0111;
															assign node6890 = (inp[8]) ? 4'b0111 : node6891;
																assign node6891 = (inp[2]) ? 4'b0110 : 4'b0111;
														assign node6895 = (inp[8]) ? node6899 : node6896;
															assign node6896 = (inp[2]) ? 4'b0111 : 4'b0110;
															assign node6899 = (inp[2]) ? 4'b0110 : 4'b0111;
													assign node6902 = (inp[12]) ? node6910 : node6903;
														assign node6903 = (inp[2]) ? node6905 : 4'b0100;
															assign node6905 = (inp[7]) ? 4'b0101 : node6906;
																assign node6906 = (inp[8]) ? 4'b0101 : 4'b0100;
														assign node6910 = (inp[2]) ? node6912 : 4'b0101;
															assign node6912 = (inp[7]) ? node6914 : 4'b0100;
																assign node6914 = (inp[8]) ? 4'b0100 : 4'b0101;
										assign node6917 = (inp[5]) ? node6973 : node6918;
											assign node6918 = (inp[7]) ? node6948 : node6919;
												assign node6919 = (inp[2]) ? node6929 : node6920;
													assign node6920 = (inp[8]) ? 4'b0000 : node6921;
														assign node6921 = (inp[4]) ? node6925 : node6922;
															assign node6922 = (inp[9]) ? 4'b0001 : 4'b0101;
															assign node6925 = (inp[9]) ? 4'b0101 : 4'b0001;
													assign node6929 = (inp[8]) ? node6937 : node6930;
														assign node6930 = (inp[4]) ? node6934 : node6931;
															assign node6931 = (inp[9]) ? 4'b0000 : 4'b0100;
															assign node6934 = (inp[9]) ? 4'b0100 : 4'b0000;
														assign node6937 = (inp[12]) ? node6943 : node6938;
															assign node6938 = (inp[4]) ? node6940 : 4'b0101;
																assign node6940 = (inp[9]) ? 4'b0101 : 4'b0001;
															assign node6943 = (inp[9]) ? 4'b0001 : node6944;
																assign node6944 = (inp[4]) ? 4'b0001 : 4'b0101;
												assign node6948 = (inp[2]) ? node6960 : node6949;
													assign node6949 = (inp[8]) ? node6955 : node6950;
														assign node6950 = (inp[4]) ? node6952 : 4'b0100;
															assign node6952 = (inp[12]) ? 4'b0000 : 4'b0100;
														assign node6955 = (inp[9]) ? node6957 : 4'b0101;
															assign node6957 = (inp[4]) ? 4'b0101 : 4'b0001;
													assign node6960 = (inp[8]) ? node6968 : node6961;
														assign node6961 = (inp[4]) ? node6965 : node6962;
															assign node6962 = (inp[9]) ? 4'b0001 : 4'b0101;
															assign node6965 = (inp[9]) ? 4'b0101 : 4'b0001;
														assign node6968 = (inp[4]) ? 4'b0100 : node6969;
															assign node6969 = (inp[9]) ? 4'b0000 : 4'b0100;
											assign node6973 = (inp[4]) ? node7007 : node6974;
												assign node6974 = (inp[9]) ? node6994 : node6975;
													assign node6975 = (inp[12]) ? node6989 : node6976;
														assign node6976 = (inp[2]) ? node6982 : node6977;
															assign node6977 = (inp[8]) ? node6979 : 4'b0100;
																assign node6979 = (inp[7]) ? 4'b0101 : 4'b0100;
															assign node6982 = (inp[7]) ? node6986 : node6983;
																assign node6983 = (inp[8]) ? 4'b0101 : 4'b0100;
																assign node6986 = (inp[8]) ? 4'b0100 : 4'b0101;
														assign node6989 = (inp[7]) ? node6991 : 4'b0101;
															assign node6991 = (inp[2]) ? 4'b0101 : 4'b0100;
													assign node6994 = (inp[7]) ? node7000 : node6995;
														assign node6995 = (inp[2]) ? 4'b0000 : node6996;
															assign node6996 = (inp[8]) ? 4'b0000 : 4'b0001;
														assign node7000 = (inp[8]) ? node7004 : node7001;
															assign node7001 = (inp[2]) ? 4'b0001 : 4'b0000;
															assign node7004 = (inp[2]) ? 4'b0000 : 4'b0001;
												assign node7007 = (inp[9]) ? node7019 : node7008;
													assign node7008 = (inp[8]) ? node7014 : node7009;
														assign node7009 = (inp[2]) ? 4'b0000 : node7010;
															assign node7010 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node7014 = (inp[7]) ? 4'b0001 : node7015;
															assign node7015 = (inp[2]) ? 4'b0001 : 4'b0000;
													assign node7019 = (inp[2]) ? node7027 : node7020;
														assign node7020 = (inp[7]) ? node7024 : node7021;
															assign node7021 = (inp[8]) ? 4'b0110 : 4'b0111;
															assign node7024 = (inp[8]) ? 4'b0111 : 4'b0110;
														assign node7027 = (inp[8]) ? 4'b0110 : node7028;
															assign node7028 = (inp[7]) ? 4'b0111 : 4'b0110;
									assign node7032 = (inp[0]) ? node7158 : node7033;
										assign node7033 = (inp[4]) ? node7095 : node7034;
											assign node7034 = (inp[9]) ? node7058 : node7035;
												assign node7035 = (inp[7]) ? node7043 : node7036;
													assign node7036 = (inp[5]) ? node7038 : 4'b0100;
														assign node7038 = (inp[2]) ? node7040 : 4'b0100;
															assign node7040 = (inp[8]) ? 4'b0101 : 4'b0100;
													assign node7043 = (inp[5]) ? node7051 : node7044;
														assign node7044 = (inp[2]) ? node7048 : node7045;
															assign node7045 = (inp[8]) ? 4'b0101 : 4'b0100;
															assign node7048 = (inp[8]) ? 4'b0100 : 4'b0101;
														assign node7051 = (inp[2]) ? node7055 : node7052;
															assign node7052 = (inp[8]) ? 4'b0101 : 4'b0100;
															assign node7055 = (inp[8]) ? 4'b0100 : 4'b0101;
												assign node7058 = (inp[5]) ? node7072 : node7059;
													assign node7059 = (inp[8]) ? node7065 : node7060;
														assign node7060 = (inp[2]) ? 4'b0000 : node7061;
															assign node7061 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node7065 = (inp[7]) ? node7069 : node7066;
															assign node7066 = (inp[2]) ? 4'b0001 : 4'b0000;
															assign node7069 = (inp[2]) ? 4'b0000 : 4'b0001;
													assign node7072 = (inp[8]) ? node7084 : node7073;
														assign node7073 = (inp[12]) ? node7079 : node7074;
															assign node7074 = (inp[2]) ? 4'b0001 : node7075;
																assign node7075 = (inp[7]) ? 4'b0000 : 4'b0001;
															assign node7079 = (inp[7]) ? 4'b0001 : node7080;
																assign node7080 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node7084 = (inp[12]) ? node7090 : node7085;
															assign node7085 = (inp[7]) ? node7087 : 4'b0000;
																assign node7087 = (inp[2]) ? 4'b0000 : 4'b0001;
															assign node7090 = (inp[7]) ? 4'b0000 : node7091;
																assign node7091 = (inp[2]) ? 4'b0001 : 4'b0000;
											assign node7095 = (inp[9]) ? node7127 : node7096;
												assign node7096 = (inp[12]) ? node7112 : node7097;
													assign node7097 = (inp[8]) ? node7105 : node7098;
														assign node7098 = (inp[2]) ? node7102 : node7099;
															assign node7099 = (inp[7]) ? 4'b0000 : 4'b0001;
															assign node7102 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node7105 = (inp[7]) ? node7109 : node7106;
															assign node7106 = (inp[2]) ? 4'b0001 : 4'b0000;
															assign node7109 = (inp[2]) ? 4'b0000 : 4'b0001;
													assign node7112 = (inp[2]) ? node7114 : 4'b0001;
														assign node7114 = (inp[5]) ? node7120 : node7115;
															assign node7115 = (inp[8]) ? 4'b0001 : node7116;
																assign node7116 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node7120 = (inp[8]) ? node7124 : node7121;
																assign node7121 = (inp[7]) ? 4'b0001 : 4'b0000;
																assign node7124 = (inp[7]) ? 4'b0000 : 4'b0001;
												assign node7127 = (inp[5]) ? node7147 : node7128;
													assign node7128 = (inp[2]) ? node7134 : node7129;
														assign node7129 = (inp[7]) ? 4'b0100 : node7130;
															assign node7130 = (inp[8]) ? 4'b0100 : 4'b0101;
														assign node7134 = (inp[12]) ? node7140 : node7135;
															assign node7135 = (inp[7]) ? 4'b0101 : node7136;
																assign node7136 = (inp[8]) ? 4'b0101 : 4'b0100;
															assign node7140 = (inp[7]) ? node7144 : node7141;
																assign node7141 = (inp[8]) ? 4'b0101 : 4'b0100;
																assign node7144 = (inp[8]) ? 4'b0100 : 4'b0101;
													assign node7147 = (inp[2]) ? node7153 : node7148;
														assign node7148 = (inp[8]) ? 4'b0110 : node7149;
															assign node7149 = (inp[7]) ? 4'b0110 : 4'b0111;
														assign node7153 = (inp[8]) ? 4'b0111 : node7154;
															assign node7154 = (inp[7]) ? 4'b0111 : 4'b0110;
										assign node7158 = (inp[9]) ? node7214 : node7159;
											assign node7159 = (inp[4]) ? node7173 : node7160;
												assign node7160 = (inp[7]) ? node7168 : node7161;
													assign node7161 = (inp[2]) ? node7165 : node7162;
														assign node7162 = (inp[8]) ? 4'b0110 : 4'b0111;
														assign node7165 = (inp[8]) ? 4'b0111 : 4'b0110;
													assign node7168 = (inp[8]) ? node7170 : 4'b0111;
														assign node7170 = (inp[2]) ? 4'b0110 : 4'b0111;
												assign node7173 = (inp[7]) ? node7193 : node7174;
													assign node7174 = (inp[5]) ? node7188 : node7175;
														assign node7175 = (inp[12]) ? node7183 : node7176;
															assign node7176 = (inp[2]) ? node7180 : node7177;
																assign node7177 = (inp[8]) ? 4'b0010 : 4'b0011;
																assign node7180 = (inp[8]) ? 4'b0011 : 4'b0010;
															assign node7183 = (inp[8]) ? 4'b0010 : node7184;
																assign node7184 = (inp[2]) ? 4'b0010 : 4'b0011;
														assign node7188 = (inp[8]) ? node7190 : 4'b0011;
															assign node7190 = (inp[2]) ? 4'b0011 : 4'b0010;
													assign node7193 = (inp[5]) ? node7205 : node7194;
														assign node7194 = (inp[12]) ? node7200 : node7195;
															assign node7195 = (inp[2]) ? node7197 : 4'b0010;
																assign node7197 = (inp[8]) ? 4'b0010 : 4'b0011;
															assign node7200 = (inp[2]) ? 4'b0010 : node7201;
																assign node7201 = (inp[8]) ? 4'b0011 : 4'b0010;
														assign node7205 = (inp[12]) ? node7209 : node7206;
															assign node7206 = (inp[2]) ? 4'b0011 : 4'b0010;
															assign node7209 = (inp[8]) ? node7211 : 4'b0010;
																assign node7211 = (inp[2]) ? 4'b0010 : 4'b0011;
											assign node7214 = (inp[4]) ? node7232 : node7215;
												assign node7215 = (inp[2]) ? node7223 : node7216;
													assign node7216 = (inp[7]) ? node7220 : node7217;
														assign node7217 = (inp[8]) ? 4'b0010 : 4'b0011;
														assign node7220 = (inp[8]) ? 4'b0011 : 4'b0010;
													assign node7223 = (inp[12]) ? node7227 : node7224;
														assign node7224 = (inp[8]) ? 4'b0010 : 4'b0011;
														assign node7227 = (inp[8]) ? 4'b0011 : node7228;
															assign node7228 = (inp[7]) ? 4'b0011 : 4'b0010;
												assign node7232 = (inp[5]) ? node7248 : node7233;
													assign node7233 = (inp[8]) ? node7241 : node7234;
														assign node7234 = (inp[2]) ? node7238 : node7235;
															assign node7235 = (inp[7]) ? 4'b0110 : 4'b0111;
															assign node7238 = (inp[7]) ? 4'b0111 : 4'b0110;
														assign node7241 = (inp[2]) ? node7245 : node7242;
															assign node7242 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node7245 = (inp[7]) ? 4'b0110 : 4'b0111;
													assign node7248 = (inp[12]) ? node7258 : node7249;
														assign node7249 = (inp[8]) ? node7251 : 4'b0100;
															assign node7251 = (inp[7]) ? node7255 : node7252;
																assign node7252 = (inp[2]) ? 4'b0101 : 4'b0100;
																assign node7255 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node7258 = (inp[2]) ? 4'b0101 : node7259;
															assign node7259 = (inp[7]) ? 4'b0100 : 4'b0101;
								assign node7263 = (inp[0]) ? node7397 : node7264;
									assign node7264 = (inp[15]) ? node7334 : node7265;
										assign node7265 = (inp[9]) ? node7295 : node7266;
											assign node7266 = (inp[4]) ? node7280 : node7267;
												assign node7267 = (inp[12]) ? node7273 : node7268;
													assign node7268 = (inp[8]) ? 4'b0111 : node7269;
														assign node7269 = (inp[7]) ? 4'b0111 : 4'b0110;
													assign node7273 = (inp[8]) ? node7277 : node7274;
														assign node7274 = (inp[7]) ? 4'b0111 : 4'b0110;
														assign node7277 = (inp[7]) ? 4'b0110 : 4'b0111;
												assign node7280 = (inp[2]) ? node7288 : node7281;
													assign node7281 = (inp[12]) ? node7283 : 4'b0010;
														assign node7283 = (inp[7]) ? node7285 : 4'b0011;
															assign node7285 = (inp[8]) ? 4'b0010 : 4'b0011;
													assign node7288 = (inp[8]) ? node7292 : node7289;
														assign node7289 = (inp[7]) ? 4'b0011 : 4'b0010;
														assign node7292 = (inp[7]) ? 4'b0010 : 4'b0011;
											assign node7295 = (inp[4]) ? node7303 : node7296;
												assign node7296 = (inp[7]) ? node7300 : node7297;
													assign node7297 = (inp[8]) ? 4'b0011 : 4'b0010;
													assign node7300 = (inp[8]) ? 4'b0010 : 4'b0011;
												assign node7303 = (inp[5]) ? node7323 : node7304;
													assign node7304 = (inp[12]) ? node7312 : node7305;
														assign node7305 = (inp[2]) ? 4'b0111 : node7306;
															assign node7306 = (inp[7]) ? node7308 : 4'b0110;
																assign node7308 = (inp[8]) ? 4'b0110 : 4'b0111;
														assign node7312 = (inp[2]) ? node7318 : node7313;
															assign node7313 = (inp[8]) ? 4'b0111 : node7314;
																assign node7314 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node7318 = (inp[8]) ? node7320 : 4'b0110;
																assign node7320 = (inp[7]) ? 4'b0110 : 4'b0111;
													assign node7323 = (inp[2]) ? node7329 : node7324;
														assign node7324 = (inp[8]) ? 4'b0101 : node7325;
															assign node7325 = (inp[7]) ? 4'b0101 : 4'b0100;
														assign node7329 = (inp[8]) ? node7331 : 4'b0101;
															assign node7331 = (inp[7]) ? 4'b0100 : 4'b0101;
										assign node7334 = (inp[9]) ? node7362 : node7335;
											assign node7335 = (inp[4]) ? node7343 : node7336;
												assign node7336 = (inp[8]) ? node7340 : node7337;
													assign node7337 = (inp[7]) ? 4'b0101 : 4'b0100;
													assign node7340 = (inp[7]) ? 4'b0100 : 4'b0101;
												assign node7343 = (inp[12]) ? node7355 : node7344;
													assign node7344 = (inp[2]) ? node7350 : node7345;
														assign node7345 = (inp[8]) ? node7347 : 4'b0001;
															assign node7347 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node7350 = (inp[8]) ? node7352 : 4'b0000;
															assign node7352 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node7355 = (inp[8]) ? node7359 : node7356;
														assign node7356 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node7359 = (inp[7]) ? 4'b0000 : 4'b0001;
											assign node7362 = (inp[4]) ? node7370 : node7363;
												assign node7363 = (inp[8]) ? node7367 : node7364;
													assign node7364 = (inp[7]) ? 4'b0001 : 4'b0000;
													assign node7367 = (inp[7]) ? 4'b0000 : 4'b0001;
												assign node7370 = (inp[5]) ? node7378 : node7371;
													assign node7371 = (inp[7]) ? node7375 : node7372;
														assign node7372 = (inp[8]) ? 4'b0101 : 4'b0100;
														assign node7375 = (inp[8]) ? 4'b0100 : 4'b0101;
													assign node7378 = (inp[2]) ? node7386 : node7379;
														assign node7379 = (inp[8]) ? node7383 : node7380;
															assign node7380 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node7383 = (inp[7]) ? 4'b0110 : 4'b0111;
														assign node7386 = (inp[12]) ? node7392 : node7387;
															assign node7387 = (inp[7]) ? 4'b0111 : node7388;
																assign node7388 = (inp[8]) ? 4'b0111 : 4'b0110;
															assign node7392 = (inp[8]) ? node7394 : 4'b0111;
																assign node7394 = (inp[7]) ? 4'b0110 : 4'b0111;
									assign node7397 = (inp[15]) ? node7499 : node7398;
										assign node7398 = (inp[5]) ? node7462 : node7399;
											assign node7399 = (inp[12]) ? node7431 : node7400;
												assign node7400 = (inp[2]) ? node7416 : node7401;
													assign node7401 = (inp[4]) ? node7411 : node7402;
														assign node7402 = (inp[9]) ? node7406 : node7403;
															assign node7403 = (inp[7]) ? 4'b0100 : 4'b0101;
															assign node7406 = (inp[8]) ? 4'b0000 : node7407;
																assign node7407 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node7411 = (inp[9]) ? node7413 : 4'b0001;
															assign node7413 = (inp[7]) ? 4'b0101 : 4'b0100;
													assign node7416 = (inp[7]) ? node7428 : node7417;
														assign node7417 = (inp[8]) ? node7423 : node7418;
															assign node7418 = (inp[4]) ? node7420 : 4'b0000;
																assign node7420 = (inp[9]) ? 4'b0100 : 4'b0000;
															assign node7423 = (inp[4]) ? node7425 : 4'b0001;
																assign node7425 = (inp[9]) ? 4'b0101 : 4'b0001;
														assign node7428 = (inp[8]) ? 4'b0000 : 4'b0001;
												assign node7431 = (inp[4]) ? node7447 : node7432;
													assign node7432 = (inp[9]) ? node7438 : node7433;
														assign node7433 = (inp[7]) ? 4'b0100 : node7434;
															assign node7434 = (inp[8]) ? 4'b0101 : 4'b0100;
														assign node7438 = (inp[2]) ? node7442 : node7439;
															assign node7439 = (inp[8]) ? 4'b0000 : 4'b0001;
															assign node7442 = (inp[7]) ? 4'b0000 : node7443;
																assign node7443 = (inp[8]) ? 4'b0001 : 4'b0000;
													assign node7447 = (inp[9]) ? node7455 : node7448;
														assign node7448 = (inp[8]) ? node7452 : node7449;
															assign node7449 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node7452 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node7455 = (inp[8]) ? node7459 : node7456;
															assign node7456 = (inp[7]) ? 4'b0101 : 4'b0100;
															assign node7459 = (inp[7]) ? 4'b0100 : 4'b0101;
											assign node7462 = (inp[4]) ? node7478 : node7463;
												assign node7463 = (inp[9]) ? node7471 : node7464;
													assign node7464 = (inp[8]) ? node7468 : node7465;
														assign node7465 = (inp[7]) ? 4'b0101 : 4'b0100;
														assign node7468 = (inp[7]) ? 4'b0100 : 4'b0101;
													assign node7471 = (inp[8]) ? node7475 : node7472;
														assign node7472 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node7475 = (inp[7]) ? 4'b0000 : 4'b0001;
												assign node7478 = (inp[9]) ? node7486 : node7479;
													assign node7479 = (inp[7]) ? node7483 : node7480;
														assign node7480 = (inp[8]) ? 4'b0001 : 4'b0000;
														assign node7483 = (inp[8]) ? 4'b0000 : 4'b0001;
													assign node7486 = (inp[12]) ? node7492 : node7487;
														assign node7487 = (inp[8]) ? 4'b0110 : node7488;
															assign node7488 = (inp[7]) ? 4'b0111 : 4'b0110;
														assign node7492 = (inp[2]) ? 4'b0111 : node7493;
															assign node7493 = (inp[7]) ? 4'b0110 : node7494;
																assign node7494 = (inp[8]) ? 4'b0111 : 4'b0110;
										assign node7499 = (inp[5]) ? node7573 : node7500;
											assign node7500 = (inp[12]) ? node7532 : node7501;
												assign node7501 = (inp[9]) ? node7517 : node7502;
													assign node7502 = (inp[4]) ? node7510 : node7503;
														assign node7503 = (inp[8]) ? node7507 : node7504;
															assign node7504 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node7507 = (inp[7]) ? 4'b0110 : 4'b0111;
														assign node7510 = (inp[8]) ? node7514 : node7511;
															assign node7511 = (inp[7]) ? 4'b0011 : 4'b0010;
															assign node7514 = (inp[7]) ? 4'b0010 : 4'b0011;
													assign node7517 = (inp[4]) ? node7523 : node7518;
														assign node7518 = (inp[8]) ? node7520 : 4'b0011;
															assign node7520 = (inp[7]) ? 4'b0010 : 4'b0011;
														assign node7523 = (inp[2]) ? node7525 : 4'b0111;
															assign node7525 = (inp[7]) ? node7529 : node7526;
																assign node7526 = (inp[8]) ? 4'b0111 : 4'b0110;
																assign node7529 = (inp[8]) ? 4'b0110 : 4'b0111;
												assign node7532 = (inp[2]) ? node7552 : node7533;
													assign node7533 = (inp[9]) ? node7541 : node7534;
														assign node7534 = (inp[8]) ? node7538 : node7535;
															assign node7535 = (inp[7]) ? 4'b0011 : 4'b0010;
															assign node7538 = (inp[7]) ? 4'b0010 : 4'b0011;
														assign node7541 = (inp[4]) ? node7549 : node7542;
															assign node7542 = (inp[8]) ? node7546 : node7543;
																assign node7543 = (inp[7]) ? 4'b0011 : 4'b0010;
																assign node7546 = (inp[7]) ? 4'b0010 : 4'b0011;
															assign node7549 = (inp[8]) ? 4'b0110 : 4'b0111;
													assign node7552 = (inp[7]) ? node7562 : node7553;
														assign node7553 = (inp[8]) ? 4'b0111 : node7554;
															assign node7554 = (inp[4]) ? node7558 : node7555;
																assign node7555 = (inp[9]) ? 4'b0010 : 4'b0110;
																assign node7558 = (inp[9]) ? 4'b0110 : 4'b0010;
														assign node7562 = (inp[8]) ? node7568 : node7563;
															assign node7563 = (inp[9]) ? 4'b0011 : node7564;
																assign node7564 = (inp[4]) ? 4'b0011 : 4'b0111;
															assign node7568 = (inp[9]) ? 4'b0010 : node7569;
																assign node7569 = (inp[4]) ? 4'b0010 : 4'b0110;
											assign node7573 = (inp[9]) ? node7599 : node7574;
												assign node7574 = (inp[4]) ? node7584 : node7575;
													assign node7575 = (inp[2]) ? 4'b0111 : node7576;
														assign node7576 = (inp[12]) ? node7580 : node7577;
															assign node7577 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node7580 = (inp[7]) ? 4'b0110 : 4'b0111;
													assign node7584 = (inp[12]) ? node7592 : node7585;
														assign node7585 = (inp[7]) ? node7589 : node7586;
															assign node7586 = (inp[8]) ? 4'b0011 : 4'b0010;
															assign node7589 = (inp[8]) ? 4'b0010 : 4'b0011;
														assign node7592 = (inp[7]) ? node7596 : node7593;
															assign node7593 = (inp[8]) ? 4'b0011 : 4'b0010;
															assign node7596 = (inp[8]) ? 4'b0010 : 4'b0011;
												assign node7599 = (inp[4]) ? node7615 : node7600;
													assign node7600 = (inp[12]) ? node7606 : node7601;
														assign node7601 = (inp[8]) ? 4'b0011 : node7602;
															assign node7602 = (inp[7]) ? 4'b0011 : 4'b0010;
														assign node7606 = (inp[2]) ? 4'b0010 : node7607;
															assign node7607 = (inp[8]) ? node7611 : node7608;
																assign node7608 = (inp[7]) ? 4'b0011 : 4'b0010;
																assign node7611 = (inp[7]) ? 4'b0010 : 4'b0011;
													assign node7615 = (inp[7]) ? node7619 : node7616;
														assign node7616 = (inp[8]) ? 4'b0101 : 4'b0100;
														assign node7619 = (inp[8]) ? 4'b0100 : 4'b0101;
							assign node7622 = (inp[12]) ? node8162 : node7623;
								assign node7623 = (inp[5]) ? node7893 : node7624;
									assign node7624 = (inp[4]) ? node7762 : node7625;
										assign node7625 = (inp[9]) ? node7699 : node7626;
											assign node7626 = (inp[8]) ? node7670 : node7627;
												assign node7627 = (inp[7]) ? node7651 : node7628;
													assign node7628 = (inp[14]) ? node7642 : node7629;
														assign node7629 = (inp[2]) ? node7637 : node7630;
															assign node7630 = (inp[15]) ? node7634 : node7631;
																assign node7631 = (inp[0]) ? 4'b0101 : 4'b0111;
																assign node7634 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node7637 = (inp[0]) ? 4'b0110 : node7638;
																assign node7638 = (inp[15]) ? 4'b0100 : 4'b0110;
														assign node7642 = (inp[2]) ? 4'b0110 : node7643;
															assign node7643 = (inp[0]) ? node7647 : node7644;
																assign node7644 = (inp[15]) ? 4'b0100 : 4'b0110;
																assign node7647 = (inp[15]) ? 4'b0110 : 4'b0100;
													assign node7651 = (inp[2]) ? node7663 : node7652;
														assign node7652 = (inp[14]) ? node7660 : node7653;
															assign node7653 = (inp[15]) ? node7657 : node7654;
																assign node7654 = (inp[0]) ? 4'b0100 : 4'b0110;
																assign node7657 = (inp[0]) ? 4'b0110 : 4'b0100;
															assign node7660 = (inp[15]) ? 4'b0111 : 4'b0101;
														assign node7663 = (inp[15]) ? node7667 : node7664;
															assign node7664 = (inp[0]) ? 4'b0101 : 4'b0111;
															assign node7667 = (inp[0]) ? 4'b0111 : 4'b0101;
												assign node7670 = (inp[7]) ? node7688 : node7671;
													assign node7671 = (inp[14]) ? node7683 : node7672;
														assign node7672 = (inp[2]) ? node7680 : node7673;
															assign node7673 = (inp[0]) ? node7677 : node7674;
																assign node7674 = (inp[15]) ? 4'b0100 : 4'b0110;
																assign node7677 = (inp[15]) ? 4'b0110 : 4'b0100;
															assign node7680 = (inp[0]) ? 4'b0101 : 4'b0111;
														assign node7683 = (inp[15]) ? 4'b0101 : node7684;
															assign node7684 = (inp[0]) ? 4'b0101 : 4'b0111;
													assign node7688 = (inp[14]) ? node7692 : node7689;
														assign node7689 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node7692 = (inp[15]) ? node7696 : node7693;
															assign node7693 = (inp[0]) ? 4'b0100 : 4'b0110;
															assign node7696 = (inp[0]) ? 4'b0110 : 4'b0100;
											assign node7699 = (inp[8]) ? node7733 : node7700;
												assign node7700 = (inp[7]) ? node7724 : node7701;
													assign node7701 = (inp[2]) ? node7715 : node7702;
														assign node7702 = (inp[14]) ? node7708 : node7703;
															assign node7703 = (inp[15]) ? 4'b0011 : node7704;
																assign node7704 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node7708 = (inp[15]) ? node7712 : node7709;
																assign node7709 = (inp[0]) ? 4'b0000 : 4'b0010;
																assign node7712 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node7715 = (inp[14]) ? 4'b0000 : node7716;
															assign node7716 = (inp[0]) ? node7720 : node7717;
																assign node7717 = (inp[15]) ? 4'b0000 : 4'b0010;
																assign node7720 = (inp[15]) ? 4'b0010 : 4'b0000;
													assign node7724 = (inp[14]) ? 4'b0001 : node7725;
														assign node7725 = (inp[2]) ? 4'b0001 : node7726;
															assign node7726 = (inp[15]) ? node7728 : 4'b0000;
																assign node7728 = (inp[0]) ? 4'b0010 : 4'b0000;
												assign node7733 = (inp[7]) ? node7745 : node7734;
													assign node7734 = (inp[2]) ? node7740 : node7735;
														assign node7735 = (inp[14]) ? node7737 : 4'b0000;
															assign node7737 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node7740 = (inp[15]) ? node7742 : 4'b0011;
															assign node7742 = (inp[0]) ? 4'b0011 : 4'b0001;
													assign node7745 = (inp[2]) ? node7753 : node7746;
														assign node7746 = (inp[14]) ? node7748 : 4'b0011;
															assign node7748 = (inp[0]) ? 4'b0000 : node7749;
																assign node7749 = (inp[15]) ? 4'b0000 : 4'b0010;
														assign node7753 = (inp[14]) ? 4'b0010 : node7754;
															assign node7754 = (inp[15]) ? node7758 : node7755;
																assign node7755 = (inp[0]) ? 4'b0000 : 4'b0010;
																assign node7758 = (inp[0]) ? 4'b0010 : 4'b0000;
										assign node7762 = (inp[9]) ? node7840 : node7763;
											assign node7763 = (inp[8]) ? node7805 : node7764;
												assign node7764 = (inp[7]) ? node7782 : node7765;
													assign node7765 = (inp[2]) ? node7775 : node7766;
														assign node7766 = (inp[14]) ? 4'b0000 : node7767;
															assign node7767 = (inp[15]) ? node7771 : node7768;
																assign node7768 = (inp[0]) ? 4'b0001 : 4'b0011;
																assign node7771 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node7775 = (inp[15]) ? node7779 : node7776;
															assign node7776 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node7779 = (inp[0]) ? 4'b0010 : 4'b0000;
													assign node7782 = (inp[2]) ? node7792 : node7783;
														assign node7783 = (inp[14]) ? node7789 : node7784;
															assign node7784 = (inp[0]) ? 4'b0000 : node7785;
																assign node7785 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node7789 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node7792 = (inp[14]) ? node7798 : node7793;
															assign node7793 = (inp[15]) ? node7795 : 4'b0001;
																assign node7795 = (inp[0]) ? 4'b0011 : 4'b0001;
															assign node7798 = (inp[0]) ? node7802 : node7799;
																assign node7799 = (inp[15]) ? 4'b0001 : 4'b0011;
																assign node7802 = (inp[15]) ? 4'b0011 : 4'b0001;
												assign node7805 = (inp[7]) ? node7821 : node7806;
													assign node7806 = (inp[14]) ? node7814 : node7807;
														assign node7807 = (inp[2]) ? 4'b0001 : node7808;
															assign node7808 = (inp[15]) ? 4'b0010 : node7809;
																assign node7809 = (inp[0]) ? 4'b0000 : 4'b0010;
														assign node7814 = (inp[0]) ? node7818 : node7815;
															assign node7815 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node7818 = (inp[15]) ? 4'b0011 : 4'b0001;
													assign node7821 = (inp[14]) ? node7827 : node7822;
														assign node7822 = (inp[2]) ? 4'b0010 : node7823;
															assign node7823 = (inp[15]) ? 4'b0001 : 4'b0011;
														assign node7827 = (inp[2]) ? node7833 : node7828;
															assign node7828 = (inp[0]) ? node7830 : 4'b0000;
																assign node7830 = (inp[15]) ? 4'b0010 : 4'b0000;
															assign node7833 = (inp[0]) ? node7837 : node7834;
																assign node7834 = (inp[15]) ? 4'b0000 : 4'b0010;
																assign node7837 = (inp[15]) ? 4'b0010 : 4'b0000;
											assign node7840 = (inp[14]) ? node7870 : node7841;
												assign node7841 = (inp[7]) ? node7855 : node7842;
													assign node7842 = (inp[2]) ? node7852 : node7843;
														assign node7843 = (inp[8]) ? node7849 : node7844;
															assign node7844 = (inp[0]) ? node7846 : 4'b0101;
																assign node7846 = (inp[15]) ? 4'b0101 : 4'b0111;
															assign node7849 = (inp[15]) ? 4'b0100 : 4'b0110;
														assign node7852 = (inp[8]) ? 4'b0111 : 4'b0110;
													assign node7855 = (inp[0]) ? node7867 : node7856;
														assign node7856 = (inp[15]) ? node7860 : node7857;
															assign node7857 = (inp[8]) ? 4'b0100 : 4'b0101;
															assign node7860 = (inp[8]) ? node7864 : node7861;
																assign node7861 = (inp[2]) ? 4'b0111 : 4'b0110;
																assign node7864 = (inp[2]) ? 4'b0110 : 4'b0111;
														assign node7867 = (inp[15]) ? 4'b0101 : 4'b0111;
												assign node7870 = (inp[8]) ? node7880 : node7871;
													assign node7871 = (inp[7]) ? 4'b0101 : node7872;
														assign node7872 = (inp[2]) ? node7874 : 4'b0100;
															assign node7874 = (inp[15]) ? node7876 : 4'b0110;
																assign node7876 = (inp[0]) ? 4'b0100 : 4'b0110;
													assign node7880 = (inp[7]) ? node7888 : node7881;
														assign node7881 = (inp[0]) ? node7885 : node7882;
															assign node7882 = (inp[15]) ? 4'b0111 : 4'b0101;
															assign node7885 = (inp[15]) ? 4'b0101 : 4'b0111;
														assign node7888 = (inp[15]) ? node7890 : 4'b0110;
															assign node7890 = (inp[0]) ? 4'b0100 : 4'b0110;
									assign node7893 = (inp[0]) ? node8021 : node7894;
										assign node7894 = (inp[15]) ? node7968 : node7895;
											assign node7895 = (inp[8]) ? node7941 : node7896;
												assign node7896 = (inp[7]) ? node7922 : node7897;
													assign node7897 = (inp[14]) ? node7913 : node7898;
														assign node7898 = (inp[2]) ? node7906 : node7899;
															assign node7899 = (inp[4]) ? node7903 : node7900;
																assign node7900 = (inp[9]) ? 4'b0001 : 4'b0101;
																assign node7903 = (inp[9]) ? 4'b0101 : 4'b0001;
															assign node7906 = (inp[4]) ? node7910 : node7907;
																assign node7907 = (inp[9]) ? 4'b0000 : 4'b0100;
																assign node7910 = (inp[9]) ? 4'b0100 : 4'b0000;
														assign node7913 = (inp[2]) ? 4'b0000 : node7914;
															assign node7914 = (inp[9]) ? node7918 : node7915;
																assign node7915 = (inp[4]) ? 4'b0000 : 4'b0100;
																assign node7918 = (inp[4]) ? 4'b0100 : 4'b0000;
													assign node7922 = (inp[14]) ? node7932 : node7923;
														assign node7923 = (inp[2]) ? node7927 : node7924;
															assign node7924 = (inp[4]) ? 4'b0100 : 4'b0000;
															assign node7927 = (inp[9]) ? node7929 : 4'b0001;
																assign node7929 = (inp[4]) ? 4'b0101 : 4'b0001;
														assign node7932 = (inp[2]) ? 4'b0101 : node7933;
															assign node7933 = (inp[9]) ? node7937 : node7934;
																assign node7934 = (inp[4]) ? 4'b0001 : 4'b0101;
																assign node7937 = (inp[4]) ? 4'b0101 : 4'b0001;
												assign node7941 = (inp[7]) ? node7957 : node7942;
													assign node7942 = (inp[2]) ? node7950 : node7943;
														assign node7943 = (inp[14]) ? 4'b0001 : node7944;
															assign node7944 = (inp[9]) ? 4'b0000 : node7945;
																assign node7945 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node7950 = (inp[4]) ? node7954 : node7951;
															assign node7951 = (inp[9]) ? 4'b0001 : 4'b0101;
															assign node7954 = (inp[14]) ? 4'b0101 : 4'b0001;
													assign node7957 = (inp[4]) ? node7965 : node7958;
														assign node7958 = (inp[9]) ? node7960 : 4'b0100;
															assign node7960 = (inp[14]) ? 4'b0000 : node7961;
																assign node7961 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node7965 = (inp[9]) ? 4'b0100 : 4'b0000;
											assign node7968 = (inp[7]) ? node7994 : node7969;
												assign node7969 = (inp[8]) ? node7983 : node7970;
													assign node7970 = (inp[14]) ? node7978 : node7971;
														assign node7971 = (inp[2]) ? node7973 : 4'b0111;
															assign node7973 = (inp[4]) ? 4'b0010 : node7974;
																assign node7974 = (inp[9]) ? 4'b0010 : 4'b0110;
														assign node7978 = (inp[9]) ? node7980 : 4'b0010;
															assign node7980 = (inp[4]) ? 4'b0110 : 4'b0010;
													assign node7983 = (inp[4]) ? node7989 : node7984;
														assign node7984 = (inp[9]) ? node7986 : 4'b0111;
															assign node7986 = (inp[14]) ? 4'b0011 : 4'b0010;
														assign node7989 = (inp[14]) ? 4'b0011 : node7990;
															assign node7990 = (inp[2]) ? 4'b0011 : 4'b0010;
												assign node7994 = (inp[8]) ? node8006 : node7995;
													assign node7995 = (inp[2]) ? node7999 : node7996;
														assign node7996 = (inp[14]) ? 4'b0011 : 4'b0010;
														assign node7999 = (inp[9]) ? node8003 : node8000;
															assign node8000 = (inp[4]) ? 4'b0011 : 4'b0111;
															assign node8003 = (inp[4]) ? 4'b0111 : 4'b0011;
													assign node8006 = (inp[14]) ? node8016 : node8007;
														assign node8007 = (inp[2]) ? node8011 : node8008;
															assign node8008 = (inp[9]) ? 4'b0011 : 4'b0111;
															assign node8011 = (inp[9]) ? 4'b0110 : node8012;
																assign node8012 = (inp[4]) ? 4'b0010 : 4'b0110;
														assign node8016 = (inp[9]) ? 4'b0010 : node8017;
															assign node8017 = (inp[4]) ? 4'b0010 : 4'b0110;
										assign node8021 = (inp[15]) ? node8083 : node8022;
											assign node8022 = (inp[2]) ? node8056 : node8023;
												assign node8023 = (inp[14]) ? node8043 : node8024;
													assign node8024 = (inp[8]) ? node8032 : node8025;
														assign node8025 = (inp[7]) ? node8027 : 4'b0111;
															assign node8027 = (inp[4]) ? 4'b0110 : node8028;
																assign node8028 = (inp[9]) ? 4'b0010 : 4'b0110;
														assign node8032 = (inp[7]) ? node8036 : node8033;
															assign node8033 = (inp[9]) ? 4'b0110 : 4'b0010;
															assign node8036 = (inp[4]) ? node8040 : node8037;
																assign node8037 = (inp[9]) ? 4'b0011 : 4'b0111;
																assign node8040 = (inp[9]) ? 4'b0111 : 4'b0011;
													assign node8043 = (inp[9]) ? node8053 : node8044;
														assign node8044 = (inp[4]) ? node8046 : 4'b0111;
															assign node8046 = (inp[7]) ? node8050 : node8047;
																assign node8047 = (inp[8]) ? 4'b0011 : 4'b0010;
																assign node8050 = (inp[8]) ? 4'b0010 : 4'b0011;
														assign node8053 = (inp[4]) ? 4'b0111 : 4'b0011;
												assign node8056 = (inp[9]) ? node8070 : node8057;
													assign node8057 = (inp[4]) ? node8063 : node8058;
														assign node8058 = (inp[8]) ? 4'b0110 : node8059;
															assign node8059 = (inp[7]) ? 4'b0111 : 4'b0110;
														assign node8063 = (inp[7]) ? node8067 : node8064;
															assign node8064 = (inp[8]) ? 4'b0011 : 4'b0010;
															assign node8067 = (inp[8]) ? 4'b0010 : 4'b0011;
													assign node8070 = (inp[4]) ? node8078 : node8071;
														assign node8071 = (inp[8]) ? node8075 : node8072;
															assign node8072 = (inp[7]) ? 4'b0011 : 4'b0010;
															assign node8075 = (inp[7]) ? 4'b0010 : 4'b0011;
														assign node8078 = (inp[8]) ? 4'b0111 : node8079;
															assign node8079 = (inp[14]) ? 4'b0111 : 4'b0110;
											assign node8083 = (inp[14]) ? node8127 : node8084;
												assign node8084 = (inp[4]) ? node8106 : node8085;
													assign node8085 = (inp[9]) ? node8099 : node8086;
														assign node8086 = (inp[8]) ? node8092 : node8087;
															assign node8087 = (inp[2]) ? node8089 : 4'b0101;
																assign node8089 = (inp[7]) ? 4'b0101 : 4'b0100;
															assign node8092 = (inp[2]) ? node8096 : node8093;
																assign node8093 = (inp[7]) ? 4'b0101 : 4'b0100;
																assign node8096 = (inp[7]) ? 4'b0100 : 4'b0101;
														assign node8099 = (inp[7]) ? node8103 : node8100;
															assign node8100 = (inp[8]) ? 4'b0001 : 4'b0000;
															assign node8103 = (inp[8]) ? 4'b0000 : 4'b0001;
													assign node8106 = (inp[9]) ? node8120 : node8107;
														assign node8107 = (inp[7]) ? node8113 : node8108;
															assign node8108 = (inp[2]) ? 4'b0001 : node8109;
																assign node8109 = (inp[8]) ? 4'b0000 : 4'b0001;
															assign node8113 = (inp[8]) ? node8117 : node8114;
																assign node8114 = (inp[2]) ? 4'b0001 : 4'b0000;
																assign node8117 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node8120 = (inp[2]) ? node8122 : 4'b0101;
															assign node8122 = (inp[7]) ? 4'b0101 : node8123;
																assign node8123 = (inp[8]) ? 4'b0101 : 4'b0100;
												assign node8127 = (inp[9]) ? node8149 : node8128;
													assign node8128 = (inp[4]) ? node8144 : node8129;
														assign node8129 = (inp[2]) ? node8137 : node8130;
															assign node8130 = (inp[8]) ? node8134 : node8131;
																assign node8131 = (inp[7]) ? 4'b0101 : 4'b0100;
																assign node8134 = (inp[7]) ? 4'b0100 : 4'b0101;
															assign node8137 = (inp[8]) ? node8141 : node8138;
																assign node8138 = (inp[7]) ? 4'b0101 : 4'b0100;
																assign node8141 = (inp[7]) ? 4'b0100 : 4'b0101;
														assign node8144 = (inp[7]) ? 4'b0000 : node8145;
															assign node8145 = (inp[8]) ? 4'b0001 : 4'b0000;
													assign node8149 = (inp[4]) ? node8157 : node8150;
														assign node8150 = (inp[8]) ? node8154 : node8151;
															assign node8151 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node8154 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node8157 = (inp[8]) ? node8159 : 4'b0100;
															assign node8159 = (inp[7]) ? 4'b0100 : 4'b0101;
								assign node8162 = (inp[5]) ? node8438 : node8163;
									assign node8163 = (inp[9]) ? node8315 : node8164;
										assign node8164 = (inp[4]) ? node8232 : node8165;
											assign node8165 = (inp[8]) ? node8199 : node8166;
												assign node8166 = (inp[7]) ? node8180 : node8167;
													assign node8167 = (inp[14]) ? 4'b0110 : node8168;
														assign node8168 = (inp[2]) ? node8174 : node8169;
															assign node8169 = (inp[0]) ? 4'b0111 : node8170;
																assign node8170 = (inp[15]) ? 4'b0101 : 4'b0111;
															assign node8174 = (inp[15]) ? node8176 : 4'b0100;
																assign node8176 = (inp[0]) ? 4'b0110 : 4'b0100;
													assign node8180 = (inp[14]) ? node8194 : node8181;
														assign node8181 = (inp[2]) ? node8189 : node8182;
															assign node8182 = (inp[15]) ? node8186 : node8183;
																assign node8183 = (inp[0]) ? 4'b0100 : 4'b0110;
																assign node8186 = (inp[0]) ? 4'b0110 : 4'b0100;
															assign node8189 = (inp[0]) ? 4'b0111 : node8190;
																assign node8190 = (inp[15]) ? 4'b0101 : 4'b0111;
														assign node8194 = (inp[0]) ? node8196 : 4'b0111;
															assign node8196 = (inp[15]) ? 4'b0111 : 4'b0101;
												assign node8199 = (inp[7]) ? node8215 : node8200;
													assign node8200 = (inp[14]) ? node8208 : node8201;
														assign node8201 = (inp[2]) ? node8203 : 4'b0100;
															assign node8203 = (inp[0]) ? node8205 : 4'b0101;
																assign node8205 = (inp[15]) ? 4'b0111 : 4'b0101;
														assign node8208 = (inp[0]) ? node8212 : node8209;
															assign node8209 = (inp[15]) ? 4'b0101 : 4'b0111;
															assign node8212 = (inp[15]) ? 4'b0111 : 4'b0101;
													assign node8215 = (inp[2]) ? node8225 : node8216;
														assign node8216 = (inp[14]) ? node8222 : node8217;
															assign node8217 = (inp[15]) ? 4'b0101 : node8218;
																assign node8218 = (inp[0]) ? 4'b0101 : 4'b0111;
															assign node8222 = (inp[0]) ? 4'b0100 : 4'b0110;
														assign node8225 = (inp[0]) ? node8229 : node8226;
															assign node8226 = (inp[15]) ? 4'b0100 : 4'b0110;
															assign node8229 = (inp[15]) ? 4'b0110 : 4'b0100;
											assign node8232 = (inp[2]) ? node8278 : node8233;
												assign node8233 = (inp[8]) ? node8261 : node8234;
													assign node8234 = (inp[7]) ? node8250 : node8235;
														assign node8235 = (inp[14]) ? node8243 : node8236;
															assign node8236 = (inp[0]) ? node8240 : node8237;
																assign node8237 = (inp[15]) ? 4'b0001 : 4'b0011;
																assign node8240 = (inp[15]) ? 4'b0011 : 4'b0001;
															assign node8243 = (inp[15]) ? node8247 : node8244;
																assign node8244 = (inp[0]) ? 4'b0000 : 4'b0010;
																assign node8247 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node8250 = (inp[14]) ? node8256 : node8251;
															assign node8251 = (inp[15]) ? 4'b0000 : node8252;
																assign node8252 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node8256 = (inp[15]) ? node8258 : 4'b0001;
																assign node8258 = (inp[0]) ? 4'b0011 : 4'b0001;
													assign node8261 = (inp[7]) ? node8269 : node8262;
														assign node8262 = (inp[14]) ? 4'b0011 : node8263;
															assign node8263 = (inp[15]) ? node8265 : 4'b0000;
																assign node8265 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node8269 = (inp[14]) ? node8273 : node8270;
															assign node8270 = (inp[15]) ? 4'b0011 : 4'b0001;
															assign node8273 = (inp[0]) ? 4'b0000 : node8274;
																assign node8274 = (inp[15]) ? 4'b0000 : 4'b0010;
												assign node8278 = (inp[7]) ? node8294 : node8279;
													assign node8279 = (inp[8]) ? node8285 : node8280;
														assign node8280 = (inp[15]) ? node8282 : 4'b0010;
															assign node8282 = (inp[14]) ? 4'b0000 : 4'b0010;
														assign node8285 = (inp[14]) ? 4'b0011 : node8286;
															assign node8286 = (inp[0]) ? node8290 : node8287;
																assign node8287 = (inp[15]) ? 4'b0001 : 4'b0011;
																assign node8290 = (inp[15]) ? 4'b0011 : 4'b0001;
													assign node8294 = (inp[8]) ? node8306 : node8295;
														assign node8295 = (inp[14]) ? node8301 : node8296;
															assign node8296 = (inp[15]) ? node8298 : 4'b0001;
																assign node8298 = (inp[0]) ? 4'b0011 : 4'b0001;
															assign node8301 = (inp[0]) ? 4'b0001 : node8302;
																assign node8302 = (inp[15]) ? 4'b0001 : 4'b0011;
														assign node8306 = (inp[14]) ? 4'b0010 : node8307;
															assign node8307 = (inp[15]) ? node8311 : node8308;
																assign node8308 = (inp[0]) ? 4'b0000 : 4'b0010;
																assign node8311 = (inp[0]) ? 4'b0010 : 4'b0000;
										assign node8315 = (inp[4]) ? node8375 : node8316;
											assign node8316 = (inp[15]) ? node8348 : node8317;
												assign node8317 = (inp[0]) ? node8329 : node8318;
													assign node8318 = (inp[7]) ? node8324 : node8319;
														assign node8319 = (inp[8]) ? node8321 : 4'b0010;
															assign node8321 = (inp[14]) ? 4'b0011 : 4'b0010;
														assign node8324 = (inp[8]) ? node8326 : 4'b0011;
															assign node8326 = (inp[2]) ? 4'b0010 : 4'b0011;
													assign node8329 = (inp[14]) ? node8343 : node8330;
														assign node8330 = (inp[7]) ? node8336 : node8331;
															assign node8331 = (inp[8]) ? node8333 : 4'b0000;
																assign node8333 = (inp[2]) ? 4'b0001 : 4'b0000;
															assign node8336 = (inp[2]) ? node8340 : node8337;
																assign node8337 = (inp[8]) ? 4'b0001 : 4'b0000;
																assign node8340 = (inp[8]) ? 4'b0000 : 4'b0001;
														assign node8343 = (inp[7]) ? node8345 : 4'b0001;
															assign node8345 = (inp[8]) ? 4'b0000 : 4'b0001;
												assign node8348 = (inp[0]) ? node8370 : node8349;
													assign node8349 = (inp[2]) ? node8363 : node8350;
														assign node8350 = (inp[8]) ? node8358 : node8351;
															assign node8351 = (inp[14]) ? node8355 : node8352;
																assign node8352 = (inp[7]) ? 4'b0000 : 4'b0001;
																assign node8355 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node8358 = (inp[14]) ? node8360 : 4'b0000;
																assign node8360 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node8363 = (inp[8]) ? node8367 : node8364;
															assign node8364 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node8367 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node8370 = (inp[14]) ? 4'b0010 : node8371;
														assign node8371 = (inp[7]) ? 4'b0011 : 4'b0010;
											assign node8375 = (inp[14]) ? node8409 : node8376;
												assign node8376 = (inp[7]) ? node8394 : node8377;
													assign node8377 = (inp[8]) ? node8385 : node8378;
														assign node8378 = (inp[2]) ? 4'b0100 : node8379;
															assign node8379 = (inp[0]) ? 4'b0101 : node8380;
																assign node8380 = (inp[15]) ? 4'b0111 : 4'b0101;
														assign node8385 = (inp[2]) ? 4'b0101 : node8386;
															assign node8386 = (inp[15]) ? node8390 : node8387;
																assign node8387 = (inp[0]) ? 4'b0110 : 4'b0100;
																assign node8390 = (inp[0]) ? 4'b0100 : 4'b0110;
													assign node8394 = (inp[2]) ? node8404 : node8395;
														assign node8395 = (inp[8]) ? 4'b0101 : node8396;
															assign node8396 = (inp[15]) ? node8400 : node8397;
																assign node8397 = (inp[0]) ? 4'b0110 : 4'b0100;
																assign node8400 = (inp[0]) ? 4'b0100 : 4'b0110;
														assign node8404 = (inp[15]) ? 4'b0110 : node8405;
															assign node8405 = (inp[0]) ? 4'b0110 : 4'b0100;
												assign node8409 = (inp[0]) ? node8425 : node8410;
													assign node8410 = (inp[15]) ? node8418 : node8411;
														assign node8411 = (inp[7]) ? node8415 : node8412;
															assign node8412 = (inp[8]) ? 4'b0101 : 4'b0100;
															assign node8415 = (inp[8]) ? 4'b0100 : 4'b0101;
														assign node8418 = (inp[8]) ? node8422 : node8419;
															assign node8419 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node8422 = (inp[7]) ? 4'b0110 : 4'b0111;
													assign node8425 = (inp[15]) ? node8433 : node8426;
														assign node8426 = (inp[8]) ? node8430 : node8427;
															assign node8427 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node8430 = (inp[2]) ? 4'b0111 : 4'b0110;
														assign node8433 = (inp[8]) ? 4'b0100 : node8434;
															assign node8434 = (inp[7]) ? 4'b0101 : 4'b0100;
									assign node8438 = (inp[8]) ? node8580 : node8439;
										assign node8439 = (inp[7]) ? node8505 : node8440;
											assign node8440 = (inp[2]) ? node8478 : node8441;
												assign node8441 = (inp[14]) ? node8457 : node8442;
													assign node8442 = (inp[4]) ? node8448 : node8443;
														assign node8443 = (inp[9]) ? 4'b0011 : node8444;
															assign node8444 = (inp[0]) ? 4'b0111 : 4'b0101;
														assign node8448 = (inp[9]) ? node8450 : 4'b0001;
															assign node8450 = (inp[15]) ? node8454 : node8451;
																assign node8451 = (inp[0]) ? 4'b0111 : 4'b0101;
																assign node8454 = (inp[0]) ? 4'b0101 : 4'b0111;
													assign node8457 = (inp[4]) ? node8465 : node8458;
														assign node8458 = (inp[9]) ? node8460 : 4'b0100;
															assign node8460 = (inp[0]) ? 4'b0000 : node8461;
																assign node8461 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node8465 = (inp[9]) ? node8473 : node8466;
															assign node8466 = (inp[0]) ? node8470 : node8467;
																assign node8467 = (inp[15]) ? 4'b0010 : 4'b0000;
																assign node8470 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node8473 = (inp[15]) ? node8475 : 4'b0100;
																assign node8475 = (inp[0]) ? 4'b0100 : 4'b0110;
												assign node8478 = (inp[9]) ? node8492 : node8479;
													assign node8479 = (inp[4]) ? node8485 : node8480;
														assign node8480 = (inp[0]) ? 4'b0110 : node8481;
															assign node8481 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node8485 = (inp[0]) ? node8489 : node8486;
															assign node8486 = (inp[15]) ? 4'b0010 : 4'b0000;
															assign node8489 = (inp[15]) ? 4'b0000 : 4'b0010;
													assign node8492 = (inp[4]) ? node8498 : node8493;
														assign node8493 = (inp[0]) ? node8495 : 4'b0010;
															assign node8495 = (inp[15]) ? 4'b0000 : 4'b0010;
														assign node8498 = (inp[0]) ? node8502 : node8499;
															assign node8499 = (inp[15]) ? 4'b0110 : 4'b0100;
															assign node8502 = (inp[15]) ? 4'b0100 : 4'b0110;
											assign node8505 = (inp[2]) ? node8547 : node8506;
												assign node8506 = (inp[14]) ? node8532 : node8507;
													assign node8507 = (inp[15]) ? node8521 : node8508;
														assign node8508 = (inp[0]) ? node8514 : node8509;
															assign node8509 = (inp[4]) ? 4'b0000 : node8510;
																assign node8510 = (inp[9]) ? 4'b0000 : 4'b0100;
															assign node8514 = (inp[4]) ? node8518 : node8515;
																assign node8515 = (inp[9]) ? 4'b0010 : 4'b0110;
																assign node8518 = (inp[9]) ? 4'b0110 : 4'b0010;
														assign node8521 = (inp[0]) ? node8527 : node8522;
															assign node8522 = (inp[4]) ? 4'b0110 : node8523;
																assign node8523 = (inp[9]) ? 4'b0010 : 4'b0110;
															assign node8527 = (inp[9]) ? node8529 : 4'b0100;
																assign node8529 = (inp[4]) ? 4'b0100 : 4'b0000;
													assign node8532 = (inp[4]) ? node8540 : node8533;
														assign node8533 = (inp[9]) ? node8535 : 4'b0111;
															assign node8535 = (inp[15]) ? 4'b0011 : node8536;
																assign node8536 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node8540 = (inp[9]) ? node8544 : node8541;
															assign node8541 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node8544 = (inp[15]) ? 4'b0101 : 4'b0111;
												assign node8547 = (inp[0]) ? node8569 : node8548;
													assign node8548 = (inp[15]) ? node8562 : node8549;
														assign node8549 = (inp[14]) ? node8555 : node8550;
															assign node8550 = (inp[4]) ? node8552 : 4'b0001;
																assign node8552 = (inp[9]) ? 4'b0101 : 4'b0001;
															assign node8555 = (inp[4]) ? node8559 : node8556;
																assign node8556 = (inp[9]) ? 4'b0001 : 4'b0101;
																assign node8559 = (inp[9]) ? 4'b0101 : 4'b0001;
														assign node8562 = (inp[4]) ? node8566 : node8563;
															assign node8563 = (inp[9]) ? 4'b0011 : 4'b0111;
															assign node8566 = (inp[9]) ? 4'b0111 : 4'b0011;
													assign node8569 = (inp[15]) ? node8573 : node8570;
														assign node8570 = (inp[4]) ? 4'b0111 : 4'b0011;
														assign node8573 = (inp[9]) ? node8577 : node8574;
															assign node8574 = (inp[4]) ? 4'b0001 : 4'b0101;
															assign node8577 = (inp[4]) ? 4'b0101 : 4'b0001;
										assign node8580 = (inp[7]) ? node8662 : node8581;
											assign node8581 = (inp[14]) ? node8625 : node8582;
												assign node8582 = (inp[2]) ? node8606 : node8583;
													assign node8583 = (inp[15]) ? node8599 : node8584;
														assign node8584 = (inp[0]) ? node8592 : node8585;
															assign node8585 = (inp[4]) ? node8589 : node8586;
																assign node8586 = (inp[9]) ? 4'b0000 : 4'b0100;
																assign node8589 = (inp[9]) ? 4'b0100 : 4'b0000;
															assign node8592 = (inp[9]) ? node8596 : node8593;
																assign node8593 = (inp[4]) ? 4'b0010 : 4'b0110;
																assign node8596 = (inp[4]) ? 4'b0110 : 4'b0010;
														assign node8599 = (inp[0]) ? 4'b0100 : node8600;
															assign node8600 = (inp[9]) ? node8602 : 4'b0110;
																assign node8602 = (inp[4]) ? 4'b0110 : 4'b0010;
													assign node8606 = (inp[9]) ? node8618 : node8607;
														assign node8607 = (inp[4]) ? node8615 : node8608;
															assign node8608 = (inp[0]) ? node8612 : node8609;
																assign node8609 = (inp[15]) ? 4'b0111 : 4'b0101;
																assign node8612 = (inp[15]) ? 4'b0101 : 4'b0111;
															assign node8615 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node8618 = (inp[0]) ? node8622 : node8619;
															assign node8619 = (inp[15]) ? 4'b0111 : 4'b0101;
															assign node8622 = (inp[15]) ? 4'b0101 : 4'b0111;
												assign node8625 = (inp[2]) ? node8643 : node8626;
													assign node8626 = (inp[0]) ? node8636 : node8627;
														assign node8627 = (inp[15]) ? node8631 : node8628;
															assign node8628 = (inp[4]) ? 4'b0001 : 4'b0101;
															assign node8631 = (inp[9]) ? node8633 : 4'b0011;
																assign node8633 = (inp[4]) ? 4'b0111 : 4'b0011;
														assign node8636 = (inp[15]) ? 4'b0101 : node8637;
															assign node8637 = (inp[4]) ? 4'b0111 : node8638;
																assign node8638 = (inp[9]) ? 4'b0011 : 4'b0111;
													assign node8643 = (inp[15]) ? node8655 : node8644;
														assign node8644 = (inp[0]) ? node8650 : node8645;
															assign node8645 = (inp[4]) ? 4'b0101 : node8646;
																assign node8646 = (inp[9]) ? 4'b0001 : 4'b0101;
															assign node8650 = (inp[4]) ? 4'b0111 : node8651;
																assign node8651 = (inp[9]) ? 4'b0011 : 4'b0111;
														assign node8655 = (inp[0]) ? node8657 : 4'b0011;
															assign node8657 = (inp[9]) ? node8659 : 4'b0001;
																assign node8659 = (inp[4]) ? 4'b0101 : 4'b0001;
											assign node8662 = (inp[2]) ? node8694 : node8663;
												assign node8663 = (inp[14]) ? node8681 : node8664;
													assign node8664 = (inp[4]) ? node8674 : node8665;
														assign node8665 = (inp[9]) ? node8671 : node8666;
															assign node8666 = (inp[15]) ? 4'b0111 : node8667;
																assign node8667 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node8671 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node8674 = (inp[9]) ? 4'b0101 : node8675;
															assign node8675 = (inp[0]) ? 4'b0001 : node8676;
																assign node8676 = (inp[15]) ? 4'b0011 : 4'b0001;
													assign node8681 = (inp[9]) ? node8687 : node8682;
														assign node8682 = (inp[15]) ? 4'b0100 : node8683;
															assign node8683 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node8687 = (inp[4]) ? node8689 : 4'b0000;
															assign node8689 = (inp[0]) ? 4'b0100 : node8690;
																assign node8690 = (inp[15]) ? 4'b0110 : 4'b0100;
												assign node8694 = (inp[0]) ? node8708 : node8695;
													assign node8695 = (inp[15]) ? node8701 : node8696;
														assign node8696 = (inp[4]) ? node8698 : 4'b0100;
															assign node8698 = (inp[9]) ? 4'b0100 : 4'b0000;
														assign node8701 = (inp[4]) ? node8705 : node8702;
															assign node8702 = (inp[9]) ? 4'b0010 : 4'b0110;
															assign node8705 = (inp[9]) ? 4'b0110 : 4'b0010;
													assign node8708 = (inp[15]) ? node8718 : node8709;
														assign node8709 = (inp[14]) ? 4'b0010 : node8710;
															assign node8710 = (inp[9]) ? node8714 : node8711;
																assign node8711 = (inp[4]) ? 4'b0010 : 4'b0110;
																assign node8714 = (inp[4]) ? 4'b0110 : 4'b0010;
														assign node8718 = (inp[9]) ? node8722 : node8719;
															assign node8719 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node8722 = (inp[4]) ? 4'b0100 : 4'b0000;
						assign node8725 = (inp[8]) ? node9647 : node8726;
							assign node8726 = (inp[7]) ? node9198 : node8727;
								assign node8727 = (inp[14]) ? node8979 : node8728;
									assign node8728 = (inp[2]) ? node8870 : node8729;
										assign node8729 = (inp[5]) ? node8803 : node8730;
											assign node8730 = (inp[12]) ? node8766 : node8731;
												assign node8731 = (inp[4]) ? node8751 : node8732;
													assign node8732 = (inp[9]) ? node8746 : node8733;
														assign node8733 = (inp[3]) ? node8739 : node8734;
															assign node8734 = (inp[15]) ? node8736 : 4'b0101;
																assign node8736 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node8739 = (inp[15]) ? node8743 : node8740;
																assign node8740 = (inp[0]) ? 4'b0101 : 4'b0111;
																assign node8743 = (inp[0]) ? 4'b0111 : 4'b0101;
														assign node8746 = (inp[0]) ? 4'b0001 : node8747;
															assign node8747 = (inp[15]) ? 4'b0001 : 4'b0011;
													assign node8751 = (inp[9]) ? node8757 : node8752;
														assign node8752 = (inp[15]) ? 4'b0011 : node8753;
															assign node8753 = (inp[0]) ? 4'b0001 : 4'b0011;
														assign node8757 = (inp[15]) ? 4'b0111 : node8758;
															assign node8758 = (inp[0]) ? node8762 : node8759;
																assign node8759 = (inp[3]) ? 4'b0101 : 4'b0111;
																assign node8762 = (inp[3]) ? 4'b0111 : 4'b0101;
												assign node8766 = (inp[15]) ? node8782 : node8767;
													assign node8767 = (inp[0]) ? node8775 : node8768;
														assign node8768 = (inp[3]) ? 4'b0011 : node8769;
															assign node8769 = (inp[4]) ? node8771 : 4'b0011;
																assign node8771 = (inp[9]) ? 4'b0111 : 4'b0011;
														assign node8775 = (inp[9]) ? node8779 : node8776;
															assign node8776 = (inp[4]) ? 4'b0001 : 4'b0101;
															assign node8779 = (inp[4]) ? 4'b0111 : 4'b0001;
													assign node8782 = (inp[0]) ? node8790 : node8783;
														assign node8783 = (inp[3]) ? 4'b0101 : node8784;
															assign node8784 = (inp[4]) ? node8786 : 4'b0001;
																assign node8786 = (inp[9]) ? 4'b0101 : 4'b0001;
														assign node8790 = (inp[3]) ? node8798 : node8791;
															assign node8791 = (inp[9]) ? node8795 : node8792;
																assign node8792 = (inp[4]) ? 4'b0011 : 4'b0111;
																assign node8795 = (inp[4]) ? 4'b0111 : 4'b0011;
															assign node8798 = (inp[4]) ? node8800 : 4'b0011;
																assign node8800 = (inp[9]) ? 4'b0101 : 4'b0011;
											assign node8803 = (inp[9]) ? node8845 : node8804;
												assign node8804 = (inp[4]) ? node8822 : node8805;
													assign node8805 = (inp[12]) ? node8817 : node8806;
														assign node8806 = (inp[15]) ? node8812 : node8807;
															assign node8807 = (inp[0]) ? node8809 : 4'b0101;
																assign node8809 = (inp[3]) ? 4'b0111 : 4'b0101;
															assign node8812 = (inp[0]) ? node8814 : 4'b0111;
																assign node8814 = (inp[3]) ? 4'b0101 : 4'b0111;
														assign node8817 = (inp[15]) ? 4'b0101 : node8818;
															assign node8818 = (inp[3]) ? 4'b0101 : 4'b0111;
													assign node8822 = (inp[15]) ? node8838 : node8823;
														assign node8823 = (inp[12]) ? node8831 : node8824;
															assign node8824 = (inp[3]) ? node8828 : node8825;
																assign node8825 = (inp[0]) ? 4'b0001 : 4'b0011;
																assign node8828 = (inp[0]) ? 4'b0011 : 4'b0001;
															assign node8831 = (inp[3]) ? node8835 : node8832;
																assign node8832 = (inp[0]) ? 4'b0001 : 4'b0011;
																assign node8835 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node8838 = (inp[3]) ? node8842 : node8839;
															assign node8839 = (inp[0]) ? 4'b0011 : 4'b0001;
															assign node8842 = (inp[0]) ? 4'b0001 : 4'b0011;
												assign node8845 = (inp[4]) ? node8861 : node8846;
													assign node8846 = (inp[15]) ? node8854 : node8847;
														assign node8847 = (inp[12]) ? 4'b0001 : node8848;
															assign node8848 = (inp[3]) ? node8850 : 4'b0001;
																assign node8850 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node8854 = (inp[3]) ? node8858 : node8855;
															assign node8855 = (inp[0]) ? 4'b0011 : 4'b0001;
															assign node8858 = (inp[0]) ? 4'b0001 : 4'b0011;
													assign node8861 = (inp[3]) ? 4'b0101 : node8862;
														assign node8862 = (inp[15]) ? node8866 : node8863;
															assign node8863 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node8866 = (inp[0]) ? 4'b0101 : 4'b0111;
										assign node8870 = (inp[9]) ? node8920 : node8871;
											assign node8871 = (inp[4]) ? node8891 : node8872;
												assign node8872 = (inp[15]) ? node8882 : node8873;
													assign node8873 = (inp[12]) ? node8875 : 4'b0110;
														assign node8875 = (inp[5]) ? node8877 : 4'b0100;
															assign node8877 = (inp[3]) ? node8879 : 4'b0110;
																assign node8879 = (inp[0]) ? 4'b0110 : 4'b0100;
													assign node8882 = (inp[12]) ? node8884 : 4'b0100;
														assign node8884 = (inp[5]) ? node8888 : node8885;
															assign node8885 = (inp[0]) ? 4'b0110 : 4'b0100;
															assign node8888 = (inp[0]) ? 4'b0100 : 4'b0110;
												assign node8891 = (inp[3]) ? node8907 : node8892;
													assign node8892 = (inp[12]) ? node8900 : node8893;
														assign node8893 = (inp[0]) ? node8897 : node8894;
															assign node8894 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node8897 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node8900 = (inp[15]) ? node8904 : node8901;
															assign node8901 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node8904 = (inp[0]) ? 4'b0010 : 4'b0000;
													assign node8907 = (inp[15]) ? node8913 : node8908;
														assign node8908 = (inp[0]) ? node8910 : 4'b0010;
															assign node8910 = (inp[5]) ? 4'b0010 : 4'b0000;
														assign node8913 = (inp[12]) ? 4'b0000 : node8914;
															assign node8914 = (inp[0]) ? node8916 : 4'b0010;
																assign node8916 = (inp[5]) ? 4'b0000 : 4'b0010;
											assign node8920 = (inp[4]) ? node8942 : node8921;
												assign node8921 = (inp[3]) ? node8927 : node8922;
													assign node8922 = (inp[15]) ? 4'b0000 : node8923;
														assign node8923 = (inp[0]) ? 4'b0000 : 4'b0010;
													assign node8927 = (inp[15]) ? node8937 : node8928;
														assign node8928 = (inp[12]) ? node8930 : 4'b0000;
															assign node8930 = (inp[5]) ? node8934 : node8931;
																assign node8931 = (inp[0]) ? 4'b0000 : 4'b0010;
																assign node8934 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node8937 = (inp[12]) ? node8939 : 4'b0010;
															assign node8939 = (inp[0]) ? 4'b0000 : 4'b0010;
												assign node8942 = (inp[12]) ? node8960 : node8943;
													assign node8943 = (inp[15]) ? node8953 : node8944;
														assign node8944 = (inp[0]) ? node8948 : node8945;
															assign node8945 = (inp[3]) ? 4'b0100 : 4'b0110;
															assign node8948 = (inp[3]) ? 4'b0110 : node8949;
																assign node8949 = (inp[5]) ? 4'b0110 : 4'b0100;
														assign node8953 = (inp[0]) ? 4'b0100 : node8954;
															assign node8954 = (inp[5]) ? 4'b0110 : node8955;
																assign node8955 = (inp[3]) ? 4'b0110 : 4'b0100;
													assign node8960 = (inp[3]) ? node8974 : node8961;
														assign node8961 = (inp[5]) ? node8967 : node8962;
															assign node8962 = (inp[0]) ? 4'b0100 : node8963;
																assign node8963 = (inp[15]) ? 4'b0100 : 4'b0110;
															assign node8967 = (inp[15]) ? node8971 : node8968;
																assign node8968 = (inp[0]) ? 4'b0110 : 4'b0100;
																assign node8971 = (inp[0]) ? 4'b0100 : 4'b0110;
														assign node8974 = (inp[0]) ? node8976 : 4'b0100;
															assign node8976 = (inp[15]) ? 4'b0100 : 4'b0110;
									assign node8979 = (inp[12]) ? node9115 : node8980;
										assign node8980 = (inp[2]) ? node9052 : node8981;
											assign node8981 = (inp[9]) ? node9015 : node8982;
												assign node8982 = (inp[4]) ? node8998 : node8983;
													assign node8983 = (inp[5]) ? node8989 : node8984;
														assign node8984 = (inp[0]) ? node8986 : 4'b0100;
															assign node8986 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node8989 = (inp[15]) ? 4'b0110 : node8990;
															assign node8990 = (inp[3]) ? node8994 : node8991;
																assign node8991 = (inp[0]) ? 4'b0100 : 4'b0110;
																assign node8994 = (inp[0]) ? 4'b0110 : 4'b0100;
													assign node8998 = (inp[3]) ? node9006 : node8999;
														assign node8999 = (inp[0]) ? node9003 : node9000;
															assign node9000 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node9003 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node9006 = (inp[15]) ? 4'b0000 : node9007;
															assign node9007 = (inp[5]) ? node9011 : node9008;
																assign node9008 = (inp[0]) ? 4'b0000 : 4'b0010;
																assign node9011 = (inp[0]) ? 4'b0010 : 4'b0000;
												assign node9015 = (inp[4]) ? node9035 : node9016;
													assign node9016 = (inp[0]) ? node9026 : node9017;
														assign node9017 = (inp[15]) ? node9023 : node9018;
															assign node9018 = (inp[5]) ? node9020 : 4'b0010;
																assign node9020 = (inp[3]) ? 4'b0000 : 4'b0010;
															assign node9023 = (inp[5]) ? 4'b0010 : 4'b0000;
														assign node9026 = (inp[15]) ? node9032 : node9027;
															assign node9027 = (inp[3]) ? node9029 : 4'b0000;
																assign node9029 = (inp[5]) ? 4'b0010 : 4'b0000;
															assign node9032 = (inp[5]) ? 4'b0000 : 4'b0010;
													assign node9035 = (inp[15]) ? node9047 : node9036;
														assign node9036 = (inp[0]) ? node9042 : node9037;
															assign node9037 = (inp[3]) ? 4'b0100 : node9038;
																assign node9038 = (inp[5]) ? 4'b0100 : 4'b0110;
															assign node9042 = (inp[5]) ? 4'b0110 : node9043;
																assign node9043 = (inp[3]) ? 4'b0110 : 4'b0100;
														assign node9047 = (inp[0]) ? node9049 : 4'b0110;
															assign node9049 = (inp[5]) ? 4'b0100 : 4'b0110;
											assign node9052 = (inp[4]) ? node9090 : node9053;
												assign node9053 = (inp[9]) ? node9075 : node9054;
													assign node9054 = (inp[5]) ? node9066 : node9055;
														assign node9055 = (inp[3]) ? node9061 : node9056;
															assign node9056 = (inp[0]) ? node9058 : 4'b0110;
																assign node9058 = (inp[15]) ? 4'b0110 : 4'b0100;
															assign node9061 = (inp[0]) ? 4'b0100 : node9062;
																assign node9062 = (inp[15]) ? 4'b0100 : 4'b0110;
														assign node9066 = (inp[0]) ? 4'b0110 : node9067;
															assign node9067 = (inp[15]) ? node9071 : node9068;
																assign node9068 = (inp[3]) ? 4'b0100 : 4'b0110;
																assign node9071 = (inp[3]) ? 4'b0110 : 4'b0100;
													assign node9075 = (inp[5]) ? node9081 : node9076;
														assign node9076 = (inp[15]) ? 4'b0010 : node9077;
															assign node9077 = (inp[0]) ? 4'b0000 : 4'b0010;
														assign node9081 = (inp[0]) ? node9083 : 4'b0000;
															assign node9083 = (inp[3]) ? node9087 : node9084;
																assign node9084 = (inp[15]) ? 4'b0010 : 4'b0000;
																assign node9087 = (inp[15]) ? 4'b0000 : 4'b0010;
												assign node9090 = (inp[9]) ? node9104 : node9091;
													assign node9091 = (inp[15]) ? node9101 : node9092;
														assign node9092 = (inp[0]) ? node9096 : node9093;
															assign node9093 = (inp[3]) ? 4'b0000 : 4'b0010;
															assign node9096 = (inp[3]) ? node9098 : 4'b0000;
																assign node9098 = (inp[5]) ? 4'b0010 : 4'b0000;
														assign node9101 = (inp[0]) ? 4'b0010 : 4'b0000;
													assign node9104 = (inp[0]) ? node9106 : 4'b0100;
														assign node9106 = (inp[15]) ? node9110 : node9107;
															assign node9107 = (inp[5]) ? 4'b0110 : 4'b0100;
															assign node9110 = (inp[5]) ? 4'b0100 : node9111;
																assign node9111 = (inp[3]) ? 4'b0100 : 4'b0110;
										assign node9115 = (inp[0]) ? node9149 : node9116;
											assign node9116 = (inp[15]) ? node9136 : node9117;
												assign node9117 = (inp[5]) ? node9123 : node9118;
													assign node9118 = (inp[9]) ? 4'b0010 : node9119;
														assign node9119 = (inp[4]) ? 4'b0010 : 4'b0110;
													assign node9123 = (inp[3]) ? node9131 : node9124;
														assign node9124 = (inp[4]) ? node9128 : node9125;
															assign node9125 = (inp[9]) ? 4'b0010 : 4'b0110;
															assign node9128 = (inp[9]) ? 4'b0100 : 4'b0010;
														assign node9131 = (inp[4]) ? node9133 : 4'b0000;
															assign node9133 = (inp[9]) ? 4'b0100 : 4'b0000;
												assign node9136 = (inp[4]) ? node9144 : node9137;
													assign node9137 = (inp[9]) ? node9139 : 4'b0100;
														assign node9139 = (inp[3]) ? node9141 : 4'b0000;
															assign node9141 = (inp[2]) ? 4'b0000 : 4'b0010;
													assign node9144 = (inp[9]) ? 4'b0110 : node9145;
														assign node9145 = (inp[5]) ? 4'b0010 : 4'b0000;
											assign node9149 = (inp[15]) ? node9175 : node9150;
												assign node9150 = (inp[5]) ? node9166 : node9151;
													assign node9151 = (inp[2]) ? node9159 : node9152;
														assign node9152 = (inp[9]) ? node9156 : node9153;
															assign node9153 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node9156 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node9159 = (inp[9]) ? node9163 : node9160;
															assign node9160 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node9163 = (inp[3]) ? 4'b0110 : 4'b0100;
													assign node9166 = (inp[4]) ? node9172 : node9167;
														assign node9167 = (inp[9]) ? node9169 : 4'b0100;
															assign node9169 = (inp[3]) ? 4'b0010 : 4'b0000;
														assign node9172 = (inp[9]) ? 4'b0110 : 4'b0010;
												assign node9175 = (inp[3]) ? node9185 : node9176;
													assign node9176 = (inp[9]) ? node9180 : node9177;
														assign node9177 = (inp[4]) ? 4'b0010 : 4'b0110;
														assign node9180 = (inp[4]) ? node9182 : 4'b0010;
															assign node9182 = (inp[5]) ? 4'b0100 : 4'b0110;
													assign node9185 = (inp[5]) ? node9191 : node9186;
														assign node9186 = (inp[4]) ? 4'b0100 : node9187;
															assign node9187 = (inp[2]) ? 4'b0010 : 4'b0110;
														assign node9191 = (inp[4]) ? node9195 : node9192;
															assign node9192 = (inp[9]) ? 4'b0000 : 4'b0100;
															assign node9195 = (inp[9]) ? 4'b0100 : 4'b0000;
								assign node9198 = (inp[14]) ? node9430 : node9199;
									assign node9199 = (inp[2]) ? node9295 : node9200;
										assign node9200 = (inp[4]) ? node9252 : node9201;
											assign node9201 = (inp[9]) ? node9231 : node9202;
												assign node9202 = (inp[3]) ? node9222 : node9203;
													assign node9203 = (inp[12]) ? node9209 : node9204;
														assign node9204 = (inp[0]) ? 4'b0110 : node9205;
															assign node9205 = (inp[15]) ? 4'b0100 : 4'b0110;
														assign node9209 = (inp[5]) ? node9217 : node9210;
															assign node9210 = (inp[0]) ? node9214 : node9211;
																assign node9211 = (inp[15]) ? 4'b0100 : 4'b0110;
																assign node9214 = (inp[15]) ? 4'b0110 : 4'b0100;
															assign node9217 = (inp[0]) ? 4'b0110 : node9218;
																assign node9218 = (inp[15]) ? 4'b0100 : 4'b0110;
													assign node9222 = (inp[12]) ? node9224 : 4'b0100;
														assign node9224 = (inp[5]) ? node9226 : 4'b0110;
															assign node9226 = (inp[15]) ? 4'b0110 : node9227;
																assign node9227 = (inp[0]) ? 4'b0110 : 4'b0100;
												assign node9231 = (inp[0]) ? node9243 : node9232;
													assign node9232 = (inp[15]) ? node9238 : node9233;
														assign node9233 = (inp[5]) ? node9235 : 4'b0010;
															assign node9235 = (inp[3]) ? 4'b0000 : 4'b0010;
														assign node9238 = (inp[3]) ? node9240 : 4'b0000;
															assign node9240 = (inp[5]) ? 4'b0010 : 4'b0000;
													assign node9243 = (inp[15]) ? node9247 : node9244;
														assign node9244 = (inp[3]) ? 4'b0010 : 4'b0000;
														assign node9247 = (inp[3]) ? node9249 : 4'b0010;
															assign node9249 = (inp[5]) ? 4'b0000 : 4'b0010;
											assign node9252 = (inp[9]) ? node9272 : node9253;
												assign node9253 = (inp[15]) ? node9265 : node9254;
													assign node9254 = (inp[0]) ? node9260 : node9255;
														assign node9255 = (inp[3]) ? node9257 : 4'b0010;
															assign node9257 = (inp[5]) ? 4'b0000 : 4'b0010;
														assign node9260 = (inp[5]) ? node9262 : 4'b0000;
															assign node9262 = (inp[3]) ? 4'b0010 : 4'b0000;
													assign node9265 = (inp[0]) ? 4'b0010 : node9266;
														assign node9266 = (inp[5]) ? node9268 : 4'b0000;
															assign node9268 = (inp[12]) ? 4'b0000 : 4'b0010;
												assign node9272 = (inp[0]) ? node9284 : node9273;
													assign node9273 = (inp[15]) ? node9279 : node9274;
														assign node9274 = (inp[12]) ? node9276 : 4'b0100;
															assign node9276 = (inp[3]) ? 4'b0100 : 4'b0110;
														assign node9279 = (inp[3]) ? 4'b0110 : node9280;
															assign node9280 = (inp[5]) ? 4'b0110 : 4'b0100;
													assign node9284 = (inp[15]) ? node9290 : node9285;
														assign node9285 = (inp[3]) ? 4'b0110 : node9286;
															assign node9286 = (inp[5]) ? 4'b0110 : 4'b0100;
														assign node9290 = (inp[5]) ? 4'b0100 : node9291;
															assign node9291 = (inp[3]) ? 4'b0100 : 4'b0110;
										assign node9295 = (inp[0]) ? node9359 : node9296;
											assign node9296 = (inp[3]) ? node9326 : node9297;
												assign node9297 = (inp[15]) ? node9311 : node9298;
													assign node9298 = (inp[12]) ? node9304 : node9299;
														assign node9299 = (inp[9]) ? node9301 : 4'b1111;
															assign node9301 = (inp[4]) ? 4'b1111 : 4'b1011;
														assign node9304 = (inp[5]) ? node9306 : 4'b1111;
															assign node9306 = (inp[4]) ? node9308 : 4'b1101;
																assign node9308 = (inp[9]) ? 4'b1001 : 4'b1101;
													assign node9311 = (inp[5]) ? node9321 : node9312;
														assign node9312 = (inp[12]) ? 4'b1001 : node9313;
															assign node9313 = (inp[4]) ? node9317 : node9314;
																assign node9314 = (inp[9]) ? 4'b1001 : 4'b1101;
																assign node9317 = (inp[9]) ? 4'b1101 : 4'b1001;
														assign node9321 = (inp[9]) ? 4'b1111 : node9322;
															assign node9322 = (inp[12]) ? 4'b1001 : 4'b1101;
												assign node9326 = (inp[15]) ? node9346 : node9327;
													assign node9327 = (inp[5]) ? node9333 : node9328;
														assign node9328 = (inp[9]) ? node9330 : 4'b1011;
															assign node9330 = (inp[12]) ? 4'b1001 : 4'b1101;
														assign node9333 = (inp[12]) ? node9341 : node9334;
															assign node9334 = (inp[9]) ? node9338 : node9335;
																assign node9335 = (inp[4]) ? 4'b1001 : 4'b1101;
																assign node9338 = (inp[4]) ? 4'b1101 : 4'b1001;
															assign node9341 = (inp[4]) ? 4'b1101 : node9342;
																assign node9342 = (inp[9]) ? 4'b1101 : 4'b1001;
													assign node9346 = (inp[5]) ? node9354 : node9347;
														assign node9347 = (inp[4]) ? 4'b1111 : node9348;
															assign node9348 = (inp[12]) ? 4'b1001 : node9349;
																assign node9349 = (inp[9]) ? 4'b1001 : 4'b1101;
														assign node9354 = (inp[4]) ? 4'b1011 : node9355;
															assign node9355 = (inp[9]) ? 4'b1011 : 4'b1111;
											assign node9359 = (inp[4]) ? node9401 : node9360;
												assign node9360 = (inp[15]) ? node9380 : node9361;
													assign node9361 = (inp[3]) ? node9371 : node9362;
														assign node9362 = (inp[5]) ? node9368 : node9363;
															assign node9363 = (inp[12]) ? node9365 : 4'b1001;
																assign node9365 = (inp[9]) ? 4'b1101 : 4'b1001;
															assign node9368 = (inp[9]) ? 4'b1111 : 4'b1101;
														assign node9371 = (inp[5]) ? node9375 : node9372;
															assign node9372 = (inp[9]) ? 4'b1111 : 4'b1101;
															assign node9375 = (inp[9]) ? node9377 : 4'b1011;
																assign node9377 = (inp[12]) ? 4'b1111 : 4'b1011;
													assign node9380 = (inp[3]) ? node9392 : node9381;
														assign node9381 = (inp[5]) ? node9387 : node9382;
															assign node9382 = (inp[12]) ? 4'b1111 : node9383;
																assign node9383 = (inp[9]) ? 4'b1011 : 4'b1111;
															assign node9387 = (inp[12]) ? 4'b1011 : node9388;
																assign node9388 = (inp[9]) ? 4'b1011 : 4'b1111;
														assign node9392 = (inp[5]) ? 4'b1001 : node9393;
															assign node9393 = (inp[12]) ? node9397 : node9394;
																assign node9394 = (inp[9]) ? 4'b1011 : 4'b1111;
																assign node9397 = (inp[9]) ? 4'b1101 : 4'b1011;
												assign node9401 = (inp[9]) ? node9417 : node9402;
													assign node9402 = (inp[12]) ? node9414 : node9403;
														assign node9403 = (inp[15]) ? node9409 : node9404;
															assign node9404 = (inp[3]) ? node9406 : 4'b1001;
																assign node9406 = (inp[5]) ? 4'b1011 : 4'b1001;
															assign node9409 = (inp[3]) ? node9411 : 4'b1011;
																assign node9411 = (inp[5]) ? 4'b1001 : 4'b1011;
														assign node9414 = (inp[5]) ? 4'b1111 : 4'b1101;
													assign node9417 = (inp[12]) ? node9423 : node9418;
														assign node9418 = (inp[15]) ? 4'b1101 : node9419;
															assign node9419 = (inp[3]) ? 4'b1111 : 4'b1101;
														assign node9423 = (inp[15]) ? 4'b1001 : node9424;
															assign node9424 = (inp[5]) ? 4'b1011 : node9425;
																assign node9425 = (inp[3]) ? 4'b1011 : 4'b1001;
									assign node9430 = (inp[5]) ? node9546 : node9431;
										assign node9431 = (inp[9]) ? node9487 : node9432;
											assign node9432 = (inp[3]) ? node9464 : node9433;
												assign node9433 = (inp[0]) ? node9447 : node9434;
													assign node9434 = (inp[15]) ? node9440 : node9435;
														assign node9435 = (inp[12]) ? 4'b1011 : node9436;
															assign node9436 = (inp[4]) ? 4'b1011 : 4'b1111;
														assign node9440 = (inp[12]) ? node9444 : node9441;
															assign node9441 = (inp[4]) ? 4'b1001 : 4'b1101;
															assign node9444 = (inp[4]) ? 4'b1101 : 4'b1001;
													assign node9447 = (inp[15]) ? node9457 : node9448;
														assign node9448 = (inp[2]) ? 4'b1101 : node9449;
															assign node9449 = (inp[4]) ? node9453 : node9450;
																assign node9450 = (inp[12]) ? 4'b1001 : 4'b1101;
																assign node9453 = (inp[12]) ? 4'b1101 : 4'b1001;
														assign node9457 = (inp[2]) ? 4'b1111 : node9458;
															assign node9458 = (inp[4]) ? node9460 : 4'b1011;
																assign node9460 = (inp[12]) ? 4'b1111 : 4'b1011;
												assign node9464 = (inp[15]) ? node9476 : node9465;
													assign node9465 = (inp[0]) ? node9471 : node9466;
														assign node9466 = (inp[4]) ? node9468 : 4'b1011;
															assign node9468 = (inp[12]) ? 4'b1101 : 4'b1011;
														assign node9471 = (inp[4]) ? 4'b1001 : node9472;
															assign node9472 = (inp[12]) ? 4'b1001 : 4'b1101;
													assign node9476 = (inp[4]) ? node9480 : node9477;
														assign node9477 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node9480 = (inp[12]) ? node9484 : node9481;
															assign node9481 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node9484 = (inp[0]) ? 4'b1101 : 4'b1111;
											assign node9487 = (inp[4]) ? node9513 : node9488;
												assign node9488 = (inp[12]) ? node9504 : node9489;
													assign node9489 = (inp[3]) ? node9497 : node9490;
														assign node9490 = (inp[15]) ? node9494 : node9491;
															assign node9491 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node9494 = (inp[2]) ? 4'b1001 : 4'b1011;
														assign node9497 = (inp[0]) ? node9501 : node9498;
															assign node9498 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node9501 = (inp[15]) ? 4'b1011 : 4'b1001;
													assign node9504 = (inp[3]) ? node9506 : 4'b1111;
														assign node9506 = (inp[0]) ? node9510 : node9507;
															assign node9507 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node9510 = (inp[15]) ? 4'b1101 : 4'b1111;
												assign node9513 = (inp[12]) ? node9531 : node9514;
													assign node9514 = (inp[0]) ? node9522 : node9515;
														assign node9515 = (inp[3]) ? node9519 : node9516;
															assign node9516 = (inp[15]) ? 4'b1101 : 4'b1111;
															assign node9519 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node9522 = (inp[2]) ? node9528 : node9523;
															assign node9523 = (inp[3]) ? 4'b1111 : node9524;
																assign node9524 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node9528 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node9531 = (inp[15]) ? node9539 : node9532;
														assign node9532 = (inp[0]) ? node9536 : node9533;
															assign node9533 = (inp[3]) ? 4'b1001 : 4'b1011;
															assign node9536 = (inp[3]) ? 4'b1011 : 4'b1001;
														assign node9539 = (inp[0]) ? node9543 : node9540;
															assign node9540 = (inp[3]) ? 4'b1011 : 4'b1001;
															assign node9543 = (inp[3]) ? 4'b1001 : 4'b1011;
										assign node9546 = (inp[0]) ? node9606 : node9547;
											assign node9547 = (inp[15]) ? node9575 : node9548;
												assign node9548 = (inp[3]) ? node9562 : node9549;
													assign node9549 = (inp[12]) ? node9557 : node9550;
														assign node9550 = (inp[9]) ? node9554 : node9551;
															assign node9551 = (inp[4]) ? 4'b1011 : 4'b1111;
															assign node9554 = (inp[4]) ? 4'b1101 : 4'b1011;
														assign node9557 = (inp[4]) ? node9559 : 4'b1101;
															assign node9559 = (inp[9]) ? 4'b1001 : 4'b1101;
													assign node9562 = (inp[12]) ? node9568 : node9563;
														assign node9563 = (inp[9]) ? node9565 : 4'b1101;
															assign node9565 = (inp[4]) ? 4'b1101 : 4'b1001;
														assign node9568 = (inp[9]) ? node9572 : node9569;
															assign node9569 = (inp[4]) ? 4'b1101 : 4'b1001;
															assign node9572 = (inp[4]) ? 4'b1001 : 4'b1101;
												assign node9575 = (inp[3]) ? node9591 : node9576;
													assign node9576 = (inp[12]) ? node9584 : node9577;
														assign node9577 = (inp[9]) ? node9581 : node9578;
															assign node9578 = (inp[4]) ? 4'b1001 : 4'b1101;
															assign node9581 = (inp[4]) ? 4'b1111 : 4'b1001;
														assign node9584 = (inp[2]) ? 4'b1111 : node9585;
															assign node9585 = (inp[9]) ? node9587 : 4'b1001;
																assign node9587 = (inp[4]) ? 4'b1011 : 4'b1111;
													assign node9591 = (inp[9]) ? node9599 : node9592;
														assign node9592 = (inp[12]) ? node9596 : node9593;
															assign node9593 = (inp[4]) ? 4'b1011 : 4'b1111;
															assign node9596 = (inp[4]) ? 4'b1111 : 4'b1011;
														assign node9599 = (inp[12]) ? node9603 : node9600;
															assign node9600 = (inp[4]) ? 4'b1111 : 4'b1011;
															assign node9603 = (inp[4]) ? 4'b1011 : 4'b1111;
											assign node9606 = (inp[15]) ? node9634 : node9607;
												assign node9607 = (inp[3]) ? node9617 : node9608;
													assign node9608 = (inp[4]) ? node9610 : 4'b1001;
														assign node9610 = (inp[12]) ? node9614 : node9611;
															assign node9611 = (inp[9]) ? 4'b1111 : 4'b1001;
															assign node9614 = (inp[9]) ? 4'b1011 : 4'b1111;
													assign node9617 = (inp[4]) ? node9627 : node9618;
														assign node9618 = (inp[2]) ? node9620 : 4'b1011;
															assign node9620 = (inp[9]) ? node9624 : node9621;
																assign node9621 = (inp[12]) ? 4'b1011 : 4'b1111;
																assign node9624 = (inp[12]) ? 4'b1111 : 4'b1011;
														assign node9627 = (inp[9]) ? node9631 : node9628;
															assign node9628 = (inp[12]) ? 4'b1111 : 4'b1011;
															assign node9631 = (inp[12]) ? 4'b1011 : 4'b1111;
												assign node9634 = (inp[3]) ? node9644 : node9635;
													assign node9635 = (inp[12]) ? node9637 : 4'b1011;
														assign node9637 = (inp[4]) ? node9641 : node9638;
															assign node9638 = (inp[9]) ? 4'b1101 : 4'b1011;
															assign node9641 = (inp[9]) ? 4'b1001 : 4'b1101;
													assign node9644 = (inp[4]) ? 4'b1101 : 4'b1001;
							assign node9647 = (inp[7]) ? node10217 : node9648;
								assign node9648 = (inp[2]) ? node9904 : node9649;
									assign node9649 = (inp[14]) ? node9757 : node9650;
										assign node9650 = (inp[15]) ? node9708 : node9651;
											assign node9651 = (inp[0]) ? node9683 : node9652;
												assign node9652 = (inp[3]) ? node9668 : node9653;
													assign node9653 = (inp[12]) ? node9661 : node9654;
														assign node9654 = (inp[9]) ? node9658 : node9655;
															assign node9655 = (inp[4]) ? 4'b0010 : 4'b0110;
															assign node9658 = (inp[4]) ? 4'b0110 : 4'b0010;
														assign node9661 = (inp[9]) ? node9665 : node9662;
															assign node9662 = (inp[4]) ? 4'b0010 : 4'b0110;
															assign node9665 = (inp[4]) ? 4'b0100 : 4'b0010;
													assign node9668 = (inp[5]) ? node9676 : node9669;
														assign node9669 = (inp[4]) ? node9673 : node9670;
															assign node9670 = (inp[9]) ? 4'b0010 : 4'b0110;
															assign node9673 = (inp[9]) ? 4'b0100 : 4'b0010;
														assign node9676 = (inp[12]) ? 4'b0000 : node9677;
															assign node9677 = (inp[9]) ? node9679 : 4'b0100;
																assign node9679 = (inp[4]) ? 4'b0100 : 4'b0000;
												assign node9683 = (inp[3]) ? node9693 : node9684;
													assign node9684 = (inp[4]) ? node9688 : node9685;
														assign node9685 = (inp[9]) ? 4'b0000 : 4'b0100;
														assign node9688 = (inp[9]) ? node9690 : 4'b0000;
															assign node9690 = (inp[5]) ? 4'b0110 : 4'b0100;
													assign node9693 = (inp[5]) ? node9701 : node9694;
														assign node9694 = (inp[4]) ? node9698 : node9695;
															assign node9695 = (inp[9]) ? 4'b0000 : 4'b0100;
															assign node9698 = (inp[9]) ? 4'b0110 : 4'b0000;
														assign node9701 = (inp[9]) ? node9705 : node9702;
															assign node9702 = (inp[4]) ? 4'b0010 : 4'b0110;
															assign node9705 = (inp[4]) ? 4'b0110 : 4'b0010;
											assign node9708 = (inp[0]) ? node9730 : node9709;
												assign node9709 = (inp[5]) ? node9717 : node9710;
													assign node9710 = (inp[4]) ? node9714 : node9711;
														assign node9711 = (inp[9]) ? 4'b0000 : 4'b0100;
														assign node9714 = (inp[9]) ? 4'b0100 : 4'b0000;
													assign node9717 = (inp[3]) ? node9723 : node9718;
														assign node9718 = (inp[9]) ? node9720 : 4'b0000;
															assign node9720 = (inp[4]) ? 4'b0110 : 4'b0000;
														assign node9723 = (inp[12]) ? node9725 : 4'b0010;
															assign node9725 = (inp[4]) ? node9727 : 4'b0110;
																assign node9727 = (inp[9]) ? 4'b0110 : 4'b0010;
												assign node9730 = (inp[3]) ? node9736 : node9731;
													assign node9731 = (inp[4]) ? 4'b0010 : node9732;
														assign node9732 = (inp[9]) ? 4'b0010 : 4'b0110;
													assign node9736 = (inp[5]) ? node9742 : node9737;
														assign node9737 = (inp[12]) ? node9739 : 4'b0010;
															assign node9739 = (inp[4]) ? 4'b0100 : 4'b0010;
														assign node9742 = (inp[12]) ? node9750 : node9743;
															assign node9743 = (inp[9]) ? node9747 : node9744;
																assign node9744 = (inp[4]) ? 4'b0000 : 4'b0100;
																assign node9747 = (inp[4]) ? 4'b0100 : 4'b0000;
															assign node9750 = (inp[9]) ? node9754 : node9751;
																assign node9751 = (inp[4]) ? 4'b0000 : 4'b0100;
																assign node9754 = (inp[4]) ? 4'b0100 : 4'b0000;
										assign node9757 = (inp[5]) ? node9829 : node9758;
											assign node9758 = (inp[15]) ? node9790 : node9759;
												assign node9759 = (inp[0]) ? node9775 : node9760;
													assign node9760 = (inp[4]) ? node9770 : node9761;
														assign node9761 = (inp[3]) ? node9765 : node9762;
															assign node9762 = (inp[12]) ? 4'b1111 : 4'b1011;
															assign node9765 = (inp[12]) ? 4'b1011 : node9766;
																assign node9766 = (inp[9]) ? 4'b1011 : 4'b1111;
														assign node9770 = (inp[3]) ? node9772 : 4'b1011;
															assign node9772 = (inp[9]) ? 4'b1001 : 4'b1101;
													assign node9775 = (inp[3]) ? node9777 : 4'b1001;
														assign node9777 = (inp[4]) ? node9783 : node9778;
															assign node9778 = (inp[9]) ? 4'b1001 : node9779;
																assign node9779 = (inp[12]) ? 4'b1001 : 4'b1101;
															assign node9783 = (inp[9]) ? node9787 : node9784;
																assign node9784 = (inp[12]) ? 4'b1111 : 4'b1001;
																assign node9787 = (inp[12]) ? 4'b1011 : 4'b1111;
												assign node9790 = (inp[0]) ? node9812 : node9791;
													assign node9791 = (inp[3]) ? node9803 : node9792;
														assign node9792 = (inp[9]) ? node9798 : node9793;
															assign node9793 = (inp[4]) ? 4'b1101 : node9794;
																assign node9794 = (inp[12]) ? 4'b1001 : 4'b1101;
															assign node9798 = (inp[12]) ? node9800 : 4'b1001;
																assign node9800 = (inp[4]) ? 4'b1001 : 4'b1101;
														assign node9803 = (inp[12]) ? 4'b1111 : node9804;
															assign node9804 = (inp[4]) ? node9808 : node9805;
																assign node9805 = (inp[9]) ? 4'b1001 : 4'b1101;
																assign node9808 = (inp[9]) ? 4'b1111 : 4'b1001;
													assign node9812 = (inp[3]) ? node9820 : node9813;
														assign node9813 = (inp[4]) ? 4'b1111 : node9814;
															assign node9814 = (inp[9]) ? 4'b1011 : node9815;
																assign node9815 = (inp[12]) ? 4'b1011 : 4'b1111;
														assign node9820 = (inp[12]) ? node9822 : 4'b1011;
															assign node9822 = (inp[9]) ? node9826 : node9823;
																assign node9823 = (inp[4]) ? 4'b1101 : 4'b1011;
																assign node9826 = (inp[4]) ? 4'b1001 : 4'b1101;
											assign node9829 = (inp[3]) ? node9871 : node9830;
												assign node9830 = (inp[15]) ? node9852 : node9831;
													assign node9831 = (inp[9]) ? node9845 : node9832;
														assign node9832 = (inp[0]) ? node9838 : node9833;
															assign node9833 = (inp[4]) ? node9835 : 4'b1011;
																assign node9835 = (inp[12]) ? 4'b1101 : 4'b1011;
															assign node9838 = (inp[4]) ? node9842 : node9839;
																assign node9839 = (inp[12]) ? 4'b1001 : 4'b1101;
																assign node9842 = (inp[12]) ? 4'b1111 : 4'b1001;
														assign node9845 = (inp[0]) ? 4'b1111 : node9846;
															assign node9846 = (inp[12]) ? node9848 : 4'b1101;
																assign node9848 = (inp[4]) ? 4'b1001 : 4'b1101;
													assign node9852 = (inp[9]) ? node9866 : node9853;
														assign node9853 = (inp[0]) ? node9861 : node9854;
															assign node9854 = (inp[4]) ? node9858 : node9855;
																assign node9855 = (inp[12]) ? 4'b1001 : 4'b1101;
																assign node9858 = (inp[12]) ? 4'b1111 : 4'b1001;
															assign node9861 = (inp[12]) ? 4'b1101 : node9862;
																assign node9862 = (inp[4]) ? 4'b1011 : 4'b1111;
														assign node9866 = (inp[12]) ? 4'b1011 : node9867;
															assign node9867 = (inp[4]) ? 4'b1111 : 4'b1011;
												assign node9871 = (inp[12]) ? node9883 : node9872;
													assign node9872 = (inp[4]) ? node9880 : node9873;
														assign node9873 = (inp[9]) ? 4'b1011 : node9874;
															assign node9874 = (inp[15]) ? node9876 : 4'b1111;
																assign node9876 = (inp[0]) ? 4'b1101 : 4'b1111;
														assign node9880 = (inp[9]) ? 4'b1111 : 4'b1011;
													assign node9883 = (inp[0]) ? node9893 : node9884;
														assign node9884 = (inp[15]) ? node9886 : 4'b1101;
															assign node9886 = (inp[9]) ? node9890 : node9887;
																assign node9887 = (inp[4]) ? 4'b1111 : 4'b1011;
																assign node9890 = (inp[4]) ? 4'b1011 : 4'b1111;
														assign node9893 = (inp[15]) ? node9899 : node9894;
															assign node9894 = (inp[4]) ? node9896 : 4'b1011;
																assign node9896 = (inp[9]) ? 4'b1011 : 4'b1111;
															assign node9899 = (inp[9]) ? node9901 : 4'b1101;
																assign node9901 = (inp[4]) ? 4'b1001 : 4'b1101;
									assign node9904 = (inp[14]) ? node10054 : node9905;
										assign node9905 = (inp[4]) ? node9975 : node9906;
											assign node9906 = (inp[12]) ? node9940 : node9907;
												assign node9907 = (inp[9]) ? node9927 : node9908;
													assign node9908 = (inp[15]) ? node9920 : node9909;
														assign node9909 = (inp[0]) ? node9915 : node9910;
															assign node9910 = (inp[5]) ? node9912 : 4'b1111;
																assign node9912 = (inp[3]) ? 4'b1101 : 4'b1111;
															assign node9915 = (inp[3]) ? node9917 : 4'b1101;
																assign node9917 = (inp[5]) ? 4'b1111 : 4'b1101;
														assign node9920 = (inp[3]) ? node9922 : 4'b1101;
															assign node9922 = (inp[5]) ? 4'b1111 : node9923;
																assign node9923 = (inp[0]) ? 4'b1111 : 4'b1101;
													assign node9927 = (inp[0]) ? node9933 : node9928;
														assign node9928 = (inp[15]) ? node9930 : 4'b1011;
															assign node9930 = (inp[5]) ? 4'b1011 : 4'b1001;
														assign node9933 = (inp[15]) ? node9935 : 4'b1001;
															assign node9935 = (inp[5]) ? node9937 : 4'b1011;
																assign node9937 = (inp[3]) ? 4'b1001 : 4'b1011;
												assign node9940 = (inp[9]) ? node9960 : node9941;
													assign node9941 = (inp[3]) ? node9949 : node9942;
														assign node9942 = (inp[5]) ? node9944 : 4'b1011;
															assign node9944 = (inp[0]) ? 4'b1011 : node9945;
																assign node9945 = (inp[15]) ? 4'b1001 : 4'b1011;
														assign node9949 = (inp[0]) ? node9955 : node9950;
															assign node9950 = (inp[15]) ? 4'b1011 : node9951;
																assign node9951 = (inp[5]) ? 4'b1001 : 4'b1011;
															assign node9955 = (inp[5]) ? node9957 : 4'b1001;
																assign node9957 = (inp[15]) ? 4'b1001 : 4'b1011;
													assign node9960 = (inp[0]) ? node9970 : node9961;
														assign node9961 = (inp[15]) ? node9965 : node9962;
															assign node9962 = (inp[3]) ? 4'b1101 : 4'b1111;
															assign node9965 = (inp[5]) ? 4'b1111 : node9966;
																assign node9966 = (inp[3]) ? 4'b1111 : 4'b1101;
														assign node9970 = (inp[15]) ? node9972 : 4'b1111;
															assign node9972 = (inp[3]) ? 4'b1101 : 4'b1111;
											assign node9975 = (inp[15]) ? node10019 : node9976;
												assign node9976 = (inp[3]) ? node10004 : node9977;
													assign node9977 = (inp[0]) ? node9989 : node9978;
														assign node9978 = (inp[5]) ? node9986 : node9979;
															assign node9979 = (inp[9]) ? node9983 : node9980;
																assign node9980 = (inp[12]) ? 4'b1111 : 4'b1011;
																assign node9983 = (inp[12]) ? 4'b1011 : 4'b1111;
															assign node9986 = (inp[9]) ? 4'b1001 : 4'b1101;
														assign node9989 = (inp[5]) ? node9997 : node9990;
															assign node9990 = (inp[12]) ? node9994 : node9991;
																assign node9991 = (inp[9]) ? 4'b1101 : 4'b1001;
																assign node9994 = (inp[9]) ? 4'b1001 : 4'b1101;
															assign node9997 = (inp[12]) ? node10001 : node9998;
																assign node9998 = (inp[9]) ? 4'b1111 : 4'b1001;
																assign node10001 = (inp[9]) ? 4'b1011 : 4'b1111;
													assign node10004 = (inp[0]) ? node10014 : node10005;
														assign node10005 = (inp[12]) ? node10011 : node10006;
															assign node10006 = (inp[9]) ? 4'b1101 : node10007;
																assign node10007 = (inp[5]) ? 4'b1001 : 4'b1011;
															assign node10011 = (inp[9]) ? 4'b1001 : 4'b1101;
														assign node10014 = (inp[9]) ? 4'b1011 : node10015;
															assign node10015 = (inp[12]) ? 4'b1111 : 4'b1011;
												assign node10019 = (inp[0]) ? node10039 : node10020;
													assign node10020 = (inp[3]) ? node10034 : node10021;
														assign node10021 = (inp[5]) ? node10029 : node10022;
															assign node10022 = (inp[9]) ? node10026 : node10023;
																assign node10023 = (inp[12]) ? 4'b1101 : 4'b1001;
																assign node10026 = (inp[12]) ? 4'b1001 : 4'b1101;
															assign node10029 = (inp[9]) ? 4'b1111 : node10030;
																assign node10030 = (inp[12]) ? 4'b1111 : 4'b1001;
														assign node10034 = (inp[12]) ? node10036 : 4'b1111;
															assign node10036 = (inp[5]) ? 4'b1111 : 4'b1011;
													assign node10039 = (inp[3]) ? node10047 : node10040;
														assign node10040 = (inp[5]) ? 4'b1001 : node10041;
															assign node10041 = (inp[9]) ? 4'b1111 : node10042;
																assign node10042 = (inp[12]) ? 4'b1111 : 4'b1011;
														assign node10047 = (inp[9]) ? node10051 : node10048;
															assign node10048 = (inp[12]) ? 4'b1101 : 4'b1001;
															assign node10051 = (inp[12]) ? 4'b1001 : 4'b1101;
										assign node10054 = (inp[3]) ? node10138 : node10055;
											assign node10055 = (inp[12]) ? node10093 : node10056;
												assign node10056 = (inp[15]) ? node10076 : node10057;
													assign node10057 = (inp[0]) ? node10071 : node10058;
														assign node10058 = (inp[5]) ? node10066 : node10059;
															assign node10059 = (inp[4]) ? node10063 : node10060;
																assign node10060 = (inp[9]) ? 4'b1011 : 4'b1111;
																assign node10063 = (inp[9]) ? 4'b1111 : 4'b1011;
															assign node10066 = (inp[4]) ? node10068 : 4'b1011;
																assign node10068 = (inp[9]) ? 4'b1101 : 4'b1011;
														assign node10071 = (inp[5]) ? node10073 : 4'b1001;
															assign node10073 = (inp[9]) ? 4'b1111 : 4'b1001;
													assign node10076 = (inp[0]) ? node10086 : node10077;
														assign node10077 = (inp[5]) ? 4'b1001 : node10078;
															assign node10078 = (inp[4]) ? node10082 : node10079;
																assign node10079 = (inp[9]) ? 4'b1001 : 4'b1101;
																assign node10082 = (inp[9]) ? 4'b1101 : 4'b1001;
														assign node10086 = (inp[5]) ? node10088 : 4'b1011;
															assign node10088 = (inp[9]) ? 4'b1101 : node10089;
																assign node10089 = (inp[4]) ? 4'b1011 : 4'b1111;
												assign node10093 = (inp[5]) ? node10113 : node10094;
													assign node10094 = (inp[15]) ? node10106 : node10095;
														assign node10095 = (inp[0]) ? node10099 : node10096;
															assign node10096 = (inp[4]) ? 4'b1111 : 4'b1011;
															assign node10099 = (inp[9]) ? node10103 : node10100;
																assign node10100 = (inp[4]) ? 4'b1101 : 4'b1001;
																assign node10103 = (inp[4]) ? 4'b1001 : 4'b1101;
														assign node10106 = (inp[0]) ? node10108 : 4'b1101;
															assign node10108 = (inp[4]) ? node10110 : 4'b1111;
																assign node10110 = (inp[9]) ? 4'b1011 : 4'b1111;
													assign node10113 = (inp[4]) ? node10127 : node10114;
														assign node10114 = (inp[9]) ? node10122 : node10115;
															assign node10115 = (inp[0]) ? node10119 : node10116;
																assign node10116 = (inp[15]) ? 4'b1001 : 4'b1011;
																assign node10119 = (inp[15]) ? 4'b1011 : 4'b1001;
															assign node10122 = (inp[15]) ? 4'b1101 : node10123;
																assign node10123 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node10127 = (inp[9]) ? node10133 : node10128;
															assign node10128 = (inp[15]) ? node10130 : 4'b1101;
																assign node10130 = (inp[0]) ? 4'b1101 : 4'b1111;
															assign node10133 = (inp[0]) ? node10135 : 4'b1011;
																assign node10135 = (inp[15]) ? 4'b1001 : 4'b1011;
											assign node10138 = (inp[0]) ? node10182 : node10139;
												assign node10139 = (inp[15]) ? node10165 : node10140;
													assign node10140 = (inp[5]) ? node10152 : node10141;
														assign node10141 = (inp[9]) ? node10147 : node10142;
															assign node10142 = (inp[4]) ? 4'b1101 : node10143;
																assign node10143 = (inp[12]) ? 4'b1011 : 4'b1111;
															assign node10147 = (inp[4]) ? node10149 : 4'b1101;
																assign node10149 = (inp[12]) ? 4'b1001 : 4'b1101;
														assign node10152 = (inp[4]) ? node10158 : node10153;
															assign node10153 = (inp[9]) ? 4'b1001 : node10154;
																assign node10154 = (inp[12]) ? 4'b1001 : 4'b1101;
															assign node10158 = (inp[12]) ? node10162 : node10159;
																assign node10159 = (inp[9]) ? 4'b1101 : 4'b1001;
																assign node10162 = (inp[9]) ? 4'b1001 : 4'b1101;
													assign node10165 = (inp[5]) ? node10175 : node10166;
														assign node10166 = (inp[9]) ? node10172 : node10167;
															assign node10167 = (inp[12]) ? 4'b1001 : node10168;
																assign node10168 = (inp[4]) ? 4'b1001 : 4'b1101;
															assign node10172 = (inp[4]) ? 4'b1111 : 4'b1001;
														assign node10175 = (inp[9]) ? 4'b1011 : node10176;
															assign node10176 = (inp[4]) ? 4'b1111 : node10177;
																assign node10177 = (inp[12]) ? 4'b1011 : 4'b1111;
												assign node10182 = (inp[15]) ? node10200 : node10183;
													assign node10183 = (inp[5]) ? node10191 : node10184;
														assign node10184 = (inp[9]) ? node10186 : 4'b1001;
															assign node10186 = (inp[4]) ? node10188 : 4'b1001;
																assign node10188 = (inp[12]) ? 4'b1011 : 4'b1111;
														assign node10191 = (inp[9]) ? 4'b1111 : node10192;
															assign node10192 = (inp[12]) ? node10196 : node10193;
																assign node10193 = (inp[4]) ? 4'b1011 : 4'b1111;
																assign node10196 = (inp[4]) ? 4'b1111 : 4'b1011;
													assign node10200 = (inp[12]) ? node10212 : node10201;
														assign node10201 = (inp[5]) ? node10207 : node10202;
															assign node10202 = (inp[4]) ? node10204 : 4'b1011;
																assign node10204 = (inp[9]) ? 4'b1101 : 4'b1011;
															assign node10207 = (inp[9]) ? node10209 : 4'b1101;
																assign node10209 = (inp[4]) ? 4'b1101 : 4'b1001;
														assign node10212 = (inp[5]) ? node10214 : 4'b1101;
															assign node10214 = (inp[9]) ? 4'b1101 : 4'b1001;
								assign node10217 = (inp[14]) ? node10485 : node10218;
									assign node10218 = (inp[2]) ? node10358 : node10219;
										assign node10219 = (inp[9]) ? node10293 : node10220;
											assign node10220 = (inp[12]) ? node10258 : node10221;
												assign node10221 = (inp[4]) ? node10239 : node10222;
													assign node10222 = (inp[3]) ? node10230 : node10223;
														assign node10223 = (inp[15]) ? node10227 : node10224;
															assign node10224 = (inp[0]) ? 4'b1101 : 4'b1111;
															assign node10227 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node10230 = (inp[5]) ? node10232 : 4'b1101;
															assign node10232 = (inp[15]) ? node10236 : node10233;
																assign node10233 = (inp[0]) ? 4'b1111 : 4'b1101;
																assign node10236 = (inp[0]) ? 4'b1101 : 4'b1111;
													assign node10239 = (inp[3]) ? node10247 : node10240;
														assign node10240 = (inp[15]) ? node10244 : node10241;
															assign node10241 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node10244 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node10247 = (inp[0]) ? node10253 : node10248;
															assign node10248 = (inp[5]) ? 4'b1011 : node10249;
																assign node10249 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node10253 = (inp[15]) ? node10255 : 4'b1001;
																assign node10255 = (inp[5]) ? 4'b1001 : 4'b1011;
												assign node10258 = (inp[4]) ? node10280 : node10259;
													assign node10259 = (inp[5]) ? node10267 : node10260;
														assign node10260 = (inp[0]) ? node10264 : node10261;
															assign node10261 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node10264 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node10267 = (inp[0]) ? node10275 : node10268;
															assign node10268 = (inp[3]) ? node10272 : node10269;
																assign node10269 = (inp[15]) ? 4'b1001 : 4'b1011;
																assign node10272 = (inp[15]) ? 4'b1011 : 4'b1001;
															assign node10275 = (inp[15]) ? node10277 : 4'b1001;
																assign node10277 = (inp[3]) ? 4'b1001 : 4'b1011;
													assign node10280 = (inp[5]) ? node10286 : node10281;
														assign node10281 = (inp[0]) ? 4'b1101 : node10282;
															assign node10282 = (inp[15]) ? 4'b1101 : 4'b1111;
														assign node10286 = (inp[0]) ? node10290 : node10287;
															assign node10287 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node10290 = (inp[15]) ? 4'b1101 : 4'b1111;
											assign node10293 = (inp[12]) ? node10327 : node10294;
												assign node10294 = (inp[4]) ? node10312 : node10295;
													assign node10295 = (inp[3]) ? node10301 : node10296;
														assign node10296 = (inp[0]) ? 4'b1011 : node10297;
															assign node10297 = (inp[15]) ? 4'b1001 : 4'b1011;
														assign node10301 = (inp[0]) ? node10307 : node10302;
															assign node10302 = (inp[15]) ? 4'b1011 : node10303;
																assign node10303 = (inp[5]) ? 4'b1001 : 4'b1011;
															assign node10307 = (inp[5]) ? 4'b1001 : node10308;
																assign node10308 = (inp[15]) ? 4'b1011 : 4'b1001;
													assign node10312 = (inp[15]) ? node10318 : node10313;
														assign node10313 = (inp[0]) ? node10315 : 4'b1101;
															assign node10315 = (inp[3]) ? 4'b1111 : 4'b1101;
														assign node10318 = (inp[0]) ? node10324 : node10319;
															assign node10319 = (inp[3]) ? 4'b1111 : node10320;
																assign node10320 = (inp[5]) ? 4'b1111 : 4'b1101;
															assign node10324 = (inp[5]) ? 4'b1101 : 4'b1111;
												assign node10327 = (inp[4]) ? node10347 : node10328;
													assign node10328 = (inp[5]) ? node10342 : node10329;
														assign node10329 = (inp[3]) ? node10335 : node10330;
															assign node10330 = (inp[0]) ? node10332 : 4'b1101;
																assign node10332 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node10335 = (inp[0]) ? node10339 : node10336;
																assign node10336 = (inp[15]) ? 4'b1111 : 4'b1101;
																assign node10339 = (inp[15]) ? 4'b1101 : 4'b1111;
														assign node10342 = (inp[0]) ? 4'b1101 : node10343;
															assign node10343 = (inp[3]) ? 4'b1101 : 4'b1111;
													assign node10347 = (inp[15]) ? node10351 : node10348;
														assign node10348 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node10351 = (inp[3]) ? 4'b1001 : node10352;
															assign node10352 = (inp[5]) ? node10354 : 4'b1011;
																assign node10354 = (inp[0]) ? 4'b1001 : 4'b1011;
										assign node10358 = (inp[15]) ? node10424 : node10359;
											assign node10359 = (inp[9]) ? node10391 : node10360;
												assign node10360 = (inp[3]) ? node10376 : node10361;
													assign node10361 = (inp[0]) ? node10371 : node10362;
														assign node10362 = (inp[12]) ? node10366 : node10363;
															assign node10363 = (inp[4]) ? 4'b1010 : 4'b1110;
															assign node10366 = (inp[4]) ? node10368 : 4'b1010;
																assign node10368 = (inp[5]) ? 4'b1100 : 4'b1110;
														assign node10371 = (inp[12]) ? 4'b1110 : node10372;
															assign node10372 = (inp[4]) ? 4'b1000 : 4'b1100;
													assign node10376 = (inp[4]) ? node10384 : node10377;
														assign node10377 = (inp[12]) ? node10379 : 4'b1110;
															assign node10379 = (inp[5]) ? node10381 : 4'b1010;
																assign node10381 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node10384 = (inp[12]) ? node10388 : node10385;
															assign node10385 = (inp[5]) ? 4'b1010 : 4'b1000;
															assign node10388 = (inp[5]) ? 4'b1100 : 4'b1110;
												assign node10391 = (inp[0]) ? node10405 : node10392;
													assign node10392 = (inp[5]) ? node10400 : node10393;
														assign node10393 = (inp[12]) ? 4'b1100 : node10394;
															assign node10394 = (inp[4]) ? node10396 : 4'b1010;
																assign node10396 = (inp[3]) ? 4'b1100 : 4'b1110;
														assign node10400 = (inp[12]) ? node10402 : 4'b1000;
															assign node10402 = (inp[4]) ? 4'b1000 : 4'b1100;
													assign node10405 = (inp[5]) ? node10419 : node10406;
														assign node10406 = (inp[3]) ? node10414 : node10407;
															assign node10407 = (inp[12]) ? node10411 : node10408;
																assign node10408 = (inp[4]) ? 4'b1100 : 4'b1000;
																assign node10411 = (inp[4]) ? 4'b1000 : 4'b1100;
															assign node10414 = (inp[4]) ? 4'b1110 : node10415;
																assign node10415 = (inp[12]) ? 4'b1110 : 4'b1000;
														assign node10419 = (inp[4]) ? node10421 : 4'b1110;
															assign node10421 = (inp[12]) ? 4'b1010 : 4'b1110;
											assign node10424 = (inp[0]) ? node10460 : node10425;
												assign node10425 = (inp[5]) ? node10447 : node10426;
													assign node10426 = (inp[12]) ? node10440 : node10427;
														assign node10427 = (inp[3]) ? node10435 : node10428;
															assign node10428 = (inp[9]) ? node10432 : node10429;
																assign node10429 = (inp[4]) ? 4'b1000 : 4'b1100;
																assign node10432 = (inp[4]) ? 4'b1100 : 4'b1000;
															assign node10435 = (inp[4]) ? 4'b1000 : node10436;
																assign node10436 = (inp[9]) ? 4'b1000 : 4'b1100;
														assign node10440 = (inp[4]) ? node10444 : node10441;
															assign node10441 = (inp[9]) ? 4'b1100 : 4'b1000;
															assign node10444 = (inp[9]) ? 4'b1010 : 4'b1110;
													assign node10447 = (inp[12]) ? node10453 : node10448;
														assign node10448 = (inp[4]) ? node10450 : 4'b1000;
															assign node10450 = (inp[9]) ? 4'b1110 : 4'b1000;
														assign node10453 = (inp[9]) ? node10457 : node10454;
															assign node10454 = (inp[4]) ? 4'b1110 : 4'b1010;
															assign node10457 = (inp[4]) ? 4'b1010 : 4'b1110;
												assign node10460 = (inp[3]) ? node10478 : node10461;
													assign node10461 = (inp[5]) ? node10469 : node10462;
														assign node10462 = (inp[9]) ? node10464 : 4'b1010;
															assign node10464 = (inp[4]) ? node10466 : 4'b1010;
																assign node10466 = (inp[12]) ? 4'b1010 : 4'b1110;
														assign node10469 = (inp[9]) ? node10475 : node10470;
															assign node10470 = (inp[4]) ? 4'b1010 : node10471;
																assign node10471 = (inp[12]) ? 4'b1010 : 4'b1110;
															assign node10475 = (inp[12]) ? 4'b1100 : 4'b1010;
													assign node10478 = (inp[5]) ? node10482 : node10479;
														assign node10479 = (inp[9]) ? 4'b1000 : 4'b1010;
														assign node10482 = (inp[9]) ? 4'b1000 : 4'b1100;
									assign node10485 = (inp[9]) ? node10587 : node10486;
										assign node10486 = (inp[3]) ? node10536 : node10487;
											assign node10487 = (inp[0]) ? node10515 : node10488;
												assign node10488 = (inp[15]) ? node10506 : node10489;
													assign node10489 = (inp[5]) ? node10499 : node10490;
														assign node10490 = (inp[2]) ? node10492 : 4'b1010;
															assign node10492 = (inp[4]) ? node10496 : node10493;
																assign node10493 = (inp[12]) ? 4'b1010 : 4'b1110;
																assign node10496 = (inp[12]) ? 4'b1110 : 4'b1010;
														assign node10499 = (inp[4]) ? node10503 : node10500;
															assign node10500 = (inp[2]) ? 4'b1110 : 4'b1010;
															assign node10503 = (inp[12]) ? 4'b1100 : 4'b1010;
													assign node10506 = (inp[12]) ? node10510 : node10507;
														assign node10507 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node10510 = (inp[4]) ? node10512 : 4'b1000;
															assign node10512 = (inp[5]) ? 4'b1110 : 4'b1100;
												assign node10515 = (inp[15]) ? node10525 : node10516;
													assign node10516 = (inp[12]) ? node10520 : node10517;
														assign node10517 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node10520 = (inp[4]) ? node10522 : 4'b1000;
															assign node10522 = (inp[5]) ? 4'b1110 : 4'b1100;
													assign node10525 = (inp[2]) ? node10527 : 4'b1110;
														assign node10527 = (inp[4]) ? node10531 : node10528;
															assign node10528 = (inp[12]) ? 4'b1010 : 4'b1110;
															assign node10531 = (inp[5]) ? 4'b1100 : node10532;
																assign node10532 = (inp[12]) ? 4'b1110 : 4'b1010;
											assign node10536 = (inp[5]) ? node10564 : node10537;
												assign node10537 = (inp[15]) ? node10551 : node10538;
													assign node10538 = (inp[0]) ? node10544 : node10539;
														assign node10539 = (inp[2]) ? 4'b1010 : node10540;
															assign node10540 = (inp[12]) ? 4'b1100 : 4'b1010;
														assign node10544 = (inp[2]) ? node10548 : node10545;
															assign node10545 = (inp[4]) ? 4'b1110 : 4'b1000;
															assign node10548 = (inp[4]) ? 4'b1000 : 4'b1100;
													assign node10551 = (inp[0]) ? node10559 : node10552;
														assign node10552 = (inp[4]) ? node10556 : node10553;
															assign node10553 = (inp[12]) ? 4'b1000 : 4'b1100;
															assign node10556 = (inp[12]) ? 4'b1110 : 4'b1000;
														assign node10559 = (inp[4]) ? 4'b1100 : node10560;
															assign node10560 = (inp[12]) ? 4'b1010 : 4'b1110;
												assign node10564 = (inp[4]) ? node10580 : node10565;
													assign node10565 = (inp[12]) ? node10573 : node10566;
														assign node10566 = (inp[15]) ? node10570 : node10567;
															assign node10567 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node10570 = (inp[0]) ? 4'b1100 : 4'b1110;
														assign node10573 = (inp[2]) ? node10575 : 4'b1000;
															assign node10575 = (inp[15]) ? node10577 : 4'b1010;
																assign node10577 = (inp[0]) ? 4'b1000 : 4'b1010;
													assign node10580 = (inp[12]) ? 4'b1110 : node10581;
														assign node10581 = (inp[2]) ? 4'b1010 : node10582;
															assign node10582 = (inp[15]) ? 4'b1000 : 4'b1010;
										assign node10587 = (inp[15]) ? node10647 : node10588;
											assign node10588 = (inp[0]) ? node10616 : node10589;
												assign node10589 = (inp[3]) ? node10607 : node10590;
													assign node10590 = (inp[5]) ? node10598 : node10591;
														assign node10591 = (inp[12]) ? node10595 : node10592;
															assign node10592 = (inp[4]) ? 4'b1110 : 4'b1010;
															assign node10595 = (inp[4]) ? 4'b1010 : 4'b1110;
														assign node10598 = (inp[2]) ? node10600 : 4'b1010;
															assign node10600 = (inp[12]) ? node10604 : node10601;
																assign node10601 = (inp[4]) ? 4'b1100 : 4'b1010;
																assign node10604 = (inp[4]) ? 4'b1000 : 4'b1100;
													assign node10607 = (inp[4]) ? node10613 : node10608;
														assign node10608 = (inp[12]) ? 4'b1100 : node10609;
															assign node10609 = (inp[5]) ? 4'b1000 : 4'b1010;
														assign node10613 = (inp[12]) ? 4'b1000 : 4'b1100;
												assign node10616 = (inp[3]) ? node10632 : node10617;
													assign node10617 = (inp[5]) ? node10625 : node10618;
														assign node10618 = (inp[12]) ? node10622 : node10619;
															assign node10619 = (inp[4]) ? 4'b1100 : 4'b1000;
															assign node10622 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node10625 = (inp[4]) ? node10629 : node10626;
															assign node10626 = (inp[12]) ? 4'b1110 : 4'b1000;
															assign node10629 = (inp[12]) ? 4'b1010 : 4'b1110;
													assign node10632 = (inp[2]) ? node10640 : node10633;
														assign node10633 = (inp[12]) ? node10637 : node10634;
															assign node10634 = (inp[5]) ? 4'b1010 : 4'b1000;
															assign node10637 = (inp[4]) ? 4'b1010 : 4'b1110;
														assign node10640 = (inp[12]) ? node10644 : node10641;
															assign node10641 = (inp[4]) ? 4'b1110 : 4'b1010;
															assign node10644 = (inp[4]) ? 4'b1010 : 4'b1110;
											assign node10647 = (inp[0]) ? node10681 : node10648;
												assign node10648 = (inp[5]) ? node10666 : node10649;
													assign node10649 = (inp[3]) ? node10657 : node10650;
														assign node10650 = (inp[2]) ? node10652 : 4'b1100;
															assign node10652 = (inp[12]) ? 4'b1000 : node10653;
																assign node10653 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node10657 = (inp[2]) ? node10659 : 4'b1110;
															assign node10659 = (inp[4]) ? node10663 : node10660;
																assign node10660 = (inp[12]) ? 4'b1110 : 4'b1000;
																assign node10663 = (inp[12]) ? 4'b1010 : 4'b1110;
													assign node10666 = (inp[3]) ? node10672 : node10667;
														assign node10667 = (inp[4]) ? node10669 : 4'b1110;
															assign node10669 = (inp[12]) ? 4'b1010 : 4'b1110;
														assign node10672 = (inp[2]) ? node10676 : node10673;
															assign node10673 = (inp[4]) ? 4'b1110 : 4'b1010;
															assign node10676 = (inp[4]) ? 4'b1010 : node10677;
																assign node10677 = (inp[12]) ? 4'b1110 : 4'b1010;
												assign node10681 = (inp[5]) ? node10697 : node10682;
													assign node10682 = (inp[3]) ? node10690 : node10683;
														assign node10683 = (inp[2]) ? 4'b1010 : node10684;
															assign node10684 = (inp[12]) ? 4'b1110 : node10685;
																assign node10685 = (inp[4]) ? 4'b1110 : 4'b1010;
														assign node10690 = (inp[4]) ? node10694 : node10691;
															assign node10691 = (inp[12]) ? 4'b1100 : 4'b1010;
															assign node10694 = (inp[12]) ? 4'b1000 : 4'b1100;
													assign node10697 = (inp[3]) ? node10705 : node10698;
														assign node10698 = (inp[4]) ? node10702 : node10699;
															assign node10699 = (inp[12]) ? 4'b1100 : 4'b1010;
															assign node10702 = (inp[12]) ? 4'b1000 : 4'b1100;
														assign node10705 = (inp[2]) ? 4'b1100 : node10706;
															assign node10706 = (inp[4]) ? node10710 : node10707;
																assign node10707 = (inp[12]) ? 4'b1100 : 4'b1000;
																assign node10710 = (inp[12]) ? 4'b1000 : 4'b1100;
					assign node10714 = (inp[1]) ? node12710 : node10715;
						assign node10715 = (inp[8]) ? node11705 : node10716;
							assign node10716 = (inp[7]) ? node11136 : node10717;
								assign node10717 = (inp[2]) ? node10957 : node10718;
									assign node10718 = (inp[14]) ? node10834 : node10719;
										assign node10719 = (inp[5]) ? node10769 : node10720;
											assign node10720 = (inp[15]) ? node10740 : node10721;
												assign node10721 = (inp[0]) ? node10731 : node10722;
													assign node10722 = (inp[4]) ? node10726 : node10723;
														assign node10723 = (inp[9]) ? 4'b0011 : 4'b0111;
														assign node10726 = (inp[9]) ? node10728 : 4'b0011;
															assign node10728 = (inp[3]) ? 4'b0101 : 4'b0111;
													assign node10731 = (inp[4]) ? node10735 : node10732;
														assign node10732 = (inp[9]) ? 4'b0001 : 4'b0101;
														assign node10735 = (inp[9]) ? node10737 : 4'b0001;
															assign node10737 = (inp[3]) ? 4'b0111 : 4'b0101;
												assign node10740 = (inp[0]) ? node10756 : node10741;
													assign node10741 = (inp[12]) ? node10749 : node10742;
														assign node10742 = (inp[4]) ? node10746 : node10743;
															assign node10743 = (inp[9]) ? 4'b0001 : 4'b0101;
															assign node10746 = (inp[9]) ? 4'b0111 : 4'b0001;
														assign node10749 = (inp[4]) ? node10753 : node10750;
															assign node10750 = (inp[9]) ? 4'b0001 : 4'b0101;
															assign node10753 = (inp[9]) ? 4'b0101 : 4'b0001;
													assign node10756 = (inp[12]) ? node10762 : node10757;
														assign node10757 = (inp[4]) ? 4'b0011 : node10758;
															assign node10758 = (inp[9]) ? 4'b0011 : 4'b0111;
														assign node10762 = (inp[4]) ? node10764 : 4'b0011;
															assign node10764 = (inp[9]) ? node10766 : 4'b0011;
																assign node10766 = (inp[3]) ? 4'b0101 : 4'b0111;
											assign node10769 = (inp[3]) ? node10799 : node10770;
												assign node10770 = (inp[0]) ? node10784 : node10771;
													assign node10771 = (inp[15]) ? node10777 : node10772;
														assign node10772 = (inp[4]) ? 4'b0101 : node10773;
															assign node10773 = (inp[12]) ? 4'b0011 : 4'b0111;
														assign node10777 = (inp[9]) ? node10781 : node10778;
															assign node10778 = (inp[4]) ? 4'b0001 : 4'b0101;
															assign node10781 = (inp[4]) ? 4'b0111 : 4'b0001;
													assign node10784 = (inp[15]) ? node10792 : node10785;
														assign node10785 = (inp[4]) ? node10789 : node10786;
															assign node10786 = (inp[9]) ? 4'b0001 : 4'b0101;
															assign node10789 = (inp[9]) ? 4'b0111 : 4'b0001;
														assign node10792 = (inp[4]) ? node10796 : node10793;
															assign node10793 = (inp[9]) ? 4'b0011 : 4'b0111;
															assign node10796 = (inp[9]) ? 4'b0101 : 4'b0011;
												assign node10799 = (inp[9]) ? node10821 : node10800;
													assign node10800 = (inp[4]) ? node10808 : node10801;
														assign node10801 = (inp[15]) ? node10805 : node10802;
															assign node10802 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node10805 = (inp[0]) ? 4'b0101 : 4'b0111;
														assign node10808 = (inp[12]) ? node10814 : node10809;
															assign node10809 = (inp[0]) ? node10811 : 4'b0011;
																assign node10811 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node10814 = (inp[15]) ? node10818 : node10815;
																assign node10815 = (inp[0]) ? 4'b0011 : 4'b0001;
																assign node10818 = (inp[0]) ? 4'b0001 : 4'b0011;
													assign node10821 = (inp[4]) ? node10829 : node10822;
														assign node10822 = (inp[0]) ? node10826 : node10823;
															assign node10823 = (inp[15]) ? 4'b0011 : 4'b0001;
															assign node10826 = (inp[15]) ? 4'b0001 : 4'b0011;
														assign node10829 = (inp[0]) ? node10831 : 4'b0101;
															assign node10831 = (inp[15]) ? 4'b0101 : 4'b0111;
										assign node10834 = (inp[15]) ? node10886 : node10835;
											assign node10835 = (inp[0]) ? node10867 : node10836;
												assign node10836 = (inp[3]) ? node10854 : node10837;
													assign node10837 = (inp[12]) ? node10849 : node10838;
														assign node10838 = (inp[5]) ? node10844 : node10839;
															assign node10839 = (inp[9]) ? node10841 : 4'b0010;
																assign node10841 = (inp[4]) ? 4'b0110 : 4'b0010;
															assign node10844 = (inp[9]) ? 4'b0100 : node10845;
																assign node10845 = (inp[4]) ? 4'b0010 : 4'b0110;
														assign node10849 = (inp[9]) ? 4'b0010 : node10850;
															assign node10850 = (inp[4]) ? 4'b0010 : 4'b0110;
													assign node10854 = (inp[5]) ? node10860 : node10855;
														assign node10855 = (inp[4]) ? node10857 : 4'b0010;
															assign node10857 = (inp[9]) ? 4'b0100 : 4'b0010;
														assign node10860 = (inp[12]) ? node10862 : 4'b0000;
															assign node10862 = (inp[4]) ? node10864 : 4'b0100;
																assign node10864 = (inp[9]) ? 4'b0100 : 4'b0000;
												assign node10867 = (inp[4]) ? node10875 : node10868;
													assign node10868 = (inp[9]) ? node10870 : 4'b0100;
														assign node10870 = (inp[3]) ? node10872 : 4'b0000;
															assign node10872 = (inp[5]) ? 4'b0010 : 4'b0000;
													assign node10875 = (inp[9]) ? node10881 : node10876;
														assign node10876 = (inp[5]) ? node10878 : 4'b0000;
															assign node10878 = (inp[3]) ? 4'b0010 : 4'b0000;
														assign node10881 = (inp[5]) ? 4'b0110 : node10882;
															assign node10882 = (inp[12]) ? 4'b0110 : 4'b0100;
											assign node10886 = (inp[0]) ? node10920 : node10887;
												assign node10887 = (inp[5]) ? node10903 : node10888;
													assign node10888 = (inp[12]) ? node10896 : node10889;
														assign node10889 = (inp[3]) ? 4'b0110 : node10890;
															assign node10890 = (inp[9]) ? 4'b0000 : node10891;
																assign node10891 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node10896 = (inp[3]) ? node10898 : 4'b0100;
															assign node10898 = (inp[9]) ? 4'b0000 : node10899;
																assign node10899 = (inp[4]) ? 4'b0000 : 4'b0100;
													assign node10903 = (inp[3]) ? node10911 : node10904;
														assign node10904 = (inp[4]) ? node10908 : node10905;
															assign node10905 = (inp[9]) ? 4'b0000 : 4'b0100;
															assign node10908 = (inp[9]) ? 4'b0110 : 4'b0000;
														assign node10911 = (inp[12]) ? node10915 : node10912;
															assign node10912 = (inp[4]) ? 4'b0010 : 4'b0110;
															assign node10915 = (inp[4]) ? 4'b0110 : node10916;
																assign node10916 = (inp[9]) ? 4'b0010 : 4'b0110;
												assign node10920 = (inp[3]) ? node10936 : node10921;
													assign node10921 = (inp[12]) ? node10927 : node10922;
														assign node10922 = (inp[4]) ? node10924 : 4'b0010;
															assign node10924 = (inp[9]) ? 4'b0110 : 4'b0010;
														assign node10927 = (inp[5]) ? node10933 : node10928;
															assign node10928 = (inp[9]) ? 4'b0110 : node10929;
																assign node10929 = (inp[4]) ? 4'b0010 : 4'b0110;
															assign node10933 = (inp[9]) ? 4'b0100 : 4'b0110;
													assign node10936 = (inp[5]) ? node10942 : node10937;
														assign node10937 = (inp[4]) ? node10939 : 4'b0010;
															assign node10939 = (inp[9]) ? 4'b0100 : 4'b0010;
														assign node10942 = (inp[12]) ? node10950 : node10943;
															assign node10943 = (inp[4]) ? node10947 : node10944;
																assign node10944 = (inp[9]) ? 4'b0000 : 4'b0100;
																assign node10947 = (inp[9]) ? 4'b0100 : 4'b0000;
															assign node10950 = (inp[4]) ? node10954 : node10951;
																assign node10951 = (inp[9]) ? 4'b0000 : 4'b0100;
																assign node10954 = (inp[9]) ? 4'b0100 : 4'b0000;
									assign node10957 = (inp[9]) ? node11053 : node10958;
										assign node10958 = (inp[4]) ? node11002 : node10959;
											assign node10959 = (inp[5]) ? node10967 : node10960;
												assign node10960 = (inp[0]) ? node10964 : node10961;
													assign node10961 = (inp[15]) ? 4'b0100 : 4'b0110;
													assign node10964 = (inp[15]) ? 4'b0110 : 4'b0100;
												assign node10967 = (inp[14]) ? node10985 : node10968;
													assign node10968 = (inp[3]) ? node10978 : node10969;
														assign node10969 = (inp[12]) ? node10973 : node10970;
															assign node10970 = (inp[0]) ? 4'b0100 : 4'b0110;
															assign node10973 = (inp[15]) ? node10975 : 4'b0110;
																assign node10975 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node10978 = (inp[15]) ? node10982 : node10979;
															assign node10979 = (inp[0]) ? 4'b0110 : 4'b0100;
															assign node10982 = (inp[0]) ? 4'b0100 : 4'b0110;
													assign node10985 = (inp[3]) ? node10993 : node10986;
														assign node10986 = (inp[0]) ? node10990 : node10987;
															assign node10987 = (inp[15]) ? 4'b0100 : 4'b0110;
															assign node10990 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node10993 = (inp[12]) ? node10999 : node10994;
															assign node10994 = (inp[0]) ? 4'b0110 : node10995;
																assign node10995 = (inp[15]) ? 4'b0110 : 4'b0100;
															assign node10999 = (inp[0]) ? 4'b0100 : 4'b0110;
											assign node11002 = (inp[14]) ? node11032 : node11003;
												assign node11003 = (inp[5]) ? node11011 : node11004;
													assign node11004 = (inp[15]) ? node11008 : node11005;
														assign node11005 = (inp[0]) ? 4'b0000 : 4'b0010;
														assign node11008 = (inp[0]) ? 4'b0010 : 4'b0000;
													assign node11011 = (inp[3]) ? node11021 : node11012;
														assign node11012 = (inp[12]) ? node11014 : 4'b0000;
															assign node11014 = (inp[15]) ? node11018 : node11015;
																assign node11015 = (inp[0]) ? 4'b0000 : 4'b0010;
																assign node11018 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node11021 = (inp[12]) ? node11027 : node11022;
															assign node11022 = (inp[0]) ? node11024 : 4'b0010;
																assign node11024 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node11027 = (inp[15]) ? node11029 : 4'b0000;
																assign node11029 = (inp[0]) ? 4'b0000 : 4'b0010;
												assign node11032 = (inp[15]) ? node11042 : node11033;
													assign node11033 = (inp[0]) ? node11037 : node11034;
														assign node11034 = (inp[3]) ? 4'b0000 : 4'b0010;
														assign node11037 = (inp[3]) ? node11039 : 4'b0000;
															assign node11039 = (inp[5]) ? 4'b0010 : 4'b0000;
													assign node11042 = (inp[0]) ? node11048 : node11043;
														assign node11043 = (inp[5]) ? node11045 : 4'b0000;
															assign node11045 = (inp[3]) ? 4'b0010 : 4'b0000;
														assign node11048 = (inp[5]) ? node11050 : 4'b0010;
															assign node11050 = (inp[3]) ? 4'b0000 : 4'b0010;
										assign node11053 = (inp[4]) ? node11105 : node11054;
											assign node11054 = (inp[5]) ? node11084 : node11055;
												assign node11055 = (inp[3]) ? node11071 : node11056;
													assign node11056 = (inp[14]) ? node11064 : node11057;
														assign node11057 = (inp[0]) ? node11061 : node11058;
															assign node11058 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node11061 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node11064 = (inp[15]) ? node11068 : node11065;
															assign node11065 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node11068 = (inp[0]) ? 4'b0010 : 4'b0000;
													assign node11071 = (inp[14]) ? node11079 : node11072;
														assign node11072 = (inp[12]) ? node11074 : 4'b0000;
															assign node11074 = (inp[0]) ? node11076 : 4'b0010;
																assign node11076 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node11079 = (inp[12]) ? 4'b0000 : node11080;
															assign node11080 = (inp[15]) ? 4'b0000 : 4'b0010;
												assign node11084 = (inp[3]) ? node11092 : node11085;
													assign node11085 = (inp[15]) ? node11089 : node11086;
														assign node11086 = (inp[0]) ? 4'b0000 : 4'b0010;
														assign node11089 = (inp[0]) ? 4'b0010 : 4'b0000;
													assign node11092 = (inp[12]) ? node11098 : node11093;
														assign node11093 = (inp[15]) ? node11095 : 4'b0010;
															assign node11095 = (inp[0]) ? 4'b0000 : 4'b0010;
														assign node11098 = (inp[15]) ? node11102 : node11099;
															assign node11099 = (inp[0]) ? 4'b0010 : 4'b0000;
															assign node11102 = (inp[0]) ? 4'b0000 : 4'b0010;
											assign node11105 = (inp[3]) ? node11129 : node11106;
												assign node11106 = (inp[14]) ? node11116 : node11107;
													assign node11107 = (inp[15]) ? 4'b0100 : node11108;
														assign node11108 = (inp[5]) ? node11112 : node11109;
															assign node11109 = (inp[0]) ? 4'b0100 : 4'b0110;
															assign node11112 = (inp[0]) ? 4'b0110 : 4'b0100;
													assign node11116 = (inp[5]) ? node11122 : node11117;
														assign node11117 = (inp[0]) ? 4'b0110 : node11118;
															assign node11118 = (inp[15]) ? 4'b0100 : 4'b0110;
														assign node11122 = (inp[15]) ? node11126 : node11123;
															assign node11123 = (inp[0]) ? 4'b0110 : 4'b0100;
															assign node11126 = (inp[0]) ? 4'b0100 : 4'b0110;
												assign node11129 = (inp[0]) ? node11133 : node11130;
													assign node11130 = (inp[15]) ? 4'b0110 : 4'b0100;
													assign node11133 = (inp[15]) ? 4'b0100 : 4'b0110;
								assign node11136 = (inp[2]) ? node11432 : node11137;
									assign node11137 = (inp[14]) ? node11271 : node11138;
										assign node11138 = (inp[12]) ? node11196 : node11139;
											assign node11139 = (inp[9]) ? node11163 : node11140;
												assign node11140 = (inp[4]) ? node11152 : node11141;
													assign node11141 = (inp[15]) ? 4'b0110 : node11142;
														assign node11142 = (inp[5]) ? node11146 : node11143;
															assign node11143 = (inp[3]) ? 4'b0110 : 4'b0100;
															assign node11146 = (inp[0]) ? 4'b0110 : node11147;
																assign node11147 = (inp[3]) ? 4'b0100 : 4'b0110;
													assign node11152 = (inp[15]) ? node11158 : node11153;
														assign node11153 = (inp[0]) ? node11155 : 4'b0010;
															assign node11155 = (inp[5]) ? 4'b0010 : 4'b0000;
														assign node11158 = (inp[5]) ? 4'b0000 : node11159;
															assign node11159 = (inp[0]) ? 4'b0010 : 4'b0000;
												assign node11163 = (inp[4]) ? node11175 : node11164;
													assign node11164 = (inp[0]) ? node11170 : node11165;
														assign node11165 = (inp[15]) ? 4'b0000 : node11166;
															assign node11166 = (inp[5]) ? 4'b0000 : 4'b0010;
														assign node11170 = (inp[15]) ? 4'b0010 : node11171;
															assign node11171 = (inp[5]) ? 4'b0010 : 4'b0000;
													assign node11175 = (inp[5]) ? node11183 : node11176;
														assign node11176 = (inp[15]) ? node11178 : 4'b0100;
															assign node11178 = (inp[3]) ? 4'b0100 : node11179;
																assign node11179 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node11183 = (inp[3]) ? node11189 : node11184;
															assign node11184 = (inp[0]) ? 4'b0110 : node11185;
																assign node11185 = (inp[15]) ? 4'b0110 : 4'b0100;
															assign node11189 = (inp[0]) ? node11193 : node11190;
																assign node11190 = (inp[15]) ? 4'b0110 : 4'b0100;
																assign node11193 = (inp[15]) ? 4'b0100 : 4'b0110;
											assign node11196 = (inp[3]) ? node11232 : node11197;
												assign node11197 = (inp[15]) ? node11215 : node11198;
													assign node11198 = (inp[0]) ? node11204 : node11199;
														assign node11199 = (inp[4]) ? 4'b0010 : node11200;
															assign node11200 = (inp[9]) ? 4'b0010 : 4'b0110;
														assign node11204 = (inp[5]) ? node11210 : node11205;
															assign node11205 = (inp[4]) ? node11207 : 4'b0000;
																assign node11207 = (inp[9]) ? 4'b0100 : 4'b0000;
															assign node11210 = (inp[4]) ? 4'b0000 : node11211;
																assign node11211 = (inp[9]) ? 4'b0000 : 4'b0100;
													assign node11215 = (inp[0]) ? node11225 : node11216;
														assign node11216 = (inp[9]) ? node11220 : node11217;
															assign node11217 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node11220 = (inp[4]) ? node11222 : 4'b0000;
																assign node11222 = (inp[5]) ? 4'b0110 : 4'b0100;
														assign node11225 = (inp[4]) ? node11229 : node11226;
															assign node11226 = (inp[9]) ? 4'b0010 : 4'b0110;
															assign node11229 = (inp[9]) ? 4'b0100 : 4'b0010;
												assign node11232 = (inp[5]) ? node11250 : node11233;
													assign node11233 = (inp[0]) ? node11241 : node11234;
														assign node11234 = (inp[15]) ? node11236 : 4'b0100;
															assign node11236 = (inp[4]) ? 4'b0000 : node11237;
																assign node11237 = (inp[9]) ? 4'b0000 : 4'b0100;
														assign node11241 = (inp[4]) ? node11247 : node11242;
															assign node11242 = (inp[9]) ? node11244 : 4'b0100;
																assign node11244 = (inp[15]) ? 4'b0010 : 4'b0000;
															assign node11247 = (inp[15]) ? 4'b0100 : 4'b0110;
													assign node11250 = (inp[15]) ? node11258 : node11251;
														assign node11251 = (inp[0]) ? node11253 : 4'b0000;
															assign node11253 = (inp[9]) ? 4'b0010 : node11254;
																assign node11254 = (inp[4]) ? 4'b0010 : 4'b0110;
														assign node11258 = (inp[0]) ? node11264 : node11259;
															assign node11259 = (inp[9]) ? node11261 : 4'b0010;
																assign node11261 = (inp[4]) ? 4'b0110 : 4'b0010;
															assign node11264 = (inp[4]) ? node11268 : node11265;
																assign node11265 = (inp[9]) ? 4'b0000 : 4'b0100;
																assign node11268 = (inp[9]) ? 4'b0100 : 4'b0000;
										assign node11271 = (inp[5]) ? node11357 : node11272;
											assign node11272 = (inp[0]) ? node11318 : node11273;
												assign node11273 = (inp[15]) ? node11295 : node11274;
													assign node11274 = (inp[3]) ? node11282 : node11275;
														assign node11275 = (inp[12]) ? node11277 : 4'b1011;
															assign node11277 = (inp[4]) ? node11279 : 4'b1011;
																assign node11279 = (inp[9]) ? 4'b1011 : 4'b1111;
														assign node11282 = (inp[9]) ? node11290 : node11283;
															assign node11283 = (inp[4]) ? node11287 : node11284;
																assign node11284 = (inp[12]) ? 4'b1011 : 4'b1111;
																assign node11287 = (inp[12]) ? 4'b1101 : 4'b1011;
															assign node11290 = (inp[4]) ? node11292 : 4'b1101;
																assign node11292 = (inp[12]) ? 4'b1001 : 4'b1101;
													assign node11295 = (inp[3]) ? node11311 : node11296;
														assign node11296 = (inp[4]) ? node11304 : node11297;
															assign node11297 = (inp[9]) ? node11301 : node11298;
																assign node11298 = (inp[12]) ? 4'b1001 : 4'b1101;
																assign node11301 = (inp[12]) ? 4'b1101 : 4'b1001;
															assign node11304 = (inp[12]) ? node11308 : node11305;
																assign node11305 = (inp[9]) ? 4'b1101 : 4'b1001;
																assign node11308 = (inp[9]) ? 4'b1001 : 4'b1101;
														assign node11311 = (inp[12]) ? node11315 : node11312;
															assign node11312 = (inp[4]) ? 4'b1001 : 4'b1101;
															assign node11315 = (inp[9]) ? 4'b1011 : 4'b1111;
												assign node11318 = (inp[15]) ? node11338 : node11319;
													assign node11319 = (inp[3]) ? node11331 : node11320;
														assign node11320 = (inp[12]) ? node11326 : node11321;
															assign node11321 = (inp[9]) ? node11323 : 4'b1101;
																assign node11323 = (inp[4]) ? 4'b1101 : 4'b1001;
															assign node11326 = (inp[9]) ? node11328 : 4'b1001;
																assign node11328 = (inp[4]) ? 4'b1001 : 4'b1101;
														assign node11331 = (inp[4]) ? 4'b1111 : node11332;
															assign node11332 = (inp[9]) ? 4'b1111 : node11333;
																assign node11333 = (inp[12]) ? 4'b1001 : 4'b1101;
													assign node11338 = (inp[3]) ? node11352 : node11339;
														assign node11339 = (inp[9]) ? node11345 : node11340;
															assign node11340 = (inp[4]) ? 4'b1111 : node11341;
																assign node11341 = (inp[12]) ? 4'b1011 : 4'b1111;
															assign node11345 = (inp[12]) ? node11349 : node11346;
																assign node11346 = (inp[4]) ? 4'b1111 : 4'b1011;
																assign node11349 = (inp[4]) ? 4'b1011 : 4'b1111;
														assign node11352 = (inp[12]) ? node11354 : 4'b1011;
															assign node11354 = (inp[4]) ? 4'b1001 : 4'b1101;
											assign node11357 = (inp[15]) ? node11397 : node11358;
												assign node11358 = (inp[0]) ? node11378 : node11359;
													assign node11359 = (inp[3]) ? node11371 : node11360;
														assign node11360 = (inp[12]) ? node11366 : node11361;
															assign node11361 = (inp[9]) ? 4'b1011 : node11362;
																assign node11362 = (inp[4]) ? 4'b1011 : 4'b1111;
															assign node11366 = (inp[4]) ? node11368 : 4'b1011;
																assign node11368 = (inp[9]) ? 4'b1001 : 4'b1101;
														assign node11371 = (inp[4]) ? node11373 : 4'b1001;
															assign node11373 = (inp[9]) ? 4'b1001 : node11374;
																assign node11374 = (inp[12]) ? 4'b1101 : 4'b1001;
													assign node11378 = (inp[3]) ? node11388 : node11379;
														assign node11379 = (inp[9]) ? node11381 : 4'b1001;
															assign node11381 = (inp[12]) ? node11385 : node11382;
																assign node11382 = (inp[4]) ? 4'b1111 : 4'b1001;
																assign node11385 = (inp[4]) ? 4'b1011 : 4'b1111;
														assign node11388 = (inp[12]) ? 4'b1011 : node11389;
															assign node11389 = (inp[9]) ? node11393 : node11390;
																assign node11390 = (inp[4]) ? 4'b1011 : 4'b1111;
																assign node11393 = (inp[4]) ? 4'b1111 : 4'b1011;
												assign node11397 = (inp[0]) ? node11411 : node11398;
													assign node11398 = (inp[12]) ? node11404 : node11399;
														assign node11399 = (inp[4]) ? 4'b1111 : node11400;
															assign node11400 = (inp[3]) ? 4'b1111 : 4'b1001;
														assign node11404 = (inp[4]) ? node11408 : node11405;
															assign node11405 = (inp[9]) ? 4'b1111 : 4'b1011;
															assign node11408 = (inp[9]) ? 4'b1011 : 4'b1111;
													assign node11411 = (inp[3]) ? node11423 : node11412;
														assign node11412 = (inp[9]) ? node11418 : node11413;
															assign node11413 = (inp[4]) ? 4'b1011 : node11414;
																assign node11414 = (inp[12]) ? 4'b1011 : 4'b1111;
															assign node11418 = (inp[12]) ? 4'b1101 : node11419;
																assign node11419 = (inp[4]) ? 4'b1101 : 4'b1011;
														assign node11423 = (inp[9]) ? node11425 : 4'b1101;
															assign node11425 = (inp[12]) ? node11429 : node11426;
																assign node11426 = (inp[4]) ? 4'b1101 : 4'b1001;
																assign node11429 = (inp[4]) ? 4'b1001 : 4'b1101;
									assign node11432 = (inp[15]) ? node11562 : node11433;
										assign node11433 = (inp[0]) ? node11499 : node11434;
											assign node11434 = (inp[5]) ? node11466 : node11435;
												assign node11435 = (inp[3]) ? node11449 : node11436;
													assign node11436 = (inp[4]) ? node11442 : node11437;
														assign node11437 = (inp[12]) ? 4'b1111 : node11438;
															assign node11438 = (inp[9]) ? 4'b1011 : 4'b1111;
														assign node11442 = (inp[12]) ? node11446 : node11443;
															assign node11443 = (inp[14]) ? 4'b1111 : 4'b1011;
															assign node11446 = (inp[14]) ? 4'b1011 : 4'b1111;
													assign node11449 = (inp[9]) ? node11459 : node11450;
														assign node11450 = (inp[14]) ? node11456 : node11451;
															assign node11451 = (inp[12]) ? 4'b1011 : node11452;
																assign node11452 = (inp[4]) ? 4'b1011 : 4'b1111;
															assign node11456 = (inp[4]) ? 4'b1101 : 4'b1111;
														assign node11459 = (inp[14]) ? node11461 : 4'b1101;
															assign node11461 = (inp[4]) ? node11463 : 4'b1011;
																assign node11463 = (inp[12]) ? 4'b1001 : 4'b1101;
												assign node11466 = (inp[9]) ? node11480 : node11467;
													assign node11467 = (inp[3]) ? node11473 : node11468;
														assign node11468 = (inp[4]) ? node11470 : 4'b1011;
															assign node11470 = (inp[12]) ? 4'b1101 : 4'b1011;
														assign node11473 = (inp[4]) ? node11477 : node11474;
															assign node11474 = (inp[12]) ? 4'b1001 : 4'b1101;
															assign node11477 = (inp[12]) ? 4'b1101 : 4'b1001;
													assign node11480 = (inp[14]) ? node11492 : node11481;
														assign node11481 = (inp[3]) ? node11487 : node11482;
															assign node11482 = (inp[4]) ? node11484 : 4'b1101;
																assign node11484 = (inp[12]) ? 4'b1001 : 4'b1101;
															assign node11487 = (inp[4]) ? 4'b1101 : node11488;
																assign node11488 = (inp[12]) ? 4'b1101 : 4'b1001;
														assign node11492 = (inp[12]) ? node11496 : node11493;
															assign node11493 = (inp[4]) ? 4'b1101 : 4'b1001;
															assign node11496 = (inp[4]) ? 4'b1001 : 4'b1101;
											assign node11499 = (inp[5]) ? node11539 : node11500;
												assign node11500 = (inp[3]) ? node11522 : node11501;
													assign node11501 = (inp[9]) ? node11507 : node11502;
														assign node11502 = (inp[14]) ? node11504 : 4'b1101;
															assign node11504 = (inp[12]) ? 4'b1101 : 4'b1001;
														assign node11507 = (inp[14]) ? node11515 : node11508;
															assign node11508 = (inp[4]) ? node11512 : node11509;
																assign node11509 = (inp[12]) ? 4'b1101 : 4'b1001;
																assign node11512 = (inp[12]) ? 4'b1001 : 4'b1101;
															assign node11515 = (inp[12]) ? node11519 : node11516;
																assign node11516 = (inp[4]) ? 4'b1101 : 4'b1001;
																assign node11519 = (inp[4]) ? 4'b1001 : 4'b1101;
													assign node11522 = (inp[9]) ? node11530 : node11523;
														assign node11523 = (inp[12]) ? node11527 : node11524;
															assign node11524 = (inp[4]) ? 4'b1001 : 4'b1101;
															assign node11527 = (inp[4]) ? 4'b1111 : 4'b1001;
														assign node11530 = (inp[14]) ? node11534 : node11531;
															assign node11531 = (inp[12]) ? 4'b1011 : 4'b1001;
															assign node11534 = (inp[4]) ? 4'b1111 : node11535;
																assign node11535 = (inp[12]) ? 4'b1111 : 4'b1001;
												assign node11539 = (inp[9]) ? node11555 : node11540;
													assign node11540 = (inp[3]) ? node11550 : node11541;
														assign node11541 = (inp[14]) ? 4'b1111 : node11542;
															assign node11542 = (inp[4]) ? node11546 : node11543;
																assign node11543 = (inp[12]) ? 4'b1001 : 4'b1101;
																assign node11546 = (inp[12]) ? 4'b1111 : 4'b1001;
														assign node11550 = (inp[14]) ? node11552 : 4'b1111;
															assign node11552 = (inp[4]) ? 4'b1011 : 4'b1111;
													assign node11555 = (inp[12]) ? node11559 : node11556;
														assign node11556 = (inp[4]) ? 4'b1111 : 4'b1011;
														assign node11559 = (inp[4]) ? 4'b1011 : 4'b1111;
										assign node11562 = (inp[5]) ? node11634 : node11563;
											assign node11563 = (inp[0]) ? node11603 : node11564;
												assign node11564 = (inp[3]) ? node11588 : node11565;
													assign node11565 = (inp[14]) ? node11579 : node11566;
														assign node11566 = (inp[9]) ? node11572 : node11567;
															assign node11567 = (inp[4]) ? node11569 : 4'b1101;
																assign node11569 = (inp[12]) ? 4'b1101 : 4'b1001;
															assign node11572 = (inp[12]) ? node11576 : node11573;
																assign node11573 = (inp[4]) ? 4'b1101 : 4'b1001;
																assign node11576 = (inp[4]) ? 4'b1001 : 4'b1101;
														assign node11579 = (inp[12]) ? 4'b1001 : node11580;
															assign node11580 = (inp[9]) ? node11584 : node11581;
																assign node11581 = (inp[4]) ? 4'b1001 : 4'b1101;
																assign node11584 = (inp[4]) ? 4'b1101 : 4'b1001;
													assign node11588 = (inp[14]) ? node11598 : node11589;
														assign node11589 = (inp[12]) ? 4'b1111 : node11590;
															assign node11590 = (inp[9]) ? node11594 : node11591;
																assign node11591 = (inp[4]) ? 4'b1001 : 4'b1101;
																assign node11594 = (inp[4]) ? 4'b1111 : 4'b1001;
														assign node11598 = (inp[12]) ? node11600 : 4'b1001;
															assign node11600 = (inp[9]) ? 4'b1011 : 4'b1001;
												assign node11603 = (inp[3]) ? node11619 : node11604;
													assign node11604 = (inp[12]) ? node11610 : node11605;
														assign node11605 = (inp[4]) ? 4'b1011 : node11606;
															assign node11606 = (inp[9]) ? 4'b1011 : 4'b1111;
														assign node11610 = (inp[14]) ? 4'b1111 : node11611;
															assign node11611 = (inp[9]) ? node11615 : node11612;
																assign node11612 = (inp[4]) ? 4'b1111 : 4'b1011;
																assign node11615 = (inp[4]) ? 4'b1011 : 4'b1111;
													assign node11619 = (inp[4]) ? node11627 : node11620;
														assign node11620 = (inp[12]) ? node11624 : node11621;
															assign node11621 = (inp[9]) ? 4'b1011 : 4'b1111;
															assign node11624 = (inp[9]) ? 4'b1101 : 4'b1011;
														assign node11627 = (inp[9]) ? node11631 : node11628;
															assign node11628 = (inp[12]) ? 4'b1101 : 4'b1011;
															assign node11631 = (inp[12]) ? 4'b1001 : 4'b1101;
											assign node11634 = (inp[0]) ? node11666 : node11635;
												assign node11635 = (inp[3]) ? node11651 : node11636;
													assign node11636 = (inp[12]) ? node11644 : node11637;
														assign node11637 = (inp[14]) ? node11639 : 4'b1001;
															assign node11639 = (inp[9]) ? 4'b1111 : node11640;
																assign node11640 = (inp[4]) ? 4'b1001 : 4'b1101;
														assign node11644 = (inp[4]) ? node11648 : node11645;
															assign node11645 = (inp[9]) ? 4'b1111 : 4'b1001;
															assign node11648 = (inp[9]) ? 4'b1011 : 4'b1111;
													assign node11651 = (inp[9]) ? node11659 : node11652;
														assign node11652 = (inp[12]) ? node11656 : node11653;
															assign node11653 = (inp[4]) ? 4'b1011 : 4'b1111;
															assign node11656 = (inp[4]) ? 4'b1111 : 4'b1011;
														assign node11659 = (inp[4]) ? node11663 : node11660;
															assign node11660 = (inp[12]) ? 4'b1111 : 4'b1011;
															assign node11663 = (inp[12]) ? 4'b1011 : 4'b1111;
												assign node11666 = (inp[3]) ? node11682 : node11667;
													assign node11667 = (inp[9]) ? node11675 : node11668;
														assign node11668 = (inp[4]) ? node11672 : node11669;
															assign node11669 = (inp[12]) ? 4'b1011 : 4'b1111;
															assign node11672 = (inp[12]) ? 4'b1101 : 4'b1011;
														assign node11675 = (inp[4]) ? node11679 : node11676;
															assign node11676 = (inp[12]) ? 4'b1101 : 4'b1011;
															assign node11679 = (inp[12]) ? 4'b1001 : 4'b1101;
													assign node11682 = (inp[14]) ? node11694 : node11683;
														assign node11683 = (inp[12]) ? node11689 : node11684;
															assign node11684 = (inp[4]) ? 4'b1001 : node11685;
																assign node11685 = (inp[9]) ? 4'b1001 : 4'b1101;
															assign node11689 = (inp[4]) ? 4'b1101 : node11690;
																assign node11690 = (inp[9]) ? 4'b1101 : 4'b1001;
														assign node11694 = (inp[12]) ? node11700 : node11695;
															assign node11695 = (inp[9]) ? 4'b1101 : node11696;
																assign node11696 = (inp[4]) ? 4'b1001 : 4'b1101;
															assign node11700 = (inp[4]) ? node11702 : 4'b1001;
																assign node11702 = (inp[9]) ? 4'b1001 : 4'b1101;
							assign node11705 = (inp[7]) ? node12193 : node11706;
								assign node11706 = (inp[2]) ? node11972 : node11707;
									assign node11707 = (inp[14]) ? node11823 : node11708;
										assign node11708 = (inp[3]) ? node11762 : node11709;
											assign node11709 = (inp[0]) ? node11737 : node11710;
												assign node11710 = (inp[15]) ? node11726 : node11711;
													assign node11711 = (inp[5]) ? node11719 : node11712;
														assign node11712 = (inp[4]) ? node11716 : node11713;
															assign node11713 = (inp[9]) ? 4'b0010 : 4'b0110;
															assign node11716 = (inp[9]) ? 4'b0110 : 4'b0010;
														assign node11719 = (inp[9]) ? node11723 : node11720;
															assign node11720 = (inp[4]) ? 4'b0010 : 4'b0110;
															assign node11723 = (inp[4]) ? 4'b0100 : 4'b0010;
													assign node11726 = (inp[5]) ? node11732 : node11727;
														assign node11727 = (inp[4]) ? 4'b0100 : node11728;
															assign node11728 = (inp[9]) ? 4'b0000 : 4'b0100;
														assign node11732 = (inp[4]) ? 4'b0000 : node11733;
															assign node11733 = (inp[9]) ? 4'b0000 : 4'b0100;
												assign node11737 = (inp[15]) ? node11755 : node11738;
													assign node11738 = (inp[5]) ? node11750 : node11739;
														assign node11739 = (inp[12]) ? node11745 : node11740;
															assign node11740 = (inp[4]) ? 4'b0100 : node11741;
																assign node11741 = (inp[9]) ? 4'b0000 : 4'b0100;
															assign node11745 = (inp[9]) ? 4'b0000 : node11746;
																assign node11746 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node11750 = (inp[9]) ? 4'b0110 : node11751;
															assign node11751 = (inp[4]) ? 4'b0000 : 4'b0100;
													assign node11755 = (inp[9]) ? node11759 : node11756;
														assign node11756 = (inp[4]) ? 4'b0010 : 4'b0110;
														assign node11759 = (inp[4]) ? 4'b0110 : 4'b0010;
											assign node11762 = (inp[15]) ? node11788 : node11763;
												assign node11763 = (inp[9]) ? node11779 : node11764;
													assign node11764 = (inp[4]) ? node11766 : 4'b0110;
														assign node11766 = (inp[12]) ? node11772 : node11767;
															assign node11767 = (inp[5]) ? 4'b0000 : node11768;
																assign node11768 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node11772 = (inp[0]) ? node11776 : node11773;
																assign node11773 = (inp[5]) ? 4'b0000 : 4'b0010;
																assign node11776 = (inp[5]) ? 4'b0010 : 4'b0000;
													assign node11779 = (inp[4]) ? node11785 : node11780;
														assign node11780 = (inp[0]) ? node11782 : 4'b0000;
															assign node11782 = (inp[5]) ? 4'b0010 : 4'b0000;
														assign node11785 = (inp[0]) ? 4'b0110 : 4'b0100;
												assign node11788 = (inp[0]) ? node11804 : node11789;
													assign node11789 = (inp[5]) ? node11797 : node11790;
														assign node11790 = (inp[9]) ? node11794 : node11791;
															assign node11791 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node11794 = (inp[4]) ? 4'b0110 : 4'b0000;
														assign node11797 = (inp[4]) ? node11801 : node11798;
															assign node11798 = (inp[9]) ? 4'b0010 : 4'b0110;
															assign node11801 = (inp[9]) ? 4'b0110 : 4'b0010;
													assign node11804 = (inp[5]) ? node11814 : node11805;
														assign node11805 = (inp[12]) ? node11807 : 4'b0010;
															assign node11807 = (inp[4]) ? node11811 : node11808;
																assign node11808 = (inp[9]) ? 4'b0010 : 4'b0110;
																assign node11811 = (inp[9]) ? 4'b0100 : 4'b0010;
														assign node11814 = (inp[12]) ? node11820 : node11815;
															assign node11815 = (inp[4]) ? 4'b0000 : node11816;
																assign node11816 = (inp[9]) ? 4'b0000 : 4'b0100;
															assign node11820 = (inp[4]) ? 4'b0100 : 4'b0000;
										assign node11823 = (inp[3]) ? node11899 : node11824;
											assign node11824 = (inp[4]) ? node11864 : node11825;
												assign node11825 = (inp[0]) ? node11847 : node11826;
													assign node11826 = (inp[15]) ? node11836 : node11827;
														assign node11827 = (inp[9]) ? node11831 : node11828;
															assign node11828 = (inp[5]) ? 4'b1111 : 4'b1011;
															assign node11831 = (inp[12]) ? node11833 : 4'b1011;
																assign node11833 = (inp[5]) ? 4'b1101 : 4'b1111;
														assign node11836 = (inp[5]) ? node11842 : node11837;
															assign node11837 = (inp[12]) ? node11839 : 4'b1101;
																assign node11839 = (inp[9]) ? 4'b1101 : 4'b1001;
															assign node11842 = (inp[9]) ? 4'b1001 : node11843;
																assign node11843 = (inp[12]) ? 4'b1001 : 4'b1101;
													assign node11847 = (inp[15]) ? node11857 : node11848;
														assign node11848 = (inp[12]) ? node11852 : node11849;
															assign node11849 = (inp[9]) ? 4'b1001 : 4'b1101;
															assign node11852 = (inp[5]) ? 4'b1111 : node11853;
																assign node11853 = (inp[9]) ? 4'b1101 : 4'b1001;
														assign node11857 = (inp[9]) ? node11861 : node11858;
															assign node11858 = (inp[12]) ? 4'b1011 : 4'b1111;
															assign node11861 = (inp[12]) ? 4'b1111 : 4'b1011;
												assign node11864 = (inp[5]) ? node11876 : node11865;
													assign node11865 = (inp[12]) ? node11869 : node11866;
														assign node11866 = (inp[9]) ? 4'b1111 : 4'b1011;
														assign node11869 = (inp[9]) ? 4'b1011 : node11870;
															assign node11870 = (inp[15]) ? node11872 : 4'b1111;
																assign node11872 = (inp[0]) ? 4'b1111 : 4'b1101;
													assign node11876 = (inp[15]) ? node11890 : node11877;
														assign node11877 = (inp[0]) ? node11883 : node11878;
															assign node11878 = (inp[12]) ? 4'b1101 : node11879;
																assign node11879 = (inp[9]) ? 4'b1101 : 4'b1011;
															assign node11883 = (inp[12]) ? node11887 : node11884;
																assign node11884 = (inp[9]) ? 4'b1111 : 4'b1001;
																assign node11887 = (inp[9]) ? 4'b1011 : 4'b1111;
														assign node11890 = (inp[0]) ? node11894 : node11891;
															assign node11891 = (inp[12]) ? 4'b1011 : 4'b1001;
															assign node11894 = (inp[9]) ? node11896 : 4'b1011;
																assign node11896 = (inp[12]) ? 4'b1001 : 4'b1101;
											assign node11899 = (inp[12]) ? node11937 : node11900;
												assign node11900 = (inp[5]) ? node11922 : node11901;
													assign node11901 = (inp[4]) ? node11909 : node11902;
														assign node11902 = (inp[9]) ? node11904 : 4'b1101;
															assign node11904 = (inp[0]) ? node11906 : 4'b1001;
																assign node11906 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node11909 = (inp[9]) ? node11917 : node11910;
															assign node11910 = (inp[15]) ? node11914 : node11911;
																assign node11911 = (inp[0]) ? 4'b1001 : 4'b1011;
																assign node11914 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node11917 = (inp[0]) ? node11919 : 4'b1111;
																assign node11919 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node11922 = (inp[9]) ? node11930 : node11923;
														assign node11923 = (inp[4]) ? 4'b1011 : node11924;
															assign node11924 = (inp[15]) ? node11926 : 4'b1111;
																assign node11926 = (inp[0]) ? 4'b1101 : 4'b1111;
														assign node11930 = (inp[4]) ? 4'b1101 : node11931;
															assign node11931 = (inp[0]) ? 4'b1011 : node11932;
																assign node11932 = (inp[15]) ? 4'b1011 : 4'b1001;
												assign node11937 = (inp[15]) ? node11959 : node11938;
													assign node11938 = (inp[0]) ? node11950 : node11939;
														assign node11939 = (inp[5]) ? node11945 : node11940;
															assign node11940 = (inp[9]) ? 4'b1101 : node11941;
																assign node11941 = (inp[4]) ? 4'b1101 : 4'b1011;
															assign node11945 = (inp[9]) ? 4'b1001 : node11946;
																assign node11946 = (inp[4]) ? 4'b1101 : 4'b1001;
														assign node11950 = (inp[5]) ? node11954 : node11951;
															assign node11951 = (inp[4]) ? 4'b1111 : 4'b1001;
															assign node11954 = (inp[9]) ? node11956 : 4'b1011;
																assign node11956 = (inp[4]) ? 4'b1011 : 4'b1111;
													assign node11959 = (inp[0]) ? node11965 : node11960;
														assign node11960 = (inp[4]) ? node11962 : 4'b1001;
															assign node11962 = (inp[9]) ? 4'b1011 : 4'b1111;
														assign node11965 = (inp[4]) ? node11969 : node11966;
															assign node11966 = (inp[9]) ? 4'b1101 : 4'b1001;
															assign node11969 = (inp[9]) ? 4'b1001 : 4'b1101;
									assign node11972 = (inp[15]) ? node12084 : node11973;
										assign node11973 = (inp[9]) ? node12027 : node11974;
											assign node11974 = (inp[0]) ? node12004 : node11975;
												assign node11975 = (inp[5]) ? node11991 : node11976;
													assign node11976 = (inp[14]) ? node11982 : node11977;
														assign node11977 = (inp[4]) ? 4'b1011 : node11978;
															assign node11978 = (inp[12]) ? 4'b1011 : 4'b1111;
														assign node11982 = (inp[12]) ? node11986 : node11983;
															assign node11983 = (inp[4]) ? 4'b1011 : 4'b1111;
															assign node11986 = (inp[3]) ? 4'b1101 : node11987;
																assign node11987 = (inp[4]) ? 4'b1111 : 4'b1011;
													assign node11991 = (inp[3]) ? node11999 : node11992;
														assign node11992 = (inp[12]) ? node11996 : node11993;
															assign node11993 = (inp[4]) ? 4'b1011 : 4'b1111;
															assign node11996 = (inp[4]) ? 4'b1101 : 4'b1011;
														assign node11999 = (inp[12]) ? node12001 : 4'b1101;
															assign node12001 = (inp[4]) ? 4'b1101 : 4'b1001;
												assign node12004 = (inp[5]) ? node12014 : node12005;
													assign node12005 = (inp[4]) ? node12009 : node12006;
														assign node12006 = (inp[12]) ? 4'b1001 : 4'b1101;
														assign node12009 = (inp[12]) ? node12011 : 4'b1001;
															assign node12011 = (inp[3]) ? 4'b1111 : 4'b1101;
													assign node12014 = (inp[3]) ? node12020 : node12015;
														assign node12015 = (inp[4]) ? 4'b1111 : node12016;
															assign node12016 = (inp[12]) ? 4'b1001 : 4'b1101;
														assign node12020 = (inp[4]) ? node12024 : node12021;
															assign node12021 = (inp[12]) ? 4'b1011 : 4'b1111;
															assign node12024 = (inp[12]) ? 4'b1111 : 4'b1011;
											assign node12027 = (inp[0]) ? node12055 : node12028;
												assign node12028 = (inp[5]) ? node12040 : node12029;
													assign node12029 = (inp[3]) ? node12035 : node12030;
														assign node12030 = (inp[14]) ? 4'b1011 : node12031;
															assign node12031 = (inp[4]) ? 4'b1011 : 4'b1111;
														assign node12035 = (inp[4]) ? node12037 : 4'b1011;
															assign node12037 = (inp[12]) ? 4'b1001 : 4'b1101;
													assign node12040 = (inp[3]) ? node12048 : node12041;
														assign node12041 = (inp[4]) ? node12045 : node12042;
															assign node12042 = (inp[12]) ? 4'b1101 : 4'b1011;
															assign node12045 = (inp[12]) ? 4'b1001 : 4'b1101;
														assign node12048 = (inp[4]) ? node12052 : node12049;
															assign node12049 = (inp[12]) ? 4'b1101 : 4'b1001;
															assign node12052 = (inp[12]) ? 4'b1001 : 4'b1101;
												assign node12055 = (inp[3]) ? node12067 : node12056;
													assign node12056 = (inp[5]) ? node12062 : node12057;
														assign node12057 = (inp[14]) ? node12059 : 4'b1001;
															assign node12059 = (inp[12]) ? 4'b1001 : 4'b1101;
														assign node12062 = (inp[12]) ? node12064 : 4'b1001;
															assign node12064 = (inp[4]) ? 4'b1011 : 4'b1111;
													assign node12067 = (inp[14]) ? node12075 : node12068;
														assign node12068 = (inp[4]) ? node12072 : node12069;
															assign node12069 = (inp[12]) ? 4'b1111 : 4'b1011;
															assign node12072 = (inp[12]) ? 4'b1011 : 4'b1111;
														assign node12075 = (inp[12]) ? node12081 : node12076;
															assign node12076 = (inp[5]) ? node12078 : 4'b1001;
																assign node12078 = (inp[4]) ? 4'b1111 : 4'b1011;
															assign node12081 = (inp[4]) ? 4'b1011 : 4'b1111;
										assign node12084 = (inp[12]) ? node12144 : node12085;
											assign node12085 = (inp[0]) ? node12119 : node12086;
												assign node12086 = (inp[3]) ? node12106 : node12087;
													assign node12087 = (inp[5]) ? node12099 : node12088;
														assign node12088 = (inp[14]) ? node12094 : node12089;
															assign node12089 = (inp[9]) ? 4'b1001 : node12090;
																assign node12090 = (inp[4]) ? 4'b1001 : 4'b1101;
															assign node12094 = (inp[9]) ? node12096 : 4'b1001;
																assign node12096 = (inp[4]) ? 4'b1101 : 4'b1001;
														assign node12099 = (inp[4]) ? node12103 : node12100;
															assign node12100 = (inp[9]) ? 4'b1001 : 4'b1101;
															assign node12103 = (inp[9]) ? 4'b1111 : 4'b1001;
													assign node12106 = (inp[5]) ? node12112 : node12107;
														assign node12107 = (inp[9]) ? 4'b1111 : node12108;
															assign node12108 = (inp[4]) ? 4'b1001 : 4'b1101;
														assign node12112 = (inp[9]) ? node12116 : node12113;
															assign node12113 = (inp[14]) ? 4'b1111 : 4'b1011;
															assign node12116 = (inp[4]) ? 4'b1111 : 4'b1011;
												assign node12119 = (inp[5]) ? node12129 : node12120;
													assign node12120 = (inp[4]) ? node12124 : node12121;
														assign node12121 = (inp[9]) ? 4'b1011 : 4'b1111;
														assign node12124 = (inp[9]) ? node12126 : 4'b1011;
															assign node12126 = (inp[3]) ? 4'b1101 : 4'b1111;
													assign node12129 = (inp[3]) ? node12137 : node12130;
														assign node12130 = (inp[9]) ? node12134 : node12131;
															assign node12131 = (inp[4]) ? 4'b1011 : 4'b1111;
															assign node12134 = (inp[4]) ? 4'b1101 : 4'b1011;
														assign node12137 = (inp[4]) ? node12141 : node12138;
															assign node12138 = (inp[9]) ? 4'b1001 : 4'b1101;
															assign node12141 = (inp[9]) ? 4'b1101 : 4'b1001;
											assign node12144 = (inp[0]) ? node12168 : node12145;
												assign node12145 = (inp[3]) ? node12161 : node12146;
													assign node12146 = (inp[5]) ? node12154 : node12147;
														assign node12147 = (inp[4]) ? node12151 : node12148;
															assign node12148 = (inp[9]) ? 4'b1101 : 4'b1001;
															assign node12151 = (inp[9]) ? 4'b1001 : 4'b1101;
														assign node12154 = (inp[14]) ? node12156 : 4'b1111;
															assign node12156 = (inp[4]) ? node12158 : 4'b1001;
																assign node12158 = (inp[9]) ? 4'b1011 : 4'b1111;
													assign node12161 = (inp[9]) ? node12165 : node12162;
														assign node12162 = (inp[4]) ? 4'b1111 : 4'b1011;
														assign node12165 = (inp[4]) ? 4'b1011 : 4'b1111;
												assign node12168 = (inp[3]) ? node12184 : node12169;
													assign node12169 = (inp[5]) ? node12177 : node12170;
														assign node12170 = (inp[4]) ? node12174 : node12171;
															assign node12171 = (inp[9]) ? 4'b1111 : 4'b1011;
															assign node12174 = (inp[9]) ? 4'b1011 : 4'b1111;
														assign node12177 = (inp[9]) ? node12181 : node12178;
															assign node12178 = (inp[4]) ? 4'b1101 : 4'b1011;
															assign node12181 = (inp[4]) ? 4'b1001 : 4'b1101;
													assign node12184 = (inp[5]) ? 4'b1101 : node12185;
														assign node12185 = (inp[4]) ? node12189 : node12186;
															assign node12186 = (inp[9]) ? 4'b1101 : 4'b1011;
															assign node12189 = (inp[9]) ? 4'b1001 : 4'b1101;
								assign node12193 = (inp[14]) ? node12465 : node12194;
									assign node12194 = (inp[2]) ? node12336 : node12195;
										assign node12195 = (inp[12]) ? node12271 : node12196;
											assign node12196 = (inp[0]) ? node12238 : node12197;
												assign node12197 = (inp[15]) ? node12209 : node12198;
													assign node12198 = (inp[5]) ? node12206 : node12199;
														assign node12199 = (inp[9]) ? node12203 : node12200;
															assign node12200 = (inp[4]) ? 4'b1011 : 4'b1111;
															assign node12203 = (inp[4]) ? 4'b1111 : 4'b1011;
														assign node12206 = (inp[3]) ? 4'b1101 : 4'b1011;
													assign node12209 = (inp[3]) ? node12225 : node12210;
														assign node12210 = (inp[5]) ? node12218 : node12211;
															assign node12211 = (inp[9]) ? node12215 : node12212;
																assign node12212 = (inp[4]) ? 4'b1001 : 4'b1101;
																assign node12215 = (inp[4]) ? 4'b1101 : 4'b1001;
															assign node12218 = (inp[9]) ? node12222 : node12219;
																assign node12219 = (inp[4]) ? 4'b1001 : 4'b1101;
																assign node12222 = (inp[4]) ? 4'b1111 : 4'b1001;
														assign node12225 = (inp[5]) ? node12231 : node12226;
															assign node12226 = (inp[4]) ? node12228 : 4'b1001;
																assign node12228 = (inp[9]) ? 4'b1111 : 4'b1001;
															assign node12231 = (inp[9]) ? node12235 : node12232;
																assign node12232 = (inp[4]) ? 4'b1011 : 4'b1111;
																assign node12235 = (inp[4]) ? 4'b1111 : 4'b1011;
												assign node12238 = (inp[15]) ? node12254 : node12239;
													assign node12239 = (inp[3]) ? node12247 : node12240;
														assign node12240 = (inp[4]) ? node12244 : node12241;
															assign node12241 = (inp[9]) ? 4'b1001 : 4'b1101;
															assign node12244 = (inp[9]) ? 4'b1101 : 4'b1001;
														assign node12247 = (inp[5]) ? 4'b1011 : node12248;
															assign node12248 = (inp[4]) ? 4'b1001 : node12249;
																assign node12249 = (inp[9]) ? 4'b1001 : 4'b1101;
													assign node12254 = (inp[3]) ? node12264 : node12255;
														assign node12255 = (inp[4]) ? node12259 : node12256;
															assign node12256 = (inp[9]) ? 4'b1011 : 4'b1111;
															assign node12259 = (inp[9]) ? node12261 : 4'b1011;
																assign node12261 = (inp[5]) ? 4'b1101 : 4'b1111;
														assign node12264 = (inp[9]) ? 4'b1101 : node12265;
															assign node12265 = (inp[5]) ? 4'b1101 : node12266;
																assign node12266 = (inp[4]) ? 4'b1011 : 4'b1111;
											assign node12271 = (inp[3]) ? node12307 : node12272;
												assign node12272 = (inp[5]) ? node12294 : node12273;
													assign node12273 = (inp[4]) ? node12283 : node12274;
														assign node12274 = (inp[9]) ? node12276 : 4'b1001;
															assign node12276 = (inp[0]) ? node12280 : node12277;
																assign node12277 = (inp[15]) ? 4'b1101 : 4'b1111;
																assign node12280 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node12283 = (inp[9]) ? node12289 : node12284;
															assign node12284 = (inp[0]) ? 4'b1111 : node12285;
																assign node12285 = (inp[15]) ? 4'b1101 : 4'b1111;
															assign node12289 = (inp[15]) ? 4'b1011 : node12290;
																assign node12290 = (inp[0]) ? 4'b1001 : 4'b1011;
													assign node12294 = (inp[4]) ? node12302 : node12295;
														assign node12295 = (inp[9]) ? 4'b1111 : node12296;
															assign node12296 = (inp[0]) ? 4'b1011 : node12297;
																assign node12297 = (inp[15]) ? 4'b1001 : 4'b1011;
														assign node12302 = (inp[9]) ? node12304 : 4'b1101;
															assign node12304 = (inp[0]) ? 4'b1001 : 4'b1011;
												assign node12307 = (inp[9]) ? node12323 : node12308;
													assign node12308 = (inp[4]) ? node12318 : node12309;
														assign node12309 = (inp[0]) ? 4'b1011 : node12310;
															assign node12310 = (inp[5]) ? node12314 : node12311;
																assign node12311 = (inp[15]) ? 4'b1001 : 4'b1011;
																assign node12314 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node12318 = (inp[5]) ? node12320 : 4'b1111;
															assign node12320 = (inp[15]) ? 4'b1111 : 4'b1101;
													assign node12323 = (inp[4]) ? node12329 : node12324;
														assign node12324 = (inp[5]) ? node12326 : 4'b1101;
															assign node12326 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node12329 = (inp[0]) ? node12333 : node12330;
															assign node12330 = (inp[15]) ? 4'b1011 : 4'b1001;
															assign node12333 = (inp[15]) ? 4'b1001 : 4'b1011;
										assign node12336 = (inp[15]) ? node12398 : node12337;
											assign node12337 = (inp[0]) ? node12375 : node12338;
												assign node12338 = (inp[3]) ? node12356 : node12339;
													assign node12339 = (inp[5]) ? node12349 : node12340;
														assign node12340 = (inp[4]) ? node12342 : 4'b1010;
															assign node12342 = (inp[12]) ? node12346 : node12343;
																assign node12343 = (inp[9]) ? 4'b1110 : 4'b1010;
																assign node12346 = (inp[9]) ? 4'b1010 : 4'b1110;
														assign node12349 = (inp[9]) ? node12353 : node12350;
															assign node12350 = (inp[12]) ? 4'b1010 : 4'b1110;
															assign node12353 = (inp[12]) ? 4'b1100 : 4'b1010;
													assign node12356 = (inp[4]) ? node12368 : node12357;
														assign node12357 = (inp[5]) ? node12363 : node12358;
															assign node12358 = (inp[12]) ? 4'b1010 : node12359;
																assign node12359 = (inp[9]) ? 4'b1010 : 4'b1110;
															assign node12363 = (inp[9]) ? node12365 : 4'b1000;
																assign node12365 = (inp[12]) ? 4'b1100 : 4'b1000;
														assign node12368 = (inp[5]) ? node12370 : 4'b1100;
															assign node12370 = (inp[12]) ? node12372 : 4'b1100;
																assign node12372 = (inp[9]) ? 4'b1000 : 4'b1100;
												assign node12375 = (inp[3]) ? node12385 : node12376;
													assign node12376 = (inp[4]) ? 4'b1000 : node12377;
														assign node12377 = (inp[9]) ? node12381 : node12378;
															assign node12378 = (inp[12]) ? 4'b1000 : 4'b1100;
															assign node12381 = (inp[12]) ? 4'b1100 : 4'b1000;
													assign node12385 = (inp[5]) ? node12391 : node12386;
														assign node12386 = (inp[9]) ? node12388 : 4'b1000;
															assign node12388 = (inp[12]) ? 4'b1110 : 4'b1000;
														assign node12391 = (inp[4]) ? 4'b1010 : node12392;
															assign node12392 = (inp[9]) ? node12394 : 4'b1110;
																assign node12394 = (inp[12]) ? 4'b1110 : 4'b1010;
											assign node12398 = (inp[0]) ? node12442 : node12399;
												assign node12399 = (inp[5]) ? node12417 : node12400;
													assign node12400 = (inp[4]) ? node12412 : node12401;
														assign node12401 = (inp[3]) ? node12407 : node12402;
															assign node12402 = (inp[9]) ? node12404 : 4'b1000;
																assign node12404 = (inp[12]) ? 4'b1100 : 4'b1000;
															assign node12407 = (inp[9]) ? 4'b1110 : node12408;
																assign node12408 = (inp[12]) ? 4'b1000 : 4'b1100;
														assign node12412 = (inp[9]) ? node12414 : 4'b1000;
															assign node12414 = (inp[3]) ? 4'b1010 : 4'b1000;
													assign node12417 = (inp[3]) ? node12431 : node12418;
														assign node12418 = (inp[12]) ? node12424 : node12419;
															assign node12419 = (inp[9]) ? 4'b1000 : node12420;
																assign node12420 = (inp[4]) ? 4'b1000 : 4'b1100;
															assign node12424 = (inp[4]) ? node12428 : node12425;
																assign node12425 = (inp[9]) ? 4'b1110 : 4'b1000;
																assign node12428 = (inp[9]) ? 4'b1010 : 4'b1110;
														assign node12431 = (inp[12]) ? node12437 : node12432;
															assign node12432 = (inp[4]) ? node12434 : 4'b1110;
																assign node12434 = (inp[9]) ? 4'b1110 : 4'b1010;
															assign node12437 = (inp[4]) ? node12439 : 4'b1010;
																assign node12439 = (inp[9]) ? 4'b1010 : 4'b1110;
												assign node12442 = (inp[3]) ? node12448 : node12443;
													assign node12443 = (inp[9]) ? node12445 : 4'b1110;
														assign node12445 = (inp[4]) ? 4'b1110 : 4'b1010;
													assign node12448 = (inp[4]) ? node12456 : node12449;
														assign node12449 = (inp[5]) ? 4'b1000 : node12450;
															assign node12450 = (inp[9]) ? 4'b1010 : node12451;
																assign node12451 = (inp[12]) ? 4'b1010 : 4'b1110;
														assign node12456 = (inp[5]) ? 4'b1100 : node12457;
															assign node12457 = (inp[9]) ? node12461 : node12458;
																assign node12458 = (inp[12]) ? 4'b1100 : 4'b1010;
																assign node12461 = (inp[12]) ? 4'b1000 : 4'b1100;
									assign node12465 = (inp[5]) ? node12583 : node12466;
										assign node12466 = (inp[12]) ? node12526 : node12467;
											assign node12467 = (inp[3]) ? node12487 : node12468;
												assign node12468 = (inp[0]) ? node12478 : node12469;
													assign node12469 = (inp[15]) ? 4'b1000 : node12470;
														assign node12470 = (inp[9]) ? node12474 : node12471;
															assign node12471 = (inp[4]) ? 4'b1010 : 4'b1110;
															assign node12474 = (inp[4]) ? 4'b1110 : 4'b1010;
													assign node12478 = (inp[15]) ? node12484 : node12479;
														assign node12479 = (inp[4]) ? 4'b1000 : node12480;
															assign node12480 = (inp[2]) ? 4'b1000 : 4'b1100;
														assign node12484 = (inp[4]) ? 4'b1110 : 4'b1010;
												assign node12487 = (inp[4]) ? node12511 : node12488;
													assign node12488 = (inp[9]) ? node12502 : node12489;
														assign node12489 = (inp[2]) ? node12495 : node12490;
															assign node12490 = (inp[15]) ? node12492 : 4'b1110;
																assign node12492 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node12495 = (inp[15]) ? node12499 : node12496;
																assign node12496 = (inp[0]) ? 4'b1100 : 4'b1110;
																assign node12499 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node12502 = (inp[2]) ? node12506 : node12503;
															assign node12503 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node12506 = (inp[15]) ? node12508 : 4'b1000;
																assign node12508 = (inp[0]) ? 4'b1010 : 4'b1000;
													assign node12511 = (inp[9]) ? node12519 : node12512;
														assign node12512 = (inp[0]) ? node12516 : node12513;
															assign node12513 = (inp[15]) ? 4'b1000 : 4'b1010;
															assign node12516 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node12519 = (inp[2]) ? 4'b1110 : node12520;
															assign node12520 = (inp[0]) ? node12522 : 4'b1100;
																assign node12522 = (inp[15]) ? 4'b1100 : 4'b1110;
											assign node12526 = (inp[9]) ? node12548 : node12527;
												assign node12527 = (inp[4]) ? node12539 : node12528;
													assign node12528 = (inp[3]) ? node12534 : node12529;
														assign node12529 = (inp[0]) ? node12531 : 4'b1010;
															assign node12531 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node12534 = (inp[0]) ? node12536 : 4'b1000;
															assign node12536 = (inp[15]) ? 4'b1010 : 4'b1000;
													assign node12539 = (inp[0]) ? node12541 : 4'b1100;
														assign node12541 = (inp[3]) ? node12545 : node12542;
															assign node12542 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node12545 = (inp[15]) ? 4'b1100 : 4'b1110;
												assign node12548 = (inp[4]) ? node12566 : node12549;
													assign node12549 = (inp[2]) ? node12559 : node12550;
														assign node12550 = (inp[15]) ? node12552 : 4'b1100;
															assign node12552 = (inp[3]) ? node12556 : node12553;
																assign node12553 = (inp[0]) ? 4'b1110 : 4'b1100;
																assign node12556 = (inp[0]) ? 4'b1100 : 4'b1110;
														assign node12559 = (inp[3]) ? 4'b1110 : node12560;
															assign node12560 = (inp[15]) ? node12562 : 4'b1110;
																assign node12562 = (inp[0]) ? 4'b1110 : 4'b1100;
													assign node12566 = (inp[2]) ? node12576 : node12567;
														assign node12567 = (inp[3]) ? node12569 : 4'b1010;
															assign node12569 = (inp[15]) ? node12573 : node12570;
																assign node12570 = (inp[0]) ? 4'b1010 : 4'b1000;
																assign node12573 = (inp[0]) ? 4'b1000 : 4'b1010;
														assign node12576 = (inp[3]) ? node12578 : 4'b1000;
															assign node12578 = (inp[0]) ? node12580 : 4'b1010;
																assign node12580 = (inp[15]) ? 4'b1000 : 4'b1010;
										assign node12583 = (inp[0]) ? node12661 : node12584;
											assign node12584 = (inp[15]) ? node12620 : node12585;
												assign node12585 = (inp[3]) ? node12597 : node12586;
													assign node12586 = (inp[4]) ? node12594 : node12587;
														assign node12587 = (inp[9]) ? node12591 : node12588;
															assign node12588 = (inp[12]) ? 4'b1010 : 4'b1110;
															assign node12591 = (inp[12]) ? 4'b1100 : 4'b1010;
														assign node12594 = (inp[12]) ? 4'b1000 : 4'b1100;
													assign node12597 = (inp[12]) ? node12611 : node12598;
														assign node12598 = (inp[2]) ? node12606 : node12599;
															assign node12599 = (inp[9]) ? node12603 : node12600;
																assign node12600 = (inp[4]) ? 4'b1000 : 4'b1100;
																assign node12603 = (inp[4]) ? 4'b1100 : 4'b1000;
															assign node12606 = (inp[9]) ? node12608 : 4'b1000;
																assign node12608 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node12611 = (inp[2]) ? 4'b1100 : node12612;
															assign node12612 = (inp[4]) ? node12616 : node12613;
																assign node12613 = (inp[9]) ? 4'b1100 : 4'b1000;
																assign node12616 = (inp[9]) ? 4'b1000 : 4'b1100;
												assign node12620 = (inp[3]) ? node12640 : node12621;
													assign node12621 = (inp[4]) ? node12629 : node12622;
														assign node12622 = (inp[9]) ? node12626 : node12623;
															assign node12623 = (inp[12]) ? 4'b1000 : 4'b1100;
															assign node12626 = (inp[12]) ? 4'b1110 : 4'b1000;
														assign node12629 = (inp[2]) ? node12635 : node12630;
															assign node12630 = (inp[9]) ? node12632 : 4'b1110;
																assign node12632 = (inp[12]) ? 4'b1010 : 4'b1110;
															assign node12635 = (inp[9]) ? node12637 : 4'b1000;
																assign node12637 = (inp[12]) ? 4'b1010 : 4'b1110;
													assign node12640 = (inp[4]) ? node12650 : node12641;
														assign node12641 = (inp[2]) ? node12643 : 4'b1110;
															assign node12643 = (inp[9]) ? node12647 : node12644;
																assign node12644 = (inp[12]) ? 4'b1010 : 4'b1110;
																assign node12647 = (inp[12]) ? 4'b1110 : 4'b1010;
														assign node12650 = (inp[2]) ? node12656 : node12651;
															assign node12651 = (inp[12]) ? node12653 : 4'b1010;
																assign node12653 = (inp[9]) ? 4'b1010 : 4'b1110;
															assign node12656 = (inp[12]) ? node12658 : 4'b1110;
																assign node12658 = (inp[9]) ? 4'b1010 : 4'b1110;
											assign node12661 = (inp[15]) ? node12675 : node12662;
												assign node12662 = (inp[3]) ? node12668 : node12663;
													assign node12663 = (inp[4]) ? node12665 : 4'b1000;
														assign node12665 = (inp[9]) ? 4'b1110 : 4'b1000;
													assign node12668 = (inp[4]) ? 4'b1110 : node12669;
														assign node12669 = (inp[2]) ? node12671 : 4'b1010;
															assign node12671 = (inp[12]) ? 4'b1010 : 4'b1110;
												assign node12675 = (inp[3]) ? node12695 : node12676;
													assign node12676 = (inp[12]) ? node12688 : node12677;
														assign node12677 = (inp[2]) ? node12683 : node12678;
															assign node12678 = (inp[9]) ? 4'b1100 : node12679;
																assign node12679 = (inp[4]) ? 4'b1010 : 4'b1110;
															assign node12683 = (inp[4]) ? 4'b1010 : node12684;
																assign node12684 = (inp[9]) ? 4'b1010 : 4'b1110;
														assign node12688 = (inp[9]) ? node12692 : node12689;
															assign node12689 = (inp[4]) ? 4'b1100 : 4'b1010;
															assign node12692 = (inp[4]) ? 4'b1000 : 4'b1100;
													assign node12695 = (inp[9]) ? node12703 : node12696;
														assign node12696 = (inp[12]) ? node12700 : node12697;
															assign node12697 = (inp[4]) ? 4'b1000 : 4'b1100;
															assign node12700 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node12703 = (inp[12]) ? node12707 : node12704;
															assign node12704 = (inp[4]) ? 4'b1100 : 4'b1000;
															assign node12707 = (inp[4]) ? 4'b1000 : 4'b1100;
						assign node12710 = (inp[14]) ? node13968 : node12711;
							assign node12711 = (inp[8]) ? node13343 : node12712;
								assign node12712 = (inp[5]) ? node13022 : node12713;
									assign node12713 = (inp[3]) ? node12875 : node12714;
										assign node12714 = (inp[2]) ? node12800 : node12715;
											assign node12715 = (inp[7]) ? node12751 : node12716;
												assign node12716 = (inp[15]) ? node12734 : node12717;
													assign node12717 = (inp[0]) ? node12727 : node12718;
														assign node12718 = (inp[4]) ? node12720 : 4'b1111;
															assign node12720 = (inp[9]) ? node12724 : node12721;
																assign node12721 = (inp[12]) ? 4'b1111 : 4'b1011;
																assign node12724 = (inp[12]) ? 4'b1011 : 4'b1111;
														assign node12727 = (inp[9]) ? node12731 : node12728;
															assign node12728 = (inp[12]) ? 4'b1001 : 4'b1101;
															assign node12731 = (inp[12]) ? 4'b1101 : 4'b1001;
													assign node12734 = (inp[0]) ? node12748 : node12735;
														assign node12735 = (inp[12]) ? node12743 : node12736;
															assign node12736 = (inp[4]) ? node12740 : node12737;
																assign node12737 = (inp[9]) ? 4'b1001 : 4'b1101;
																assign node12740 = (inp[9]) ? 4'b1101 : 4'b1001;
															assign node12743 = (inp[4]) ? node12745 : 4'b1001;
																assign node12745 = (inp[9]) ? 4'b1001 : 4'b1101;
														assign node12748 = (inp[9]) ? 4'b1111 : 4'b1011;
												assign node12751 = (inp[9]) ? node12773 : node12752;
													assign node12752 = (inp[0]) ? node12760 : node12753;
														assign node12753 = (inp[15]) ? node12755 : 4'b1010;
															assign node12755 = (inp[4]) ? 4'b1000 : node12756;
																assign node12756 = (inp[12]) ? 4'b1000 : 4'b1100;
														assign node12760 = (inp[15]) ? node12768 : node12761;
															assign node12761 = (inp[4]) ? node12765 : node12762;
																assign node12762 = (inp[12]) ? 4'b1000 : 4'b1100;
																assign node12765 = (inp[12]) ? 4'b1100 : 4'b1000;
															assign node12768 = (inp[12]) ? node12770 : 4'b1110;
																assign node12770 = (inp[4]) ? 4'b1110 : 4'b1010;
													assign node12773 = (inp[4]) ? node12785 : node12774;
														assign node12774 = (inp[12]) ? node12780 : node12775;
															assign node12775 = (inp[15]) ? node12777 : 4'b1010;
																assign node12777 = (inp[0]) ? 4'b1010 : 4'b1000;
															assign node12780 = (inp[0]) ? 4'b1110 : node12781;
																assign node12781 = (inp[15]) ? 4'b1100 : 4'b1110;
														assign node12785 = (inp[12]) ? node12793 : node12786;
															assign node12786 = (inp[0]) ? node12790 : node12787;
																assign node12787 = (inp[15]) ? 4'b1100 : 4'b1110;
																assign node12790 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node12793 = (inp[0]) ? node12797 : node12794;
																assign node12794 = (inp[15]) ? 4'b1000 : 4'b1010;
																assign node12797 = (inp[15]) ? 4'b1010 : 4'b1000;
											assign node12800 = (inp[7]) ? node12832 : node12801;
												assign node12801 = (inp[9]) ? node12817 : node12802;
													assign node12802 = (inp[0]) ? node12806 : node12803;
														assign node12803 = (inp[15]) ? 4'b1100 : 4'b1110;
														assign node12806 = (inp[15]) ? node12810 : node12807;
															assign node12807 = (inp[4]) ? 4'b1000 : 4'b1100;
															assign node12810 = (inp[12]) ? node12814 : node12811;
																assign node12811 = (inp[4]) ? 4'b1010 : 4'b1110;
																assign node12814 = (inp[4]) ? 4'b1110 : 4'b1010;
													assign node12817 = (inp[15]) ? node12825 : node12818;
														assign node12818 = (inp[0]) ? node12820 : 4'b1110;
															assign node12820 = (inp[12]) ? node12822 : 4'b1100;
																assign node12822 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node12825 = (inp[0]) ? 4'b1010 : node12826;
															assign node12826 = (inp[4]) ? node12828 : 4'b1000;
																assign node12828 = (inp[12]) ? 4'b1000 : 4'b1100;
												assign node12832 = (inp[4]) ? node12860 : node12833;
													assign node12833 = (inp[0]) ? node12845 : node12834;
														assign node12834 = (inp[15]) ? node12838 : node12835;
															assign node12835 = (inp[9]) ? 4'b1011 : 4'b1111;
															assign node12838 = (inp[12]) ? node12842 : node12839;
																assign node12839 = (inp[9]) ? 4'b1001 : 4'b1101;
																assign node12842 = (inp[9]) ? 4'b1101 : 4'b1001;
														assign node12845 = (inp[15]) ? node12853 : node12846;
															assign node12846 = (inp[9]) ? node12850 : node12847;
																assign node12847 = (inp[12]) ? 4'b1001 : 4'b1101;
																assign node12850 = (inp[12]) ? 4'b1101 : 4'b1001;
															assign node12853 = (inp[12]) ? node12857 : node12854;
																assign node12854 = (inp[9]) ? 4'b1011 : 4'b1111;
																assign node12857 = (inp[9]) ? 4'b1111 : 4'b1011;
													assign node12860 = (inp[0]) ? node12868 : node12861;
														assign node12861 = (inp[15]) ? 4'b1101 : node12862;
															assign node12862 = (inp[9]) ? 4'b1111 : node12863;
																assign node12863 = (inp[12]) ? 4'b1111 : 4'b1011;
														assign node12868 = (inp[15]) ? node12870 : 4'b1101;
															assign node12870 = (inp[9]) ? 4'b1011 : node12871;
																assign node12871 = (inp[12]) ? 4'b1111 : 4'b1011;
										assign node12875 = (inp[2]) ? node12941 : node12876;
											assign node12876 = (inp[7]) ? node12916 : node12877;
												assign node12877 = (inp[15]) ? node12895 : node12878;
													assign node12878 = (inp[4]) ? node12890 : node12879;
														assign node12879 = (inp[0]) ? node12887 : node12880;
															assign node12880 = (inp[12]) ? node12884 : node12881;
																assign node12881 = (inp[9]) ? 4'b1011 : 4'b1111;
																assign node12884 = (inp[9]) ? 4'b1101 : 4'b1011;
															assign node12887 = (inp[9]) ? 4'b1111 : 4'b1101;
														assign node12890 = (inp[12]) ? 4'b1011 : node12891;
															assign node12891 = (inp[0]) ? 4'b1111 : 4'b1011;
													assign node12895 = (inp[9]) ? node12903 : node12896;
														assign node12896 = (inp[0]) ? node12900 : node12897;
															assign node12897 = (inp[12]) ? 4'b1111 : 4'b1001;
															assign node12900 = (inp[12]) ? 4'b1011 : 4'b1111;
														assign node12903 = (inp[0]) ? node12909 : node12904;
															assign node12904 = (inp[12]) ? 4'b1111 : node12905;
																assign node12905 = (inp[4]) ? 4'b1111 : 4'b1001;
															assign node12909 = (inp[12]) ? node12913 : node12910;
																assign node12910 = (inp[4]) ? 4'b1101 : 4'b1011;
																assign node12913 = (inp[4]) ? 4'b1001 : 4'b1101;
												assign node12916 = (inp[15]) ? node12928 : node12917;
													assign node12917 = (inp[9]) ? node12923 : node12918;
														assign node12918 = (inp[12]) ? node12920 : 4'b1100;
															assign node12920 = (inp[0]) ? 4'b1000 : 4'b1010;
														assign node12923 = (inp[12]) ? 4'b1010 : node12924;
															assign node12924 = (inp[0]) ? 4'b1110 : 4'b1010;
													assign node12928 = (inp[9]) ? node12938 : node12929;
														assign node12929 = (inp[0]) ? node12933 : node12930;
															assign node12930 = (inp[12]) ? 4'b1110 : 4'b1100;
															assign node12933 = (inp[4]) ? 4'b1010 : node12934;
																assign node12934 = (inp[12]) ? 4'b1010 : 4'b1110;
														assign node12938 = (inp[0]) ? 4'b1100 : 4'b1110;
											assign node12941 = (inp[7]) ? node12979 : node12942;
												assign node12942 = (inp[4]) ? node12960 : node12943;
													assign node12943 = (inp[12]) ? node12949 : node12944;
														assign node12944 = (inp[0]) ? 4'b1110 : node12945;
															assign node12945 = (inp[15]) ? 4'b1100 : 4'b1110;
														assign node12949 = (inp[9]) ? node12955 : node12950;
															assign node12950 = (inp[15]) ? node12952 : 4'b1010;
																assign node12952 = (inp[0]) ? 4'b1010 : 4'b1000;
															assign node12955 = (inp[15]) ? 4'b1110 : node12956;
																assign node12956 = (inp[0]) ? 4'b1110 : 4'b1100;
													assign node12960 = (inp[9]) ? node12968 : node12961;
														assign node12961 = (inp[12]) ? 4'b1100 : node12962;
															assign node12962 = (inp[0]) ? node12964 : 4'b1000;
																assign node12964 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node12968 = (inp[12]) ? node12974 : node12969;
															assign node12969 = (inp[0]) ? node12971 : 4'b1110;
																assign node12971 = (inp[15]) ? 4'b1100 : 4'b1110;
															assign node12974 = (inp[0]) ? 4'b1000 : node12975;
																assign node12975 = (inp[15]) ? 4'b1010 : 4'b1000;
												assign node12979 = (inp[4]) ? node13001 : node12980;
													assign node12980 = (inp[12]) ? node12990 : node12981;
														assign node12981 = (inp[9]) ? 4'b1001 : node12982;
															assign node12982 = (inp[0]) ? node12986 : node12983;
																assign node12983 = (inp[15]) ? 4'b1101 : 4'b1111;
																assign node12986 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node12990 = (inp[9]) ? node12996 : node12991;
															assign node12991 = (inp[15]) ? node12993 : 4'b1001;
																assign node12993 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node12996 = (inp[0]) ? 4'b1101 : node12997;
																assign node12997 = (inp[15]) ? 4'b1111 : 4'b1101;
													assign node13001 = (inp[12]) ? node13011 : node13002;
														assign node13002 = (inp[9]) ? node13008 : node13003;
															assign node13003 = (inp[15]) ? 4'b1001 : node13004;
																assign node13004 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node13008 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node13011 = (inp[9]) ? node13017 : node13012;
															assign node13012 = (inp[0]) ? node13014 : 4'b1111;
																assign node13014 = (inp[15]) ? 4'b1101 : 4'b1111;
															assign node13017 = (inp[15]) ? node13019 : 4'b1011;
																assign node13019 = (inp[0]) ? 4'b1001 : 4'b1011;
									assign node13022 = (inp[9]) ? node13198 : node13023;
										assign node13023 = (inp[0]) ? node13107 : node13024;
											assign node13024 = (inp[15]) ? node13068 : node13025;
												assign node13025 = (inp[3]) ? node13041 : node13026;
													assign node13026 = (inp[4]) ? node13036 : node13027;
														assign node13027 = (inp[12]) ? node13029 : 4'b1110;
															assign node13029 = (inp[2]) ? node13033 : node13030;
																assign node13030 = (inp[7]) ? 4'b1010 : 4'b1011;
																assign node13033 = (inp[7]) ? 4'b1011 : 4'b1010;
														assign node13036 = (inp[12]) ? node13038 : 4'b1011;
															assign node13038 = (inp[2]) ? 4'b1101 : 4'b1100;
													assign node13041 = (inp[12]) ? node13053 : node13042;
														assign node13042 = (inp[4]) ? node13048 : node13043;
															assign node13043 = (inp[2]) ? node13045 : 4'b1100;
																assign node13045 = (inp[7]) ? 4'b1101 : 4'b1100;
															assign node13048 = (inp[2]) ? 4'b1000 : node13049;
																assign node13049 = (inp[7]) ? 4'b1000 : 4'b1001;
														assign node13053 = (inp[4]) ? node13061 : node13054;
															assign node13054 = (inp[7]) ? node13058 : node13055;
																assign node13055 = (inp[2]) ? 4'b1000 : 4'b1001;
																assign node13058 = (inp[2]) ? 4'b1001 : 4'b1000;
															assign node13061 = (inp[2]) ? node13065 : node13062;
																assign node13062 = (inp[7]) ? 4'b1100 : 4'b1101;
																assign node13065 = (inp[7]) ? 4'b1101 : 4'b1100;
												assign node13068 = (inp[3]) ? node13088 : node13069;
													assign node13069 = (inp[4]) ? node13081 : node13070;
														assign node13070 = (inp[12]) ? node13078 : node13071;
															assign node13071 = (inp[7]) ? node13075 : node13072;
																assign node13072 = (inp[2]) ? 4'b1100 : 4'b1101;
																assign node13075 = (inp[2]) ? 4'b1101 : 4'b1100;
															assign node13078 = (inp[2]) ? 4'b1001 : 4'b1000;
														assign node13081 = (inp[12]) ? 4'b1111 : node13082;
															assign node13082 = (inp[7]) ? node13084 : 4'b1000;
																assign node13084 = (inp[2]) ? 4'b1001 : 4'b1000;
													assign node13088 = (inp[4]) ? node13100 : node13089;
														assign node13089 = (inp[12]) ? node13093 : node13090;
															assign node13090 = (inp[2]) ? 4'b1111 : 4'b1110;
															assign node13093 = (inp[2]) ? node13097 : node13094;
																assign node13094 = (inp[7]) ? 4'b1010 : 4'b1011;
																assign node13097 = (inp[7]) ? 4'b1011 : 4'b1010;
														assign node13100 = (inp[12]) ? node13102 : 4'b1010;
															assign node13102 = (inp[7]) ? node13104 : 4'b1110;
																assign node13104 = (inp[2]) ? 4'b1111 : 4'b1110;
											assign node13107 = (inp[15]) ? node13155 : node13108;
												assign node13108 = (inp[3]) ? node13134 : node13109;
													assign node13109 = (inp[4]) ? node13123 : node13110;
														assign node13110 = (inp[12]) ? node13118 : node13111;
															assign node13111 = (inp[7]) ? node13115 : node13112;
																assign node13112 = (inp[2]) ? 4'b1100 : 4'b1101;
																assign node13115 = (inp[2]) ? 4'b1101 : 4'b1100;
															assign node13118 = (inp[7]) ? node13120 : 4'b1001;
																assign node13120 = (inp[2]) ? 4'b1001 : 4'b1000;
														assign node13123 = (inp[12]) ? node13129 : node13124;
															assign node13124 = (inp[2]) ? 4'b1000 : node13125;
																assign node13125 = (inp[7]) ? 4'b1000 : 4'b1001;
															assign node13129 = (inp[7]) ? node13131 : 4'b1110;
																assign node13131 = (inp[2]) ? 4'b1111 : 4'b1110;
													assign node13134 = (inp[7]) ? node13144 : node13135;
														assign node13135 = (inp[2]) ? node13139 : node13136;
															assign node13136 = (inp[4]) ? 4'b1111 : 4'b1011;
															assign node13139 = (inp[4]) ? node13141 : 4'b1110;
																assign node13141 = (inp[12]) ? 4'b1110 : 4'b1010;
														assign node13144 = (inp[2]) ? node13148 : node13145;
															assign node13145 = (inp[4]) ? 4'b1110 : 4'b1010;
															assign node13148 = (inp[4]) ? node13152 : node13149;
																assign node13149 = (inp[12]) ? 4'b1011 : 4'b1111;
																assign node13152 = (inp[12]) ? 4'b1111 : 4'b1011;
												assign node13155 = (inp[3]) ? node13179 : node13156;
													assign node13156 = (inp[12]) ? node13168 : node13157;
														assign node13157 = (inp[4]) ? node13161 : node13158;
															assign node13158 = (inp[7]) ? 4'b1110 : 4'b1111;
															assign node13161 = (inp[2]) ? node13165 : node13162;
																assign node13162 = (inp[7]) ? 4'b1010 : 4'b1011;
																assign node13165 = (inp[7]) ? 4'b1011 : 4'b1010;
														assign node13168 = (inp[4]) ? node13172 : node13169;
															assign node13169 = (inp[2]) ? 4'b1010 : 4'b1011;
															assign node13172 = (inp[7]) ? node13176 : node13173;
																assign node13173 = (inp[2]) ? 4'b1100 : 4'b1101;
																assign node13176 = (inp[2]) ? 4'b1101 : 4'b1100;
													assign node13179 = (inp[4]) ? node13191 : node13180;
														assign node13180 = (inp[12]) ? node13186 : node13181;
															assign node13181 = (inp[2]) ? node13183 : 4'b1101;
																assign node13183 = (inp[7]) ? 4'b1101 : 4'b1100;
															assign node13186 = (inp[7]) ? 4'b1000 : node13187;
																assign node13187 = (inp[2]) ? 4'b1000 : 4'b1001;
														assign node13191 = (inp[12]) ? node13193 : 4'b1001;
															assign node13193 = (inp[7]) ? node13195 : 4'b1101;
																assign node13195 = (inp[2]) ? 4'b1101 : 4'b1100;
										assign node13198 = (inp[0]) ? node13264 : node13199;
											assign node13199 = (inp[15]) ? node13231 : node13200;
												assign node13200 = (inp[2]) ? node13218 : node13201;
													assign node13201 = (inp[7]) ? node13211 : node13202;
														assign node13202 = (inp[3]) ? 4'b1001 : node13203;
															assign node13203 = (inp[4]) ? node13207 : node13204;
																assign node13204 = (inp[12]) ? 4'b1101 : 4'b1011;
																assign node13207 = (inp[12]) ? 4'b1001 : 4'b1101;
														assign node13211 = (inp[4]) ? node13215 : node13212;
															assign node13212 = (inp[12]) ? 4'b1100 : 4'b1010;
															assign node13215 = (inp[12]) ? 4'b1000 : 4'b1100;
													assign node13218 = (inp[7]) ? node13220 : 4'b1100;
														assign node13220 = (inp[3]) ? node13224 : node13221;
															assign node13221 = (inp[4]) ? 4'b1101 : 4'b1011;
															assign node13224 = (inp[4]) ? node13228 : node13225;
																assign node13225 = (inp[12]) ? 4'b1101 : 4'b1001;
																assign node13228 = (inp[12]) ? 4'b1001 : 4'b1101;
												assign node13231 = (inp[4]) ? node13251 : node13232;
													assign node13232 = (inp[12]) ? node13246 : node13233;
														assign node13233 = (inp[3]) ? node13239 : node13234;
															assign node13234 = (inp[7]) ? 4'b1000 : node13235;
																assign node13235 = (inp[2]) ? 4'b1000 : 4'b1001;
															assign node13239 = (inp[7]) ? node13243 : node13240;
																assign node13240 = (inp[2]) ? 4'b1010 : 4'b1011;
																assign node13243 = (inp[2]) ? 4'b1011 : 4'b1010;
														assign node13246 = (inp[2]) ? node13248 : 4'b1111;
															assign node13248 = (inp[7]) ? 4'b1111 : 4'b1110;
													assign node13251 = (inp[12]) ? node13259 : node13252;
														assign node13252 = (inp[2]) ? node13256 : node13253;
															assign node13253 = (inp[7]) ? 4'b1110 : 4'b1111;
															assign node13256 = (inp[7]) ? 4'b1111 : 4'b1110;
														assign node13259 = (inp[2]) ? node13261 : 4'b1011;
															assign node13261 = (inp[7]) ? 4'b1011 : 4'b1010;
											assign node13264 = (inp[15]) ? node13302 : node13265;
												assign node13265 = (inp[12]) ? node13283 : node13266;
													assign node13266 = (inp[4]) ? node13278 : node13267;
														assign node13267 = (inp[3]) ? node13275 : node13268;
															assign node13268 = (inp[2]) ? node13272 : node13269;
																assign node13269 = (inp[7]) ? 4'b1000 : 4'b1001;
																assign node13272 = (inp[7]) ? 4'b1001 : 4'b1000;
															assign node13275 = (inp[7]) ? 4'b1011 : 4'b1010;
														assign node13278 = (inp[7]) ? 4'b1110 : node13279;
															assign node13279 = (inp[2]) ? 4'b1110 : 4'b1111;
													assign node13283 = (inp[4]) ? node13297 : node13284;
														assign node13284 = (inp[3]) ? node13292 : node13285;
															assign node13285 = (inp[2]) ? node13289 : node13286;
																assign node13286 = (inp[7]) ? 4'b1110 : 4'b1111;
																assign node13289 = (inp[7]) ? 4'b1111 : 4'b1110;
															assign node13292 = (inp[2]) ? 4'b1111 : node13293;
																assign node13293 = (inp[7]) ? 4'b1110 : 4'b1111;
														assign node13297 = (inp[7]) ? 4'b1011 : node13298;
															assign node13298 = (inp[2]) ? 4'b1010 : 4'b1011;
												assign node13302 = (inp[12]) ? node13326 : node13303;
													assign node13303 = (inp[4]) ? node13317 : node13304;
														assign node13304 = (inp[3]) ? node13310 : node13305;
															assign node13305 = (inp[7]) ? node13307 : 4'b1011;
																assign node13307 = (inp[2]) ? 4'b1011 : 4'b1010;
															assign node13310 = (inp[7]) ? node13314 : node13311;
																assign node13311 = (inp[2]) ? 4'b1000 : 4'b1001;
																assign node13314 = (inp[2]) ? 4'b1001 : 4'b1000;
														assign node13317 = (inp[3]) ? node13319 : 4'b1101;
															assign node13319 = (inp[2]) ? node13323 : node13320;
																assign node13320 = (inp[7]) ? 4'b1100 : 4'b1101;
																assign node13323 = (inp[7]) ? 4'b1101 : 4'b1100;
													assign node13326 = (inp[4]) ? node13336 : node13327;
														assign node13327 = (inp[3]) ? 4'b1100 : node13328;
															assign node13328 = (inp[7]) ? node13332 : node13329;
																assign node13329 = (inp[2]) ? 4'b1100 : 4'b1101;
																assign node13332 = (inp[2]) ? 4'b1101 : 4'b1100;
														assign node13336 = (inp[7]) ? node13340 : node13337;
															assign node13337 = (inp[2]) ? 4'b1000 : 4'b1001;
															assign node13340 = (inp[2]) ? 4'b1001 : 4'b1000;
								assign node13343 = (inp[2]) ? node13659 : node13344;
									assign node13344 = (inp[7]) ? node13488 : node13345;
										assign node13345 = (inp[9]) ? node13421 : node13346;
											assign node13346 = (inp[5]) ? node13380 : node13347;
												assign node13347 = (inp[3]) ? node13361 : node13348;
													assign node13348 = (inp[12]) ? node13358 : node13349;
														assign node13349 = (inp[4]) ? node13355 : node13350;
															assign node13350 = (inp[0]) ? node13352 : 4'b1100;
																assign node13352 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node13355 = (inp[15]) ? 4'b1000 : 4'b1010;
														assign node13358 = (inp[4]) ? 4'b1110 : 4'b1010;
													assign node13361 = (inp[0]) ? node13373 : node13362;
														assign node13362 = (inp[15]) ? node13366 : node13363;
															assign node13363 = (inp[4]) ? 4'b1100 : 4'b1110;
															assign node13366 = (inp[4]) ? node13370 : node13367;
																assign node13367 = (inp[12]) ? 4'b1000 : 4'b1100;
																assign node13370 = (inp[12]) ? 4'b1110 : 4'b1000;
														assign node13373 = (inp[15]) ? 4'b1010 : node13374;
															assign node13374 = (inp[4]) ? 4'b1000 : node13375;
																assign node13375 = (inp[12]) ? 4'b1000 : 4'b1100;
												assign node13380 = (inp[15]) ? node13400 : node13381;
													assign node13381 = (inp[0]) ? node13391 : node13382;
														assign node13382 = (inp[3]) ? 4'b1000 : node13383;
															assign node13383 = (inp[12]) ? node13387 : node13384;
																assign node13384 = (inp[4]) ? 4'b1010 : 4'b1110;
																assign node13387 = (inp[4]) ? 4'b1100 : 4'b1010;
														assign node13391 = (inp[3]) ? node13393 : 4'b1000;
															assign node13393 = (inp[12]) ? node13397 : node13394;
																assign node13394 = (inp[4]) ? 4'b1010 : 4'b1110;
																assign node13397 = (inp[4]) ? 4'b1110 : 4'b1010;
													assign node13400 = (inp[0]) ? node13412 : node13401;
														assign node13401 = (inp[3]) ? node13407 : node13402;
															assign node13402 = (inp[4]) ? 4'b1000 : node13403;
																assign node13403 = (inp[12]) ? 4'b1000 : 4'b1100;
															assign node13407 = (inp[12]) ? 4'b1110 : node13408;
																assign node13408 = (inp[4]) ? 4'b1010 : 4'b1110;
														assign node13412 = (inp[4]) ? node13418 : node13413;
															assign node13413 = (inp[3]) ? 4'b1000 : node13414;
																assign node13414 = (inp[12]) ? 4'b1010 : 4'b1110;
															assign node13418 = (inp[12]) ? 4'b1100 : 4'b1000;
											assign node13421 = (inp[3]) ? node13449 : node13422;
												assign node13422 = (inp[12]) ? node13432 : node13423;
													assign node13423 = (inp[4]) ? 4'b1110 : node13424;
														assign node13424 = (inp[5]) ? 4'b1010 : node13425;
															assign node13425 = (inp[0]) ? 4'b1000 : node13426;
																assign node13426 = (inp[15]) ? 4'b1000 : 4'b1010;
													assign node13432 = (inp[4]) ? node13440 : node13433;
														assign node13433 = (inp[0]) ? node13435 : 4'b1100;
															assign node13435 = (inp[15]) ? node13437 : 4'b1110;
																assign node13437 = (inp[5]) ? 4'b1100 : 4'b1110;
														assign node13440 = (inp[15]) ? node13442 : 4'b1000;
															assign node13442 = (inp[5]) ? node13446 : node13443;
																assign node13443 = (inp[0]) ? 4'b1010 : 4'b1000;
																assign node13446 = (inp[0]) ? 4'b1000 : 4'b1010;
												assign node13449 = (inp[5]) ? node13473 : node13450;
													assign node13450 = (inp[0]) ? node13460 : node13451;
														assign node13451 = (inp[12]) ? node13457 : node13452;
															assign node13452 = (inp[4]) ? 4'b1100 : node13453;
																assign node13453 = (inp[15]) ? 4'b1000 : 4'b1010;
															assign node13457 = (inp[4]) ? 4'b1010 : 4'b1110;
														assign node13460 = (inp[15]) ? node13466 : node13461;
															assign node13461 = (inp[4]) ? node13463 : 4'b1000;
																assign node13463 = (inp[12]) ? 4'b1010 : 4'b1110;
															assign node13466 = (inp[4]) ? node13470 : node13467;
																assign node13467 = (inp[12]) ? 4'b1100 : 4'b1010;
																assign node13470 = (inp[12]) ? 4'b1000 : 4'b1100;
													assign node13473 = (inp[0]) ? node13485 : node13474;
														assign node13474 = (inp[15]) ? node13478 : node13475;
															assign node13475 = (inp[12]) ? 4'b1100 : 4'b1000;
															assign node13478 = (inp[12]) ? node13482 : node13479;
																assign node13479 = (inp[4]) ? 4'b1110 : 4'b1010;
																assign node13482 = (inp[4]) ? 4'b1010 : 4'b1110;
														assign node13485 = (inp[15]) ? 4'b1100 : 4'b1110;
										assign node13488 = (inp[3]) ? node13572 : node13489;
											assign node13489 = (inp[15]) ? node13529 : node13490;
												assign node13490 = (inp[0]) ? node13512 : node13491;
													assign node13491 = (inp[5]) ? node13499 : node13492;
														assign node13492 = (inp[9]) ? 4'b1111 : node13493;
															assign node13493 = (inp[4]) ? 4'b1011 : node13494;
																assign node13494 = (inp[12]) ? 4'b1011 : 4'b1111;
														assign node13499 = (inp[4]) ? node13507 : node13500;
															assign node13500 = (inp[12]) ? node13504 : node13501;
																assign node13501 = (inp[9]) ? 4'b1011 : 4'b1111;
																assign node13504 = (inp[9]) ? 4'b1101 : 4'b1011;
															assign node13507 = (inp[12]) ? node13509 : 4'b1101;
																assign node13509 = (inp[9]) ? 4'b1001 : 4'b1101;
													assign node13512 = (inp[9]) ? node13520 : node13513;
														assign node13513 = (inp[5]) ? 4'b1001 : node13514;
															assign node13514 = (inp[4]) ? 4'b1001 : node13515;
																assign node13515 = (inp[12]) ? 4'b1001 : 4'b1101;
														assign node13520 = (inp[5]) ? node13524 : node13521;
															assign node13521 = (inp[4]) ? 4'b1001 : 4'b1101;
															assign node13524 = (inp[4]) ? 4'b1111 : node13525;
																assign node13525 = (inp[12]) ? 4'b1111 : 4'b1001;
												assign node13529 = (inp[0]) ? node13551 : node13530;
													assign node13530 = (inp[5]) ? node13538 : node13531;
														assign node13531 = (inp[12]) ? 4'b1001 : node13532;
															assign node13532 = (inp[9]) ? node13534 : 4'b1101;
																assign node13534 = (inp[4]) ? 4'b1101 : 4'b1001;
														assign node13538 = (inp[4]) ? node13546 : node13539;
															assign node13539 = (inp[12]) ? node13543 : node13540;
																assign node13540 = (inp[9]) ? 4'b1001 : 4'b1101;
																assign node13543 = (inp[9]) ? 4'b1111 : 4'b1001;
															assign node13546 = (inp[9]) ? node13548 : 4'b1111;
																assign node13548 = (inp[12]) ? 4'b1011 : 4'b1111;
													assign node13551 = (inp[5]) ? node13561 : node13552;
														assign node13552 = (inp[4]) ? node13554 : 4'b1111;
															assign node13554 = (inp[9]) ? node13558 : node13555;
																assign node13555 = (inp[12]) ? 4'b1111 : 4'b1011;
																assign node13558 = (inp[12]) ? 4'b1011 : 4'b1111;
														assign node13561 = (inp[4]) ? node13567 : node13562;
															assign node13562 = (inp[9]) ? 4'b1011 : node13563;
																assign node13563 = (inp[12]) ? 4'b1011 : 4'b1111;
															assign node13567 = (inp[9]) ? node13569 : 4'b1011;
																assign node13569 = (inp[12]) ? 4'b1001 : 4'b1101;
											assign node13572 = (inp[15]) ? node13624 : node13573;
												assign node13573 = (inp[0]) ? node13599 : node13574;
													assign node13574 = (inp[5]) ? node13584 : node13575;
														assign node13575 = (inp[12]) ? node13577 : 4'b1011;
															assign node13577 = (inp[4]) ? node13581 : node13578;
																assign node13578 = (inp[9]) ? 4'b1101 : 4'b1011;
																assign node13581 = (inp[9]) ? 4'b1001 : 4'b1101;
														assign node13584 = (inp[4]) ? node13592 : node13585;
															assign node13585 = (inp[9]) ? node13589 : node13586;
																assign node13586 = (inp[12]) ? 4'b1001 : 4'b1101;
																assign node13589 = (inp[12]) ? 4'b1101 : 4'b1001;
															assign node13592 = (inp[9]) ? node13596 : node13593;
																assign node13593 = (inp[12]) ? 4'b1101 : 4'b1001;
																assign node13596 = (inp[12]) ? 4'b1001 : 4'b1101;
													assign node13599 = (inp[5]) ? node13611 : node13600;
														assign node13600 = (inp[9]) ? node13604 : node13601;
															assign node13601 = (inp[12]) ? 4'b1001 : 4'b1101;
															assign node13604 = (inp[4]) ? node13608 : node13605;
																assign node13605 = (inp[12]) ? 4'b1111 : 4'b1001;
																assign node13608 = (inp[12]) ? 4'b1011 : 4'b1111;
														assign node13611 = (inp[4]) ? node13617 : node13612;
															assign node13612 = (inp[9]) ? node13614 : 4'b1011;
																assign node13614 = (inp[12]) ? 4'b1111 : 4'b1011;
															assign node13617 = (inp[12]) ? node13621 : node13618;
																assign node13618 = (inp[9]) ? 4'b1111 : 4'b1011;
																assign node13621 = (inp[9]) ? 4'b1011 : 4'b1111;
												assign node13624 = (inp[0]) ? node13640 : node13625;
													assign node13625 = (inp[5]) ? node13637 : node13626;
														assign node13626 = (inp[4]) ? node13632 : node13627;
															assign node13627 = (inp[9]) ? 4'b1001 : node13628;
																assign node13628 = (inp[12]) ? 4'b1001 : 4'b1101;
															assign node13632 = (inp[9]) ? 4'b1111 : node13633;
																assign node13633 = (inp[12]) ? 4'b1111 : 4'b1001;
														assign node13637 = (inp[12]) ? 4'b1011 : 4'b1111;
													assign node13640 = (inp[9]) ? node13654 : node13641;
														assign node13641 = (inp[5]) ? node13647 : node13642;
															assign node13642 = (inp[4]) ? node13644 : 4'b1011;
																assign node13644 = (inp[12]) ? 4'b1101 : 4'b1011;
															assign node13647 = (inp[12]) ? node13651 : node13648;
																assign node13648 = (inp[4]) ? 4'b1001 : 4'b1101;
																assign node13651 = (inp[4]) ? 4'b1101 : 4'b1001;
														assign node13654 = (inp[12]) ? node13656 : 4'b1101;
															assign node13656 = (inp[4]) ? 4'b1001 : 4'b1101;
									assign node13659 = (inp[7]) ? node13807 : node13660;
										assign node13660 = (inp[9]) ? node13740 : node13661;
											assign node13661 = (inp[5]) ? node13697 : node13662;
												assign node13662 = (inp[0]) ? node13684 : node13663;
													assign node13663 = (inp[15]) ? node13677 : node13664;
														assign node13664 = (inp[3]) ? node13672 : node13665;
															assign node13665 = (inp[4]) ? node13669 : node13666;
																assign node13666 = (inp[12]) ? 4'b1011 : 4'b1111;
																assign node13669 = (inp[12]) ? 4'b1111 : 4'b1011;
															assign node13672 = (inp[12]) ? 4'b1101 : node13673;
																assign node13673 = (inp[4]) ? 4'b1011 : 4'b1111;
														assign node13677 = (inp[12]) ? node13679 : 4'b1001;
															assign node13679 = (inp[4]) ? node13681 : 4'b1001;
																assign node13681 = (inp[3]) ? 4'b1111 : 4'b1101;
													assign node13684 = (inp[15]) ? node13690 : node13685;
														assign node13685 = (inp[12]) ? node13687 : 4'b1001;
															assign node13687 = (inp[4]) ? 4'b1111 : 4'b1001;
														assign node13690 = (inp[4]) ? node13694 : node13691;
															assign node13691 = (inp[12]) ? 4'b1011 : 4'b1111;
															assign node13694 = (inp[12]) ? 4'b1111 : 4'b1011;
												assign node13697 = (inp[12]) ? node13719 : node13698;
													assign node13698 = (inp[4]) ? node13712 : node13699;
														assign node13699 = (inp[3]) ? node13707 : node13700;
															assign node13700 = (inp[0]) ? node13704 : node13701;
																assign node13701 = (inp[15]) ? 4'b1101 : 4'b1111;
																assign node13704 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node13707 = (inp[15]) ? node13709 : 4'b1101;
																assign node13709 = (inp[0]) ? 4'b1101 : 4'b1111;
														assign node13712 = (inp[15]) ? node13716 : node13713;
															assign node13713 = (inp[3]) ? 4'b1001 : 4'b1011;
															assign node13716 = (inp[3]) ? 4'b1011 : 4'b1001;
													assign node13719 = (inp[4]) ? node13733 : node13720;
														assign node13720 = (inp[15]) ? node13728 : node13721;
															assign node13721 = (inp[0]) ? node13725 : node13722;
																assign node13722 = (inp[3]) ? 4'b1001 : 4'b1011;
																assign node13725 = (inp[3]) ? 4'b1011 : 4'b1001;
															assign node13728 = (inp[3]) ? node13730 : 4'b1001;
																assign node13730 = (inp[0]) ? 4'b1001 : 4'b1011;
														assign node13733 = (inp[3]) ? 4'b1111 : node13734;
															assign node13734 = (inp[15]) ? node13736 : 4'b1101;
																assign node13736 = (inp[0]) ? 4'b1101 : 4'b1111;
											assign node13740 = (inp[12]) ? node13772 : node13741;
												assign node13741 = (inp[4]) ? node13763 : node13742;
													assign node13742 = (inp[3]) ? node13750 : node13743;
														assign node13743 = (inp[15]) ? node13747 : node13744;
															assign node13744 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node13747 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node13750 = (inp[15]) ? node13758 : node13751;
															assign node13751 = (inp[5]) ? node13755 : node13752;
																assign node13752 = (inp[0]) ? 4'b1001 : 4'b1011;
																assign node13755 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node13758 = (inp[0]) ? 4'b1001 : node13759;
																assign node13759 = (inp[5]) ? 4'b1011 : 4'b1001;
													assign node13763 = (inp[5]) ? node13765 : 4'b1111;
														assign node13765 = (inp[15]) ? node13769 : node13766;
															assign node13766 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node13769 = (inp[0]) ? 4'b1101 : 4'b1111;
												assign node13772 = (inp[4]) ? node13782 : node13773;
													assign node13773 = (inp[5]) ? node13779 : node13774;
														assign node13774 = (inp[3]) ? node13776 : 4'b1101;
															assign node13776 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node13779 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node13782 = (inp[5]) ? node13798 : node13783;
														assign node13783 = (inp[15]) ? node13791 : node13784;
															assign node13784 = (inp[3]) ? node13788 : node13785;
																assign node13785 = (inp[0]) ? 4'b1001 : 4'b1011;
																assign node13788 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node13791 = (inp[0]) ? node13795 : node13792;
																assign node13792 = (inp[3]) ? 4'b1011 : 4'b1001;
																assign node13795 = (inp[3]) ? 4'b1001 : 4'b1011;
														assign node13798 = (inp[3]) ? node13804 : node13799;
															assign node13799 = (inp[15]) ? node13801 : 4'b1001;
																assign node13801 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node13804 = (inp[15]) ? 4'b1001 : 4'b1011;
										assign node13807 = (inp[9]) ? node13891 : node13808;
											assign node13808 = (inp[15]) ? node13854 : node13809;
												assign node13809 = (inp[0]) ? node13831 : node13810;
													assign node13810 = (inp[3]) ? node13818 : node13811;
														assign node13811 = (inp[12]) ? node13815 : node13812;
															assign node13812 = (inp[4]) ? 4'b1010 : 4'b1110;
															assign node13815 = (inp[4]) ? 4'b1100 : 4'b1010;
														assign node13818 = (inp[5]) ? node13824 : node13819;
															assign node13819 = (inp[12]) ? 4'b1100 : node13820;
																assign node13820 = (inp[4]) ? 4'b1010 : 4'b1110;
															assign node13824 = (inp[4]) ? node13828 : node13825;
																assign node13825 = (inp[12]) ? 4'b1000 : 4'b1100;
																assign node13828 = (inp[12]) ? 4'b1100 : 4'b1000;
													assign node13831 = (inp[5]) ? node13847 : node13832;
														assign node13832 = (inp[3]) ? node13840 : node13833;
															assign node13833 = (inp[12]) ? node13837 : node13834;
																assign node13834 = (inp[4]) ? 4'b1000 : 4'b1100;
																assign node13837 = (inp[4]) ? 4'b1100 : 4'b1000;
															assign node13840 = (inp[12]) ? node13844 : node13841;
																assign node13841 = (inp[4]) ? 4'b1000 : 4'b1100;
																assign node13844 = (inp[4]) ? 4'b1110 : 4'b1000;
														assign node13847 = (inp[12]) ? node13851 : node13848;
															assign node13848 = (inp[3]) ? 4'b1010 : 4'b1000;
															assign node13851 = (inp[4]) ? 4'b1110 : 4'b1010;
												assign node13854 = (inp[0]) ? node13872 : node13855;
													assign node13855 = (inp[3]) ? node13861 : node13856;
														assign node13856 = (inp[5]) ? node13858 : 4'b1100;
															assign node13858 = (inp[12]) ? 4'b1000 : 4'b1100;
														assign node13861 = (inp[5]) ? node13867 : node13862;
															assign node13862 = (inp[12]) ? node13864 : 4'b1000;
																assign node13864 = (inp[4]) ? 4'b1110 : 4'b1000;
															assign node13867 = (inp[12]) ? node13869 : 4'b1110;
																assign node13869 = (inp[4]) ? 4'b1110 : 4'b1010;
													assign node13872 = (inp[3]) ? node13878 : node13873;
														assign node13873 = (inp[4]) ? 4'b1010 : node13874;
															assign node13874 = (inp[12]) ? 4'b1010 : 4'b1110;
														assign node13878 = (inp[5]) ? node13886 : node13879;
															assign node13879 = (inp[12]) ? node13883 : node13880;
																assign node13880 = (inp[4]) ? 4'b1010 : 4'b1110;
																assign node13883 = (inp[4]) ? 4'b1100 : 4'b1010;
															assign node13886 = (inp[4]) ? 4'b1100 : node13887;
																assign node13887 = (inp[12]) ? 4'b1000 : 4'b1100;
											assign node13891 = (inp[15]) ? node13931 : node13892;
												assign node13892 = (inp[0]) ? node13912 : node13893;
													assign node13893 = (inp[3]) ? node13905 : node13894;
														assign node13894 = (inp[5]) ? node13898 : node13895;
															assign node13895 = (inp[12]) ? 4'b1010 : 4'b1110;
															assign node13898 = (inp[12]) ? node13902 : node13899;
																assign node13899 = (inp[4]) ? 4'b1100 : 4'b1010;
																assign node13902 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node13905 = (inp[12]) ? node13909 : node13906;
															assign node13906 = (inp[4]) ? 4'b1100 : 4'b1000;
															assign node13909 = (inp[4]) ? 4'b1000 : 4'b1100;
													assign node13912 = (inp[5]) ? node13922 : node13913;
														assign node13913 = (inp[3]) ? 4'b1000 : node13914;
															assign node13914 = (inp[4]) ? node13918 : node13915;
																assign node13915 = (inp[12]) ? 4'b1100 : 4'b1000;
																assign node13918 = (inp[12]) ? 4'b1000 : 4'b1100;
														assign node13922 = (inp[4]) ? node13928 : node13923;
															assign node13923 = (inp[3]) ? node13925 : 4'b1000;
																assign node13925 = (inp[12]) ? 4'b1110 : 4'b1010;
															assign node13928 = (inp[12]) ? 4'b1010 : 4'b1110;
												assign node13931 = (inp[0]) ? node13945 : node13932;
													assign node13932 = (inp[12]) ? node13938 : node13933;
														assign node13933 = (inp[4]) ? node13935 : 4'b1000;
															assign node13935 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node13938 = (inp[4]) ? 4'b1010 : node13939;
															assign node13939 = (inp[5]) ? 4'b1110 : node13940;
																assign node13940 = (inp[3]) ? 4'b1110 : 4'b1100;
													assign node13945 = (inp[5]) ? node13959 : node13946;
														assign node13946 = (inp[3]) ? node13952 : node13947;
															assign node13947 = (inp[12]) ? node13949 : 4'b1010;
																assign node13949 = (inp[4]) ? 4'b1010 : 4'b1110;
															assign node13952 = (inp[4]) ? node13956 : node13953;
																assign node13953 = (inp[12]) ? 4'b1100 : 4'b1010;
																assign node13956 = (inp[12]) ? 4'b1000 : 4'b1100;
														assign node13959 = (inp[12]) ? node13965 : node13960;
															assign node13960 = (inp[4]) ? 4'b1100 : node13961;
																assign node13961 = (inp[3]) ? 4'b1000 : 4'b1010;
															assign node13965 = (inp[4]) ? 4'b1000 : 4'b1100;
							assign node13968 = (inp[4]) ? node14456 : node13969;
								assign node13969 = (inp[8]) ? node14205 : node13970;
									assign node13970 = (inp[7]) ? node14116 : node13971;
										assign node13971 = (inp[3]) ? node14043 : node13972;
											assign node13972 = (inp[2]) ? node14002 : node13973;
												assign node13973 = (inp[9]) ? node13987 : node13974;
													assign node13974 = (inp[12]) ? node13982 : node13975;
														assign node13975 = (inp[0]) ? node13979 : node13976;
															assign node13976 = (inp[15]) ? 4'b1100 : 4'b1110;
															assign node13979 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node13982 = (inp[5]) ? 4'b1000 : node13983;
															assign node13983 = (inp[0]) ? 4'b1010 : 4'b1000;
													assign node13987 = (inp[12]) ? node13995 : node13988;
														assign node13988 = (inp[5]) ? 4'b1010 : node13989;
															assign node13989 = (inp[15]) ? 4'b1010 : node13990;
																assign node13990 = (inp[0]) ? 4'b1000 : 4'b1010;
														assign node13995 = (inp[0]) ? 4'b1110 : node13996;
															assign node13996 = (inp[15]) ? 4'b1100 : node13997;
																assign node13997 = (inp[5]) ? 4'b1100 : 4'b1110;
												assign node14002 = (inp[5]) ? node14024 : node14003;
													assign node14003 = (inp[9]) ? node14013 : node14004;
														assign node14004 = (inp[12]) ? node14006 : 4'b1100;
															assign node14006 = (inp[0]) ? node14010 : node14007;
																assign node14007 = (inp[15]) ? 4'b1000 : 4'b1010;
																assign node14010 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node14013 = (inp[12]) ? node14019 : node14014;
															assign node14014 = (inp[0]) ? node14016 : 4'b1000;
																assign node14016 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node14019 = (inp[0]) ? node14021 : 4'b1100;
																assign node14021 = (inp[15]) ? 4'b1110 : 4'b1100;
													assign node14024 = (inp[15]) ? node14038 : node14025;
														assign node14025 = (inp[0]) ? node14033 : node14026;
															assign node14026 = (inp[9]) ? node14030 : node14027;
																assign node14027 = (inp[12]) ? 4'b1010 : 4'b1110;
																assign node14030 = (inp[12]) ? 4'b1100 : 4'b1010;
															assign node14033 = (inp[9]) ? 4'b1110 : node14034;
																assign node14034 = (inp[12]) ? 4'b1000 : 4'b1100;
														assign node14038 = (inp[0]) ? 4'b1100 : node14039;
															assign node14039 = (inp[12]) ? 4'b1000 : 4'b1100;
											assign node14043 = (inp[5]) ? node14071 : node14044;
												assign node14044 = (inp[9]) ? node14058 : node14045;
													assign node14045 = (inp[12]) ? node14051 : node14046;
														assign node14046 = (inp[2]) ? node14048 : 4'b1110;
															assign node14048 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node14051 = (inp[2]) ? 4'b1010 : node14052;
															assign node14052 = (inp[15]) ? node14054 : 4'b1010;
																assign node14054 = (inp[0]) ? 4'b1010 : 4'b1000;
													assign node14058 = (inp[12]) ? node14066 : node14059;
														assign node14059 = (inp[0]) ? node14063 : node14060;
															assign node14060 = (inp[15]) ? 4'b1000 : 4'b1010;
															assign node14063 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node14066 = (inp[15]) ? 4'b1110 : node14067;
															assign node14067 = (inp[0]) ? 4'b1110 : 4'b1100;
												assign node14071 = (inp[0]) ? node14095 : node14072;
													assign node14072 = (inp[15]) ? node14080 : node14073;
														assign node14073 = (inp[9]) ? node14077 : node14074;
															assign node14074 = (inp[12]) ? 4'b1000 : 4'b1100;
															assign node14077 = (inp[12]) ? 4'b1100 : 4'b1000;
														assign node14080 = (inp[2]) ? node14088 : node14081;
															assign node14081 = (inp[9]) ? node14085 : node14082;
																assign node14082 = (inp[12]) ? 4'b1010 : 4'b1110;
																assign node14085 = (inp[12]) ? 4'b1110 : 4'b1010;
															assign node14088 = (inp[12]) ? node14092 : node14089;
																assign node14089 = (inp[9]) ? 4'b1010 : 4'b1110;
																assign node14092 = (inp[9]) ? 4'b1110 : 4'b1010;
													assign node14095 = (inp[15]) ? node14103 : node14096;
														assign node14096 = (inp[12]) ? node14100 : node14097;
															assign node14097 = (inp[9]) ? 4'b1010 : 4'b1110;
															assign node14100 = (inp[9]) ? 4'b1110 : 4'b1010;
														assign node14103 = (inp[2]) ? node14111 : node14104;
															assign node14104 = (inp[12]) ? node14108 : node14105;
																assign node14105 = (inp[9]) ? 4'b1000 : 4'b1100;
																assign node14108 = (inp[9]) ? 4'b1100 : 4'b1000;
															assign node14111 = (inp[12]) ? node14113 : 4'b1100;
																assign node14113 = (inp[9]) ? 4'b1100 : 4'b1000;
										assign node14116 = (inp[0]) ? node14164 : node14117;
											assign node14117 = (inp[15]) ? node14141 : node14118;
												assign node14118 = (inp[5]) ? node14128 : node14119;
													assign node14119 = (inp[9]) ? node14123 : node14120;
														assign node14120 = (inp[12]) ? 4'b1011 : 4'b1111;
														assign node14123 = (inp[12]) ? node14125 : 4'b1011;
															assign node14125 = (inp[3]) ? 4'b1101 : 4'b1111;
													assign node14128 = (inp[3]) ? node14134 : node14129;
														assign node14129 = (inp[12]) ? 4'b1101 : node14130;
															assign node14130 = (inp[9]) ? 4'b1011 : 4'b1111;
														assign node14134 = (inp[9]) ? node14138 : node14135;
															assign node14135 = (inp[12]) ? 4'b1001 : 4'b1101;
															assign node14138 = (inp[12]) ? 4'b1101 : 4'b1001;
												assign node14141 = (inp[3]) ? node14153 : node14142;
													assign node14142 = (inp[2]) ? node14148 : node14143;
														assign node14143 = (inp[12]) ? node14145 : 4'b1101;
															assign node14145 = (inp[9]) ? 4'b1101 : 4'b1001;
														assign node14148 = (inp[5]) ? 4'b1001 : node14149;
															assign node14149 = (inp[9]) ? 4'b1101 : 4'b1001;
													assign node14153 = (inp[5]) ? node14157 : node14154;
														assign node14154 = (inp[9]) ? 4'b1001 : 4'b1101;
														assign node14157 = (inp[12]) ? node14161 : node14158;
															assign node14158 = (inp[9]) ? 4'b1011 : 4'b1111;
															assign node14161 = (inp[9]) ? 4'b1111 : 4'b1011;
											assign node14164 = (inp[12]) ? node14182 : node14165;
												assign node14165 = (inp[9]) ? node14171 : node14166;
													assign node14166 = (inp[15]) ? node14168 : 4'b1101;
														assign node14168 = (inp[5]) ? 4'b1101 : 4'b1111;
													assign node14171 = (inp[15]) ? node14177 : node14172;
														assign node14172 = (inp[3]) ? node14174 : 4'b1001;
															assign node14174 = (inp[5]) ? 4'b1011 : 4'b1001;
														assign node14177 = (inp[2]) ? 4'b1011 : node14178;
															assign node14178 = (inp[5]) ? 4'b1001 : 4'b1011;
												assign node14182 = (inp[9]) ? node14194 : node14183;
													assign node14183 = (inp[15]) ? node14189 : node14184;
														assign node14184 = (inp[3]) ? node14186 : 4'b1001;
															assign node14186 = (inp[5]) ? 4'b1011 : 4'b1001;
														assign node14189 = (inp[5]) ? node14191 : 4'b1011;
															assign node14191 = (inp[3]) ? 4'b1001 : 4'b1011;
													assign node14194 = (inp[15]) ? node14200 : node14195;
														assign node14195 = (inp[5]) ? 4'b1111 : node14196;
															assign node14196 = (inp[3]) ? 4'b1111 : 4'b1101;
														assign node14200 = (inp[3]) ? 4'b1101 : node14201;
															assign node14201 = (inp[2]) ? 4'b1101 : 4'b1111;
									assign node14205 = (inp[7]) ? node14325 : node14206;
										assign node14206 = (inp[9]) ? node14268 : node14207;
											assign node14207 = (inp[12]) ? node14229 : node14208;
												assign node14208 = (inp[5]) ? node14216 : node14209;
													assign node14209 = (inp[0]) ? node14213 : node14210;
														assign node14210 = (inp[15]) ? 4'b1101 : 4'b1111;
														assign node14213 = (inp[15]) ? 4'b1111 : 4'b1101;
													assign node14216 = (inp[0]) ? node14224 : node14217;
														assign node14217 = (inp[15]) ? node14221 : node14218;
															assign node14218 = (inp[3]) ? 4'b1101 : 4'b1111;
															assign node14221 = (inp[3]) ? 4'b1111 : 4'b1101;
														assign node14224 = (inp[3]) ? node14226 : 4'b1111;
															assign node14226 = (inp[15]) ? 4'b1101 : 4'b1111;
												assign node14229 = (inp[3]) ? node14245 : node14230;
													assign node14230 = (inp[5]) ? node14240 : node14231;
														assign node14231 = (inp[2]) ? node14237 : node14232;
															assign node14232 = (inp[15]) ? node14234 : 4'b1011;
																assign node14234 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node14237 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node14240 = (inp[2]) ? 4'b1011 : node14241;
															assign node14241 = (inp[15]) ? 4'b1001 : 4'b1011;
													assign node14245 = (inp[2]) ? node14255 : node14246;
														assign node14246 = (inp[15]) ? node14248 : 4'b1001;
															assign node14248 = (inp[0]) ? node14252 : node14249;
																assign node14249 = (inp[5]) ? 4'b1011 : 4'b1001;
																assign node14252 = (inp[5]) ? 4'b1001 : 4'b1011;
														assign node14255 = (inp[0]) ? node14263 : node14256;
															assign node14256 = (inp[15]) ? node14260 : node14257;
																assign node14257 = (inp[5]) ? 4'b1001 : 4'b1011;
																assign node14260 = (inp[5]) ? 4'b1011 : 4'b1001;
															assign node14263 = (inp[5]) ? node14265 : 4'b1001;
																assign node14265 = (inp[15]) ? 4'b1001 : 4'b1011;
											assign node14268 = (inp[12]) ? node14288 : node14269;
												assign node14269 = (inp[15]) ? node14279 : node14270;
													assign node14270 = (inp[0]) ? node14276 : node14271;
														assign node14271 = (inp[5]) ? node14273 : 4'b1011;
															assign node14273 = (inp[2]) ? 4'b1011 : 4'b1001;
														assign node14276 = (inp[5]) ? 4'b1011 : 4'b1001;
													assign node14279 = (inp[0]) ? node14283 : node14280;
														assign node14280 = (inp[3]) ? 4'b1011 : 4'b1001;
														assign node14283 = (inp[3]) ? node14285 : 4'b1011;
															assign node14285 = (inp[5]) ? 4'b1001 : 4'b1011;
												assign node14288 = (inp[5]) ? node14302 : node14289;
													assign node14289 = (inp[0]) ? node14297 : node14290;
														assign node14290 = (inp[3]) ? node14294 : node14291;
															assign node14291 = (inp[15]) ? 4'b1101 : 4'b1111;
															assign node14294 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node14297 = (inp[3]) ? node14299 : 4'b1111;
															assign node14299 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node14302 = (inp[3]) ? node14310 : node14303;
														assign node14303 = (inp[0]) ? node14307 : node14304;
															assign node14304 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node14307 = (inp[15]) ? 4'b1101 : 4'b1111;
														assign node14310 = (inp[2]) ? node14318 : node14311;
															assign node14311 = (inp[0]) ? node14315 : node14312;
																assign node14312 = (inp[15]) ? 4'b1111 : 4'b1101;
																assign node14315 = (inp[15]) ? 4'b1101 : 4'b1111;
															assign node14318 = (inp[0]) ? node14322 : node14319;
																assign node14319 = (inp[15]) ? 4'b1111 : 4'b1101;
																assign node14322 = (inp[15]) ? 4'b1101 : 4'b1111;
										assign node14325 = (inp[3]) ? node14391 : node14326;
											assign node14326 = (inp[2]) ? node14364 : node14327;
												assign node14327 = (inp[12]) ? node14345 : node14328;
													assign node14328 = (inp[9]) ? node14340 : node14329;
														assign node14329 = (inp[5]) ? node14335 : node14330;
															assign node14330 = (inp[15]) ? node14332 : 4'b1100;
																assign node14332 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node14335 = (inp[0]) ? node14337 : 4'b1110;
																assign node14337 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node14340 = (inp[5]) ? node14342 : 4'b1010;
															assign node14342 = (inp[0]) ? 4'b1000 : 4'b1010;
													assign node14345 = (inp[9]) ? node14353 : node14346;
														assign node14346 = (inp[0]) ? node14350 : node14347;
															assign node14347 = (inp[15]) ? 4'b1000 : 4'b1010;
															assign node14350 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node14353 = (inp[5]) ? node14359 : node14354;
															assign node14354 = (inp[15]) ? 4'b1100 : node14355;
																assign node14355 = (inp[0]) ? 4'b1100 : 4'b1110;
															assign node14359 = (inp[15]) ? node14361 : 4'b1110;
																assign node14361 = (inp[0]) ? 4'b1100 : 4'b1110;
												assign node14364 = (inp[15]) ? node14378 : node14365;
													assign node14365 = (inp[0]) ? node14373 : node14366;
														assign node14366 = (inp[12]) ? node14370 : node14367;
															assign node14367 = (inp[9]) ? 4'b1010 : 4'b1110;
															assign node14370 = (inp[5]) ? 4'b1100 : 4'b1110;
														assign node14373 = (inp[12]) ? node14375 : 4'b1100;
															assign node14375 = (inp[5]) ? 4'b1110 : 4'b1100;
													assign node14378 = (inp[0]) ? node14386 : node14379;
														assign node14379 = (inp[9]) ? node14383 : node14380;
															assign node14380 = (inp[12]) ? 4'b1000 : 4'b1100;
															assign node14383 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node14386 = (inp[9]) ? 4'b1100 : node14387;
															assign node14387 = (inp[12]) ? 4'b1010 : 4'b1110;
											assign node14391 = (inp[15]) ? node14429 : node14392;
												assign node14392 = (inp[0]) ? node14412 : node14393;
													assign node14393 = (inp[5]) ? node14399 : node14394;
														assign node14394 = (inp[2]) ? node14396 : 4'b1010;
															assign node14396 = (inp[9]) ? 4'b1010 : 4'b1110;
														assign node14399 = (inp[2]) ? node14405 : node14400;
															assign node14400 = (inp[12]) ? node14402 : 4'b1000;
																assign node14402 = (inp[9]) ? 4'b1100 : 4'b1000;
															assign node14405 = (inp[9]) ? node14409 : node14406;
																assign node14406 = (inp[12]) ? 4'b1000 : 4'b1100;
																assign node14409 = (inp[12]) ? 4'b1100 : 4'b1000;
													assign node14412 = (inp[5]) ? node14420 : node14413;
														assign node14413 = (inp[12]) ? node14417 : node14414;
															assign node14414 = (inp[9]) ? 4'b1000 : 4'b1100;
															assign node14417 = (inp[9]) ? 4'b1110 : 4'b1000;
														assign node14420 = (inp[2]) ? 4'b1010 : node14421;
															assign node14421 = (inp[9]) ? node14425 : node14422;
																assign node14422 = (inp[12]) ? 4'b1010 : 4'b1110;
																assign node14425 = (inp[12]) ? 4'b1110 : 4'b1010;
												assign node14429 = (inp[0]) ? node14445 : node14430;
													assign node14430 = (inp[5]) ? node14434 : node14431;
														assign node14431 = (inp[9]) ? 4'b1110 : 4'b1100;
														assign node14434 = (inp[2]) ? node14440 : node14435;
															assign node14435 = (inp[12]) ? 4'b1110 : node14436;
																assign node14436 = (inp[9]) ? 4'b1010 : 4'b1110;
															assign node14440 = (inp[9]) ? 4'b1010 : node14441;
																assign node14441 = (inp[12]) ? 4'b1010 : 4'b1110;
													assign node14445 = (inp[5]) ? node14453 : node14446;
														assign node14446 = (inp[12]) ? node14450 : node14447;
															assign node14447 = (inp[9]) ? 4'b1010 : 4'b1110;
															assign node14450 = (inp[9]) ? 4'b1100 : 4'b1010;
														assign node14453 = (inp[12]) ? 4'b1100 : 4'b1000;
								assign node14456 = (inp[7]) ? node14654 : node14457;
									assign node14457 = (inp[8]) ? node14569 : node14458;
										assign node14458 = (inp[0]) ? node14516 : node14459;
											assign node14459 = (inp[15]) ? node14483 : node14460;
												assign node14460 = (inp[3]) ? node14474 : node14461;
													assign node14461 = (inp[5]) ? node14467 : node14462;
														assign node14462 = (inp[9]) ? node14464 : 4'b1110;
															assign node14464 = (inp[12]) ? 4'b1010 : 4'b1110;
														assign node14467 = (inp[2]) ? node14469 : 4'b1100;
															assign node14469 = (inp[12]) ? node14471 : 4'b1010;
																assign node14471 = (inp[9]) ? 4'b1000 : 4'b1100;
													assign node14474 = (inp[12]) ? node14480 : node14475;
														assign node14475 = (inp[9]) ? 4'b1100 : node14476;
															assign node14476 = (inp[5]) ? 4'b1000 : 4'b1010;
														assign node14480 = (inp[9]) ? 4'b1000 : 4'b1100;
												assign node14483 = (inp[3]) ? node14499 : node14484;
													assign node14484 = (inp[5]) ? node14492 : node14485;
														assign node14485 = (inp[9]) ? node14489 : node14486;
															assign node14486 = (inp[12]) ? 4'b1100 : 4'b1000;
															assign node14489 = (inp[12]) ? 4'b1000 : 4'b1100;
														assign node14492 = (inp[2]) ? 4'b1110 : node14493;
															assign node14493 = (inp[9]) ? node14495 : 4'b1000;
																assign node14495 = (inp[12]) ? 4'b1010 : 4'b1110;
													assign node14499 = (inp[5]) ? node14507 : node14500;
														assign node14500 = (inp[2]) ? 4'b1110 : node14501;
															assign node14501 = (inp[12]) ? node14503 : 4'b1000;
																assign node14503 = (inp[9]) ? 4'b1010 : 4'b1110;
														assign node14507 = (inp[2]) ? 4'b1010 : node14508;
															assign node14508 = (inp[12]) ? node14512 : node14509;
																assign node14509 = (inp[9]) ? 4'b1110 : 4'b1010;
																assign node14512 = (inp[9]) ? 4'b1010 : 4'b1110;
											assign node14516 = (inp[15]) ? node14536 : node14517;
												assign node14517 = (inp[3]) ? node14527 : node14518;
													assign node14518 = (inp[5]) ? node14522 : node14519;
														assign node14519 = (inp[2]) ? 4'b1000 : 4'b1100;
														assign node14522 = (inp[12]) ? node14524 : 4'b1000;
															assign node14524 = (inp[9]) ? 4'b1010 : 4'b1110;
													assign node14527 = (inp[9]) ? node14533 : node14528;
														assign node14528 = (inp[12]) ? 4'b1110 : node14529;
															assign node14529 = (inp[5]) ? 4'b1010 : 4'b1000;
														assign node14533 = (inp[12]) ? 4'b1010 : 4'b1110;
												assign node14536 = (inp[5]) ? node14550 : node14537;
													assign node14537 = (inp[3]) ? node14543 : node14538;
														assign node14538 = (inp[12]) ? 4'b1110 : node14539;
															assign node14539 = (inp[9]) ? 4'b1110 : 4'b1010;
														assign node14543 = (inp[2]) ? node14547 : node14544;
															assign node14544 = (inp[12]) ? 4'b1100 : 4'b1010;
															assign node14547 = (inp[12]) ? 4'b1000 : 4'b1100;
													assign node14550 = (inp[3]) ? node14558 : node14551;
														assign node14551 = (inp[9]) ? node14555 : node14552;
															assign node14552 = (inp[12]) ? 4'b1100 : 4'b1010;
															assign node14555 = (inp[12]) ? 4'b1000 : 4'b1100;
														assign node14558 = (inp[2]) ? node14564 : node14559;
															assign node14559 = (inp[12]) ? node14561 : 4'b1100;
																assign node14561 = (inp[9]) ? 4'b1000 : 4'b1100;
															assign node14564 = (inp[12]) ? 4'b1100 : node14565;
																assign node14565 = (inp[9]) ? 4'b1100 : 4'b1000;
										assign node14569 = (inp[12]) ? node14611 : node14570;
											assign node14570 = (inp[9]) ? node14588 : node14571;
												assign node14571 = (inp[15]) ? node14579 : node14572;
													assign node14572 = (inp[0]) ? node14574 : 4'b1011;
														assign node14574 = (inp[5]) ? node14576 : 4'b1001;
															assign node14576 = (inp[3]) ? 4'b1011 : 4'b1001;
													assign node14579 = (inp[0]) ? node14585 : node14580;
														assign node14580 = (inp[5]) ? node14582 : 4'b1001;
															assign node14582 = (inp[2]) ? 4'b1011 : 4'b1001;
														assign node14585 = (inp[3]) ? 4'b1001 : 4'b1011;
												assign node14588 = (inp[0]) ? node14600 : node14589;
													assign node14589 = (inp[15]) ? node14595 : node14590;
														assign node14590 = (inp[5]) ? 4'b1101 : node14591;
															assign node14591 = (inp[3]) ? 4'b1101 : 4'b1111;
														assign node14595 = (inp[3]) ? 4'b1111 : node14596;
															assign node14596 = (inp[5]) ? 4'b1111 : 4'b1101;
													assign node14600 = (inp[15]) ? node14608 : node14601;
														assign node14601 = (inp[2]) ? node14603 : 4'b1111;
															assign node14603 = (inp[3]) ? 4'b1111 : node14604;
																assign node14604 = (inp[5]) ? 4'b1111 : 4'b1101;
														assign node14608 = (inp[3]) ? 4'b1101 : 4'b1111;
											assign node14611 = (inp[9]) ? node14631 : node14612;
												assign node14612 = (inp[0]) ? node14622 : node14613;
													assign node14613 = (inp[15]) ? node14619 : node14614;
														assign node14614 = (inp[3]) ? 4'b1101 : node14615;
															assign node14615 = (inp[5]) ? 4'b1101 : 4'b1111;
														assign node14619 = (inp[5]) ? 4'b1111 : 4'b1101;
													assign node14622 = (inp[15]) ? node14626 : node14623;
														assign node14623 = (inp[3]) ? 4'b1111 : 4'b1101;
														assign node14626 = (inp[5]) ? 4'b1101 : node14627;
															assign node14627 = (inp[3]) ? 4'b1101 : 4'b1111;
												assign node14631 = (inp[2]) ? node14643 : node14632;
													assign node14632 = (inp[5]) ? 4'b1001 : node14633;
														assign node14633 = (inp[0]) ? 4'b1001 : node14634;
															assign node14634 = (inp[3]) ? node14638 : node14635;
																assign node14635 = (inp[15]) ? 4'b1001 : 4'b1011;
																assign node14638 = (inp[15]) ? 4'b1011 : 4'b1001;
													assign node14643 = (inp[3]) ? 4'b1011 : node14644;
														assign node14644 = (inp[5]) ? node14646 : 4'b1001;
															assign node14646 = (inp[0]) ? node14650 : node14647;
																assign node14647 = (inp[15]) ? 4'b1011 : 4'b1001;
																assign node14650 = (inp[15]) ? 4'b1001 : 4'b1011;
									assign node14654 = (inp[8]) ? node14802 : node14655;
										assign node14655 = (inp[2]) ? node14731 : node14656;
											assign node14656 = (inp[0]) ? node14696 : node14657;
												assign node14657 = (inp[15]) ? node14677 : node14658;
													assign node14658 = (inp[5]) ? node14670 : node14659;
														assign node14659 = (inp[3]) ? node14665 : node14660;
															assign node14660 = (inp[9]) ? node14662 : 4'b1111;
																assign node14662 = (inp[12]) ? 4'b1011 : 4'b1111;
															assign node14665 = (inp[12]) ? 4'b1101 : node14666;
																assign node14666 = (inp[9]) ? 4'b1101 : 4'b1011;
														assign node14670 = (inp[9]) ? node14674 : node14671;
															assign node14671 = (inp[3]) ? 4'b1001 : 4'b1101;
															assign node14674 = (inp[12]) ? 4'b1001 : 4'b1101;
													assign node14677 = (inp[5]) ? node14689 : node14678;
														assign node14678 = (inp[3]) ? node14684 : node14679;
															assign node14679 = (inp[9]) ? 4'b1001 : node14680;
																assign node14680 = (inp[12]) ? 4'b1101 : 4'b1001;
															assign node14684 = (inp[9]) ? 4'b1111 : node14685;
																assign node14685 = (inp[12]) ? 4'b1111 : 4'b1001;
														assign node14689 = (inp[9]) ? node14693 : node14690;
															assign node14690 = (inp[12]) ? 4'b1111 : 4'b1001;
															assign node14693 = (inp[12]) ? 4'b1011 : 4'b1111;
												assign node14696 = (inp[15]) ? node14714 : node14697;
													assign node14697 = (inp[3]) ? node14707 : node14698;
														assign node14698 = (inp[5]) ? node14700 : 4'b1001;
															assign node14700 = (inp[12]) ? node14704 : node14701;
																assign node14701 = (inp[9]) ? 4'b1111 : 4'b1001;
																assign node14704 = (inp[9]) ? 4'b1011 : 4'b1111;
														assign node14707 = (inp[12]) ? node14711 : node14708;
															assign node14708 = (inp[9]) ? 4'b1111 : 4'b1011;
															assign node14711 = (inp[9]) ? 4'b1011 : 4'b1111;
													assign node14714 = (inp[3]) ? node14724 : node14715;
														assign node14715 = (inp[5]) ? node14721 : node14716;
															assign node14716 = (inp[12]) ? node14718 : 4'b1011;
																assign node14718 = (inp[9]) ? 4'b1011 : 4'b1111;
															assign node14721 = (inp[12]) ? 4'b1001 : 4'b1011;
														assign node14724 = (inp[5]) ? 4'b1101 : node14725;
															assign node14725 = (inp[9]) ? node14727 : 4'b1011;
																assign node14727 = (inp[12]) ? 4'b1001 : 4'b1101;
											assign node14731 = (inp[9]) ? node14767 : node14732;
												assign node14732 = (inp[12]) ? node14748 : node14733;
													assign node14733 = (inp[3]) ? node14741 : node14734;
														assign node14734 = (inp[5]) ? 4'b1011 : node14735;
															assign node14735 = (inp[15]) ? 4'b1001 : node14736;
																assign node14736 = (inp[0]) ? 4'b1001 : 4'b1011;
														assign node14741 = (inp[5]) ? node14743 : 4'b1001;
															assign node14743 = (inp[15]) ? node14745 : 4'b1001;
																assign node14745 = (inp[0]) ? 4'b1001 : 4'b1011;
													assign node14748 = (inp[15]) ? node14756 : node14749;
														assign node14749 = (inp[0]) ? node14751 : 4'b1101;
															assign node14751 = (inp[5]) ? 4'b1111 : node14752;
																assign node14752 = (inp[3]) ? 4'b1111 : 4'b1101;
														assign node14756 = (inp[0]) ? node14762 : node14757;
															assign node14757 = (inp[5]) ? 4'b1111 : node14758;
																assign node14758 = (inp[3]) ? 4'b1111 : 4'b1101;
															assign node14762 = (inp[3]) ? 4'b1101 : node14763;
																assign node14763 = (inp[5]) ? 4'b1101 : 4'b1111;
												assign node14767 = (inp[12]) ? node14783 : node14768;
													assign node14768 = (inp[3]) ? node14776 : node14769;
														assign node14769 = (inp[0]) ? 4'b1111 : node14770;
															assign node14770 = (inp[5]) ? 4'b1111 : node14771;
																assign node14771 = (inp[15]) ? 4'b1101 : 4'b1111;
														assign node14776 = (inp[0]) ? node14780 : node14777;
															assign node14777 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node14780 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node14783 = (inp[15]) ? node14793 : node14784;
														assign node14784 = (inp[0]) ? node14790 : node14785;
															assign node14785 = (inp[5]) ? 4'b1001 : node14786;
																assign node14786 = (inp[3]) ? 4'b1001 : 4'b1011;
															assign node14790 = (inp[3]) ? 4'b1011 : 4'b1001;
														assign node14793 = (inp[5]) ? 4'b1011 : node14794;
															assign node14794 = (inp[3]) ? node14798 : node14795;
																assign node14795 = (inp[0]) ? 4'b1011 : 4'b1001;
																assign node14798 = (inp[0]) ? 4'b1001 : 4'b1011;
										assign node14802 = (inp[12]) ? node14860 : node14803;
											assign node14803 = (inp[9]) ? node14833 : node14804;
												assign node14804 = (inp[5]) ? node14820 : node14805;
													assign node14805 = (inp[3]) ? node14815 : node14806;
														assign node14806 = (inp[2]) ? node14810 : node14807;
															assign node14807 = (inp[0]) ? 4'b1010 : 4'b1000;
															assign node14810 = (inp[0]) ? node14812 : 4'b1010;
																assign node14812 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node14815 = (inp[15]) ? 4'b1000 : node14816;
															assign node14816 = (inp[0]) ? 4'b1000 : 4'b1010;
													assign node14820 = (inp[3]) ? node14826 : node14821;
														assign node14821 = (inp[0]) ? 4'b1010 : node14822;
															assign node14822 = (inp[15]) ? 4'b1000 : 4'b1010;
														assign node14826 = (inp[0]) ? node14830 : node14827;
															assign node14827 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node14830 = (inp[15]) ? 4'b1000 : 4'b1010;
												assign node14833 = (inp[5]) ? node14847 : node14834;
													assign node14834 = (inp[15]) ? node14840 : node14835;
														assign node14835 = (inp[0]) ? 4'b1110 : node14836;
															assign node14836 = (inp[3]) ? 4'b1100 : 4'b1110;
														assign node14840 = (inp[3]) ? node14844 : node14841;
															assign node14841 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node14844 = (inp[0]) ? 4'b1100 : 4'b1110;
													assign node14847 = (inp[2]) ? node14855 : node14848;
														assign node14848 = (inp[0]) ? node14852 : node14849;
															assign node14849 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node14852 = (inp[15]) ? 4'b1100 : 4'b1110;
														assign node14855 = (inp[15]) ? 4'b1100 : node14856;
															assign node14856 = (inp[0]) ? 4'b1110 : 4'b1100;
											assign node14860 = (inp[9]) ? node14884 : node14861;
												assign node14861 = (inp[0]) ? node14873 : node14862;
													assign node14862 = (inp[15]) ? node14868 : node14863;
														assign node14863 = (inp[3]) ? 4'b1100 : node14864;
															assign node14864 = (inp[5]) ? 4'b1100 : 4'b1110;
														assign node14868 = (inp[3]) ? 4'b1110 : node14869;
															assign node14869 = (inp[5]) ? 4'b1110 : 4'b1100;
													assign node14873 = (inp[15]) ? node14879 : node14874;
														assign node14874 = (inp[5]) ? 4'b1110 : node14875;
															assign node14875 = (inp[3]) ? 4'b1110 : 4'b1100;
														assign node14879 = (inp[2]) ? 4'b1100 : node14880;
															assign node14880 = (inp[5]) ? 4'b1100 : 4'b1110;
												assign node14884 = (inp[2]) ? node14898 : node14885;
													assign node14885 = (inp[15]) ? node14891 : node14886;
														assign node14886 = (inp[0]) ? 4'b1010 : node14887;
															assign node14887 = (inp[5]) ? 4'b1000 : 4'b1010;
														assign node14891 = (inp[0]) ? 4'b1000 : node14892;
															assign node14892 = (inp[5]) ? 4'b1010 : node14893;
																assign node14893 = (inp[3]) ? 4'b1010 : 4'b1000;
													assign node14898 = (inp[5]) ? node14908 : node14899;
														assign node14899 = (inp[15]) ? 4'b1000 : node14900;
															assign node14900 = (inp[0]) ? node14904 : node14901;
																assign node14901 = (inp[3]) ? 4'b1000 : 4'b1010;
																assign node14904 = (inp[3]) ? 4'b1010 : 4'b1000;
														assign node14908 = (inp[3]) ? node14916 : node14909;
															assign node14909 = (inp[15]) ? node14913 : node14910;
																assign node14910 = (inp[0]) ? 4'b1010 : 4'b1000;
																assign node14913 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node14916 = (inp[15]) ? node14920 : node14917;
																assign node14917 = (inp[0]) ? 4'b1010 : 4'b1000;
																assign node14920 = (inp[0]) ? 4'b1000 : 4'b1010;
			assign node14923 = (inp[11]) ? node22797 : node14924;
				assign node14924 = (inp[1]) ? node18668 : node14925;
					assign node14925 = (inp[13]) ? node16721 : node14926;
						assign node14926 = (inp[3]) ? node15772 : node14927;
							assign node14927 = (inp[14]) ? node15473 : node14928;
								assign node14928 = (inp[12]) ? node15190 : node14929;
									assign node14929 = (inp[2]) ? node15055 : node14930;
										assign node14930 = (inp[0]) ? node14990 : node14931;
											assign node14931 = (inp[15]) ? node14955 : node14932;
												assign node14932 = (inp[4]) ? node14944 : node14933;
													assign node14933 = (inp[9]) ? node14939 : node14934;
														assign node14934 = (inp[5]) ? node14936 : 4'b0111;
															assign node14936 = (inp[7]) ? 4'b0110 : 4'b0111;
														assign node14939 = (inp[7]) ? node14941 : 4'b0011;
															assign node14941 = (inp[8]) ? 4'b0011 : 4'b0010;
													assign node14944 = (inp[9]) ? node14950 : node14945;
														assign node14945 = (inp[7]) ? node14947 : 4'b0010;
															assign node14947 = (inp[5]) ? 4'b0011 : 4'b0010;
														assign node14950 = (inp[5]) ? 4'b0100 : node14951;
															assign node14951 = (inp[7]) ? 4'b0110 : 4'b0111;
												assign node14955 = (inp[7]) ? node14971 : node14956;
													assign node14956 = (inp[8]) ? node14966 : node14957;
														assign node14957 = (inp[4]) ? node14961 : node14958;
															assign node14958 = (inp[9]) ? 4'b0001 : 4'b0101;
															assign node14961 = (inp[9]) ? node14963 : 4'b0001;
																assign node14963 = (inp[5]) ? 4'b0111 : 4'b0101;
														assign node14966 = (inp[9]) ? 4'b0000 : node14967;
															assign node14967 = (inp[4]) ? 4'b0000 : 4'b0100;
													assign node14971 = (inp[8]) ? node14981 : node14972;
														assign node14972 = (inp[5]) ? node14978 : node14973;
															assign node14973 = (inp[4]) ? 4'b0100 : node14974;
																assign node14974 = (inp[9]) ? 4'b0000 : 4'b0100;
															assign node14978 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node14981 = (inp[5]) ? 4'b0111 : node14982;
															assign node14982 = (inp[9]) ? node14986 : node14983;
																assign node14983 = (inp[4]) ? 4'b0001 : 4'b0101;
																assign node14986 = (inp[4]) ? 4'b0101 : 4'b0001;
											assign node14990 = (inp[15]) ? node15026 : node14991;
												assign node14991 = (inp[4]) ? node15009 : node14992;
													assign node14992 = (inp[9]) ? node15002 : node14993;
														assign node14993 = (inp[5]) ? node14995 : 4'b0101;
															assign node14995 = (inp[8]) ? node14999 : node14996;
																assign node14996 = (inp[7]) ? 4'b0100 : 4'b0101;
																assign node14999 = (inp[7]) ? 4'b0101 : 4'b0100;
														assign node15002 = (inp[8]) ? node15006 : node15003;
															assign node15003 = (inp[7]) ? 4'b0000 : 4'b0001;
															assign node15006 = (inp[7]) ? 4'b0001 : 4'b0000;
													assign node15009 = (inp[9]) ? node15015 : node15010;
														assign node15010 = (inp[7]) ? node15012 : 4'b0001;
															assign node15012 = (inp[8]) ? 4'b0001 : 4'b0000;
														assign node15015 = (inp[5]) ? node15021 : node15016;
															assign node15016 = (inp[7]) ? 4'b0100 : node15017;
																assign node15017 = (inp[8]) ? 4'b0100 : 4'b0101;
															assign node15021 = (inp[7]) ? node15023 : 4'b0110;
																assign node15023 = (inp[8]) ? 4'b0111 : 4'b0110;
												assign node15026 = (inp[8]) ? node15036 : node15027;
													assign node15027 = (inp[7]) ? 4'b0010 : node15028;
														assign node15028 = (inp[4]) ? node15032 : node15029;
															assign node15029 = (inp[9]) ? 4'b0011 : 4'b0111;
															assign node15032 = (inp[9]) ? 4'b0111 : 4'b0011;
													assign node15036 = (inp[7]) ? node15046 : node15037;
														assign node15037 = (inp[5]) ? 4'b0010 : node15038;
															assign node15038 = (inp[4]) ? node15042 : node15039;
																assign node15039 = (inp[9]) ? 4'b0010 : 4'b0110;
																assign node15042 = (inp[9]) ? 4'b0110 : 4'b0010;
														assign node15046 = (inp[9]) ? node15050 : node15047;
															assign node15047 = (inp[4]) ? 4'b0011 : 4'b0111;
															assign node15050 = (inp[5]) ? 4'b0101 : node15051;
																assign node15051 = (inp[4]) ? 4'b0111 : 4'b0011;
										assign node15055 = (inp[9]) ? node15123 : node15056;
											assign node15056 = (inp[4]) ? node15082 : node15057;
												assign node15057 = (inp[8]) ? node15071 : node15058;
													assign node15058 = (inp[7]) ? node15064 : node15059;
														assign node15059 = (inp[15]) ? node15061 : 4'b0100;
															assign node15061 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node15064 = (inp[15]) ? node15068 : node15065;
															assign node15065 = (inp[0]) ? 4'b0101 : 4'b0111;
															assign node15068 = (inp[0]) ? 4'b0111 : 4'b0101;
													assign node15071 = (inp[7]) ? node15075 : node15072;
														assign node15072 = (inp[0]) ? 4'b0101 : 4'b0111;
														assign node15075 = (inp[5]) ? 4'b0110 : node15076;
															assign node15076 = (inp[15]) ? node15078 : 4'b0100;
																assign node15078 = (inp[0]) ? 4'b0110 : 4'b0100;
												assign node15082 = (inp[5]) ? node15108 : node15083;
													assign node15083 = (inp[7]) ? node15097 : node15084;
														assign node15084 = (inp[8]) ? node15092 : node15085;
															assign node15085 = (inp[15]) ? node15089 : node15086;
																assign node15086 = (inp[0]) ? 4'b0000 : 4'b0010;
																assign node15089 = (inp[0]) ? 4'b0010 : 4'b0000;
															assign node15092 = (inp[0]) ? 4'b0001 : node15093;
																assign node15093 = (inp[15]) ? 4'b0001 : 4'b0011;
														assign node15097 = (inp[8]) ? node15101 : node15098;
															assign node15098 = (inp[0]) ? 4'b0011 : 4'b0001;
															assign node15101 = (inp[15]) ? node15105 : node15102;
																assign node15102 = (inp[0]) ? 4'b0000 : 4'b0010;
																assign node15105 = (inp[0]) ? 4'b0010 : 4'b0000;
													assign node15108 = (inp[15]) ? node15116 : node15109;
														assign node15109 = (inp[0]) ? 4'b0001 : node15110;
															assign node15110 = (inp[7]) ? 4'b0011 : node15111;
																assign node15111 = (inp[8]) ? 4'b0011 : 4'b0010;
														assign node15116 = (inp[0]) ? node15118 : 4'b0001;
															assign node15118 = (inp[8]) ? 4'b0010 : node15119;
																assign node15119 = (inp[7]) ? 4'b0011 : 4'b0010;
											assign node15123 = (inp[4]) ? node15149 : node15124;
												assign node15124 = (inp[0]) ? node15140 : node15125;
													assign node15125 = (inp[15]) ? node15131 : node15126;
														assign node15126 = (inp[8]) ? 4'b0010 : node15127;
															assign node15127 = (inp[7]) ? 4'b0011 : 4'b0010;
														assign node15131 = (inp[5]) ? node15133 : 4'b0000;
															assign node15133 = (inp[8]) ? node15137 : node15134;
																assign node15134 = (inp[7]) ? 4'b0001 : 4'b0000;
																assign node15137 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node15140 = (inp[15]) ? 4'b0011 : node15141;
														assign node15141 = (inp[8]) ? node15145 : node15142;
															assign node15142 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node15145 = (inp[7]) ? 4'b0000 : 4'b0001;
												assign node15149 = (inp[0]) ? node15171 : node15150;
													assign node15150 = (inp[5]) ? node15160 : node15151;
														assign node15151 = (inp[15]) ? 4'b0101 : node15152;
															assign node15152 = (inp[7]) ? node15156 : node15153;
																assign node15153 = (inp[8]) ? 4'b0111 : 4'b0110;
																assign node15156 = (inp[8]) ? 4'b0110 : 4'b0111;
														assign node15160 = (inp[15]) ? node15168 : node15161;
															assign node15161 = (inp[7]) ? node15165 : node15162;
																assign node15162 = (inp[8]) ? 4'b0101 : 4'b0100;
																assign node15165 = (inp[8]) ? 4'b0100 : 4'b0101;
															assign node15168 = (inp[8]) ? 4'b0110 : 4'b0111;
													assign node15171 = (inp[15]) ? node15183 : node15172;
														assign node15172 = (inp[5]) ? node15178 : node15173;
															assign node15173 = (inp[8]) ? node15175 : 4'b0100;
																assign node15175 = (inp[7]) ? 4'b0100 : 4'b0101;
															assign node15178 = (inp[7]) ? 4'b0110 : node15179;
																assign node15179 = (inp[8]) ? 4'b0111 : 4'b0110;
														assign node15183 = (inp[5]) ? node15185 : 4'b0110;
															assign node15185 = (inp[7]) ? node15187 : 4'b0100;
																assign node15187 = (inp[8]) ? 4'b0100 : 4'b0101;
									assign node15190 = (inp[15]) ? node15344 : node15191;
										assign node15191 = (inp[0]) ? node15263 : node15192;
											assign node15192 = (inp[4]) ? node15232 : node15193;
												assign node15193 = (inp[9]) ? node15215 : node15194;
													assign node15194 = (inp[8]) ? node15208 : node15195;
														assign node15195 = (inp[5]) ? node15201 : node15196;
															assign node15196 = (inp[7]) ? 4'b0110 : node15197;
																assign node15197 = (inp[2]) ? 4'b0110 : 4'b0111;
															assign node15201 = (inp[2]) ? node15205 : node15202;
																assign node15202 = (inp[7]) ? 4'b0110 : 4'b0111;
																assign node15205 = (inp[7]) ? 4'b0111 : 4'b0110;
														assign node15208 = (inp[7]) ? node15212 : node15209;
															assign node15209 = (inp[2]) ? 4'b0111 : 4'b0110;
															assign node15212 = (inp[2]) ? 4'b0110 : 4'b0111;
													assign node15215 = (inp[5]) ? node15225 : node15216;
														assign node15216 = (inp[7]) ? node15218 : 4'b0011;
															assign node15218 = (inp[2]) ? node15222 : node15219;
																assign node15219 = (inp[8]) ? 4'b0011 : 4'b0010;
																assign node15222 = (inp[8]) ? 4'b0010 : 4'b0011;
														assign node15225 = (inp[2]) ? 4'b0010 : node15226;
															assign node15226 = (inp[7]) ? 4'b0011 : node15227;
																assign node15227 = (inp[8]) ? 4'b0010 : 4'b0011;
												assign node15232 = (inp[9]) ? node15246 : node15233;
													assign node15233 = (inp[2]) ? node15239 : node15234;
														assign node15234 = (inp[8]) ? node15236 : 4'b0011;
															assign node15236 = (inp[7]) ? 4'b0011 : 4'b0010;
														assign node15239 = (inp[8]) ? node15243 : node15240;
															assign node15240 = (inp[7]) ? 4'b0011 : 4'b0010;
															assign node15243 = (inp[7]) ? 4'b0010 : 4'b0011;
													assign node15246 = (inp[5]) ? node15248 : 4'b0110;
														assign node15248 = (inp[2]) ? node15256 : node15249;
															assign node15249 = (inp[8]) ? node15253 : node15250;
																assign node15250 = (inp[7]) ? 4'b0100 : 4'b0101;
																assign node15253 = (inp[7]) ? 4'b0101 : 4'b0100;
															assign node15256 = (inp[8]) ? node15260 : node15257;
																assign node15257 = (inp[7]) ? 4'b0101 : 4'b0100;
																assign node15260 = (inp[7]) ? 4'b0100 : 4'b0101;
											assign node15263 = (inp[9]) ? node15301 : node15264;
												assign node15264 = (inp[4]) ? node15282 : node15265;
													assign node15265 = (inp[7]) ? node15273 : node15266;
														assign node15266 = (inp[2]) ? node15270 : node15267;
															assign node15267 = (inp[8]) ? 4'b0100 : 4'b0101;
															assign node15270 = (inp[8]) ? 4'b0101 : 4'b0100;
														assign node15273 = (inp[5]) ? node15275 : 4'b0101;
															assign node15275 = (inp[8]) ? node15279 : node15276;
																assign node15276 = (inp[2]) ? 4'b0101 : 4'b0100;
																assign node15279 = (inp[2]) ? 4'b0100 : 4'b0101;
													assign node15282 = (inp[5]) ? node15292 : node15283;
														assign node15283 = (inp[2]) ? 4'b0000 : node15284;
															assign node15284 = (inp[7]) ? node15288 : node15285;
																assign node15285 = (inp[8]) ? 4'b0000 : 4'b0001;
																assign node15288 = (inp[8]) ? 4'b0001 : 4'b0000;
														assign node15292 = (inp[8]) ? 4'b0001 : node15293;
															assign node15293 = (inp[7]) ? node15297 : node15294;
																assign node15294 = (inp[2]) ? 4'b0000 : 4'b0001;
																assign node15297 = (inp[2]) ? 4'b0001 : 4'b0000;
												assign node15301 = (inp[4]) ? node15313 : node15302;
													assign node15302 = (inp[2]) ? node15308 : node15303;
														assign node15303 = (inp[5]) ? 4'b0000 : node15304;
															assign node15304 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node15308 = (inp[7]) ? 4'b0001 : node15309;
															assign node15309 = (inp[8]) ? 4'b0001 : 4'b0000;
													assign node15313 = (inp[5]) ? node15329 : node15314;
														assign node15314 = (inp[7]) ? node15322 : node15315;
															assign node15315 = (inp[8]) ? node15319 : node15316;
																assign node15316 = (inp[2]) ? 4'b0100 : 4'b0101;
																assign node15319 = (inp[2]) ? 4'b0101 : 4'b0100;
															assign node15322 = (inp[8]) ? node15326 : node15323;
																assign node15323 = (inp[2]) ? 4'b0101 : 4'b0100;
																assign node15326 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node15329 = (inp[2]) ? node15337 : node15330;
															assign node15330 = (inp[7]) ? node15334 : node15331;
																assign node15331 = (inp[8]) ? 4'b0110 : 4'b0111;
																assign node15334 = (inp[8]) ? 4'b0111 : 4'b0110;
															assign node15337 = (inp[7]) ? node15341 : node15338;
																assign node15338 = (inp[8]) ? 4'b0111 : 4'b0110;
																assign node15341 = (inp[8]) ? 4'b0110 : 4'b0111;
										assign node15344 = (inp[0]) ? node15400 : node15345;
											assign node15345 = (inp[4]) ? node15365 : node15346;
												assign node15346 = (inp[9]) ? node15352 : node15347;
													assign node15347 = (inp[8]) ? node15349 : 4'b0100;
														assign node15349 = (inp[5]) ? 4'b0100 : 4'b0101;
													assign node15352 = (inp[8]) ? node15358 : node15353;
														assign node15353 = (inp[2]) ? node15355 : 4'b0000;
															assign node15355 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node15358 = (inp[5]) ? node15362 : node15359;
															assign node15359 = (inp[7]) ? 4'b0000 : 4'b0001;
															assign node15362 = (inp[7]) ? 4'b0001 : 4'b0000;
												assign node15365 = (inp[9]) ? node15381 : node15366;
													assign node15366 = (inp[7]) ? node15376 : node15367;
														assign node15367 = (inp[5]) ? node15373 : node15368;
															assign node15368 = (inp[8]) ? node15370 : 4'b0000;
																assign node15370 = (inp[2]) ? 4'b0001 : 4'b0000;
															assign node15373 = (inp[8]) ? 4'b0000 : 4'b0001;
														assign node15376 = (inp[5]) ? 4'b0001 : node15377;
															assign node15377 = (inp[8]) ? 4'b0001 : 4'b0000;
													assign node15381 = (inp[5]) ? node15393 : node15382;
														assign node15382 = (inp[7]) ? node15388 : node15383;
															assign node15383 = (inp[2]) ? node15385 : 4'b0100;
																assign node15385 = (inp[8]) ? 4'b0101 : 4'b0100;
															assign node15388 = (inp[2]) ? node15390 : 4'b0101;
																assign node15390 = (inp[8]) ? 4'b0100 : 4'b0101;
														assign node15393 = (inp[7]) ? 4'b0110 : node15394;
															assign node15394 = (inp[8]) ? 4'b0111 : node15395;
																assign node15395 = (inp[2]) ? 4'b0110 : 4'b0111;
											assign node15400 = (inp[5]) ? node15440 : node15401;
												assign node15401 = (inp[8]) ? node15415 : node15402;
													assign node15402 = (inp[9]) ? node15412 : node15403;
														assign node15403 = (inp[4]) ? node15409 : node15404;
															assign node15404 = (inp[2]) ? node15406 : 4'b0110;
																assign node15406 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node15409 = (inp[2]) ? 4'b0011 : 4'b0010;
														assign node15412 = (inp[4]) ? 4'b0111 : 4'b0011;
													assign node15415 = (inp[2]) ? node15431 : node15416;
														assign node15416 = (inp[7]) ? node15424 : node15417;
															assign node15417 = (inp[9]) ? node15421 : node15418;
																assign node15418 = (inp[4]) ? 4'b0010 : 4'b0110;
																assign node15421 = (inp[4]) ? 4'b0110 : 4'b0010;
															assign node15424 = (inp[9]) ? node15428 : node15425;
																assign node15425 = (inp[4]) ? 4'b0011 : 4'b0111;
																assign node15428 = (inp[4]) ? 4'b0111 : 4'b0011;
														assign node15431 = (inp[7]) ? node15433 : 4'b0111;
															assign node15433 = (inp[9]) ? node15437 : node15434;
																assign node15434 = (inp[4]) ? 4'b0010 : 4'b0110;
																assign node15437 = (inp[4]) ? 4'b0110 : 4'b0010;
												assign node15440 = (inp[4]) ? node15456 : node15441;
													assign node15441 = (inp[9]) ? node15449 : node15442;
														assign node15442 = (inp[2]) ? node15444 : 4'b0110;
															assign node15444 = (inp[7]) ? 4'b0110 : node15445;
																assign node15445 = (inp[8]) ? 4'b0111 : 4'b0110;
														assign node15449 = (inp[7]) ? node15451 : 4'b0010;
															assign node15451 = (inp[2]) ? node15453 : 4'b0010;
																assign node15453 = (inp[8]) ? 4'b0010 : 4'b0011;
													assign node15456 = (inp[9]) ? node15462 : node15457;
														assign node15457 = (inp[7]) ? 4'b0010 : node15458;
															assign node15458 = (inp[2]) ? 4'b0010 : 4'b0011;
														assign node15462 = (inp[8]) ? node15468 : node15463;
															assign node15463 = (inp[7]) ? node15465 : 4'b0100;
																assign node15465 = (inp[2]) ? 4'b0101 : 4'b0100;
															assign node15468 = (inp[7]) ? 4'b0101 : node15469;
																assign node15469 = (inp[2]) ? 4'b0101 : 4'b0100;
								assign node15473 = (inp[9]) ? node15637 : node15474;
									assign node15474 = (inp[4]) ? node15546 : node15475;
										assign node15475 = (inp[0]) ? node15499 : node15476;
											assign node15476 = (inp[15]) ? node15492 : node15477;
												assign node15477 = (inp[2]) ? node15485 : node15478;
													assign node15478 = (inp[7]) ? node15482 : node15479;
														assign node15479 = (inp[8]) ? 4'b0111 : 4'b0110;
														assign node15482 = (inp[8]) ? 4'b0110 : 4'b0111;
													assign node15485 = (inp[8]) ? node15489 : node15486;
														assign node15486 = (inp[7]) ? 4'b0111 : 4'b0110;
														assign node15489 = (inp[7]) ? 4'b0110 : 4'b0111;
												assign node15492 = (inp[8]) ? node15496 : node15493;
													assign node15493 = (inp[7]) ? 4'b0101 : 4'b0100;
													assign node15496 = (inp[7]) ? 4'b0100 : 4'b0101;
											assign node15499 = (inp[15]) ? node15515 : node15500;
												assign node15500 = (inp[12]) ? node15508 : node15501;
													assign node15501 = (inp[7]) ? node15505 : node15502;
														assign node15502 = (inp[8]) ? 4'b0101 : 4'b0100;
														assign node15505 = (inp[8]) ? 4'b0100 : 4'b0101;
													assign node15508 = (inp[7]) ? node15512 : node15509;
														assign node15509 = (inp[8]) ? 4'b0101 : 4'b0100;
														assign node15512 = (inp[8]) ? 4'b0100 : 4'b0101;
												assign node15515 = (inp[5]) ? node15529 : node15516;
													assign node15516 = (inp[2]) ? node15524 : node15517;
														assign node15517 = (inp[8]) ? node15521 : node15518;
															assign node15518 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node15521 = (inp[7]) ? 4'b0110 : 4'b0111;
														assign node15524 = (inp[8]) ? node15526 : 4'b0110;
															assign node15526 = (inp[7]) ? 4'b0110 : 4'b0111;
													assign node15529 = (inp[2]) ? node15535 : node15530;
														assign node15530 = (inp[8]) ? 4'b0110 : node15531;
															assign node15531 = (inp[7]) ? 4'b0111 : 4'b0110;
														assign node15535 = (inp[12]) ? node15541 : node15536;
															assign node15536 = (inp[8]) ? 4'b0111 : node15537;
																assign node15537 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node15541 = (inp[7]) ? node15543 : 4'b0111;
																assign node15543 = (inp[8]) ? 4'b0110 : 4'b0111;
										assign node15546 = (inp[7]) ? node15598 : node15547;
											assign node15547 = (inp[8]) ? node15581 : node15548;
												assign node15548 = (inp[5]) ? node15564 : node15549;
													assign node15549 = (inp[2]) ? node15557 : node15550;
														assign node15550 = (inp[15]) ? node15554 : node15551;
															assign node15551 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node15554 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node15557 = (inp[0]) ? node15561 : node15558;
															assign node15558 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node15561 = (inp[15]) ? 4'b0010 : 4'b0000;
													assign node15564 = (inp[12]) ? node15574 : node15565;
														assign node15565 = (inp[2]) ? node15567 : 4'b0010;
															assign node15567 = (inp[15]) ? node15571 : node15568;
																assign node15568 = (inp[0]) ? 4'b0000 : 4'b0010;
																assign node15571 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node15574 = (inp[15]) ? node15578 : node15575;
															assign node15575 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node15578 = (inp[0]) ? 4'b0010 : 4'b0000;
												assign node15581 = (inp[12]) ? node15591 : node15582;
													assign node15582 = (inp[5]) ? node15584 : 4'b0001;
														assign node15584 = (inp[0]) ? node15588 : node15585;
															assign node15585 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node15588 = (inp[15]) ? 4'b0011 : 4'b0001;
													assign node15591 = (inp[0]) ? node15595 : node15592;
														assign node15592 = (inp[15]) ? 4'b0001 : 4'b0011;
														assign node15595 = (inp[15]) ? 4'b0011 : 4'b0001;
											assign node15598 = (inp[8]) ? node15622 : node15599;
												assign node15599 = (inp[12]) ? node15615 : node15600;
													assign node15600 = (inp[2]) ? node15608 : node15601;
														assign node15601 = (inp[15]) ? node15605 : node15602;
															assign node15602 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node15605 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node15608 = (inp[0]) ? node15612 : node15609;
															assign node15609 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node15612 = (inp[15]) ? 4'b0011 : 4'b0001;
													assign node15615 = (inp[15]) ? node15619 : node15616;
														assign node15616 = (inp[0]) ? 4'b0001 : 4'b0011;
														assign node15619 = (inp[0]) ? 4'b0011 : 4'b0001;
												assign node15622 = (inp[5]) ? node15630 : node15623;
													assign node15623 = (inp[2]) ? node15625 : 4'b0010;
														assign node15625 = (inp[0]) ? node15627 : 4'b0000;
															assign node15627 = (inp[15]) ? 4'b0010 : 4'b0000;
													assign node15630 = (inp[15]) ? node15634 : node15631;
														assign node15631 = (inp[0]) ? 4'b0000 : 4'b0010;
														assign node15634 = (inp[0]) ? 4'b0010 : 4'b0000;
									assign node15637 = (inp[4]) ? node15681 : node15638;
										assign node15638 = (inp[15]) ? node15666 : node15639;
											assign node15639 = (inp[0]) ? node15647 : node15640;
												assign node15640 = (inp[8]) ? node15644 : node15641;
													assign node15641 = (inp[7]) ? 4'b0011 : 4'b0010;
													assign node15644 = (inp[7]) ? 4'b0010 : 4'b0011;
												assign node15647 = (inp[5]) ? node15659 : node15648;
													assign node15648 = (inp[2]) ? node15654 : node15649;
														assign node15649 = (inp[12]) ? 4'b0000 : node15650;
															assign node15650 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node15654 = (inp[8]) ? 4'b0001 : node15655;
															assign node15655 = (inp[7]) ? 4'b0001 : 4'b0000;
													assign node15659 = (inp[7]) ? node15663 : node15660;
														assign node15660 = (inp[8]) ? 4'b0001 : 4'b0000;
														assign node15663 = (inp[8]) ? 4'b0000 : 4'b0001;
											assign node15666 = (inp[0]) ? node15674 : node15667;
												assign node15667 = (inp[7]) ? node15671 : node15668;
													assign node15668 = (inp[8]) ? 4'b0001 : 4'b0000;
													assign node15671 = (inp[8]) ? 4'b0000 : 4'b0001;
												assign node15674 = (inp[7]) ? node15678 : node15675;
													assign node15675 = (inp[8]) ? 4'b0011 : 4'b0010;
													assign node15678 = (inp[8]) ? 4'b0010 : 4'b0011;
										assign node15681 = (inp[5]) ? node15733 : node15682;
											assign node15682 = (inp[12]) ? node15712 : node15683;
												assign node15683 = (inp[15]) ? node15699 : node15684;
													assign node15684 = (inp[0]) ? node15692 : node15685;
														assign node15685 = (inp[8]) ? node15689 : node15686;
															assign node15686 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node15689 = (inp[7]) ? 4'b0110 : 4'b0111;
														assign node15692 = (inp[8]) ? node15696 : node15693;
															assign node15693 = (inp[7]) ? 4'b0101 : 4'b0100;
															assign node15696 = (inp[7]) ? 4'b0100 : 4'b0101;
													assign node15699 = (inp[0]) ? node15705 : node15700;
														assign node15700 = (inp[7]) ? 4'b0101 : node15701;
															assign node15701 = (inp[8]) ? 4'b0101 : 4'b0100;
														assign node15705 = (inp[7]) ? node15709 : node15706;
															assign node15706 = (inp[8]) ? 4'b0111 : 4'b0110;
															assign node15709 = (inp[8]) ? 4'b0110 : 4'b0111;
												assign node15712 = (inp[8]) ? node15724 : node15713;
													assign node15713 = (inp[7]) ? node15717 : node15714;
														assign node15714 = (inp[15]) ? 4'b0100 : 4'b0110;
														assign node15717 = (inp[2]) ? 4'b0101 : node15718;
															assign node15718 = (inp[0]) ? 4'b0111 : node15719;
																assign node15719 = (inp[15]) ? 4'b0101 : 4'b0111;
													assign node15724 = (inp[7]) ? 4'b0100 : node15725;
														assign node15725 = (inp[0]) ? node15729 : node15726;
															assign node15726 = (inp[15]) ? 4'b0101 : 4'b0111;
															assign node15729 = (inp[15]) ? 4'b0111 : 4'b0101;
											assign node15733 = (inp[0]) ? node15749 : node15734;
												assign node15734 = (inp[15]) ? node15742 : node15735;
													assign node15735 = (inp[8]) ? node15739 : node15736;
														assign node15736 = (inp[7]) ? 4'b0101 : 4'b0100;
														assign node15739 = (inp[7]) ? 4'b0100 : 4'b0101;
													assign node15742 = (inp[7]) ? node15746 : node15743;
														assign node15743 = (inp[8]) ? 4'b0111 : 4'b0110;
														assign node15746 = (inp[8]) ? 4'b0110 : 4'b0111;
												assign node15749 = (inp[15]) ? node15765 : node15750;
													assign node15750 = (inp[2]) ? node15760 : node15751;
														assign node15751 = (inp[12]) ? 4'b0111 : node15752;
															assign node15752 = (inp[7]) ? node15756 : node15753;
																assign node15753 = (inp[8]) ? 4'b0111 : 4'b0110;
																assign node15756 = (inp[8]) ? 4'b0110 : 4'b0111;
														assign node15760 = (inp[7]) ? node15762 : 4'b0110;
															assign node15762 = (inp[8]) ? 4'b0110 : 4'b0111;
													assign node15765 = (inp[7]) ? node15769 : node15766;
														assign node15766 = (inp[8]) ? 4'b0101 : 4'b0100;
														assign node15769 = (inp[8]) ? 4'b0100 : 4'b0101;
							assign node15772 = (inp[4]) ? node16302 : node15773;
								assign node15773 = (inp[9]) ? node16007 : node15774;
									assign node15774 = (inp[12]) ? node15876 : node15775;
										assign node15775 = (inp[5]) ? node15821 : node15776;
											assign node15776 = (inp[15]) ? node15800 : node15777;
												assign node15777 = (inp[0]) ? node15787 : node15778;
													assign node15778 = (inp[14]) ? node15780 : 4'b0111;
														assign node15780 = (inp[8]) ? node15784 : node15781;
															assign node15781 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node15784 = (inp[7]) ? 4'b0110 : 4'b0111;
													assign node15787 = (inp[7]) ? 4'b0101 : node15788;
														assign node15788 = (inp[8]) ? node15794 : node15789;
															assign node15789 = (inp[14]) ? 4'b0100 : node15790;
																assign node15790 = (inp[2]) ? 4'b0100 : 4'b0101;
															assign node15794 = (inp[14]) ? 4'b0101 : node15795;
																assign node15795 = (inp[2]) ? 4'b0101 : 4'b0100;
												assign node15800 = (inp[0]) ? node15816 : node15801;
													assign node15801 = (inp[7]) ? node15811 : node15802;
														assign node15802 = (inp[8]) ? node15808 : node15803;
															assign node15803 = (inp[14]) ? 4'b0100 : node15804;
																assign node15804 = (inp[2]) ? 4'b0100 : 4'b0101;
															assign node15808 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node15811 = (inp[8]) ? node15813 : 4'b0101;
															assign node15813 = (inp[14]) ? 4'b0100 : 4'b0101;
													assign node15816 = (inp[8]) ? node15818 : 4'b0110;
														assign node15818 = (inp[2]) ? 4'b0110 : 4'b0111;
											assign node15821 = (inp[7]) ? node15845 : node15822;
												assign node15822 = (inp[8]) ? node15834 : node15823;
													assign node15823 = (inp[14]) ? node15831 : node15824;
														assign node15824 = (inp[2]) ? 4'b0100 : node15825;
															assign node15825 = (inp[15]) ? node15827 : 4'b0111;
																assign node15827 = (inp[0]) ? 4'b0101 : 4'b0111;
														assign node15831 = (inp[0]) ? 4'b0110 : 4'b0100;
													assign node15834 = (inp[15]) ? node15838 : node15835;
														assign node15835 = (inp[0]) ? 4'b0111 : 4'b0101;
														assign node15838 = (inp[0]) ? node15842 : node15839;
															assign node15839 = (inp[14]) ? 4'b0111 : 4'b0110;
															assign node15842 = (inp[2]) ? 4'b0101 : 4'b0100;
												assign node15845 = (inp[8]) ? node15859 : node15846;
													assign node15846 = (inp[14]) ? node15854 : node15847;
														assign node15847 = (inp[2]) ? 4'b0111 : node15848;
															assign node15848 = (inp[0]) ? 4'b0110 : node15849;
																assign node15849 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node15854 = (inp[0]) ? node15856 : 4'b0111;
															assign node15856 = (inp[15]) ? 4'b0101 : 4'b0111;
													assign node15859 = (inp[2]) ? node15869 : node15860;
														assign node15860 = (inp[14]) ? node15866 : node15861;
															assign node15861 = (inp[0]) ? 4'b0111 : node15862;
																assign node15862 = (inp[15]) ? 4'b0111 : 4'b0101;
															assign node15866 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node15869 = (inp[0]) ? node15873 : node15870;
															assign node15870 = (inp[15]) ? 4'b0110 : 4'b0100;
															assign node15873 = (inp[15]) ? 4'b0100 : 4'b0110;
										assign node15876 = (inp[5]) ? node15930 : node15877;
											assign node15877 = (inp[8]) ? node15907 : node15878;
												assign node15878 = (inp[7]) ? node15894 : node15879;
													assign node15879 = (inp[2]) ? node15887 : node15880;
														assign node15880 = (inp[14]) ? 4'b0110 : node15881;
															assign node15881 = (inp[15]) ? node15883 : 4'b0101;
																assign node15883 = (inp[0]) ? 4'b0111 : 4'b0101;
														assign node15887 = (inp[0]) ? node15891 : node15888;
															assign node15888 = (inp[15]) ? 4'b0100 : 4'b0110;
															assign node15891 = (inp[15]) ? 4'b0110 : 4'b0100;
													assign node15894 = (inp[2]) ? node15902 : node15895;
														assign node15895 = (inp[14]) ? 4'b0111 : node15896;
															assign node15896 = (inp[15]) ? 4'b0100 : node15897;
																assign node15897 = (inp[0]) ? 4'b0100 : 4'b0110;
														assign node15902 = (inp[0]) ? node15904 : 4'b0101;
															assign node15904 = (inp[15]) ? 4'b0111 : 4'b0101;
												assign node15907 = (inp[7]) ? node15915 : node15908;
													assign node15908 = (inp[15]) ? node15912 : node15909;
														assign node15909 = (inp[0]) ? 4'b0101 : 4'b0111;
														assign node15912 = (inp[0]) ? 4'b0110 : 4'b0100;
													assign node15915 = (inp[2]) ? node15923 : node15916;
														assign node15916 = (inp[14]) ? node15918 : 4'b0101;
															assign node15918 = (inp[0]) ? node15920 : 4'b0100;
																assign node15920 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node15923 = (inp[0]) ? node15927 : node15924;
															assign node15924 = (inp[15]) ? 4'b0100 : 4'b0110;
															assign node15927 = (inp[15]) ? 4'b0110 : 4'b0100;
											assign node15930 = (inp[2]) ? node15976 : node15931;
												assign node15931 = (inp[8]) ? node15955 : node15932;
													assign node15932 = (inp[15]) ? node15944 : node15933;
														assign node15933 = (inp[0]) ? node15939 : node15934;
															assign node15934 = (inp[14]) ? node15936 : 4'b0101;
																assign node15936 = (inp[7]) ? 4'b0101 : 4'b0100;
															assign node15939 = (inp[7]) ? 4'b0111 : node15940;
																assign node15940 = (inp[14]) ? 4'b0110 : 4'b0111;
														assign node15944 = (inp[0]) ? node15950 : node15945;
															assign node15945 = (inp[14]) ? node15947 : 4'b0110;
																assign node15947 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node15950 = (inp[7]) ? 4'b0100 : node15951;
																assign node15951 = (inp[14]) ? 4'b0100 : 4'b0101;
													assign node15955 = (inp[15]) ? node15965 : node15956;
														assign node15956 = (inp[0]) ? 4'b0110 : node15957;
															assign node15957 = (inp[14]) ? node15961 : node15958;
																assign node15958 = (inp[7]) ? 4'b0101 : 4'b0100;
																assign node15961 = (inp[7]) ? 4'b0100 : 4'b0101;
														assign node15965 = (inp[0]) ? node15969 : node15966;
															assign node15966 = (inp[14]) ? 4'b0111 : 4'b0110;
															assign node15969 = (inp[14]) ? node15973 : node15970;
																assign node15970 = (inp[7]) ? 4'b0101 : 4'b0100;
																assign node15973 = (inp[7]) ? 4'b0100 : 4'b0101;
												assign node15976 = (inp[8]) ? node15994 : node15977;
													assign node15977 = (inp[7]) ? node15985 : node15978;
														assign node15978 = (inp[0]) ? node15982 : node15979;
															assign node15979 = (inp[15]) ? 4'b0110 : 4'b0100;
															assign node15982 = (inp[15]) ? 4'b0100 : 4'b0110;
														assign node15985 = (inp[14]) ? 4'b0101 : node15986;
															assign node15986 = (inp[15]) ? node15990 : node15987;
																assign node15987 = (inp[0]) ? 4'b0111 : 4'b0101;
																assign node15990 = (inp[0]) ? 4'b0101 : 4'b0111;
													assign node15994 = (inp[7]) ? node16002 : node15995;
														assign node15995 = (inp[14]) ? node15997 : 4'b0111;
															assign node15997 = (inp[15]) ? 4'b0111 : node15998;
																assign node15998 = (inp[0]) ? 4'b0111 : 4'b0101;
														assign node16002 = (inp[0]) ? node16004 : 4'b0110;
															assign node16004 = (inp[15]) ? 4'b0100 : 4'b0110;
									assign node16007 = (inp[0]) ? node16167 : node16008;
										assign node16008 = (inp[2]) ? node16086 : node16009;
											assign node16009 = (inp[14]) ? node16047 : node16010;
												assign node16010 = (inp[5]) ? node16032 : node16011;
													assign node16011 = (inp[15]) ? node16019 : node16012;
														assign node16012 = (inp[7]) ? node16016 : node16013;
															assign node16013 = (inp[8]) ? 4'b0010 : 4'b0011;
															assign node16016 = (inp[8]) ? 4'b0011 : 4'b0010;
														assign node16019 = (inp[12]) ? node16025 : node16020;
															assign node16020 = (inp[7]) ? 4'b0001 : node16021;
																assign node16021 = (inp[8]) ? 4'b0000 : 4'b0001;
															assign node16025 = (inp[8]) ? node16029 : node16026;
																assign node16026 = (inp[7]) ? 4'b0000 : 4'b0001;
																assign node16029 = (inp[7]) ? 4'b0001 : 4'b0000;
													assign node16032 = (inp[15]) ? node16040 : node16033;
														assign node16033 = (inp[7]) ? node16037 : node16034;
															assign node16034 = (inp[8]) ? 4'b0000 : 4'b0001;
															assign node16037 = (inp[8]) ? 4'b0001 : 4'b0000;
														assign node16040 = (inp[8]) ? node16044 : node16041;
															assign node16041 = (inp[7]) ? 4'b0010 : 4'b0011;
															assign node16044 = (inp[7]) ? 4'b0011 : 4'b0010;
												assign node16047 = (inp[12]) ? node16065 : node16048;
													assign node16048 = (inp[8]) ? node16056 : node16049;
														assign node16049 = (inp[15]) ? node16053 : node16050;
															assign node16050 = (inp[5]) ? 4'b0000 : 4'b0010;
															assign node16053 = (inp[5]) ? 4'b0010 : 4'b0000;
														assign node16056 = (inp[7]) ? 4'b0000 : node16057;
															assign node16057 = (inp[15]) ? node16061 : node16058;
																assign node16058 = (inp[5]) ? 4'b0001 : 4'b0011;
																assign node16061 = (inp[5]) ? 4'b0011 : 4'b0001;
													assign node16065 = (inp[5]) ? node16073 : node16066;
														assign node16066 = (inp[15]) ? node16068 : 4'b0011;
															assign node16068 = (inp[8]) ? 4'b0001 : node16069;
																assign node16069 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node16073 = (inp[15]) ? node16081 : node16074;
															assign node16074 = (inp[7]) ? node16078 : node16075;
																assign node16075 = (inp[8]) ? 4'b0001 : 4'b0000;
																assign node16078 = (inp[8]) ? 4'b0000 : 4'b0001;
															assign node16081 = (inp[7]) ? node16083 : 4'b0011;
																assign node16083 = (inp[8]) ? 4'b0010 : 4'b0011;
											assign node16086 = (inp[5]) ? node16130 : node16087;
												assign node16087 = (inp[15]) ? node16109 : node16088;
													assign node16088 = (inp[12]) ? node16104 : node16089;
														assign node16089 = (inp[14]) ? node16097 : node16090;
															assign node16090 = (inp[7]) ? node16094 : node16091;
																assign node16091 = (inp[8]) ? 4'b0011 : 4'b0010;
																assign node16094 = (inp[8]) ? 4'b0010 : 4'b0011;
															assign node16097 = (inp[7]) ? node16101 : node16098;
																assign node16098 = (inp[8]) ? 4'b0011 : 4'b0010;
																assign node16101 = (inp[8]) ? 4'b0010 : 4'b0011;
														assign node16104 = (inp[7]) ? node16106 : 4'b0010;
															assign node16106 = (inp[8]) ? 4'b0010 : 4'b0011;
													assign node16109 = (inp[12]) ? node16123 : node16110;
														assign node16110 = (inp[14]) ? node16116 : node16111;
															assign node16111 = (inp[8]) ? node16113 : 4'b0000;
																assign node16113 = (inp[7]) ? 4'b0000 : 4'b0001;
															assign node16116 = (inp[8]) ? node16120 : node16117;
																assign node16117 = (inp[7]) ? 4'b0001 : 4'b0000;
																assign node16120 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node16123 = (inp[7]) ? node16127 : node16124;
															assign node16124 = (inp[8]) ? 4'b0001 : 4'b0000;
															assign node16127 = (inp[8]) ? 4'b0000 : 4'b0001;
												assign node16130 = (inp[15]) ? node16144 : node16131;
													assign node16131 = (inp[14]) ? node16133 : 4'b0001;
														assign node16133 = (inp[12]) ? node16139 : node16134;
															assign node16134 = (inp[7]) ? 4'b0001 : node16135;
																assign node16135 = (inp[8]) ? 4'b0001 : 4'b0000;
															assign node16139 = (inp[8]) ? node16141 : 4'b0000;
																assign node16141 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node16144 = (inp[12]) ? node16160 : node16145;
														assign node16145 = (inp[14]) ? node16153 : node16146;
															assign node16146 = (inp[8]) ? node16150 : node16147;
																assign node16147 = (inp[7]) ? 4'b0011 : 4'b0010;
																assign node16150 = (inp[7]) ? 4'b0010 : 4'b0011;
															assign node16153 = (inp[7]) ? node16157 : node16154;
																assign node16154 = (inp[8]) ? 4'b0011 : 4'b0010;
																assign node16157 = (inp[8]) ? 4'b0010 : 4'b0011;
														assign node16160 = (inp[7]) ? node16164 : node16161;
															assign node16161 = (inp[14]) ? 4'b0010 : 4'b0011;
															assign node16164 = (inp[8]) ? 4'b0010 : 4'b0011;
										assign node16167 = (inp[2]) ? node16251 : node16168;
											assign node16168 = (inp[12]) ? node16220 : node16169;
												assign node16169 = (inp[15]) ? node16197 : node16170;
													assign node16170 = (inp[5]) ? node16184 : node16171;
														assign node16171 = (inp[14]) ? node16179 : node16172;
															assign node16172 = (inp[7]) ? node16176 : node16173;
																assign node16173 = (inp[8]) ? 4'b0000 : 4'b0001;
																assign node16176 = (inp[8]) ? 4'b0001 : 4'b0000;
															assign node16179 = (inp[8]) ? node16181 : 4'b0000;
																assign node16181 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node16184 = (inp[8]) ? node16192 : node16185;
															assign node16185 = (inp[14]) ? node16189 : node16186;
																assign node16186 = (inp[7]) ? 4'b0010 : 4'b0011;
																assign node16189 = (inp[7]) ? 4'b0011 : 4'b0010;
															assign node16192 = (inp[14]) ? node16194 : 4'b0011;
																assign node16194 = (inp[7]) ? 4'b0010 : 4'b0011;
													assign node16197 = (inp[5]) ? node16205 : node16198;
														assign node16198 = (inp[7]) ? 4'b0011 : node16199;
															assign node16199 = (inp[8]) ? node16201 : 4'b0010;
																assign node16201 = (inp[14]) ? 4'b0011 : 4'b0010;
														assign node16205 = (inp[14]) ? node16213 : node16206;
															assign node16206 = (inp[7]) ? node16210 : node16207;
																assign node16207 = (inp[8]) ? 4'b0000 : 4'b0001;
																assign node16210 = (inp[8]) ? 4'b0001 : 4'b0000;
															assign node16213 = (inp[7]) ? node16217 : node16214;
																assign node16214 = (inp[8]) ? 4'b0001 : 4'b0000;
																assign node16217 = (inp[8]) ? 4'b0000 : 4'b0001;
												assign node16220 = (inp[7]) ? node16234 : node16221;
													assign node16221 = (inp[5]) ? node16229 : node16222;
														assign node16222 = (inp[15]) ? 4'b0011 : node16223;
															assign node16223 = (inp[8]) ? 4'b0001 : node16224;
																assign node16224 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node16229 = (inp[8]) ? node16231 : 4'b0011;
															assign node16231 = (inp[14]) ? 4'b0011 : 4'b0010;
													assign node16234 = (inp[5]) ? node16240 : node16235;
														assign node16235 = (inp[15]) ? node16237 : 4'b0000;
															assign node16237 = (inp[8]) ? 4'b0010 : 4'b0011;
														assign node16240 = (inp[15]) ? node16246 : node16241;
															assign node16241 = (inp[8]) ? 4'b0011 : node16242;
																assign node16242 = (inp[14]) ? 4'b0011 : 4'b0010;
															assign node16246 = (inp[14]) ? 4'b0000 : node16247;
																assign node16247 = (inp[8]) ? 4'b0001 : 4'b0000;
											assign node16251 = (inp[15]) ? node16265 : node16252;
												assign node16252 = (inp[5]) ? node16258 : node16253;
													assign node16253 = (inp[7]) ? node16255 : 4'b0001;
														assign node16255 = (inp[8]) ? 4'b0000 : 4'b0001;
													assign node16258 = (inp[8]) ? node16262 : node16259;
														assign node16259 = (inp[7]) ? 4'b0011 : 4'b0010;
														assign node16262 = (inp[7]) ? 4'b0010 : 4'b0011;
												assign node16265 = (inp[5]) ? node16281 : node16266;
													assign node16266 = (inp[12]) ? node16274 : node16267;
														assign node16267 = (inp[8]) ? node16271 : node16268;
															assign node16268 = (inp[7]) ? 4'b0011 : 4'b0010;
															assign node16271 = (inp[7]) ? 4'b0010 : 4'b0011;
														assign node16274 = (inp[7]) ? node16278 : node16275;
															assign node16275 = (inp[8]) ? 4'b0011 : 4'b0010;
															assign node16278 = (inp[8]) ? 4'b0010 : 4'b0011;
													assign node16281 = (inp[14]) ? node16291 : node16282;
														assign node16282 = (inp[12]) ? node16284 : 4'b0000;
															assign node16284 = (inp[7]) ? node16288 : node16285;
																assign node16285 = (inp[8]) ? 4'b0001 : 4'b0000;
																assign node16288 = (inp[8]) ? 4'b0000 : 4'b0001;
														assign node16291 = (inp[12]) ? node16297 : node16292;
															assign node16292 = (inp[7]) ? 4'b0001 : node16293;
																assign node16293 = (inp[8]) ? 4'b0001 : 4'b0000;
															assign node16297 = (inp[7]) ? node16299 : 4'b0000;
																assign node16299 = (inp[8]) ? 4'b0000 : 4'b0001;
								assign node16302 = (inp[9]) ? node16594 : node16303;
									assign node16303 = (inp[2]) ? node16457 : node16304;
										assign node16304 = (inp[8]) ? node16380 : node16305;
											assign node16305 = (inp[12]) ? node16339 : node16306;
												assign node16306 = (inp[15]) ? node16320 : node16307;
													assign node16307 = (inp[5]) ? node16317 : node16308;
														assign node16308 = (inp[0]) ? node16310 : 4'b0010;
															assign node16310 = (inp[7]) ? node16314 : node16311;
																assign node16311 = (inp[14]) ? 4'b0000 : 4'b0001;
																assign node16314 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node16317 = (inp[0]) ? 4'b0010 : 4'b0000;
													assign node16320 = (inp[0]) ? node16330 : node16321;
														assign node16321 = (inp[5]) ? node16323 : 4'b0000;
															assign node16323 = (inp[7]) ? node16327 : node16324;
																assign node16324 = (inp[14]) ? 4'b0010 : 4'b0011;
																assign node16327 = (inp[14]) ? 4'b0011 : 4'b0010;
														assign node16330 = (inp[5]) ? 4'b0000 : node16331;
															assign node16331 = (inp[7]) ? node16335 : node16332;
																assign node16332 = (inp[14]) ? 4'b0010 : 4'b0011;
																assign node16335 = (inp[14]) ? 4'b0011 : 4'b0010;
												assign node16339 = (inp[14]) ? node16363 : node16340;
													assign node16340 = (inp[7]) ? node16350 : node16341;
														assign node16341 = (inp[15]) ? 4'b0001 : node16342;
															assign node16342 = (inp[5]) ? node16346 : node16343;
																assign node16343 = (inp[0]) ? 4'b0001 : 4'b0011;
																assign node16346 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node16350 = (inp[15]) ? node16358 : node16351;
															assign node16351 = (inp[0]) ? node16355 : node16352;
																assign node16352 = (inp[5]) ? 4'b0000 : 4'b0010;
																assign node16355 = (inp[5]) ? 4'b0010 : 4'b0000;
															assign node16358 = (inp[0]) ? 4'b0010 : node16359;
																assign node16359 = (inp[5]) ? 4'b0010 : 4'b0000;
													assign node16363 = (inp[7]) ? node16369 : node16364;
														assign node16364 = (inp[0]) ? node16366 : 4'b0010;
															assign node16366 = (inp[15]) ? 4'b0000 : 4'b0010;
														assign node16369 = (inp[5]) ? node16375 : node16370;
															assign node16370 = (inp[15]) ? node16372 : 4'b0001;
																assign node16372 = (inp[0]) ? 4'b0011 : 4'b0001;
															assign node16375 = (inp[15]) ? node16377 : 4'b0011;
																assign node16377 = (inp[0]) ? 4'b0001 : 4'b0011;
											assign node16380 = (inp[15]) ? node16410 : node16381;
												assign node16381 = (inp[14]) ? node16397 : node16382;
													assign node16382 = (inp[7]) ? node16390 : node16383;
														assign node16383 = (inp[5]) ? node16387 : node16384;
															assign node16384 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node16387 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node16390 = (inp[0]) ? node16394 : node16391;
															assign node16391 = (inp[5]) ? 4'b0001 : 4'b0011;
															assign node16394 = (inp[5]) ? 4'b0011 : 4'b0001;
													assign node16397 = (inp[7]) ? node16403 : node16398;
														assign node16398 = (inp[0]) ? 4'b0001 : node16399;
															assign node16399 = (inp[12]) ? 4'b0011 : 4'b0001;
														assign node16403 = (inp[0]) ? node16407 : node16404;
															assign node16404 = (inp[5]) ? 4'b0000 : 4'b0010;
															assign node16407 = (inp[5]) ? 4'b0010 : 4'b0000;
												assign node16410 = (inp[12]) ? node16436 : node16411;
													assign node16411 = (inp[14]) ? node16423 : node16412;
														assign node16412 = (inp[7]) ? node16416 : node16413;
															assign node16413 = (inp[5]) ? 4'b0000 : 4'b0010;
															assign node16416 = (inp[5]) ? node16420 : node16417;
																assign node16417 = (inp[0]) ? 4'b0011 : 4'b0001;
																assign node16420 = (inp[0]) ? 4'b0001 : 4'b0011;
														assign node16423 = (inp[7]) ? node16429 : node16424;
															assign node16424 = (inp[0]) ? node16426 : 4'b0011;
																assign node16426 = (inp[5]) ? 4'b0001 : 4'b0011;
															assign node16429 = (inp[0]) ? node16433 : node16430;
																assign node16430 = (inp[5]) ? 4'b0010 : 4'b0000;
																assign node16433 = (inp[5]) ? 4'b0000 : 4'b0010;
													assign node16436 = (inp[7]) ? node16450 : node16437;
														assign node16437 = (inp[14]) ? node16445 : node16438;
															assign node16438 = (inp[0]) ? node16442 : node16439;
																assign node16439 = (inp[5]) ? 4'b0010 : 4'b0000;
																assign node16442 = (inp[5]) ? 4'b0000 : 4'b0010;
															assign node16445 = (inp[0]) ? 4'b0001 : node16446;
																assign node16446 = (inp[5]) ? 4'b0011 : 4'b0001;
														assign node16450 = (inp[14]) ? 4'b0000 : node16451;
															assign node16451 = (inp[0]) ? node16453 : 4'b0001;
																assign node16453 = (inp[5]) ? 4'b0001 : 4'b0011;
										assign node16457 = (inp[5]) ? node16539 : node16458;
											assign node16458 = (inp[12]) ? node16506 : node16459;
												assign node16459 = (inp[14]) ? node16481 : node16460;
													assign node16460 = (inp[15]) ? node16470 : node16461;
														assign node16461 = (inp[0]) ? node16463 : 4'b0011;
															assign node16463 = (inp[8]) ? node16467 : node16464;
																assign node16464 = (inp[7]) ? 4'b0001 : 4'b0000;
																assign node16467 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node16470 = (inp[0]) ? node16476 : node16471;
															assign node16471 = (inp[7]) ? 4'b0001 : node16472;
																assign node16472 = (inp[8]) ? 4'b0001 : 4'b0000;
															assign node16476 = (inp[8]) ? 4'b0011 : node16477;
																assign node16477 = (inp[7]) ? 4'b0011 : 4'b0010;
													assign node16481 = (inp[7]) ? node16493 : node16482;
														assign node16482 = (inp[8]) ? node16486 : node16483;
															assign node16483 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node16486 = (inp[15]) ? node16490 : node16487;
																assign node16487 = (inp[0]) ? 4'b0001 : 4'b0011;
																assign node16490 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node16493 = (inp[8]) ? node16499 : node16494;
															assign node16494 = (inp[15]) ? 4'b0001 : node16495;
																assign node16495 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node16499 = (inp[15]) ? node16503 : node16500;
																assign node16500 = (inp[0]) ? 4'b0000 : 4'b0010;
																assign node16503 = (inp[0]) ? 4'b0010 : 4'b0000;
												assign node16506 = (inp[7]) ? node16520 : node16507;
													assign node16507 = (inp[8]) ? node16515 : node16508;
														assign node16508 = (inp[14]) ? 4'b0010 : node16509;
															assign node16509 = (inp[15]) ? node16511 : 4'b0000;
																assign node16511 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node16515 = (inp[15]) ? 4'b0011 : node16516;
															assign node16516 = (inp[0]) ? 4'b0001 : 4'b0011;
													assign node16520 = (inp[8]) ? node16532 : node16521;
														assign node16521 = (inp[14]) ? node16527 : node16522;
															assign node16522 = (inp[15]) ? node16524 : 4'b0011;
																assign node16524 = (inp[0]) ? 4'b0011 : 4'b0001;
															assign node16527 = (inp[0]) ? node16529 : 4'b0001;
																assign node16529 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node16532 = (inp[15]) ? node16536 : node16533;
															assign node16533 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node16536 = (inp[0]) ? 4'b0010 : 4'b0000;
											assign node16539 = (inp[15]) ? node16561 : node16540;
												assign node16540 = (inp[0]) ? node16548 : node16541;
													assign node16541 = (inp[14]) ? node16543 : 4'b0000;
														assign node16543 = (inp[12]) ? node16545 : 4'b0001;
															assign node16545 = (inp[7]) ? 4'b0001 : 4'b0000;
													assign node16548 = (inp[12]) ? node16554 : node16549;
														assign node16549 = (inp[7]) ? node16551 : 4'b0010;
															assign node16551 = (inp[8]) ? 4'b0010 : 4'b0011;
														assign node16554 = (inp[8]) ? node16558 : node16555;
															assign node16555 = (inp[7]) ? 4'b0011 : 4'b0010;
															assign node16558 = (inp[7]) ? 4'b0010 : 4'b0011;
												assign node16561 = (inp[0]) ? node16581 : node16562;
													assign node16562 = (inp[14]) ? node16572 : node16563;
														assign node16563 = (inp[12]) ? 4'b0010 : node16564;
															assign node16564 = (inp[8]) ? node16568 : node16565;
																assign node16565 = (inp[7]) ? 4'b0011 : 4'b0010;
																assign node16568 = (inp[7]) ? 4'b0010 : 4'b0011;
														assign node16572 = (inp[12]) ? 4'b0011 : node16573;
															assign node16573 = (inp[8]) ? node16577 : node16574;
																assign node16574 = (inp[7]) ? 4'b0011 : 4'b0010;
																assign node16577 = (inp[7]) ? 4'b0010 : 4'b0011;
													assign node16581 = (inp[12]) ? node16587 : node16582;
														assign node16582 = (inp[7]) ? 4'b0000 : node16583;
															assign node16583 = (inp[8]) ? 4'b0001 : 4'b0000;
														assign node16587 = (inp[8]) ? node16591 : node16588;
															assign node16588 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node16591 = (inp[7]) ? 4'b0000 : 4'b0001;
									assign node16594 = (inp[7]) ? node16662 : node16595;
										assign node16595 = (inp[8]) ? node16635 : node16596;
											assign node16596 = (inp[14]) ? node16620 : node16597;
												assign node16597 = (inp[2]) ? node16613 : node16598;
													assign node16598 = (inp[5]) ? node16606 : node16599;
														assign node16599 = (inp[15]) ? node16603 : node16600;
															assign node16600 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node16603 = (inp[0]) ? 4'b0101 : 4'b0111;
														assign node16606 = (inp[15]) ? node16610 : node16607;
															assign node16607 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node16610 = (inp[12]) ? 4'b0101 : 4'b0111;
													assign node16613 = (inp[0]) ? node16617 : node16614;
														assign node16614 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node16617 = (inp[15]) ? 4'b0100 : 4'b0110;
												assign node16620 = (inp[2]) ? node16628 : node16621;
													assign node16621 = (inp[15]) ? node16625 : node16622;
														assign node16622 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node16625 = (inp[0]) ? 4'b0100 : 4'b0110;
													assign node16628 = (inp[15]) ? node16632 : node16629;
														assign node16629 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node16632 = (inp[0]) ? 4'b0100 : 4'b0110;
											assign node16635 = (inp[2]) ? node16655 : node16636;
												assign node16636 = (inp[14]) ? node16644 : node16637;
													assign node16637 = (inp[0]) ? node16641 : node16638;
														assign node16638 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node16641 = (inp[15]) ? 4'b0100 : 4'b0110;
													assign node16644 = (inp[5]) ? node16650 : node16645;
														assign node16645 = (inp[15]) ? 4'b0101 : node16646;
															assign node16646 = (inp[0]) ? 4'b0111 : 4'b0101;
														assign node16650 = (inp[0]) ? 4'b0101 : node16651;
															assign node16651 = (inp[15]) ? 4'b0111 : 4'b0101;
												assign node16655 = (inp[0]) ? node16659 : node16656;
													assign node16656 = (inp[15]) ? 4'b0111 : 4'b0101;
													assign node16659 = (inp[15]) ? 4'b0101 : 4'b0111;
										assign node16662 = (inp[8]) ? node16696 : node16663;
											assign node16663 = (inp[14]) ? node16677 : node16664;
												assign node16664 = (inp[2]) ? node16672 : node16665;
													assign node16665 = (inp[15]) ? node16669 : node16666;
														assign node16666 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node16669 = (inp[0]) ? 4'b0100 : 4'b0110;
													assign node16672 = (inp[0]) ? 4'b0111 : node16673;
														assign node16673 = (inp[15]) ? 4'b0111 : 4'b0101;
												assign node16677 = (inp[2]) ? node16687 : node16678;
													assign node16678 = (inp[5]) ? node16680 : 4'b0111;
														assign node16680 = (inp[15]) ? node16684 : node16681;
															assign node16681 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node16684 = (inp[0]) ? 4'b0101 : 4'b0111;
													assign node16687 = (inp[5]) ? node16693 : node16688;
														assign node16688 = (inp[15]) ? node16690 : 4'b0101;
															assign node16690 = (inp[0]) ? 4'b0101 : 4'b0111;
														assign node16693 = (inp[15]) ? 4'b0101 : 4'b0111;
											assign node16696 = (inp[14]) ? node16714 : node16697;
												assign node16697 = (inp[2]) ? node16707 : node16698;
													assign node16698 = (inp[12]) ? node16702 : node16699;
														assign node16699 = (inp[15]) ? 4'b0101 : 4'b0111;
														assign node16702 = (inp[15]) ? 4'b0111 : node16703;
															assign node16703 = (inp[0]) ? 4'b0111 : 4'b0101;
													assign node16707 = (inp[0]) ? node16711 : node16708;
														assign node16708 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node16711 = (inp[15]) ? 4'b0100 : 4'b0110;
												assign node16714 = (inp[15]) ? node16718 : node16715;
													assign node16715 = (inp[0]) ? 4'b0110 : 4'b0100;
													assign node16718 = (inp[0]) ? 4'b0100 : 4'b0110;
						assign node16721 = (inp[8]) ? node17641 : node16722;
							assign node16722 = (inp[7]) ? node17102 : node16723;
								assign node16723 = (inp[2]) ? node16929 : node16724;
									assign node16724 = (inp[14]) ? node16808 : node16725;
										assign node16725 = (inp[15]) ? node16773 : node16726;
											assign node16726 = (inp[0]) ? node16748 : node16727;
												assign node16727 = (inp[3]) ? node16739 : node16728;
													assign node16728 = (inp[5]) ? node16736 : node16729;
														assign node16729 = (inp[4]) ? node16733 : node16730;
															assign node16730 = (inp[9]) ? 4'b0011 : 4'b0111;
															assign node16733 = (inp[9]) ? 4'b0111 : 4'b0011;
														assign node16736 = (inp[9]) ? 4'b0101 : 4'b0011;
													assign node16739 = (inp[4]) ? 4'b0101 : node16740;
														assign node16740 = (inp[12]) ? node16744 : node16741;
															assign node16741 = (inp[9]) ? 4'b0011 : 4'b0111;
															assign node16744 = (inp[9]) ? 4'b0001 : 4'b0101;
												assign node16748 = (inp[3]) ? node16758 : node16749;
													assign node16749 = (inp[9]) ? node16753 : node16750;
														assign node16750 = (inp[4]) ? 4'b0001 : 4'b0101;
														assign node16753 = (inp[4]) ? node16755 : 4'b0001;
															assign node16755 = (inp[5]) ? 4'b0111 : 4'b0101;
													assign node16758 = (inp[5]) ? node16766 : node16759;
														assign node16759 = (inp[9]) ? node16763 : node16760;
															assign node16760 = (inp[4]) ? 4'b0001 : 4'b0101;
															assign node16763 = (inp[4]) ? 4'b0111 : 4'b0001;
														assign node16766 = (inp[4]) ? node16770 : node16767;
															assign node16767 = (inp[9]) ? 4'b0011 : 4'b0111;
															assign node16770 = (inp[9]) ? 4'b0111 : 4'b0011;
											assign node16773 = (inp[0]) ? node16789 : node16774;
												assign node16774 = (inp[3]) ? node16782 : node16775;
													assign node16775 = (inp[4]) ? node16779 : node16776;
														assign node16776 = (inp[9]) ? 4'b0001 : 4'b0101;
														assign node16779 = (inp[9]) ? 4'b0101 : 4'b0001;
													assign node16782 = (inp[5]) ? node16784 : 4'b0001;
														assign node16784 = (inp[9]) ? 4'b0011 : node16785;
															assign node16785 = (inp[4]) ? 4'b0011 : 4'b0111;
												assign node16789 = (inp[5]) ? node16797 : node16790;
													assign node16790 = (inp[4]) ? node16794 : node16791;
														assign node16791 = (inp[9]) ? 4'b0011 : 4'b0111;
														assign node16794 = (inp[9]) ? 4'b0111 : 4'b0011;
													assign node16797 = (inp[3]) ? node16803 : node16798;
														assign node16798 = (inp[4]) ? node16800 : 4'b0011;
															assign node16800 = (inp[9]) ? 4'b0101 : 4'b0011;
														assign node16803 = (inp[4]) ? 4'b0101 : node16804;
															assign node16804 = (inp[9]) ? 4'b0001 : 4'b0101;
										assign node16808 = (inp[5]) ? node16866 : node16809;
											assign node16809 = (inp[4]) ? node16833 : node16810;
												assign node16810 = (inp[9]) ? node16818 : node16811;
													assign node16811 = (inp[15]) ? node16815 : node16812;
														assign node16812 = (inp[0]) ? 4'b0100 : 4'b0110;
														assign node16815 = (inp[0]) ? 4'b0110 : 4'b0100;
													assign node16818 = (inp[12]) ? node16826 : node16819;
														assign node16819 = (inp[0]) ? node16823 : node16820;
															assign node16820 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node16823 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node16826 = (inp[0]) ? node16830 : node16827;
															assign node16827 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node16830 = (inp[15]) ? 4'b0010 : 4'b0000;
												assign node16833 = (inp[9]) ? node16847 : node16834;
													assign node16834 = (inp[3]) ? node16840 : node16835;
														assign node16835 = (inp[12]) ? node16837 : 4'b0000;
															assign node16837 = (inp[15]) ? 4'b0000 : 4'b0010;
														assign node16840 = (inp[15]) ? node16844 : node16841;
															assign node16841 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node16844 = (inp[0]) ? 4'b0010 : 4'b0000;
													assign node16847 = (inp[15]) ? node16853 : node16848;
														assign node16848 = (inp[0]) ? node16850 : 4'b0100;
															assign node16850 = (inp[3]) ? 4'b0110 : 4'b0100;
														assign node16853 = (inp[12]) ? node16861 : node16854;
															assign node16854 = (inp[3]) ? node16858 : node16855;
																assign node16855 = (inp[0]) ? 4'b0110 : 4'b0100;
																assign node16858 = (inp[0]) ? 4'b0100 : 4'b0110;
															assign node16861 = (inp[3]) ? node16863 : 4'b0100;
																assign node16863 = (inp[0]) ? 4'b0100 : 4'b0110;
											assign node16866 = (inp[0]) ? node16896 : node16867;
												assign node16867 = (inp[15]) ? node16887 : node16868;
													assign node16868 = (inp[3]) ? node16876 : node16869;
														assign node16869 = (inp[9]) ? node16873 : node16870;
															assign node16870 = (inp[4]) ? 4'b0010 : 4'b0110;
															assign node16873 = (inp[4]) ? 4'b0100 : 4'b0010;
														assign node16876 = (inp[12]) ? node16882 : node16877;
															assign node16877 = (inp[9]) ? 4'b0000 : node16878;
																assign node16878 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node16882 = (inp[9]) ? 4'b0100 : node16883;
																assign node16883 = (inp[4]) ? 4'b0000 : 4'b0100;
													assign node16887 = (inp[3]) ? node16889 : 4'b0000;
														assign node16889 = (inp[4]) ? node16893 : node16890;
															assign node16890 = (inp[9]) ? 4'b0010 : 4'b0110;
															assign node16893 = (inp[9]) ? 4'b0110 : 4'b0010;
												assign node16896 = (inp[15]) ? node16910 : node16897;
													assign node16897 = (inp[3]) ? node16903 : node16898;
														assign node16898 = (inp[4]) ? 4'b0110 : node16899;
															assign node16899 = (inp[9]) ? 4'b0000 : 4'b0100;
														assign node16903 = (inp[4]) ? node16907 : node16904;
															assign node16904 = (inp[9]) ? 4'b0010 : 4'b0110;
															assign node16907 = (inp[9]) ? 4'b0110 : 4'b0010;
													assign node16910 = (inp[3]) ? node16918 : node16911;
														assign node16911 = (inp[12]) ? 4'b0010 : node16912;
															assign node16912 = (inp[4]) ? 4'b0100 : node16913;
																assign node16913 = (inp[9]) ? 4'b0010 : 4'b0110;
														assign node16918 = (inp[12]) ? node16924 : node16919;
															assign node16919 = (inp[4]) ? 4'b0100 : node16920;
																assign node16920 = (inp[9]) ? 4'b0000 : 4'b0100;
															assign node16924 = (inp[9]) ? 4'b0100 : node16925;
																assign node16925 = (inp[4]) ? 4'b0000 : 4'b0100;
									assign node16929 = (inp[3]) ? node17039 : node16930;
										assign node16930 = (inp[5]) ? node17008 : node16931;
											assign node16931 = (inp[14]) ? node16971 : node16932;
												assign node16932 = (inp[9]) ? node16946 : node16933;
													assign node16933 = (inp[4]) ? node16939 : node16934;
														assign node16934 = (inp[15]) ? 4'b0110 : node16935;
															assign node16935 = (inp[0]) ? 4'b0100 : 4'b0110;
														assign node16939 = (inp[15]) ? node16943 : node16940;
															assign node16940 = (inp[12]) ? 4'b0010 : 4'b0000;
															assign node16943 = (inp[0]) ? 4'b0010 : 4'b0000;
													assign node16946 = (inp[4]) ? node16958 : node16947;
														assign node16947 = (inp[12]) ? node16953 : node16948;
															assign node16948 = (inp[15]) ? 4'b0000 : node16949;
																assign node16949 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node16953 = (inp[0]) ? 4'b0010 : node16954;
																assign node16954 = (inp[15]) ? 4'b0000 : 4'b0010;
														assign node16958 = (inp[12]) ? node16966 : node16959;
															assign node16959 = (inp[15]) ? node16963 : node16960;
																assign node16960 = (inp[0]) ? 4'b0100 : 4'b0110;
																assign node16963 = (inp[0]) ? 4'b0110 : 4'b0100;
															assign node16966 = (inp[15]) ? 4'b0100 : node16967;
																assign node16967 = (inp[0]) ? 4'b0100 : 4'b0110;
												assign node16971 = (inp[0]) ? node16985 : node16972;
													assign node16972 = (inp[15]) ? node16980 : node16973;
														assign node16973 = (inp[4]) ? node16977 : node16974;
															assign node16974 = (inp[9]) ? 4'b0010 : 4'b0110;
															assign node16977 = (inp[9]) ? 4'b0110 : 4'b0010;
														assign node16980 = (inp[9]) ? node16982 : 4'b0000;
															assign node16982 = (inp[4]) ? 4'b0100 : 4'b0000;
													assign node16985 = (inp[15]) ? node16993 : node16986;
														assign node16986 = (inp[9]) ? node16990 : node16987;
															assign node16987 = (inp[12]) ? 4'b0000 : 4'b0100;
															assign node16990 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node16993 = (inp[12]) ? node17001 : node16994;
															assign node16994 = (inp[4]) ? node16998 : node16995;
																assign node16995 = (inp[9]) ? 4'b0010 : 4'b0110;
																assign node16998 = (inp[9]) ? 4'b0110 : 4'b0010;
															assign node17001 = (inp[9]) ? node17005 : node17002;
																assign node17002 = (inp[4]) ? 4'b0010 : 4'b0110;
																assign node17005 = (inp[4]) ? 4'b0110 : 4'b0010;
											assign node17008 = (inp[0]) ? node17024 : node17009;
												assign node17009 = (inp[15]) ? node17017 : node17010;
													assign node17010 = (inp[4]) ? node17014 : node17011;
														assign node17011 = (inp[9]) ? 4'b0010 : 4'b0110;
														assign node17014 = (inp[9]) ? 4'b0100 : 4'b0010;
													assign node17017 = (inp[4]) ? node17021 : node17018;
														assign node17018 = (inp[9]) ? 4'b0000 : 4'b0100;
														assign node17021 = (inp[9]) ? 4'b0110 : 4'b0000;
												assign node17024 = (inp[15]) ? node17032 : node17025;
													assign node17025 = (inp[12]) ? 4'b0000 : node17026;
														assign node17026 = (inp[4]) ? node17028 : 4'b0000;
															assign node17028 = (inp[9]) ? 4'b0110 : 4'b0000;
													assign node17032 = (inp[4]) ? node17036 : node17033;
														assign node17033 = (inp[9]) ? 4'b0010 : 4'b0110;
														assign node17036 = (inp[9]) ? 4'b0100 : 4'b0010;
										assign node17039 = (inp[15]) ? node17071 : node17040;
											assign node17040 = (inp[0]) ? node17056 : node17041;
												assign node17041 = (inp[5]) ? node17049 : node17042;
													assign node17042 = (inp[4]) ? node17046 : node17043;
														assign node17043 = (inp[9]) ? 4'b0010 : 4'b0110;
														assign node17046 = (inp[9]) ? 4'b0100 : 4'b0010;
													assign node17049 = (inp[9]) ? node17053 : node17050;
														assign node17050 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node17053 = (inp[4]) ? 4'b0100 : 4'b0000;
												assign node17056 = (inp[5]) ? node17064 : node17057;
													assign node17057 = (inp[9]) ? node17061 : node17058;
														assign node17058 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node17061 = (inp[4]) ? 4'b0110 : 4'b0000;
													assign node17064 = (inp[4]) ? node17068 : node17065;
														assign node17065 = (inp[9]) ? 4'b0010 : 4'b0110;
														assign node17068 = (inp[9]) ? 4'b0110 : 4'b0010;
											assign node17071 = (inp[0]) ? node17087 : node17072;
												assign node17072 = (inp[5]) ? node17080 : node17073;
													assign node17073 = (inp[4]) ? node17077 : node17074;
														assign node17074 = (inp[9]) ? 4'b0000 : 4'b0100;
														assign node17077 = (inp[9]) ? 4'b0110 : 4'b0000;
													assign node17080 = (inp[4]) ? node17084 : node17081;
														assign node17081 = (inp[9]) ? 4'b0010 : 4'b0110;
														assign node17084 = (inp[9]) ? 4'b0110 : 4'b0010;
												assign node17087 = (inp[5]) ? node17095 : node17088;
													assign node17088 = (inp[4]) ? node17092 : node17089;
														assign node17089 = (inp[9]) ? 4'b0010 : 4'b0110;
														assign node17092 = (inp[9]) ? 4'b0100 : 4'b0010;
													assign node17095 = (inp[9]) ? node17099 : node17096;
														assign node17096 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node17099 = (inp[4]) ? 4'b0100 : 4'b0000;
								assign node17102 = (inp[2]) ? node17352 : node17103;
									assign node17103 = (inp[14]) ? node17217 : node17104;
										assign node17104 = (inp[0]) ? node17156 : node17105;
											assign node17105 = (inp[15]) ? node17129 : node17106;
												assign node17106 = (inp[5]) ? node17116 : node17107;
													assign node17107 = (inp[9]) ? node17111 : node17108;
														assign node17108 = (inp[4]) ? 4'b0010 : 4'b0110;
														assign node17111 = (inp[4]) ? node17113 : 4'b0010;
															assign node17113 = (inp[3]) ? 4'b0100 : 4'b0110;
													assign node17116 = (inp[3]) ? node17124 : node17117;
														assign node17117 = (inp[4]) ? node17121 : node17118;
															assign node17118 = (inp[9]) ? 4'b0010 : 4'b0110;
															assign node17121 = (inp[9]) ? 4'b0100 : 4'b0010;
														assign node17124 = (inp[9]) ? node17126 : 4'b0100;
															assign node17126 = (inp[4]) ? 4'b0100 : 4'b0000;
												assign node17129 = (inp[3]) ? node17139 : node17130;
													assign node17130 = (inp[4]) ? node17134 : node17131;
														assign node17131 = (inp[9]) ? 4'b0000 : 4'b0100;
														assign node17134 = (inp[9]) ? node17136 : 4'b0000;
															assign node17136 = (inp[5]) ? 4'b0110 : 4'b0100;
													assign node17139 = (inp[5]) ? node17147 : node17140;
														assign node17140 = (inp[4]) ? node17144 : node17141;
															assign node17141 = (inp[9]) ? 4'b0000 : 4'b0100;
															assign node17144 = (inp[9]) ? 4'b0110 : 4'b0000;
														assign node17147 = (inp[12]) ? node17149 : 4'b0110;
															assign node17149 = (inp[9]) ? node17153 : node17150;
																assign node17150 = (inp[4]) ? 4'b0010 : 4'b0110;
																assign node17153 = (inp[4]) ? 4'b0110 : 4'b0010;
											assign node17156 = (inp[15]) ? node17194 : node17157;
												assign node17157 = (inp[5]) ? node17173 : node17158;
													assign node17158 = (inp[12]) ? node17166 : node17159;
														assign node17159 = (inp[4]) ? node17163 : node17160;
															assign node17160 = (inp[9]) ? 4'b0000 : 4'b0100;
															assign node17163 = (inp[9]) ? 4'b0100 : 4'b0000;
														assign node17166 = (inp[4]) ? node17168 : 4'b0000;
															assign node17168 = (inp[9]) ? node17170 : 4'b0000;
																assign node17170 = (inp[3]) ? 4'b0110 : 4'b0100;
													assign node17173 = (inp[3]) ? node17181 : node17174;
														assign node17174 = (inp[4]) ? node17178 : node17175;
															assign node17175 = (inp[9]) ? 4'b0000 : 4'b0100;
															assign node17178 = (inp[9]) ? 4'b0110 : 4'b0000;
														assign node17181 = (inp[12]) ? node17187 : node17182;
															assign node17182 = (inp[4]) ? 4'b0010 : node17183;
																assign node17183 = (inp[9]) ? 4'b0010 : 4'b0110;
															assign node17187 = (inp[9]) ? node17191 : node17188;
																assign node17188 = (inp[4]) ? 4'b0010 : 4'b0110;
																assign node17191 = (inp[4]) ? 4'b0110 : 4'b0010;
												assign node17194 = (inp[3]) ? node17204 : node17195;
													assign node17195 = (inp[4]) ? node17199 : node17196;
														assign node17196 = (inp[9]) ? 4'b0010 : 4'b0110;
														assign node17199 = (inp[9]) ? node17201 : 4'b0010;
															assign node17201 = (inp[5]) ? 4'b0100 : 4'b0110;
													assign node17204 = (inp[5]) ? node17212 : node17205;
														assign node17205 = (inp[9]) ? node17209 : node17206;
															assign node17206 = (inp[4]) ? 4'b0010 : 4'b0110;
															assign node17209 = (inp[4]) ? 4'b0100 : 4'b0010;
														assign node17212 = (inp[4]) ? 4'b0000 : node17213;
															assign node17213 = (inp[9]) ? 4'b0000 : 4'b0100;
										assign node17217 = (inp[0]) ? node17297 : node17218;
											assign node17218 = (inp[5]) ? node17256 : node17219;
												assign node17219 = (inp[15]) ? node17237 : node17220;
													assign node17220 = (inp[3]) ? node17228 : node17221;
														assign node17221 = (inp[12]) ? node17223 : 4'b1011;
															assign node17223 = (inp[4]) ? 4'b1111 : node17224;
																assign node17224 = (inp[9]) ? 4'b1111 : 4'b1011;
														assign node17228 = (inp[12]) ? 4'b1101 : node17229;
															assign node17229 = (inp[9]) ? node17233 : node17230;
																assign node17230 = (inp[4]) ? 4'b1011 : 4'b1111;
																assign node17233 = (inp[4]) ? 4'b1101 : 4'b1011;
													assign node17237 = (inp[3]) ? node17251 : node17238;
														assign node17238 = (inp[9]) ? node17246 : node17239;
															assign node17239 = (inp[12]) ? node17243 : node17240;
																assign node17240 = (inp[4]) ? 4'b1001 : 4'b1101;
																assign node17243 = (inp[4]) ? 4'b1101 : 4'b1001;
															assign node17246 = (inp[4]) ? 4'b1101 : node17247;
																assign node17247 = (inp[12]) ? 4'b1101 : 4'b1001;
														assign node17251 = (inp[9]) ? 4'b1001 : node17252;
															assign node17252 = (inp[4]) ? 4'b1001 : 4'b1101;
												assign node17256 = (inp[15]) ? node17280 : node17257;
													assign node17257 = (inp[3]) ? node17273 : node17258;
														assign node17258 = (inp[4]) ? node17266 : node17259;
															assign node17259 = (inp[9]) ? node17263 : node17260;
																assign node17260 = (inp[12]) ? 4'b1011 : 4'b1111;
																assign node17263 = (inp[12]) ? 4'b1101 : 4'b1011;
															assign node17266 = (inp[12]) ? node17270 : node17267;
																assign node17267 = (inp[9]) ? 4'b1101 : 4'b1011;
																assign node17270 = (inp[9]) ? 4'b1001 : 4'b1101;
														assign node17273 = (inp[9]) ? node17275 : 4'b1001;
															assign node17275 = (inp[4]) ? 4'b1001 : node17276;
																assign node17276 = (inp[12]) ? 4'b1101 : 4'b1001;
													assign node17280 = (inp[3]) ? node17290 : node17281;
														assign node17281 = (inp[9]) ? 4'b1111 : node17282;
															assign node17282 = (inp[4]) ? node17286 : node17283;
																assign node17283 = (inp[12]) ? 4'b1001 : 4'b1101;
																assign node17286 = (inp[12]) ? 4'b1111 : 4'b1001;
														assign node17290 = (inp[9]) ? node17292 : 4'b1111;
															assign node17292 = (inp[12]) ? 4'b1011 : node17293;
																assign node17293 = (inp[4]) ? 4'b1111 : 4'b1011;
											assign node17297 = (inp[4]) ? node17327 : node17298;
												assign node17298 = (inp[15]) ? node17310 : node17299;
													assign node17299 = (inp[12]) ? node17303 : node17300;
														assign node17300 = (inp[9]) ? 4'b1001 : 4'b1101;
														assign node17303 = (inp[9]) ? 4'b1111 : node17304;
															assign node17304 = (inp[5]) ? node17306 : 4'b1001;
																assign node17306 = (inp[3]) ? 4'b1011 : 4'b1001;
													assign node17310 = (inp[3]) ? node17320 : node17311;
														assign node17311 = (inp[5]) ? 4'b1111 : node17312;
															assign node17312 = (inp[12]) ? node17316 : node17313;
																assign node17313 = (inp[9]) ? 4'b1011 : 4'b1111;
																assign node17316 = (inp[9]) ? 4'b1111 : 4'b1011;
														assign node17320 = (inp[5]) ? node17322 : 4'b1111;
															assign node17322 = (inp[12]) ? node17324 : 4'b1101;
																assign node17324 = (inp[9]) ? 4'b1101 : 4'b1001;
												assign node17327 = (inp[5]) ? node17337 : node17328;
													assign node17328 = (inp[15]) ? node17330 : 4'b1001;
														assign node17330 = (inp[3]) ? node17332 : 4'b1011;
															assign node17332 = (inp[12]) ? node17334 : 4'b1011;
																assign node17334 = (inp[9]) ? 4'b1001 : 4'b1101;
													assign node17337 = (inp[15]) ? node17345 : node17338;
														assign node17338 = (inp[12]) ? node17342 : node17339;
															assign node17339 = (inp[3]) ? 4'b1011 : 4'b1001;
															assign node17342 = (inp[9]) ? 4'b1011 : 4'b1111;
														assign node17345 = (inp[9]) ? node17349 : node17346;
															assign node17346 = (inp[3]) ? 4'b1001 : 4'b1011;
															assign node17349 = (inp[12]) ? 4'b1001 : 4'b1101;
									assign node17352 = (inp[5]) ? node17502 : node17353;
										assign node17353 = (inp[14]) ? node17433 : node17354;
											assign node17354 = (inp[0]) ? node17396 : node17355;
												assign node17355 = (inp[15]) ? node17377 : node17356;
													assign node17356 = (inp[3]) ? node17368 : node17357;
														assign node17357 = (inp[9]) ? node17363 : node17358;
															assign node17358 = (inp[4]) ? node17360 : 4'b1111;
																assign node17360 = (inp[12]) ? 4'b1111 : 4'b1011;
															assign node17363 = (inp[12]) ? 4'b1011 : node17364;
																assign node17364 = (inp[4]) ? 4'b1111 : 4'b1011;
														assign node17368 = (inp[9]) ? node17370 : 4'b1011;
															assign node17370 = (inp[4]) ? node17374 : node17371;
																assign node17371 = (inp[12]) ? 4'b1101 : 4'b1011;
																assign node17374 = (inp[12]) ? 4'b1001 : 4'b1101;
													assign node17377 = (inp[3]) ? node17387 : node17378;
														assign node17378 = (inp[9]) ? 4'b1101 : node17379;
															assign node17379 = (inp[12]) ? node17383 : node17380;
																assign node17380 = (inp[4]) ? 4'b1001 : 4'b1101;
																assign node17383 = (inp[4]) ? 4'b1101 : 4'b1001;
														assign node17387 = (inp[12]) ? node17389 : 4'b1001;
															assign node17389 = (inp[4]) ? node17393 : node17390;
																assign node17390 = (inp[9]) ? 4'b1111 : 4'b1001;
																assign node17393 = (inp[9]) ? 4'b1011 : 4'b1111;
												assign node17396 = (inp[15]) ? node17420 : node17397;
													assign node17397 = (inp[3]) ? node17409 : node17398;
														assign node17398 = (inp[9]) ? node17404 : node17399;
															assign node17399 = (inp[4]) ? node17401 : 4'b1001;
																assign node17401 = (inp[12]) ? 4'b1101 : 4'b1001;
															assign node17404 = (inp[4]) ? 4'b1101 : node17405;
																assign node17405 = (inp[12]) ? 4'b1101 : 4'b1001;
														assign node17409 = (inp[9]) ? node17413 : node17410;
															assign node17410 = (inp[4]) ? 4'b1001 : 4'b1101;
															assign node17413 = (inp[12]) ? node17417 : node17414;
																assign node17414 = (inp[4]) ? 4'b1111 : 4'b1001;
																assign node17417 = (inp[4]) ? 4'b1011 : 4'b1111;
													assign node17420 = (inp[4]) ? node17426 : node17421;
														assign node17421 = (inp[9]) ? 4'b1011 : node17422;
															assign node17422 = (inp[12]) ? 4'b1011 : 4'b1111;
														assign node17426 = (inp[3]) ? node17428 : 4'b1011;
															assign node17428 = (inp[9]) ? node17430 : 4'b1101;
																assign node17430 = (inp[12]) ? 4'b1001 : 4'b1101;
											assign node17433 = (inp[0]) ? node17475 : node17434;
												assign node17434 = (inp[15]) ? node17454 : node17435;
													assign node17435 = (inp[3]) ? node17445 : node17436;
														assign node17436 = (inp[9]) ? 4'b1011 : node17437;
															assign node17437 = (inp[4]) ? node17441 : node17438;
																assign node17438 = (inp[12]) ? 4'b1011 : 4'b1111;
																assign node17441 = (inp[12]) ? 4'b1111 : 4'b1011;
														assign node17445 = (inp[12]) ? node17447 : 4'b1011;
															assign node17447 = (inp[4]) ? node17451 : node17448;
																assign node17448 = (inp[9]) ? 4'b1101 : 4'b1011;
																assign node17451 = (inp[9]) ? 4'b1001 : 4'b1101;
													assign node17454 = (inp[3]) ? node17464 : node17455;
														assign node17455 = (inp[12]) ? node17457 : 4'b1001;
															assign node17457 = (inp[4]) ? node17461 : node17458;
																assign node17458 = (inp[9]) ? 4'b1101 : 4'b1001;
																assign node17461 = (inp[9]) ? 4'b1001 : 4'b1101;
														assign node17464 = (inp[12]) ? node17468 : node17465;
															assign node17465 = (inp[9]) ? 4'b1001 : 4'b1101;
															assign node17468 = (inp[4]) ? node17472 : node17469;
																assign node17469 = (inp[9]) ? 4'b1111 : 4'b1001;
																assign node17472 = (inp[9]) ? 4'b1011 : 4'b1111;
												assign node17475 = (inp[15]) ? node17493 : node17476;
													assign node17476 = (inp[3]) ? node17484 : node17477;
														assign node17477 = (inp[9]) ? 4'b1001 : node17478;
															assign node17478 = (inp[4]) ? 4'b1001 : node17479;
																assign node17479 = (inp[12]) ? 4'b1001 : 4'b1101;
														assign node17484 = (inp[9]) ? node17486 : 4'b1001;
															assign node17486 = (inp[4]) ? node17490 : node17487;
																assign node17487 = (inp[12]) ? 4'b1111 : 4'b1001;
																assign node17490 = (inp[12]) ? 4'b1011 : 4'b1111;
													assign node17493 = (inp[9]) ? node17499 : node17494;
														assign node17494 = (inp[3]) ? 4'b1011 : node17495;
															assign node17495 = (inp[12]) ? 4'b1011 : 4'b1111;
														assign node17499 = (inp[3]) ? 4'b1001 : 4'b1011;
										assign node17502 = (inp[3]) ? node17578 : node17503;
											assign node17503 = (inp[15]) ? node17545 : node17504;
												assign node17504 = (inp[14]) ? node17524 : node17505;
													assign node17505 = (inp[9]) ? node17519 : node17506;
														assign node17506 = (inp[0]) ? node17514 : node17507;
															assign node17507 = (inp[4]) ? node17511 : node17508;
																assign node17508 = (inp[12]) ? 4'b1011 : 4'b1111;
																assign node17511 = (inp[12]) ? 4'b1101 : 4'b1011;
															assign node17514 = (inp[4]) ? node17516 : 4'b1001;
																assign node17516 = (inp[12]) ? 4'b1111 : 4'b1001;
														assign node17519 = (inp[4]) ? node17521 : 4'b1011;
															assign node17521 = (inp[0]) ? 4'b1011 : 4'b1001;
													assign node17524 = (inp[12]) ? node17534 : node17525;
														assign node17525 = (inp[9]) ? node17531 : node17526;
															assign node17526 = (inp[4]) ? 4'b1001 : node17527;
																assign node17527 = (inp[0]) ? 4'b1101 : 4'b1111;
															assign node17531 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node17534 = (inp[0]) ? node17538 : node17535;
															assign node17535 = (inp[4]) ? 4'b1001 : 4'b1011;
															assign node17538 = (inp[9]) ? node17542 : node17539;
																assign node17539 = (inp[4]) ? 4'b1111 : 4'b1001;
																assign node17542 = (inp[4]) ? 4'b1011 : 4'b1111;
												assign node17545 = (inp[4]) ? node17561 : node17546;
													assign node17546 = (inp[0]) ? node17554 : node17547;
														assign node17547 = (inp[12]) ? node17551 : node17548;
															assign node17548 = (inp[9]) ? 4'b1001 : 4'b1101;
															assign node17551 = (inp[9]) ? 4'b1111 : 4'b1001;
														assign node17554 = (inp[9]) ? node17558 : node17555;
															assign node17555 = (inp[12]) ? 4'b1011 : 4'b1111;
															assign node17558 = (inp[12]) ? 4'b1101 : 4'b1011;
													assign node17561 = (inp[0]) ? node17569 : node17562;
														assign node17562 = (inp[14]) ? node17564 : 4'b1111;
															assign node17564 = (inp[12]) ? node17566 : 4'b1111;
																assign node17566 = (inp[9]) ? 4'b1011 : 4'b1111;
														assign node17569 = (inp[14]) ? node17575 : node17570;
															assign node17570 = (inp[12]) ? node17572 : 4'b1101;
																assign node17572 = (inp[9]) ? 4'b1001 : 4'b1101;
															assign node17575 = (inp[12]) ? 4'b1101 : 4'b1011;
											assign node17578 = (inp[12]) ? node17612 : node17579;
												assign node17579 = (inp[4]) ? node17597 : node17580;
													assign node17580 = (inp[9]) ? node17588 : node17581;
														assign node17581 = (inp[0]) ? node17585 : node17582;
															assign node17582 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node17585 = (inp[15]) ? 4'b1101 : 4'b1111;
														assign node17588 = (inp[14]) ? node17592 : node17589;
															assign node17589 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node17592 = (inp[0]) ? 4'b1011 : node17593;
																assign node17593 = (inp[15]) ? 4'b1011 : 4'b1001;
													assign node17597 = (inp[9]) ? node17607 : node17598;
														assign node17598 = (inp[14]) ? 4'b1001 : node17599;
															assign node17599 = (inp[0]) ? node17603 : node17600;
																assign node17600 = (inp[15]) ? 4'b1011 : 4'b1001;
																assign node17603 = (inp[15]) ? 4'b1001 : 4'b1011;
														assign node17607 = (inp[15]) ? node17609 : 4'b1101;
															assign node17609 = (inp[0]) ? 4'b1101 : 4'b1111;
												assign node17612 = (inp[9]) ? node17630 : node17613;
													assign node17613 = (inp[4]) ? node17623 : node17614;
														assign node17614 = (inp[14]) ? node17618 : node17615;
															assign node17615 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node17618 = (inp[15]) ? 4'b1001 : node17619;
																assign node17619 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node17623 = (inp[15]) ? node17627 : node17624;
															assign node17624 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node17627 = (inp[0]) ? 4'b1101 : 4'b1111;
													assign node17630 = (inp[4]) ? node17638 : node17631;
														assign node17631 = (inp[15]) ? node17635 : node17632;
															assign node17632 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node17635 = (inp[0]) ? 4'b1101 : 4'b1111;
														assign node17638 = (inp[15]) ? 4'b1011 : 4'b1001;
							assign node17641 = (inp[7]) ? node18093 : node17642;
								assign node17642 = (inp[2]) ? node17884 : node17643;
									assign node17643 = (inp[14]) ? node17753 : node17644;
										assign node17644 = (inp[5]) ? node17694 : node17645;
											assign node17645 = (inp[9]) ? node17667 : node17646;
												assign node17646 = (inp[4]) ? node17656 : node17647;
													assign node17647 = (inp[12]) ? node17649 : 4'b0110;
														assign node17649 = (inp[0]) ? node17653 : node17650;
															assign node17650 = (inp[15]) ? 4'b0100 : 4'b0110;
															assign node17653 = (inp[15]) ? 4'b0110 : 4'b0100;
													assign node17656 = (inp[12]) ? node17662 : node17657;
														assign node17657 = (inp[15]) ? 4'b0010 : node17658;
															assign node17658 = (inp[0]) ? 4'b0000 : 4'b0010;
														assign node17662 = (inp[15]) ? node17664 : 4'b0010;
															assign node17664 = (inp[0]) ? 4'b0010 : 4'b0000;
												assign node17667 = (inp[4]) ? node17679 : node17668;
													assign node17668 = (inp[3]) ? node17674 : node17669;
														assign node17669 = (inp[0]) ? 4'b0010 : node17670;
															assign node17670 = (inp[15]) ? 4'b0000 : 4'b0010;
														assign node17674 = (inp[0]) ? 4'b0000 : node17675;
															assign node17675 = (inp[15]) ? 4'b0000 : 4'b0010;
													assign node17679 = (inp[0]) ? node17687 : node17680;
														assign node17680 = (inp[3]) ? node17684 : node17681;
															assign node17681 = (inp[15]) ? 4'b0100 : 4'b0110;
															assign node17684 = (inp[12]) ? 4'b0110 : 4'b0100;
														assign node17687 = (inp[12]) ? node17689 : 4'b0110;
															assign node17689 = (inp[15]) ? 4'b0110 : node17690;
																assign node17690 = (inp[3]) ? 4'b0110 : 4'b0100;
											assign node17694 = (inp[15]) ? node17724 : node17695;
												assign node17695 = (inp[3]) ? node17713 : node17696;
													assign node17696 = (inp[12]) ? node17708 : node17697;
														assign node17697 = (inp[4]) ? node17701 : node17698;
															assign node17698 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node17701 = (inp[9]) ? node17705 : node17702;
																assign node17702 = (inp[0]) ? 4'b0000 : 4'b0010;
																assign node17705 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node17708 = (inp[4]) ? 4'b0000 : node17709;
															assign node17709 = (inp[9]) ? 4'b0000 : 4'b0100;
													assign node17713 = (inp[0]) ? node17717 : node17714;
														assign node17714 = (inp[9]) ? 4'b0100 : 4'b0000;
														assign node17717 = (inp[12]) ? node17719 : 4'b0010;
															assign node17719 = (inp[9]) ? 4'b0010 : node17720;
																assign node17720 = (inp[4]) ? 4'b0010 : 4'b0110;
												assign node17724 = (inp[3]) ? node17738 : node17725;
													assign node17725 = (inp[0]) ? node17733 : node17726;
														assign node17726 = (inp[4]) ? node17730 : node17727;
															assign node17727 = (inp[9]) ? 4'b0000 : 4'b0100;
															assign node17730 = (inp[9]) ? 4'b0110 : 4'b0000;
														assign node17733 = (inp[4]) ? 4'b0010 : node17734;
															assign node17734 = (inp[9]) ? 4'b0010 : 4'b0110;
													assign node17738 = (inp[0]) ? node17746 : node17739;
														assign node17739 = (inp[12]) ? 4'b0110 : node17740;
															assign node17740 = (inp[4]) ? 4'b0010 : node17741;
																assign node17741 = (inp[9]) ? 4'b0010 : 4'b0110;
														assign node17746 = (inp[9]) ? node17750 : node17747;
															assign node17747 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node17750 = (inp[4]) ? 4'b0100 : 4'b0000;
										assign node17753 = (inp[0]) ? node17835 : node17754;
											assign node17754 = (inp[5]) ? node17796 : node17755;
												assign node17755 = (inp[15]) ? node17781 : node17756;
													assign node17756 = (inp[3]) ? node17768 : node17757;
														assign node17757 = (inp[12]) ? node17763 : node17758;
															assign node17758 = (inp[9]) ? 4'b1111 : node17759;
																assign node17759 = (inp[4]) ? 4'b1011 : 4'b1111;
															assign node17763 = (inp[9]) ? 4'b1011 : node17764;
																assign node17764 = (inp[4]) ? 4'b1111 : 4'b1011;
														assign node17768 = (inp[4]) ? node17774 : node17769;
															assign node17769 = (inp[9]) ? 4'b1011 : node17770;
																assign node17770 = (inp[12]) ? 4'b1011 : 4'b1111;
															assign node17774 = (inp[9]) ? node17778 : node17775;
																assign node17775 = (inp[12]) ? 4'b1101 : 4'b1011;
																assign node17778 = (inp[12]) ? 4'b1001 : 4'b1101;
													assign node17781 = (inp[9]) ? node17789 : node17782;
														assign node17782 = (inp[3]) ? node17784 : 4'b1101;
															assign node17784 = (inp[12]) ? 4'b1001 : node17785;
																assign node17785 = (inp[4]) ? 4'b1001 : 4'b1101;
														assign node17789 = (inp[3]) ? node17791 : 4'b1101;
															assign node17791 = (inp[4]) ? 4'b1111 : node17792;
																assign node17792 = (inp[12]) ? 4'b1111 : 4'b1001;
												assign node17796 = (inp[15]) ? node17814 : node17797;
													assign node17797 = (inp[3]) ? node17809 : node17798;
														assign node17798 = (inp[4]) ? node17804 : node17799;
															assign node17799 = (inp[12]) ? 4'b1011 : node17800;
																assign node17800 = (inp[9]) ? 4'b1011 : 4'b1111;
															assign node17804 = (inp[12]) ? node17806 : 4'b1011;
																assign node17806 = (inp[9]) ? 4'b1001 : 4'b1101;
														assign node17809 = (inp[9]) ? 4'b1001 : node17810;
															assign node17810 = (inp[12]) ? 4'b1001 : 4'b1101;
													assign node17814 = (inp[3]) ? node17824 : node17815;
														assign node17815 = (inp[12]) ? node17817 : 4'b1001;
															assign node17817 = (inp[9]) ? node17821 : node17818;
																assign node17818 = (inp[4]) ? 4'b1111 : 4'b1001;
																assign node17821 = (inp[4]) ? 4'b1011 : 4'b1111;
														assign node17824 = (inp[12]) ? node17830 : node17825;
															assign node17825 = (inp[9]) ? 4'b1111 : node17826;
																assign node17826 = (inp[4]) ? 4'b1011 : 4'b1111;
															assign node17830 = (inp[9]) ? 4'b1011 : node17831;
																assign node17831 = (inp[4]) ? 4'b1111 : 4'b1011;
											assign node17835 = (inp[12]) ? node17851 : node17836;
												assign node17836 = (inp[15]) ? node17844 : node17837;
													assign node17837 = (inp[9]) ? node17841 : node17838;
														assign node17838 = (inp[4]) ? 4'b1001 : 4'b1101;
														assign node17841 = (inp[4]) ? 4'b1111 : 4'b1001;
													assign node17844 = (inp[5]) ? node17846 : 4'b1111;
														assign node17846 = (inp[9]) ? 4'b1101 : node17847;
															assign node17847 = (inp[3]) ? 4'b1001 : 4'b1011;
												assign node17851 = (inp[15]) ? node17871 : node17852;
													assign node17852 = (inp[3]) ? node17864 : node17853;
														assign node17853 = (inp[5]) ? node17857 : node17854;
															assign node17854 = (inp[4]) ? 4'b1101 : 4'b1001;
															assign node17857 = (inp[4]) ? node17861 : node17858;
																assign node17858 = (inp[9]) ? 4'b1111 : 4'b1001;
																assign node17861 = (inp[9]) ? 4'b1011 : 4'b1111;
														assign node17864 = (inp[9]) ? node17868 : node17865;
															assign node17865 = (inp[4]) ? 4'b1111 : 4'b1011;
															assign node17868 = (inp[4]) ? 4'b1011 : 4'b1111;
													assign node17871 = (inp[5]) ? node17879 : node17872;
														assign node17872 = (inp[9]) ? 4'b1011 : node17873;
															assign node17873 = (inp[4]) ? node17875 : 4'b1011;
																assign node17875 = (inp[3]) ? 4'b1101 : 4'b1111;
														assign node17879 = (inp[4]) ? node17881 : 4'b1101;
															assign node17881 = (inp[9]) ? 4'b1001 : 4'b1101;
									assign node17884 = (inp[9]) ? node17990 : node17885;
										assign node17885 = (inp[5]) ? node17925 : node17886;
											assign node17886 = (inp[12]) ? node17910 : node17887;
												assign node17887 = (inp[4]) ? node17895 : node17888;
													assign node17888 = (inp[15]) ? node17892 : node17889;
														assign node17889 = (inp[0]) ? 4'b1101 : 4'b1111;
														assign node17892 = (inp[0]) ? 4'b1111 : 4'b1101;
													assign node17895 = (inp[14]) ? node17903 : node17896;
														assign node17896 = (inp[0]) ? node17900 : node17897;
															assign node17897 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node17900 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node17903 = (inp[0]) ? node17907 : node17904;
															assign node17904 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node17907 = (inp[15]) ? 4'b1011 : 4'b1001;
												assign node17910 = (inp[4]) ? node17916 : node17911;
													assign node17911 = (inp[15]) ? node17913 : 4'b1001;
														assign node17913 = (inp[0]) ? 4'b1011 : 4'b1001;
													assign node17916 = (inp[15]) ? 4'b1101 : node17917;
														assign node17917 = (inp[3]) ? node17921 : node17918;
															assign node17918 = (inp[0]) ? 4'b1101 : 4'b1111;
															assign node17921 = (inp[0]) ? 4'b1111 : 4'b1101;
											assign node17925 = (inp[15]) ? node17959 : node17926;
												assign node17926 = (inp[14]) ? node17940 : node17927;
													assign node17927 = (inp[12]) ? node17933 : node17928;
														assign node17928 = (inp[0]) ? 4'b1001 : node17929;
															assign node17929 = (inp[3]) ? 4'b1001 : 4'b1011;
														assign node17933 = (inp[4]) ? node17937 : node17934;
															assign node17934 = (inp[3]) ? 4'b1011 : 4'b1001;
															assign node17937 = (inp[0]) ? 4'b1111 : 4'b1101;
													assign node17940 = (inp[3]) ? node17952 : node17941;
														assign node17941 = (inp[0]) ? node17947 : node17942;
															assign node17942 = (inp[12]) ? 4'b1011 : node17943;
																assign node17943 = (inp[4]) ? 4'b1011 : 4'b1111;
															assign node17947 = (inp[12]) ? node17949 : 4'b1001;
																assign node17949 = (inp[4]) ? 4'b1111 : 4'b1001;
														assign node17952 = (inp[0]) ? node17954 : 4'b1001;
															assign node17954 = (inp[12]) ? 4'b1011 : node17955;
																assign node17955 = (inp[4]) ? 4'b1011 : 4'b1111;
												assign node17959 = (inp[0]) ? node17975 : node17960;
													assign node17960 = (inp[3]) ? node17968 : node17961;
														assign node17961 = (inp[4]) ? node17965 : node17962;
															assign node17962 = (inp[12]) ? 4'b1001 : 4'b1101;
															assign node17965 = (inp[12]) ? 4'b1111 : 4'b1001;
														assign node17968 = (inp[14]) ? 4'b1111 : node17969;
															assign node17969 = (inp[4]) ? node17971 : 4'b1011;
																assign node17971 = (inp[12]) ? 4'b1111 : 4'b1011;
													assign node17975 = (inp[3]) ? node17983 : node17976;
														assign node17976 = (inp[12]) ? node17980 : node17977;
															assign node17977 = (inp[4]) ? 4'b1011 : 4'b1111;
															assign node17980 = (inp[4]) ? 4'b1101 : 4'b1011;
														assign node17983 = (inp[4]) ? node17987 : node17984;
															assign node17984 = (inp[12]) ? 4'b1001 : 4'b1101;
															assign node17987 = (inp[12]) ? 4'b1101 : 4'b1001;
										assign node17990 = (inp[0]) ? node18044 : node17991;
											assign node17991 = (inp[15]) ? node18015 : node17992;
												assign node17992 = (inp[5]) ? node18006 : node17993;
													assign node17993 = (inp[3]) ? node17999 : node17994;
														assign node17994 = (inp[12]) ? node17996 : 4'b1111;
															assign node17996 = (inp[4]) ? 4'b1011 : 4'b1111;
														assign node17999 = (inp[4]) ? node18003 : node18000;
															assign node18000 = (inp[12]) ? 4'b1101 : 4'b1011;
															assign node18003 = (inp[12]) ? 4'b1001 : 4'b1101;
													assign node18006 = (inp[4]) ? node18012 : node18007;
														assign node18007 = (inp[12]) ? 4'b1101 : node18008;
															assign node18008 = (inp[3]) ? 4'b1001 : 4'b1011;
														assign node18012 = (inp[12]) ? 4'b1001 : 4'b1101;
												assign node18015 = (inp[5]) ? node18029 : node18016;
													assign node18016 = (inp[3]) ? node18022 : node18017;
														assign node18017 = (inp[12]) ? 4'b1001 : node18018;
															assign node18018 = (inp[4]) ? 4'b1101 : 4'b1001;
														assign node18022 = (inp[12]) ? node18026 : node18023;
															assign node18023 = (inp[4]) ? 4'b1111 : 4'b1001;
															assign node18026 = (inp[4]) ? 4'b1011 : 4'b1111;
													assign node18029 = (inp[3]) ? node18031 : 4'b1111;
														assign node18031 = (inp[14]) ? node18039 : node18032;
															assign node18032 = (inp[12]) ? node18036 : node18033;
																assign node18033 = (inp[4]) ? 4'b1111 : 4'b1011;
																assign node18036 = (inp[4]) ? 4'b1011 : 4'b1111;
															assign node18039 = (inp[4]) ? node18041 : 4'b1011;
																assign node18041 = (inp[12]) ? 4'b1011 : 4'b1111;
											assign node18044 = (inp[15]) ? node18060 : node18045;
												assign node18045 = (inp[12]) ? node18057 : node18046;
													assign node18046 = (inp[4]) ? node18052 : node18047;
														assign node18047 = (inp[3]) ? node18049 : 4'b1001;
															assign node18049 = (inp[5]) ? 4'b1011 : 4'b1001;
														assign node18052 = (inp[3]) ? 4'b1111 : node18053;
															assign node18053 = (inp[5]) ? 4'b1111 : 4'b1101;
													assign node18057 = (inp[4]) ? 4'b1011 : 4'b1111;
												assign node18060 = (inp[5]) ? node18078 : node18061;
													assign node18061 = (inp[3]) ? node18071 : node18062;
														assign node18062 = (inp[14]) ? node18064 : 4'b1011;
															assign node18064 = (inp[12]) ? node18068 : node18065;
																assign node18065 = (inp[4]) ? 4'b1111 : 4'b1011;
																assign node18068 = (inp[4]) ? 4'b1011 : 4'b1111;
														assign node18071 = (inp[4]) ? node18075 : node18072;
															assign node18072 = (inp[12]) ? 4'b1101 : 4'b1011;
															assign node18075 = (inp[12]) ? 4'b1001 : 4'b1101;
													assign node18078 = (inp[3]) ? node18086 : node18079;
														assign node18079 = (inp[12]) ? node18083 : node18080;
															assign node18080 = (inp[4]) ? 4'b1101 : 4'b1011;
															assign node18083 = (inp[14]) ? 4'b1101 : 4'b1001;
														assign node18086 = (inp[12]) ? node18090 : node18087;
															assign node18087 = (inp[4]) ? 4'b1101 : 4'b1001;
															assign node18090 = (inp[4]) ? 4'b1001 : 4'b1101;
								assign node18093 = (inp[2]) ? node18379 : node18094;
									assign node18094 = (inp[14]) ? node18234 : node18095;
										assign node18095 = (inp[15]) ? node18159 : node18096;
											assign node18096 = (inp[4]) ? node18128 : node18097;
												assign node18097 = (inp[5]) ? node18109 : node18098;
													assign node18098 = (inp[0]) ? node18106 : node18099;
														assign node18099 = (inp[3]) ? node18103 : node18100;
															assign node18100 = (inp[9]) ? 4'b1111 : 4'b1011;
															assign node18103 = (inp[12]) ? 4'b1101 : 4'b1111;
														assign node18106 = (inp[9]) ? 4'b1001 : 4'b1101;
													assign node18109 = (inp[12]) ? node18117 : node18110;
														assign node18110 = (inp[9]) ? 4'b1011 : node18111;
															assign node18111 = (inp[3]) ? 4'b1111 : node18112;
																assign node18112 = (inp[0]) ? 4'b1101 : 4'b1111;
														assign node18117 = (inp[9]) ? node18125 : node18118;
															assign node18118 = (inp[3]) ? node18122 : node18119;
																assign node18119 = (inp[0]) ? 4'b1001 : 4'b1011;
																assign node18122 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node18125 = (inp[3]) ? 4'b1111 : 4'b1101;
												assign node18128 = (inp[0]) ? node18144 : node18129;
													assign node18129 = (inp[9]) ? node18135 : node18130;
														assign node18130 = (inp[12]) ? node18132 : 4'b1011;
															assign node18132 = (inp[5]) ? 4'b1101 : 4'b1111;
														assign node18135 = (inp[12]) ? node18139 : node18136;
															assign node18136 = (inp[3]) ? 4'b1101 : 4'b1111;
															assign node18139 = (inp[5]) ? 4'b1001 : node18140;
																assign node18140 = (inp[3]) ? 4'b1001 : 4'b1011;
													assign node18144 = (inp[9]) ? node18152 : node18145;
														assign node18145 = (inp[12]) ? 4'b1111 : node18146;
															assign node18146 = (inp[3]) ? node18148 : 4'b1001;
																assign node18148 = (inp[5]) ? 4'b1011 : 4'b1001;
														assign node18152 = (inp[12]) ? node18154 : 4'b1111;
															assign node18154 = (inp[5]) ? 4'b1011 : node18155;
																assign node18155 = (inp[3]) ? 4'b1011 : 4'b1001;
											assign node18159 = (inp[3]) ? node18193 : node18160;
												assign node18160 = (inp[0]) ? node18180 : node18161;
													assign node18161 = (inp[5]) ? node18169 : node18162;
														assign node18162 = (inp[12]) ? 4'b1001 : node18163;
															assign node18163 = (inp[4]) ? 4'b1101 : node18164;
																assign node18164 = (inp[9]) ? 4'b1001 : 4'b1101;
														assign node18169 = (inp[9]) ? node18175 : node18170;
															assign node18170 = (inp[12]) ? node18172 : 4'b1001;
																assign node18172 = (inp[4]) ? 4'b1111 : 4'b1001;
															assign node18175 = (inp[12]) ? node18177 : 4'b1111;
																assign node18177 = (inp[4]) ? 4'b1011 : 4'b1111;
													assign node18180 = (inp[5]) ? node18188 : node18181;
														assign node18181 = (inp[9]) ? 4'b1111 : node18182;
															assign node18182 = (inp[12]) ? node18184 : 4'b1011;
																assign node18184 = (inp[4]) ? 4'b1111 : 4'b1011;
														assign node18188 = (inp[9]) ? node18190 : 4'b1101;
															assign node18190 = (inp[4]) ? 4'b1001 : 4'b1011;
												assign node18193 = (inp[0]) ? node18209 : node18194;
													assign node18194 = (inp[5]) ? node18204 : node18195;
														assign node18195 = (inp[12]) ? 4'b1011 : node18196;
															assign node18196 = (inp[9]) ? node18200 : node18197;
																assign node18197 = (inp[4]) ? 4'b1001 : 4'b1101;
																assign node18200 = (inp[4]) ? 4'b1111 : 4'b1001;
														assign node18204 = (inp[9]) ? node18206 : 4'b1011;
															assign node18206 = (inp[12]) ? 4'b1111 : 4'b1011;
													assign node18209 = (inp[5]) ? node18219 : node18210;
														assign node18210 = (inp[9]) ? node18212 : 4'b1011;
															assign node18212 = (inp[4]) ? node18216 : node18213;
																assign node18213 = (inp[12]) ? 4'b1101 : 4'b1011;
																assign node18216 = (inp[12]) ? 4'b1001 : 4'b1101;
														assign node18219 = (inp[9]) ? node18227 : node18220;
															assign node18220 = (inp[12]) ? node18224 : node18221;
																assign node18221 = (inp[4]) ? 4'b1001 : 4'b1101;
																assign node18224 = (inp[4]) ? 4'b1101 : 4'b1001;
															assign node18227 = (inp[4]) ? node18231 : node18228;
																assign node18228 = (inp[12]) ? 4'b1101 : 4'b1001;
																assign node18231 = (inp[12]) ? 4'b1001 : 4'b1101;
										assign node18234 = (inp[9]) ? node18304 : node18235;
											assign node18235 = (inp[3]) ? node18261 : node18236;
												assign node18236 = (inp[12]) ? node18248 : node18237;
													assign node18237 = (inp[4]) ? node18239 : 4'b1110;
														assign node18239 = (inp[5]) ? 4'b1000 : node18240;
															assign node18240 = (inp[0]) ? node18244 : node18241;
																assign node18241 = (inp[15]) ? 4'b1000 : 4'b1010;
																assign node18244 = (inp[15]) ? 4'b1010 : 4'b1000;
													assign node18248 = (inp[4]) ? node18256 : node18249;
														assign node18249 = (inp[5]) ? 4'b1000 : node18250;
															assign node18250 = (inp[0]) ? 4'b1010 : node18251;
																assign node18251 = (inp[15]) ? 4'b1000 : 4'b1010;
														assign node18256 = (inp[0]) ? 4'b1110 : node18257;
															assign node18257 = (inp[5]) ? 4'b1110 : 4'b1100;
												assign node18261 = (inp[5]) ? node18285 : node18262;
													assign node18262 = (inp[0]) ? node18274 : node18263;
														assign node18263 = (inp[15]) ? node18269 : node18264;
															assign node18264 = (inp[12]) ? 4'b1100 : node18265;
																assign node18265 = (inp[4]) ? 4'b1010 : 4'b1110;
															assign node18269 = (inp[4]) ? 4'b1110 : node18270;
																assign node18270 = (inp[12]) ? 4'b1000 : 4'b1100;
														assign node18274 = (inp[4]) ? node18278 : node18275;
															assign node18275 = (inp[12]) ? 4'b1010 : 4'b1110;
															assign node18278 = (inp[12]) ? node18282 : node18279;
																assign node18279 = (inp[15]) ? 4'b1010 : 4'b1000;
																assign node18282 = (inp[15]) ? 4'b1100 : 4'b1110;
													assign node18285 = (inp[12]) ? node18295 : node18286;
														assign node18286 = (inp[4]) ? 4'b1000 : node18287;
															assign node18287 = (inp[0]) ? node18291 : node18288;
																assign node18288 = (inp[15]) ? 4'b1110 : 4'b1100;
																assign node18291 = (inp[15]) ? 4'b1100 : 4'b1110;
														assign node18295 = (inp[4]) ? 4'b1110 : node18296;
															assign node18296 = (inp[15]) ? node18300 : node18297;
																assign node18297 = (inp[0]) ? 4'b1010 : 4'b1000;
																assign node18300 = (inp[0]) ? 4'b1000 : 4'b1010;
											assign node18304 = (inp[15]) ? node18350 : node18305;
												assign node18305 = (inp[0]) ? node18331 : node18306;
													assign node18306 = (inp[3]) ? node18318 : node18307;
														assign node18307 = (inp[5]) ? node18311 : node18308;
															assign node18308 = (inp[12]) ? 4'b1110 : 4'b1010;
															assign node18311 = (inp[4]) ? node18315 : node18312;
																assign node18312 = (inp[12]) ? 4'b1100 : 4'b1010;
																assign node18315 = (inp[12]) ? 4'b1000 : 4'b1100;
														assign node18318 = (inp[5]) ? node18324 : node18319;
															assign node18319 = (inp[12]) ? node18321 : 4'b1100;
																assign node18321 = (inp[4]) ? 4'b1000 : 4'b1100;
															assign node18324 = (inp[12]) ? node18328 : node18325;
																assign node18325 = (inp[4]) ? 4'b1100 : 4'b1000;
																assign node18328 = (inp[4]) ? 4'b1000 : 4'b1100;
													assign node18331 = (inp[5]) ? node18343 : node18332;
														assign node18332 = (inp[3]) ? node18340 : node18333;
															assign node18333 = (inp[4]) ? node18337 : node18334;
																assign node18334 = (inp[12]) ? 4'b1100 : 4'b1000;
																assign node18337 = (inp[12]) ? 4'b1000 : 4'b1100;
															assign node18340 = (inp[12]) ? 4'b1010 : 4'b1000;
														assign node18343 = (inp[12]) ? node18347 : node18344;
															assign node18344 = (inp[4]) ? 4'b1110 : 4'b1000;
															assign node18347 = (inp[4]) ? 4'b1010 : 4'b1110;
												assign node18350 = (inp[0]) ? node18366 : node18351;
													assign node18351 = (inp[3]) ? node18357 : node18352;
														assign node18352 = (inp[12]) ? node18354 : 4'b1000;
															assign node18354 = (inp[5]) ? 4'b1110 : 4'b1000;
														assign node18357 = (inp[5]) ? 4'b1010 : node18358;
															assign node18358 = (inp[4]) ? node18362 : node18359;
																assign node18359 = (inp[12]) ? 4'b1110 : 4'b1000;
																assign node18362 = (inp[12]) ? 4'b1010 : 4'b1110;
													assign node18366 = (inp[4]) ? node18372 : node18367;
														assign node18367 = (inp[12]) ? node18369 : 4'b1010;
															assign node18369 = (inp[3]) ? 4'b1100 : 4'b1110;
														assign node18372 = (inp[12]) ? 4'b1000 : node18373;
															assign node18373 = (inp[3]) ? 4'b1100 : node18374;
																assign node18374 = (inp[5]) ? 4'b1100 : 4'b1110;
									assign node18379 = (inp[3]) ? node18525 : node18380;
										assign node18380 = (inp[5]) ? node18468 : node18381;
											assign node18381 = (inp[14]) ? node18423 : node18382;
												assign node18382 = (inp[4]) ? node18406 : node18383;
													assign node18383 = (inp[9]) ? node18393 : node18384;
														assign node18384 = (inp[12]) ? node18390 : node18385;
															assign node18385 = (inp[0]) ? 4'b1100 : node18386;
																assign node18386 = (inp[15]) ? 4'b1100 : 4'b1110;
															assign node18390 = (inp[0]) ? 4'b1000 : 4'b1010;
														assign node18393 = (inp[12]) ? node18401 : node18394;
															assign node18394 = (inp[15]) ? node18398 : node18395;
																assign node18395 = (inp[0]) ? 4'b1000 : 4'b1010;
																assign node18398 = (inp[0]) ? 4'b1010 : 4'b1000;
															assign node18401 = (inp[15]) ? node18403 : 4'b1100;
																assign node18403 = (inp[0]) ? 4'b1110 : 4'b1100;
													assign node18406 = (inp[12]) ? node18414 : node18407;
														assign node18407 = (inp[9]) ? 4'b1110 : node18408;
															assign node18408 = (inp[15]) ? node18410 : 4'b1010;
																assign node18410 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node18414 = (inp[9]) ? node18416 : 4'b1110;
															assign node18416 = (inp[15]) ? node18420 : node18417;
																assign node18417 = (inp[0]) ? 4'b1000 : 4'b1010;
																assign node18420 = (inp[0]) ? 4'b1010 : 4'b1000;
												assign node18423 = (inp[0]) ? node18445 : node18424;
													assign node18424 = (inp[15]) ? node18432 : node18425;
														assign node18425 = (inp[12]) ? 4'b1010 : node18426;
															assign node18426 = (inp[4]) ? 4'b1110 : node18427;
																assign node18427 = (inp[9]) ? 4'b1010 : 4'b1110;
														assign node18432 = (inp[9]) ? node18440 : node18433;
															assign node18433 = (inp[12]) ? node18437 : node18434;
																assign node18434 = (inp[4]) ? 4'b1000 : 4'b1100;
																assign node18437 = (inp[4]) ? 4'b1100 : 4'b1000;
															assign node18440 = (inp[4]) ? 4'b1100 : node18441;
																assign node18441 = (inp[12]) ? 4'b1100 : 4'b1000;
													assign node18445 = (inp[15]) ? node18453 : node18446;
														assign node18446 = (inp[12]) ? 4'b1100 : node18447;
															assign node18447 = (inp[9]) ? 4'b1100 : node18448;
																assign node18448 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node18453 = (inp[12]) ? node18461 : node18454;
															assign node18454 = (inp[9]) ? node18458 : node18455;
																assign node18455 = (inp[4]) ? 4'b1010 : 4'b1110;
																assign node18458 = (inp[4]) ? 4'b1110 : 4'b1010;
															assign node18461 = (inp[9]) ? node18465 : node18462;
																assign node18462 = (inp[4]) ? 4'b1110 : 4'b1010;
																assign node18465 = (inp[4]) ? 4'b1010 : 4'b1110;
											assign node18468 = (inp[15]) ? node18494 : node18469;
												assign node18469 = (inp[0]) ? node18485 : node18470;
													assign node18470 = (inp[9]) ? node18478 : node18471;
														assign node18471 = (inp[4]) ? node18475 : node18472;
															assign node18472 = (inp[12]) ? 4'b1010 : 4'b1110;
															assign node18475 = (inp[12]) ? 4'b1100 : 4'b1010;
														assign node18478 = (inp[4]) ? node18482 : node18479;
															assign node18479 = (inp[12]) ? 4'b1100 : 4'b1010;
															assign node18482 = (inp[12]) ? 4'b1000 : 4'b1100;
													assign node18485 = (inp[12]) ? 4'b1110 : node18486;
														assign node18486 = (inp[4]) ? node18490 : node18487;
															assign node18487 = (inp[9]) ? 4'b1000 : 4'b1100;
															assign node18490 = (inp[9]) ? 4'b1110 : 4'b1000;
												assign node18494 = (inp[12]) ? node18510 : node18495;
													assign node18495 = (inp[0]) ? node18503 : node18496;
														assign node18496 = (inp[4]) ? node18500 : node18497;
															assign node18497 = (inp[9]) ? 4'b1000 : 4'b1100;
															assign node18500 = (inp[9]) ? 4'b1110 : 4'b1000;
														assign node18503 = (inp[9]) ? node18507 : node18504;
															assign node18504 = (inp[4]) ? 4'b1010 : 4'b1110;
															assign node18507 = (inp[4]) ? 4'b1100 : 4'b1010;
													assign node18510 = (inp[0]) ? node18518 : node18511;
														assign node18511 = (inp[14]) ? 4'b1110 : node18512;
															assign node18512 = (inp[9]) ? node18514 : 4'b1000;
																assign node18514 = (inp[4]) ? 4'b1010 : 4'b1110;
														assign node18518 = (inp[4]) ? node18522 : node18519;
															assign node18519 = (inp[9]) ? 4'b1100 : 4'b1010;
															assign node18522 = (inp[9]) ? 4'b1000 : 4'b1100;
										assign node18525 = (inp[14]) ? node18601 : node18526;
											assign node18526 = (inp[0]) ? node18562 : node18527;
												assign node18527 = (inp[15]) ? node18543 : node18528;
													assign node18528 = (inp[5]) ? node18538 : node18529;
														assign node18529 = (inp[9]) ? node18535 : node18530;
															assign node18530 = (inp[4]) ? 4'b1010 : node18531;
																assign node18531 = (inp[12]) ? 4'b1010 : 4'b1110;
															assign node18535 = (inp[12]) ? 4'b1100 : 4'b1010;
														assign node18538 = (inp[4]) ? 4'b1000 : node18539;
															assign node18539 = (inp[12]) ? 4'b1000 : 4'b1100;
													assign node18543 = (inp[5]) ? node18553 : node18544;
														assign node18544 = (inp[4]) ? node18546 : 4'b1000;
															assign node18546 = (inp[9]) ? node18550 : node18547;
																assign node18547 = (inp[12]) ? 4'b1110 : 4'b1000;
																assign node18550 = (inp[12]) ? 4'b1010 : 4'b1110;
														assign node18553 = (inp[4]) ? 4'b1010 : node18554;
															assign node18554 = (inp[9]) ? node18558 : node18555;
																assign node18555 = (inp[12]) ? 4'b1010 : 4'b1110;
																assign node18558 = (inp[12]) ? 4'b1110 : 4'b1010;
												assign node18562 = (inp[15]) ? node18580 : node18563;
													assign node18563 = (inp[12]) ? node18571 : node18564;
														assign node18564 = (inp[9]) ? node18566 : 4'b1000;
															assign node18566 = (inp[4]) ? 4'b1110 : node18567;
																assign node18567 = (inp[5]) ? 4'b1010 : 4'b1000;
														assign node18571 = (inp[5]) ? node18575 : node18572;
															assign node18572 = (inp[4]) ? 4'b1010 : 4'b1110;
															assign node18575 = (inp[4]) ? 4'b1110 : node18576;
																assign node18576 = (inp[9]) ? 4'b1110 : 4'b1010;
													assign node18580 = (inp[5]) ? node18594 : node18581;
														assign node18581 = (inp[4]) ? node18587 : node18582;
															assign node18582 = (inp[12]) ? 4'b1010 : node18583;
																assign node18583 = (inp[9]) ? 4'b1010 : 4'b1110;
															assign node18587 = (inp[12]) ? node18591 : node18588;
																assign node18588 = (inp[9]) ? 4'b1100 : 4'b1010;
																assign node18591 = (inp[9]) ? 4'b1000 : 4'b1100;
														assign node18594 = (inp[4]) ? 4'b1100 : node18595;
															assign node18595 = (inp[9]) ? 4'b1000 : node18596;
																assign node18596 = (inp[12]) ? 4'b1000 : 4'b1100;
											assign node18601 = (inp[5]) ? node18639 : node18602;
												assign node18602 = (inp[12]) ? node18620 : node18603;
													assign node18603 = (inp[4]) ? node18613 : node18604;
														assign node18604 = (inp[9]) ? 4'b1010 : node18605;
															assign node18605 = (inp[0]) ? node18609 : node18606;
																assign node18606 = (inp[15]) ? 4'b1100 : 4'b1110;
																assign node18609 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node18613 = (inp[15]) ? node18617 : node18614;
															assign node18614 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node18617 = (inp[0]) ? 4'b1100 : 4'b1110;
													assign node18620 = (inp[15]) ? node18632 : node18621;
														assign node18621 = (inp[9]) ? node18629 : node18622;
															assign node18622 = (inp[4]) ? node18626 : node18623;
																assign node18623 = (inp[0]) ? 4'b1000 : 4'b1010;
																assign node18626 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node18629 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node18632 = (inp[0]) ? 4'b1000 : node18633;
															assign node18633 = (inp[4]) ? node18635 : 4'b1110;
																assign node18635 = (inp[9]) ? 4'b1010 : 4'b1110;
												assign node18639 = (inp[4]) ? node18651 : node18640;
													assign node18640 = (inp[15]) ? node18644 : node18641;
														assign node18641 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node18644 = (inp[0]) ? 4'b1000 : node18645;
															assign node18645 = (inp[9]) ? node18647 : 4'b1110;
																assign node18647 = (inp[12]) ? 4'b1110 : 4'b1010;
													assign node18651 = (inp[0]) ? node18665 : node18652;
														assign node18652 = (inp[15]) ? node18658 : node18653;
															assign node18653 = (inp[9]) ? node18655 : 4'b1000;
																assign node18655 = (inp[12]) ? 4'b1000 : 4'b1100;
															assign node18658 = (inp[12]) ? node18662 : node18659;
																assign node18659 = (inp[9]) ? 4'b1110 : 4'b1010;
																assign node18662 = (inp[9]) ? 4'b1010 : 4'b1110;
														assign node18665 = (inp[15]) ? 4'b1000 : 4'b1010;
					assign node18668 = (inp[13]) ? node20686 : node18669;
						assign node18669 = (inp[7]) ? node19653 : node18670;
							assign node18670 = (inp[8]) ? node19148 : node18671;
								assign node18671 = (inp[14]) ? node18889 : node18672;
									assign node18672 = (inp[2]) ? node18774 : node18673;
										assign node18673 = (inp[15]) ? node18723 : node18674;
											assign node18674 = (inp[0]) ? node18700 : node18675;
												assign node18675 = (inp[5]) ? node18685 : node18676;
													assign node18676 = (inp[9]) ? node18680 : node18677;
														assign node18677 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node18680 = (inp[4]) ? node18682 : 4'b0011;
															assign node18682 = (inp[3]) ? 4'b0101 : 4'b0111;
													assign node18685 = (inp[3]) ? node18691 : node18686;
														assign node18686 = (inp[4]) ? node18688 : 4'b0011;
															assign node18688 = (inp[9]) ? 4'b0101 : 4'b0011;
														assign node18691 = (inp[12]) ? node18693 : 4'b0101;
															assign node18693 = (inp[9]) ? node18697 : node18694;
																assign node18694 = (inp[4]) ? 4'b0001 : 4'b0101;
																assign node18697 = (inp[4]) ? 4'b0101 : 4'b0001;
												assign node18700 = (inp[5]) ? node18710 : node18701;
													assign node18701 = (inp[4]) ? node18705 : node18702;
														assign node18702 = (inp[9]) ? 4'b0001 : 4'b0101;
														assign node18705 = (inp[9]) ? node18707 : 4'b0001;
															assign node18707 = (inp[3]) ? 4'b0111 : 4'b0101;
													assign node18710 = (inp[3]) ? node18716 : node18711;
														assign node18711 = (inp[4]) ? 4'b0111 : node18712;
															assign node18712 = (inp[9]) ? 4'b0001 : 4'b0101;
														assign node18716 = (inp[9]) ? node18720 : node18717;
															assign node18717 = (inp[12]) ? 4'b0111 : 4'b0011;
															assign node18720 = (inp[4]) ? 4'b0111 : 4'b0011;
											assign node18723 = (inp[0]) ? node18749 : node18724;
												assign node18724 = (inp[3]) ? node18732 : node18725;
													assign node18725 = (inp[9]) ? node18729 : node18726;
														assign node18726 = (inp[4]) ? 4'b0001 : 4'b0101;
														assign node18729 = (inp[4]) ? 4'b0101 : 4'b0001;
													assign node18732 = (inp[5]) ? node18742 : node18733;
														assign node18733 = (inp[12]) ? node18735 : 4'b0111;
															assign node18735 = (inp[9]) ? node18739 : node18736;
																assign node18736 = (inp[4]) ? 4'b0001 : 4'b0101;
																assign node18739 = (inp[4]) ? 4'b0111 : 4'b0001;
														assign node18742 = (inp[9]) ? node18746 : node18743;
															assign node18743 = (inp[4]) ? 4'b0011 : 4'b0111;
															assign node18746 = (inp[4]) ? 4'b0111 : 4'b0011;
												assign node18749 = (inp[3]) ? node18757 : node18750;
													assign node18750 = (inp[4]) ? node18754 : node18751;
														assign node18751 = (inp[9]) ? 4'b0011 : 4'b0111;
														assign node18754 = (inp[9]) ? 4'b0111 : 4'b0011;
													assign node18757 = (inp[5]) ? node18765 : node18758;
														assign node18758 = (inp[9]) ? node18762 : node18759;
															assign node18759 = (inp[4]) ? 4'b0011 : 4'b0111;
															assign node18762 = (inp[4]) ? 4'b0101 : 4'b0011;
														assign node18765 = (inp[12]) ? node18767 : 4'b0001;
															assign node18767 = (inp[4]) ? node18771 : node18768;
																assign node18768 = (inp[9]) ? 4'b0001 : 4'b0101;
																assign node18771 = (inp[9]) ? 4'b0101 : 4'b0001;
										assign node18774 = (inp[3]) ? node18822 : node18775;
											assign node18775 = (inp[4]) ? node18799 : node18776;
												assign node18776 = (inp[9]) ? node18784 : node18777;
													assign node18777 = (inp[15]) ? node18781 : node18778;
														assign node18778 = (inp[0]) ? 4'b0100 : 4'b0110;
														assign node18781 = (inp[0]) ? 4'b0110 : 4'b0100;
													assign node18784 = (inp[12]) ? node18792 : node18785;
														assign node18785 = (inp[5]) ? 4'b0000 : node18786;
															assign node18786 = (inp[0]) ? node18788 : 4'b0000;
																assign node18788 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node18792 = (inp[15]) ? node18796 : node18793;
															assign node18793 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node18796 = (inp[0]) ? 4'b0010 : 4'b0000;
												assign node18799 = (inp[9]) ? node18807 : node18800;
													assign node18800 = (inp[15]) ? node18804 : node18801;
														assign node18801 = (inp[0]) ? 4'b0000 : 4'b0010;
														assign node18804 = (inp[0]) ? 4'b0010 : 4'b0000;
													assign node18807 = (inp[5]) ? node18815 : node18808;
														assign node18808 = (inp[15]) ? node18812 : node18809;
															assign node18809 = (inp[0]) ? 4'b0100 : 4'b0110;
															assign node18812 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node18815 = (inp[15]) ? node18819 : node18816;
															assign node18816 = (inp[0]) ? 4'b0110 : 4'b0100;
															assign node18819 = (inp[0]) ? 4'b0100 : 4'b0110;
											assign node18822 = (inp[15]) ? node18852 : node18823;
												assign node18823 = (inp[0]) ? node18837 : node18824;
													assign node18824 = (inp[5]) ? node18832 : node18825;
														assign node18825 = (inp[12]) ? 4'b0010 : node18826;
															assign node18826 = (inp[9]) ? node18828 : 4'b0010;
																assign node18828 = (inp[4]) ? 4'b0100 : 4'b0010;
														assign node18832 = (inp[9]) ? node18834 : 4'b0000;
															assign node18834 = (inp[4]) ? 4'b0100 : 4'b0000;
													assign node18837 = (inp[5]) ? node18843 : node18838;
														assign node18838 = (inp[12]) ? node18840 : 4'b0000;
															assign node18840 = (inp[4]) ? 4'b0110 : 4'b0100;
														assign node18843 = (inp[12]) ? 4'b0010 : node18844;
															assign node18844 = (inp[4]) ? node18848 : node18845;
																assign node18845 = (inp[9]) ? 4'b0010 : 4'b0110;
																assign node18848 = (inp[9]) ? 4'b0110 : 4'b0010;
												assign node18852 = (inp[12]) ? node18868 : node18853;
													assign node18853 = (inp[9]) ? node18865 : node18854;
														assign node18854 = (inp[4]) ? node18860 : node18855;
															assign node18855 = (inp[0]) ? node18857 : 4'b0110;
																assign node18857 = (inp[5]) ? 4'b0100 : 4'b0110;
															assign node18860 = (inp[5]) ? 4'b0000 : node18861;
																assign node18861 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node18865 = (inp[4]) ? 4'b0110 : 4'b0010;
													assign node18868 = (inp[9]) ? node18880 : node18869;
														assign node18869 = (inp[4]) ? node18875 : node18870;
															assign node18870 = (inp[5]) ? 4'b0110 : node18871;
																assign node18871 = (inp[0]) ? 4'b0110 : 4'b0100;
															assign node18875 = (inp[5]) ? 4'b0010 : node18876;
																assign node18876 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node18880 = (inp[4]) ? node18886 : node18881;
															assign node18881 = (inp[0]) ? node18883 : 4'b0000;
																assign node18883 = (inp[5]) ? 4'b0000 : 4'b0010;
															assign node18886 = (inp[0]) ? 4'b0100 : 4'b0110;
									assign node18889 = (inp[2]) ? node19049 : node18890;
										assign node18890 = (inp[12]) ? node18972 : node18891;
											assign node18891 = (inp[3]) ? node18931 : node18892;
												assign node18892 = (inp[0]) ? node18914 : node18893;
													assign node18893 = (inp[15]) ? node18907 : node18894;
														assign node18894 = (inp[5]) ? node18900 : node18895;
															assign node18895 = (inp[4]) ? node18897 : 4'b0010;
																assign node18897 = (inp[9]) ? 4'b0110 : 4'b0010;
															assign node18900 = (inp[4]) ? node18904 : node18901;
																assign node18901 = (inp[9]) ? 4'b0010 : 4'b0110;
																assign node18904 = (inp[9]) ? 4'b0100 : 4'b0010;
														assign node18907 = (inp[9]) ? node18911 : node18908;
															assign node18908 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node18911 = (inp[4]) ? 4'b0110 : 4'b0000;
													assign node18914 = (inp[15]) ? node18922 : node18915;
														assign node18915 = (inp[9]) ? node18919 : node18916;
															assign node18916 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node18919 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node18922 = (inp[4]) ? node18926 : node18923;
															assign node18923 = (inp[9]) ? 4'b0010 : 4'b0110;
															assign node18926 = (inp[9]) ? node18928 : 4'b0010;
																assign node18928 = (inp[5]) ? 4'b0100 : 4'b0110;
												assign node18931 = (inp[4]) ? node18957 : node18932;
													assign node18932 = (inp[9]) ? node18944 : node18933;
														assign node18933 = (inp[5]) ? node18939 : node18934;
															assign node18934 = (inp[15]) ? 4'b0110 : node18935;
																assign node18935 = (inp[0]) ? 4'b0100 : 4'b0110;
															assign node18939 = (inp[15]) ? 4'b0100 : node18940;
																assign node18940 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node18944 = (inp[5]) ? node18952 : node18945;
															assign node18945 = (inp[0]) ? node18949 : node18946;
																assign node18946 = (inp[15]) ? 4'b0000 : 4'b0010;
																assign node18949 = (inp[15]) ? 4'b0010 : 4'b0000;
															assign node18952 = (inp[0]) ? node18954 : 4'b0000;
																assign node18954 = (inp[15]) ? 4'b0000 : 4'b0010;
													assign node18957 = (inp[15]) ? node18965 : node18958;
														assign node18958 = (inp[5]) ? node18962 : node18959;
															assign node18959 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node18962 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node18965 = (inp[0]) ? node18969 : node18966;
															assign node18966 = (inp[5]) ? 4'b0010 : 4'b0000;
															assign node18969 = (inp[5]) ? 4'b0000 : 4'b0010;
											assign node18972 = (inp[0]) ? node19012 : node18973;
												assign node18973 = (inp[15]) ? node18995 : node18974;
													assign node18974 = (inp[5]) ? node18982 : node18975;
														assign node18975 = (inp[3]) ? node18977 : 4'b0110;
															assign node18977 = (inp[9]) ? 4'b0010 : node18978;
																assign node18978 = (inp[4]) ? 4'b0010 : 4'b0110;
														assign node18982 = (inp[3]) ? node18988 : node18983;
															assign node18983 = (inp[9]) ? 4'b0100 : node18984;
																assign node18984 = (inp[4]) ? 4'b0010 : 4'b0110;
															assign node18988 = (inp[9]) ? node18992 : node18989;
																assign node18989 = (inp[4]) ? 4'b0000 : 4'b0100;
																assign node18992 = (inp[4]) ? 4'b0100 : 4'b0000;
													assign node18995 = (inp[3]) ? node19007 : node18996;
														assign node18996 = (inp[5]) ? node19002 : node18997;
															assign node18997 = (inp[4]) ? node18999 : 4'b0100;
																assign node18999 = (inp[9]) ? 4'b0100 : 4'b0000;
															assign node19002 = (inp[4]) ? 4'b0110 : node19003;
																assign node19003 = (inp[9]) ? 4'b0000 : 4'b0100;
														assign node19007 = (inp[4]) ? node19009 : 4'b0110;
															assign node19009 = (inp[9]) ? 4'b0110 : 4'b0000;
												assign node19012 = (inp[15]) ? node19032 : node19013;
													assign node19013 = (inp[3]) ? node19021 : node19014;
														assign node19014 = (inp[4]) ? node19018 : node19015;
															assign node19015 = (inp[9]) ? 4'b0000 : 4'b0100;
															assign node19018 = (inp[5]) ? 4'b0110 : 4'b0100;
														assign node19021 = (inp[5]) ? node19027 : node19022;
															assign node19022 = (inp[9]) ? node19024 : 4'b0000;
																assign node19024 = (inp[4]) ? 4'b0110 : 4'b0000;
															assign node19027 = (inp[9]) ? 4'b0110 : node19028;
																assign node19028 = (inp[4]) ? 4'b0010 : 4'b0110;
													assign node19032 = (inp[5]) ? node19040 : node19033;
														assign node19033 = (inp[4]) ? node19037 : node19034;
															assign node19034 = (inp[9]) ? 4'b0010 : 4'b0110;
															assign node19037 = (inp[9]) ? 4'b0110 : 4'b0010;
														assign node19040 = (inp[3]) ? node19046 : node19041;
															assign node19041 = (inp[4]) ? 4'b0010 : node19042;
																assign node19042 = (inp[9]) ? 4'b0010 : 4'b0110;
															assign node19046 = (inp[9]) ? 4'b0000 : 4'b0100;
										assign node19049 = (inp[15]) ? node19101 : node19050;
											assign node19050 = (inp[0]) ? node19086 : node19051;
												assign node19051 = (inp[5]) ? node19073 : node19052;
													assign node19052 = (inp[3]) ? node19066 : node19053;
														assign node19053 = (inp[12]) ? node19059 : node19054;
															assign node19054 = (inp[9]) ? 4'b0110 : node19055;
																assign node19055 = (inp[4]) ? 4'b0010 : 4'b0110;
															assign node19059 = (inp[9]) ? node19063 : node19060;
																assign node19060 = (inp[4]) ? 4'b0010 : 4'b0110;
																assign node19063 = (inp[4]) ? 4'b0110 : 4'b0010;
														assign node19066 = (inp[4]) ? node19070 : node19067;
															assign node19067 = (inp[9]) ? 4'b0010 : 4'b0110;
															assign node19070 = (inp[9]) ? 4'b0100 : 4'b0010;
													assign node19073 = (inp[3]) ? node19081 : node19074;
														assign node19074 = (inp[4]) ? node19078 : node19075;
															assign node19075 = (inp[9]) ? 4'b0010 : 4'b0110;
															assign node19078 = (inp[9]) ? 4'b0100 : 4'b0010;
														assign node19081 = (inp[4]) ? node19083 : 4'b0100;
															assign node19083 = (inp[9]) ? 4'b0100 : 4'b0000;
												assign node19086 = (inp[5]) ? node19094 : node19087;
													assign node19087 = (inp[12]) ? 4'b0100 : node19088;
														assign node19088 = (inp[4]) ? 4'b0000 : node19089;
															assign node19089 = (inp[9]) ? 4'b0000 : 4'b0100;
													assign node19094 = (inp[4]) ? node19098 : node19095;
														assign node19095 = (inp[9]) ? 4'b0000 : 4'b0110;
														assign node19098 = (inp[9]) ? 4'b0110 : 4'b0010;
											assign node19101 = (inp[0]) ? node19133 : node19102;
												assign node19102 = (inp[3]) ? node19112 : node19103;
													assign node19103 = (inp[9]) ? node19107 : node19104;
														assign node19104 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node19107 = (inp[4]) ? node19109 : 4'b0000;
															assign node19109 = (inp[12]) ? 4'b0110 : 4'b0100;
													assign node19112 = (inp[5]) ? node19120 : node19113;
														assign node19113 = (inp[12]) ? node19115 : 4'b0110;
															assign node19115 = (inp[4]) ? 4'b0000 : node19116;
																assign node19116 = (inp[9]) ? 4'b0000 : 4'b0100;
														assign node19120 = (inp[12]) ? node19128 : node19121;
															assign node19121 = (inp[9]) ? node19125 : node19122;
																assign node19122 = (inp[4]) ? 4'b0010 : 4'b0110;
																assign node19125 = (inp[4]) ? 4'b0110 : 4'b0010;
															assign node19128 = (inp[4]) ? node19130 : 4'b0110;
																assign node19130 = (inp[9]) ? 4'b0110 : 4'b0010;
												assign node19133 = (inp[9]) ? node19137 : node19134;
													assign node19134 = (inp[4]) ? 4'b0010 : 4'b0110;
													assign node19137 = (inp[4]) ? node19143 : node19138;
														assign node19138 = (inp[5]) ? node19140 : 4'b0010;
															assign node19140 = (inp[3]) ? 4'b0000 : 4'b0010;
														assign node19143 = (inp[3]) ? 4'b0100 : node19144;
															assign node19144 = (inp[5]) ? 4'b0100 : 4'b0110;
								assign node19148 = (inp[2]) ? node19366 : node19149;
									assign node19149 = (inp[14]) ? node19255 : node19150;
										assign node19150 = (inp[15]) ? node19204 : node19151;
											assign node19151 = (inp[3]) ? node19171 : node19152;
												assign node19152 = (inp[0]) ? node19162 : node19153;
													assign node19153 = (inp[9]) ? node19157 : node19154;
														assign node19154 = (inp[4]) ? 4'b0010 : 4'b0110;
														assign node19157 = (inp[4]) ? node19159 : 4'b0010;
															assign node19159 = (inp[5]) ? 4'b0100 : 4'b0110;
													assign node19162 = (inp[9]) ? node19166 : node19163;
														assign node19163 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node19166 = (inp[4]) ? node19168 : 4'b0000;
															assign node19168 = (inp[5]) ? 4'b0110 : 4'b0100;
												assign node19171 = (inp[0]) ? node19185 : node19172;
													assign node19172 = (inp[5]) ? node19180 : node19173;
														assign node19173 = (inp[4]) ? node19177 : node19174;
															assign node19174 = (inp[9]) ? 4'b0010 : 4'b0110;
															assign node19177 = (inp[9]) ? 4'b0100 : 4'b0010;
														assign node19180 = (inp[4]) ? 4'b0000 : node19181;
															assign node19181 = (inp[9]) ? 4'b0000 : 4'b0100;
													assign node19185 = (inp[5]) ? node19189 : node19186;
														assign node19186 = (inp[4]) ? 4'b0110 : 4'b0100;
														assign node19189 = (inp[12]) ? node19197 : node19190;
															assign node19190 = (inp[9]) ? node19194 : node19191;
																assign node19191 = (inp[4]) ? 4'b0010 : 4'b0110;
																assign node19194 = (inp[4]) ? 4'b0110 : 4'b0010;
															assign node19197 = (inp[9]) ? node19201 : node19198;
																assign node19198 = (inp[4]) ? 4'b0010 : 4'b0110;
																assign node19201 = (inp[4]) ? 4'b0110 : 4'b0010;
											assign node19204 = (inp[0]) ? node19230 : node19205;
												assign node19205 = (inp[5]) ? node19215 : node19206;
													assign node19206 = (inp[3]) ? 4'b0000 : node19207;
														assign node19207 = (inp[9]) ? node19211 : node19208;
															assign node19208 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node19211 = (inp[4]) ? 4'b0100 : 4'b0000;
													assign node19215 = (inp[3]) ? node19223 : node19216;
														assign node19216 = (inp[12]) ? node19218 : 4'b0000;
															assign node19218 = (inp[9]) ? 4'b0110 : node19219;
																assign node19219 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node19223 = (inp[9]) ? node19227 : node19224;
															assign node19224 = (inp[4]) ? 4'b0010 : 4'b0110;
															assign node19227 = (inp[4]) ? 4'b0110 : 4'b0010;
												assign node19230 = (inp[3]) ? node19240 : node19231;
													assign node19231 = (inp[9]) ? node19235 : node19232;
														assign node19232 = (inp[4]) ? 4'b0010 : 4'b0110;
														assign node19235 = (inp[4]) ? node19237 : 4'b0010;
															assign node19237 = (inp[5]) ? 4'b0100 : 4'b0110;
													assign node19240 = (inp[5]) ? node19250 : node19241;
														assign node19241 = (inp[12]) ? node19243 : 4'b0010;
															assign node19243 = (inp[9]) ? node19247 : node19244;
																assign node19244 = (inp[4]) ? 4'b0010 : 4'b0110;
																assign node19247 = (inp[4]) ? 4'b0100 : 4'b0010;
														assign node19250 = (inp[4]) ? 4'b0000 : node19251;
															assign node19251 = (inp[9]) ? 4'b0000 : 4'b0100;
										assign node19255 = (inp[4]) ? node19307 : node19256;
											assign node19256 = (inp[9]) ? node19282 : node19257;
												assign node19257 = (inp[12]) ? node19267 : node19258;
													assign node19258 = (inp[0]) ? node19260 : 4'b1111;
														assign node19260 = (inp[3]) ? node19262 : 4'b1111;
															assign node19262 = (inp[15]) ? 4'b1101 : node19263;
																assign node19263 = (inp[5]) ? 4'b1111 : 4'b1101;
													assign node19267 = (inp[5]) ? node19275 : node19268;
														assign node19268 = (inp[0]) ? node19272 : node19269;
															assign node19269 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node19272 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node19275 = (inp[0]) ? 4'b1011 : node19276;
															assign node19276 = (inp[3]) ? 4'b1011 : node19277;
																assign node19277 = (inp[15]) ? 4'b1001 : 4'b1011;
												assign node19282 = (inp[12]) ? node19298 : node19283;
													assign node19283 = (inp[15]) ? node19293 : node19284;
														assign node19284 = (inp[5]) ? node19286 : 4'b1011;
															assign node19286 = (inp[3]) ? node19290 : node19287;
																assign node19287 = (inp[0]) ? 4'b1001 : 4'b1011;
																assign node19290 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node19293 = (inp[0]) ? node19295 : 4'b1001;
															assign node19295 = (inp[3]) ? 4'b1001 : 4'b1011;
													assign node19298 = (inp[0]) ? 4'b1101 : node19299;
														assign node19299 = (inp[5]) ? 4'b1101 : node19300;
															assign node19300 = (inp[15]) ? 4'b1111 : node19301;
																assign node19301 = (inp[3]) ? 4'b1101 : 4'b1111;
											assign node19307 = (inp[12]) ? node19335 : node19308;
												assign node19308 = (inp[9]) ? node19314 : node19309;
													assign node19309 = (inp[5]) ? 4'b1001 : node19310;
														assign node19310 = (inp[0]) ? 4'b1001 : 4'b1011;
													assign node19314 = (inp[5]) ? node19324 : node19315;
														assign node19315 = (inp[0]) ? node19317 : 4'b1111;
															assign node19317 = (inp[3]) ? node19321 : node19318;
																assign node19318 = (inp[15]) ? 4'b1111 : 4'b1101;
																assign node19321 = (inp[15]) ? 4'b1101 : 4'b1111;
														assign node19324 = (inp[3]) ? node19330 : node19325;
															assign node19325 = (inp[15]) ? 4'b1111 : node19326;
																assign node19326 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node19330 = (inp[15]) ? 4'b1101 : node19331;
																assign node19331 = (inp[0]) ? 4'b1111 : 4'b1101;
												assign node19335 = (inp[9]) ? node19351 : node19336;
													assign node19336 = (inp[15]) ? node19342 : node19337;
														assign node19337 = (inp[5]) ? node19339 : 4'b1111;
															assign node19339 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node19342 = (inp[0]) ? node19346 : node19343;
															assign node19343 = (inp[3]) ? 4'b1111 : 4'b1101;
															assign node19346 = (inp[5]) ? 4'b1101 : node19347;
																assign node19347 = (inp[3]) ? 4'b1101 : 4'b1111;
													assign node19351 = (inp[5]) ? node19361 : node19352;
														assign node19352 = (inp[15]) ? node19354 : 4'b1001;
															assign node19354 = (inp[0]) ? node19358 : node19355;
																assign node19355 = (inp[3]) ? 4'b1011 : 4'b1001;
																assign node19358 = (inp[3]) ? 4'b1001 : 4'b1011;
														assign node19361 = (inp[0]) ? node19363 : 4'b1011;
															assign node19363 = (inp[15]) ? 4'b1001 : 4'b1011;
									assign node19366 = (inp[14]) ? node19520 : node19367;
										assign node19367 = (inp[15]) ? node19441 : node19368;
											assign node19368 = (inp[4]) ? node19406 : node19369;
												assign node19369 = (inp[3]) ? node19387 : node19370;
													assign node19370 = (inp[0]) ? node19382 : node19371;
														assign node19371 = (inp[5]) ? node19379 : node19372;
															assign node19372 = (inp[12]) ? node19376 : node19373;
																assign node19373 = (inp[9]) ? 4'b1011 : 4'b1111;
																assign node19376 = (inp[9]) ? 4'b1111 : 4'b1011;
															assign node19379 = (inp[12]) ? 4'b1101 : 4'b1111;
														assign node19382 = (inp[9]) ? node19384 : 4'b1101;
															assign node19384 = (inp[12]) ? 4'b1101 : 4'b1001;
													assign node19387 = (inp[0]) ? node19397 : node19388;
														assign node19388 = (inp[5]) ? 4'b1101 : node19389;
															assign node19389 = (inp[9]) ? node19393 : node19390;
																assign node19390 = (inp[12]) ? 4'b1011 : 4'b1111;
																assign node19393 = (inp[12]) ? 4'b1101 : 4'b1011;
														assign node19397 = (inp[5]) ? node19399 : 4'b1111;
															assign node19399 = (inp[9]) ? node19403 : node19400;
																assign node19400 = (inp[12]) ? 4'b1011 : 4'b1111;
																assign node19403 = (inp[12]) ? 4'b1111 : 4'b1011;
												assign node19406 = (inp[5]) ? node19424 : node19407;
													assign node19407 = (inp[12]) ? node19417 : node19408;
														assign node19408 = (inp[9]) ? node19412 : node19409;
															assign node19409 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node19412 = (inp[0]) ? 4'b1101 : node19413;
																assign node19413 = (inp[3]) ? 4'b1101 : 4'b1111;
														assign node19417 = (inp[3]) ? node19421 : node19418;
															assign node19418 = (inp[0]) ? 4'b1101 : 4'b1111;
															assign node19421 = (inp[0]) ? 4'b1111 : 4'b1101;
													assign node19424 = (inp[0]) ? node19434 : node19425;
														assign node19425 = (inp[3]) ? node19429 : node19426;
															assign node19426 = (inp[12]) ? 4'b1001 : 4'b1011;
															assign node19429 = (inp[12]) ? 4'b1001 : node19430;
																assign node19430 = (inp[9]) ? 4'b1101 : 4'b1001;
														assign node19434 = (inp[12]) ? node19438 : node19435;
															assign node19435 = (inp[9]) ? 4'b1111 : 4'b1001;
															assign node19438 = (inp[9]) ? 4'b1011 : 4'b1111;
											assign node19441 = (inp[0]) ? node19487 : node19442;
												assign node19442 = (inp[3]) ? node19466 : node19443;
													assign node19443 = (inp[4]) ? node19457 : node19444;
														assign node19444 = (inp[5]) ? node19452 : node19445;
															assign node19445 = (inp[9]) ? node19449 : node19446;
																assign node19446 = (inp[12]) ? 4'b1001 : 4'b1101;
																assign node19449 = (inp[12]) ? 4'b1101 : 4'b1001;
															assign node19452 = (inp[9]) ? 4'b1001 : node19453;
																assign node19453 = (inp[12]) ? 4'b1001 : 4'b1101;
														assign node19457 = (inp[9]) ? node19459 : 4'b1001;
															assign node19459 = (inp[12]) ? node19463 : node19460;
																assign node19460 = (inp[5]) ? 4'b1111 : 4'b1101;
																assign node19463 = (inp[5]) ? 4'b1011 : 4'b1001;
													assign node19466 = (inp[5]) ? node19480 : node19467;
														assign node19467 = (inp[4]) ? node19473 : node19468;
															assign node19468 = (inp[12]) ? 4'b1001 : node19469;
																assign node19469 = (inp[9]) ? 4'b1001 : 4'b1101;
															assign node19473 = (inp[9]) ? node19477 : node19474;
																assign node19474 = (inp[12]) ? 4'b1111 : 4'b1001;
																assign node19477 = (inp[12]) ? 4'b1011 : 4'b1111;
														assign node19480 = (inp[12]) ? node19482 : 4'b1111;
															assign node19482 = (inp[9]) ? 4'b1011 : node19483;
																assign node19483 = (inp[4]) ? 4'b1111 : 4'b1011;
												assign node19487 = (inp[5]) ? node19503 : node19488;
													assign node19488 = (inp[3]) ? node19498 : node19489;
														assign node19489 = (inp[12]) ? node19491 : 4'b1111;
															assign node19491 = (inp[4]) ? node19495 : node19492;
																assign node19492 = (inp[9]) ? 4'b1111 : 4'b1011;
																assign node19495 = (inp[9]) ? 4'b1011 : 4'b1111;
														assign node19498 = (inp[12]) ? 4'b1101 : node19499;
															assign node19499 = (inp[9]) ? 4'b1011 : 4'b1111;
													assign node19503 = (inp[12]) ? node19515 : node19504;
														assign node19504 = (inp[3]) ? node19510 : node19505;
															assign node19505 = (inp[4]) ? node19507 : 4'b1011;
																assign node19507 = (inp[9]) ? 4'b1101 : 4'b1011;
															assign node19510 = (inp[4]) ? node19512 : 4'b1101;
																assign node19512 = (inp[9]) ? 4'b1101 : 4'b1001;
														assign node19515 = (inp[4]) ? node19517 : 4'b1101;
															assign node19517 = (inp[9]) ? 4'b1001 : 4'b1101;
										assign node19520 = (inp[15]) ? node19582 : node19521;
											assign node19521 = (inp[5]) ? node19553 : node19522;
												assign node19522 = (inp[0]) ? node19534 : node19523;
													assign node19523 = (inp[12]) ? node19527 : node19524;
														assign node19524 = (inp[3]) ? 4'b1011 : 4'b1111;
														assign node19527 = (inp[3]) ? node19529 : 4'b1011;
															assign node19529 = (inp[9]) ? node19531 : 4'b1101;
																assign node19531 = (inp[4]) ? 4'b1001 : 4'b1101;
													assign node19534 = (inp[3]) ? node19544 : node19535;
														assign node19535 = (inp[4]) ? node19537 : 4'b1001;
															assign node19537 = (inp[9]) ? node19541 : node19538;
																assign node19538 = (inp[12]) ? 4'b1101 : 4'b1001;
																assign node19541 = (inp[12]) ? 4'b1001 : 4'b1101;
														assign node19544 = (inp[9]) ? 4'b1011 : node19545;
															assign node19545 = (inp[4]) ? node19549 : node19546;
																assign node19546 = (inp[12]) ? 4'b1001 : 4'b1101;
																assign node19549 = (inp[12]) ? 4'b1111 : 4'b1001;
												assign node19553 = (inp[0]) ? node19569 : node19554;
													assign node19554 = (inp[9]) ? node19562 : node19555;
														assign node19555 = (inp[3]) ? node19557 : 4'b1011;
															assign node19557 = (inp[4]) ? 4'b1101 : node19558;
																assign node19558 = (inp[12]) ? 4'b1001 : 4'b1101;
														assign node19562 = (inp[12]) ? node19566 : node19563;
															assign node19563 = (inp[4]) ? 4'b1101 : 4'b1001;
															assign node19566 = (inp[4]) ? 4'b1001 : 4'b1101;
													assign node19569 = (inp[3]) ? node19577 : node19570;
														assign node19570 = (inp[9]) ? node19572 : 4'b1001;
															assign node19572 = (inp[12]) ? 4'b1111 : node19573;
																assign node19573 = (inp[4]) ? 4'b1111 : 4'b1001;
														assign node19577 = (inp[9]) ? 4'b1111 : node19578;
															assign node19578 = (inp[4]) ? 4'b1111 : 4'b1011;
											assign node19582 = (inp[4]) ? node19614 : node19583;
												assign node19583 = (inp[3]) ? node19597 : node19584;
													assign node19584 = (inp[12]) ? node19588 : node19585;
														assign node19585 = (inp[9]) ? 4'b1001 : 4'b1101;
														assign node19588 = (inp[9]) ? node19590 : 4'b1001;
															assign node19590 = (inp[0]) ? node19594 : node19591;
																assign node19591 = (inp[5]) ? 4'b1111 : 4'b1101;
																assign node19594 = (inp[5]) ? 4'b1101 : 4'b1111;
													assign node19597 = (inp[5]) ? node19607 : node19598;
														assign node19598 = (inp[9]) ? node19604 : node19599;
															assign node19599 = (inp[0]) ? node19601 : 4'b1101;
																assign node19601 = (inp[12]) ? 4'b1011 : 4'b1111;
															assign node19604 = (inp[12]) ? 4'b1101 : 4'b1001;
														assign node19607 = (inp[9]) ? node19611 : node19608;
															assign node19608 = (inp[12]) ? 4'b1011 : 4'b1111;
															assign node19611 = (inp[12]) ? 4'b1111 : 4'b1011;
												assign node19614 = (inp[0]) ? node19632 : node19615;
													assign node19615 = (inp[3]) ? node19623 : node19616;
														assign node19616 = (inp[12]) ? node19618 : 4'b1001;
															assign node19618 = (inp[9]) ? 4'b1001 : node19619;
																assign node19619 = (inp[5]) ? 4'b1111 : 4'b1101;
														assign node19623 = (inp[9]) ? node19629 : node19624;
															assign node19624 = (inp[12]) ? 4'b1111 : node19625;
																assign node19625 = (inp[5]) ? 4'b1011 : 4'b1001;
															assign node19629 = (inp[12]) ? 4'b1011 : 4'b1111;
													assign node19632 = (inp[5]) ? node19642 : node19633;
														assign node19633 = (inp[3]) ? node19639 : node19634;
															assign node19634 = (inp[12]) ? 4'b1011 : node19635;
																assign node19635 = (inp[9]) ? 4'b1111 : 4'b1011;
															assign node19639 = (inp[9]) ? 4'b1001 : 4'b1011;
														assign node19642 = (inp[3]) ? node19646 : node19643;
															assign node19643 = (inp[12]) ? 4'b1001 : 4'b1011;
															assign node19646 = (inp[12]) ? node19650 : node19647;
																assign node19647 = (inp[9]) ? 4'b1101 : 4'b1001;
																assign node19650 = (inp[9]) ? 4'b1001 : 4'b1101;
							assign node19653 = (inp[8]) ? node20171 : node19654;
								assign node19654 = (inp[2]) ? node19912 : node19655;
									assign node19655 = (inp[14]) ? node19775 : node19656;
										assign node19656 = (inp[15]) ? node19720 : node19657;
											assign node19657 = (inp[0]) ? node19695 : node19658;
												assign node19658 = (inp[5]) ? node19674 : node19659;
													assign node19659 = (inp[12]) ? node19665 : node19660;
														assign node19660 = (inp[9]) ? 4'b0010 : node19661;
															assign node19661 = (inp[4]) ? 4'b0010 : 4'b0110;
														assign node19665 = (inp[9]) ? node19669 : node19666;
															assign node19666 = (inp[4]) ? 4'b0010 : 4'b0110;
															assign node19669 = (inp[4]) ? node19671 : 4'b0010;
																assign node19671 = (inp[3]) ? 4'b0100 : 4'b0110;
													assign node19674 = (inp[3]) ? node19682 : node19675;
														assign node19675 = (inp[9]) ? node19679 : node19676;
															assign node19676 = (inp[4]) ? 4'b0010 : 4'b0110;
															assign node19679 = (inp[4]) ? 4'b0100 : 4'b0010;
														assign node19682 = (inp[12]) ? node19690 : node19683;
															assign node19683 = (inp[9]) ? node19687 : node19684;
																assign node19684 = (inp[4]) ? 4'b0000 : 4'b0100;
																assign node19687 = (inp[4]) ? 4'b0100 : 4'b0000;
															assign node19690 = (inp[4]) ? 4'b0100 : node19691;
																assign node19691 = (inp[9]) ? 4'b0000 : 4'b0100;
												assign node19695 = (inp[5]) ? node19705 : node19696;
													assign node19696 = (inp[3]) ? 4'b0000 : node19697;
														assign node19697 = (inp[4]) ? node19701 : node19698;
															assign node19698 = (inp[9]) ? 4'b0000 : 4'b0100;
															assign node19701 = (inp[9]) ? 4'b0100 : 4'b0000;
													assign node19705 = (inp[3]) ? node19715 : node19706;
														assign node19706 = (inp[12]) ? node19708 : 4'b0000;
															assign node19708 = (inp[9]) ? node19712 : node19709;
																assign node19709 = (inp[4]) ? 4'b0000 : 4'b0100;
																assign node19712 = (inp[4]) ? 4'b0110 : 4'b0000;
														assign node19715 = (inp[4]) ? 4'b0110 : node19716;
															assign node19716 = (inp[12]) ? 4'b0010 : 4'b0110;
											assign node19720 = (inp[0]) ? node19750 : node19721;
												assign node19721 = (inp[3]) ? node19737 : node19722;
													assign node19722 = (inp[5]) ? node19730 : node19723;
														assign node19723 = (inp[4]) ? node19727 : node19724;
															assign node19724 = (inp[9]) ? 4'b0000 : 4'b0100;
															assign node19727 = (inp[9]) ? 4'b0100 : 4'b0000;
														assign node19730 = (inp[12]) ? node19734 : node19731;
															assign node19731 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node19734 = (inp[4]) ? 4'b0110 : 4'b0000;
													assign node19737 = (inp[5]) ? node19745 : node19738;
														assign node19738 = (inp[9]) ? node19742 : node19739;
															assign node19739 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node19742 = (inp[4]) ? 4'b0110 : 4'b0000;
														assign node19745 = (inp[9]) ? node19747 : 4'b0110;
															assign node19747 = (inp[4]) ? 4'b0110 : 4'b0010;
												assign node19750 = (inp[3]) ? node19766 : node19751;
													assign node19751 = (inp[5]) ? node19759 : node19752;
														assign node19752 = (inp[9]) ? node19756 : node19753;
															assign node19753 = (inp[4]) ? 4'b0010 : 4'b0110;
															assign node19756 = (inp[4]) ? 4'b0110 : 4'b0010;
														assign node19759 = (inp[9]) ? node19763 : node19760;
															assign node19760 = (inp[4]) ? 4'b0010 : 4'b0110;
															assign node19763 = (inp[4]) ? 4'b0100 : 4'b0010;
													assign node19766 = (inp[4]) ? 4'b0100 : node19767;
														assign node19767 = (inp[5]) ? node19771 : node19768;
															assign node19768 = (inp[9]) ? 4'b0010 : 4'b0110;
															assign node19771 = (inp[9]) ? 4'b0000 : 4'b0100;
										assign node19775 = (inp[12]) ? node19839 : node19776;
											assign node19776 = (inp[0]) ? node19802 : node19777;
												assign node19777 = (inp[3]) ? node19785 : node19778;
													assign node19778 = (inp[15]) ? 4'b1001 : node19779;
														assign node19779 = (inp[4]) ? 4'b1011 : node19780;
															assign node19780 = (inp[9]) ? 4'b1011 : 4'b1111;
													assign node19785 = (inp[15]) ? node19793 : node19786;
														assign node19786 = (inp[9]) ? node19790 : node19787;
															assign node19787 = (inp[5]) ? 4'b1001 : 4'b1011;
															assign node19790 = (inp[4]) ? 4'b1101 : 4'b1001;
														assign node19793 = (inp[5]) ? node19795 : 4'b1001;
															assign node19795 = (inp[4]) ? node19799 : node19796;
																assign node19796 = (inp[9]) ? 4'b1011 : 4'b1111;
																assign node19799 = (inp[9]) ? 4'b1111 : 4'b1011;
												assign node19802 = (inp[15]) ? node19820 : node19803;
													assign node19803 = (inp[5]) ? node19809 : node19804;
														assign node19804 = (inp[4]) ? 4'b1001 : node19805;
															assign node19805 = (inp[9]) ? 4'b1001 : 4'b1101;
														assign node19809 = (inp[3]) ? node19817 : node19810;
															assign node19810 = (inp[4]) ? node19814 : node19811;
																assign node19811 = (inp[9]) ? 4'b1001 : 4'b1101;
																assign node19814 = (inp[9]) ? 4'b1111 : 4'b1001;
															assign node19817 = (inp[4]) ? 4'b1011 : 4'b1111;
													assign node19820 = (inp[5]) ? node19826 : node19821;
														assign node19821 = (inp[4]) ? 4'b1111 : node19822;
															assign node19822 = (inp[9]) ? 4'b1011 : 4'b1111;
														assign node19826 = (inp[3]) ? node19832 : node19827;
															assign node19827 = (inp[9]) ? 4'b1101 : node19828;
																assign node19828 = (inp[4]) ? 4'b1011 : 4'b1111;
															assign node19832 = (inp[9]) ? node19836 : node19833;
																assign node19833 = (inp[4]) ? 4'b1001 : 4'b1101;
																assign node19836 = (inp[4]) ? 4'b1101 : 4'b1001;
											assign node19839 = (inp[15]) ? node19877 : node19840;
												assign node19840 = (inp[0]) ? node19856 : node19841;
													assign node19841 = (inp[5]) ? node19851 : node19842;
														assign node19842 = (inp[3]) ? node19848 : node19843;
															assign node19843 = (inp[4]) ? node19845 : 4'b1111;
																assign node19845 = (inp[9]) ? 4'b1011 : 4'b1111;
															assign node19848 = (inp[4]) ? 4'b1001 : 4'b1011;
														assign node19851 = (inp[9]) ? node19853 : 4'b1101;
															assign node19853 = (inp[4]) ? 4'b1001 : 4'b1101;
													assign node19856 = (inp[3]) ? node19864 : node19857;
														assign node19857 = (inp[5]) ? node19859 : 4'b1001;
															assign node19859 = (inp[9]) ? node19861 : 4'b1111;
																assign node19861 = (inp[4]) ? 4'b1011 : 4'b1111;
														assign node19864 = (inp[5]) ? node19870 : node19865;
															assign node19865 = (inp[4]) ? node19867 : 4'b1111;
																assign node19867 = (inp[9]) ? 4'b1011 : 4'b1111;
															assign node19870 = (inp[9]) ? node19874 : node19871;
																assign node19871 = (inp[4]) ? 4'b1111 : 4'b1011;
																assign node19874 = (inp[4]) ? 4'b1011 : 4'b1111;
												assign node19877 = (inp[0]) ? node19897 : node19878;
													assign node19878 = (inp[5]) ? node19890 : node19879;
														assign node19879 = (inp[3]) ? node19885 : node19880;
															assign node19880 = (inp[9]) ? 4'b1101 : node19881;
																assign node19881 = (inp[4]) ? 4'b1101 : 4'b1001;
															assign node19885 = (inp[4]) ? 4'b1111 : node19886;
																assign node19886 = (inp[9]) ? 4'b1111 : 4'b1001;
														assign node19890 = (inp[4]) ? node19894 : node19891;
															assign node19891 = (inp[9]) ? 4'b1111 : 4'b1001;
															assign node19894 = (inp[9]) ? 4'b1011 : 4'b1111;
													assign node19897 = (inp[4]) ? node19905 : node19898;
														assign node19898 = (inp[9]) ? node19900 : 4'b1011;
															assign node19900 = (inp[3]) ? 4'b1101 : node19901;
																assign node19901 = (inp[5]) ? 4'b1101 : 4'b1111;
														assign node19905 = (inp[9]) ? node19907 : 4'b1101;
															assign node19907 = (inp[3]) ? 4'b1001 : node19908;
																assign node19908 = (inp[5]) ? 4'b1001 : 4'b1011;
									assign node19912 = (inp[15]) ? node20036 : node19913;
										assign node19913 = (inp[5]) ? node19973 : node19914;
											assign node19914 = (inp[0]) ? node19944 : node19915;
												assign node19915 = (inp[3]) ? node19933 : node19916;
													assign node19916 = (inp[14]) ? node19924 : node19917;
														assign node19917 = (inp[9]) ? node19919 : 4'b1111;
															assign node19919 = (inp[4]) ? node19921 : 4'b1111;
																assign node19921 = (inp[12]) ? 4'b1011 : 4'b1111;
														assign node19924 = (inp[12]) ? 4'b1011 : node19925;
															assign node19925 = (inp[9]) ? node19929 : node19926;
																assign node19926 = (inp[4]) ? 4'b1011 : 4'b1111;
																assign node19929 = (inp[4]) ? 4'b1111 : 4'b1011;
													assign node19933 = (inp[12]) ? node19939 : node19934;
														assign node19934 = (inp[4]) ? 4'b1101 : node19935;
															assign node19935 = (inp[9]) ? 4'b1011 : 4'b1111;
														assign node19939 = (inp[9]) ? node19941 : 4'b1101;
															assign node19941 = (inp[4]) ? 4'b1001 : 4'b1101;
												assign node19944 = (inp[3]) ? node19958 : node19945;
													assign node19945 = (inp[12]) ? node19953 : node19946;
														assign node19946 = (inp[4]) ? node19950 : node19947;
															assign node19947 = (inp[9]) ? 4'b1001 : 4'b1101;
															assign node19950 = (inp[9]) ? 4'b1101 : 4'b1001;
														assign node19953 = (inp[14]) ? node19955 : 4'b1101;
															assign node19955 = (inp[4]) ? 4'b1001 : 4'b1101;
													assign node19958 = (inp[9]) ? node19966 : node19959;
														assign node19959 = (inp[12]) ? node19963 : node19960;
															assign node19960 = (inp[4]) ? 4'b1001 : 4'b1101;
															assign node19963 = (inp[4]) ? 4'b1111 : 4'b1001;
														assign node19966 = (inp[4]) ? node19970 : node19967;
															assign node19967 = (inp[12]) ? 4'b1111 : 4'b1001;
															assign node19970 = (inp[12]) ? 4'b1011 : 4'b1111;
											assign node19973 = (inp[0]) ? node20011 : node19974;
												assign node19974 = (inp[3]) ? node19988 : node19975;
													assign node19975 = (inp[9]) ? node19983 : node19976;
														assign node19976 = (inp[4]) ? node19980 : node19977;
															assign node19977 = (inp[12]) ? 4'b1011 : 4'b1111;
															assign node19980 = (inp[12]) ? 4'b1101 : 4'b1011;
														assign node19983 = (inp[4]) ? node19985 : 4'b1101;
															assign node19985 = (inp[12]) ? 4'b1001 : 4'b1101;
													assign node19988 = (inp[14]) ? node20004 : node19989;
														assign node19989 = (inp[4]) ? node19997 : node19990;
															assign node19990 = (inp[9]) ? node19994 : node19991;
																assign node19991 = (inp[12]) ? 4'b1001 : 4'b1101;
																assign node19994 = (inp[12]) ? 4'b1101 : 4'b1001;
															assign node19997 = (inp[9]) ? node20001 : node19998;
																assign node19998 = (inp[12]) ? 4'b1101 : 4'b1001;
																assign node20001 = (inp[12]) ? 4'b1001 : 4'b1101;
														assign node20004 = (inp[4]) ? 4'b1001 : node20005;
															assign node20005 = (inp[12]) ? node20007 : 4'b1001;
																assign node20007 = (inp[9]) ? 4'b1101 : 4'b1001;
												assign node20011 = (inp[3]) ? node20021 : node20012;
													assign node20012 = (inp[9]) ? node20018 : node20013;
														assign node20013 = (inp[4]) ? 4'b1001 : node20014;
															assign node20014 = (inp[12]) ? 4'b1001 : 4'b1101;
														assign node20018 = (inp[14]) ? 4'b1001 : 4'b1111;
													assign node20021 = (inp[14]) ? node20031 : node20022;
														assign node20022 = (inp[12]) ? node20024 : 4'b1011;
															assign node20024 = (inp[9]) ? node20028 : node20025;
																assign node20025 = (inp[4]) ? 4'b1111 : 4'b1011;
																assign node20028 = (inp[4]) ? 4'b1011 : 4'b1111;
														assign node20031 = (inp[4]) ? 4'b1111 : node20032;
															assign node20032 = (inp[12]) ? 4'b1111 : 4'b1011;
										assign node20036 = (inp[0]) ? node20104 : node20037;
											assign node20037 = (inp[5]) ? node20067 : node20038;
												assign node20038 = (inp[3]) ? node20054 : node20039;
													assign node20039 = (inp[12]) ? node20047 : node20040;
														assign node20040 = (inp[4]) ? node20044 : node20041;
															assign node20041 = (inp[9]) ? 4'b1001 : 4'b1101;
															assign node20044 = (inp[9]) ? 4'b1101 : 4'b1001;
														assign node20047 = (inp[4]) ? node20051 : node20048;
															assign node20048 = (inp[9]) ? 4'b1101 : 4'b1001;
															assign node20051 = (inp[9]) ? 4'b1001 : 4'b1101;
													assign node20054 = (inp[9]) ? node20062 : node20055;
														assign node20055 = (inp[12]) ? node20059 : node20056;
															assign node20056 = (inp[4]) ? 4'b1001 : 4'b1101;
															assign node20059 = (inp[4]) ? 4'b1111 : 4'b1001;
														assign node20062 = (inp[12]) ? node20064 : 4'b1111;
															assign node20064 = (inp[4]) ? 4'b1011 : 4'b1111;
												assign node20067 = (inp[3]) ? node20083 : node20068;
													assign node20068 = (inp[12]) ? node20076 : node20069;
														assign node20069 = (inp[9]) ? node20073 : node20070;
															assign node20070 = (inp[4]) ? 4'b1001 : 4'b1101;
															assign node20073 = (inp[4]) ? 4'b1111 : 4'b1001;
														assign node20076 = (inp[14]) ? node20078 : 4'b1111;
															assign node20078 = (inp[9]) ? node20080 : 4'b1111;
																assign node20080 = (inp[4]) ? 4'b1011 : 4'b1111;
													assign node20083 = (inp[9]) ? node20091 : node20084;
														assign node20084 = (inp[12]) ? node20088 : node20085;
															assign node20085 = (inp[4]) ? 4'b1011 : 4'b1111;
															assign node20088 = (inp[4]) ? 4'b1111 : 4'b1011;
														assign node20091 = (inp[14]) ? node20097 : node20092;
															assign node20092 = (inp[4]) ? node20094 : 4'b1011;
																assign node20094 = (inp[12]) ? 4'b1011 : 4'b1111;
															assign node20097 = (inp[12]) ? node20101 : node20098;
																assign node20098 = (inp[4]) ? 4'b1111 : 4'b1011;
																assign node20101 = (inp[4]) ? 4'b1011 : 4'b1111;
											assign node20104 = (inp[3]) ? node20138 : node20105;
												assign node20105 = (inp[5]) ? node20123 : node20106;
													assign node20106 = (inp[14]) ? node20114 : node20107;
														assign node20107 = (inp[4]) ? node20111 : node20108;
															assign node20108 = (inp[12]) ? 4'b1011 : 4'b1111;
															assign node20111 = (inp[12]) ? 4'b1111 : 4'b1011;
														assign node20114 = (inp[9]) ? node20116 : 4'b1011;
															assign node20116 = (inp[12]) ? node20120 : node20117;
																assign node20117 = (inp[4]) ? 4'b1111 : 4'b1011;
																assign node20120 = (inp[4]) ? 4'b1011 : 4'b1111;
													assign node20123 = (inp[4]) ? node20131 : node20124;
														assign node20124 = (inp[9]) ? node20128 : node20125;
															assign node20125 = (inp[12]) ? 4'b1011 : 4'b1111;
															assign node20128 = (inp[12]) ? 4'b1101 : 4'b1011;
														assign node20131 = (inp[9]) ? node20135 : node20132;
															assign node20132 = (inp[12]) ? 4'b1101 : 4'b1011;
															assign node20135 = (inp[12]) ? 4'b1001 : 4'b1101;
												assign node20138 = (inp[5]) ? node20152 : node20139;
													assign node20139 = (inp[9]) ? node20147 : node20140;
														assign node20140 = (inp[4]) ? node20144 : node20141;
															assign node20141 = (inp[12]) ? 4'b1011 : 4'b1111;
															assign node20144 = (inp[12]) ? 4'b1101 : 4'b1011;
														assign node20147 = (inp[12]) ? node20149 : 4'b1101;
															assign node20149 = (inp[4]) ? 4'b1001 : 4'b1101;
													assign node20152 = (inp[14]) ? node20166 : node20153;
														assign node20153 = (inp[9]) ? node20161 : node20154;
															assign node20154 = (inp[4]) ? node20158 : node20155;
																assign node20155 = (inp[12]) ? 4'b1001 : 4'b1101;
																assign node20158 = (inp[12]) ? 4'b1101 : 4'b1001;
															assign node20161 = (inp[4]) ? node20163 : 4'b1001;
																assign node20163 = (inp[12]) ? 4'b1001 : 4'b1101;
														assign node20166 = (inp[4]) ? node20168 : 4'b1101;
															assign node20168 = (inp[12]) ? 4'b1101 : 4'b1001;
								assign node20171 = (inp[14]) ? node20455 : node20172;
									assign node20172 = (inp[2]) ? node20334 : node20173;
										assign node20173 = (inp[3]) ? node20245 : node20174;
											assign node20174 = (inp[4]) ? node20206 : node20175;
												assign node20175 = (inp[0]) ? node20191 : node20176;
													assign node20176 = (inp[15]) ? node20184 : node20177;
														assign node20177 = (inp[9]) ? node20181 : node20178;
															assign node20178 = (inp[12]) ? 4'b1011 : 4'b1111;
															assign node20181 = (inp[12]) ? 4'b1101 : 4'b1011;
														assign node20184 = (inp[12]) ? node20188 : node20185;
															assign node20185 = (inp[9]) ? 4'b1001 : 4'b1101;
															assign node20188 = (inp[9]) ? 4'b1101 : 4'b1001;
													assign node20191 = (inp[15]) ? node20197 : node20192;
														assign node20192 = (inp[12]) ? node20194 : 4'b1101;
															assign node20194 = (inp[9]) ? 4'b1101 : 4'b1001;
														assign node20197 = (inp[5]) ? node20199 : 4'b1111;
															assign node20199 = (inp[9]) ? node20203 : node20200;
																assign node20200 = (inp[12]) ? 4'b1011 : 4'b1111;
																assign node20203 = (inp[12]) ? 4'b1101 : 4'b1011;
												assign node20206 = (inp[0]) ? node20232 : node20207;
													assign node20207 = (inp[15]) ? node20221 : node20208;
														assign node20208 = (inp[5]) ? node20214 : node20209;
															assign node20209 = (inp[12]) ? node20211 : 4'b1011;
																assign node20211 = (inp[9]) ? 4'b1011 : 4'b1111;
															assign node20214 = (inp[12]) ? node20218 : node20215;
																assign node20215 = (inp[9]) ? 4'b1101 : 4'b1011;
																assign node20218 = (inp[9]) ? 4'b1001 : 4'b1101;
														assign node20221 = (inp[5]) ? node20227 : node20222;
															assign node20222 = (inp[12]) ? node20224 : 4'b1001;
																assign node20224 = (inp[9]) ? 4'b1001 : 4'b1101;
															assign node20227 = (inp[9]) ? 4'b1111 : node20228;
																assign node20228 = (inp[12]) ? 4'b1111 : 4'b1001;
													assign node20232 = (inp[15]) ? node20240 : node20233;
														assign node20233 = (inp[12]) ? node20235 : 4'b1001;
															assign node20235 = (inp[5]) ? node20237 : 4'b1001;
																assign node20237 = (inp[9]) ? 4'b1011 : 4'b1111;
														assign node20240 = (inp[12]) ? 4'b1001 : node20241;
															assign node20241 = (inp[9]) ? 4'b1111 : 4'b1011;
											assign node20245 = (inp[9]) ? node20291 : node20246;
												assign node20246 = (inp[4]) ? node20270 : node20247;
													assign node20247 = (inp[12]) ? node20261 : node20248;
														assign node20248 = (inp[5]) ? node20256 : node20249;
															assign node20249 = (inp[0]) ? node20253 : node20250;
																assign node20250 = (inp[15]) ? 4'b1101 : 4'b1111;
																assign node20253 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node20256 = (inp[15]) ? node20258 : 4'b1101;
																assign node20258 = (inp[0]) ? 4'b1101 : 4'b1111;
														assign node20261 = (inp[5]) ? node20263 : 4'b1001;
															assign node20263 = (inp[15]) ? node20267 : node20264;
																assign node20264 = (inp[0]) ? 4'b1011 : 4'b1001;
																assign node20267 = (inp[0]) ? 4'b1001 : 4'b1011;
													assign node20270 = (inp[12]) ? node20276 : node20271;
														assign node20271 = (inp[0]) ? node20273 : 4'b1011;
															assign node20273 = (inp[5]) ? 4'b1011 : 4'b1001;
														assign node20276 = (inp[5]) ? node20284 : node20277;
															assign node20277 = (inp[0]) ? node20281 : node20278;
																assign node20278 = (inp[15]) ? 4'b1111 : 4'b1101;
																assign node20281 = (inp[15]) ? 4'b1101 : 4'b1111;
															assign node20284 = (inp[15]) ? node20288 : node20285;
																assign node20285 = (inp[0]) ? 4'b1111 : 4'b1101;
																assign node20288 = (inp[0]) ? 4'b1101 : 4'b1111;
												assign node20291 = (inp[5]) ? node20313 : node20292;
													assign node20292 = (inp[12]) ? node20300 : node20293;
														assign node20293 = (inp[4]) ? 4'b1111 : node20294;
															assign node20294 = (inp[15]) ? node20296 : 4'b1011;
																assign node20296 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node20300 = (inp[4]) ? node20308 : node20301;
															assign node20301 = (inp[15]) ? node20305 : node20302;
																assign node20302 = (inp[0]) ? 4'b1111 : 4'b1101;
																assign node20305 = (inp[0]) ? 4'b1101 : 4'b1111;
															assign node20308 = (inp[0]) ? 4'b1011 : node20309;
																assign node20309 = (inp[15]) ? 4'b1011 : 4'b1001;
													assign node20313 = (inp[0]) ? node20327 : node20314;
														assign node20314 = (inp[15]) ? node20320 : node20315;
															assign node20315 = (inp[4]) ? node20317 : 4'b1001;
																assign node20317 = (inp[12]) ? 4'b1001 : 4'b1101;
															assign node20320 = (inp[12]) ? node20324 : node20321;
																assign node20321 = (inp[4]) ? 4'b1111 : 4'b1011;
																assign node20324 = (inp[4]) ? 4'b1011 : 4'b1111;
														assign node20327 = (inp[15]) ? node20329 : 4'b1111;
															assign node20329 = (inp[4]) ? 4'b1101 : node20330;
																assign node20330 = (inp[12]) ? 4'b1101 : 4'b1001;
										assign node20334 = (inp[15]) ? node20398 : node20335;
											assign node20335 = (inp[5]) ? node20367 : node20336;
												assign node20336 = (inp[0]) ? node20354 : node20337;
													assign node20337 = (inp[3]) ? node20343 : node20338;
														assign node20338 = (inp[9]) ? 4'b1110 : node20339;
															assign node20339 = (inp[4]) ? 4'b1110 : 4'b1010;
														assign node20343 = (inp[12]) ? node20349 : node20344;
															assign node20344 = (inp[4]) ? 4'b1010 : node20345;
																assign node20345 = (inp[9]) ? 4'b1010 : 4'b1110;
															assign node20349 = (inp[4]) ? node20351 : 4'b1100;
																assign node20351 = (inp[9]) ? 4'b1000 : 4'b1100;
													assign node20354 = (inp[9]) ? node20360 : node20355;
														assign node20355 = (inp[12]) ? 4'b1000 : node20356;
															assign node20356 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node20360 = (inp[3]) ? node20362 : 4'b1000;
															assign node20362 = (inp[4]) ? node20364 : 4'b1000;
																assign node20364 = (inp[12]) ? 4'b1010 : 4'b1110;
												assign node20367 = (inp[0]) ? node20385 : node20368;
													assign node20368 = (inp[3]) ? node20380 : node20369;
														assign node20369 = (inp[12]) ? node20375 : node20370;
															assign node20370 = (inp[9]) ? 4'b1010 : node20371;
																assign node20371 = (inp[4]) ? 4'b1010 : 4'b1110;
															assign node20375 = (inp[9]) ? 4'b1100 : node20376;
																assign node20376 = (inp[4]) ? 4'b1100 : 4'b1010;
														assign node20380 = (inp[12]) ? node20382 : 4'b1100;
															assign node20382 = (inp[4]) ? 4'b1000 : 4'b1100;
													assign node20385 = (inp[9]) ? node20391 : node20386;
														assign node20386 = (inp[12]) ? 4'b1110 : node20387;
															assign node20387 = (inp[4]) ? 4'b1000 : 4'b1110;
														assign node20391 = (inp[12]) ? node20395 : node20392;
															assign node20392 = (inp[3]) ? 4'b1010 : 4'b1110;
															assign node20395 = (inp[4]) ? 4'b1010 : 4'b1110;
											assign node20398 = (inp[12]) ? node20424 : node20399;
												assign node20399 = (inp[0]) ? node20411 : node20400;
													assign node20400 = (inp[3]) ? node20408 : node20401;
														assign node20401 = (inp[4]) ? node20405 : node20402;
															assign node20402 = (inp[9]) ? 4'b1000 : 4'b1100;
															assign node20405 = (inp[9]) ? 4'b1100 : 4'b1000;
														assign node20408 = (inp[5]) ? 4'b1010 : 4'b1000;
													assign node20411 = (inp[3]) ? node20413 : 4'b1010;
														assign node20413 = (inp[5]) ? node20419 : node20414;
															assign node20414 = (inp[9]) ? node20416 : 4'b1010;
																assign node20416 = (inp[4]) ? 4'b1100 : 4'b1010;
															assign node20419 = (inp[9]) ? 4'b1100 : node20420;
																assign node20420 = (inp[4]) ? 4'b1000 : 4'b1100;
												assign node20424 = (inp[0]) ? node20440 : node20425;
													assign node20425 = (inp[3]) ? node20433 : node20426;
														assign node20426 = (inp[4]) ? node20430 : node20427;
															assign node20427 = (inp[9]) ? 4'b1100 : 4'b1000;
															assign node20430 = (inp[5]) ? 4'b1110 : 4'b1000;
														assign node20433 = (inp[9]) ? node20437 : node20434;
															assign node20434 = (inp[5]) ? 4'b1010 : 4'b1000;
															assign node20437 = (inp[4]) ? 4'b1010 : 4'b1110;
													assign node20440 = (inp[3]) ? node20446 : node20441;
														assign node20441 = (inp[5]) ? node20443 : 4'b1110;
															assign node20443 = (inp[4]) ? 4'b1000 : 4'b1010;
														assign node20446 = (inp[4]) ? node20452 : node20447;
															assign node20447 = (inp[9]) ? 4'b1100 : node20448;
																assign node20448 = (inp[5]) ? 4'b1000 : 4'b1010;
															assign node20452 = (inp[9]) ? 4'b1000 : 4'b1100;
									assign node20455 = (inp[0]) ? node20591 : node20456;
										assign node20456 = (inp[5]) ? node20522 : node20457;
											assign node20457 = (inp[15]) ? node20493 : node20458;
												assign node20458 = (inp[3]) ? node20476 : node20459;
													assign node20459 = (inp[12]) ? node20467 : node20460;
														assign node20460 = (inp[9]) ? node20464 : node20461;
															assign node20461 = (inp[4]) ? 4'b1010 : 4'b1110;
															assign node20464 = (inp[4]) ? 4'b1110 : 4'b1010;
														assign node20467 = (inp[2]) ? 4'b1110 : node20468;
															assign node20468 = (inp[9]) ? node20472 : node20469;
																assign node20469 = (inp[4]) ? 4'b1110 : 4'b1010;
																assign node20472 = (inp[4]) ? 4'b1010 : 4'b1110;
													assign node20476 = (inp[9]) ? node20484 : node20477;
														assign node20477 = (inp[12]) ? node20481 : node20478;
															assign node20478 = (inp[4]) ? 4'b1010 : 4'b1110;
															assign node20481 = (inp[4]) ? 4'b1100 : 4'b1010;
														assign node20484 = (inp[2]) ? node20490 : node20485;
															assign node20485 = (inp[4]) ? node20487 : 4'b1100;
																assign node20487 = (inp[12]) ? 4'b1000 : 4'b1100;
															assign node20490 = (inp[12]) ? 4'b1100 : 4'b1010;
												assign node20493 = (inp[3]) ? node20507 : node20494;
													assign node20494 = (inp[12]) ? node20502 : node20495;
														assign node20495 = (inp[9]) ? node20499 : node20496;
															assign node20496 = (inp[4]) ? 4'b1000 : 4'b1100;
															assign node20499 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node20502 = (inp[4]) ? node20504 : 4'b1000;
															assign node20504 = (inp[9]) ? 4'b1000 : 4'b1100;
													assign node20507 = (inp[4]) ? node20515 : node20508;
														assign node20508 = (inp[2]) ? node20510 : 4'b1000;
															assign node20510 = (inp[9]) ? node20512 : 4'b1000;
																assign node20512 = (inp[12]) ? 4'b1110 : 4'b1000;
														assign node20515 = (inp[12]) ? node20519 : node20516;
															assign node20516 = (inp[9]) ? 4'b1110 : 4'b1000;
															assign node20519 = (inp[9]) ? 4'b1010 : 4'b1110;
											assign node20522 = (inp[15]) ? node20552 : node20523;
												assign node20523 = (inp[3]) ? node20539 : node20524;
													assign node20524 = (inp[12]) ? node20530 : node20525;
														assign node20525 = (inp[4]) ? 4'b1010 : node20526;
															assign node20526 = (inp[9]) ? 4'b1010 : 4'b1110;
														assign node20530 = (inp[2]) ? node20536 : node20531;
															assign node20531 = (inp[4]) ? 4'b1100 : node20532;
																assign node20532 = (inp[9]) ? 4'b1100 : 4'b1010;
															assign node20536 = (inp[9]) ? 4'b1000 : 4'b1010;
													assign node20539 = (inp[4]) ? node20547 : node20540;
														assign node20540 = (inp[9]) ? node20544 : node20541;
															assign node20541 = (inp[12]) ? 4'b1000 : 4'b1100;
															assign node20544 = (inp[12]) ? 4'b1100 : 4'b1000;
														assign node20547 = (inp[9]) ? 4'b1100 : node20548;
															assign node20548 = (inp[12]) ? 4'b1100 : 4'b1000;
												assign node20552 = (inp[3]) ? node20566 : node20553;
													assign node20553 = (inp[12]) ? node20561 : node20554;
														assign node20554 = (inp[4]) ? node20558 : node20555;
															assign node20555 = (inp[9]) ? 4'b1000 : 4'b1100;
															assign node20558 = (inp[9]) ? 4'b1110 : 4'b1000;
														assign node20561 = (inp[4]) ? node20563 : 4'b1110;
															assign node20563 = (inp[9]) ? 4'b1010 : 4'b1110;
													assign node20566 = (inp[12]) ? node20576 : node20567;
														assign node20567 = (inp[2]) ? node20571 : node20568;
															assign node20568 = (inp[4]) ? 4'b1110 : 4'b1010;
															assign node20571 = (inp[4]) ? 4'b1010 : node20572;
																assign node20572 = (inp[9]) ? 4'b1010 : 4'b1110;
														assign node20576 = (inp[2]) ? node20584 : node20577;
															assign node20577 = (inp[9]) ? node20581 : node20578;
																assign node20578 = (inp[4]) ? 4'b1110 : 4'b1010;
																assign node20581 = (inp[4]) ? 4'b1010 : 4'b1110;
															assign node20584 = (inp[9]) ? node20588 : node20585;
																assign node20585 = (inp[4]) ? 4'b1110 : 4'b1010;
																assign node20588 = (inp[4]) ? 4'b1010 : 4'b1110;
										assign node20591 = (inp[15]) ? node20641 : node20592;
											assign node20592 = (inp[5]) ? node20614 : node20593;
												assign node20593 = (inp[3]) ? node20601 : node20594;
													assign node20594 = (inp[2]) ? node20596 : 4'b1100;
														assign node20596 = (inp[9]) ? 4'b1000 : node20597;
															assign node20597 = (inp[4]) ? 4'b1100 : 4'b1000;
													assign node20601 = (inp[12]) ? node20609 : node20602;
														assign node20602 = (inp[4]) ? node20606 : node20603;
															assign node20603 = (inp[9]) ? 4'b1000 : 4'b1100;
															assign node20606 = (inp[9]) ? 4'b1110 : 4'b1000;
														assign node20609 = (inp[9]) ? 4'b1110 : node20610;
															assign node20610 = (inp[4]) ? 4'b1110 : 4'b1000;
												assign node20614 = (inp[3]) ? node20630 : node20615;
													assign node20615 = (inp[4]) ? node20623 : node20616;
														assign node20616 = (inp[9]) ? node20620 : node20617;
															assign node20617 = (inp[12]) ? 4'b1000 : 4'b1100;
															assign node20620 = (inp[12]) ? 4'b1110 : 4'b1000;
														assign node20623 = (inp[12]) ? node20627 : node20624;
															assign node20624 = (inp[9]) ? 4'b1110 : 4'b1000;
															assign node20627 = (inp[9]) ? 4'b1010 : 4'b1110;
													assign node20630 = (inp[9]) ? node20634 : node20631;
														assign node20631 = (inp[2]) ? 4'b1010 : 4'b1110;
														assign node20634 = (inp[4]) ? node20638 : node20635;
															assign node20635 = (inp[12]) ? 4'b1110 : 4'b1010;
															assign node20638 = (inp[12]) ? 4'b1010 : 4'b1110;
											assign node20641 = (inp[3]) ? node20657 : node20642;
												assign node20642 = (inp[9]) ? node20648 : node20643;
													assign node20643 = (inp[4]) ? 4'b1010 : node20644;
														assign node20644 = (inp[12]) ? 4'b1010 : 4'b1110;
													assign node20648 = (inp[2]) ? node20654 : node20649;
														assign node20649 = (inp[4]) ? 4'b1010 : node20650;
															assign node20650 = (inp[12]) ? 4'b1100 : 4'b1010;
														assign node20654 = (inp[5]) ? 4'b1100 : 4'b1110;
												assign node20657 = (inp[5]) ? node20671 : node20658;
													assign node20658 = (inp[12]) ? node20666 : node20659;
														assign node20659 = (inp[9]) ? node20663 : node20660;
															assign node20660 = (inp[4]) ? 4'b1010 : 4'b1110;
															assign node20663 = (inp[4]) ? 4'b1100 : 4'b1010;
														assign node20666 = (inp[4]) ? node20668 : 4'b1100;
															assign node20668 = (inp[9]) ? 4'b1000 : 4'b1100;
													assign node20671 = (inp[4]) ? node20679 : node20672;
														assign node20672 = (inp[9]) ? node20676 : node20673;
															assign node20673 = (inp[12]) ? 4'b1000 : 4'b1100;
															assign node20676 = (inp[12]) ? 4'b1100 : 4'b1000;
														assign node20679 = (inp[2]) ? 4'b1000 : node20680;
															assign node20680 = (inp[9]) ? 4'b1100 : node20681;
																assign node20681 = (inp[12]) ? 4'b1100 : 4'b1000;
						assign node20686 = (inp[2]) ? node21888 : node20687;
							assign node20687 = (inp[15]) ? node21277 : node20688;
								assign node20688 = (inp[4]) ? node20984 : node20689;
									assign node20689 = (inp[0]) ? node20853 : node20690;
										assign node20690 = (inp[3]) ? node20764 : node20691;
											assign node20691 = (inp[5]) ? node20733 : node20692;
												assign node20692 = (inp[14]) ? node20716 : node20693;
													assign node20693 = (inp[12]) ? node20703 : node20694;
														assign node20694 = (inp[9]) ? node20696 : 4'b1110;
															assign node20696 = (inp[8]) ? node20700 : node20697;
																assign node20697 = (inp[7]) ? 4'b1010 : 4'b1011;
																assign node20700 = (inp[7]) ? 4'b1011 : 4'b1010;
														assign node20703 = (inp[9]) ? node20709 : node20704;
															assign node20704 = (inp[7]) ? 4'b1011 : node20705;
																assign node20705 = (inp[8]) ? 4'b1010 : 4'b1011;
															assign node20709 = (inp[7]) ? node20713 : node20710;
																assign node20710 = (inp[8]) ? 4'b1110 : 4'b1111;
																assign node20713 = (inp[8]) ? 4'b1111 : 4'b1110;
													assign node20716 = (inp[9]) ? node20724 : node20717;
														assign node20717 = (inp[12]) ? 4'b1010 : node20718;
															assign node20718 = (inp[7]) ? 4'b1110 : node20719;
																assign node20719 = (inp[8]) ? 4'b1111 : 4'b1110;
														assign node20724 = (inp[12]) ? 4'b1110 : node20725;
															assign node20725 = (inp[8]) ? node20729 : node20726;
																assign node20726 = (inp[7]) ? 4'b1011 : 4'b1010;
																assign node20729 = (inp[7]) ? 4'b1010 : 4'b1011;
												assign node20733 = (inp[12]) ? node20751 : node20734;
													assign node20734 = (inp[9]) ? node20744 : node20735;
														assign node20735 = (inp[8]) ? node20737 : 4'b1111;
															assign node20737 = (inp[7]) ? node20741 : node20738;
																assign node20738 = (inp[14]) ? 4'b1111 : 4'b1110;
																assign node20741 = (inp[14]) ? 4'b1110 : 4'b1111;
														assign node20744 = (inp[7]) ? 4'b1011 : node20745;
															assign node20745 = (inp[14]) ? node20747 : 4'b1010;
																assign node20747 = (inp[8]) ? 4'b1011 : 4'b1010;
													assign node20751 = (inp[9]) ? node20761 : node20752;
														assign node20752 = (inp[7]) ? node20754 : 4'b1011;
															assign node20754 = (inp[14]) ? node20758 : node20755;
																assign node20755 = (inp[8]) ? 4'b1011 : 4'b1010;
																assign node20758 = (inp[8]) ? 4'b1010 : 4'b1011;
														assign node20761 = (inp[8]) ? 4'b1100 : 4'b1101;
											assign node20764 = (inp[5]) ? node20810 : node20765;
												assign node20765 = (inp[12]) ? node20791 : node20766;
													assign node20766 = (inp[9]) ? node20778 : node20767;
														assign node20767 = (inp[14]) ? node20773 : node20768;
															assign node20768 = (inp[7]) ? node20770 : 4'b1111;
																assign node20770 = (inp[8]) ? 4'b1111 : 4'b1110;
															assign node20773 = (inp[7]) ? node20775 : 4'b1110;
																assign node20775 = (inp[8]) ? 4'b1110 : 4'b1111;
														assign node20778 = (inp[14]) ? node20786 : node20779;
															assign node20779 = (inp[8]) ? node20783 : node20780;
																assign node20780 = (inp[7]) ? 4'b1010 : 4'b1011;
																assign node20783 = (inp[7]) ? 4'b1011 : 4'b1010;
															assign node20786 = (inp[8]) ? 4'b1011 : node20787;
																assign node20787 = (inp[7]) ? 4'b1011 : 4'b1010;
													assign node20791 = (inp[9]) ? node20799 : node20792;
														assign node20792 = (inp[14]) ? 4'b1011 : node20793;
															assign node20793 = (inp[7]) ? node20795 : 4'b1010;
																assign node20795 = (inp[8]) ? 4'b1011 : 4'b1010;
														assign node20799 = (inp[8]) ? node20805 : node20800;
															assign node20800 = (inp[14]) ? node20802 : 4'b1101;
																assign node20802 = (inp[7]) ? 4'b1101 : 4'b1100;
															assign node20805 = (inp[7]) ? 4'b1100 : node20806;
																assign node20806 = (inp[14]) ? 4'b1101 : 4'b1100;
												assign node20810 = (inp[9]) ? node20828 : node20811;
													assign node20811 = (inp[12]) ? node20817 : node20812;
														assign node20812 = (inp[14]) ? 4'b1100 : node20813;
															assign node20813 = (inp[8]) ? 4'b1101 : 4'b1100;
														assign node20817 = (inp[14]) ? node20823 : node20818;
															assign node20818 = (inp[7]) ? node20820 : 4'b1000;
																assign node20820 = (inp[8]) ? 4'b1001 : 4'b1000;
															assign node20823 = (inp[8]) ? node20825 : 4'b1001;
																assign node20825 = (inp[7]) ? 4'b1000 : 4'b1001;
													assign node20828 = (inp[12]) ? node20838 : node20829;
														assign node20829 = (inp[7]) ? 4'b1001 : node20830;
															assign node20830 = (inp[14]) ? node20834 : node20831;
																assign node20831 = (inp[8]) ? 4'b1000 : 4'b1001;
																assign node20834 = (inp[8]) ? 4'b1001 : 4'b1000;
														assign node20838 = (inp[14]) ? node20846 : node20839;
															assign node20839 = (inp[7]) ? node20843 : node20840;
																assign node20840 = (inp[8]) ? 4'b1100 : 4'b1101;
																assign node20843 = (inp[8]) ? 4'b1101 : 4'b1100;
															assign node20846 = (inp[8]) ? node20850 : node20847;
																assign node20847 = (inp[7]) ? 4'b1101 : 4'b1100;
																assign node20850 = (inp[7]) ? 4'b1100 : 4'b1101;
										assign node20853 = (inp[3]) ? node20909 : node20854;
											assign node20854 = (inp[9]) ? node20882 : node20855;
												assign node20855 = (inp[12]) ? node20869 : node20856;
													assign node20856 = (inp[8]) ? node20864 : node20857;
														assign node20857 = (inp[7]) ? node20861 : node20858;
															assign node20858 = (inp[14]) ? 4'b1100 : 4'b1101;
															assign node20861 = (inp[14]) ? 4'b1101 : 4'b1100;
														assign node20864 = (inp[14]) ? node20866 : 4'b1101;
															assign node20866 = (inp[7]) ? 4'b1100 : 4'b1101;
													assign node20869 = (inp[7]) ? node20877 : node20870;
														assign node20870 = (inp[8]) ? node20874 : node20871;
															assign node20871 = (inp[14]) ? 4'b1000 : 4'b1001;
															assign node20874 = (inp[14]) ? 4'b1001 : 4'b1000;
														assign node20877 = (inp[5]) ? node20879 : 4'b1000;
															assign node20879 = (inp[14]) ? 4'b1000 : 4'b1001;
												assign node20882 = (inp[12]) ? node20896 : node20883;
													assign node20883 = (inp[8]) ? node20891 : node20884;
														assign node20884 = (inp[14]) ? node20888 : node20885;
															assign node20885 = (inp[7]) ? 4'b1000 : 4'b1001;
															assign node20888 = (inp[7]) ? 4'b1001 : 4'b1000;
														assign node20891 = (inp[7]) ? 4'b1000 : node20892;
															assign node20892 = (inp[14]) ? 4'b1001 : 4'b1000;
													assign node20896 = (inp[5]) ? node20902 : node20897;
														assign node20897 = (inp[8]) ? node20899 : 4'b1101;
															assign node20899 = (inp[7]) ? 4'b1100 : 4'b1101;
														assign node20902 = (inp[7]) ? node20904 : 4'b1111;
															assign node20904 = (inp[14]) ? node20906 : 4'b1111;
																assign node20906 = (inp[8]) ? 4'b1110 : 4'b1111;
											assign node20909 = (inp[5]) ? node20943 : node20910;
												assign node20910 = (inp[12]) ? node20922 : node20911;
													assign node20911 = (inp[9]) ? node20915 : node20912;
														assign node20912 = (inp[8]) ? 4'b1101 : 4'b1100;
														assign node20915 = (inp[7]) ? node20917 : 4'b1001;
															assign node20917 = (inp[8]) ? 4'b1000 : node20918;
																assign node20918 = (inp[14]) ? 4'b1001 : 4'b1000;
													assign node20922 = (inp[9]) ? node20930 : node20923;
														assign node20923 = (inp[14]) ? node20925 : 4'b1000;
															assign node20925 = (inp[8]) ? 4'b1001 : node20926;
																assign node20926 = (inp[7]) ? 4'b1001 : 4'b1000;
														assign node20930 = (inp[8]) ? node20938 : node20931;
															assign node20931 = (inp[14]) ? node20935 : node20932;
																assign node20932 = (inp[7]) ? 4'b1110 : 4'b1111;
																assign node20935 = (inp[7]) ? 4'b1111 : 4'b1110;
															assign node20938 = (inp[14]) ? node20940 : 4'b1111;
																assign node20940 = (inp[7]) ? 4'b1110 : 4'b1111;
												assign node20943 = (inp[9]) ? node20967 : node20944;
													assign node20944 = (inp[12]) ? node20956 : node20945;
														assign node20945 = (inp[14]) ? node20951 : node20946;
															assign node20946 = (inp[8]) ? 4'b1110 : node20947;
																assign node20947 = (inp[7]) ? 4'b1110 : 4'b1111;
															assign node20951 = (inp[7]) ? 4'b1111 : node20952;
																assign node20952 = (inp[8]) ? 4'b1111 : 4'b1110;
														assign node20956 = (inp[8]) ? node20962 : node20957;
															assign node20957 = (inp[7]) ? 4'b1010 : node20958;
																assign node20958 = (inp[14]) ? 4'b1010 : 4'b1011;
															assign node20962 = (inp[7]) ? 4'b1011 : node20963;
																assign node20963 = (inp[14]) ? 4'b1011 : 4'b1010;
													assign node20967 = (inp[12]) ? node20981 : node20968;
														assign node20968 = (inp[7]) ? node20976 : node20969;
															assign node20969 = (inp[14]) ? node20973 : node20970;
																assign node20970 = (inp[8]) ? 4'b1010 : 4'b1011;
																assign node20973 = (inp[8]) ? 4'b1011 : 4'b1010;
															assign node20976 = (inp[14]) ? node20978 : 4'b1010;
																assign node20978 = (inp[8]) ? 4'b1010 : 4'b1011;
														assign node20981 = (inp[7]) ? 4'b1111 : 4'b1110;
									assign node20984 = (inp[0]) ? node21120 : node20985;
										assign node20985 = (inp[5]) ? node21047 : node20986;
											assign node20986 = (inp[3]) ? node21018 : node20987;
												assign node20987 = (inp[7]) ? node21007 : node20988;
													assign node20988 = (inp[8]) ? node20996 : node20989;
														assign node20989 = (inp[14]) ? node20991 : 4'b1111;
															assign node20991 = (inp[9]) ? node20993 : 4'b1010;
																assign node20993 = (inp[12]) ? 4'b1010 : 4'b1110;
														assign node20996 = (inp[14]) ? node21002 : node20997;
															assign node20997 = (inp[9]) ? 4'b1010 : node20998;
																assign node20998 = (inp[12]) ? 4'b1110 : 4'b1010;
															assign node21002 = (inp[12]) ? node21004 : 4'b1111;
																assign node21004 = (inp[9]) ? 4'b1011 : 4'b1111;
													assign node21007 = (inp[9]) ? node21011 : node21008;
														assign node21008 = (inp[12]) ? 4'b1111 : 4'b1011;
														assign node21011 = (inp[12]) ? node21015 : node21012;
															assign node21012 = (inp[8]) ? 4'b1111 : 4'b1110;
															assign node21015 = (inp[14]) ? 4'b1011 : 4'b1010;
												assign node21018 = (inp[9]) ? node21028 : node21019;
													assign node21019 = (inp[12]) ? node21025 : node21020;
														assign node21020 = (inp[14]) ? node21022 : 4'b1010;
															assign node21022 = (inp[7]) ? 4'b1011 : 4'b1010;
														assign node21025 = (inp[14]) ? 4'b1101 : 4'b1100;
													assign node21028 = (inp[12]) ? node21040 : node21029;
														assign node21029 = (inp[14]) ? node21035 : node21030;
															assign node21030 = (inp[7]) ? 4'b1100 : node21031;
																assign node21031 = (inp[8]) ? 4'b1100 : 4'b1101;
															assign node21035 = (inp[8]) ? 4'b1101 : node21036;
																assign node21036 = (inp[7]) ? 4'b1101 : 4'b1100;
														assign node21040 = (inp[14]) ? node21042 : 4'b1001;
															assign node21042 = (inp[8]) ? node21044 : 4'b1000;
																assign node21044 = (inp[7]) ? 4'b1000 : 4'b1001;
											assign node21047 = (inp[14]) ? node21093 : node21048;
												assign node21048 = (inp[3]) ? node21070 : node21049;
													assign node21049 = (inp[12]) ? node21063 : node21050;
														assign node21050 = (inp[9]) ? node21058 : node21051;
															assign node21051 = (inp[7]) ? node21055 : node21052;
																assign node21052 = (inp[8]) ? 4'b1010 : 4'b1011;
																assign node21055 = (inp[8]) ? 4'b1011 : 4'b1010;
															assign node21058 = (inp[8]) ? 4'b1100 : node21059;
																assign node21059 = (inp[7]) ? 4'b1100 : 4'b1101;
														assign node21063 = (inp[9]) ? 4'b1001 : node21064;
															assign node21064 = (inp[7]) ? node21066 : 4'b1101;
																assign node21066 = (inp[8]) ? 4'b1101 : 4'b1100;
													assign node21070 = (inp[7]) ? node21084 : node21071;
														assign node21071 = (inp[8]) ? node21079 : node21072;
															assign node21072 = (inp[9]) ? node21076 : node21073;
																assign node21073 = (inp[12]) ? 4'b1101 : 4'b1001;
																assign node21076 = (inp[12]) ? 4'b1001 : 4'b1101;
															assign node21079 = (inp[12]) ? node21081 : 4'b1100;
																assign node21081 = (inp[9]) ? 4'b1000 : 4'b1100;
														assign node21084 = (inp[8]) ? 4'b1001 : node21085;
															assign node21085 = (inp[12]) ? node21089 : node21086;
																assign node21086 = (inp[9]) ? 4'b1100 : 4'b1000;
																assign node21089 = (inp[9]) ? 4'b1000 : 4'b1100;
												assign node21093 = (inp[9]) ? node21107 : node21094;
													assign node21094 = (inp[12]) ? node21100 : node21095;
														assign node21095 = (inp[8]) ? 4'b1001 : node21096;
															assign node21096 = (inp[7]) ? 4'b1001 : 4'b1000;
														assign node21100 = (inp[7]) ? node21104 : node21101;
															assign node21101 = (inp[8]) ? 4'b1101 : 4'b1100;
															assign node21104 = (inp[8]) ? 4'b1100 : 4'b1101;
													assign node21107 = (inp[12]) ? node21115 : node21108;
														assign node21108 = (inp[7]) ? node21112 : node21109;
															assign node21109 = (inp[3]) ? 4'b1100 : 4'b1101;
															assign node21112 = (inp[8]) ? 4'b1100 : 4'b1101;
														assign node21115 = (inp[8]) ? node21117 : 4'b1001;
															assign node21117 = (inp[7]) ? 4'b1000 : 4'b1001;
										assign node21120 = (inp[3]) ? node21208 : node21121;
											assign node21121 = (inp[5]) ? node21169 : node21122;
												assign node21122 = (inp[7]) ? node21146 : node21123;
													assign node21123 = (inp[12]) ? node21135 : node21124;
														assign node21124 = (inp[9]) ? node21130 : node21125;
															assign node21125 = (inp[14]) ? node21127 : 4'b1001;
																assign node21127 = (inp[8]) ? 4'b1001 : 4'b1000;
															assign node21130 = (inp[8]) ? node21132 : 4'b1101;
																assign node21132 = (inp[14]) ? 4'b1101 : 4'b1100;
														assign node21135 = (inp[9]) ? node21143 : node21136;
															assign node21136 = (inp[14]) ? node21140 : node21137;
																assign node21137 = (inp[8]) ? 4'b1100 : 4'b1101;
																assign node21140 = (inp[8]) ? 4'b1101 : 4'b1100;
															assign node21143 = (inp[14]) ? 4'b1001 : 4'b1000;
													assign node21146 = (inp[14]) ? node21160 : node21147;
														assign node21147 = (inp[8]) ? node21155 : node21148;
															assign node21148 = (inp[9]) ? node21152 : node21149;
																assign node21149 = (inp[12]) ? 4'b1100 : 4'b1000;
																assign node21152 = (inp[12]) ? 4'b1000 : 4'b1100;
															assign node21155 = (inp[9]) ? 4'b1001 : node21156;
																assign node21156 = (inp[12]) ? 4'b1101 : 4'b1001;
														assign node21160 = (inp[8]) ? node21162 : 4'b1101;
															assign node21162 = (inp[9]) ? node21166 : node21163;
																assign node21163 = (inp[12]) ? 4'b1100 : 4'b1000;
																assign node21166 = (inp[12]) ? 4'b1000 : 4'b1100;
												assign node21169 = (inp[12]) ? node21187 : node21170;
													assign node21170 = (inp[9]) ? node21184 : node21171;
														assign node21171 = (inp[7]) ? node21177 : node21172;
															assign node21172 = (inp[8]) ? node21174 : 4'b1001;
																assign node21174 = (inp[14]) ? 4'b1001 : 4'b1000;
															assign node21177 = (inp[14]) ? node21181 : node21178;
																assign node21178 = (inp[8]) ? 4'b1001 : 4'b1000;
																assign node21181 = (inp[8]) ? 4'b1000 : 4'b1001;
														assign node21184 = (inp[8]) ? 4'b1110 : 4'b1111;
													assign node21187 = (inp[9]) ? node21195 : node21188;
														assign node21188 = (inp[14]) ? node21190 : 4'b1111;
															assign node21190 = (inp[7]) ? node21192 : 4'b1111;
																assign node21192 = (inp[8]) ? 4'b1110 : 4'b1111;
														assign node21195 = (inp[7]) ? node21201 : node21196;
															assign node21196 = (inp[8]) ? 4'b1010 : node21197;
																assign node21197 = (inp[14]) ? 4'b1010 : 4'b1011;
															assign node21201 = (inp[8]) ? node21205 : node21202;
																assign node21202 = (inp[14]) ? 4'b1011 : 4'b1010;
																assign node21205 = (inp[14]) ? 4'b1010 : 4'b1011;
											assign node21208 = (inp[9]) ? node21242 : node21209;
												assign node21209 = (inp[12]) ? node21227 : node21210;
													assign node21210 = (inp[5]) ? node21220 : node21211;
														assign node21211 = (inp[8]) ? 4'b1000 : node21212;
															assign node21212 = (inp[7]) ? node21216 : node21213;
																assign node21213 = (inp[14]) ? 4'b1000 : 4'b1001;
																assign node21216 = (inp[14]) ? 4'b1001 : 4'b1000;
														assign node21220 = (inp[14]) ? node21222 : 4'b1011;
															assign node21222 = (inp[7]) ? 4'b1010 : node21223;
																assign node21223 = (inp[8]) ? 4'b1011 : 4'b1010;
													assign node21227 = (inp[14]) ? node21229 : 4'b1111;
														assign node21229 = (inp[5]) ? node21235 : node21230;
															assign node21230 = (inp[8]) ? 4'b1111 : node21231;
																assign node21231 = (inp[7]) ? 4'b1111 : 4'b1110;
															assign node21235 = (inp[7]) ? node21239 : node21236;
																assign node21236 = (inp[8]) ? 4'b1111 : 4'b1110;
																assign node21239 = (inp[8]) ? 4'b1110 : 4'b1111;
												assign node21242 = (inp[12]) ? node21256 : node21243;
													assign node21243 = (inp[7]) ? node21249 : node21244;
														assign node21244 = (inp[8]) ? 4'b1111 : node21245;
															assign node21245 = (inp[14]) ? 4'b1110 : 4'b1111;
														assign node21249 = (inp[8]) ? node21253 : node21250;
															assign node21250 = (inp[14]) ? 4'b1111 : 4'b1110;
															assign node21253 = (inp[14]) ? 4'b1110 : 4'b1111;
													assign node21256 = (inp[5]) ? node21270 : node21257;
														assign node21257 = (inp[7]) ? node21263 : node21258;
															assign node21258 = (inp[8]) ? node21260 : 4'b1011;
																assign node21260 = (inp[14]) ? 4'b1011 : 4'b1010;
															assign node21263 = (inp[14]) ? node21267 : node21264;
																assign node21264 = (inp[8]) ? 4'b1011 : 4'b1010;
																assign node21267 = (inp[8]) ? 4'b1010 : 4'b1011;
														assign node21270 = (inp[14]) ? node21272 : 4'b1010;
															assign node21272 = (inp[7]) ? 4'b1010 : node21273;
																assign node21273 = (inp[8]) ? 4'b1011 : 4'b1010;
								assign node21277 = (inp[8]) ? node21623 : node21278;
									assign node21278 = (inp[3]) ? node21452 : node21279;
										assign node21279 = (inp[0]) ? node21357 : node21280;
											assign node21280 = (inp[5]) ? node21320 : node21281;
												assign node21281 = (inp[7]) ? node21305 : node21282;
													assign node21282 = (inp[14]) ? node21292 : node21283;
														assign node21283 = (inp[12]) ? node21285 : 4'b1101;
															assign node21285 = (inp[9]) ? node21289 : node21286;
																assign node21286 = (inp[4]) ? 4'b1101 : 4'b1001;
																assign node21289 = (inp[4]) ? 4'b1001 : 4'b1101;
														assign node21292 = (inp[4]) ? node21298 : node21293;
															assign node21293 = (inp[9]) ? 4'b1100 : node21294;
																assign node21294 = (inp[12]) ? 4'b1000 : 4'b1100;
															assign node21298 = (inp[12]) ? node21302 : node21299;
																assign node21299 = (inp[9]) ? 4'b1100 : 4'b1000;
																assign node21302 = (inp[9]) ? 4'b1000 : 4'b1100;
													assign node21305 = (inp[14]) ? node21315 : node21306;
														assign node21306 = (inp[4]) ? node21308 : 4'b1000;
															assign node21308 = (inp[9]) ? node21312 : node21309;
																assign node21309 = (inp[12]) ? 4'b1100 : 4'b1000;
																assign node21312 = (inp[12]) ? 4'b1000 : 4'b1100;
														assign node21315 = (inp[12]) ? 4'b1001 : node21316;
															assign node21316 = (inp[9]) ? 4'b1101 : 4'b1001;
												assign node21320 = (inp[12]) ? node21342 : node21321;
													assign node21321 = (inp[9]) ? node21333 : node21322;
														assign node21322 = (inp[4]) ? node21328 : node21323;
															assign node21323 = (inp[14]) ? 4'b1100 : node21324;
																assign node21324 = (inp[7]) ? 4'b1100 : 4'b1101;
															assign node21328 = (inp[7]) ? node21330 : 4'b1000;
																assign node21330 = (inp[14]) ? 4'b1001 : 4'b1000;
														assign node21333 = (inp[4]) ? node21335 : 4'b1001;
															assign node21335 = (inp[14]) ? node21339 : node21336;
																assign node21336 = (inp[7]) ? 4'b1110 : 4'b1111;
																assign node21339 = (inp[7]) ? 4'b1111 : 4'b1110;
													assign node21342 = (inp[9]) ? node21350 : node21343;
														assign node21343 = (inp[4]) ? node21345 : 4'b1001;
															assign node21345 = (inp[14]) ? node21347 : 4'b1111;
																assign node21347 = (inp[7]) ? 4'b1111 : 4'b1110;
														assign node21350 = (inp[4]) ? 4'b1010 : node21351;
															assign node21351 = (inp[14]) ? node21353 : 4'b1110;
																assign node21353 = (inp[7]) ? 4'b1111 : 4'b1110;
											assign node21357 = (inp[5]) ? node21405 : node21358;
												assign node21358 = (inp[14]) ? node21384 : node21359;
													assign node21359 = (inp[7]) ? node21371 : node21360;
														assign node21360 = (inp[9]) ? node21366 : node21361;
															assign node21361 = (inp[12]) ? node21363 : 4'b1111;
																assign node21363 = (inp[4]) ? 4'b1111 : 4'b1011;
															assign node21366 = (inp[4]) ? 4'b1011 : node21367;
																assign node21367 = (inp[12]) ? 4'b1111 : 4'b1011;
														assign node21371 = (inp[12]) ? node21377 : node21372;
															assign node21372 = (inp[4]) ? node21374 : 4'b1010;
																assign node21374 = (inp[9]) ? 4'b1110 : 4'b1010;
															assign node21377 = (inp[4]) ? node21381 : node21378;
																assign node21378 = (inp[9]) ? 4'b1110 : 4'b1010;
																assign node21381 = (inp[9]) ? 4'b1010 : 4'b1110;
													assign node21384 = (inp[7]) ? node21392 : node21385;
														assign node21385 = (inp[4]) ? node21387 : 4'b1110;
															assign node21387 = (inp[9]) ? 4'b1110 : node21388;
																assign node21388 = (inp[12]) ? 4'b1110 : 4'b1010;
														assign node21392 = (inp[12]) ? node21398 : node21393;
															assign node21393 = (inp[4]) ? 4'b1111 : node21394;
																assign node21394 = (inp[9]) ? 4'b1011 : 4'b1111;
															assign node21398 = (inp[4]) ? node21402 : node21399;
																assign node21399 = (inp[9]) ? 4'b1111 : 4'b1011;
																assign node21402 = (inp[9]) ? 4'b1011 : 4'b1111;
												assign node21405 = (inp[12]) ? node21431 : node21406;
													assign node21406 = (inp[4]) ? node21420 : node21407;
														assign node21407 = (inp[9]) ? node21415 : node21408;
															assign node21408 = (inp[7]) ? node21412 : node21409;
																assign node21409 = (inp[14]) ? 4'b1110 : 4'b1111;
																assign node21412 = (inp[14]) ? 4'b1111 : 4'b1110;
															assign node21415 = (inp[7]) ? 4'b1011 : node21416;
																assign node21416 = (inp[14]) ? 4'b1010 : 4'b1011;
														assign node21420 = (inp[9]) ? node21426 : node21421;
															assign node21421 = (inp[7]) ? node21423 : 4'b1011;
																assign node21423 = (inp[14]) ? 4'b1011 : 4'b1010;
															assign node21426 = (inp[14]) ? 4'b1100 : node21427;
																assign node21427 = (inp[7]) ? 4'b1100 : 4'b1101;
													assign node21431 = (inp[9]) ? node21443 : node21432;
														assign node21432 = (inp[4]) ? node21438 : node21433;
															assign node21433 = (inp[14]) ? 4'b1010 : node21434;
																assign node21434 = (inp[7]) ? 4'b1010 : 4'b1011;
															assign node21438 = (inp[14]) ? 4'b1100 : node21439;
																assign node21439 = (inp[7]) ? 4'b1100 : 4'b1101;
														assign node21443 = (inp[4]) ? node21449 : node21444;
															assign node21444 = (inp[7]) ? node21446 : 4'b1101;
																assign node21446 = (inp[14]) ? 4'b1101 : 4'b1100;
															assign node21449 = (inp[14]) ? 4'b1001 : 4'b1000;
										assign node21452 = (inp[0]) ? node21546 : node21453;
											assign node21453 = (inp[5]) ? node21499 : node21454;
												assign node21454 = (inp[4]) ? node21476 : node21455;
													assign node21455 = (inp[12]) ? node21463 : node21456;
														assign node21456 = (inp[9]) ? node21458 : 4'b1100;
															assign node21458 = (inp[7]) ? node21460 : 4'b1000;
																assign node21460 = (inp[14]) ? 4'b1001 : 4'b1000;
														assign node21463 = (inp[9]) ? node21469 : node21464;
															assign node21464 = (inp[7]) ? node21466 : 4'b1000;
																assign node21466 = (inp[14]) ? 4'b1001 : 4'b1000;
															assign node21469 = (inp[7]) ? node21473 : node21470;
																assign node21470 = (inp[14]) ? 4'b1110 : 4'b1111;
																assign node21473 = (inp[14]) ? 4'b1111 : 4'b1110;
													assign node21476 = (inp[9]) ? node21486 : node21477;
														assign node21477 = (inp[12]) ? node21481 : node21478;
															assign node21478 = (inp[7]) ? 4'b1001 : 4'b1000;
															assign node21481 = (inp[7]) ? 4'b1111 : node21482;
																assign node21482 = (inp[14]) ? 4'b1110 : 4'b1111;
														assign node21486 = (inp[12]) ? node21494 : node21487;
															assign node21487 = (inp[14]) ? node21491 : node21488;
																assign node21488 = (inp[7]) ? 4'b1110 : 4'b1111;
																assign node21491 = (inp[7]) ? 4'b1111 : 4'b1110;
															assign node21494 = (inp[14]) ? 4'b1010 : node21495;
																assign node21495 = (inp[7]) ? 4'b1010 : 4'b1011;
												assign node21499 = (inp[14]) ? node21521 : node21500;
													assign node21500 = (inp[7]) ? node21506 : node21501;
														assign node21501 = (inp[9]) ? node21503 : 4'b1111;
															assign node21503 = (inp[4]) ? 4'b1011 : 4'b1111;
														assign node21506 = (inp[4]) ? node21514 : node21507;
															assign node21507 = (inp[9]) ? node21511 : node21508;
																assign node21508 = (inp[12]) ? 4'b1010 : 4'b1110;
																assign node21511 = (inp[12]) ? 4'b1110 : 4'b1010;
															assign node21514 = (inp[12]) ? node21518 : node21515;
																assign node21515 = (inp[9]) ? 4'b1110 : 4'b1010;
																assign node21518 = (inp[9]) ? 4'b1010 : 4'b1110;
													assign node21521 = (inp[7]) ? node21535 : node21522;
														assign node21522 = (inp[4]) ? node21530 : node21523;
															assign node21523 = (inp[12]) ? node21527 : node21524;
																assign node21524 = (inp[9]) ? 4'b1010 : 4'b1110;
																assign node21527 = (inp[9]) ? 4'b1110 : 4'b1010;
															assign node21530 = (inp[12]) ? 4'b1010 : node21531;
																assign node21531 = (inp[9]) ? 4'b1110 : 4'b1010;
														assign node21535 = (inp[9]) ? node21541 : node21536;
															assign node21536 = (inp[12]) ? 4'b1111 : node21537;
																assign node21537 = (inp[4]) ? 4'b1011 : 4'b1111;
															assign node21541 = (inp[4]) ? node21543 : 4'b1011;
																assign node21543 = (inp[12]) ? 4'b1011 : 4'b1111;
											assign node21546 = (inp[5]) ? node21584 : node21547;
												assign node21547 = (inp[12]) ? node21571 : node21548;
													assign node21548 = (inp[9]) ? node21560 : node21549;
														assign node21549 = (inp[4]) ? node21555 : node21550;
															assign node21550 = (inp[14]) ? node21552 : 4'b1111;
																assign node21552 = (inp[7]) ? 4'b1111 : 4'b1110;
															assign node21555 = (inp[7]) ? 4'b1011 : node21556;
																assign node21556 = (inp[14]) ? 4'b1010 : 4'b1011;
														assign node21560 = (inp[4]) ? node21568 : node21561;
															assign node21561 = (inp[14]) ? node21565 : node21562;
																assign node21562 = (inp[7]) ? 4'b1010 : 4'b1011;
																assign node21565 = (inp[7]) ? 4'b1011 : 4'b1010;
															assign node21568 = (inp[7]) ? 4'b1101 : 4'b1100;
													assign node21571 = (inp[4]) ? node21579 : node21572;
														assign node21572 = (inp[9]) ? node21574 : 4'b1011;
															assign node21574 = (inp[14]) ? 4'b1101 : node21575;
																assign node21575 = (inp[7]) ? 4'b1100 : 4'b1101;
														assign node21579 = (inp[9]) ? node21581 : 4'b1100;
															assign node21581 = (inp[14]) ? 4'b1001 : 4'b1000;
												assign node21584 = (inp[9]) ? node21610 : node21585;
													assign node21585 = (inp[12]) ? node21597 : node21586;
														assign node21586 = (inp[4]) ? node21594 : node21587;
															assign node21587 = (inp[7]) ? node21591 : node21588;
																assign node21588 = (inp[14]) ? 4'b1100 : 4'b1101;
																assign node21591 = (inp[14]) ? 4'b1101 : 4'b1100;
															assign node21594 = (inp[7]) ? 4'b1000 : 4'b1001;
														assign node21597 = (inp[4]) ? node21605 : node21598;
															assign node21598 = (inp[7]) ? node21602 : node21599;
																assign node21599 = (inp[14]) ? 4'b1000 : 4'b1001;
																assign node21602 = (inp[14]) ? 4'b1001 : 4'b1000;
															assign node21605 = (inp[14]) ? node21607 : 4'b1100;
																assign node21607 = (inp[7]) ? 4'b1101 : 4'b1100;
													assign node21610 = (inp[7]) ? node21614 : node21611;
														assign node21611 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node21614 = (inp[14]) ? node21620 : node21615;
															assign node21615 = (inp[4]) ? node21617 : 4'b1000;
																assign node21617 = (inp[12]) ? 4'b1000 : 4'b1100;
															assign node21620 = (inp[4]) ? 4'b1101 : 4'b1001;
									assign node21623 = (inp[14]) ? node21751 : node21624;
										assign node21624 = (inp[7]) ? node21678 : node21625;
											assign node21625 = (inp[12]) ? node21657 : node21626;
												assign node21626 = (inp[0]) ? node21640 : node21627;
													assign node21627 = (inp[9]) ? node21631 : node21628;
														assign node21628 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node21631 = (inp[4]) ? node21635 : node21632;
															assign node21632 = (inp[5]) ? 4'b1010 : 4'b1000;
															assign node21635 = (inp[3]) ? 4'b1110 : node21636;
																assign node21636 = (inp[5]) ? 4'b1110 : 4'b1100;
													assign node21640 = (inp[5]) ? node21648 : node21641;
														assign node21641 = (inp[9]) ? node21645 : node21642;
															assign node21642 = (inp[4]) ? 4'b1010 : 4'b1110;
															assign node21645 = (inp[4]) ? 4'b1110 : 4'b1010;
														assign node21648 = (inp[3]) ? node21654 : node21649;
															assign node21649 = (inp[4]) ? node21651 : 4'b1010;
																assign node21651 = (inp[9]) ? 4'b1100 : 4'b1010;
															assign node21654 = (inp[4]) ? 4'b1000 : 4'b1100;
												assign node21657 = (inp[4]) ? node21667 : node21658;
													assign node21658 = (inp[9]) ? node21662 : node21659;
														assign node21659 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node21662 = (inp[3]) ? node21664 : 4'b1100;
															assign node21664 = (inp[5]) ? 4'b1110 : 4'b1100;
													assign node21667 = (inp[9]) ? node21669 : 4'b1100;
														assign node21669 = (inp[3]) ? node21675 : node21670;
															assign node21670 = (inp[0]) ? node21672 : 4'b1000;
																assign node21672 = (inp[5]) ? 4'b1000 : 4'b1010;
															assign node21675 = (inp[0]) ? 4'b1000 : 4'b1010;
											assign node21678 = (inp[4]) ? node21706 : node21679;
												assign node21679 = (inp[3]) ? node21697 : node21680;
													assign node21680 = (inp[0]) ? node21690 : node21681;
														assign node21681 = (inp[5]) ? node21683 : 4'b1101;
															assign node21683 = (inp[12]) ? node21687 : node21684;
																assign node21684 = (inp[9]) ? 4'b1001 : 4'b1101;
																assign node21687 = (inp[9]) ? 4'b1111 : 4'b1001;
														assign node21690 = (inp[5]) ? 4'b1011 : node21691;
															assign node21691 = (inp[12]) ? 4'b1111 : node21692;
																assign node21692 = (inp[9]) ? 4'b1011 : 4'b1111;
													assign node21697 = (inp[0]) ? 4'b1101 : node21698;
														assign node21698 = (inp[5]) ? 4'b1111 : node21699;
															assign node21699 = (inp[12]) ? 4'b1111 : node21700;
																assign node21700 = (inp[9]) ? 4'b1001 : 4'b1101;
												assign node21706 = (inp[0]) ? node21736 : node21707;
													assign node21707 = (inp[3]) ? node21723 : node21708;
														assign node21708 = (inp[5]) ? node21716 : node21709;
															assign node21709 = (inp[12]) ? node21713 : node21710;
																assign node21710 = (inp[9]) ? 4'b1101 : 4'b1001;
																assign node21713 = (inp[9]) ? 4'b1001 : 4'b1101;
															assign node21716 = (inp[9]) ? node21720 : node21717;
																assign node21717 = (inp[12]) ? 4'b1111 : 4'b1001;
																assign node21720 = (inp[12]) ? 4'b1011 : 4'b1111;
														assign node21723 = (inp[5]) ? node21729 : node21724;
															assign node21724 = (inp[9]) ? node21726 : 4'b1111;
																assign node21726 = (inp[12]) ? 4'b1011 : 4'b1111;
															assign node21729 = (inp[9]) ? node21733 : node21730;
																assign node21730 = (inp[12]) ? 4'b1111 : 4'b1011;
																assign node21733 = (inp[12]) ? 4'b1011 : 4'b1111;
													assign node21736 = (inp[9]) ? node21744 : node21737;
														assign node21737 = (inp[12]) ? node21739 : 4'b1011;
															assign node21739 = (inp[3]) ? 4'b1101 : node21740;
																assign node21740 = (inp[5]) ? 4'b1101 : 4'b1111;
														assign node21744 = (inp[12]) ? 4'b1001 : node21745;
															assign node21745 = (inp[5]) ? 4'b1101 : node21746;
																assign node21746 = (inp[3]) ? 4'b1101 : 4'b1111;
										assign node21751 = (inp[7]) ? node21821 : node21752;
											assign node21752 = (inp[12]) ? node21788 : node21753;
												assign node21753 = (inp[9]) ? node21771 : node21754;
													assign node21754 = (inp[4]) ? node21762 : node21755;
														assign node21755 = (inp[3]) ? node21757 : 4'b1111;
															assign node21757 = (inp[0]) ? 4'b1101 : node21758;
																assign node21758 = (inp[5]) ? 4'b1111 : 4'b1101;
														assign node21762 = (inp[5]) ? node21766 : node21763;
															assign node21763 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node21766 = (inp[0]) ? 4'b1001 : node21767;
																assign node21767 = (inp[3]) ? 4'b1011 : 4'b1001;
													assign node21771 = (inp[4]) ? node21777 : node21772;
														assign node21772 = (inp[5]) ? 4'b1011 : node21773;
															assign node21773 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node21777 = (inp[0]) ? node21783 : node21778;
															assign node21778 = (inp[3]) ? 4'b1111 : node21779;
																assign node21779 = (inp[5]) ? 4'b1111 : 4'b1101;
															assign node21783 = (inp[5]) ? 4'b1101 : node21784;
																assign node21784 = (inp[3]) ? 4'b1101 : 4'b1111;
												assign node21788 = (inp[5]) ? node21808 : node21789;
													assign node21789 = (inp[3]) ? node21799 : node21790;
														assign node21790 = (inp[0]) ? 4'b1111 : node21791;
															assign node21791 = (inp[4]) ? node21795 : node21792;
																assign node21792 = (inp[9]) ? 4'b1101 : 4'b1001;
																assign node21795 = (inp[9]) ? 4'b1001 : 4'b1101;
														assign node21799 = (inp[4]) ? node21805 : node21800;
															assign node21800 = (inp[9]) ? 4'b1111 : node21801;
																assign node21801 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node21805 = (inp[0]) ? 4'b1001 : 4'b1011;
													assign node21808 = (inp[0]) ? node21816 : node21809;
														assign node21809 = (inp[4]) ? node21813 : node21810;
															assign node21810 = (inp[3]) ? 4'b1011 : 4'b1001;
															assign node21813 = (inp[9]) ? 4'b1011 : 4'b1111;
														assign node21816 = (inp[3]) ? 4'b1101 : node21817;
															assign node21817 = (inp[9]) ? 4'b1001 : 4'b1011;
											assign node21821 = (inp[9]) ? node21857 : node21822;
												assign node21822 = (inp[0]) ? node21844 : node21823;
													assign node21823 = (inp[3]) ? node21833 : node21824;
														assign node21824 = (inp[4]) ? node21828 : node21825;
															assign node21825 = (inp[12]) ? 4'b1000 : 4'b1100;
															assign node21828 = (inp[12]) ? node21830 : 4'b1000;
																assign node21830 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node21833 = (inp[5]) ? node21839 : node21834;
															assign node21834 = (inp[4]) ? node21836 : 4'b1000;
																assign node21836 = (inp[12]) ? 4'b1110 : 4'b1000;
															assign node21839 = (inp[12]) ? node21841 : 4'b1110;
																assign node21841 = (inp[4]) ? 4'b1110 : 4'b1010;
													assign node21844 = (inp[4]) ? node21848 : node21845;
														assign node21845 = (inp[12]) ? 4'b1010 : 4'b1110;
														assign node21848 = (inp[12]) ? node21852 : node21849;
															assign node21849 = (inp[3]) ? 4'b1000 : 4'b1010;
															assign node21852 = (inp[5]) ? 4'b1100 : node21853;
																assign node21853 = (inp[3]) ? 4'b1100 : 4'b1110;
												assign node21857 = (inp[0]) ? node21877 : node21858;
													assign node21858 = (inp[3]) ? node21870 : node21859;
														assign node21859 = (inp[5]) ? node21863 : node21860;
															assign node21860 = (inp[12]) ? 4'b1100 : 4'b1000;
															assign node21863 = (inp[4]) ? node21867 : node21864;
																assign node21864 = (inp[12]) ? 4'b1110 : 4'b1000;
																assign node21867 = (inp[12]) ? 4'b1010 : 4'b1110;
														assign node21870 = (inp[5]) ? 4'b1010 : node21871;
															assign node21871 = (inp[4]) ? node21873 : 4'b1110;
																assign node21873 = (inp[12]) ? 4'b1010 : 4'b1110;
													assign node21877 = (inp[4]) ? node21885 : node21878;
														assign node21878 = (inp[12]) ? 4'b1100 : node21879;
															assign node21879 = (inp[3]) ? node21881 : 4'b1010;
																assign node21881 = (inp[5]) ? 4'b1000 : 4'b1010;
														assign node21885 = (inp[12]) ? 4'b1000 : 4'b1100;
							assign node21888 = (inp[9]) ? node22304 : node21889;
								assign node21889 = (inp[4]) ? node22117 : node21890;
									assign node21890 = (inp[12]) ? node22006 : node21891;
										assign node21891 = (inp[15]) ? node21957 : node21892;
											assign node21892 = (inp[0]) ? node21926 : node21893;
												assign node21893 = (inp[3]) ? node21911 : node21894;
													assign node21894 = (inp[14]) ? node21902 : node21895;
														assign node21895 = (inp[7]) ? node21899 : node21896;
															assign node21896 = (inp[8]) ? 4'b1111 : 4'b1110;
															assign node21899 = (inp[8]) ? 4'b1110 : 4'b1111;
														assign node21902 = (inp[5]) ? node21904 : 4'b1111;
															assign node21904 = (inp[7]) ? node21908 : node21905;
																assign node21905 = (inp[8]) ? 4'b1111 : 4'b1110;
																assign node21908 = (inp[8]) ? 4'b1110 : 4'b1111;
													assign node21911 = (inp[5]) ? node21919 : node21912;
														assign node21912 = (inp[7]) ? node21916 : node21913;
															assign node21913 = (inp[8]) ? 4'b1111 : 4'b1110;
															assign node21916 = (inp[14]) ? 4'b1110 : 4'b1111;
														assign node21919 = (inp[14]) ? node21921 : 4'b1101;
															assign node21921 = (inp[8]) ? node21923 : 4'b1100;
																assign node21923 = (inp[7]) ? 4'b1100 : 4'b1101;
												assign node21926 = (inp[5]) ? node21944 : node21927;
													assign node21927 = (inp[14]) ? node21937 : node21928;
														assign node21928 = (inp[3]) ? node21932 : node21929;
															assign node21929 = (inp[8]) ? 4'b1100 : 4'b1101;
															assign node21932 = (inp[7]) ? 4'b1101 : node21933;
																assign node21933 = (inp[8]) ? 4'b1101 : 4'b1100;
														assign node21937 = (inp[7]) ? node21941 : node21938;
															assign node21938 = (inp[8]) ? 4'b1101 : 4'b1100;
															assign node21941 = (inp[8]) ? 4'b1100 : 4'b1101;
													assign node21944 = (inp[3]) ? node21950 : node21945;
														assign node21945 = (inp[7]) ? node21947 : 4'b1101;
															assign node21947 = (inp[8]) ? 4'b1100 : 4'b1101;
														assign node21950 = (inp[8]) ? node21954 : node21951;
															assign node21951 = (inp[7]) ? 4'b1111 : 4'b1110;
															assign node21954 = (inp[7]) ? 4'b1110 : 4'b1111;
											assign node21957 = (inp[0]) ? node21987 : node21958;
												assign node21958 = (inp[3]) ? node21974 : node21959;
													assign node21959 = (inp[14]) ? node21967 : node21960;
														assign node21960 = (inp[5]) ? node21962 : 4'b1100;
															assign node21962 = (inp[7]) ? node21964 : 4'b1100;
																assign node21964 = (inp[8]) ? 4'b1100 : 4'b1101;
														assign node21967 = (inp[7]) ? node21971 : node21968;
															assign node21968 = (inp[8]) ? 4'b1101 : 4'b1100;
															assign node21971 = (inp[8]) ? 4'b1100 : 4'b1101;
													assign node21974 = (inp[5]) ? node21980 : node21975;
														assign node21975 = (inp[8]) ? node21977 : 4'b1101;
															assign node21977 = (inp[14]) ? 4'b1100 : 4'b1101;
														assign node21980 = (inp[8]) ? node21984 : node21981;
															assign node21981 = (inp[7]) ? 4'b1111 : 4'b1110;
															assign node21984 = (inp[7]) ? 4'b1110 : 4'b1111;
												assign node21987 = (inp[3]) ? node21999 : node21988;
													assign node21988 = (inp[5]) ? node21994 : node21989;
														assign node21989 = (inp[8]) ? node21991 : 4'b1110;
															assign node21991 = (inp[7]) ? 4'b1110 : 4'b1111;
														assign node21994 = (inp[8]) ? 4'b1111 : node21995;
															assign node21995 = (inp[7]) ? 4'b1111 : 4'b1110;
													assign node21999 = (inp[5]) ? 4'b1100 : node22000;
														assign node22000 = (inp[7]) ? 4'b1110 : node22001;
															assign node22001 = (inp[14]) ? 4'b1111 : 4'b1110;
										assign node22006 = (inp[5]) ? node22044 : node22007;
											assign node22007 = (inp[0]) ? node22029 : node22008;
												assign node22008 = (inp[15]) ? node22022 : node22009;
													assign node22009 = (inp[3]) ? node22017 : node22010;
														assign node22010 = (inp[8]) ? node22014 : node22011;
															assign node22011 = (inp[7]) ? 4'b1011 : 4'b1010;
															assign node22014 = (inp[7]) ? 4'b1010 : 4'b1011;
														assign node22017 = (inp[7]) ? 4'b1010 : node22018;
															assign node22018 = (inp[8]) ? 4'b1011 : 4'b1010;
													assign node22022 = (inp[8]) ? node22026 : node22023;
														assign node22023 = (inp[7]) ? 4'b1001 : 4'b1000;
														assign node22026 = (inp[7]) ? 4'b1000 : 4'b1001;
												assign node22029 = (inp[15]) ? node22037 : node22030;
													assign node22030 = (inp[8]) ? node22034 : node22031;
														assign node22031 = (inp[7]) ? 4'b1001 : 4'b1000;
														assign node22034 = (inp[7]) ? 4'b1000 : 4'b1001;
													assign node22037 = (inp[7]) ? node22041 : node22038;
														assign node22038 = (inp[8]) ? 4'b1011 : 4'b1010;
														assign node22041 = (inp[8]) ? 4'b1010 : 4'b1011;
											assign node22044 = (inp[0]) ? node22084 : node22045;
												assign node22045 = (inp[14]) ? node22065 : node22046;
													assign node22046 = (inp[7]) ? node22054 : node22047;
														assign node22047 = (inp[8]) ? node22049 : 4'b1010;
															assign node22049 = (inp[3]) ? node22051 : 4'b1011;
																assign node22051 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node22054 = (inp[8]) ? node22060 : node22055;
															assign node22055 = (inp[3]) ? 4'b1011 : node22056;
																assign node22056 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node22060 = (inp[3]) ? node22062 : 4'b1010;
																assign node22062 = (inp[15]) ? 4'b1010 : 4'b1000;
													assign node22065 = (inp[3]) ? node22077 : node22066;
														assign node22066 = (inp[15]) ? node22070 : node22067;
															assign node22067 = (inp[7]) ? 4'b1011 : 4'b1010;
															assign node22070 = (inp[8]) ? node22074 : node22071;
																assign node22071 = (inp[7]) ? 4'b1001 : 4'b1000;
																assign node22074 = (inp[7]) ? 4'b1000 : 4'b1001;
														assign node22077 = (inp[15]) ? 4'b1011 : node22078;
															assign node22078 = (inp[7]) ? node22080 : 4'b1001;
																assign node22080 = (inp[8]) ? 4'b1000 : 4'b1001;
												assign node22084 = (inp[3]) ? node22104 : node22085;
													assign node22085 = (inp[15]) ? node22099 : node22086;
														assign node22086 = (inp[14]) ? node22092 : node22087;
															assign node22087 = (inp[8]) ? 4'b1001 : node22088;
																assign node22088 = (inp[7]) ? 4'b1001 : 4'b1000;
															assign node22092 = (inp[8]) ? node22096 : node22093;
																assign node22093 = (inp[7]) ? 4'b1001 : 4'b1000;
																assign node22096 = (inp[7]) ? 4'b1000 : 4'b1001;
														assign node22099 = (inp[8]) ? node22101 : 4'b1011;
															assign node22101 = (inp[7]) ? 4'b1010 : 4'b1011;
													assign node22104 = (inp[15]) ? node22110 : node22105;
														assign node22105 = (inp[14]) ? 4'b1011 : node22106;
															assign node22106 = (inp[7]) ? 4'b1011 : 4'b1010;
														assign node22110 = (inp[7]) ? node22114 : node22111;
															assign node22111 = (inp[8]) ? 4'b1001 : 4'b1000;
															assign node22114 = (inp[8]) ? 4'b1000 : 4'b1001;
									assign node22117 = (inp[12]) ? node22203 : node22118;
										assign node22118 = (inp[7]) ? node22160 : node22119;
											assign node22119 = (inp[8]) ? node22137 : node22120;
												assign node22120 = (inp[3]) ? node22128 : node22121;
													assign node22121 = (inp[15]) ? node22125 : node22122;
														assign node22122 = (inp[0]) ? 4'b1000 : 4'b1010;
														assign node22125 = (inp[0]) ? 4'b1010 : 4'b1000;
													assign node22128 = (inp[5]) ? node22130 : 4'b1000;
														assign node22130 = (inp[0]) ? node22134 : node22131;
															assign node22131 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node22134 = (inp[15]) ? 4'b1000 : 4'b1010;
												assign node22137 = (inp[3]) ? node22145 : node22138;
													assign node22138 = (inp[15]) ? node22142 : node22139;
														assign node22139 = (inp[0]) ? 4'b1001 : 4'b1011;
														assign node22142 = (inp[0]) ? 4'b1011 : 4'b1001;
													assign node22145 = (inp[15]) ? node22153 : node22146;
														assign node22146 = (inp[0]) ? node22150 : node22147;
															assign node22147 = (inp[5]) ? 4'b1001 : 4'b1011;
															assign node22150 = (inp[5]) ? 4'b1011 : 4'b1001;
														assign node22153 = (inp[0]) ? node22157 : node22154;
															assign node22154 = (inp[5]) ? 4'b1011 : 4'b1001;
															assign node22157 = (inp[5]) ? 4'b1001 : 4'b1011;
											assign node22160 = (inp[8]) ? node22182 : node22161;
												assign node22161 = (inp[0]) ? node22173 : node22162;
													assign node22162 = (inp[15]) ? node22168 : node22163;
														assign node22163 = (inp[5]) ? node22165 : 4'b1011;
															assign node22165 = (inp[3]) ? 4'b1001 : 4'b1011;
														assign node22168 = (inp[3]) ? node22170 : 4'b1001;
															assign node22170 = (inp[5]) ? 4'b1011 : 4'b1001;
													assign node22173 = (inp[15]) ? node22179 : node22174;
														assign node22174 = (inp[5]) ? node22176 : 4'b1001;
															assign node22176 = (inp[3]) ? 4'b1011 : 4'b1001;
														assign node22179 = (inp[5]) ? 4'b1001 : 4'b1011;
												assign node22182 = (inp[0]) ? node22192 : node22183;
													assign node22183 = (inp[15]) ? node22187 : node22184;
														assign node22184 = (inp[3]) ? 4'b1000 : 4'b1010;
														assign node22187 = (inp[5]) ? node22189 : 4'b1000;
															assign node22189 = (inp[3]) ? 4'b1010 : 4'b1000;
													assign node22192 = (inp[15]) ? node22198 : node22193;
														assign node22193 = (inp[3]) ? node22195 : 4'b1000;
															assign node22195 = (inp[5]) ? 4'b1010 : 4'b1000;
														assign node22198 = (inp[5]) ? node22200 : 4'b1010;
															assign node22200 = (inp[3]) ? 4'b1000 : 4'b1010;
										assign node22203 = (inp[14]) ? node22253 : node22204;
											assign node22204 = (inp[15]) ? node22224 : node22205;
												assign node22205 = (inp[0]) ? node22213 : node22206;
													assign node22206 = (inp[8]) ? node22210 : node22207;
														assign node22207 = (inp[7]) ? 4'b1101 : 4'b1100;
														assign node22210 = (inp[7]) ? 4'b1100 : 4'b1101;
													assign node22213 = (inp[5]) ? node22215 : 4'b1101;
														assign node22215 = (inp[3]) ? 4'b1111 : node22216;
															assign node22216 = (inp[7]) ? node22220 : node22217;
																assign node22217 = (inp[8]) ? 4'b1111 : 4'b1110;
																assign node22220 = (inp[8]) ? 4'b1110 : 4'b1111;
												assign node22224 = (inp[0]) ? node22244 : node22225;
													assign node22225 = (inp[5]) ? node22239 : node22226;
														assign node22226 = (inp[3]) ? node22234 : node22227;
															assign node22227 = (inp[8]) ? node22231 : node22228;
																assign node22228 = (inp[7]) ? 4'b1101 : 4'b1100;
																assign node22231 = (inp[7]) ? 4'b1100 : 4'b1101;
															assign node22234 = (inp[7]) ? node22236 : 4'b1110;
																assign node22236 = (inp[8]) ? 4'b1110 : 4'b1111;
														assign node22239 = (inp[8]) ? node22241 : 4'b1111;
															assign node22241 = (inp[7]) ? 4'b1110 : 4'b1111;
													assign node22244 = (inp[5]) ? node22246 : 4'b1110;
														assign node22246 = (inp[8]) ? node22250 : node22247;
															assign node22247 = (inp[7]) ? 4'b1101 : 4'b1100;
															assign node22250 = (inp[7]) ? 4'b1100 : 4'b1101;
											assign node22253 = (inp[7]) ? node22281 : node22254;
												assign node22254 = (inp[8]) ? node22270 : node22255;
													assign node22255 = (inp[5]) ? node22263 : node22256;
														assign node22256 = (inp[15]) ? 4'b1110 : node22257;
															assign node22257 = (inp[3]) ? node22259 : 4'b1110;
																assign node22259 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node22263 = (inp[0]) ? node22267 : node22264;
															assign node22264 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node22267 = (inp[15]) ? 4'b1100 : 4'b1110;
													assign node22270 = (inp[0]) ? node22278 : node22271;
														assign node22271 = (inp[3]) ? 4'b1111 : node22272;
															assign node22272 = (inp[5]) ? 4'b1111 : node22273;
																assign node22273 = (inp[15]) ? 4'b1101 : 4'b1111;
														assign node22278 = (inp[5]) ? 4'b1101 : 4'b1111;
												assign node22281 = (inp[8]) ? node22293 : node22282;
													assign node22282 = (inp[3]) ? node22286 : node22283;
														assign node22283 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node22286 = (inp[15]) ? node22290 : node22287;
															assign node22287 = (inp[5]) ? 4'b1111 : 4'b1101;
															assign node22290 = (inp[0]) ? 4'b1101 : 4'b1111;
													assign node22293 = (inp[15]) ? node22295 : 4'b1100;
														assign node22295 = (inp[5]) ? node22301 : node22296;
															assign node22296 = (inp[0]) ? 4'b1110 : node22297;
																assign node22297 = (inp[3]) ? 4'b1110 : 4'b1100;
															assign node22301 = (inp[0]) ? 4'b1100 : 4'b1110;
								assign node22304 = (inp[15]) ? node22544 : node22305;
									assign node22305 = (inp[0]) ? node22407 : node22306;
										assign node22306 = (inp[3]) ? node22370 : node22307;
											assign node22307 = (inp[5]) ? node22333 : node22308;
												assign node22308 = (inp[4]) ? node22322 : node22309;
													assign node22309 = (inp[12]) ? node22315 : node22310;
														assign node22310 = (inp[14]) ? 4'b1011 : node22311;
															assign node22311 = (inp[8]) ? 4'b1010 : 4'b1011;
														assign node22315 = (inp[14]) ? 4'b1111 : node22316;
															assign node22316 = (inp[7]) ? node22318 : 4'b1110;
																assign node22318 = (inp[8]) ? 4'b1110 : 4'b1111;
													assign node22322 = (inp[12]) ? node22328 : node22323;
														assign node22323 = (inp[8]) ? 4'b1110 : node22324;
															assign node22324 = (inp[7]) ? 4'b1111 : 4'b1110;
														assign node22328 = (inp[7]) ? node22330 : 4'b1010;
															assign node22330 = (inp[8]) ? 4'b1010 : 4'b1011;
												assign node22333 = (inp[12]) ? node22355 : node22334;
													assign node22334 = (inp[4]) ? node22348 : node22335;
														assign node22335 = (inp[14]) ? node22343 : node22336;
															assign node22336 = (inp[8]) ? node22340 : node22337;
																assign node22337 = (inp[7]) ? 4'b1011 : 4'b1010;
																assign node22340 = (inp[7]) ? 4'b1010 : 4'b1011;
															assign node22343 = (inp[7]) ? node22345 : 4'b1010;
																assign node22345 = (inp[8]) ? 4'b1010 : 4'b1011;
														assign node22348 = (inp[8]) ? node22352 : node22349;
															assign node22349 = (inp[7]) ? 4'b1101 : 4'b1100;
															assign node22352 = (inp[14]) ? 4'b1100 : 4'b1101;
													assign node22355 = (inp[4]) ? node22363 : node22356;
														assign node22356 = (inp[8]) ? node22360 : node22357;
															assign node22357 = (inp[7]) ? 4'b1101 : 4'b1100;
															assign node22360 = (inp[7]) ? 4'b1100 : 4'b1101;
														assign node22363 = (inp[8]) ? node22367 : node22364;
															assign node22364 = (inp[7]) ? 4'b1001 : 4'b1000;
															assign node22367 = (inp[7]) ? 4'b1000 : 4'b1001;
											assign node22370 = (inp[4]) ? node22386 : node22371;
												assign node22371 = (inp[12]) ? node22379 : node22372;
													assign node22372 = (inp[5]) ? node22374 : 4'b1010;
														assign node22374 = (inp[8]) ? node22376 : 4'b1001;
															assign node22376 = (inp[7]) ? 4'b1000 : 4'b1001;
													assign node22379 = (inp[7]) ? node22383 : node22380;
														assign node22380 = (inp[8]) ? 4'b1101 : 4'b1100;
														assign node22383 = (inp[8]) ? 4'b1100 : 4'b1101;
												assign node22386 = (inp[12]) ? node22394 : node22387;
													assign node22387 = (inp[7]) ? node22391 : node22388;
														assign node22388 = (inp[8]) ? 4'b1101 : 4'b1100;
														assign node22391 = (inp[8]) ? 4'b1100 : 4'b1101;
													assign node22394 = (inp[14]) ? node22400 : node22395;
														assign node22395 = (inp[8]) ? node22397 : 4'b1000;
															assign node22397 = (inp[7]) ? 4'b1000 : 4'b1001;
														assign node22400 = (inp[7]) ? node22404 : node22401;
															assign node22401 = (inp[8]) ? 4'b1001 : 4'b1000;
															assign node22404 = (inp[8]) ? 4'b1000 : 4'b1001;
										assign node22407 = (inp[3]) ? node22467 : node22408;
											assign node22408 = (inp[5]) ? node22436 : node22409;
												assign node22409 = (inp[4]) ? node22425 : node22410;
													assign node22410 = (inp[12]) ? 4'b1100 : node22411;
														assign node22411 = (inp[14]) ? node22419 : node22412;
															assign node22412 = (inp[8]) ? node22416 : node22413;
																assign node22413 = (inp[7]) ? 4'b1001 : 4'b1000;
																assign node22416 = (inp[7]) ? 4'b1000 : 4'b1001;
															assign node22419 = (inp[8]) ? 4'b1000 : node22420;
																assign node22420 = (inp[7]) ? 4'b1001 : 4'b1000;
													assign node22425 = (inp[12]) ? node22433 : node22426;
														assign node22426 = (inp[7]) ? node22430 : node22427;
															assign node22427 = (inp[8]) ? 4'b1101 : 4'b1100;
															assign node22430 = (inp[8]) ? 4'b1100 : 4'b1101;
														assign node22433 = (inp[8]) ? 4'b1001 : 4'b1000;
												assign node22436 = (inp[12]) ? node22452 : node22437;
													assign node22437 = (inp[4]) ? node22447 : node22438;
														assign node22438 = (inp[14]) ? node22444 : node22439;
															assign node22439 = (inp[8]) ? 4'b1000 : node22440;
																assign node22440 = (inp[7]) ? 4'b1001 : 4'b1000;
															assign node22444 = (inp[7]) ? 4'b1000 : 4'b1001;
														assign node22447 = (inp[8]) ? node22449 : 4'b1110;
															assign node22449 = (inp[7]) ? 4'b1110 : 4'b1111;
													assign node22452 = (inp[4]) ? node22464 : node22453;
														assign node22453 = (inp[14]) ? node22459 : node22454;
															assign node22454 = (inp[7]) ? node22456 : 4'b1111;
																assign node22456 = (inp[8]) ? 4'b1110 : 4'b1111;
															assign node22459 = (inp[8]) ? 4'b1110 : node22460;
																assign node22460 = (inp[7]) ? 4'b1111 : 4'b1110;
														assign node22464 = (inp[7]) ? 4'b1010 : 4'b1011;
											assign node22467 = (inp[5]) ? node22495 : node22468;
												assign node22468 = (inp[12]) ? node22480 : node22469;
													assign node22469 = (inp[4]) ? node22475 : node22470;
														assign node22470 = (inp[8]) ? node22472 : 4'b1000;
															assign node22472 = (inp[7]) ? 4'b1000 : 4'b1001;
														assign node22475 = (inp[8]) ? node22477 : 4'b1111;
															assign node22477 = (inp[7]) ? 4'b1110 : 4'b1111;
													assign node22480 = (inp[4]) ? node22488 : node22481;
														assign node22481 = (inp[8]) ? node22485 : node22482;
															assign node22482 = (inp[7]) ? 4'b1111 : 4'b1110;
															assign node22485 = (inp[7]) ? 4'b1110 : 4'b1111;
														assign node22488 = (inp[14]) ? node22490 : 4'b1010;
															assign node22490 = (inp[7]) ? 4'b1011 : node22491;
																assign node22491 = (inp[8]) ? 4'b1011 : 4'b1010;
												assign node22495 = (inp[14]) ? node22519 : node22496;
													assign node22496 = (inp[12]) ? node22510 : node22497;
														assign node22497 = (inp[4]) ? node22505 : node22498;
															assign node22498 = (inp[7]) ? node22502 : node22499;
																assign node22499 = (inp[8]) ? 4'b1011 : 4'b1010;
																assign node22502 = (inp[8]) ? 4'b1010 : 4'b1011;
															assign node22505 = (inp[8]) ? 4'b1111 : node22506;
																assign node22506 = (inp[7]) ? 4'b1111 : 4'b1110;
														assign node22510 = (inp[4]) ? node22512 : 4'b1110;
															assign node22512 = (inp[7]) ? node22516 : node22513;
																assign node22513 = (inp[8]) ? 4'b1011 : 4'b1010;
																assign node22516 = (inp[8]) ? 4'b1010 : 4'b1011;
													assign node22519 = (inp[4]) ? node22533 : node22520;
														assign node22520 = (inp[12]) ? node22526 : node22521;
															assign node22521 = (inp[7]) ? node22523 : 4'b1010;
																assign node22523 = (inp[8]) ? 4'b1010 : 4'b1011;
															assign node22526 = (inp[8]) ? node22530 : node22527;
																assign node22527 = (inp[7]) ? 4'b1111 : 4'b1110;
																assign node22530 = (inp[7]) ? 4'b1110 : 4'b1111;
														assign node22533 = (inp[12]) ? node22539 : node22534;
															assign node22534 = (inp[7]) ? node22536 : 4'b1111;
																assign node22536 = (inp[8]) ? 4'b1110 : 4'b1111;
															assign node22539 = (inp[7]) ? node22541 : 4'b1011;
																assign node22541 = (inp[8]) ? 4'b1010 : 4'b1011;
									assign node22544 = (inp[0]) ? node22662 : node22545;
										assign node22545 = (inp[5]) ? node22599 : node22546;
											assign node22546 = (inp[3]) ? node22578 : node22547;
												assign node22547 = (inp[14]) ? node22567 : node22548;
													assign node22548 = (inp[12]) ? node22558 : node22549;
														assign node22549 = (inp[4]) ? 4'b1101 : node22550;
															assign node22550 = (inp[8]) ? node22554 : node22551;
																assign node22551 = (inp[7]) ? 4'b1001 : 4'b1000;
																assign node22554 = (inp[7]) ? 4'b1000 : 4'b1001;
														assign node22558 = (inp[4]) ? node22560 : 4'b1101;
															assign node22560 = (inp[8]) ? node22564 : node22561;
																assign node22561 = (inp[7]) ? 4'b1001 : 4'b1000;
																assign node22564 = (inp[7]) ? 4'b1000 : 4'b1001;
													assign node22567 = (inp[4]) ? node22575 : node22568;
														assign node22568 = (inp[12]) ? node22570 : 4'b1000;
															assign node22570 = (inp[8]) ? 4'b1101 : node22571;
																assign node22571 = (inp[7]) ? 4'b1101 : 4'b1100;
														assign node22575 = (inp[12]) ? 4'b1000 : 4'b1100;
												assign node22578 = (inp[4]) ? node22590 : node22579;
													assign node22579 = (inp[12]) ? node22587 : node22580;
														assign node22580 = (inp[8]) ? node22584 : node22581;
															assign node22581 = (inp[7]) ? 4'b1001 : 4'b1000;
															assign node22584 = (inp[7]) ? 4'b1000 : 4'b1001;
														assign node22587 = (inp[8]) ? 4'b1111 : 4'b1110;
													assign node22590 = (inp[12]) ? node22592 : 4'b1110;
														assign node22592 = (inp[7]) ? node22596 : node22593;
															assign node22593 = (inp[8]) ? 4'b1011 : 4'b1010;
															assign node22596 = (inp[8]) ? 4'b1010 : 4'b1011;
											assign node22599 = (inp[4]) ? node22635 : node22600;
												assign node22600 = (inp[12]) ? node22624 : node22601;
													assign node22601 = (inp[3]) ? node22613 : node22602;
														assign node22602 = (inp[14]) ? node22608 : node22603;
															assign node22603 = (inp[8]) ? 4'b1001 : node22604;
																assign node22604 = (inp[7]) ? 4'b1001 : 4'b1000;
															assign node22608 = (inp[8]) ? 4'b1000 : node22609;
																assign node22609 = (inp[7]) ? 4'b1001 : 4'b1000;
														assign node22613 = (inp[14]) ? node22619 : node22614;
															assign node22614 = (inp[8]) ? 4'b1011 : node22615;
																assign node22615 = (inp[7]) ? 4'b1011 : 4'b1010;
															assign node22619 = (inp[8]) ? node22621 : 4'b1010;
																assign node22621 = (inp[7]) ? 4'b1010 : 4'b1011;
													assign node22624 = (inp[14]) ? node22630 : node22625;
														assign node22625 = (inp[3]) ? node22627 : 4'b1110;
															assign node22627 = (inp[8]) ? 4'b1110 : 4'b1111;
														assign node22630 = (inp[7]) ? 4'b1111 : node22631;
															assign node22631 = (inp[8]) ? 4'b1111 : 4'b1110;
												assign node22635 = (inp[12]) ? node22643 : node22636;
													assign node22636 = (inp[8]) ? node22640 : node22637;
														assign node22637 = (inp[7]) ? 4'b1111 : 4'b1110;
														assign node22640 = (inp[7]) ? 4'b1110 : 4'b1111;
													assign node22643 = (inp[3]) ? node22657 : node22644;
														assign node22644 = (inp[14]) ? node22650 : node22645;
															assign node22645 = (inp[7]) ? node22647 : 4'b1011;
																assign node22647 = (inp[8]) ? 4'b1010 : 4'b1011;
															assign node22650 = (inp[7]) ? node22654 : node22651;
																assign node22651 = (inp[8]) ? 4'b1011 : 4'b1010;
																assign node22654 = (inp[8]) ? 4'b1010 : 4'b1011;
														assign node22657 = (inp[7]) ? 4'b1011 : node22658;
															assign node22658 = (inp[8]) ? 4'b1011 : 4'b1010;
										assign node22662 = (inp[5]) ? node22726 : node22663;
											assign node22663 = (inp[3]) ? node22697 : node22664;
												assign node22664 = (inp[4]) ? node22684 : node22665;
													assign node22665 = (inp[12]) ? node22671 : node22666;
														assign node22666 = (inp[8]) ? node22668 : 4'b1010;
															assign node22668 = (inp[7]) ? 4'b1010 : 4'b1011;
														assign node22671 = (inp[14]) ? node22679 : node22672;
															assign node22672 = (inp[7]) ? node22676 : node22673;
																assign node22673 = (inp[8]) ? 4'b1111 : 4'b1110;
																assign node22676 = (inp[8]) ? 4'b1110 : 4'b1111;
															assign node22679 = (inp[8]) ? node22681 : 4'b1111;
																assign node22681 = (inp[7]) ? 4'b1110 : 4'b1111;
													assign node22684 = (inp[12]) ? node22686 : 4'b1111;
														assign node22686 = (inp[14]) ? node22692 : node22687;
															assign node22687 = (inp[8]) ? node22689 : 4'b1011;
																assign node22689 = (inp[7]) ? 4'b1010 : 4'b1011;
															assign node22692 = (inp[7]) ? 4'b1010 : node22693;
																assign node22693 = (inp[8]) ? 4'b1011 : 4'b1010;
												assign node22697 = (inp[4]) ? node22711 : node22698;
													assign node22698 = (inp[12]) ? node22706 : node22699;
														assign node22699 = (inp[8]) ? node22703 : node22700;
															assign node22700 = (inp[7]) ? 4'b1011 : 4'b1010;
															assign node22703 = (inp[7]) ? 4'b1010 : 4'b1011;
														assign node22706 = (inp[7]) ? node22708 : 4'b1101;
															assign node22708 = (inp[8]) ? 4'b1100 : 4'b1101;
													assign node22711 = (inp[12]) ? node22719 : node22712;
														assign node22712 = (inp[7]) ? node22716 : node22713;
															assign node22713 = (inp[8]) ? 4'b1101 : 4'b1100;
															assign node22716 = (inp[8]) ? 4'b1100 : 4'b1101;
														assign node22719 = (inp[14]) ? node22721 : 4'b1001;
															assign node22721 = (inp[7]) ? node22723 : 4'b1000;
																assign node22723 = (inp[8]) ? 4'b1000 : 4'b1001;
											assign node22726 = (inp[3]) ? node22760 : node22727;
												assign node22727 = (inp[4]) ? node22745 : node22728;
													assign node22728 = (inp[12]) ? node22738 : node22729;
														assign node22729 = (inp[14]) ? 4'b1011 : node22730;
															assign node22730 = (inp[8]) ? node22734 : node22731;
																assign node22731 = (inp[7]) ? 4'b1011 : 4'b1010;
																assign node22734 = (inp[7]) ? 4'b1010 : 4'b1011;
														assign node22738 = (inp[7]) ? node22742 : node22739;
															assign node22739 = (inp[8]) ? 4'b1101 : 4'b1100;
															assign node22742 = (inp[8]) ? 4'b1100 : 4'b1101;
													assign node22745 = (inp[12]) ? node22751 : node22746;
														assign node22746 = (inp[7]) ? node22748 : 4'b1100;
															assign node22748 = (inp[14]) ? 4'b1101 : 4'b1100;
														assign node22751 = (inp[14]) ? node22753 : 4'b1000;
															assign node22753 = (inp[7]) ? node22757 : node22754;
																assign node22754 = (inp[8]) ? 4'b1001 : 4'b1000;
																assign node22757 = (inp[8]) ? 4'b1000 : 4'b1001;
												assign node22760 = (inp[7]) ? node22782 : node22761;
													assign node22761 = (inp[8]) ? node22769 : node22762;
														assign node22762 = (inp[4]) ? node22766 : node22763;
															assign node22763 = (inp[12]) ? 4'b1100 : 4'b1000;
															assign node22766 = (inp[12]) ? 4'b1000 : 4'b1100;
														assign node22769 = (inp[14]) ? node22775 : node22770;
															assign node22770 = (inp[12]) ? node22772 : 4'b1001;
																assign node22772 = (inp[4]) ? 4'b1001 : 4'b1101;
															assign node22775 = (inp[12]) ? node22779 : node22776;
																assign node22776 = (inp[4]) ? 4'b1101 : 4'b1001;
																assign node22779 = (inp[4]) ? 4'b1001 : 4'b1101;
													assign node22782 = (inp[8]) ? node22784 : 4'b1001;
														assign node22784 = (inp[14]) ? node22790 : node22785;
															assign node22785 = (inp[4]) ? 4'b1000 : node22786;
																assign node22786 = (inp[12]) ? 4'b1100 : 4'b1000;
															assign node22790 = (inp[12]) ? node22794 : node22791;
																assign node22791 = (inp[4]) ? 4'b1100 : 4'b1000;
																assign node22794 = (inp[4]) ? 4'b1000 : 4'b1100;
				assign node22797 = (inp[1]) ? node27015 : node22798;
					assign node22798 = (inp[13]) ? node24998 : node22799;
						assign node22799 = (inp[5]) ? node23985 : node22800;
							assign node22800 = (inp[2]) ? node23462 : node22801;
								assign node22801 = (inp[7]) ? node23127 : node22802;
									assign node22802 = (inp[0]) ? node22962 : node22803;
										assign node22803 = (inp[15]) ? node22881 : node22804;
											assign node22804 = (inp[3]) ? node22844 : node22805;
												assign node22805 = (inp[8]) ? node22827 : node22806;
													assign node22806 = (inp[14]) ? node22820 : node22807;
														assign node22807 = (inp[9]) ? node22815 : node22808;
															assign node22808 = (inp[4]) ? node22812 : node22809;
																assign node22809 = (inp[12]) ? 4'b1011 : 4'b1111;
																assign node22812 = (inp[12]) ? 4'b1111 : 4'b1011;
															assign node22815 = (inp[12]) ? 4'b1111 : node22816;
																assign node22816 = (inp[4]) ? 4'b1111 : 4'b1011;
														assign node22820 = (inp[12]) ? 4'b1110 : node22821;
															assign node22821 = (inp[4]) ? node22823 : 4'b1010;
																assign node22823 = (inp[9]) ? 4'b1110 : 4'b1010;
													assign node22827 = (inp[14]) ? node22837 : node22828;
														assign node22828 = (inp[4]) ? 4'b1010 : node22829;
															assign node22829 = (inp[12]) ? node22833 : node22830;
																assign node22830 = (inp[9]) ? 4'b1010 : 4'b1110;
																assign node22833 = (inp[9]) ? 4'b1110 : 4'b1010;
														assign node22837 = (inp[9]) ? node22841 : node22838;
															assign node22838 = (inp[12]) ? 4'b1011 : 4'b1111;
															assign node22841 = (inp[12]) ? 4'b1111 : 4'b1011;
												assign node22844 = (inp[9]) ? node22864 : node22845;
													assign node22845 = (inp[4]) ? node22857 : node22846;
														assign node22846 = (inp[12]) ? node22850 : node22847;
															assign node22847 = (inp[14]) ? 4'b1110 : 4'b1111;
															assign node22850 = (inp[14]) ? node22854 : node22851;
																assign node22851 = (inp[8]) ? 4'b1010 : 4'b1011;
																assign node22854 = (inp[8]) ? 4'b1011 : 4'b1010;
														assign node22857 = (inp[12]) ? node22859 : 4'b1010;
															assign node22859 = (inp[8]) ? node22861 : 4'b1101;
																assign node22861 = (inp[14]) ? 4'b1101 : 4'b1100;
													assign node22864 = (inp[4]) ? node22874 : node22865;
														assign node22865 = (inp[12]) ? node22867 : 4'b1011;
															assign node22867 = (inp[8]) ? node22871 : node22868;
																assign node22868 = (inp[14]) ? 4'b1100 : 4'b1101;
																assign node22871 = (inp[14]) ? 4'b1101 : 4'b1100;
														assign node22874 = (inp[12]) ? node22876 : 4'b1100;
															assign node22876 = (inp[8]) ? 4'b1000 : node22877;
																assign node22877 = (inp[14]) ? 4'b1000 : 4'b1001;
											assign node22881 = (inp[3]) ? node22925 : node22882;
												assign node22882 = (inp[4]) ? node22902 : node22883;
													assign node22883 = (inp[8]) ? node22893 : node22884;
														assign node22884 = (inp[14]) ? node22886 : 4'b1101;
															assign node22886 = (inp[12]) ? node22890 : node22887;
																assign node22887 = (inp[9]) ? 4'b1000 : 4'b1100;
																assign node22890 = (inp[9]) ? 4'b1100 : 4'b1000;
														assign node22893 = (inp[14]) ? 4'b1001 : node22894;
															assign node22894 = (inp[12]) ? node22898 : node22895;
																assign node22895 = (inp[9]) ? 4'b1000 : 4'b1100;
																assign node22898 = (inp[9]) ? 4'b1100 : 4'b1000;
													assign node22902 = (inp[9]) ? node22918 : node22903;
														assign node22903 = (inp[12]) ? node22911 : node22904;
															assign node22904 = (inp[14]) ? node22908 : node22905;
																assign node22905 = (inp[8]) ? 4'b1000 : 4'b1001;
																assign node22908 = (inp[8]) ? 4'b1001 : 4'b1000;
															assign node22911 = (inp[8]) ? node22915 : node22912;
																assign node22912 = (inp[14]) ? 4'b1100 : 4'b1101;
																assign node22915 = (inp[14]) ? 4'b1101 : 4'b1100;
														assign node22918 = (inp[12]) ? node22920 : 4'b1101;
															assign node22920 = (inp[8]) ? 4'b1001 : node22921;
																assign node22921 = (inp[14]) ? 4'b1000 : 4'b1001;
												assign node22925 = (inp[4]) ? node22941 : node22926;
													assign node22926 = (inp[12]) ? node22938 : node22927;
														assign node22927 = (inp[9]) ? node22933 : node22928;
															assign node22928 = (inp[14]) ? 4'b1100 : node22929;
																assign node22929 = (inp[8]) ? 4'b1100 : 4'b1101;
															assign node22933 = (inp[14]) ? 4'b1001 : node22934;
																assign node22934 = (inp[8]) ? 4'b1000 : 4'b1001;
														assign node22938 = (inp[9]) ? 4'b1111 : 4'b1001;
													assign node22941 = (inp[12]) ? node22951 : node22942;
														assign node22942 = (inp[9]) ? node22944 : 4'b1001;
															assign node22944 = (inp[14]) ? node22948 : node22945;
																assign node22945 = (inp[8]) ? 4'b1110 : 4'b1111;
																assign node22948 = (inp[8]) ? 4'b1111 : 4'b1110;
														assign node22951 = (inp[9]) ? node22955 : node22952;
															assign node22952 = (inp[14]) ? 4'b1111 : 4'b1110;
															assign node22955 = (inp[14]) ? node22959 : node22956;
																assign node22956 = (inp[8]) ? 4'b1010 : 4'b1011;
																assign node22959 = (inp[8]) ? 4'b1011 : 4'b1010;
										assign node22962 = (inp[15]) ? node23058 : node22963;
											assign node22963 = (inp[3]) ? node23007 : node22964;
												assign node22964 = (inp[4]) ? node22984 : node22965;
													assign node22965 = (inp[9]) ? node22973 : node22966;
														assign node22966 = (inp[12]) ? node22968 : 4'b1100;
															assign node22968 = (inp[14]) ? node22970 : 4'b1001;
																assign node22970 = (inp[8]) ? 4'b1001 : 4'b1000;
														assign node22973 = (inp[12]) ? node22979 : node22974;
															assign node22974 = (inp[8]) ? node22976 : 4'b1001;
																assign node22976 = (inp[14]) ? 4'b1001 : 4'b1000;
															assign node22979 = (inp[14]) ? 4'b1101 : node22980;
																assign node22980 = (inp[8]) ? 4'b1100 : 4'b1101;
													assign node22984 = (inp[9]) ? node22994 : node22985;
														assign node22985 = (inp[12]) ? node22987 : 4'b1001;
															assign node22987 = (inp[14]) ? node22991 : node22988;
																assign node22988 = (inp[8]) ? 4'b1100 : 4'b1101;
																assign node22991 = (inp[8]) ? 4'b1101 : 4'b1100;
														assign node22994 = (inp[12]) ? node23002 : node22995;
															assign node22995 = (inp[14]) ? node22999 : node22996;
																assign node22996 = (inp[8]) ? 4'b1100 : 4'b1101;
																assign node22999 = (inp[8]) ? 4'b1101 : 4'b1100;
															assign node23002 = (inp[8]) ? node23004 : 4'b1000;
																assign node23004 = (inp[14]) ? 4'b1001 : 4'b1000;
												assign node23007 = (inp[9]) ? node23033 : node23008;
													assign node23008 = (inp[12]) ? node23018 : node23009;
														assign node23009 = (inp[4]) ? node23011 : 4'b1100;
															assign node23011 = (inp[8]) ? node23015 : node23012;
																assign node23012 = (inp[14]) ? 4'b1000 : 4'b1001;
																assign node23015 = (inp[14]) ? 4'b1001 : 4'b1000;
														assign node23018 = (inp[4]) ? node23026 : node23019;
															assign node23019 = (inp[8]) ? node23023 : node23020;
																assign node23020 = (inp[14]) ? 4'b1000 : 4'b1001;
																assign node23023 = (inp[14]) ? 4'b1001 : 4'b1000;
															assign node23026 = (inp[8]) ? node23030 : node23027;
																assign node23027 = (inp[14]) ? 4'b1110 : 4'b1111;
																assign node23030 = (inp[14]) ? 4'b1111 : 4'b1110;
													assign node23033 = (inp[4]) ? node23047 : node23034;
														assign node23034 = (inp[12]) ? node23040 : node23035;
															assign node23035 = (inp[14]) ? node23037 : 4'b1000;
																assign node23037 = (inp[8]) ? 4'b1001 : 4'b1000;
															assign node23040 = (inp[8]) ? node23044 : node23041;
																assign node23041 = (inp[14]) ? 4'b1110 : 4'b1111;
																assign node23044 = (inp[14]) ? 4'b1111 : 4'b1110;
														assign node23047 = (inp[12]) ? node23055 : node23048;
															assign node23048 = (inp[8]) ? node23052 : node23049;
																assign node23049 = (inp[14]) ? 4'b1110 : 4'b1111;
																assign node23052 = (inp[14]) ? 4'b1111 : 4'b1110;
															assign node23055 = (inp[8]) ? 4'b1011 : 4'b1010;
											assign node23058 = (inp[3]) ? node23092 : node23059;
												assign node23059 = (inp[4]) ? node23071 : node23060;
													assign node23060 = (inp[8]) ? node23064 : node23061;
														assign node23061 = (inp[14]) ? 4'b1110 : 4'b1111;
														assign node23064 = (inp[14]) ? 4'b1111 : node23065;
															assign node23065 = (inp[9]) ? 4'b1110 : node23066;
																assign node23066 = (inp[12]) ? 4'b1010 : 4'b1110;
													assign node23071 = (inp[12]) ? node23083 : node23072;
														assign node23072 = (inp[9]) ? node23076 : node23073;
															assign node23073 = (inp[14]) ? 4'b1011 : 4'b1010;
															assign node23076 = (inp[14]) ? node23080 : node23077;
																assign node23077 = (inp[8]) ? 4'b1110 : 4'b1111;
																assign node23080 = (inp[8]) ? 4'b1111 : 4'b1110;
														assign node23083 = (inp[9]) ? node23087 : node23084;
															assign node23084 = (inp[14]) ? 4'b1111 : 4'b1110;
															assign node23087 = (inp[14]) ? 4'b1010 : node23088;
																assign node23088 = (inp[8]) ? 4'b1010 : 4'b1011;
												assign node23092 = (inp[4]) ? node23112 : node23093;
													assign node23093 = (inp[12]) ? node23107 : node23094;
														assign node23094 = (inp[9]) ? node23102 : node23095;
															assign node23095 = (inp[8]) ? node23099 : node23096;
																assign node23096 = (inp[14]) ? 4'b1110 : 4'b1111;
																assign node23099 = (inp[14]) ? 4'b1111 : 4'b1110;
															assign node23102 = (inp[14]) ? node23104 : 4'b1010;
																assign node23104 = (inp[8]) ? 4'b1011 : 4'b1010;
														assign node23107 = (inp[9]) ? node23109 : 4'b1011;
															assign node23109 = (inp[8]) ? 4'b1101 : 4'b1100;
													assign node23112 = (inp[8]) ? node23124 : node23113;
														assign node23113 = (inp[14]) ? node23119 : node23114;
															assign node23114 = (inp[9]) ? node23116 : 4'b1101;
																assign node23116 = (inp[12]) ? 4'b1001 : 4'b1101;
															assign node23119 = (inp[12]) ? 4'b1100 : node23120;
																assign node23120 = (inp[9]) ? 4'b1100 : 4'b1010;
														assign node23124 = (inp[14]) ? 4'b1101 : 4'b1100;
									assign node23127 = (inp[14]) ? node23289 : node23128;
										assign node23128 = (inp[8]) ? node23210 : node23129;
											assign node23129 = (inp[12]) ? node23177 : node23130;
												assign node23130 = (inp[3]) ? node23154 : node23131;
													assign node23131 = (inp[9]) ? node23143 : node23132;
														assign node23132 = (inp[4]) ? node23138 : node23133;
															assign node23133 = (inp[15]) ? node23135 : 4'b1110;
																assign node23135 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node23138 = (inp[0]) ? 4'b1010 : node23139;
																assign node23139 = (inp[15]) ? 4'b1000 : 4'b1010;
														assign node23143 = (inp[4]) ? node23149 : node23144;
															assign node23144 = (inp[15]) ? 4'b1010 : node23145;
																assign node23145 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node23149 = (inp[0]) ? node23151 : 4'b1110;
																assign node23151 = (inp[15]) ? 4'b1110 : 4'b1100;
													assign node23154 = (inp[15]) ? node23166 : node23155;
														assign node23155 = (inp[0]) ? node23161 : node23156;
															assign node23156 = (inp[4]) ? node23158 : 4'b1010;
																assign node23158 = (inp[9]) ? 4'b1100 : 4'b1010;
															assign node23161 = (inp[4]) ? 4'b1000 : node23162;
																assign node23162 = (inp[9]) ? 4'b1000 : 4'b1100;
														assign node23166 = (inp[0]) ? node23172 : node23167;
															assign node23167 = (inp[4]) ? node23169 : 4'b1000;
																assign node23169 = (inp[9]) ? 4'b1110 : 4'b1000;
															assign node23172 = (inp[4]) ? 4'b1010 : node23173;
																assign node23173 = (inp[9]) ? 4'b1010 : 4'b1110;
												assign node23177 = (inp[0]) ? node23191 : node23178;
													assign node23178 = (inp[9]) ? node23184 : node23179;
														assign node23179 = (inp[4]) ? 4'b1100 : node23180;
															assign node23180 = (inp[15]) ? 4'b1000 : 4'b1010;
														assign node23184 = (inp[4]) ? node23186 : 4'b1110;
															assign node23186 = (inp[15]) ? node23188 : 4'b1000;
																assign node23188 = (inp[3]) ? 4'b1010 : 4'b1000;
													assign node23191 = (inp[3]) ? node23199 : node23192;
														assign node23192 = (inp[15]) ? node23194 : 4'b1000;
															assign node23194 = (inp[9]) ? 4'b1010 : node23195;
																assign node23195 = (inp[4]) ? 4'b1110 : 4'b1010;
														assign node23199 = (inp[15]) ? node23207 : node23200;
															assign node23200 = (inp[9]) ? node23204 : node23201;
																assign node23201 = (inp[4]) ? 4'b1110 : 4'b1000;
																assign node23204 = (inp[4]) ? 4'b1010 : 4'b1110;
															assign node23207 = (inp[4]) ? 4'b1000 : 4'b1100;
											assign node23210 = (inp[0]) ? node23250 : node23211;
												assign node23211 = (inp[15]) ? node23231 : node23212;
													assign node23212 = (inp[3]) ? node23220 : node23213;
														assign node23213 = (inp[4]) ? node23215 : 4'b1111;
															assign node23215 = (inp[12]) ? node23217 : 4'b1011;
																assign node23217 = (inp[9]) ? 4'b1011 : 4'b1111;
														assign node23220 = (inp[12]) ? node23228 : node23221;
															assign node23221 = (inp[4]) ? node23225 : node23222;
																assign node23222 = (inp[9]) ? 4'b1011 : 4'b1111;
																assign node23225 = (inp[9]) ? 4'b1101 : 4'b1011;
															assign node23228 = (inp[4]) ? 4'b1001 : 4'b1101;
													assign node23231 = (inp[3]) ? node23237 : node23232;
														assign node23232 = (inp[4]) ? node23234 : 4'b1101;
															assign node23234 = (inp[9]) ? 4'b1101 : 4'b1001;
														assign node23237 = (inp[4]) ? node23243 : node23238;
															assign node23238 = (inp[12]) ? 4'b1001 : node23239;
																assign node23239 = (inp[9]) ? 4'b1001 : 4'b1101;
															assign node23243 = (inp[9]) ? node23247 : node23244;
																assign node23244 = (inp[12]) ? 4'b1111 : 4'b1001;
																assign node23247 = (inp[12]) ? 4'b1011 : 4'b1111;
												assign node23250 = (inp[15]) ? node23268 : node23251;
													assign node23251 = (inp[3]) ? node23261 : node23252;
														assign node23252 = (inp[9]) ? 4'b1001 : node23253;
															assign node23253 = (inp[4]) ? node23257 : node23254;
																assign node23254 = (inp[12]) ? 4'b1001 : 4'b1101;
																assign node23257 = (inp[12]) ? 4'b1101 : 4'b1001;
														assign node23261 = (inp[4]) ? node23263 : 4'b1001;
															assign node23263 = (inp[9]) ? node23265 : 4'b1001;
																assign node23265 = (inp[12]) ? 4'b1011 : 4'b1111;
													assign node23268 = (inp[3]) ? node23282 : node23269;
														assign node23269 = (inp[12]) ? node23275 : node23270;
															assign node23270 = (inp[4]) ? 4'b1011 : node23271;
																assign node23271 = (inp[9]) ? 4'b1011 : 4'b1111;
															assign node23275 = (inp[9]) ? node23279 : node23276;
																assign node23276 = (inp[4]) ? 4'b1111 : 4'b1011;
																assign node23279 = (inp[4]) ? 4'b1011 : 4'b1111;
														assign node23282 = (inp[12]) ? node23286 : node23283;
															assign node23283 = (inp[4]) ? 4'b1101 : 4'b1011;
															assign node23286 = (inp[4]) ? 4'b1001 : 4'b1101;
										assign node23289 = (inp[8]) ? node23377 : node23290;
											assign node23290 = (inp[4]) ? node23334 : node23291;
												assign node23291 = (inp[3]) ? node23315 : node23292;
													assign node23292 = (inp[0]) ? node23302 : node23293;
														assign node23293 = (inp[15]) ? 4'b1001 : node23294;
															assign node23294 = (inp[9]) ? node23298 : node23295;
																assign node23295 = (inp[12]) ? 4'b1011 : 4'b1111;
																assign node23298 = (inp[12]) ? 4'b1111 : 4'b1011;
														assign node23302 = (inp[15]) ? node23310 : node23303;
															assign node23303 = (inp[9]) ? node23307 : node23304;
																assign node23304 = (inp[12]) ? 4'b1001 : 4'b1101;
																assign node23307 = (inp[12]) ? 4'b1101 : 4'b1001;
															assign node23310 = (inp[12]) ? node23312 : 4'b1111;
																assign node23312 = (inp[9]) ? 4'b1111 : 4'b1011;
													assign node23315 = (inp[15]) ? node23321 : node23316;
														assign node23316 = (inp[9]) ? 4'b1101 : node23317;
															assign node23317 = (inp[0]) ? 4'b1101 : 4'b1111;
														assign node23321 = (inp[0]) ? node23329 : node23322;
															assign node23322 = (inp[9]) ? node23326 : node23323;
																assign node23323 = (inp[12]) ? 4'b1001 : 4'b1101;
																assign node23326 = (inp[12]) ? 4'b1111 : 4'b1001;
															assign node23329 = (inp[9]) ? 4'b1101 : node23330;
																assign node23330 = (inp[12]) ? 4'b1011 : 4'b1111;
												assign node23334 = (inp[0]) ? node23352 : node23335;
													assign node23335 = (inp[3]) ? node23343 : node23336;
														assign node23336 = (inp[15]) ? node23338 : 4'b1111;
															assign node23338 = (inp[9]) ? 4'b1001 : node23339;
																assign node23339 = (inp[12]) ? 4'b1101 : 4'b1001;
														assign node23343 = (inp[15]) ? node23347 : node23344;
															assign node23344 = (inp[12]) ? 4'b1001 : 4'b1011;
															assign node23347 = (inp[9]) ? node23349 : 4'b1001;
																assign node23349 = (inp[12]) ? 4'b1011 : 4'b1111;
													assign node23352 = (inp[15]) ? node23364 : node23353;
														assign node23353 = (inp[3]) ? node23361 : node23354;
															assign node23354 = (inp[9]) ? node23358 : node23355;
																assign node23355 = (inp[12]) ? 4'b1101 : 4'b1001;
																assign node23358 = (inp[12]) ? 4'b1001 : 4'b1101;
															assign node23361 = (inp[9]) ? 4'b1111 : 4'b1001;
														assign node23364 = (inp[3]) ? node23372 : node23365;
															assign node23365 = (inp[12]) ? node23369 : node23366;
																assign node23366 = (inp[9]) ? 4'b1111 : 4'b1011;
																assign node23369 = (inp[9]) ? 4'b1011 : 4'b1111;
															assign node23372 = (inp[12]) ? node23374 : 4'b1101;
																assign node23374 = (inp[9]) ? 4'b1001 : 4'b1101;
											assign node23377 = (inp[15]) ? node23421 : node23378;
												assign node23378 = (inp[0]) ? node23404 : node23379;
													assign node23379 = (inp[4]) ? node23393 : node23380;
														assign node23380 = (inp[3]) ? node23388 : node23381;
															assign node23381 = (inp[12]) ? node23385 : node23382;
																assign node23382 = (inp[9]) ? 4'b1010 : 4'b1110;
																assign node23385 = (inp[9]) ? 4'b1110 : 4'b1010;
															assign node23388 = (inp[12]) ? 4'b1010 : node23389;
																assign node23389 = (inp[9]) ? 4'b1010 : 4'b1110;
														assign node23393 = (inp[3]) ? node23397 : node23394;
															assign node23394 = (inp[9]) ? 4'b1010 : 4'b1110;
															assign node23397 = (inp[9]) ? node23401 : node23398;
																assign node23398 = (inp[12]) ? 4'b1100 : 4'b1010;
																assign node23401 = (inp[12]) ? 4'b1000 : 4'b1100;
													assign node23404 = (inp[3]) ? node23412 : node23405;
														assign node23405 = (inp[9]) ? node23407 : 4'b1000;
															assign node23407 = (inp[12]) ? 4'b1100 : node23408;
																assign node23408 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node23412 = (inp[4]) ? node23416 : node23413;
															assign node23413 = (inp[12]) ? 4'b1110 : 4'b1100;
															assign node23416 = (inp[12]) ? node23418 : 4'b1110;
																assign node23418 = (inp[9]) ? 4'b1010 : 4'b1110;
												assign node23421 = (inp[0]) ? node23447 : node23422;
													assign node23422 = (inp[3]) ? node23436 : node23423;
														assign node23423 = (inp[12]) ? node23429 : node23424;
															assign node23424 = (inp[4]) ? 4'b1000 : node23425;
																assign node23425 = (inp[9]) ? 4'b1000 : 4'b1100;
															assign node23429 = (inp[9]) ? node23433 : node23430;
																assign node23430 = (inp[4]) ? 4'b1100 : 4'b1000;
																assign node23433 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node23436 = (inp[12]) ? node23442 : node23437;
															assign node23437 = (inp[4]) ? 4'b1000 : node23438;
																assign node23438 = (inp[9]) ? 4'b1000 : 4'b1100;
															assign node23442 = (inp[9]) ? node23444 : 4'b1110;
																assign node23444 = (inp[4]) ? 4'b1010 : 4'b1110;
													assign node23447 = (inp[3]) ? node23455 : node23448;
														assign node23448 = (inp[12]) ? node23450 : 4'b1110;
															assign node23450 = (inp[9]) ? node23452 : 4'b1010;
																assign node23452 = (inp[4]) ? 4'b1010 : 4'b1110;
														assign node23455 = (inp[9]) ? 4'b1100 : node23456;
															assign node23456 = (inp[12]) ? node23458 : 4'b1010;
																assign node23458 = (inp[4]) ? 4'b1100 : 4'b1010;
								assign node23462 = (inp[0]) ? node23706 : node23463;
									assign node23463 = (inp[15]) ? node23603 : node23464;
										assign node23464 = (inp[3]) ? node23520 : node23465;
											assign node23465 = (inp[4]) ? node23495 : node23466;
												assign node23466 = (inp[7]) ? node23482 : node23467;
													assign node23467 = (inp[8]) ? node23475 : node23468;
														assign node23468 = (inp[12]) ? node23472 : node23469;
															assign node23469 = (inp[9]) ? 4'b1010 : 4'b1110;
															assign node23472 = (inp[9]) ? 4'b1110 : 4'b1010;
														assign node23475 = (inp[9]) ? node23479 : node23476;
															assign node23476 = (inp[12]) ? 4'b1011 : 4'b1111;
															assign node23479 = (inp[12]) ? 4'b1111 : 4'b1011;
													assign node23482 = (inp[8]) ? node23488 : node23483;
														assign node23483 = (inp[9]) ? 4'b1111 : node23484;
															assign node23484 = (inp[12]) ? 4'b1011 : 4'b1111;
														assign node23488 = (inp[12]) ? node23492 : node23489;
															assign node23489 = (inp[9]) ? 4'b1010 : 4'b1110;
															assign node23492 = (inp[9]) ? 4'b1110 : 4'b1010;
												assign node23495 = (inp[12]) ? node23507 : node23496;
													assign node23496 = (inp[9]) ? node23502 : node23497;
														assign node23497 = (inp[7]) ? 4'b1011 : node23498;
															assign node23498 = (inp[8]) ? 4'b1011 : 4'b1010;
														assign node23502 = (inp[7]) ? 4'b1111 : node23503;
															assign node23503 = (inp[8]) ? 4'b1111 : 4'b1110;
													assign node23507 = (inp[9]) ? node23515 : node23508;
														assign node23508 = (inp[8]) ? node23512 : node23509;
															assign node23509 = (inp[7]) ? 4'b1111 : 4'b1110;
															assign node23512 = (inp[7]) ? 4'b1110 : 4'b1111;
														assign node23515 = (inp[7]) ? node23517 : 4'b1011;
															assign node23517 = (inp[8]) ? 4'b1010 : 4'b1011;
											assign node23520 = (inp[4]) ? node23562 : node23521;
												assign node23521 = (inp[12]) ? node23541 : node23522;
													assign node23522 = (inp[9]) ? node23530 : node23523;
														assign node23523 = (inp[8]) ? node23527 : node23524;
															assign node23524 = (inp[7]) ? 4'b1111 : 4'b1110;
															assign node23527 = (inp[7]) ? 4'b1110 : 4'b1111;
														assign node23530 = (inp[14]) ? node23536 : node23531;
															assign node23531 = (inp[7]) ? 4'b1010 : node23532;
																assign node23532 = (inp[8]) ? 4'b1011 : 4'b1010;
															assign node23536 = (inp[8]) ? 4'b1011 : node23537;
																assign node23537 = (inp[7]) ? 4'b1011 : 4'b1010;
													assign node23541 = (inp[9]) ? node23549 : node23542;
														assign node23542 = (inp[7]) ? node23546 : node23543;
															assign node23543 = (inp[8]) ? 4'b1011 : 4'b1010;
															assign node23546 = (inp[8]) ? 4'b1010 : 4'b1011;
														assign node23549 = (inp[14]) ? node23557 : node23550;
															assign node23550 = (inp[8]) ? node23554 : node23551;
																assign node23551 = (inp[7]) ? 4'b1101 : 4'b1100;
																assign node23554 = (inp[7]) ? 4'b1100 : 4'b1101;
															assign node23557 = (inp[8]) ? 4'b1100 : node23558;
																assign node23558 = (inp[7]) ? 4'b1101 : 4'b1100;
												assign node23562 = (inp[12]) ? node23582 : node23563;
													assign node23563 = (inp[9]) ? node23571 : node23564;
														assign node23564 = (inp[14]) ? node23566 : 4'b1011;
															assign node23566 = (inp[8]) ? 4'b1010 : node23567;
																assign node23567 = (inp[7]) ? 4'b1011 : 4'b1010;
														assign node23571 = (inp[14]) ? node23577 : node23572;
															assign node23572 = (inp[8]) ? 4'b1101 : node23573;
																assign node23573 = (inp[7]) ? 4'b1101 : 4'b1100;
															assign node23577 = (inp[7]) ? 4'b1100 : node23578;
																assign node23578 = (inp[8]) ? 4'b1101 : 4'b1100;
													assign node23582 = (inp[9]) ? node23596 : node23583;
														assign node23583 = (inp[14]) ? node23591 : node23584;
															assign node23584 = (inp[7]) ? node23588 : node23585;
																assign node23585 = (inp[8]) ? 4'b1101 : 4'b1100;
																assign node23588 = (inp[8]) ? 4'b1100 : 4'b1101;
															assign node23591 = (inp[7]) ? node23593 : 4'b1101;
																assign node23593 = (inp[8]) ? 4'b1100 : 4'b1101;
														assign node23596 = (inp[7]) ? node23600 : node23597;
															assign node23597 = (inp[8]) ? 4'b1001 : 4'b1000;
															assign node23600 = (inp[8]) ? 4'b1000 : 4'b1001;
										assign node23603 = (inp[3]) ? node23649 : node23604;
											assign node23604 = (inp[7]) ? node23624 : node23605;
												assign node23605 = (inp[8]) ? node23609 : node23606;
													assign node23606 = (inp[12]) ? 4'b1000 : 4'b1100;
													assign node23609 = (inp[4]) ? node23617 : node23610;
														assign node23610 = (inp[9]) ? node23614 : node23611;
															assign node23611 = (inp[12]) ? 4'b1001 : 4'b1101;
															assign node23614 = (inp[12]) ? 4'b1101 : 4'b1001;
														assign node23617 = (inp[12]) ? node23621 : node23618;
															assign node23618 = (inp[9]) ? 4'b1101 : 4'b1001;
															assign node23621 = (inp[9]) ? 4'b1001 : 4'b1101;
												assign node23624 = (inp[8]) ? node23636 : node23625;
													assign node23625 = (inp[12]) ? node23631 : node23626;
														assign node23626 = (inp[9]) ? node23628 : 4'b1001;
															assign node23628 = (inp[4]) ? 4'b1101 : 4'b1001;
														assign node23631 = (inp[4]) ? 4'b1101 : node23632;
															assign node23632 = (inp[9]) ? 4'b1101 : 4'b1001;
													assign node23636 = (inp[14]) ? node23642 : node23637;
														assign node23637 = (inp[12]) ? node23639 : 4'b1000;
															assign node23639 = (inp[9]) ? 4'b1000 : 4'b1100;
														assign node23642 = (inp[9]) ? 4'b1100 : node23643;
															assign node23643 = (inp[4]) ? 4'b1000 : node23644;
																assign node23644 = (inp[12]) ? 4'b1000 : 4'b1100;
											assign node23649 = (inp[9]) ? node23675 : node23650;
												assign node23650 = (inp[12]) ? node23664 : node23651;
													assign node23651 = (inp[4]) ? node23659 : node23652;
														assign node23652 = (inp[8]) ? node23656 : node23653;
															assign node23653 = (inp[7]) ? 4'b1101 : 4'b1100;
															assign node23656 = (inp[7]) ? 4'b1100 : 4'b1101;
														assign node23659 = (inp[8]) ? node23661 : 4'b1001;
															assign node23661 = (inp[7]) ? 4'b1000 : 4'b1001;
													assign node23664 = (inp[4]) ? node23672 : node23665;
														assign node23665 = (inp[7]) ? node23669 : node23666;
															assign node23666 = (inp[8]) ? 4'b1001 : 4'b1000;
															assign node23669 = (inp[8]) ? 4'b1000 : 4'b1001;
														assign node23672 = (inp[14]) ? 4'b1110 : 4'b1111;
												assign node23675 = (inp[4]) ? node23691 : node23676;
													assign node23676 = (inp[12]) ? node23684 : node23677;
														assign node23677 = (inp[8]) ? node23681 : node23678;
															assign node23678 = (inp[7]) ? 4'b1001 : 4'b1000;
															assign node23681 = (inp[7]) ? 4'b1000 : 4'b1001;
														assign node23684 = (inp[14]) ? 4'b1111 : node23685;
															assign node23685 = (inp[8]) ? 4'b1110 : node23686;
																assign node23686 = (inp[7]) ? 4'b1111 : 4'b1110;
													assign node23691 = (inp[12]) ? node23701 : node23692;
														assign node23692 = (inp[14]) ? node23698 : node23693;
															assign node23693 = (inp[8]) ? node23695 : 4'b1111;
																assign node23695 = (inp[7]) ? 4'b1110 : 4'b1111;
															assign node23698 = (inp[7]) ? 4'b1111 : 4'b1110;
														assign node23701 = (inp[7]) ? node23703 : 4'b1011;
															assign node23703 = (inp[8]) ? 4'b1010 : 4'b1011;
									assign node23706 = (inp[15]) ? node23860 : node23707;
										assign node23707 = (inp[3]) ? node23797 : node23708;
											assign node23708 = (inp[14]) ? node23746 : node23709;
												assign node23709 = (inp[12]) ? node23731 : node23710;
													assign node23710 = (inp[9]) ? node23722 : node23711;
														assign node23711 = (inp[4]) ? node23717 : node23712;
															assign node23712 = (inp[8]) ? 4'b1101 : node23713;
																assign node23713 = (inp[7]) ? 4'b1101 : 4'b1100;
															assign node23717 = (inp[8]) ? 4'b1001 : node23718;
																assign node23718 = (inp[7]) ? 4'b1001 : 4'b1000;
														assign node23722 = (inp[4]) ? node23728 : node23723;
															assign node23723 = (inp[8]) ? node23725 : 4'b1001;
																assign node23725 = (inp[7]) ? 4'b1000 : 4'b1001;
															assign node23728 = (inp[7]) ? 4'b1100 : 4'b1101;
													assign node23731 = (inp[7]) ? node23739 : node23732;
														assign node23732 = (inp[8]) ? 4'b1001 : node23733;
															assign node23733 = (inp[4]) ? node23735 : 4'b1000;
																assign node23735 = (inp[9]) ? 4'b1000 : 4'b1100;
														assign node23739 = (inp[8]) ? 4'b1000 : node23740;
															assign node23740 = (inp[9]) ? node23742 : 4'b1001;
																assign node23742 = (inp[4]) ? 4'b1001 : 4'b1101;
												assign node23746 = (inp[12]) ? node23774 : node23747;
													assign node23747 = (inp[9]) ? node23761 : node23748;
														assign node23748 = (inp[4]) ? node23754 : node23749;
															assign node23749 = (inp[7]) ? node23751 : 4'b1100;
																assign node23751 = (inp[8]) ? 4'b1100 : 4'b1101;
															assign node23754 = (inp[8]) ? node23758 : node23755;
																assign node23755 = (inp[7]) ? 4'b1001 : 4'b1000;
																assign node23758 = (inp[7]) ? 4'b1000 : 4'b1001;
														assign node23761 = (inp[4]) ? node23767 : node23762;
															assign node23762 = (inp[8]) ? node23764 : 4'b1001;
																assign node23764 = (inp[7]) ? 4'b1000 : 4'b1001;
															assign node23767 = (inp[7]) ? node23771 : node23768;
																assign node23768 = (inp[8]) ? 4'b1101 : 4'b1100;
																assign node23771 = (inp[8]) ? 4'b1100 : 4'b1101;
													assign node23774 = (inp[7]) ? node23790 : node23775;
														assign node23775 = (inp[8]) ? node23783 : node23776;
															assign node23776 = (inp[9]) ? node23780 : node23777;
																assign node23777 = (inp[4]) ? 4'b1100 : 4'b1000;
																assign node23780 = (inp[4]) ? 4'b1000 : 4'b1100;
															assign node23783 = (inp[9]) ? node23787 : node23784;
																assign node23784 = (inp[4]) ? 4'b1101 : 4'b1001;
																assign node23787 = (inp[4]) ? 4'b1001 : 4'b1101;
														assign node23790 = (inp[8]) ? 4'b1100 : node23791;
															assign node23791 = (inp[9]) ? 4'b1101 : node23792;
																assign node23792 = (inp[4]) ? 4'b1101 : 4'b1001;
											assign node23797 = (inp[4]) ? node23829 : node23798;
												assign node23798 = (inp[12]) ? node23812 : node23799;
													assign node23799 = (inp[9]) ? node23805 : node23800;
														assign node23800 = (inp[8]) ? node23802 : 4'b1100;
															assign node23802 = (inp[7]) ? 4'b1100 : 4'b1101;
														assign node23805 = (inp[7]) ? node23809 : node23806;
															assign node23806 = (inp[8]) ? 4'b1001 : 4'b1000;
															assign node23809 = (inp[8]) ? 4'b1000 : 4'b1001;
													assign node23812 = (inp[9]) ? node23824 : node23813;
														assign node23813 = (inp[14]) ? node23819 : node23814;
															assign node23814 = (inp[7]) ? 4'b1001 : node23815;
																assign node23815 = (inp[8]) ? 4'b1001 : 4'b1000;
															assign node23819 = (inp[8]) ? node23821 : 4'b1000;
																assign node23821 = (inp[7]) ? 4'b1000 : 4'b1001;
														assign node23824 = (inp[8]) ? node23826 : 4'b1111;
															assign node23826 = (inp[7]) ? 4'b1110 : 4'b1111;
												assign node23829 = (inp[12]) ? node23843 : node23830;
													assign node23830 = (inp[9]) ? node23838 : node23831;
														assign node23831 = (inp[14]) ? 4'b1001 : node23832;
															assign node23832 = (inp[8]) ? node23834 : 4'b1000;
																assign node23834 = (inp[7]) ? 4'b1000 : 4'b1001;
														assign node23838 = (inp[7]) ? node23840 : 4'b1111;
															assign node23840 = (inp[8]) ? 4'b1110 : 4'b1111;
													assign node23843 = (inp[9]) ? node23853 : node23844;
														assign node23844 = (inp[14]) ? 4'b1110 : node23845;
															assign node23845 = (inp[8]) ? node23849 : node23846;
																assign node23846 = (inp[7]) ? 4'b1111 : 4'b1110;
																assign node23849 = (inp[7]) ? 4'b1110 : 4'b1111;
														assign node23853 = (inp[8]) ? node23857 : node23854;
															assign node23854 = (inp[7]) ? 4'b1011 : 4'b1010;
															assign node23857 = (inp[7]) ? 4'b1010 : 4'b1011;
										assign node23860 = (inp[3]) ? node23928 : node23861;
											assign node23861 = (inp[9]) ? node23897 : node23862;
												assign node23862 = (inp[12]) ? node23880 : node23863;
													assign node23863 = (inp[4]) ? node23875 : node23864;
														assign node23864 = (inp[14]) ? node23870 : node23865;
															assign node23865 = (inp[8]) ? node23867 : 4'b1110;
																assign node23867 = (inp[7]) ? 4'b1110 : 4'b1111;
															assign node23870 = (inp[8]) ? 4'b1110 : node23871;
																assign node23871 = (inp[7]) ? 4'b1111 : 4'b1110;
														assign node23875 = (inp[7]) ? 4'b1010 : node23876;
															assign node23876 = (inp[8]) ? 4'b1011 : 4'b1010;
													assign node23880 = (inp[4]) ? node23892 : node23881;
														assign node23881 = (inp[14]) ? node23887 : node23882;
															assign node23882 = (inp[8]) ? 4'b1010 : node23883;
																assign node23883 = (inp[7]) ? 4'b1011 : 4'b1010;
															assign node23887 = (inp[7]) ? 4'b1011 : node23888;
																assign node23888 = (inp[8]) ? 4'b1011 : 4'b1010;
														assign node23892 = (inp[7]) ? node23894 : 4'b1110;
															assign node23894 = (inp[8]) ? 4'b1110 : 4'b1111;
												assign node23897 = (inp[12]) ? node23913 : node23898;
													assign node23898 = (inp[4]) ? node23906 : node23899;
														assign node23899 = (inp[8]) ? node23903 : node23900;
															assign node23900 = (inp[7]) ? 4'b1011 : 4'b1010;
															assign node23903 = (inp[7]) ? 4'b1010 : 4'b1011;
														assign node23906 = (inp[14]) ? 4'b1110 : node23907;
															assign node23907 = (inp[8]) ? node23909 : 4'b1111;
																assign node23909 = (inp[7]) ? 4'b1110 : 4'b1111;
													assign node23913 = (inp[4]) ? node23921 : node23914;
														assign node23914 = (inp[7]) ? node23918 : node23915;
															assign node23915 = (inp[8]) ? 4'b1111 : 4'b1110;
															assign node23918 = (inp[8]) ? 4'b1110 : 4'b1111;
														assign node23921 = (inp[14]) ? node23923 : 4'b1010;
															assign node23923 = (inp[8]) ? node23925 : 4'b1011;
																assign node23925 = (inp[7]) ? 4'b1010 : 4'b1011;
											assign node23928 = (inp[9]) ? node23962 : node23929;
												assign node23929 = (inp[12]) ? node23947 : node23930;
													assign node23930 = (inp[4]) ? node23940 : node23931;
														assign node23931 = (inp[14]) ? 4'b1110 : node23932;
															assign node23932 = (inp[8]) ? node23936 : node23933;
																assign node23933 = (inp[7]) ? 4'b1111 : 4'b1110;
																assign node23936 = (inp[7]) ? 4'b1110 : 4'b1111;
														assign node23940 = (inp[7]) ? node23944 : node23941;
															assign node23941 = (inp[8]) ? 4'b1011 : 4'b1010;
															assign node23944 = (inp[8]) ? 4'b1010 : 4'b1011;
													assign node23947 = (inp[4]) ? node23955 : node23948;
														assign node23948 = (inp[8]) ? node23952 : node23949;
															assign node23949 = (inp[7]) ? 4'b1011 : 4'b1010;
															assign node23952 = (inp[7]) ? 4'b1010 : 4'b1011;
														assign node23955 = (inp[7]) ? node23959 : node23956;
															assign node23956 = (inp[8]) ? 4'b1101 : 4'b1100;
															assign node23959 = (inp[8]) ? 4'b1100 : 4'b1101;
												assign node23962 = (inp[12]) ? node23974 : node23963;
													assign node23963 = (inp[4]) ? node23969 : node23964;
														assign node23964 = (inp[7]) ? node23966 : 4'b1011;
															assign node23966 = (inp[8]) ? 4'b1010 : 4'b1011;
														assign node23969 = (inp[8]) ? node23971 : 4'b1101;
															assign node23971 = (inp[7]) ? 4'b1100 : 4'b1101;
													assign node23974 = (inp[4]) ? node23978 : node23975;
														assign node23975 = (inp[14]) ? 4'b1101 : 4'b1100;
														assign node23978 = (inp[14]) ? 4'b1000 : node23979;
															assign node23979 = (inp[7]) ? node23981 : 4'b1001;
																assign node23981 = (inp[8]) ? 4'b1000 : 4'b1001;
							assign node23985 = (inp[15]) ? node24513 : node23986;
								assign node23986 = (inp[0]) ? node24258 : node23987;
									assign node23987 = (inp[3]) ? node24113 : node23988;
										assign node23988 = (inp[9]) ? node24050 : node23989;
											assign node23989 = (inp[12]) ? node24027 : node23990;
												assign node23990 = (inp[4]) ? node24008 : node23991;
													assign node23991 = (inp[2]) ? node24001 : node23992;
														assign node23992 = (inp[8]) ? 4'b1111 : node23993;
															assign node23993 = (inp[7]) ? node23997 : node23994;
																assign node23994 = (inp[14]) ? 4'b1110 : 4'b1111;
																assign node23997 = (inp[14]) ? 4'b1111 : 4'b1110;
														assign node24001 = (inp[8]) ? node24005 : node24002;
															assign node24002 = (inp[7]) ? 4'b1111 : 4'b1110;
															assign node24005 = (inp[7]) ? 4'b1110 : 4'b1111;
													assign node24008 = (inp[14]) ? node24018 : node24009;
														assign node24009 = (inp[8]) ? node24011 : 4'b1010;
															assign node24011 = (inp[7]) ? node24015 : node24012;
																assign node24012 = (inp[2]) ? 4'b1011 : 4'b1010;
																assign node24015 = (inp[2]) ? 4'b1010 : 4'b1011;
														assign node24018 = (inp[2]) ? node24024 : node24019;
															assign node24019 = (inp[7]) ? 4'b1011 : node24020;
																assign node24020 = (inp[8]) ? 4'b1011 : 4'b1010;
															assign node24024 = (inp[8]) ? 4'b1010 : 4'b1011;
												assign node24027 = (inp[4]) ? node24039 : node24028;
													assign node24028 = (inp[2]) ? node24034 : node24029;
														assign node24029 = (inp[7]) ? node24031 : 4'b1011;
															assign node24031 = (inp[8]) ? 4'b1011 : 4'b1010;
														assign node24034 = (inp[7]) ? node24036 : 4'b1010;
															assign node24036 = (inp[8]) ? 4'b1010 : 4'b1011;
													assign node24039 = (inp[8]) ? node24041 : 4'b1101;
														assign node24041 = (inp[2]) ? node24047 : node24042;
															assign node24042 = (inp[14]) ? 4'b1100 : node24043;
																assign node24043 = (inp[7]) ? 4'b1101 : 4'b1100;
															assign node24047 = (inp[7]) ? 4'b1100 : 4'b1101;
											assign node24050 = (inp[4]) ? node24086 : node24051;
												assign node24051 = (inp[12]) ? node24067 : node24052;
													assign node24052 = (inp[8]) ? node24058 : node24053;
														assign node24053 = (inp[7]) ? 4'b1011 : node24054;
															assign node24054 = (inp[14]) ? 4'b1010 : 4'b1011;
														assign node24058 = (inp[14]) ? 4'b1010 : node24059;
															assign node24059 = (inp[2]) ? node24063 : node24060;
																assign node24060 = (inp[7]) ? 4'b1011 : 4'b1010;
																assign node24063 = (inp[7]) ? 4'b1010 : 4'b1011;
													assign node24067 = (inp[14]) ? node24077 : node24068;
														assign node24068 = (inp[2]) ? 4'b1101 : node24069;
															assign node24069 = (inp[7]) ? node24073 : node24070;
																assign node24070 = (inp[8]) ? 4'b1100 : 4'b1101;
																assign node24073 = (inp[8]) ? 4'b1101 : 4'b1100;
														assign node24077 = (inp[2]) ? node24079 : 4'b1100;
															assign node24079 = (inp[8]) ? node24083 : node24080;
																assign node24080 = (inp[7]) ? 4'b1101 : 4'b1100;
																assign node24083 = (inp[7]) ? 4'b1100 : 4'b1101;
												assign node24086 = (inp[12]) ? node24100 : node24087;
													assign node24087 = (inp[7]) ? node24095 : node24088;
														assign node24088 = (inp[8]) ? node24090 : 4'b1100;
															assign node24090 = (inp[2]) ? 4'b1101 : node24091;
																assign node24091 = (inp[14]) ? 4'b1101 : 4'b1100;
														assign node24095 = (inp[8]) ? node24097 : 4'b1101;
															assign node24097 = (inp[14]) ? 4'b1100 : 4'b1101;
													assign node24100 = (inp[2]) ? node24106 : node24101;
														assign node24101 = (inp[7]) ? node24103 : 4'b1001;
															assign node24103 = (inp[14]) ? 4'b1001 : 4'b1000;
														assign node24106 = (inp[7]) ? node24110 : node24107;
															assign node24107 = (inp[8]) ? 4'b1001 : 4'b1000;
															assign node24110 = (inp[8]) ? 4'b1000 : 4'b1001;
										assign node24113 = (inp[9]) ? node24185 : node24114;
											assign node24114 = (inp[7]) ? node24150 : node24115;
												assign node24115 = (inp[8]) ? node24135 : node24116;
													assign node24116 = (inp[2]) ? node24124 : node24117;
														assign node24117 = (inp[14]) ? node24119 : 4'b1101;
															assign node24119 = (inp[4]) ? node24121 : 4'b1100;
																assign node24121 = (inp[12]) ? 4'b1100 : 4'b1000;
														assign node24124 = (inp[14]) ? node24130 : node24125;
															assign node24125 = (inp[12]) ? node24127 : 4'b1100;
																assign node24127 = (inp[4]) ? 4'b1100 : 4'b1000;
															assign node24130 = (inp[12]) ? 4'b1100 : node24131;
																assign node24131 = (inp[4]) ? 4'b1000 : 4'b1100;
													assign node24135 = (inp[2]) ? node24143 : node24136;
														assign node24136 = (inp[14]) ? 4'b1101 : node24137;
															assign node24137 = (inp[12]) ? 4'b1000 : node24138;
																assign node24138 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node24143 = (inp[4]) ? node24147 : node24144;
															assign node24144 = (inp[12]) ? 4'b1001 : 4'b1101;
															assign node24147 = (inp[12]) ? 4'b1101 : 4'b1001;
												assign node24150 = (inp[8]) ? node24170 : node24151;
													assign node24151 = (inp[14]) ? node24163 : node24152;
														assign node24152 = (inp[2]) ? node24160 : node24153;
															assign node24153 = (inp[12]) ? node24157 : node24154;
																assign node24154 = (inp[4]) ? 4'b1000 : 4'b1100;
																assign node24157 = (inp[4]) ? 4'b1100 : 4'b1000;
															assign node24160 = (inp[12]) ? 4'b1101 : 4'b1001;
														assign node24163 = (inp[4]) ? node24167 : node24164;
															assign node24164 = (inp[12]) ? 4'b1001 : 4'b1101;
															assign node24167 = (inp[12]) ? 4'b1101 : 4'b1001;
													assign node24170 = (inp[2]) ? node24178 : node24171;
														assign node24171 = (inp[14]) ? 4'b1100 : node24172;
															assign node24172 = (inp[4]) ? 4'b1101 : node24173;
																assign node24173 = (inp[12]) ? 4'b1001 : 4'b1101;
														assign node24178 = (inp[4]) ? node24182 : node24179;
															assign node24179 = (inp[12]) ? 4'b1000 : 4'b1100;
															assign node24182 = (inp[12]) ? 4'b1100 : 4'b1000;
											assign node24185 = (inp[14]) ? node24229 : node24186;
												assign node24186 = (inp[7]) ? node24206 : node24187;
													assign node24187 = (inp[8]) ? node24199 : node24188;
														assign node24188 = (inp[2]) ? node24194 : node24189;
															assign node24189 = (inp[4]) ? 4'b1001 : node24190;
																assign node24190 = (inp[12]) ? 4'b1101 : 4'b1001;
															assign node24194 = (inp[12]) ? node24196 : 4'b1000;
																assign node24196 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node24199 = (inp[2]) ? node24201 : 4'b1100;
															assign node24201 = (inp[4]) ? 4'b1001 : node24202;
																assign node24202 = (inp[12]) ? 4'b1101 : 4'b1001;
													assign node24206 = (inp[8]) ? node24218 : node24207;
														assign node24207 = (inp[2]) ? node24215 : node24208;
															assign node24208 = (inp[4]) ? node24212 : node24209;
																assign node24209 = (inp[12]) ? 4'b1100 : 4'b1000;
																assign node24212 = (inp[12]) ? 4'b1000 : 4'b1100;
															assign node24215 = (inp[12]) ? 4'b1001 : 4'b1101;
														assign node24218 = (inp[2]) ? node24224 : node24219;
															assign node24219 = (inp[12]) ? node24221 : 4'b1001;
																assign node24221 = (inp[4]) ? 4'b1001 : 4'b1101;
															assign node24224 = (inp[12]) ? 4'b1000 : node24225;
																assign node24225 = (inp[4]) ? 4'b1100 : 4'b1000;
												assign node24229 = (inp[4]) ? node24241 : node24230;
													assign node24230 = (inp[12]) ? node24236 : node24231;
														assign node24231 = (inp[7]) ? node24233 : 4'b1000;
															assign node24233 = (inp[8]) ? 4'b1000 : 4'b1001;
														assign node24236 = (inp[8]) ? node24238 : 4'b1100;
															assign node24238 = (inp[7]) ? 4'b1100 : 4'b1101;
													assign node24241 = (inp[12]) ? node24251 : node24242;
														assign node24242 = (inp[2]) ? 4'b1101 : node24243;
															assign node24243 = (inp[7]) ? node24247 : node24244;
																assign node24244 = (inp[8]) ? 4'b1101 : 4'b1100;
																assign node24247 = (inp[8]) ? 4'b1100 : 4'b1101;
														assign node24251 = (inp[2]) ? node24253 : 4'b1000;
															assign node24253 = (inp[7]) ? 4'b1001 : node24254;
																assign node24254 = (inp[8]) ? 4'b1001 : 4'b1000;
									assign node24258 = (inp[3]) ? node24376 : node24259;
										assign node24259 = (inp[9]) ? node24321 : node24260;
											assign node24260 = (inp[12]) ? node24286 : node24261;
												assign node24261 = (inp[4]) ? node24269 : node24262;
													assign node24262 = (inp[2]) ? node24264 : 4'b1100;
														assign node24264 = (inp[7]) ? node24266 : 4'b1101;
															assign node24266 = (inp[8]) ? 4'b1100 : 4'b1101;
													assign node24269 = (inp[2]) ? 4'b1001 : node24270;
														assign node24270 = (inp[14]) ? node24278 : node24271;
															assign node24271 = (inp[7]) ? node24275 : node24272;
																assign node24272 = (inp[8]) ? 4'b1000 : 4'b1001;
																assign node24275 = (inp[8]) ? 4'b1001 : 4'b1000;
															assign node24278 = (inp[8]) ? node24282 : node24279;
																assign node24279 = (inp[7]) ? 4'b1001 : 4'b1000;
																assign node24282 = (inp[7]) ? 4'b1000 : 4'b1001;
												assign node24286 = (inp[4]) ? node24302 : node24287;
													assign node24287 = (inp[2]) ? node24295 : node24288;
														assign node24288 = (inp[7]) ? node24290 : 4'b1000;
															assign node24290 = (inp[14]) ? node24292 : 4'b1001;
																assign node24292 = (inp[8]) ? 4'b1000 : 4'b1001;
														assign node24295 = (inp[7]) ? node24299 : node24296;
															assign node24296 = (inp[8]) ? 4'b1001 : 4'b1000;
															assign node24299 = (inp[8]) ? 4'b1000 : 4'b1001;
													assign node24302 = (inp[8]) ? node24310 : node24303;
														assign node24303 = (inp[7]) ? 4'b1111 : node24304;
															assign node24304 = (inp[14]) ? 4'b1110 : node24305;
																assign node24305 = (inp[2]) ? 4'b1110 : 4'b1111;
														assign node24310 = (inp[7]) ? node24316 : node24311;
															assign node24311 = (inp[14]) ? 4'b1111 : node24312;
																assign node24312 = (inp[2]) ? 4'b1111 : 4'b1110;
															assign node24316 = (inp[14]) ? 4'b1110 : node24317;
																assign node24317 = (inp[2]) ? 4'b1110 : 4'b1111;
											assign node24321 = (inp[4]) ? node24349 : node24322;
												assign node24322 = (inp[12]) ? node24336 : node24323;
													assign node24323 = (inp[14]) ? node24329 : node24324;
														assign node24324 = (inp[7]) ? node24326 : 4'b1000;
															assign node24326 = (inp[8]) ? 4'b1001 : 4'b1000;
														assign node24329 = (inp[7]) ? node24333 : node24330;
															assign node24330 = (inp[8]) ? 4'b1001 : 4'b1000;
															assign node24333 = (inp[8]) ? 4'b1000 : 4'b1001;
													assign node24336 = (inp[8]) ? node24344 : node24337;
														assign node24337 = (inp[7]) ? 4'b1111 : node24338;
															assign node24338 = (inp[2]) ? 4'b1110 : node24339;
																assign node24339 = (inp[14]) ? 4'b1110 : 4'b1111;
														assign node24344 = (inp[7]) ? 4'b1110 : node24345;
															assign node24345 = (inp[2]) ? 4'b1111 : 4'b1110;
												assign node24349 = (inp[12]) ? node24363 : node24350;
													assign node24350 = (inp[7]) ? node24356 : node24351;
														assign node24351 = (inp[8]) ? node24353 : 4'b1110;
															assign node24353 = (inp[14]) ? 4'b1111 : 4'b1110;
														assign node24356 = (inp[8]) ? 4'b1110 : node24357;
															assign node24357 = (inp[14]) ? 4'b1111 : node24358;
																assign node24358 = (inp[2]) ? 4'b1111 : 4'b1110;
													assign node24363 = (inp[8]) ? node24371 : node24364;
														assign node24364 = (inp[14]) ? 4'b1011 : node24365;
															assign node24365 = (inp[2]) ? node24367 : 4'b1010;
																assign node24367 = (inp[7]) ? 4'b1011 : 4'b1010;
														assign node24371 = (inp[14]) ? 4'b1010 : node24372;
															assign node24372 = (inp[2]) ? 4'b1011 : 4'b1010;
										assign node24376 = (inp[2]) ? node24450 : node24377;
											assign node24377 = (inp[14]) ? node24415 : node24378;
												assign node24378 = (inp[9]) ? node24398 : node24379;
													assign node24379 = (inp[4]) ? node24389 : node24380;
														assign node24380 = (inp[12]) ? node24386 : node24381;
															assign node24381 = (inp[7]) ? node24383 : 4'b1111;
																assign node24383 = (inp[8]) ? 4'b1111 : 4'b1110;
															assign node24386 = (inp[7]) ? 4'b1010 : 4'b1011;
														assign node24389 = (inp[12]) ? 4'b1110 : node24390;
															assign node24390 = (inp[7]) ? node24394 : node24391;
																assign node24391 = (inp[8]) ? 4'b1010 : 4'b1011;
																assign node24394 = (inp[8]) ? 4'b1011 : 4'b1010;
													assign node24398 = (inp[12]) ? node24408 : node24399;
														assign node24399 = (inp[4]) ? node24403 : node24400;
															assign node24400 = (inp[8]) ? 4'b1010 : 4'b1011;
															assign node24403 = (inp[7]) ? node24405 : 4'b1110;
																assign node24405 = (inp[8]) ? 4'b1111 : 4'b1110;
														assign node24408 = (inp[4]) ? 4'b1011 : node24409;
															assign node24409 = (inp[8]) ? node24411 : 4'b1111;
																assign node24411 = (inp[7]) ? 4'b1111 : 4'b1110;
												assign node24415 = (inp[4]) ? node24437 : node24416;
													assign node24416 = (inp[7]) ? node24424 : node24417;
														assign node24417 = (inp[8]) ? 4'b1111 : node24418;
															assign node24418 = (inp[9]) ? 4'b1010 : node24419;
																assign node24419 = (inp[12]) ? 4'b1010 : 4'b1110;
														assign node24424 = (inp[8]) ? node24432 : node24425;
															assign node24425 = (inp[12]) ? node24429 : node24426;
																assign node24426 = (inp[9]) ? 4'b1011 : 4'b1111;
																assign node24429 = (inp[9]) ? 4'b1111 : 4'b1011;
															assign node24432 = (inp[9]) ? node24434 : 4'b1010;
																assign node24434 = (inp[12]) ? 4'b1110 : 4'b1010;
													assign node24437 = (inp[9]) ? node24443 : node24438;
														assign node24438 = (inp[12]) ? 4'b1111 : node24439;
															assign node24439 = (inp[7]) ? 4'b1010 : 4'b1011;
														assign node24443 = (inp[12]) ? node24445 : 4'b1111;
															assign node24445 = (inp[7]) ? 4'b1011 : node24446;
																assign node24446 = (inp[8]) ? 4'b1011 : 4'b1010;
											assign node24450 = (inp[12]) ? node24488 : node24451;
												assign node24451 = (inp[14]) ? node24473 : node24452;
													assign node24452 = (inp[7]) ? node24466 : node24453;
														assign node24453 = (inp[8]) ? node24459 : node24454;
															assign node24454 = (inp[4]) ? node24456 : 4'b1110;
																assign node24456 = (inp[9]) ? 4'b1110 : 4'b1010;
															assign node24459 = (inp[4]) ? node24463 : node24460;
																assign node24460 = (inp[9]) ? 4'b1011 : 4'b1111;
																assign node24463 = (inp[9]) ? 4'b1111 : 4'b1011;
														assign node24466 = (inp[8]) ? node24468 : 4'b1011;
															assign node24468 = (inp[4]) ? 4'b1110 : node24469;
																assign node24469 = (inp[9]) ? 4'b1010 : 4'b1110;
													assign node24473 = (inp[4]) ? node24481 : node24474;
														assign node24474 = (inp[9]) ? 4'b1010 : node24475;
															assign node24475 = (inp[7]) ? node24477 : 4'b1110;
																assign node24477 = (inp[8]) ? 4'b1110 : 4'b1111;
														assign node24481 = (inp[7]) ? node24485 : node24482;
															assign node24482 = (inp[8]) ? 4'b1011 : 4'b1010;
															assign node24485 = (inp[8]) ? 4'b1010 : 4'b1011;
												assign node24488 = (inp[9]) ? node24504 : node24489;
													assign node24489 = (inp[4]) ? node24497 : node24490;
														assign node24490 = (inp[8]) ? node24494 : node24491;
															assign node24491 = (inp[7]) ? 4'b1011 : 4'b1010;
															assign node24494 = (inp[7]) ? 4'b1010 : 4'b1011;
														assign node24497 = (inp[8]) ? node24501 : node24498;
															assign node24498 = (inp[7]) ? 4'b1111 : 4'b1110;
															assign node24501 = (inp[7]) ? 4'b1110 : 4'b1111;
													assign node24504 = (inp[4]) ? 4'b1010 : node24505;
														assign node24505 = (inp[7]) ? node24509 : node24506;
															assign node24506 = (inp[8]) ? 4'b1111 : 4'b1110;
															assign node24509 = (inp[8]) ? 4'b1110 : 4'b1111;
								assign node24513 = (inp[0]) ? node24789 : node24514;
									assign node24514 = (inp[3]) ? node24658 : node24515;
										assign node24515 = (inp[4]) ? node24589 : node24516;
											assign node24516 = (inp[12]) ? node24554 : node24517;
												assign node24517 = (inp[9]) ? node24531 : node24518;
													assign node24518 = (inp[14]) ? node24524 : node24519;
														assign node24519 = (inp[2]) ? 4'b1101 : node24520;
															assign node24520 = (inp[8]) ? 4'b1100 : 4'b1101;
														assign node24524 = (inp[7]) ? node24528 : node24525;
															assign node24525 = (inp[8]) ? 4'b1101 : 4'b1100;
															assign node24528 = (inp[8]) ? 4'b1100 : 4'b1101;
													assign node24531 = (inp[14]) ? node24547 : node24532;
														assign node24532 = (inp[7]) ? node24540 : node24533;
															assign node24533 = (inp[2]) ? node24537 : node24534;
																assign node24534 = (inp[8]) ? 4'b1000 : 4'b1001;
																assign node24537 = (inp[8]) ? 4'b1001 : 4'b1000;
															assign node24540 = (inp[2]) ? node24544 : node24541;
																assign node24541 = (inp[8]) ? 4'b1001 : 4'b1000;
																assign node24544 = (inp[8]) ? 4'b1000 : 4'b1001;
														assign node24547 = (inp[8]) ? node24551 : node24548;
															assign node24548 = (inp[7]) ? 4'b1001 : 4'b1000;
															assign node24551 = (inp[7]) ? 4'b1000 : 4'b1001;
												assign node24554 = (inp[9]) ? node24570 : node24555;
													assign node24555 = (inp[8]) ? node24561 : node24556;
														assign node24556 = (inp[7]) ? node24558 : 4'b1000;
															assign node24558 = (inp[14]) ? 4'b1001 : 4'b1000;
														assign node24561 = (inp[14]) ? 4'b1000 : node24562;
															assign node24562 = (inp[2]) ? node24566 : node24563;
																assign node24563 = (inp[7]) ? 4'b1001 : 4'b1000;
																assign node24566 = (inp[7]) ? 4'b1000 : 4'b1001;
													assign node24570 = (inp[7]) ? node24578 : node24571;
														assign node24571 = (inp[8]) ? 4'b1111 : node24572;
															assign node24572 = (inp[14]) ? 4'b1110 : node24573;
																assign node24573 = (inp[2]) ? 4'b1110 : 4'b1111;
														assign node24578 = (inp[8]) ? node24584 : node24579;
															assign node24579 = (inp[2]) ? 4'b1111 : node24580;
																assign node24580 = (inp[14]) ? 4'b1111 : 4'b1110;
															assign node24584 = (inp[14]) ? 4'b1110 : node24585;
																assign node24585 = (inp[2]) ? 4'b1110 : 4'b1111;
											assign node24589 = (inp[12]) ? node24617 : node24590;
												assign node24590 = (inp[9]) ? node24602 : node24591;
													assign node24591 = (inp[8]) ? node24597 : node24592;
														assign node24592 = (inp[7]) ? 4'b1001 : node24593;
															assign node24593 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node24597 = (inp[7]) ? 4'b1000 : node24598;
															assign node24598 = (inp[2]) ? 4'b1001 : 4'b1000;
													assign node24602 = (inp[14]) ? node24610 : node24603;
														assign node24603 = (inp[8]) ? 4'b1111 : node24604;
															assign node24604 = (inp[2]) ? 4'b1111 : node24605;
																assign node24605 = (inp[7]) ? 4'b1110 : 4'b1111;
														assign node24610 = (inp[8]) ? node24614 : node24611;
															assign node24611 = (inp[7]) ? 4'b1111 : 4'b1110;
															assign node24614 = (inp[7]) ? 4'b1110 : 4'b1111;
												assign node24617 = (inp[9]) ? node24637 : node24618;
													assign node24618 = (inp[8]) ? node24628 : node24619;
														assign node24619 = (inp[7]) ? node24625 : node24620;
															assign node24620 = (inp[2]) ? 4'b1110 : node24621;
																assign node24621 = (inp[14]) ? 4'b1110 : 4'b1111;
															assign node24625 = (inp[2]) ? 4'b1111 : 4'b1110;
														assign node24628 = (inp[14]) ? 4'b1111 : node24629;
															assign node24629 = (inp[2]) ? node24633 : node24630;
																assign node24630 = (inp[7]) ? 4'b1111 : 4'b1110;
																assign node24633 = (inp[7]) ? 4'b1110 : 4'b1111;
													assign node24637 = (inp[8]) ? node24649 : node24638;
														assign node24638 = (inp[7]) ? node24644 : node24639;
															assign node24639 = (inp[14]) ? 4'b1010 : node24640;
																assign node24640 = (inp[2]) ? 4'b1010 : 4'b1011;
															assign node24644 = (inp[14]) ? 4'b1011 : node24645;
																assign node24645 = (inp[2]) ? 4'b1011 : 4'b1010;
														assign node24649 = (inp[7]) ? node24653 : node24650;
															assign node24650 = (inp[14]) ? 4'b1011 : 4'b1010;
															assign node24653 = (inp[14]) ? 4'b1010 : node24654;
																assign node24654 = (inp[2]) ? 4'b1010 : 4'b1011;
										assign node24658 = (inp[7]) ? node24728 : node24659;
											assign node24659 = (inp[8]) ? node24693 : node24660;
												assign node24660 = (inp[2]) ? node24672 : node24661;
													assign node24661 = (inp[14]) ? node24667 : node24662;
														assign node24662 = (inp[9]) ? node24664 : 4'b1111;
															assign node24664 = (inp[4]) ? 4'b1111 : 4'b1011;
														assign node24667 = (inp[12]) ? 4'b1010 : node24668;
															assign node24668 = (inp[4]) ? 4'b1110 : 4'b1010;
													assign node24672 = (inp[4]) ? node24686 : node24673;
														assign node24673 = (inp[14]) ? node24679 : node24674;
															assign node24674 = (inp[12]) ? node24676 : 4'b1110;
																assign node24676 = (inp[9]) ? 4'b1110 : 4'b1010;
															assign node24679 = (inp[9]) ? node24683 : node24680;
																assign node24680 = (inp[12]) ? 4'b1010 : 4'b1110;
																assign node24683 = (inp[12]) ? 4'b1110 : 4'b1010;
														assign node24686 = (inp[12]) ? node24690 : node24687;
															assign node24687 = (inp[9]) ? 4'b1110 : 4'b1010;
															assign node24690 = (inp[9]) ? 4'b1010 : 4'b1110;
												assign node24693 = (inp[14]) ? node24711 : node24694;
													assign node24694 = (inp[2]) ? node24702 : node24695;
														assign node24695 = (inp[4]) ? node24697 : 4'b1010;
															assign node24697 = (inp[12]) ? 4'b1010 : node24698;
																assign node24698 = (inp[9]) ? 4'b1110 : 4'b1010;
														assign node24702 = (inp[9]) ? node24704 : 4'b1011;
															assign node24704 = (inp[4]) ? node24708 : node24705;
																assign node24705 = (inp[12]) ? 4'b1111 : 4'b1011;
																assign node24708 = (inp[12]) ? 4'b1011 : 4'b1111;
													assign node24711 = (inp[4]) ? node24719 : node24712;
														assign node24712 = (inp[9]) ? node24716 : node24713;
															assign node24713 = (inp[12]) ? 4'b1011 : 4'b1111;
															assign node24716 = (inp[12]) ? 4'b1111 : 4'b1011;
														assign node24719 = (inp[2]) ? 4'b1011 : node24720;
															assign node24720 = (inp[9]) ? node24724 : node24721;
																assign node24721 = (inp[12]) ? 4'b1111 : 4'b1011;
																assign node24724 = (inp[12]) ? 4'b1011 : 4'b1111;
											assign node24728 = (inp[8]) ? node24764 : node24729;
												assign node24729 = (inp[2]) ? node24743 : node24730;
													assign node24730 = (inp[14]) ? node24732 : 4'b1010;
														assign node24732 = (inp[4]) ? node24738 : node24733;
															assign node24733 = (inp[9]) ? 4'b1011 : node24734;
																assign node24734 = (inp[12]) ? 4'b1011 : 4'b1111;
															assign node24738 = (inp[9]) ? 4'b1111 : node24739;
																assign node24739 = (inp[12]) ? 4'b1111 : 4'b1011;
													assign node24743 = (inp[9]) ? node24751 : node24744;
														assign node24744 = (inp[4]) ? node24748 : node24745;
															assign node24745 = (inp[12]) ? 4'b1011 : 4'b1111;
															assign node24748 = (inp[12]) ? 4'b1111 : 4'b1011;
														assign node24751 = (inp[14]) ? node24759 : node24752;
															assign node24752 = (inp[12]) ? node24756 : node24753;
																assign node24753 = (inp[4]) ? 4'b1111 : 4'b1011;
																assign node24756 = (inp[4]) ? 4'b1011 : 4'b1111;
															assign node24759 = (inp[4]) ? node24761 : 4'b1011;
																assign node24761 = (inp[12]) ? 4'b1011 : 4'b1111;
												assign node24764 = (inp[14]) ? node24776 : node24765;
													assign node24765 = (inp[2]) ? node24771 : node24766;
														assign node24766 = (inp[12]) ? node24768 : 4'b1111;
															assign node24768 = (inp[4]) ? 4'b1011 : 4'b1111;
														assign node24771 = (inp[9]) ? node24773 : 4'b1110;
															assign node24773 = (inp[12]) ? 4'b1110 : 4'b1010;
													assign node24776 = (inp[4]) ? node24784 : node24777;
														assign node24777 = (inp[12]) ? node24781 : node24778;
															assign node24778 = (inp[9]) ? 4'b1010 : 4'b1110;
															assign node24781 = (inp[9]) ? 4'b1110 : 4'b1010;
														assign node24784 = (inp[12]) ? 4'b1110 : node24785;
															assign node24785 = (inp[2]) ? 4'b1010 : 4'b1110;
									assign node24789 = (inp[3]) ? node24881 : node24790;
										assign node24790 = (inp[12]) ? node24846 : node24791;
											assign node24791 = (inp[4]) ? node24825 : node24792;
												assign node24792 = (inp[9]) ? node24808 : node24793;
													assign node24793 = (inp[7]) ? node24803 : node24794;
														assign node24794 = (inp[8]) ? node24800 : node24795;
															assign node24795 = (inp[14]) ? 4'b1110 : node24796;
																assign node24796 = (inp[2]) ? 4'b1110 : 4'b1111;
															assign node24800 = (inp[2]) ? 4'b1111 : 4'b1110;
														assign node24803 = (inp[8]) ? node24805 : 4'b1111;
															assign node24805 = (inp[14]) ? 4'b1110 : 4'b1111;
													assign node24808 = (inp[8]) ? node24814 : node24809;
														assign node24809 = (inp[7]) ? 4'b1011 : node24810;
															assign node24810 = (inp[14]) ? 4'b1010 : 4'b1011;
														assign node24814 = (inp[7]) ? node24820 : node24815;
															assign node24815 = (inp[2]) ? 4'b1011 : node24816;
																assign node24816 = (inp[14]) ? 4'b1011 : 4'b1010;
															assign node24820 = (inp[2]) ? 4'b1010 : node24821;
																assign node24821 = (inp[14]) ? 4'b1010 : 4'b1011;
												assign node24825 = (inp[9]) ? node24839 : node24826;
													assign node24826 = (inp[7]) ? node24832 : node24827;
														assign node24827 = (inp[2]) ? 4'b1011 : node24828;
															assign node24828 = (inp[14]) ? 4'b1010 : 4'b1011;
														assign node24832 = (inp[8]) ? 4'b1010 : node24833;
															assign node24833 = (inp[14]) ? 4'b1011 : node24834;
																assign node24834 = (inp[2]) ? 4'b1011 : 4'b1010;
													assign node24839 = (inp[8]) ? node24843 : node24840;
														assign node24840 = (inp[14]) ? 4'b1101 : 4'b1100;
														assign node24843 = (inp[2]) ? 4'b1100 : 4'b1101;
											assign node24846 = (inp[4]) ? node24860 : node24847;
												assign node24847 = (inp[9]) ? node24857 : node24848;
													assign node24848 = (inp[7]) ? 4'b1010 : node24849;
														assign node24849 = (inp[8]) ? node24851 : 4'b1010;
															assign node24851 = (inp[14]) ? 4'b1011 : node24852;
																assign node24852 = (inp[2]) ? 4'b1011 : 4'b1010;
													assign node24857 = (inp[7]) ? 4'b1100 : 4'b1101;
												assign node24860 = (inp[9]) ? node24874 : node24861;
													assign node24861 = (inp[7]) ? node24867 : node24862;
														assign node24862 = (inp[8]) ? node24864 : 4'b1100;
															assign node24864 = (inp[14]) ? 4'b1101 : 4'b1100;
														assign node24867 = (inp[8]) ? 4'b1100 : node24868;
															assign node24868 = (inp[14]) ? 4'b1101 : node24869;
																assign node24869 = (inp[2]) ? 4'b1101 : 4'b1100;
													assign node24874 = (inp[8]) ? node24876 : 4'b1000;
														assign node24876 = (inp[7]) ? node24878 : 4'b1001;
															assign node24878 = (inp[14]) ? 4'b1000 : 4'b1001;
										assign node24881 = (inp[8]) ? node24941 : node24882;
											assign node24882 = (inp[7]) ? node24912 : node24883;
												assign node24883 = (inp[2]) ? node24899 : node24884;
													assign node24884 = (inp[14]) ? node24892 : node24885;
														assign node24885 = (inp[4]) ? 4'b1101 : node24886;
															assign node24886 = (inp[12]) ? 4'b1001 : node24887;
																assign node24887 = (inp[9]) ? 4'b1001 : 4'b1101;
														assign node24892 = (inp[12]) ? 4'b1000 : node24893;
															assign node24893 = (inp[4]) ? 4'b1100 : node24894;
																assign node24894 = (inp[9]) ? 4'b1000 : 4'b1100;
													assign node24899 = (inp[9]) ? node24905 : node24900;
														assign node24900 = (inp[4]) ? 4'b1000 : node24901;
															assign node24901 = (inp[12]) ? 4'b1000 : 4'b1100;
														assign node24905 = (inp[14]) ? 4'b1100 : node24906;
															assign node24906 = (inp[12]) ? 4'b1000 : node24907;
																assign node24907 = (inp[4]) ? 4'b1100 : 4'b1000;
												assign node24912 = (inp[14]) ? node24926 : node24913;
													assign node24913 = (inp[2]) ? node24923 : node24914;
														assign node24914 = (inp[4]) ? node24916 : 4'b1100;
															assign node24916 = (inp[9]) ? node24920 : node24917;
																assign node24917 = (inp[12]) ? 4'b1100 : 4'b1000;
																assign node24920 = (inp[12]) ? 4'b1000 : 4'b1100;
														assign node24923 = (inp[12]) ? 4'b1101 : 4'b1001;
													assign node24926 = (inp[12]) ? node24934 : node24927;
														assign node24927 = (inp[4]) ? node24931 : node24928;
															assign node24928 = (inp[9]) ? 4'b1001 : 4'b1101;
															assign node24931 = (inp[9]) ? 4'b1101 : 4'b1001;
														assign node24934 = (inp[4]) ? node24938 : node24935;
															assign node24935 = (inp[9]) ? 4'b1101 : 4'b1001;
															assign node24938 = (inp[9]) ? 4'b1001 : 4'b1101;
											assign node24941 = (inp[7]) ? node24965 : node24942;
												assign node24942 = (inp[14]) ? node24954 : node24943;
													assign node24943 = (inp[2]) ? node24951 : node24944;
														assign node24944 = (inp[12]) ? node24946 : 4'b1100;
															assign node24946 = (inp[4]) ? 4'b1100 : node24947;
																assign node24947 = (inp[9]) ? 4'b1100 : 4'b1000;
														assign node24951 = (inp[4]) ? 4'b1001 : 4'b1101;
													assign node24954 = (inp[9]) ? node24958 : node24955;
														assign node24955 = (inp[4]) ? 4'b1001 : 4'b1101;
														assign node24958 = (inp[2]) ? node24960 : 4'b1001;
															assign node24960 = (inp[4]) ? node24962 : 4'b1001;
																assign node24962 = (inp[12]) ? 4'b1001 : 4'b1101;
												assign node24965 = (inp[14]) ? node24977 : node24966;
													assign node24966 = (inp[2]) ? node24974 : node24967;
														assign node24967 = (inp[12]) ? node24969 : 4'b1001;
															assign node24969 = (inp[4]) ? node24971 : 4'b1001;
																assign node24971 = (inp[9]) ? 4'b1001 : 4'b1101;
														assign node24974 = (inp[4]) ? 4'b1100 : 4'b1000;
													assign node24977 = (inp[2]) ? node24991 : node24978;
														assign node24978 = (inp[9]) ? node24984 : node24979;
															assign node24979 = (inp[12]) ? 4'b1100 : node24980;
																assign node24980 = (inp[4]) ? 4'b1000 : 4'b1100;
															assign node24984 = (inp[12]) ? node24988 : node24985;
																assign node24985 = (inp[4]) ? 4'b1100 : 4'b1000;
																assign node24988 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node24991 = (inp[9]) ? node24993 : 4'b1000;
															assign node24993 = (inp[12]) ? node24995 : 4'b1000;
																assign node24995 = (inp[4]) ? 4'b1000 : 4'b1100;
						assign node24998 = (inp[8]) ? node25940 : node24999;
							assign node24999 = (inp[7]) ? node25493 : node25000;
								assign node25000 = (inp[14]) ? node25276 : node25001;
									assign node25001 = (inp[2]) ? node25135 : node25002;
										assign node25002 = (inp[0]) ? node25074 : node25003;
											assign node25003 = (inp[5]) ? node25043 : node25004;
												assign node25004 = (inp[15]) ? node25026 : node25005;
													assign node25005 = (inp[9]) ? node25015 : node25006;
														assign node25006 = (inp[3]) ? node25012 : node25007;
															assign node25007 = (inp[4]) ? node25009 : 4'b1011;
																assign node25009 = (inp[12]) ? 4'b1111 : 4'b1011;
															assign node25012 = (inp[12]) ? 4'b1011 : 4'b1111;
														assign node25015 = (inp[3]) ? node25019 : node25016;
															assign node25016 = (inp[12]) ? 4'b1011 : 4'b1111;
															assign node25019 = (inp[4]) ? node25023 : node25020;
																assign node25020 = (inp[12]) ? 4'b1101 : 4'b1011;
																assign node25023 = (inp[12]) ? 4'b1001 : 4'b1101;
													assign node25026 = (inp[4]) ? node25028 : 4'b1001;
														assign node25028 = (inp[3]) ? node25036 : node25029;
															assign node25029 = (inp[12]) ? node25033 : node25030;
																assign node25030 = (inp[9]) ? 4'b1101 : 4'b1001;
																assign node25033 = (inp[9]) ? 4'b1001 : 4'b1101;
															assign node25036 = (inp[9]) ? node25040 : node25037;
																assign node25037 = (inp[12]) ? 4'b1111 : 4'b1001;
																assign node25040 = (inp[12]) ? 4'b1011 : 4'b1111;
												assign node25043 = (inp[15]) ? node25059 : node25044;
													assign node25044 = (inp[3]) ? node25056 : node25045;
														assign node25045 = (inp[4]) ? node25051 : node25046;
															assign node25046 = (inp[12]) ? node25048 : 4'b1011;
																assign node25048 = (inp[9]) ? 4'b1101 : 4'b1011;
															assign node25051 = (inp[12]) ? 4'b1101 : node25052;
																assign node25052 = (inp[9]) ? 4'b1101 : 4'b1011;
														assign node25056 = (inp[4]) ? 4'b1001 : 4'b1101;
													assign node25059 = (inp[3]) ? node25067 : node25060;
														assign node25060 = (inp[9]) ? node25062 : 4'b1101;
															assign node25062 = (inp[4]) ? node25064 : 4'b1111;
																assign node25064 = (inp[12]) ? 4'b1011 : 4'b1111;
														assign node25067 = (inp[12]) ? 4'b1011 : node25068;
															assign node25068 = (inp[4]) ? node25070 : 4'b1011;
																assign node25070 = (inp[9]) ? 4'b1111 : 4'b1011;
											assign node25074 = (inp[4]) ? node25096 : node25075;
												assign node25075 = (inp[15]) ? node25087 : node25076;
													assign node25076 = (inp[9]) ? node25082 : node25077;
														assign node25077 = (inp[5]) ? node25079 : 4'b1101;
															assign node25079 = (inp[3]) ? 4'b1111 : 4'b1101;
														assign node25082 = (inp[12]) ? 4'b1111 : node25083;
															assign node25083 = (inp[3]) ? 4'b1011 : 4'b1001;
													assign node25087 = (inp[9]) ? node25091 : node25088;
														assign node25088 = (inp[12]) ? 4'b1011 : 4'b1111;
														assign node25091 = (inp[12]) ? node25093 : 4'b1011;
															assign node25093 = (inp[3]) ? 4'b1101 : 4'b1111;
												assign node25096 = (inp[15]) ? node25116 : node25097;
													assign node25097 = (inp[5]) ? node25107 : node25098;
														assign node25098 = (inp[3]) ? 4'b1111 : node25099;
															assign node25099 = (inp[12]) ? node25103 : node25100;
																assign node25100 = (inp[9]) ? 4'b1101 : 4'b1001;
																assign node25103 = (inp[9]) ? 4'b1001 : 4'b1101;
														assign node25107 = (inp[3]) ? node25109 : 4'b1111;
															assign node25109 = (inp[12]) ? node25113 : node25110;
																assign node25110 = (inp[9]) ? 4'b1111 : 4'b1011;
																assign node25113 = (inp[9]) ? 4'b1011 : 4'b1111;
													assign node25116 = (inp[5]) ? node25130 : node25117;
														assign node25117 = (inp[3]) ? node25123 : node25118;
															assign node25118 = (inp[12]) ? 4'b1111 : node25119;
																assign node25119 = (inp[9]) ? 4'b1111 : 4'b1011;
															assign node25123 = (inp[12]) ? node25127 : node25124;
																assign node25124 = (inp[9]) ? 4'b1101 : 4'b1011;
																assign node25127 = (inp[9]) ? 4'b1001 : 4'b1101;
														assign node25130 = (inp[3]) ? 4'b1101 : node25131;
															assign node25131 = (inp[9]) ? 4'b1001 : 4'b1101;
										assign node25135 = (inp[5]) ? node25209 : node25136;
											assign node25136 = (inp[15]) ? node25184 : node25137;
												assign node25137 = (inp[0]) ? node25155 : node25138;
													assign node25138 = (inp[3]) ? node25150 : node25139;
														assign node25139 = (inp[12]) ? node25145 : node25140;
															assign node25140 = (inp[9]) ? 4'b1110 : node25141;
																assign node25141 = (inp[4]) ? 4'b1010 : 4'b1110;
															assign node25145 = (inp[4]) ? node25147 : 4'b1010;
																assign node25147 = (inp[9]) ? 4'b1010 : 4'b1110;
														assign node25150 = (inp[12]) ? 4'b1100 : node25151;
															assign node25151 = (inp[9]) ? 4'b1010 : 4'b1110;
													assign node25155 = (inp[3]) ? node25169 : node25156;
														assign node25156 = (inp[9]) ? node25164 : node25157;
															assign node25157 = (inp[4]) ? node25161 : node25158;
																assign node25158 = (inp[12]) ? 4'b1000 : 4'b1100;
																assign node25161 = (inp[12]) ? 4'b1100 : 4'b1000;
															assign node25164 = (inp[12]) ? 4'b1000 : node25165;
																assign node25165 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node25169 = (inp[4]) ? node25177 : node25170;
															assign node25170 = (inp[9]) ? node25174 : node25171;
																assign node25171 = (inp[12]) ? 4'b1000 : 4'b1100;
																assign node25174 = (inp[12]) ? 4'b1110 : 4'b1000;
															assign node25177 = (inp[12]) ? node25181 : node25178;
																assign node25178 = (inp[9]) ? 4'b1110 : 4'b1000;
																assign node25181 = (inp[9]) ? 4'b1010 : 4'b1110;
												assign node25184 = (inp[0]) ? node25200 : node25185;
													assign node25185 = (inp[4]) ? node25191 : node25186;
														assign node25186 = (inp[12]) ? 4'b1000 : node25187;
															assign node25187 = (inp[9]) ? 4'b1000 : 4'b1100;
														assign node25191 = (inp[3]) ? node25195 : node25192;
															assign node25192 = (inp[12]) ? 4'b1000 : 4'b1100;
															assign node25195 = (inp[9]) ? node25197 : 4'b1110;
																assign node25197 = (inp[12]) ? 4'b1010 : 4'b1110;
													assign node25200 = (inp[9]) ? 4'b1010 : node25201;
														assign node25201 = (inp[12]) ? node25205 : node25202;
															assign node25202 = (inp[4]) ? 4'b1010 : 4'b1110;
															assign node25205 = (inp[4]) ? 4'b1110 : 4'b1010;
											assign node25209 = (inp[4]) ? node25253 : node25210;
												assign node25210 = (inp[12]) ? node25228 : node25211;
													assign node25211 = (inp[9]) ? 4'b1000 : node25212;
														assign node25212 = (inp[0]) ? node25220 : node25213;
															assign node25213 = (inp[15]) ? node25217 : node25214;
																assign node25214 = (inp[3]) ? 4'b1100 : 4'b1110;
																assign node25217 = (inp[3]) ? 4'b1110 : 4'b1100;
															assign node25220 = (inp[3]) ? node25224 : node25221;
																assign node25221 = (inp[15]) ? 4'b1110 : 4'b1100;
																assign node25224 = (inp[15]) ? 4'b1100 : 4'b1110;
													assign node25228 = (inp[9]) ? node25240 : node25229;
														assign node25229 = (inp[3]) ? node25235 : node25230;
															assign node25230 = (inp[0]) ? node25232 : 4'b1010;
																assign node25232 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node25235 = (inp[15]) ? 4'b1000 : node25236;
																assign node25236 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node25240 = (inp[3]) ? node25246 : node25241;
															assign node25241 = (inp[15]) ? node25243 : 4'b1110;
																assign node25243 = (inp[0]) ? 4'b1100 : 4'b1110;
															assign node25246 = (inp[0]) ? node25250 : node25247;
																assign node25247 = (inp[15]) ? 4'b1110 : 4'b1100;
																assign node25250 = (inp[15]) ? 4'b1100 : 4'b1110;
												assign node25253 = (inp[3]) ? node25265 : node25254;
													assign node25254 = (inp[9]) ? node25260 : node25255;
														assign node25255 = (inp[12]) ? 4'b1110 : node25256;
															assign node25256 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node25260 = (inp[12]) ? 4'b1000 : node25261;
															assign node25261 = (inp[0]) ? 4'b1110 : 4'b1100;
													assign node25265 = (inp[9]) ? node25273 : node25266;
														assign node25266 = (inp[12]) ? 4'b1100 : node25267;
															assign node25267 = (inp[0]) ? node25269 : 4'b1000;
																assign node25269 = (inp[15]) ? 4'b1000 : 4'b1010;
														assign node25273 = (inp[12]) ? 4'b1000 : 4'b1100;
									assign node25276 = (inp[0]) ? node25382 : node25277;
										assign node25277 = (inp[12]) ? node25319 : node25278;
											assign node25278 = (inp[15]) ? node25300 : node25279;
												assign node25279 = (inp[5]) ? node25289 : node25280;
													assign node25280 = (inp[9]) ? node25284 : node25281;
														assign node25281 = (inp[4]) ? 4'b1010 : 4'b1110;
														assign node25284 = (inp[3]) ? 4'b1100 : node25285;
															assign node25285 = (inp[2]) ? 4'b1110 : 4'b1010;
													assign node25289 = (inp[4]) ? node25297 : node25290;
														assign node25290 = (inp[3]) ? node25294 : node25291;
															assign node25291 = (inp[9]) ? 4'b1010 : 4'b1110;
															assign node25294 = (inp[2]) ? 4'b1100 : 4'b1000;
														assign node25297 = (inp[9]) ? 4'b1100 : 4'b1000;
												assign node25300 = (inp[3]) ? node25310 : node25301;
													assign node25301 = (inp[9]) ? node25305 : node25302;
														assign node25302 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node25305 = (inp[4]) ? node25307 : 4'b1000;
															assign node25307 = (inp[5]) ? 4'b1110 : 4'b1100;
													assign node25310 = (inp[5]) ? 4'b1110 : node25311;
														assign node25311 = (inp[4]) ? node25315 : node25312;
															assign node25312 = (inp[9]) ? 4'b1000 : 4'b1100;
															assign node25315 = (inp[9]) ? 4'b1110 : 4'b1000;
											assign node25319 = (inp[15]) ? node25351 : node25320;
												assign node25320 = (inp[5]) ? node25332 : node25321;
													assign node25321 = (inp[3]) ? node25327 : node25322;
														assign node25322 = (inp[9]) ? 4'b1010 : node25323;
															assign node25323 = (inp[4]) ? 4'b1110 : 4'b1010;
														assign node25327 = (inp[4]) ? node25329 : 4'b1010;
															assign node25329 = (inp[9]) ? 4'b1000 : 4'b1100;
													assign node25332 = (inp[2]) ? node25340 : node25333;
														assign node25333 = (inp[9]) ? node25337 : node25334;
															assign node25334 = (inp[4]) ? 4'b1100 : 4'b1000;
															assign node25337 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node25340 = (inp[3]) ? node25344 : node25341;
															assign node25341 = (inp[4]) ? 4'b1000 : 4'b1010;
															assign node25344 = (inp[9]) ? node25348 : node25345;
																assign node25345 = (inp[4]) ? 4'b1100 : 4'b1000;
																assign node25348 = (inp[4]) ? 4'b1000 : 4'b1100;
												assign node25351 = (inp[5]) ? node25373 : node25352;
													assign node25352 = (inp[3]) ? node25366 : node25353;
														assign node25353 = (inp[2]) ? node25361 : node25354;
															assign node25354 = (inp[4]) ? node25358 : node25355;
																assign node25355 = (inp[9]) ? 4'b1100 : 4'b1000;
																assign node25358 = (inp[9]) ? 4'b1000 : 4'b1100;
															assign node25361 = (inp[4]) ? node25363 : 4'b1100;
																assign node25363 = (inp[9]) ? 4'b1000 : 4'b1100;
														assign node25366 = (inp[9]) ? node25370 : node25367;
															assign node25367 = (inp[4]) ? 4'b1110 : 4'b1000;
															assign node25370 = (inp[4]) ? 4'b1010 : 4'b1110;
													assign node25373 = (inp[4]) ? node25379 : node25374;
														assign node25374 = (inp[9]) ? 4'b1110 : node25375;
															assign node25375 = (inp[3]) ? 4'b1010 : 4'b1000;
														assign node25379 = (inp[9]) ? 4'b1010 : 4'b1110;
										assign node25382 = (inp[4]) ? node25432 : node25383;
											assign node25383 = (inp[15]) ? node25411 : node25384;
												assign node25384 = (inp[3]) ? node25396 : node25385;
													assign node25385 = (inp[5]) ? node25387 : 4'b1100;
														assign node25387 = (inp[2]) ? 4'b1000 : node25388;
															assign node25388 = (inp[9]) ? node25392 : node25389;
																assign node25389 = (inp[12]) ? 4'b1000 : 4'b1100;
																assign node25392 = (inp[12]) ? 4'b1110 : 4'b1000;
													assign node25396 = (inp[5]) ? node25404 : node25397;
														assign node25397 = (inp[9]) ? node25401 : node25398;
															assign node25398 = (inp[12]) ? 4'b1000 : 4'b1100;
															assign node25401 = (inp[12]) ? 4'b1110 : 4'b1000;
														assign node25404 = (inp[12]) ? node25408 : node25405;
															assign node25405 = (inp[9]) ? 4'b1010 : 4'b1110;
															assign node25408 = (inp[9]) ? 4'b1110 : 4'b1010;
												assign node25411 = (inp[3]) ? node25421 : node25412;
													assign node25412 = (inp[9]) ? node25416 : node25413;
														assign node25413 = (inp[12]) ? 4'b1010 : 4'b1110;
														assign node25416 = (inp[12]) ? node25418 : 4'b1010;
															assign node25418 = (inp[5]) ? 4'b1100 : 4'b1110;
													assign node25421 = (inp[5]) ? node25427 : node25422;
														assign node25422 = (inp[12]) ? node25424 : 4'b1010;
															assign node25424 = (inp[9]) ? 4'b1100 : 4'b1010;
														assign node25427 = (inp[9]) ? 4'b1100 : node25428;
															assign node25428 = (inp[12]) ? 4'b1000 : 4'b1100;
											assign node25432 = (inp[15]) ? node25464 : node25433;
												assign node25433 = (inp[5]) ? node25455 : node25434;
													assign node25434 = (inp[3]) ? node25448 : node25435;
														assign node25435 = (inp[2]) ? node25441 : node25436;
															assign node25436 = (inp[9]) ? node25438 : 4'b1100;
																assign node25438 = (inp[12]) ? 4'b1000 : 4'b1100;
															assign node25441 = (inp[12]) ? node25445 : node25442;
																assign node25442 = (inp[9]) ? 4'b1100 : 4'b1000;
																assign node25445 = (inp[9]) ? 4'b1000 : 4'b1100;
														assign node25448 = (inp[9]) ? node25452 : node25449;
															assign node25449 = (inp[12]) ? 4'b1110 : 4'b1000;
															assign node25452 = (inp[12]) ? 4'b1010 : 4'b1110;
													assign node25455 = (inp[9]) ? node25461 : node25456;
														assign node25456 = (inp[12]) ? 4'b1110 : node25457;
															assign node25457 = (inp[3]) ? 4'b1010 : 4'b1000;
														assign node25461 = (inp[12]) ? 4'b1010 : 4'b1110;
												assign node25464 = (inp[5]) ? node25478 : node25465;
													assign node25465 = (inp[3]) ? node25471 : node25466;
														assign node25466 = (inp[12]) ? 4'b1110 : node25467;
															assign node25467 = (inp[9]) ? 4'b1110 : 4'b1010;
														assign node25471 = (inp[9]) ? node25475 : node25472;
															assign node25472 = (inp[12]) ? 4'b1100 : 4'b1010;
															assign node25475 = (inp[12]) ? 4'b1000 : 4'b1100;
													assign node25478 = (inp[2]) ? node25484 : node25479;
														assign node25479 = (inp[12]) ? 4'b1100 : node25480;
															assign node25480 = (inp[9]) ? 4'b1100 : 4'b1000;
														assign node25484 = (inp[12]) ? node25490 : node25485;
															assign node25485 = (inp[9]) ? 4'b1100 : node25486;
																assign node25486 = (inp[3]) ? 4'b1000 : 4'b1010;
															assign node25490 = (inp[9]) ? 4'b1000 : 4'b1100;
								assign node25493 = (inp[2]) ? node25731 : node25494;
									assign node25494 = (inp[14]) ? node25614 : node25495;
										assign node25495 = (inp[4]) ? node25551 : node25496;
											assign node25496 = (inp[12]) ? node25524 : node25497;
												assign node25497 = (inp[9]) ? node25503 : node25498;
													assign node25498 = (inp[5]) ? node25500 : 4'b1110;
														assign node25500 = (inp[15]) ? 4'b1100 : 4'b1110;
													assign node25503 = (inp[15]) ? node25515 : node25504;
														assign node25504 = (inp[0]) ? node25510 : node25505;
															assign node25505 = (inp[3]) ? node25507 : 4'b1010;
																assign node25507 = (inp[5]) ? 4'b1000 : 4'b1010;
															assign node25510 = (inp[3]) ? node25512 : 4'b1000;
																assign node25512 = (inp[5]) ? 4'b1010 : 4'b1000;
														assign node25515 = (inp[0]) ? node25521 : node25516;
															assign node25516 = (inp[5]) ? node25518 : 4'b1000;
																assign node25518 = (inp[3]) ? 4'b1010 : 4'b1000;
															assign node25521 = (inp[3]) ? 4'b1000 : 4'b1010;
												assign node25524 = (inp[9]) ? node25538 : node25525;
													assign node25525 = (inp[15]) ? node25533 : node25526;
														assign node25526 = (inp[0]) ? node25528 : 4'b1010;
															assign node25528 = (inp[3]) ? node25530 : 4'b1000;
																assign node25530 = (inp[5]) ? 4'b1010 : 4'b1000;
														assign node25533 = (inp[5]) ? 4'b1000 : node25534;
															assign node25534 = (inp[0]) ? 4'b1010 : 4'b1000;
													assign node25538 = (inp[15]) ? node25546 : node25539;
														assign node25539 = (inp[5]) ? 4'b1100 : node25540;
															assign node25540 = (inp[3]) ? 4'b1100 : node25541;
																assign node25541 = (inp[0]) ? 4'b1100 : 4'b1110;
														assign node25546 = (inp[0]) ? node25548 : 4'b1110;
															assign node25548 = (inp[5]) ? 4'b1100 : 4'b1110;
											assign node25551 = (inp[9]) ? node25583 : node25552;
												assign node25552 = (inp[12]) ? node25570 : node25553;
													assign node25553 = (inp[15]) ? node25565 : node25554;
														assign node25554 = (inp[0]) ? node25560 : node25555;
															assign node25555 = (inp[5]) ? node25557 : 4'b1010;
																assign node25557 = (inp[3]) ? 4'b1000 : 4'b1010;
															assign node25560 = (inp[3]) ? node25562 : 4'b1000;
																assign node25562 = (inp[5]) ? 4'b1010 : 4'b1000;
														assign node25565 = (inp[0]) ? 4'b1010 : node25566;
															assign node25566 = (inp[5]) ? 4'b1010 : 4'b1000;
													assign node25570 = (inp[0]) ? node25578 : node25571;
														assign node25571 = (inp[15]) ? node25573 : 4'b1110;
															assign node25573 = (inp[3]) ? 4'b1110 : node25574;
																assign node25574 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node25578 = (inp[15]) ? 4'b1100 : node25579;
															assign node25579 = (inp[3]) ? 4'b1110 : 4'b1100;
												assign node25583 = (inp[12]) ? node25605 : node25584;
													assign node25584 = (inp[0]) ? node25596 : node25585;
														assign node25585 = (inp[15]) ? node25591 : node25586;
															assign node25586 = (inp[5]) ? 4'b1100 : node25587;
																assign node25587 = (inp[3]) ? 4'b1100 : 4'b1110;
															assign node25591 = (inp[5]) ? 4'b1110 : node25592;
																assign node25592 = (inp[3]) ? 4'b1110 : 4'b1100;
														assign node25596 = (inp[15]) ? node25600 : node25597;
															assign node25597 = (inp[5]) ? 4'b1110 : 4'b1100;
															assign node25600 = (inp[5]) ? 4'b1100 : node25601;
																assign node25601 = (inp[3]) ? 4'b1100 : 4'b1110;
													assign node25605 = (inp[3]) ? 4'b1010 : node25606;
														assign node25606 = (inp[15]) ? 4'b1000 : node25607;
															assign node25607 = (inp[0]) ? 4'b1010 : node25608;
																assign node25608 = (inp[5]) ? 4'b1000 : 4'b1010;
										assign node25614 = (inp[9]) ? node25668 : node25615;
											assign node25615 = (inp[12]) ? node25645 : node25616;
												assign node25616 = (inp[4]) ? node25628 : node25617;
													assign node25617 = (inp[0]) ? node25621 : node25618;
														assign node25618 = (inp[15]) ? 4'b0101 : 4'b0111;
														assign node25621 = (inp[15]) ? node25623 : 4'b0101;
															assign node25623 = (inp[5]) ? node25625 : 4'b0111;
																assign node25625 = (inp[3]) ? 4'b0101 : 4'b0111;
													assign node25628 = (inp[5]) ? node25634 : node25629;
														assign node25629 = (inp[0]) ? node25631 : 4'b0011;
															assign node25631 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node25634 = (inp[3]) ? node25640 : node25635;
															assign node25635 = (inp[0]) ? node25637 : 4'b0001;
																assign node25637 = (inp[15]) ? 4'b0011 : 4'b0001;
															assign node25640 = (inp[0]) ? node25642 : 4'b0011;
																assign node25642 = (inp[15]) ? 4'b0001 : 4'b0011;
												assign node25645 = (inp[4]) ? node25655 : node25646;
													assign node25646 = (inp[3]) ? 4'b0011 : node25647;
														assign node25647 = (inp[0]) ? node25651 : node25648;
															assign node25648 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node25651 = (inp[15]) ? 4'b0011 : 4'b0001;
													assign node25655 = (inp[5]) ? node25661 : node25656;
														assign node25656 = (inp[15]) ? node25658 : 4'b0111;
															assign node25658 = (inp[0]) ? 4'b0101 : 4'b0111;
														assign node25661 = (inp[0]) ? node25665 : node25662;
															assign node25662 = (inp[15]) ? 4'b0111 : 4'b0101;
															assign node25665 = (inp[15]) ? 4'b0101 : 4'b0111;
											assign node25668 = (inp[3]) ? node25706 : node25669;
												assign node25669 = (inp[5]) ? node25687 : node25670;
													assign node25670 = (inp[4]) ? node25678 : node25671;
														assign node25671 = (inp[12]) ? node25673 : 4'b0001;
															assign node25673 = (inp[15]) ? 4'b0101 : node25674;
																assign node25674 = (inp[0]) ? 4'b0101 : 4'b0111;
														assign node25678 = (inp[12]) ? 4'b0011 : node25679;
															assign node25679 = (inp[0]) ? node25683 : node25680;
																assign node25680 = (inp[15]) ? 4'b0101 : 4'b0111;
																assign node25683 = (inp[15]) ? 4'b0111 : 4'b0101;
													assign node25687 = (inp[0]) ? node25695 : node25688;
														assign node25688 = (inp[15]) ? 4'b0111 : node25689;
															assign node25689 = (inp[12]) ? node25691 : 4'b0101;
																assign node25691 = (inp[4]) ? 4'b0001 : 4'b0101;
														assign node25695 = (inp[4]) ? node25703 : node25696;
															assign node25696 = (inp[12]) ? node25700 : node25697;
																assign node25697 = (inp[15]) ? 4'b0011 : 4'b0001;
																assign node25700 = (inp[15]) ? 4'b0101 : 4'b0111;
															assign node25703 = (inp[12]) ? 4'b0001 : 4'b0101;
												assign node25706 = (inp[12]) ? node25718 : node25707;
													assign node25707 = (inp[4]) ? node25715 : node25708;
														assign node25708 = (inp[0]) ? node25710 : 4'b0001;
															assign node25710 = (inp[5]) ? node25712 : 4'b0001;
																assign node25712 = (inp[15]) ? 4'b0001 : 4'b0011;
														assign node25715 = (inp[0]) ? 4'b0111 : 4'b0101;
													assign node25718 = (inp[4]) ? node25722 : node25719;
														assign node25719 = (inp[0]) ? 4'b0101 : 4'b0111;
														assign node25722 = (inp[5]) ? 4'b0001 : node25723;
															assign node25723 = (inp[0]) ? node25727 : node25724;
																assign node25724 = (inp[15]) ? 4'b0011 : 4'b0001;
																assign node25727 = (inp[15]) ? 4'b0001 : 4'b0011;
									assign node25731 = (inp[12]) ? node25823 : node25732;
										assign node25732 = (inp[4]) ? node25774 : node25733;
											assign node25733 = (inp[9]) ? node25759 : node25734;
												assign node25734 = (inp[3]) ? node25750 : node25735;
													assign node25735 = (inp[14]) ? node25743 : node25736;
														assign node25736 = (inp[15]) ? node25740 : node25737;
															assign node25737 = (inp[0]) ? 4'b0101 : 4'b0111;
															assign node25740 = (inp[0]) ? 4'b0111 : 4'b0101;
														assign node25743 = (inp[15]) ? node25747 : node25744;
															assign node25744 = (inp[0]) ? 4'b0101 : 4'b0111;
															assign node25747 = (inp[0]) ? 4'b0111 : 4'b0101;
													assign node25750 = (inp[15]) ? 4'b0101 : node25751;
														assign node25751 = (inp[0]) ? node25755 : node25752;
															assign node25752 = (inp[5]) ? 4'b0101 : 4'b0111;
															assign node25755 = (inp[5]) ? 4'b0111 : 4'b0101;
												assign node25759 = (inp[0]) ? node25767 : node25760;
													assign node25760 = (inp[15]) ? 4'b0001 : node25761;
														assign node25761 = (inp[3]) ? node25763 : 4'b0011;
															assign node25763 = (inp[5]) ? 4'b0001 : 4'b0011;
													assign node25767 = (inp[15]) ? node25769 : 4'b0001;
														assign node25769 = (inp[3]) ? node25771 : 4'b0011;
															assign node25771 = (inp[5]) ? 4'b0001 : 4'b0011;
											assign node25774 = (inp[9]) ? node25798 : node25775;
												assign node25775 = (inp[0]) ? node25787 : node25776;
													assign node25776 = (inp[15]) ? node25782 : node25777;
														assign node25777 = (inp[5]) ? node25779 : 4'b0011;
															assign node25779 = (inp[3]) ? 4'b0001 : 4'b0011;
														assign node25782 = (inp[5]) ? node25784 : 4'b0001;
															assign node25784 = (inp[14]) ? 4'b0011 : 4'b0001;
													assign node25787 = (inp[15]) ? node25793 : node25788;
														assign node25788 = (inp[3]) ? node25790 : 4'b0001;
															assign node25790 = (inp[5]) ? 4'b0011 : 4'b0001;
														assign node25793 = (inp[3]) ? node25795 : 4'b0011;
															assign node25795 = (inp[5]) ? 4'b0001 : 4'b0011;
												assign node25798 = (inp[14]) ? node25810 : node25799;
													assign node25799 = (inp[5]) ? node25805 : node25800;
														assign node25800 = (inp[15]) ? node25802 : 4'b0111;
															assign node25802 = (inp[0]) ? 4'b0101 : 4'b0111;
														assign node25805 = (inp[15]) ? 4'b0111 : node25806;
															assign node25806 = (inp[0]) ? 4'b0111 : 4'b0101;
													assign node25810 = (inp[5]) ? 4'b0101 : node25811;
														assign node25811 = (inp[15]) ? node25817 : node25812;
															assign node25812 = (inp[3]) ? node25814 : 4'b0101;
																assign node25814 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node25817 = (inp[0]) ? node25819 : 4'b0111;
																assign node25819 = (inp[3]) ? 4'b0101 : 4'b0111;
										assign node25823 = (inp[5]) ? node25885 : node25824;
											assign node25824 = (inp[0]) ? node25856 : node25825;
												assign node25825 = (inp[15]) ? node25841 : node25826;
													assign node25826 = (inp[3]) ? node25834 : node25827;
														assign node25827 = (inp[9]) ? node25831 : node25828;
															assign node25828 = (inp[4]) ? 4'b0111 : 4'b0011;
															assign node25831 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node25834 = (inp[9]) ? node25838 : node25835;
															assign node25835 = (inp[4]) ? 4'b0101 : 4'b0011;
															assign node25838 = (inp[4]) ? 4'b0001 : 4'b0101;
													assign node25841 = (inp[3]) ? node25849 : node25842;
														assign node25842 = (inp[14]) ? node25844 : 4'b0101;
															assign node25844 = (inp[9]) ? 4'b0001 : node25845;
																assign node25845 = (inp[4]) ? 4'b0101 : 4'b0001;
														assign node25849 = (inp[4]) ? node25853 : node25850;
															assign node25850 = (inp[9]) ? 4'b0111 : 4'b0001;
															assign node25853 = (inp[9]) ? 4'b0011 : 4'b0111;
												assign node25856 = (inp[15]) ? node25870 : node25857;
													assign node25857 = (inp[3]) ? node25863 : node25858;
														assign node25858 = (inp[9]) ? node25860 : 4'b0101;
															assign node25860 = (inp[4]) ? 4'b0001 : 4'b0101;
														assign node25863 = (inp[9]) ? node25867 : node25864;
															assign node25864 = (inp[4]) ? 4'b0111 : 4'b0001;
															assign node25867 = (inp[4]) ? 4'b0011 : 4'b0111;
													assign node25870 = (inp[3]) ? node25878 : node25871;
														assign node25871 = (inp[4]) ? node25875 : node25872;
															assign node25872 = (inp[9]) ? 4'b0111 : 4'b0011;
															assign node25875 = (inp[9]) ? 4'b0011 : 4'b0111;
														assign node25878 = (inp[9]) ? node25882 : node25879;
															assign node25879 = (inp[4]) ? 4'b0101 : 4'b0011;
															assign node25882 = (inp[4]) ? 4'b0001 : 4'b0101;
											assign node25885 = (inp[4]) ? node25917 : node25886;
												assign node25886 = (inp[9]) ? node25906 : node25887;
													assign node25887 = (inp[14]) ? node25897 : node25888;
														assign node25888 = (inp[3]) ? 4'b0011 : node25889;
															assign node25889 = (inp[0]) ? node25893 : node25890;
																assign node25890 = (inp[15]) ? 4'b0001 : 4'b0011;
																assign node25893 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node25897 = (inp[0]) ? node25899 : 4'b0001;
															assign node25899 = (inp[15]) ? node25903 : node25900;
																assign node25900 = (inp[3]) ? 4'b0011 : 4'b0001;
																assign node25903 = (inp[3]) ? 4'b0001 : 4'b0011;
													assign node25906 = (inp[3]) ? node25912 : node25907;
														assign node25907 = (inp[15]) ? node25909 : 4'b0101;
															assign node25909 = (inp[0]) ? 4'b0101 : 4'b0111;
														assign node25912 = (inp[0]) ? node25914 : 4'b0111;
															assign node25914 = (inp[15]) ? 4'b0101 : 4'b0111;
												assign node25917 = (inp[9]) ? node25931 : node25918;
													assign node25918 = (inp[3]) ? node25924 : node25919;
														assign node25919 = (inp[0]) ? node25921 : 4'b0101;
															assign node25921 = (inp[15]) ? 4'b0101 : 4'b0111;
														assign node25924 = (inp[14]) ? 4'b0111 : node25925;
															assign node25925 = (inp[0]) ? 4'b0101 : node25926;
																assign node25926 = (inp[15]) ? 4'b0111 : 4'b0101;
													assign node25931 = (inp[3]) ? 4'b0001 : node25932;
														assign node25932 = (inp[15]) ? node25936 : node25933;
															assign node25933 = (inp[0]) ? 4'b0011 : 4'b0001;
															assign node25936 = (inp[0]) ? 4'b0001 : 4'b0011;
							assign node25940 = (inp[7]) ? node26522 : node25941;
								assign node25941 = (inp[14]) ? node26203 : node25942;
									assign node25942 = (inp[2]) ? node26084 : node25943;
										assign node25943 = (inp[15]) ? node26027 : node25944;
											assign node25944 = (inp[3]) ? node25990 : node25945;
												assign node25945 = (inp[0]) ? node25965 : node25946;
													assign node25946 = (inp[9]) ? node25956 : node25947;
														assign node25947 = (inp[5]) ? 4'b1010 : node25948;
															assign node25948 = (inp[12]) ? node25952 : node25949;
																assign node25949 = (inp[4]) ? 4'b1010 : 4'b1110;
																assign node25952 = (inp[4]) ? 4'b1110 : 4'b1010;
														assign node25956 = (inp[4]) ? node25962 : node25957;
															assign node25957 = (inp[12]) ? node25959 : 4'b1010;
																assign node25959 = (inp[5]) ? 4'b1100 : 4'b1110;
															assign node25962 = (inp[12]) ? 4'b1000 : 4'b1100;
													assign node25965 = (inp[5]) ? node25979 : node25966;
														assign node25966 = (inp[9]) ? node25974 : node25967;
															assign node25967 = (inp[4]) ? node25971 : node25968;
																assign node25968 = (inp[12]) ? 4'b1000 : 4'b1100;
																assign node25971 = (inp[12]) ? 4'b1100 : 4'b1000;
															assign node25974 = (inp[4]) ? 4'b1100 : node25975;
																assign node25975 = (inp[12]) ? 4'b1100 : 4'b1000;
														assign node25979 = (inp[9]) ? node25985 : node25980;
															assign node25980 = (inp[4]) ? 4'b1110 : node25981;
																assign node25981 = (inp[12]) ? 4'b1000 : 4'b1100;
															assign node25985 = (inp[12]) ? node25987 : 4'b1110;
																assign node25987 = (inp[4]) ? 4'b1010 : 4'b1110;
												assign node25990 = (inp[0]) ? node26010 : node25991;
													assign node25991 = (inp[4]) ? node26005 : node25992;
														assign node25992 = (inp[5]) ? node25998 : node25993;
															assign node25993 = (inp[9]) ? node25995 : 4'b1010;
																assign node25995 = (inp[12]) ? 4'b1100 : 4'b1010;
															assign node25998 = (inp[12]) ? node26002 : node25999;
																assign node25999 = (inp[9]) ? 4'b1000 : 4'b1100;
																assign node26002 = (inp[9]) ? 4'b1100 : 4'b1000;
														assign node26005 = (inp[9]) ? node26007 : 4'b1100;
															assign node26007 = (inp[12]) ? 4'b1000 : 4'b1100;
													assign node26010 = (inp[9]) ? node26022 : node26011;
														assign node26011 = (inp[5]) ? node26017 : node26012;
															assign node26012 = (inp[12]) ? 4'b1000 : node26013;
																assign node26013 = (inp[4]) ? 4'b1000 : 4'b1100;
															assign node26017 = (inp[12]) ? 4'b1110 : node26018;
																assign node26018 = (inp[4]) ? 4'b1010 : 4'b1110;
														assign node26022 = (inp[12]) ? node26024 : 4'b1110;
															assign node26024 = (inp[4]) ? 4'b1010 : 4'b1110;
											assign node26027 = (inp[12]) ? node26049 : node26028;
												assign node26028 = (inp[4]) ? node26040 : node26029;
													assign node26029 = (inp[9]) ? node26037 : node26030;
														assign node26030 = (inp[3]) ? node26032 : 4'b1110;
															assign node26032 = (inp[0]) ? 4'b1100 : node26033;
																assign node26033 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node26037 = (inp[0]) ? 4'b1010 : 4'b1000;
													assign node26040 = (inp[9]) ? 4'b1110 : node26041;
														assign node26041 = (inp[3]) ? node26043 : 4'b1010;
															assign node26043 = (inp[5]) ? node26045 : 4'b1010;
																assign node26045 = (inp[0]) ? 4'b1000 : 4'b1010;
												assign node26049 = (inp[0]) ? node26065 : node26050;
													assign node26050 = (inp[3]) ? node26058 : node26051;
														assign node26051 = (inp[4]) ? node26053 : 4'b1000;
															assign node26053 = (inp[9]) ? 4'b1000 : node26054;
																assign node26054 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node26058 = (inp[9]) ? node26062 : node26059;
															assign node26059 = (inp[4]) ? 4'b1110 : 4'b1010;
															assign node26062 = (inp[4]) ? 4'b1010 : 4'b1110;
													assign node26065 = (inp[5]) ? node26075 : node26066;
														assign node26066 = (inp[3]) ? 4'b1000 : node26067;
															assign node26067 = (inp[4]) ? node26071 : node26068;
																assign node26068 = (inp[9]) ? 4'b1110 : 4'b1010;
																assign node26071 = (inp[9]) ? 4'b1010 : 4'b1110;
														assign node26075 = (inp[4]) ? node26081 : node26076;
															assign node26076 = (inp[9]) ? 4'b1100 : node26077;
																assign node26077 = (inp[3]) ? 4'b1000 : 4'b1010;
															assign node26081 = (inp[9]) ? 4'b1000 : 4'b1100;
										assign node26084 = (inp[0]) ? node26150 : node26085;
											assign node26085 = (inp[15]) ? node26119 : node26086;
												assign node26086 = (inp[5]) ? node26102 : node26087;
													assign node26087 = (inp[3]) ? node26089 : 4'b0011;
														assign node26089 = (inp[4]) ? node26095 : node26090;
															assign node26090 = (inp[12]) ? node26092 : 4'b0011;
																assign node26092 = (inp[9]) ? 4'b0101 : 4'b0011;
															assign node26095 = (inp[9]) ? node26099 : node26096;
																assign node26096 = (inp[12]) ? 4'b0101 : 4'b0011;
																assign node26099 = (inp[12]) ? 4'b0001 : 4'b0101;
													assign node26102 = (inp[3]) ? node26110 : node26103;
														assign node26103 = (inp[9]) ? 4'b0101 : node26104;
															assign node26104 = (inp[4]) ? 4'b0101 : node26105;
																assign node26105 = (inp[12]) ? 4'b0011 : 4'b0111;
														assign node26110 = (inp[4]) ? 4'b0001 : node26111;
															assign node26111 = (inp[12]) ? node26115 : node26112;
																assign node26112 = (inp[9]) ? 4'b0001 : 4'b0101;
																assign node26115 = (inp[9]) ? 4'b0101 : 4'b0001;
												assign node26119 = (inp[5]) ? node26139 : node26120;
													assign node26120 = (inp[3]) ? node26130 : node26121;
														assign node26121 = (inp[9]) ? 4'b0101 : node26122;
															assign node26122 = (inp[12]) ? node26126 : node26123;
																assign node26123 = (inp[4]) ? 4'b0001 : 4'b0101;
																assign node26126 = (inp[4]) ? 4'b0101 : 4'b0001;
														assign node26130 = (inp[12]) ? 4'b0111 : node26131;
															assign node26131 = (inp[9]) ? node26135 : node26132;
																assign node26132 = (inp[4]) ? 4'b0001 : 4'b0101;
																assign node26135 = (inp[4]) ? 4'b0111 : 4'b0001;
													assign node26139 = (inp[9]) ? node26145 : node26140;
														assign node26140 = (inp[12]) ? 4'b0111 : node26141;
															assign node26141 = (inp[3]) ? 4'b0111 : 4'b0101;
														assign node26145 = (inp[4]) ? node26147 : 4'b0011;
															assign node26147 = (inp[12]) ? 4'b0011 : 4'b0111;
											assign node26150 = (inp[12]) ? node26166 : node26151;
												assign node26151 = (inp[5]) ? node26155 : node26152;
													assign node26152 = (inp[15]) ? 4'b0011 : 4'b0001;
													assign node26155 = (inp[15]) ? node26157 : 4'b0111;
														assign node26157 = (inp[3]) ? 4'b0001 : node26158;
															assign node26158 = (inp[9]) ? node26162 : node26159;
																assign node26159 = (inp[4]) ? 4'b0011 : 4'b0111;
																assign node26162 = (inp[4]) ? 4'b0101 : 4'b0011;
												assign node26166 = (inp[15]) ? node26184 : node26167;
													assign node26167 = (inp[3]) ? node26175 : node26168;
														assign node26168 = (inp[5]) ? node26170 : 4'b0001;
															assign node26170 = (inp[9]) ? 4'b0111 : node26171;
																assign node26171 = (inp[4]) ? 4'b0111 : 4'b0001;
														assign node26175 = (inp[5]) ? node26177 : 4'b0111;
															assign node26177 = (inp[4]) ? node26181 : node26178;
																assign node26178 = (inp[9]) ? 4'b0111 : 4'b0011;
																assign node26181 = (inp[9]) ? 4'b0011 : 4'b0111;
													assign node26184 = (inp[5]) ? node26196 : node26185;
														assign node26185 = (inp[3]) ? node26193 : node26186;
															assign node26186 = (inp[4]) ? node26190 : node26187;
																assign node26187 = (inp[9]) ? 4'b0111 : 4'b0011;
																assign node26190 = (inp[9]) ? 4'b0011 : 4'b0111;
															assign node26193 = (inp[4]) ? 4'b0101 : 4'b0011;
														assign node26196 = (inp[9]) ? node26200 : node26197;
															assign node26197 = (inp[3]) ? 4'b0001 : 4'b0011;
															assign node26200 = (inp[4]) ? 4'b0001 : 4'b0101;
									assign node26203 = (inp[9]) ? node26359 : node26204;
										assign node26204 = (inp[2]) ? node26278 : node26205;
											assign node26205 = (inp[0]) ? node26239 : node26206;
												assign node26206 = (inp[15]) ? node26220 : node26207;
													assign node26207 = (inp[3]) ? node26215 : node26208;
														assign node26208 = (inp[12]) ? node26212 : node26209;
															assign node26209 = (inp[4]) ? 4'b0011 : 4'b0111;
															assign node26212 = (inp[4]) ? 4'b0111 : 4'b0011;
														assign node26215 = (inp[12]) ? 4'b0101 : node26216;
															assign node26216 = (inp[5]) ? 4'b0001 : 4'b0011;
													assign node26220 = (inp[4]) ? node26228 : node26221;
														assign node26221 = (inp[12]) ? node26223 : 4'b0101;
															assign node26223 = (inp[5]) ? node26225 : 4'b0001;
																assign node26225 = (inp[3]) ? 4'b0011 : 4'b0001;
														assign node26228 = (inp[12]) ? node26234 : node26229;
															assign node26229 = (inp[3]) ? node26231 : 4'b0001;
																assign node26231 = (inp[5]) ? 4'b0011 : 4'b0001;
															assign node26234 = (inp[5]) ? 4'b0111 : node26235;
																assign node26235 = (inp[3]) ? 4'b0111 : 4'b0101;
												assign node26239 = (inp[15]) ? node26259 : node26240;
													assign node26240 = (inp[3]) ? node26250 : node26241;
														assign node26241 = (inp[4]) ? node26245 : node26242;
															assign node26242 = (inp[12]) ? 4'b0001 : 4'b0101;
															assign node26245 = (inp[12]) ? node26247 : 4'b0001;
																assign node26247 = (inp[5]) ? 4'b0111 : 4'b0101;
														assign node26250 = (inp[5]) ? node26256 : node26251;
															assign node26251 = (inp[12]) ? node26253 : 4'b0001;
																assign node26253 = (inp[4]) ? 4'b0111 : 4'b0001;
															assign node26256 = (inp[4]) ? 4'b0011 : 4'b0111;
													assign node26259 = (inp[3]) ? node26267 : node26260;
														assign node26260 = (inp[12]) ? node26264 : node26261;
															assign node26261 = (inp[4]) ? 4'b0011 : 4'b0111;
															assign node26264 = (inp[4]) ? 4'b0101 : 4'b0011;
														assign node26267 = (inp[5]) ? node26273 : node26268;
															assign node26268 = (inp[4]) ? 4'b0101 : node26269;
																assign node26269 = (inp[12]) ? 4'b0011 : 4'b0111;
															assign node26273 = (inp[4]) ? 4'b0001 : node26274;
																assign node26274 = (inp[12]) ? 4'b0001 : 4'b0101;
											assign node26278 = (inp[5]) ? node26308 : node26279;
												assign node26279 = (inp[3]) ? node26295 : node26280;
													assign node26280 = (inp[4]) ? node26290 : node26281;
														assign node26281 = (inp[12]) ? 4'b0011 : node26282;
															assign node26282 = (inp[0]) ? node26286 : node26283;
																assign node26283 = (inp[15]) ? 4'b0101 : 4'b0111;
																assign node26286 = (inp[15]) ? 4'b0111 : 4'b0101;
														assign node26290 = (inp[12]) ? 4'b0101 : node26291;
															assign node26291 = (inp[15]) ? 4'b0001 : 4'b0011;
													assign node26295 = (inp[4]) ? node26305 : node26296;
														assign node26296 = (inp[12]) ? node26298 : 4'b0111;
															assign node26298 = (inp[0]) ? node26302 : node26299;
																assign node26299 = (inp[15]) ? 4'b0001 : 4'b0011;
																assign node26302 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node26305 = (inp[12]) ? 4'b0111 : 4'b0011;
												assign node26308 = (inp[15]) ? node26340 : node26309;
													assign node26309 = (inp[0]) ? node26325 : node26310;
														assign node26310 = (inp[3]) ? node26318 : node26311;
															assign node26311 = (inp[4]) ? node26315 : node26312;
																assign node26312 = (inp[12]) ? 4'b0011 : 4'b0111;
																assign node26315 = (inp[12]) ? 4'b0101 : 4'b0011;
															assign node26318 = (inp[4]) ? node26322 : node26319;
																assign node26319 = (inp[12]) ? 4'b0001 : 4'b0101;
																assign node26322 = (inp[12]) ? 4'b0101 : 4'b0001;
														assign node26325 = (inp[3]) ? node26333 : node26326;
															assign node26326 = (inp[12]) ? node26330 : node26327;
																assign node26327 = (inp[4]) ? 4'b0001 : 4'b0101;
																assign node26330 = (inp[4]) ? 4'b0111 : 4'b0001;
															assign node26333 = (inp[12]) ? node26337 : node26334;
																assign node26334 = (inp[4]) ? 4'b0011 : 4'b0111;
																assign node26337 = (inp[4]) ? 4'b0111 : 4'b0011;
													assign node26340 = (inp[12]) ? node26350 : node26341;
														assign node26341 = (inp[4]) ? 4'b0011 : node26342;
															assign node26342 = (inp[0]) ? node26346 : node26343;
																assign node26343 = (inp[3]) ? 4'b0111 : 4'b0101;
																assign node26346 = (inp[3]) ? 4'b0101 : 4'b0111;
														assign node26350 = (inp[4]) ? node26356 : node26351;
															assign node26351 = (inp[3]) ? 4'b0011 : node26352;
																assign node26352 = (inp[0]) ? 4'b0011 : 4'b0001;
															assign node26356 = (inp[0]) ? 4'b0101 : 4'b0111;
										assign node26359 = (inp[2]) ? node26441 : node26360;
											assign node26360 = (inp[5]) ? node26402 : node26361;
												assign node26361 = (inp[0]) ? node26381 : node26362;
													assign node26362 = (inp[3]) ? node26370 : node26363;
														assign node26363 = (inp[15]) ? node26365 : 4'b0011;
															assign node26365 = (inp[4]) ? 4'b0001 : node26366;
																assign node26366 = (inp[12]) ? 4'b0101 : 4'b0001;
														assign node26370 = (inp[12]) ? node26378 : node26371;
															assign node26371 = (inp[4]) ? node26375 : node26372;
																assign node26372 = (inp[15]) ? 4'b0001 : 4'b0011;
																assign node26375 = (inp[15]) ? 4'b0111 : 4'b0101;
															assign node26378 = (inp[4]) ? 4'b0001 : 4'b0101;
													assign node26381 = (inp[15]) ? node26391 : node26382;
														assign node26382 = (inp[12]) ? node26386 : node26383;
															assign node26383 = (inp[4]) ? 4'b0101 : 4'b0001;
															assign node26386 = (inp[3]) ? node26388 : 4'b0101;
																assign node26388 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node26391 = (inp[3]) ? node26399 : node26392;
															assign node26392 = (inp[12]) ? node26396 : node26393;
																assign node26393 = (inp[4]) ? 4'b0111 : 4'b0011;
																assign node26396 = (inp[4]) ? 4'b0011 : 4'b0111;
															assign node26399 = (inp[12]) ? 4'b0101 : 4'b0011;
												assign node26402 = (inp[3]) ? node26424 : node26403;
													assign node26403 = (inp[0]) ? node26417 : node26404;
														assign node26404 = (inp[15]) ? node26410 : node26405;
															assign node26405 = (inp[12]) ? node26407 : 4'b0101;
																assign node26407 = (inp[4]) ? 4'b0001 : 4'b0101;
															assign node26410 = (inp[4]) ? node26414 : node26411;
																assign node26411 = (inp[12]) ? 4'b0111 : 4'b0001;
																assign node26414 = (inp[12]) ? 4'b0011 : 4'b0111;
														assign node26417 = (inp[15]) ? 4'b0101 : node26418;
															assign node26418 = (inp[4]) ? 4'b0111 : node26419;
																assign node26419 = (inp[12]) ? 4'b0111 : 4'b0001;
													assign node26424 = (inp[0]) ? node26432 : node26425;
														assign node26425 = (inp[15]) ? node26427 : 4'b0101;
															assign node26427 = (inp[4]) ? 4'b0111 : node26428;
																assign node26428 = (inp[12]) ? 4'b0111 : 4'b0011;
														assign node26432 = (inp[15]) ? node26438 : node26433;
															assign node26433 = (inp[12]) ? node26435 : 4'b0011;
																assign node26435 = (inp[4]) ? 4'b0011 : 4'b0111;
															assign node26438 = (inp[4]) ? 4'b0001 : 4'b0101;
											assign node26441 = (inp[0]) ? node26485 : node26442;
												assign node26442 = (inp[15]) ? node26462 : node26443;
													assign node26443 = (inp[5]) ? node26453 : node26444;
														assign node26444 = (inp[4]) ? node26448 : node26445;
															assign node26445 = (inp[12]) ? 4'b0111 : 4'b0011;
															assign node26448 = (inp[12]) ? node26450 : 4'b0101;
																assign node26450 = (inp[3]) ? 4'b0001 : 4'b0011;
														assign node26453 = (inp[12]) ? node26459 : node26454;
															assign node26454 = (inp[4]) ? 4'b0101 : node26455;
																assign node26455 = (inp[3]) ? 4'b0001 : 4'b0011;
															assign node26459 = (inp[4]) ? 4'b0001 : 4'b0101;
													assign node26462 = (inp[5]) ? node26474 : node26463;
														assign node26463 = (inp[3]) ? node26471 : node26464;
															assign node26464 = (inp[4]) ? node26468 : node26465;
																assign node26465 = (inp[12]) ? 4'b0101 : 4'b0001;
																assign node26468 = (inp[12]) ? 4'b0001 : 4'b0101;
															assign node26471 = (inp[4]) ? 4'b0111 : 4'b0001;
														assign node26474 = (inp[3]) ? node26480 : node26475;
															assign node26475 = (inp[4]) ? 4'b0111 : node26476;
																assign node26476 = (inp[12]) ? 4'b0111 : 4'b0001;
															assign node26480 = (inp[4]) ? node26482 : 4'b0011;
																assign node26482 = (inp[12]) ? 4'b0011 : 4'b0111;
												assign node26485 = (inp[15]) ? node26503 : node26486;
													assign node26486 = (inp[3]) ? node26496 : node26487;
														assign node26487 = (inp[5]) ? node26493 : node26488;
															assign node26488 = (inp[12]) ? node26490 : 4'b0101;
																assign node26490 = (inp[4]) ? 4'b0001 : 4'b0101;
															assign node26493 = (inp[12]) ? 4'b0111 : 4'b0001;
														assign node26496 = (inp[4]) ? 4'b0111 : node26497;
															assign node26497 = (inp[12]) ? 4'b0111 : node26498;
																assign node26498 = (inp[5]) ? 4'b0011 : 4'b0001;
													assign node26503 = (inp[3]) ? node26515 : node26504;
														assign node26504 = (inp[5]) ? node26508 : node26505;
															assign node26505 = (inp[12]) ? 4'b0011 : 4'b0111;
															assign node26508 = (inp[4]) ? node26512 : node26509;
																assign node26509 = (inp[12]) ? 4'b0101 : 4'b0011;
																assign node26512 = (inp[12]) ? 4'b0001 : 4'b0101;
														assign node26515 = (inp[12]) ? node26519 : node26516;
															assign node26516 = (inp[4]) ? 4'b0101 : 4'b0001;
															assign node26519 = (inp[4]) ? 4'b0001 : 4'b0101;
								assign node26522 = (inp[2]) ? node26782 : node26523;
									assign node26523 = (inp[14]) ? node26651 : node26524;
										assign node26524 = (inp[12]) ? node26586 : node26525;
											assign node26525 = (inp[9]) ? node26557 : node26526;
												assign node26526 = (inp[4]) ? node26536 : node26527;
													assign node26527 = (inp[15]) ? node26529 : 4'b0101;
														assign node26529 = (inp[0]) ? 4'b0111 : node26530;
															assign node26530 = (inp[3]) ? node26532 : 4'b0101;
																assign node26532 = (inp[5]) ? 4'b0111 : 4'b0101;
													assign node26536 = (inp[3]) ? node26544 : node26537;
														assign node26537 = (inp[5]) ? node26539 : 4'b0011;
															assign node26539 = (inp[0]) ? node26541 : 4'b0001;
																assign node26541 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node26544 = (inp[15]) ? node26552 : node26545;
															assign node26545 = (inp[0]) ? node26549 : node26546;
																assign node26546 = (inp[5]) ? 4'b0001 : 4'b0011;
																assign node26549 = (inp[5]) ? 4'b0011 : 4'b0001;
															assign node26552 = (inp[0]) ? 4'b0001 : node26553;
																assign node26553 = (inp[5]) ? 4'b0011 : 4'b0001;
												assign node26557 = (inp[4]) ? node26573 : node26558;
													assign node26558 = (inp[0]) ? node26568 : node26559;
														assign node26559 = (inp[5]) ? node26563 : node26560;
															assign node26560 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node26563 = (inp[3]) ? node26565 : 4'b0011;
																assign node26565 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node26568 = (inp[15]) ? 4'b0011 : node26569;
															assign node26569 = (inp[3]) ? 4'b0011 : 4'b0001;
													assign node26573 = (inp[15]) ? node26579 : node26574;
														assign node26574 = (inp[5]) ? node26576 : 4'b0111;
															assign node26576 = (inp[0]) ? 4'b0111 : 4'b0101;
														assign node26579 = (inp[0]) ? node26581 : 4'b0111;
															assign node26581 = (inp[3]) ? 4'b0101 : node26582;
																assign node26582 = (inp[5]) ? 4'b0101 : 4'b0111;
											assign node26586 = (inp[9]) ? node26618 : node26587;
												assign node26587 = (inp[4]) ? node26601 : node26588;
													assign node26588 = (inp[0]) ? node26596 : node26589;
														assign node26589 = (inp[15]) ? node26591 : 4'b0011;
															assign node26591 = (inp[3]) ? node26593 : 4'b0001;
																assign node26593 = (inp[5]) ? 4'b0011 : 4'b0001;
														assign node26596 = (inp[15]) ? 4'b0011 : node26597;
															assign node26597 = (inp[3]) ? 4'b0011 : 4'b0001;
													assign node26601 = (inp[5]) ? node26613 : node26602;
														assign node26602 = (inp[0]) ? node26608 : node26603;
															assign node26603 = (inp[3]) ? node26605 : 4'b0111;
																assign node26605 = (inp[15]) ? 4'b0111 : 4'b0101;
															assign node26608 = (inp[3]) ? node26610 : 4'b0101;
																assign node26610 = (inp[15]) ? 4'b0101 : 4'b0111;
														assign node26613 = (inp[0]) ? 4'b0111 : node26614;
															assign node26614 = (inp[15]) ? 4'b0111 : 4'b0101;
												assign node26618 = (inp[4]) ? node26638 : node26619;
													assign node26619 = (inp[0]) ? node26629 : node26620;
														assign node26620 = (inp[15]) ? node26626 : node26621;
															assign node26621 = (inp[5]) ? 4'b0101 : node26622;
																assign node26622 = (inp[3]) ? 4'b0101 : 4'b0111;
															assign node26626 = (inp[5]) ? 4'b0111 : 4'b0101;
														assign node26629 = (inp[3]) ? 4'b0111 : node26630;
															assign node26630 = (inp[5]) ? node26634 : node26631;
																assign node26631 = (inp[15]) ? 4'b0111 : 4'b0101;
																assign node26634 = (inp[15]) ? 4'b0101 : 4'b0111;
													assign node26638 = (inp[0]) ? node26646 : node26639;
														assign node26639 = (inp[5]) ? 4'b0001 : node26640;
															assign node26640 = (inp[15]) ? 4'b0011 : node26641;
																assign node26641 = (inp[3]) ? 4'b0001 : 4'b0011;
														assign node26646 = (inp[15]) ? 4'b0001 : node26647;
															assign node26647 = (inp[5]) ? 4'b0011 : 4'b0001;
										assign node26651 = (inp[12]) ? node26711 : node26652;
											assign node26652 = (inp[4]) ? node26682 : node26653;
												assign node26653 = (inp[9]) ? node26661 : node26654;
													assign node26654 = (inp[15]) ? node26656 : 4'b0110;
														assign node26656 = (inp[5]) ? node26658 : 4'b0100;
															assign node26658 = (inp[0]) ? 4'b0100 : 4'b0110;
													assign node26661 = (inp[5]) ? node26669 : node26662;
														assign node26662 = (inp[15]) ? node26666 : node26663;
															assign node26663 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node26666 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node26669 = (inp[15]) ? node26675 : node26670;
															assign node26670 = (inp[3]) ? 4'b0000 : node26671;
																assign node26671 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node26675 = (inp[3]) ? node26679 : node26676;
																assign node26676 = (inp[0]) ? 4'b0010 : 4'b0000;
																assign node26679 = (inp[0]) ? 4'b0000 : 4'b0010;
												assign node26682 = (inp[9]) ? node26696 : node26683;
													assign node26683 = (inp[3]) ? node26689 : node26684;
														assign node26684 = (inp[0]) ? 4'b0010 : node26685;
															assign node26685 = (inp[15]) ? 4'b0000 : 4'b0010;
														assign node26689 = (inp[5]) ? 4'b0000 : node26690;
															assign node26690 = (inp[15]) ? 4'b0010 : node26691;
																assign node26691 = (inp[0]) ? 4'b0000 : 4'b0010;
													assign node26696 = (inp[3]) ? node26704 : node26697;
														assign node26697 = (inp[15]) ? 4'b0110 : node26698;
															assign node26698 = (inp[5]) ? node26700 : 4'b0110;
																assign node26700 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node26704 = (inp[15]) ? node26708 : node26705;
															assign node26705 = (inp[0]) ? 4'b0110 : 4'b0100;
															assign node26708 = (inp[0]) ? 4'b0100 : 4'b0110;
											assign node26711 = (inp[3]) ? node26745 : node26712;
												assign node26712 = (inp[4]) ? node26726 : node26713;
													assign node26713 = (inp[9]) ? node26719 : node26714;
														assign node26714 = (inp[0]) ? 4'b0000 : node26715;
															assign node26715 = (inp[15]) ? 4'b0000 : 4'b0010;
														assign node26719 = (inp[0]) ? 4'b0100 : node26720;
															assign node26720 = (inp[15]) ? 4'b0100 : node26721;
																assign node26721 = (inp[5]) ? 4'b0100 : 4'b0110;
													assign node26726 = (inp[9]) ? node26738 : node26727;
														assign node26727 = (inp[15]) ? node26733 : node26728;
															assign node26728 = (inp[0]) ? node26730 : 4'b0100;
																assign node26730 = (inp[5]) ? 4'b0110 : 4'b0100;
															assign node26733 = (inp[0]) ? node26735 : 4'b0110;
																assign node26735 = (inp[5]) ? 4'b0100 : 4'b0110;
														assign node26738 = (inp[5]) ? 4'b0000 : node26739;
															assign node26739 = (inp[0]) ? 4'b0010 : node26740;
																assign node26740 = (inp[15]) ? 4'b0000 : 4'b0010;
												assign node26745 = (inp[9]) ? node26761 : node26746;
													assign node26746 = (inp[4]) ? node26754 : node26747;
														assign node26747 = (inp[15]) ? 4'b0000 : node26748;
															assign node26748 = (inp[5]) ? node26750 : 4'b0010;
																assign node26750 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node26754 = (inp[0]) ? node26758 : node26755;
															assign node26755 = (inp[15]) ? 4'b0110 : 4'b0100;
															assign node26758 = (inp[15]) ? 4'b0100 : 4'b0110;
													assign node26761 = (inp[4]) ? node26769 : node26762;
														assign node26762 = (inp[5]) ? node26764 : 4'b0110;
															assign node26764 = (inp[15]) ? 4'b0100 : node26765;
																assign node26765 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node26769 = (inp[5]) ? node26775 : node26770;
															assign node26770 = (inp[15]) ? node26772 : 4'b0000;
																assign node26772 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node26775 = (inp[0]) ? node26779 : node26776;
																assign node26776 = (inp[15]) ? 4'b0010 : 4'b0000;
																assign node26779 = (inp[15]) ? 4'b0000 : 4'b0010;
									assign node26782 = (inp[9]) ? node26882 : node26783;
										assign node26783 = (inp[12]) ? node26823 : node26784;
											assign node26784 = (inp[4]) ? node26808 : node26785;
												assign node26785 = (inp[15]) ? node26797 : node26786;
													assign node26786 = (inp[0]) ? node26792 : node26787;
														assign node26787 = (inp[5]) ? node26789 : 4'b0110;
															assign node26789 = (inp[3]) ? 4'b0100 : 4'b0110;
														assign node26792 = (inp[3]) ? node26794 : 4'b0100;
															assign node26794 = (inp[5]) ? 4'b0110 : 4'b0100;
													assign node26797 = (inp[0]) ? node26803 : node26798;
														assign node26798 = (inp[5]) ? node26800 : 4'b0100;
															assign node26800 = (inp[3]) ? 4'b0110 : 4'b0100;
														assign node26803 = (inp[5]) ? node26805 : 4'b0110;
															assign node26805 = (inp[3]) ? 4'b0100 : 4'b0110;
												assign node26808 = (inp[15]) ? node26816 : node26809;
													assign node26809 = (inp[0]) ? node26811 : 4'b0010;
														assign node26811 = (inp[3]) ? node26813 : 4'b0000;
															assign node26813 = (inp[5]) ? 4'b0010 : 4'b0000;
													assign node26816 = (inp[0]) ? node26818 : 4'b0000;
														assign node26818 = (inp[5]) ? node26820 : 4'b0010;
															assign node26820 = (inp[3]) ? 4'b0000 : 4'b0010;
											assign node26823 = (inp[4]) ? node26845 : node26824;
												assign node26824 = (inp[5]) ? node26832 : node26825;
													assign node26825 = (inp[0]) ? node26829 : node26826;
														assign node26826 = (inp[15]) ? 4'b0000 : 4'b0010;
														assign node26829 = (inp[15]) ? 4'b0010 : 4'b0000;
													assign node26832 = (inp[15]) ? node26840 : node26833;
														assign node26833 = (inp[0]) ? node26837 : node26834;
															assign node26834 = (inp[3]) ? 4'b0000 : 4'b0010;
															assign node26837 = (inp[3]) ? 4'b0010 : 4'b0000;
														assign node26840 = (inp[3]) ? 4'b0000 : node26841;
															assign node26841 = (inp[0]) ? 4'b0010 : 4'b0000;
												assign node26845 = (inp[3]) ? node26859 : node26846;
													assign node26846 = (inp[0]) ? node26854 : node26847;
														assign node26847 = (inp[15]) ? node26851 : node26848;
															assign node26848 = (inp[5]) ? 4'b0100 : 4'b0110;
															assign node26851 = (inp[5]) ? 4'b0110 : 4'b0100;
														assign node26854 = (inp[5]) ? 4'b0110 : node26855;
															assign node26855 = (inp[15]) ? 4'b0110 : 4'b0100;
													assign node26859 = (inp[14]) ? node26867 : node26860;
														assign node26860 = (inp[0]) ? node26864 : node26861;
															assign node26861 = (inp[15]) ? 4'b0110 : 4'b0100;
															assign node26864 = (inp[15]) ? 4'b0100 : 4'b0110;
														assign node26867 = (inp[5]) ? node26875 : node26868;
															assign node26868 = (inp[0]) ? node26872 : node26869;
																assign node26869 = (inp[15]) ? 4'b0110 : 4'b0100;
																assign node26872 = (inp[15]) ? 4'b0100 : 4'b0110;
															assign node26875 = (inp[0]) ? node26879 : node26876;
																assign node26876 = (inp[15]) ? 4'b0110 : 4'b0100;
																assign node26879 = (inp[15]) ? 4'b0100 : 4'b0110;
										assign node26882 = (inp[3]) ? node26952 : node26883;
											assign node26883 = (inp[4]) ? node26917 : node26884;
												assign node26884 = (inp[12]) ? node26906 : node26885;
													assign node26885 = (inp[14]) ? node26893 : node26886;
														assign node26886 = (inp[0]) ? node26890 : node26887;
															assign node26887 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node26890 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node26893 = (inp[5]) ? node26899 : node26894;
															assign node26894 = (inp[15]) ? node26896 : 4'b0000;
																assign node26896 = (inp[0]) ? 4'b0010 : 4'b0000;
															assign node26899 = (inp[0]) ? node26903 : node26900;
																assign node26900 = (inp[15]) ? 4'b0000 : 4'b0010;
																assign node26903 = (inp[15]) ? 4'b0010 : 4'b0000;
													assign node26906 = (inp[14]) ? 4'b0110 : node26907;
														assign node26907 = (inp[0]) ? 4'b0100 : node26908;
															assign node26908 = (inp[5]) ? node26912 : node26909;
																assign node26909 = (inp[15]) ? 4'b0100 : 4'b0110;
																assign node26912 = (inp[15]) ? 4'b0110 : 4'b0100;
												assign node26917 = (inp[12]) ? node26931 : node26918;
													assign node26918 = (inp[0]) ? node26924 : node26919;
														assign node26919 = (inp[5]) ? node26921 : 4'b0110;
															assign node26921 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node26924 = (inp[15]) ? node26928 : node26925;
															assign node26925 = (inp[5]) ? 4'b0110 : 4'b0100;
															assign node26928 = (inp[5]) ? 4'b0100 : 4'b0110;
													assign node26931 = (inp[0]) ? node26947 : node26932;
														assign node26932 = (inp[14]) ? node26940 : node26933;
															assign node26933 = (inp[15]) ? node26937 : node26934;
																assign node26934 = (inp[5]) ? 4'b0000 : 4'b0010;
																assign node26937 = (inp[5]) ? 4'b0010 : 4'b0000;
															assign node26940 = (inp[15]) ? node26944 : node26941;
																assign node26941 = (inp[5]) ? 4'b0000 : 4'b0010;
																assign node26944 = (inp[5]) ? 4'b0010 : 4'b0000;
														assign node26947 = (inp[5]) ? node26949 : 4'b0000;
															assign node26949 = (inp[15]) ? 4'b0000 : 4'b0010;
											assign node26952 = (inp[5]) ? node26980 : node26953;
												assign node26953 = (inp[4]) ? node26967 : node26954;
													assign node26954 = (inp[12]) ? node26960 : node26955;
														assign node26955 = (inp[15]) ? node26957 : 4'b0010;
															assign node26957 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node26960 = (inp[0]) ? node26964 : node26961;
															assign node26961 = (inp[15]) ? 4'b0110 : 4'b0100;
															assign node26964 = (inp[15]) ? 4'b0100 : 4'b0110;
													assign node26967 = (inp[12]) ? node26973 : node26968;
														assign node26968 = (inp[15]) ? node26970 : 4'b0100;
															assign node26970 = (inp[0]) ? 4'b0100 : 4'b0110;
														assign node26973 = (inp[15]) ? node26977 : node26974;
															assign node26974 = (inp[0]) ? 4'b0010 : 4'b0000;
															assign node26977 = (inp[0]) ? 4'b0000 : 4'b0010;
												assign node26980 = (inp[0]) ? node27000 : node26981;
													assign node26981 = (inp[15]) ? node26997 : node26982;
														assign node26982 = (inp[14]) ? node26990 : node26983;
															assign node26983 = (inp[4]) ? node26987 : node26984;
																assign node26984 = (inp[12]) ? 4'b0100 : 4'b0000;
																assign node26987 = (inp[12]) ? 4'b0000 : 4'b0100;
															assign node26990 = (inp[12]) ? node26994 : node26991;
																assign node26991 = (inp[4]) ? 4'b0100 : 4'b0000;
																assign node26994 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node26997 = (inp[14]) ? 4'b0110 : 4'b0010;
													assign node27000 = (inp[15]) ? node27008 : node27001;
														assign node27001 = (inp[12]) ? node27005 : node27002;
															assign node27002 = (inp[4]) ? 4'b0110 : 4'b0010;
															assign node27005 = (inp[4]) ? 4'b0010 : 4'b0110;
														assign node27008 = (inp[4]) ? node27012 : node27009;
															assign node27009 = (inp[12]) ? 4'b0100 : 4'b0000;
															assign node27012 = (inp[12]) ? 4'b0000 : 4'b0100;
					assign node27015 = (inp[13]) ? node29131 : node27016;
						assign node27016 = (inp[8]) ? node28050 : node27017;
							assign node27017 = (inp[7]) ? node27517 : node27018;
								assign node27018 = (inp[14]) ? node27278 : node27019;
									assign node27019 = (inp[2]) ? node27151 : node27020;
										assign node27020 = (inp[4]) ? node27082 : node27021;
											assign node27021 = (inp[5]) ? node27053 : node27022;
												assign node27022 = (inp[15]) ? node27038 : node27023;
													assign node27023 = (inp[0]) ? node27031 : node27024;
														assign node27024 = (inp[9]) ? node27026 : 4'b1011;
															assign node27026 = (inp[12]) ? node27028 : 4'b1011;
																assign node27028 = (inp[3]) ? 4'b1101 : 4'b1111;
														assign node27031 = (inp[9]) ? node27035 : node27032;
															assign node27032 = (inp[12]) ? 4'b1001 : 4'b1101;
															assign node27035 = (inp[12]) ? 4'b1111 : 4'b1001;
													assign node27038 = (inp[0]) ? node27046 : node27039;
														assign node27039 = (inp[12]) ? node27043 : node27040;
															assign node27040 = (inp[9]) ? 4'b1001 : 4'b1101;
															assign node27043 = (inp[9]) ? 4'b1111 : 4'b1001;
														assign node27046 = (inp[9]) ? node27050 : node27047;
															assign node27047 = (inp[12]) ? 4'b1011 : 4'b1111;
															assign node27050 = (inp[12]) ? 4'b1101 : 4'b1011;
												assign node27053 = (inp[15]) ? node27065 : node27054;
													assign node27054 = (inp[9]) ? node27060 : node27055;
														assign node27055 = (inp[3]) ? 4'b1101 : node27056;
															assign node27056 = (inp[0]) ? 4'b1101 : 4'b1111;
														assign node27060 = (inp[12]) ? node27062 : 4'b1011;
															assign node27062 = (inp[0]) ? 4'b1111 : 4'b1101;
													assign node27065 = (inp[9]) ? node27075 : node27066;
														assign node27066 = (inp[12]) ? node27068 : 4'b1101;
															assign node27068 = (inp[0]) ? node27072 : node27069;
																assign node27069 = (inp[3]) ? 4'b1011 : 4'b1001;
																assign node27072 = (inp[3]) ? 4'b1001 : 4'b1011;
														assign node27075 = (inp[12]) ? node27079 : node27076;
															assign node27076 = (inp[3]) ? 4'b1001 : 4'b1011;
															assign node27079 = (inp[0]) ? 4'b1101 : 4'b1111;
											assign node27082 = (inp[15]) ? node27116 : node27083;
												assign node27083 = (inp[5]) ? node27103 : node27084;
													assign node27084 = (inp[12]) ? node27096 : node27085;
														assign node27085 = (inp[9]) ? node27089 : node27086;
															assign node27086 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node27089 = (inp[3]) ? node27093 : node27090;
																assign node27090 = (inp[0]) ? 4'b1101 : 4'b1111;
																assign node27093 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node27096 = (inp[9]) ? node27098 : 4'b1101;
															assign node27098 = (inp[0]) ? 4'b1001 : node27099;
																assign node27099 = (inp[3]) ? 4'b1001 : 4'b1011;
													assign node27103 = (inp[0]) ? node27111 : node27104;
														assign node27104 = (inp[9]) ? node27108 : node27105;
															assign node27105 = (inp[12]) ? 4'b1101 : 4'b1001;
															assign node27108 = (inp[12]) ? 4'b1001 : 4'b1101;
														assign node27111 = (inp[3]) ? node27113 : 4'b1001;
															assign node27113 = (inp[9]) ? 4'b1011 : 4'b1111;
												assign node27116 = (inp[0]) ? node27136 : node27117;
													assign node27117 = (inp[3]) ? node27131 : node27118;
														assign node27118 = (inp[5]) ? node27126 : node27119;
															assign node27119 = (inp[9]) ? node27123 : node27120;
																assign node27120 = (inp[12]) ? 4'b1101 : 4'b1001;
																assign node27123 = (inp[12]) ? 4'b1001 : 4'b1101;
															assign node27126 = (inp[12]) ? 4'b1111 : node27127;
																assign node27127 = (inp[9]) ? 4'b1111 : 4'b1001;
														assign node27131 = (inp[9]) ? 4'b1011 : node27132;
															assign node27132 = (inp[12]) ? 4'b1111 : 4'b1011;
													assign node27136 = (inp[5]) ? node27144 : node27137;
														assign node27137 = (inp[9]) ? node27141 : node27138;
															assign node27138 = (inp[3]) ? 4'b1011 : 4'b1111;
															assign node27141 = (inp[3]) ? 4'b1101 : 4'b1111;
														assign node27144 = (inp[9]) ? node27148 : node27145;
															assign node27145 = (inp[12]) ? 4'b1101 : 4'b1001;
															assign node27148 = (inp[12]) ? 4'b1001 : 4'b1101;
										assign node27151 = (inp[4]) ? node27225 : node27152;
											assign node27152 = (inp[5]) ? node27194 : node27153;
												assign node27153 = (inp[3]) ? node27175 : node27154;
													assign node27154 = (inp[9]) ? node27166 : node27155;
														assign node27155 = (inp[12]) ? node27161 : node27156;
															assign node27156 = (inp[15]) ? 4'b1100 : node27157;
																assign node27157 = (inp[0]) ? 4'b1100 : 4'b1110;
															assign node27161 = (inp[0]) ? 4'b1010 : node27162;
																assign node27162 = (inp[15]) ? 4'b1000 : 4'b1010;
														assign node27166 = (inp[12]) ? node27168 : 4'b1010;
															assign node27168 = (inp[15]) ? node27172 : node27169;
																assign node27169 = (inp[0]) ? 4'b1100 : 4'b1110;
																assign node27172 = (inp[0]) ? 4'b1110 : 4'b1100;
													assign node27175 = (inp[15]) ? node27183 : node27176;
														assign node27176 = (inp[0]) ? node27178 : 4'b1100;
															assign node27178 = (inp[12]) ? 4'b1000 : node27179;
																assign node27179 = (inp[9]) ? 4'b1000 : 4'b1100;
														assign node27183 = (inp[9]) ? node27189 : node27184;
															assign node27184 = (inp[12]) ? 4'b1010 : node27185;
																assign node27185 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node27189 = (inp[12]) ? node27191 : 4'b1000;
																assign node27191 = (inp[0]) ? 4'b1100 : 4'b1110;
												assign node27194 = (inp[9]) ? node27210 : node27195;
													assign node27195 = (inp[12]) ? node27205 : node27196;
														assign node27196 = (inp[0]) ? node27198 : 4'b1100;
															assign node27198 = (inp[15]) ? node27202 : node27199;
																assign node27199 = (inp[3]) ? 4'b1110 : 4'b1100;
																assign node27202 = (inp[3]) ? 4'b1100 : 4'b1110;
														assign node27205 = (inp[0]) ? node27207 : 4'b1010;
															assign node27207 = (inp[15]) ? 4'b1010 : 4'b1000;
													assign node27210 = (inp[12]) ? node27212 : 4'b1010;
														assign node27212 = (inp[3]) ? node27220 : node27213;
															assign node27213 = (inp[0]) ? node27217 : node27214;
																assign node27214 = (inp[15]) ? 4'b1110 : 4'b1100;
																assign node27217 = (inp[15]) ? 4'b1100 : 4'b1110;
															assign node27220 = (inp[15]) ? 4'b1110 : node27221;
																assign node27221 = (inp[0]) ? 4'b1110 : 4'b1100;
											assign node27225 = (inp[15]) ? node27257 : node27226;
												assign node27226 = (inp[0]) ? node27240 : node27227;
													assign node27227 = (inp[5]) ? node27235 : node27228;
														assign node27228 = (inp[12]) ? node27232 : node27229;
															assign node27229 = (inp[9]) ? 4'b1110 : 4'b1010;
															assign node27232 = (inp[3]) ? 4'b1000 : 4'b1010;
														assign node27235 = (inp[12]) ? 4'b1000 : node27236;
															assign node27236 = (inp[3]) ? 4'b1000 : 4'b1010;
													assign node27240 = (inp[3]) ? node27250 : node27241;
														assign node27241 = (inp[5]) ? 4'b1110 : node27242;
															assign node27242 = (inp[12]) ? node27246 : node27243;
																assign node27243 = (inp[9]) ? 4'b1100 : 4'b1000;
																assign node27246 = (inp[9]) ? 4'b1000 : 4'b1100;
														assign node27250 = (inp[5]) ? node27252 : 4'b1110;
															assign node27252 = (inp[9]) ? node27254 : 4'b1010;
																assign node27254 = (inp[12]) ? 4'b1010 : 4'b1110;
												assign node27257 = (inp[9]) ? node27271 : node27258;
													assign node27258 = (inp[12]) ? node27262 : node27259;
														assign node27259 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node27262 = (inp[5]) ? 4'b1100 : node27263;
															assign node27263 = (inp[0]) ? node27267 : node27264;
																assign node27264 = (inp[3]) ? 4'b1110 : 4'b1100;
																assign node27267 = (inp[3]) ? 4'b1100 : 4'b1110;
													assign node27271 = (inp[12]) ? 4'b1000 : node27272;
														assign node27272 = (inp[5]) ? node27274 : 4'b1100;
															assign node27274 = (inp[3]) ? 4'b1100 : 4'b1110;
									assign node27278 = (inp[15]) ? node27390 : node27279;
										assign node27279 = (inp[12]) ? node27317 : node27280;
											assign node27280 = (inp[9]) ? node27298 : node27281;
												assign node27281 = (inp[4]) ? node27291 : node27282;
													assign node27282 = (inp[0]) ? node27288 : node27283;
														assign node27283 = (inp[3]) ? node27285 : 4'b1110;
															assign node27285 = (inp[5]) ? 4'b1100 : 4'b1110;
														assign node27288 = (inp[5]) ? 4'b1110 : 4'b1100;
													assign node27291 = (inp[3]) ? node27293 : 4'b1010;
														assign node27293 = (inp[0]) ? node27295 : 4'b1000;
															assign node27295 = (inp[5]) ? 4'b1010 : 4'b1000;
												assign node27298 = (inp[4]) ? node27308 : node27299;
													assign node27299 = (inp[0]) ? node27303 : node27300;
														assign node27300 = (inp[5]) ? 4'b1000 : 4'b1010;
														assign node27303 = (inp[5]) ? node27305 : 4'b1000;
															assign node27305 = (inp[3]) ? 4'b1010 : 4'b1000;
													assign node27308 = (inp[0]) ? node27314 : node27309;
														assign node27309 = (inp[5]) ? 4'b1100 : node27310;
															assign node27310 = (inp[3]) ? 4'b1100 : 4'b1110;
														assign node27314 = (inp[2]) ? 4'b1110 : 4'b1100;
											assign node27317 = (inp[0]) ? node27355 : node27318;
												assign node27318 = (inp[3]) ? node27334 : node27319;
													assign node27319 = (inp[5]) ? node27329 : node27320;
														assign node27320 = (inp[2]) ? node27324 : node27321;
															assign node27321 = (inp[4]) ? 4'b1010 : 4'b1110;
															assign node27324 = (inp[9]) ? 4'b1010 : node27325;
																assign node27325 = (inp[4]) ? 4'b1110 : 4'b1010;
														assign node27329 = (inp[9]) ? node27331 : 4'b1010;
															assign node27331 = (inp[4]) ? 4'b1000 : 4'b1100;
													assign node27334 = (inp[5]) ? node27342 : node27335;
														assign node27335 = (inp[9]) ? node27339 : node27336;
															assign node27336 = (inp[4]) ? 4'b1100 : 4'b1010;
															assign node27339 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node27342 = (inp[2]) ? node27350 : node27343;
															assign node27343 = (inp[9]) ? node27347 : node27344;
																assign node27344 = (inp[4]) ? 4'b1100 : 4'b1000;
																assign node27347 = (inp[4]) ? 4'b1000 : 4'b1100;
															assign node27350 = (inp[9]) ? 4'b1100 : node27351;
																assign node27351 = (inp[4]) ? 4'b1100 : 4'b1000;
												assign node27355 = (inp[3]) ? node27373 : node27356;
													assign node27356 = (inp[5]) ? node27368 : node27357;
														assign node27357 = (inp[2]) ? node27363 : node27358;
															assign node27358 = (inp[9]) ? node27360 : 4'b1100;
																assign node27360 = (inp[4]) ? 4'b1000 : 4'b1100;
															assign node27363 = (inp[4]) ? node27365 : 4'b1000;
																assign node27365 = (inp[9]) ? 4'b1000 : 4'b1100;
														assign node27368 = (inp[9]) ? node27370 : 4'b1000;
															assign node27370 = (inp[4]) ? 4'b1010 : 4'b1110;
													assign node27373 = (inp[5]) ? node27383 : node27374;
														assign node27374 = (inp[2]) ? node27378 : node27375;
															assign node27375 = (inp[9]) ? 4'b1010 : 4'b1000;
															assign node27378 = (inp[4]) ? node27380 : 4'b1110;
																assign node27380 = (inp[9]) ? 4'b1010 : 4'b1110;
														assign node27383 = (inp[9]) ? node27387 : node27384;
															assign node27384 = (inp[4]) ? 4'b1110 : 4'b1010;
															assign node27387 = (inp[4]) ? 4'b1010 : 4'b1110;
										assign node27390 = (inp[5]) ? node27448 : node27391;
											assign node27391 = (inp[0]) ? node27415 : node27392;
												assign node27392 = (inp[9]) ? node27400 : node27393;
													assign node27393 = (inp[4]) ? node27397 : node27394;
														assign node27394 = (inp[12]) ? 4'b1000 : 4'b1100;
														assign node27397 = (inp[12]) ? 4'b1100 : 4'b1000;
													assign node27400 = (inp[3]) ? node27408 : node27401;
														assign node27401 = (inp[2]) ? node27403 : 4'b1100;
															assign node27403 = (inp[4]) ? 4'b1000 : node27404;
																assign node27404 = (inp[12]) ? 4'b1100 : 4'b1000;
														assign node27408 = (inp[12]) ? node27412 : node27409;
															assign node27409 = (inp[4]) ? 4'b1110 : 4'b1000;
															assign node27412 = (inp[4]) ? 4'b1010 : 4'b1110;
												assign node27415 = (inp[3]) ? node27431 : node27416;
													assign node27416 = (inp[4]) ? node27424 : node27417;
														assign node27417 = (inp[12]) ? node27421 : node27418;
															assign node27418 = (inp[9]) ? 4'b1010 : 4'b1110;
															assign node27421 = (inp[9]) ? 4'b1110 : 4'b1010;
														assign node27424 = (inp[12]) ? node27428 : node27425;
															assign node27425 = (inp[2]) ? 4'b1010 : 4'b1110;
															assign node27428 = (inp[9]) ? 4'b1010 : 4'b1110;
													assign node27431 = (inp[9]) ? node27441 : node27432;
														assign node27432 = (inp[2]) ? node27438 : node27433;
															assign node27433 = (inp[12]) ? 4'b1010 : node27434;
																assign node27434 = (inp[4]) ? 4'b1010 : 4'b1110;
															assign node27438 = (inp[12]) ? 4'b1100 : 4'b1110;
														assign node27441 = (inp[4]) ? node27445 : node27442;
															assign node27442 = (inp[12]) ? 4'b1100 : 4'b1010;
															assign node27445 = (inp[12]) ? 4'b1000 : 4'b1100;
											assign node27448 = (inp[0]) ? node27484 : node27449;
												assign node27449 = (inp[3]) ? node27463 : node27450;
													assign node27450 = (inp[12]) ? node27458 : node27451;
														assign node27451 = (inp[4]) ? node27455 : node27452;
															assign node27452 = (inp[9]) ? 4'b1000 : 4'b1100;
															assign node27455 = (inp[9]) ? 4'b1110 : 4'b1000;
														assign node27458 = (inp[4]) ? 4'b1110 : node27459;
															assign node27459 = (inp[9]) ? 4'b1110 : 4'b1000;
													assign node27463 = (inp[9]) ? node27477 : node27464;
														assign node27464 = (inp[2]) ? node27470 : node27465;
															assign node27465 = (inp[12]) ? 4'b1110 : node27466;
																assign node27466 = (inp[4]) ? 4'b1010 : 4'b1110;
															assign node27470 = (inp[4]) ? node27474 : node27471;
																assign node27471 = (inp[12]) ? 4'b1010 : 4'b1110;
																assign node27474 = (inp[12]) ? 4'b1110 : 4'b1010;
														assign node27477 = (inp[12]) ? node27481 : node27478;
															assign node27478 = (inp[4]) ? 4'b1110 : 4'b1010;
															assign node27481 = (inp[4]) ? 4'b1010 : 4'b1110;
												assign node27484 = (inp[3]) ? node27502 : node27485;
													assign node27485 = (inp[4]) ? node27495 : node27486;
														assign node27486 = (inp[2]) ? node27488 : 4'b1010;
															assign node27488 = (inp[9]) ? node27492 : node27489;
																assign node27489 = (inp[12]) ? 4'b1010 : 4'b1110;
																assign node27492 = (inp[12]) ? 4'b1100 : 4'b1010;
														assign node27495 = (inp[12]) ? node27499 : node27496;
															assign node27496 = (inp[9]) ? 4'b1100 : 4'b1010;
															assign node27499 = (inp[9]) ? 4'b1000 : 4'b1100;
													assign node27502 = (inp[12]) ? node27510 : node27503;
														assign node27503 = (inp[4]) ? node27507 : node27504;
															assign node27504 = (inp[9]) ? 4'b1000 : 4'b1100;
															assign node27507 = (inp[9]) ? 4'b1100 : 4'b1000;
														assign node27510 = (inp[9]) ? node27514 : node27511;
															assign node27511 = (inp[4]) ? 4'b1100 : 4'b1000;
															assign node27514 = (inp[4]) ? 4'b1000 : 4'b1100;
								assign node27517 = (inp[2]) ? node27777 : node27518;
									assign node27518 = (inp[14]) ? node27644 : node27519;
										assign node27519 = (inp[4]) ? node27581 : node27520;
											assign node27520 = (inp[9]) ? node27552 : node27521;
												assign node27521 = (inp[12]) ? node27531 : node27522;
													assign node27522 = (inp[3]) ? node27524 : 4'b1110;
														assign node27524 = (inp[5]) ? node27526 : 4'b1110;
															assign node27526 = (inp[0]) ? 4'b1100 : node27527;
																assign node27527 = (inp[15]) ? 4'b1110 : 4'b1100;
													assign node27531 = (inp[5]) ? node27539 : node27532;
														assign node27532 = (inp[3]) ? node27534 : 4'b1010;
															assign node27534 = (inp[15]) ? 4'b1010 : node27535;
																assign node27535 = (inp[0]) ? 4'b1000 : 4'b1010;
														assign node27539 = (inp[3]) ? node27547 : node27540;
															assign node27540 = (inp[0]) ? node27544 : node27541;
																assign node27541 = (inp[15]) ? 4'b1000 : 4'b1010;
																assign node27544 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node27547 = (inp[15]) ? 4'b1010 : node27548;
																assign node27548 = (inp[0]) ? 4'b1010 : 4'b1000;
												assign node27552 = (inp[12]) ? node27566 : node27553;
													assign node27553 = (inp[15]) ? node27559 : node27554;
														assign node27554 = (inp[0]) ? node27556 : 4'b1010;
															assign node27556 = (inp[5]) ? 4'b1010 : 4'b1000;
														assign node27559 = (inp[0]) ? 4'b1010 : node27560;
															assign node27560 = (inp[5]) ? node27562 : 4'b1000;
																assign node27562 = (inp[3]) ? 4'b1010 : 4'b1000;
													assign node27566 = (inp[15]) ? node27578 : node27567;
														assign node27567 = (inp[0]) ? node27573 : node27568;
															assign node27568 = (inp[3]) ? 4'b1100 : node27569;
																assign node27569 = (inp[5]) ? 4'b1100 : 4'b1110;
															assign node27573 = (inp[3]) ? 4'b1110 : node27574;
																assign node27574 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node27578 = (inp[0]) ? 4'b1100 : 4'b1110;
											assign node27581 = (inp[15]) ? node27609 : node27582;
												assign node27582 = (inp[0]) ? node27598 : node27583;
													assign node27583 = (inp[5]) ? node27593 : node27584;
														assign node27584 = (inp[3]) ? node27588 : node27585;
															assign node27585 = (inp[9]) ? 4'b1010 : 4'b1110;
															assign node27588 = (inp[9]) ? node27590 : 4'b1010;
																assign node27590 = (inp[12]) ? 4'b1000 : 4'b1100;
														assign node27593 = (inp[12]) ? 4'b1100 : node27594;
															assign node27594 = (inp[9]) ? 4'b1100 : 4'b1000;
													assign node27598 = (inp[5]) ? 4'b1110 : node27599;
														assign node27599 = (inp[3]) ? node27603 : node27600;
															assign node27600 = (inp[12]) ? 4'b1000 : 4'b1100;
															assign node27603 = (inp[9]) ? 4'b1110 : node27604;
																assign node27604 = (inp[12]) ? 4'b1110 : 4'b1000;
												assign node27609 = (inp[0]) ? node27625 : node27610;
													assign node27610 = (inp[3]) ? node27616 : node27611;
														assign node27611 = (inp[9]) ? 4'b1000 : node27612;
															assign node27612 = (inp[12]) ? 4'b1100 : 4'b1000;
														assign node27616 = (inp[9]) ? node27622 : node27617;
															assign node27617 = (inp[5]) ? node27619 : 4'b1000;
																assign node27619 = (inp[12]) ? 4'b1110 : 4'b1010;
															assign node27622 = (inp[12]) ? 4'b1010 : 4'b1110;
													assign node27625 = (inp[3]) ? node27637 : node27626;
														assign node27626 = (inp[5]) ? node27630 : node27627;
															assign node27627 = (inp[12]) ? 4'b1010 : 4'b1110;
															assign node27630 = (inp[12]) ? node27634 : node27631;
																assign node27631 = (inp[9]) ? 4'b1100 : 4'b1010;
																assign node27634 = (inp[9]) ? 4'b1000 : 4'b1100;
														assign node27637 = (inp[9]) ? node27641 : node27638;
															assign node27638 = (inp[12]) ? 4'b1100 : 4'b1000;
															assign node27641 = (inp[12]) ? 4'b1000 : 4'b1100;
										assign node27644 = (inp[5]) ? node27718 : node27645;
											assign node27645 = (inp[9]) ? node27681 : node27646;
												assign node27646 = (inp[12]) ? node27658 : node27647;
													assign node27647 = (inp[4]) ? node27653 : node27648;
														assign node27648 = (inp[0]) ? node27650 : 4'b0111;
															assign node27650 = (inp[15]) ? 4'b0111 : 4'b0101;
														assign node27653 = (inp[0]) ? 4'b0011 : node27654;
															assign node27654 = (inp[15]) ? 4'b0001 : 4'b0011;
													assign node27658 = (inp[4]) ? node27674 : node27659;
														assign node27659 = (inp[3]) ? node27667 : node27660;
															assign node27660 = (inp[0]) ? node27664 : node27661;
																assign node27661 = (inp[15]) ? 4'b0001 : 4'b0011;
																assign node27664 = (inp[15]) ? 4'b0011 : 4'b0001;
															assign node27667 = (inp[15]) ? node27671 : node27668;
																assign node27668 = (inp[0]) ? 4'b0001 : 4'b0011;
																assign node27671 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node27674 = (inp[3]) ? node27676 : 4'b0101;
															assign node27676 = (inp[0]) ? 4'b0111 : node27677;
																assign node27677 = (inp[15]) ? 4'b0111 : 4'b0101;
												assign node27681 = (inp[15]) ? node27697 : node27682;
													assign node27682 = (inp[3]) ? node27688 : node27683;
														assign node27683 = (inp[4]) ? 4'b0001 : node27684;
															assign node27684 = (inp[12]) ? 4'b0101 : 4'b0001;
														assign node27688 = (inp[4]) ? node27692 : node27689;
															assign node27689 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node27692 = (inp[0]) ? 4'b0011 : node27693;
																assign node27693 = (inp[12]) ? 4'b0001 : 4'b0101;
													assign node27697 = (inp[3]) ? node27707 : node27698;
														assign node27698 = (inp[0]) ? node27700 : 4'b0001;
															assign node27700 = (inp[12]) ? node27704 : node27701;
																assign node27701 = (inp[4]) ? 4'b0111 : 4'b0011;
																assign node27704 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node27707 = (inp[0]) ? node27713 : node27708;
															assign node27708 = (inp[12]) ? 4'b0111 : node27709;
																assign node27709 = (inp[4]) ? 4'b0111 : 4'b0001;
															assign node27713 = (inp[12]) ? node27715 : 4'b0101;
																assign node27715 = (inp[4]) ? 4'b0001 : 4'b0101;
											assign node27718 = (inp[4]) ? node27746 : node27719;
												assign node27719 = (inp[12]) ? node27731 : node27720;
													assign node27720 = (inp[9]) ? 4'b0011 : node27721;
														assign node27721 = (inp[15]) ? node27723 : 4'b0111;
															assign node27723 = (inp[3]) ? node27727 : node27724;
																assign node27724 = (inp[0]) ? 4'b0111 : 4'b0101;
																assign node27727 = (inp[0]) ? 4'b0101 : 4'b0111;
													assign node27731 = (inp[9]) ? node27739 : node27732;
														assign node27732 = (inp[0]) ? 4'b0011 : node27733;
															assign node27733 = (inp[3]) ? node27735 : 4'b0011;
																assign node27735 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node27739 = (inp[0]) ? node27743 : node27740;
															assign node27740 = (inp[15]) ? 4'b0111 : 4'b0101;
															assign node27743 = (inp[15]) ? 4'b0101 : 4'b0111;
												assign node27746 = (inp[3]) ? node27760 : node27747;
													assign node27747 = (inp[0]) ? node27757 : node27748;
														assign node27748 = (inp[15]) ? node27754 : node27749;
															assign node27749 = (inp[12]) ? node27751 : 4'b0101;
																assign node27751 = (inp[9]) ? 4'b0001 : 4'b0101;
															assign node27754 = (inp[12]) ? 4'b0111 : 4'b0001;
														assign node27757 = (inp[15]) ? 4'b0101 : 4'b0111;
													assign node27760 = (inp[15]) ? node27766 : node27761;
														assign node27761 = (inp[0]) ? node27763 : 4'b0101;
															assign node27763 = (inp[9]) ? 4'b0011 : 4'b0111;
														assign node27766 = (inp[0]) ? node27772 : node27767;
															assign node27767 = (inp[9]) ? node27769 : 4'b0011;
																assign node27769 = (inp[12]) ? 4'b0011 : 4'b0111;
															assign node27772 = (inp[12]) ? 4'b0101 : node27773;
																assign node27773 = (inp[9]) ? 4'b0101 : 4'b0001;
									assign node27777 = (inp[15]) ? node27899 : node27778;
										assign node27778 = (inp[12]) ? node27832 : node27779;
											assign node27779 = (inp[0]) ? node27811 : node27780;
												assign node27780 = (inp[5]) ? node27788 : node27781;
													assign node27781 = (inp[9]) ? node27785 : node27782;
														assign node27782 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node27785 = (inp[4]) ? 4'b0101 : 4'b0011;
													assign node27788 = (inp[3]) ? node27796 : node27789;
														assign node27789 = (inp[4]) ? node27793 : node27790;
															assign node27790 = (inp[14]) ? 4'b0111 : 4'b0011;
															assign node27793 = (inp[9]) ? 4'b0101 : 4'b0011;
														assign node27796 = (inp[14]) ? node27804 : node27797;
															assign node27797 = (inp[9]) ? node27801 : node27798;
																assign node27798 = (inp[4]) ? 4'b0001 : 4'b0101;
																assign node27801 = (inp[4]) ? 4'b0101 : 4'b0001;
															assign node27804 = (inp[4]) ? node27808 : node27805;
																assign node27805 = (inp[9]) ? 4'b0001 : 4'b0101;
																assign node27808 = (inp[9]) ? 4'b0101 : 4'b0001;
												assign node27811 = (inp[5]) ? node27821 : node27812;
													assign node27812 = (inp[4]) ? node27816 : node27813;
														assign node27813 = (inp[9]) ? 4'b0001 : 4'b0101;
														assign node27816 = (inp[9]) ? node27818 : 4'b0001;
															assign node27818 = (inp[3]) ? 4'b0111 : 4'b0101;
													assign node27821 = (inp[3]) ? node27827 : node27822;
														assign node27822 = (inp[4]) ? node27824 : 4'b0001;
															assign node27824 = (inp[9]) ? 4'b0111 : 4'b0001;
														assign node27827 = (inp[4]) ? node27829 : 4'b0011;
															assign node27829 = (inp[9]) ? 4'b0111 : 4'b0011;
											assign node27832 = (inp[0]) ? node27872 : node27833;
												assign node27833 = (inp[5]) ? node27849 : node27834;
													assign node27834 = (inp[3]) ? node27842 : node27835;
														assign node27835 = (inp[4]) ? node27839 : node27836;
															assign node27836 = (inp[9]) ? 4'b0111 : 4'b0011;
															assign node27839 = (inp[9]) ? 4'b0011 : 4'b0111;
														assign node27842 = (inp[9]) ? node27846 : node27843;
															assign node27843 = (inp[4]) ? 4'b0101 : 4'b0011;
															assign node27846 = (inp[14]) ? 4'b0001 : 4'b0101;
													assign node27849 = (inp[14]) ? node27861 : node27850;
														assign node27850 = (inp[3]) ? node27856 : node27851;
															assign node27851 = (inp[9]) ? node27853 : 4'b0101;
																assign node27853 = (inp[4]) ? 4'b0001 : 4'b0101;
															assign node27856 = (inp[4]) ? 4'b0001 : node27857;
																assign node27857 = (inp[9]) ? 4'b0101 : 4'b0001;
														assign node27861 = (inp[3]) ? node27865 : node27862;
															assign node27862 = (inp[9]) ? 4'b0001 : 4'b0011;
															assign node27865 = (inp[4]) ? node27869 : node27866;
																assign node27866 = (inp[9]) ? 4'b0101 : 4'b0001;
																assign node27869 = (inp[9]) ? 4'b0001 : 4'b0101;
												assign node27872 = (inp[5]) ? node27882 : node27873;
													assign node27873 = (inp[3]) ? node27879 : node27874;
														assign node27874 = (inp[4]) ? node27876 : 4'b0001;
															assign node27876 = (inp[9]) ? 4'b0001 : 4'b0101;
														assign node27879 = (inp[4]) ? 4'b0011 : 4'b0001;
													assign node27882 = (inp[14]) ? node27892 : node27883;
														assign node27883 = (inp[3]) ? node27885 : 4'b0111;
															assign node27885 = (inp[9]) ? node27889 : node27886;
																assign node27886 = (inp[4]) ? 4'b0111 : 4'b0011;
																assign node27889 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node27892 = (inp[9]) ? node27896 : node27893;
															assign node27893 = (inp[4]) ? 4'b0111 : 4'b0001;
															assign node27896 = (inp[4]) ? 4'b0011 : 4'b0111;
										assign node27899 = (inp[14]) ? node27963 : node27900;
											assign node27900 = (inp[0]) ? node27934 : node27901;
												assign node27901 = (inp[3]) ? node27919 : node27902;
													assign node27902 = (inp[5]) ? node27912 : node27903;
														assign node27903 = (inp[4]) ? node27905 : 4'b0001;
															assign node27905 = (inp[9]) ? node27909 : node27906;
																assign node27906 = (inp[12]) ? 4'b0101 : 4'b0001;
																assign node27909 = (inp[12]) ? 4'b0001 : 4'b0101;
														assign node27912 = (inp[12]) ? 4'b0111 : node27913;
															assign node27913 = (inp[9]) ? node27915 : 4'b0001;
																assign node27915 = (inp[4]) ? 4'b0111 : 4'b0001;
													assign node27919 = (inp[4]) ? 4'b0111 : node27920;
														assign node27920 = (inp[5]) ? node27926 : node27921;
															assign node27921 = (inp[9]) ? 4'b0111 : node27922;
																assign node27922 = (inp[12]) ? 4'b0001 : 4'b0101;
															assign node27926 = (inp[9]) ? node27930 : node27927;
																assign node27927 = (inp[12]) ? 4'b0011 : 4'b0111;
																assign node27930 = (inp[12]) ? 4'b0111 : 4'b0011;
												assign node27934 = (inp[3]) ? node27950 : node27935;
													assign node27935 = (inp[9]) ? node27941 : node27936;
														assign node27936 = (inp[5]) ? node27938 : 4'b0111;
															assign node27938 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node27941 = (inp[5]) ? 4'b0011 : node27942;
															assign node27942 = (inp[4]) ? node27946 : node27943;
																assign node27943 = (inp[12]) ? 4'b0111 : 4'b0011;
																assign node27946 = (inp[12]) ? 4'b0011 : 4'b0111;
													assign node27950 = (inp[12]) ? node27958 : node27951;
														assign node27951 = (inp[5]) ? 4'b0101 : node27952;
															assign node27952 = (inp[4]) ? 4'b0011 : node27953;
																assign node27953 = (inp[9]) ? 4'b0011 : 4'b0111;
														assign node27958 = (inp[5]) ? 4'b0001 : node27959;
															assign node27959 = (inp[4]) ? 4'b0001 : 4'b0101;
											assign node27963 = (inp[5]) ? node28009 : node27964;
												assign node27964 = (inp[0]) ? node27986 : node27965;
													assign node27965 = (inp[3]) ? node27975 : node27966;
														assign node27966 = (inp[9]) ? 4'b0001 : node27967;
															assign node27967 = (inp[12]) ? node27971 : node27968;
																assign node27968 = (inp[4]) ? 4'b0001 : 4'b0101;
																assign node27971 = (inp[4]) ? 4'b0101 : 4'b0001;
														assign node27975 = (inp[12]) ? node27981 : node27976;
															assign node27976 = (inp[4]) ? 4'b0111 : node27977;
																assign node27977 = (inp[9]) ? 4'b0001 : 4'b0101;
															assign node27981 = (inp[9]) ? node27983 : 4'b0111;
																assign node27983 = (inp[4]) ? 4'b0011 : 4'b0111;
													assign node27986 = (inp[3]) ? node27996 : node27987;
														assign node27987 = (inp[12]) ? 4'b0111 : node27988;
															assign node27988 = (inp[9]) ? node27992 : node27989;
																assign node27989 = (inp[4]) ? 4'b0011 : 4'b0111;
																assign node27992 = (inp[4]) ? 4'b0111 : 4'b0011;
														assign node27996 = (inp[9]) ? node28004 : node27997;
															assign node27997 = (inp[4]) ? node28001 : node27998;
																assign node27998 = (inp[12]) ? 4'b0011 : 4'b0111;
																assign node28001 = (inp[12]) ? 4'b0101 : 4'b0011;
															assign node28004 = (inp[12]) ? node28006 : 4'b0101;
																assign node28006 = (inp[4]) ? 4'b0001 : 4'b0101;
												assign node28009 = (inp[0]) ? node28027 : node28010;
													assign node28010 = (inp[3]) ? node28020 : node28011;
														assign node28011 = (inp[9]) ? 4'b0011 : node28012;
															assign node28012 = (inp[12]) ? node28016 : node28013;
																assign node28013 = (inp[4]) ? 4'b0001 : 4'b0101;
																assign node28016 = (inp[4]) ? 4'b0111 : 4'b0001;
														assign node28020 = (inp[12]) ? 4'b0111 : node28021;
															assign node28021 = (inp[4]) ? node28023 : 4'b0011;
																assign node28023 = (inp[9]) ? 4'b0111 : 4'b0011;
													assign node28027 = (inp[3]) ? node28037 : node28028;
														assign node28028 = (inp[12]) ? node28032 : node28029;
															assign node28029 = (inp[9]) ? 4'b0011 : 4'b0111;
															assign node28032 = (inp[4]) ? node28034 : 4'b0101;
																assign node28034 = (inp[9]) ? 4'b0001 : 4'b0101;
														assign node28037 = (inp[9]) ? node28045 : node28038;
															assign node28038 = (inp[4]) ? node28042 : node28039;
																assign node28039 = (inp[12]) ? 4'b0001 : 4'b0101;
																assign node28042 = (inp[12]) ? 4'b0101 : 4'b0001;
															assign node28045 = (inp[4]) ? 4'b0101 : node28046;
																assign node28046 = (inp[12]) ? 4'b0101 : 4'b0001;
							assign node28050 = (inp[7]) ? node28612 : node28051;
								assign node28051 = (inp[14]) ? node28327 : node28052;
									assign node28052 = (inp[2]) ? node28180 : node28053;
										assign node28053 = (inp[15]) ? node28109 : node28054;
											assign node28054 = (inp[5]) ? node28082 : node28055;
												assign node28055 = (inp[0]) ? node28067 : node28056;
													assign node28056 = (inp[3]) ? node28064 : node28057;
														assign node28057 = (inp[12]) ? 4'b1110 : node28058;
															assign node28058 = (inp[4]) ? node28060 : 4'b1010;
																assign node28060 = (inp[9]) ? 4'b1110 : 4'b1010;
														assign node28064 = (inp[9]) ? 4'b1000 : 4'b1010;
													assign node28067 = (inp[9]) ? node28075 : node28068;
														assign node28068 = (inp[3]) ? node28070 : 4'b1000;
															assign node28070 = (inp[12]) ? 4'b1000 : node28071;
																assign node28071 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node28075 = (inp[4]) ? node28079 : node28076;
															assign node28076 = (inp[12]) ? 4'b1100 : 4'b1000;
															assign node28079 = (inp[12]) ? 4'b1000 : 4'b1110;
												assign node28082 = (inp[0]) ? node28096 : node28083;
													assign node28083 = (inp[4]) ? node28091 : node28084;
														assign node28084 = (inp[3]) ? node28086 : 4'b1010;
															assign node28086 = (inp[9]) ? 4'b1000 : node28087;
																assign node28087 = (inp[12]) ? 4'b1000 : 4'b1100;
														assign node28091 = (inp[9]) ? node28093 : 4'b1100;
															assign node28093 = (inp[12]) ? 4'b1000 : 4'b1100;
													assign node28096 = (inp[3]) ? node28104 : node28097;
														assign node28097 = (inp[12]) ? node28099 : 4'b1000;
															assign node28099 = (inp[9]) ? node28101 : 4'b1110;
																assign node28101 = (inp[4]) ? 4'b1010 : 4'b1110;
														assign node28104 = (inp[12]) ? node28106 : 4'b1110;
															assign node28106 = (inp[4]) ? 4'b1010 : 4'b1110;
											assign node28109 = (inp[0]) ? node28143 : node28110;
												assign node28110 = (inp[5]) ? node28122 : node28111;
													assign node28111 = (inp[4]) ? node28117 : node28112;
														assign node28112 = (inp[9]) ? 4'b1000 : node28113;
															assign node28113 = (inp[12]) ? 4'b1000 : 4'b1100;
														assign node28117 = (inp[9]) ? 4'b1010 : node28118;
															assign node28118 = (inp[3]) ? 4'b1110 : 4'b1100;
													assign node28122 = (inp[3]) ? node28136 : node28123;
														assign node28123 = (inp[12]) ? node28129 : node28124;
															assign node28124 = (inp[4]) ? 4'b1000 : node28125;
																assign node28125 = (inp[9]) ? 4'b1000 : 4'b1100;
															assign node28129 = (inp[9]) ? node28133 : node28130;
																assign node28130 = (inp[4]) ? 4'b1110 : 4'b1000;
																assign node28133 = (inp[4]) ? 4'b1010 : 4'b1110;
														assign node28136 = (inp[9]) ? 4'b1110 : node28137;
															assign node28137 = (inp[4]) ? 4'b1010 : node28138;
																assign node28138 = (inp[12]) ? 4'b1010 : 4'b1110;
												assign node28143 = (inp[3]) ? node28163 : node28144;
													assign node28144 = (inp[5]) ? node28154 : node28145;
														assign node28145 = (inp[12]) ? node28147 : 4'b1110;
															assign node28147 = (inp[9]) ? node28151 : node28148;
																assign node28148 = (inp[4]) ? 4'b1110 : 4'b1010;
																assign node28151 = (inp[4]) ? 4'b1010 : 4'b1110;
														assign node28154 = (inp[12]) ? 4'b1100 : node28155;
															assign node28155 = (inp[9]) ? node28159 : node28156;
																assign node28156 = (inp[4]) ? 4'b1010 : 4'b1110;
																assign node28159 = (inp[4]) ? 4'b1100 : 4'b1010;
													assign node28163 = (inp[4]) ? node28173 : node28164;
														assign node28164 = (inp[5]) ? 4'b1000 : node28165;
															assign node28165 = (inp[12]) ? node28169 : node28166;
																assign node28166 = (inp[9]) ? 4'b1010 : 4'b1110;
																assign node28169 = (inp[9]) ? 4'b1100 : 4'b1010;
														assign node28173 = (inp[12]) ? node28177 : node28174;
															assign node28174 = (inp[9]) ? 4'b1100 : 4'b1000;
															assign node28177 = (inp[9]) ? 4'b1000 : 4'b1100;
										assign node28180 = (inp[9]) ? node28242 : node28181;
											assign node28181 = (inp[15]) ? node28211 : node28182;
												assign node28182 = (inp[12]) ? node28196 : node28183;
													assign node28183 = (inp[4]) ? 4'b0011 : node28184;
														assign node28184 = (inp[0]) ? node28190 : node28185;
															assign node28185 = (inp[3]) ? node28187 : 4'b0111;
																assign node28187 = (inp[5]) ? 4'b0101 : 4'b0111;
															assign node28190 = (inp[5]) ? node28192 : 4'b0101;
																assign node28192 = (inp[3]) ? 4'b0111 : 4'b0101;
													assign node28196 = (inp[4]) ? node28202 : node28197;
														assign node28197 = (inp[0]) ? node28199 : 4'b0011;
															assign node28199 = (inp[3]) ? 4'b0011 : 4'b0001;
														assign node28202 = (inp[5]) ? node28208 : node28203;
															assign node28203 = (inp[3]) ? 4'b0111 : node28204;
																assign node28204 = (inp[0]) ? 4'b0101 : 4'b0111;
															assign node28208 = (inp[0]) ? 4'b0111 : 4'b0101;
												assign node28211 = (inp[3]) ? node28221 : node28212;
													assign node28212 = (inp[0]) ? node28216 : node28213;
														assign node28213 = (inp[4]) ? 4'b0111 : 4'b0101;
														assign node28216 = (inp[4]) ? 4'b0011 : node28217;
															assign node28217 = (inp[12]) ? 4'b0011 : 4'b0111;
													assign node28221 = (inp[12]) ? node28233 : node28222;
														assign node28222 = (inp[4]) ? node28228 : node28223;
															assign node28223 = (inp[5]) ? 4'b0101 : node28224;
																assign node28224 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node28228 = (inp[5]) ? node28230 : 4'b0001;
																assign node28230 = (inp[0]) ? 4'b0001 : 4'b0011;
														assign node28233 = (inp[4]) ? 4'b0111 : node28234;
															assign node28234 = (inp[5]) ? node28238 : node28235;
																assign node28235 = (inp[0]) ? 4'b0011 : 4'b0001;
																assign node28238 = (inp[0]) ? 4'b0001 : 4'b0011;
											assign node28242 = (inp[5]) ? node28286 : node28243;
												assign node28243 = (inp[3]) ? node28265 : node28244;
													assign node28244 = (inp[15]) ? node28254 : node28245;
														assign node28245 = (inp[0]) ? 4'b0001 : node28246;
															assign node28246 = (inp[12]) ? node28250 : node28247;
																assign node28247 = (inp[4]) ? 4'b0111 : 4'b0011;
																assign node28250 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node28254 = (inp[0]) ? node28260 : node28255;
															assign node28255 = (inp[4]) ? node28257 : 4'b0101;
																assign node28257 = (inp[12]) ? 4'b0001 : 4'b0101;
															assign node28260 = (inp[4]) ? node28262 : 4'b0111;
																assign node28262 = (inp[12]) ? 4'b0011 : 4'b0111;
													assign node28265 = (inp[15]) ? node28279 : node28266;
														assign node28266 = (inp[0]) ? node28274 : node28267;
															assign node28267 = (inp[4]) ? node28271 : node28268;
																assign node28268 = (inp[12]) ? 4'b0101 : 4'b0011;
																assign node28271 = (inp[12]) ? 4'b0001 : 4'b0101;
															assign node28274 = (inp[4]) ? node28276 : 4'b0001;
																assign node28276 = (inp[12]) ? 4'b0011 : 4'b0111;
														assign node28279 = (inp[4]) ? node28283 : node28280;
															assign node28280 = (inp[0]) ? 4'b0011 : 4'b0001;
															assign node28283 = (inp[0]) ? 4'b0001 : 4'b0011;
												assign node28286 = (inp[3]) ? node28312 : node28287;
													assign node28287 = (inp[12]) ? node28299 : node28288;
														assign node28288 = (inp[4]) ? node28294 : node28289;
															assign node28289 = (inp[15]) ? 4'b0001 : node28290;
																assign node28290 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node28294 = (inp[0]) ? 4'b0101 : node28295;
																assign node28295 = (inp[15]) ? 4'b0111 : 4'b0101;
														assign node28299 = (inp[4]) ? node28305 : node28300;
															assign node28300 = (inp[15]) ? 4'b0101 : node28301;
																assign node28301 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node28305 = (inp[0]) ? node28309 : node28306;
																assign node28306 = (inp[15]) ? 4'b0011 : 4'b0001;
																assign node28309 = (inp[15]) ? 4'b0001 : 4'b0011;
													assign node28312 = (inp[0]) ? node28320 : node28313;
														assign node28313 = (inp[15]) ? 4'b0111 : node28314;
															assign node28314 = (inp[4]) ? node28316 : 4'b0001;
																assign node28316 = (inp[12]) ? 4'b0001 : 4'b0101;
														assign node28320 = (inp[15]) ? node28322 : 4'b0111;
															assign node28322 = (inp[4]) ? node28324 : 4'b0101;
																assign node28324 = (inp[12]) ? 4'b0001 : 4'b0101;
									assign node28327 = (inp[2]) ? node28471 : node28328;
										assign node28328 = (inp[9]) ? node28410 : node28329;
											assign node28329 = (inp[3]) ? node28373 : node28330;
												assign node28330 = (inp[4]) ? node28354 : node28331;
													assign node28331 = (inp[12]) ? node28345 : node28332;
														assign node28332 = (inp[5]) ? node28338 : node28333;
															assign node28333 = (inp[15]) ? node28335 : 4'b0101;
																assign node28335 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node28338 = (inp[15]) ? node28342 : node28339;
																assign node28339 = (inp[0]) ? 4'b0101 : 4'b0111;
																assign node28342 = (inp[0]) ? 4'b0111 : 4'b0101;
														assign node28345 = (inp[5]) ? node28347 : 4'b0011;
															assign node28347 = (inp[15]) ? node28351 : node28348;
																assign node28348 = (inp[0]) ? 4'b0001 : 4'b0011;
																assign node28351 = (inp[0]) ? 4'b0011 : 4'b0001;
													assign node28354 = (inp[12]) ? node28364 : node28355;
														assign node28355 = (inp[5]) ? 4'b0011 : node28356;
															assign node28356 = (inp[0]) ? node28360 : node28357;
																assign node28357 = (inp[15]) ? 4'b0001 : 4'b0011;
																assign node28360 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node28364 = (inp[0]) ? 4'b0111 : node28365;
															assign node28365 = (inp[5]) ? node28369 : node28366;
																assign node28366 = (inp[15]) ? 4'b0101 : 4'b0111;
																assign node28369 = (inp[15]) ? 4'b0111 : 4'b0101;
												assign node28373 = (inp[15]) ? node28393 : node28374;
													assign node28374 = (inp[4]) ? node28384 : node28375;
														assign node28375 = (inp[12]) ? node28377 : 4'b0111;
															assign node28377 = (inp[5]) ? node28381 : node28378;
																assign node28378 = (inp[0]) ? 4'b0001 : 4'b0011;
																assign node28381 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node28384 = (inp[12]) ? node28390 : node28385;
															assign node28385 = (inp[5]) ? node28387 : 4'b0001;
																assign node28387 = (inp[0]) ? 4'b0011 : 4'b0001;
															assign node28390 = (inp[0]) ? 4'b0111 : 4'b0101;
													assign node28393 = (inp[0]) ? node28405 : node28394;
														assign node28394 = (inp[5]) ? node28400 : node28395;
															assign node28395 = (inp[12]) ? node28397 : 4'b0001;
																assign node28397 = (inp[4]) ? 4'b0111 : 4'b0001;
															assign node28400 = (inp[12]) ? 4'b0111 : node28401;
																assign node28401 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node28405 = (inp[5]) ? 4'b0001 : node28406;
															assign node28406 = (inp[4]) ? 4'b0101 : 4'b0111;
											assign node28410 = (inp[15]) ? node28440 : node28411;
												assign node28411 = (inp[0]) ? node28425 : node28412;
													assign node28412 = (inp[3]) ? 4'b0101 : node28413;
														assign node28413 = (inp[5]) ? node28419 : node28414;
															assign node28414 = (inp[12]) ? node28416 : 4'b0111;
																assign node28416 = (inp[4]) ? 4'b0011 : 4'b0111;
															assign node28419 = (inp[12]) ? node28421 : 4'b0011;
																assign node28421 = (inp[4]) ? 4'b0001 : 4'b0101;
													assign node28425 = (inp[3]) ? node28433 : node28426;
														assign node28426 = (inp[4]) ? node28430 : node28427;
															assign node28427 = (inp[12]) ? 4'b0111 : 4'b0001;
															assign node28430 = (inp[12]) ? 4'b0011 : 4'b0111;
														assign node28433 = (inp[4]) ? node28437 : node28434;
															assign node28434 = (inp[12]) ? 4'b0111 : 4'b0011;
															assign node28437 = (inp[12]) ? 4'b0011 : 4'b0111;
												assign node28440 = (inp[0]) ? node28460 : node28441;
													assign node28441 = (inp[5]) ? node28451 : node28442;
														assign node28442 = (inp[12]) ? node28448 : node28443;
															assign node28443 = (inp[4]) ? node28445 : 4'b0001;
																assign node28445 = (inp[3]) ? 4'b0111 : 4'b0101;
															assign node28448 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node28451 = (inp[3]) ? node28455 : node28452;
															assign node28452 = (inp[12]) ? 4'b0011 : 4'b0111;
															assign node28455 = (inp[4]) ? 4'b0111 : node28456;
																assign node28456 = (inp[12]) ? 4'b0111 : 4'b0011;
													assign node28460 = (inp[4]) ? node28464 : node28461;
														assign node28461 = (inp[12]) ? 4'b0101 : 4'b0001;
														assign node28464 = (inp[12]) ? node28466 : 4'b0101;
															assign node28466 = (inp[5]) ? 4'b0001 : node28467;
																assign node28467 = (inp[3]) ? 4'b0001 : 4'b0011;
										assign node28471 = (inp[15]) ? node28555 : node28472;
											assign node28472 = (inp[9]) ? node28518 : node28473;
												assign node28473 = (inp[0]) ? node28497 : node28474;
													assign node28474 = (inp[3]) ? node28484 : node28475;
														assign node28475 = (inp[4]) ? node28479 : node28476;
															assign node28476 = (inp[12]) ? 4'b0011 : 4'b0111;
															assign node28479 = (inp[12]) ? node28481 : 4'b0011;
																assign node28481 = (inp[5]) ? 4'b0101 : 4'b0111;
														assign node28484 = (inp[5]) ? node28490 : node28485;
															assign node28485 = (inp[4]) ? 4'b0101 : node28486;
																assign node28486 = (inp[12]) ? 4'b0011 : 4'b0111;
															assign node28490 = (inp[4]) ? node28494 : node28491;
																assign node28491 = (inp[12]) ? 4'b0001 : 4'b0101;
																assign node28494 = (inp[12]) ? 4'b0101 : 4'b0001;
													assign node28497 = (inp[3]) ? node28505 : node28498;
														assign node28498 = (inp[4]) ? node28502 : node28499;
															assign node28499 = (inp[12]) ? 4'b0001 : 4'b0101;
															assign node28502 = (inp[12]) ? 4'b0101 : 4'b0001;
														assign node28505 = (inp[5]) ? node28513 : node28506;
															assign node28506 = (inp[12]) ? node28510 : node28507;
																assign node28507 = (inp[4]) ? 4'b0001 : 4'b0101;
																assign node28510 = (inp[4]) ? 4'b0111 : 4'b0001;
															assign node28513 = (inp[12]) ? 4'b0111 : node28514;
																assign node28514 = (inp[4]) ? 4'b0011 : 4'b0111;
												assign node28518 = (inp[0]) ? node28534 : node28519;
													assign node28519 = (inp[3]) ? node28529 : node28520;
														assign node28520 = (inp[5]) ? node28526 : node28521;
															assign node28521 = (inp[4]) ? 4'b0011 : node28522;
																assign node28522 = (inp[12]) ? 4'b0111 : 4'b0011;
															assign node28526 = (inp[12]) ? 4'b0001 : 4'b0011;
														assign node28529 = (inp[4]) ? node28531 : 4'b0101;
															assign node28531 = (inp[12]) ? 4'b0001 : 4'b0101;
													assign node28534 = (inp[3]) ? node28548 : node28535;
														assign node28535 = (inp[5]) ? node28541 : node28536;
															assign node28536 = (inp[4]) ? node28538 : 4'b0001;
																assign node28538 = (inp[12]) ? 4'b0001 : 4'b0101;
															assign node28541 = (inp[4]) ? node28545 : node28542;
																assign node28542 = (inp[12]) ? 4'b0111 : 4'b0001;
																assign node28545 = (inp[12]) ? 4'b0011 : 4'b0111;
														assign node28548 = (inp[4]) ? node28552 : node28549;
															assign node28549 = (inp[12]) ? 4'b0111 : 4'b0011;
															assign node28552 = (inp[12]) ? 4'b0011 : 4'b0111;
											assign node28555 = (inp[5]) ? node28585 : node28556;
												assign node28556 = (inp[0]) ? node28574 : node28557;
													assign node28557 = (inp[4]) ? node28567 : node28558;
														assign node28558 = (inp[3]) ? node28560 : 4'b0001;
															assign node28560 = (inp[12]) ? node28564 : node28561;
																assign node28561 = (inp[9]) ? 4'b0001 : 4'b0101;
																assign node28564 = (inp[9]) ? 4'b0111 : 4'b0001;
														assign node28567 = (inp[3]) ? node28569 : 4'b0101;
															assign node28569 = (inp[9]) ? 4'b0111 : node28570;
																assign node28570 = (inp[12]) ? 4'b0111 : 4'b0001;
													assign node28574 = (inp[9]) ? node28580 : node28575;
														assign node28575 = (inp[4]) ? 4'b0011 : node28576;
															assign node28576 = (inp[12]) ? 4'b0011 : 4'b0111;
														assign node28580 = (inp[4]) ? 4'b0001 : node28581;
															assign node28581 = (inp[3]) ? 4'b0101 : 4'b0111;
												assign node28585 = (inp[0]) ? node28597 : node28586;
													assign node28586 = (inp[3]) ? node28592 : node28587;
														assign node28587 = (inp[12]) ? node28589 : 4'b0001;
															assign node28589 = (inp[9]) ? 4'b0011 : 4'b0001;
														assign node28592 = (inp[12]) ? 4'b0011 : node28593;
															assign node28593 = (inp[4]) ? 4'b0011 : 4'b0111;
													assign node28597 = (inp[3]) ? node28603 : node28598;
														assign node28598 = (inp[12]) ? node28600 : 4'b0011;
															assign node28600 = (inp[9]) ? 4'b0101 : 4'b0011;
														assign node28603 = (inp[12]) ? 4'b0001 : node28604;
															assign node28604 = (inp[4]) ? node28608 : node28605;
																assign node28605 = (inp[9]) ? 4'b0001 : 4'b0101;
																assign node28608 = (inp[9]) ? 4'b0101 : 4'b0001;
								assign node28612 = (inp[14]) ? node28914 : node28613;
									assign node28613 = (inp[2]) ? node28761 : node28614;
										assign node28614 = (inp[12]) ? node28694 : node28615;
											assign node28615 = (inp[5]) ? node28661 : node28616;
												assign node28616 = (inp[3]) ? node28640 : node28617;
													assign node28617 = (inp[15]) ? node28627 : node28618;
														assign node28618 = (inp[0]) ? 4'b0101 : node28619;
															assign node28619 = (inp[9]) ? node28623 : node28620;
																assign node28620 = (inp[4]) ? 4'b0011 : 4'b0111;
																assign node28623 = (inp[4]) ? 4'b0111 : 4'b0011;
														assign node28627 = (inp[0]) ? node28633 : node28628;
															assign node28628 = (inp[4]) ? 4'b0001 : node28629;
																assign node28629 = (inp[9]) ? 4'b0001 : 4'b0101;
															assign node28633 = (inp[9]) ? node28637 : node28634;
																assign node28634 = (inp[4]) ? 4'b0011 : 4'b0111;
																assign node28637 = (inp[4]) ? 4'b0111 : 4'b0011;
													assign node28640 = (inp[9]) ? node28650 : node28641;
														assign node28641 = (inp[4]) ? 4'b0011 : node28642;
															assign node28642 = (inp[15]) ? node28646 : node28643;
																assign node28643 = (inp[0]) ? 4'b0101 : 4'b0111;
																assign node28646 = (inp[0]) ? 4'b0111 : 4'b0101;
														assign node28650 = (inp[4]) ? node28656 : node28651;
															assign node28651 = (inp[15]) ? 4'b0011 : node28652;
																assign node28652 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node28656 = (inp[0]) ? node28658 : 4'b0101;
																assign node28658 = (inp[15]) ? 4'b0101 : 4'b0111;
												assign node28661 = (inp[9]) ? node28681 : node28662;
													assign node28662 = (inp[4]) ? node28668 : node28663;
														assign node28663 = (inp[0]) ? 4'b0111 : node28664;
															assign node28664 = (inp[3]) ? 4'b0101 : 4'b0111;
														assign node28668 = (inp[3]) ? node28674 : node28669;
															assign node28669 = (inp[15]) ? 4'b0001 : node28670;
																assign node28670 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node28674 = (inp[15]) ? node28678 : node28675;
																assign node28675 = (inp[0]) ? 4'b0011 : 4'b0001;
																assign node28678 = (inp[0]) ? 4'b0001 : 4'b0011;
													assign node28681 = (inp[4]) ? node28687 : node28682;
														assign node28682 = (inp[0]) ? node28684 : 4'b0001;
															assign node28684 = (inp[3]) ? 4'b0011 : 4'b0001;
														assign node28687 = (inp[15]) ? node28691 : node28688;
															assign node28688 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node28691 = (inp[0]) ? 4'b0101 : 4'b0111;
											assign node28694 = (inp[0]) ? node28728 : node28695;
												assign node28695 = (inp[4]) ? node28709 : node28696;
													assign node28696 = (inp[9]) ? node28702 : node28697;
														assign node28697 = (inp[15]) ? node28699 : 4'b0011;
															assign node28699 = (inp[3]) ? 4'b0011 : 4'b0001;
														assign node28702 = (inp[5]) ? 4'b0111 : node28703;
															assign node28703 = (inp[3]) ? node28705 : 4'b0101;
																assign node28705 = (inp[15]) ? 4'b0111 : 4'b0101;
													assign node28709 = (inp[9]) ? node28719 : node28710;
														assign node28710 = (inp[3]) ? 4'b0101 : node28711;
															assign node28711 = (inp[5]) ? node28715 : node28712;
																assign node28712 = (inp[15]) ? 4'b0101 : 4'b0111;
																assign node28715 = (inp[15]) ? 4'b0111 : 4'b0101;
														assign node28719 = (inp[3]) ? node28725 : node28720;
															assign node28720 = (inp[15]) ? node28722 : 4'b0011;
																assign node28722 = (inp[5]) ? 4'b0011 : 4'b0001;
															assign node28725 = (inp[15]) ? 4'b0011 : 4'b0001;
												assign node28728 = (inp[5]) ? node28748 : node28729;
													assign node28729 = (inp[9]) ? node28737 : node28730;
														assign node28730 = (inp[4]) ? node28732 : 4'b0001;
															assign node28732 = (inp[3]) ? node28734 : 4'b0101;
																assign node28734 = (inp[15]) ? 4'b0101 : 4'b0111;
														assign node28737 = (inp[4]) ? node28745 : node28738;
															assign node28738 = (inp[3]) ? node28742 : node28739;
																assign node28739 = (inp[15]) ? 4'b0111 : 4'b0101;
																assign node28742 = (inp[15]) ? 4'b0101 : 4'b0111;
															assign node28745 = (inp[15]) ? 4'b0011 : 4'b0001;
													assign node28748 = (inp[15]) ? node28754 : node28749;
														assign node28749 = (inp[3]) ? 4'b0111 : node28750;
															assign node28750 = (inp[4]) ? 4'b0011 : 4'b0001;
														assign node28754 = (inp[9]) ? node28758 : node28755;
															assign node28755 = (inp[4]) ? 4'b0101 : 4'b0001;
															assign node28758 = (inp[4]) ? 4'b0001 : 4'b0101;
										assign node28761 = (inp[0]) ? node28839 : node28762;
											assign node28762 = (inp[5]) ? node28810 : node28763;
												assign node28763 = (inp[15]) ? node28785 : node28764;
													assign node28764 = (inp[3]) ? node28772 : node28765;
														assign node28765 = (inp[4]) ? node28767 : 4'b0110;
															assign node28767 = (inp[12]) ? 4'b0010 : node28768;
																assign node28768 = (inp[9]) ? 4'b0110 : 4'b0010;
														assign node28772 = (inp[9]) ? node28780 : node28773;
															assign node28773 = (inp[12]) ? node28777 : node28774;
																assign node28774 = (inp[4]) ? 4'b0010 : 4'b0110;
																assign node28777 = (inp[4]) ? 4'b0100 : 4'b0010;
															assign node28780 = (inp[12]) ? node28782 : 4'b0100;
																assign node28782 = (inp[4]) ? 4'b0000 : 4'b0100;
													assign node28785 = (inp[3]) ? node28797 : node28786;
														assign node28786 = (inp[4]) ? node28792 : node28787;
															assign node28787 = (inp[9]) ? 4'b0000 : node28788;
																assign node28788 = (inp[12]) ? 4'b0000 : 4'b0100;
															assign node28792 = (inp[9]) ? 4'b0100 : node28793;
																assign node28793 = (inp[12]) ? 4'b0100 : 4'b0000;
														assign node28797 = (inp[12]) ? node28803 : node28798;
															assign node28798 = (inp[4]) ? node28800 : 4'b0000;
																assign node28800 = (inp[9]) ? 4'b0110 : 4'b0000;
															assign node28803 = (inp[9]) ? node28807 : node28804;
																assign node28804 = (inp[4]) ? 4'b0110 : 4'b0000;
																assign node28807 = (inp[4]) ? 4'b0010 : 4'b0110;
												assign node28810 = (inp[15]) ? node28834 : node28811;
													assign node28811 = (inp[3]) ? node28821 : node28812;
														assign node28812 = (inp[9]) ? 4'b0100 : node28813;
															assign node28813 = (inp[4]) ? node28817 : node28814;
																assign node28814 = (inp[12]) ? 4'b0010 : 4'b0110;
																assign node28817 = (inp[12]) ? 4'b0100 : 4'b0010;
														assign node28821 = (inp[12]) ? node28829 : node28822;
															assign node28822 = (inp[4]) ? node28826 : node28823;
																assign node28823 = (inp[9]) ? 4'b0000 : 4'b0100;
																assign node28826 = (inp[9]) ? 4'b0100 : 4'b0000;
															assign node28829 = (inp[4]) ? node28831 : 4'b0000;
																assign node28831 = (inp[9]) ? 4'b0000 : 4'b0100;
													assign node28834 = (inp[12]) ? 4'b0110 : node28835;
														assign node28835 = (inp[3]) ? 4'b0110 : 4'b0100;
											assign node28839 = (inp[5]) ? node28869 : node28840;
												assign node28840 = (inp[15]) ? node28856 : node28841;
													assign node28841 = (inp[3]) ? 4'b0110 : node28842;
														assign node28842 = (inp[9]) ? node28848 : node28843;
															assign node28843 = (inp[4]) ? node28845 : 4'b0100;
																assign node28845 = (inp[12]) ? 4'b0100 : 4'b0000;
															assign node28848 = (inp[4]) ? node28852 : node28849;
																assign node28849 = (inp[12]) ? 4'b0100 : 4'b0000;
																assign node28852 = (inp[12]) ? 4'b0000 : 4'b0100;
													assign node28856 = (inp[9]) ? node28862 : node28857;
														assign node28857 = (inp[12]) ? node28859 : 4'b0110;
															assign node28859 = (inp[3]) ? 4'b0100 : 4'b0110;
														assign node28862 = (inp[3]) ? 4'b0010 : node28863;
															assign node28863 = (inp[12]) ? node28865 : 4'b0110;
																assign node28865 = (inp[4]) ? 4'b0010 : 4'b0110;
												assign node28869 = (inp[15]) ? node28895 : node28870;
													assign node28870 = (inp[3]) ? node28882 : node28871;
														assign node28871 = (inp[4]) ? node28879 : node28872;
															assign node28872 = (inp[12]) ? node28876 : node28873;
																assign node28873 = (inp[9]) ? 4'b0000 : 4'b0100;
																assign node28876 = (inp[9]) ? 4'b0110 : 4'b0000;
															assign node28879 = (inp[12]) ? 4'b0010 : 4'b0110;
														assign node28882 = (inp[4]) ? node28888 : node28883;
															assign node28883 = (inp[9]) ? 4'b0010 : node28884;
																assign node28884 = (inp[12]) ? 4'b0010 : 4'b0110;
															assign node28888 = (inp[9]) ? node28892 : node28889;
																assign node28889 = (inp[12]) ? 4'b0110 : 4'b0010;
																assign node28892 = (inp[12]) ? 4'b0010 : 4'b0110;
													assign node28895 = (inp[3]) ? node28905 : node28896;
														assign node28896 = (inp[4]) ? 4'b0000 : node28897;
															assign node28897 = (inp[9]) ? node28901 : node28898;
																assign node28898 = (inp[12]) ? 4'b0010 : 4'b0110;
																assign node28901 = (inp[12]) ? 4'b0100 : 4'b0010;
														assign node28905 = (inp[4]) ? 4'b0100 : node28906;
															assign node28906 = (inp[9]) ? node28910 : node28907;
																assign node28907 = (inp[12]) ? 4'b0000 : 4'b0100;
																assign node28910 = (inp[12]) ? 4'b0100 : 4'b0000;
									assign node28914 = (inp[12]) ? node29020 : node28915;
										assign node28915 = (inp[9]) ? node28963 : node28916;
											assign node28916 = (inp[4]) ? node28940 : node28917;
												assign node28917 = (inp[0]) ? node28929 : node28918;
													assign node28918 = (inp[15]) ? node28924 : node28919;
														assign node28919 = (inp[3]) ? node28921 : 4'b0110;
															assign node28921 = (inp[5]) ? 4'b0100 : 4'b0110;
														assign node28924 = (inp[5]) ? node28926 : 4'b0100;
															assign node28926 = (inp[3]) ? 4'b0110 : 4'b0100;
													assign node28929 = (inp[15]) ? node28933 : node28930;
														assign node28930 = (inp[5]) ? 4'b0110 : 4'b0100;
														assign node28933 = (inp[2]) ? 4'b0110 : node28934;
															assign node28934 = (inp[3]) ? node28936 : 4'b0110;
																assign node28936 = (inp[5]) ? 4'b0100 : 4'b0110;
												assign node28940 = (inp[15]) ? node28952 : node28941;
													assign node28941 = (inp[0]) ? node28947 : node28942;
														assign node28942 = (inp[3]) ? node28944 : 4'b0010;
															assign node28944 = (inp[5]) ? 4'b0000 : 4'b0010;
														assign node28947 = (inp[3]) ? node28949 : 4'b0000;
															assign node28949 = (inp[5]) ? 4'b0010 : 4'b0000;
													assign node28952 = (inp[0]) ? node28958 : node28953;
														assign node28953 = (inp[5]) ? node28955 : 4'b0000;
															assign node28955 = (inp[3]) ? 4'b0010 : 4'b0000;
														assign node28958 = (inp[5]) ? node28960 : 4'b0010;
															assign node28960 = (inp[3]) ? 4'b0000 : 4'b0010;
											assign node28963 = (inp[4]) ? node28985 : node28964;
												assign node28964 = (inp[2]) ? node28972 : node28965;
													assign node28965 = (inp[3]) ? 4'b0010 : node28966;
														assign node28966 = (inp[0]) ? 4'b0010 : node28967;
															assign node28967 = (inp[15]) ? 4'b0000 : 4'b0010;
													assign node28972 = (inp[5]) ? node28978 : node28973;
														assign node28973 = (inp[15]) ? 4'b0000 : node28974;
															assign node28974 = (inp[0]) ? 4'b0000 : 4'b0010;
														assign node28978 = (inp[15]) ? 4'b0010 : node28979;
															assign node28979 = (inp[3]) ? node28981 : 4'b0000;
																assign node28981 = (inp[0]) ? 4'b0010 : 4'b0000;
												assign node28985 = (inp[3]) ? node29007 : node28986;
													assign node28986 = (inp[5]) ? node28994 : node28987;
														assign node28987 = (inp[0]) ? node28991 : node28988;
															assign node28988 = (inp[15]) ? 4'b0100 : 4'b0110;
															assign node28991 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node28994 = (inp[2]) ? node29002 : node28995;
															assign node28995 = (inp[0]) ? node28999 : node28996;
																assign node28996 = (inp[15]) ? 4'b0110 : 4'b0100;
																assign node28999 = (inp[15]) ? 4'b0100 : 4'b0110;
															assign node29002 = (inp[0]) ? 4'b0110 : node29003;
																assign node29003 = (inp[15]) ? 4'b0110 : 4'b0100;
													assign node29007 = (inp[5]) ? node29013 : node29008;
														assign node29008 = (inp[15]) ? node29010 : 4'b0110;
															assign node29010 = (inp[0]) ? 4'b0100 : 4'b0110;
														assign node29013 = (inp[0]) ? node29017 : node29014;
															assign node29014 = (inp[15]) ? 4'b0110 : 4'b0100;
															assign node29017 = (inp[15]) ? 4'b0100 : 4'b0110;
										assign node29020 = (inp[5]) ? node29074 : node29021;
											assign node29021 = (inp[9]) ? node29043 : node29022;
												assign node29022 = (inp[4]) ? node29030 : node29023;
													assign node29023 = (inp[15]) ? node29027 : node29024;
														assign node29024 = (inp[0]) ? 4'b0000 : 4'b0010;
														assign node29027 = (inp[0]) ? 4'b0010 : 4'b0000;
													assign node29030 = (inp[2]) ? node29038 : node29031;
														assign node29031 = (inp[0]) ? 4'b0100 : node29032;
															assign node29032 = (inp[15]) ? node29034 : 4'b0110;
																assign node29034 = (inp[3]) ? 4'b0110 : 4'b0100;
														assign node29038 = (inp[3]) ? node29040 : 4'b0110;
															assign node29040 = (inp[0]) ? 4'b0110 : 4'b0100;
												assign node29043 = (inp[4]) ? node29059 : node29044;
													assign node29044 = (inp[3]) ? node29052 : node29045;
														assign node29045 = (inp[2]) ? 4'b0100 : node29046;
															assign node29046 = (inp[0]) ? 4'b0110 : node29047;
																assign node29047 = (inp[15]) ? 4'b0100 : 4'b0110;
														assign node29052 = (inp[2]) ? node29054 : 4'b0110;
															assign node29054 = (inp[0]) ? 4'b0110 : node29055;
																assign node29055 = (inp[15]) ? 4'b0110 : 4'b0100;
													assign node29059 = (inp[15]) ? node29065 : node29060;
														assign node29060 = (inp[3]) ? node29062 : 4'b0010;
															assign node29062 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node29065 = (inp[2]) ? node29067 : 4'b0000;
															assign node29067 = (inp[0]) ? node29071 : node29068;
																assign node29068 = (inp[3]) ? 4'b0010 : 4'b0000;
																assign node29071 = (inp[3]) ? 4'b0000 : 4'b0010;
											assign node29074 = (inp[0]) ? node29106 : node29075;
												assign node29075 = (inp[15]) ? node29091 : node29076;
													assign node29076 = (inp[3]) ? node29084 : node29077;
														assign node29077 = (inp[4]) ? node29081 : node29078;
															assign node29078 = (inp[9]) ? 4'b0100 : 4'b0010;
															assign node29081 = (inp[9]) ? 4'b0000 : 4'b0100;
														assign node29084 = (inp[2]) ? 4'b0000 : node29085;
															assign node29085 = (inp[9]) ? node29087 : 4'b0000;
																assign node29087 = (inp[4]) ? 4'b0000 : 4'b0100;
													assign node29091 = (inp[3]) ? node29097 : node29092;
														assign node29092 = (inp[9]) ? node29094 : 4'b0000;
															assign node29094 = (inp[4]) ? 4'b0010 : 4'b0110;
														assign node29097 = (inp[2]) ? 4'b0010 : node29098;
															assign node29098 = (inp[4]) ? node29102 : node29099;
																assign node29099 = (inp[9]) ? 4'b0110 : 4'b0010;
																assign node29102 = (inp[9]) ? 4'b0010 : 4'b0110;
												assign node29106 = (inp[15]) ? node29116 : node29107;
													assign node29107 = (inp[3]) ? 4'b0110 : node29108;
														assign node29108 = (inp[9]) ? node29112 : node29109;
															assign node29109 = (inp[4]) ? 4'b0110 : 4'b0000;
															assign node29112 = (inp[4]) ? 4'b0010 : 4'b0110;
													assign node29116 = (inp[3]) ? node29124 : node29117;
														assign node29117 = (inp[4]) ? node29121 : node29118;
															assign node29118 = (inp[9]) ? 4'b0100 : 4'b0010;
															assign node29121 = (inp[9]) ? 4'b0000 : 4'b0100;
														assign node29124 = (inp[9]) ? node29128 : node29125;
															assign node29125 = (inp[4]) ? 4'b0100 : 4'b0000;
															assign node29128 = (inp[4]) ? 4'b0000 : 4'b0100;
						assign node29131 = (inp[0]) ? node30099 : node29132;
							assign node29132 = (inp[9]) ? node29600 : node29133;
								assign node29133 = (inp[15]) ? node29355 : node29134;
									assign node29134 = (inp[3]) ? node29244 : node29135;
										assign node29135 = (inp[12]) ? node29187 : node29136;
											assign node29136 = (inp[4]) ? node29170 : node29137;
												assign node29137 = (inp[2]) ? node29153 : node29138;
													assign node29138 = (inp[8]) ? node29146 : node29139;
														assign node29139 = (inp[14]) ? node29143 : node29140;
															assign node29140 = (inp[7]) ? 4'b0110 : 4'b0111;
															assign node29143 = (inp[7]) ? 4'b0111 : 4'b0110;
														assign node29146 = (inp[14]) ? node29150 : node29147;
															assign node29147 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node29150 = (inp[7]) ? 4'b0110 : 4'b0111;
													assign node29153 = (inp[14]) ? node29163 : node29154;
														assign node29154 = (inp[5]) ? node29156 : 4'b0110;
															assign node29156 = (inp[8]) ? node29160 : node29157;
																assign node29157 = (inp[7]) ? 4'b0111 : 4'b0110;
																assign node29160 = (inp[7]) ? 4'b0110 : 4'b0111;
														assign node29163 = (inp[5]) ? 4'b0111 : node29164;
															assign node29164 = (inp[8]) ? 4'b0111 : node29165;
																assign node29165 = (inp[7]) ? 4'b0111 : 4'b0110;
												assign node29170 = (inp[8]) ? node29182 : node29171;
													assign node29171 = (inp[7]) ? node29177 : node29172;
														assign node29172 = (inp[14]) ? 4'b0010 : node29173;
															assign node29173 = (inp[2]) ? 4'b0010 : 4'b0011;
														assign node29177 = (inp[2]) ? 4'b0011 : node29178;
															assign node29178 = (inp[14]) ? 4'b0011 : 4'b0010;
													assign node29182 = (inp[7]) ? 4'b0010 : node29183;
														assign node29183 = (inp[2]) ? 4'b0011 : 4'b0010;
											assign node29187 = (inp[4]) ? node29205 : node29188;
												assign node29188 = (inp[14]) ? node29198 : node29189;
													assign node29189 = (inp[5]) ? 4'b0011 : node29190;
														assign node29190 = (inp[2]) ? node29192 : 4'b0011;
															assign node29192 = (inp[8]) ? 4'b0011 : node29193;
																assign node29193 = (inp[7]) ? 4'b0011 : 4'b0010;
													assign node29198 = (inp[8]) ? node29202 : node29199;
														assign node29199 = (inp[7]) ? 4'b0011 : 4'b0010;
														assign node29202 = (inp[7]) ? 4'b0010 : 4'b0011;
												assign node29205 = (inp[5]) ? node29229 : node29206;
													assign node29206 = (inp[7]) ? node29218 : node29207;
														assign node29207 = (inp[8]) ? node29213 : node29208;
															assign node29208 = (inp[2]) ? 4'b0110 : node29209;
																assign node29209 = (inp[14]) ? 4'b0110 : 4'b0111;
															assign node29213 = (inp[14]) ? 4'b0111 : node29214;
																assign node29214 = (inp[2]) ? 4'b0111 : 4'b0110;
														assign node29218 = (inp[8]) ? node29224 : node29219;
															assign node29219 = (inp[2]) ? 4'b0111 : node29220;
																assign node29220 = (inp[14]) ? 4'b0111 : 4'b0110;
															assign node29224 = (inp[14]) ? 4'b0110 : node29225;
																assign node29225 = (inp[2]) ? 4'b0110 : 4'b0111;
													assign node29229 = (inp[8]) ? node29241 : node29230;
														assign node29230 = (inp[7]) ? node29236 : node29231;
															assign node29231 = (inp[2]) ? 4'b0100 : node29232;
																assign node29232 = (inp[14]) ? 4'b0100 : 4'b0101;
															assign node29236 = (inp[2]) ? 4'b0101 : node29237;
																assign node29237 = (inp[14]) ? 4'b0101 : 4'b0100;
														assign node29241 = (inp[7]) ? 4'b0100 : 4'b0101;
										assign node29244 = (inp[5]) ? node29290 : node29245;
											assign node29245 = (inp[4]) ? node29265 : node29246;
												assign node29246 = (inp[12]) ? node29256 : node29247;
													assign node29247 = (inp[8]) ? 4'b0110 : node29248;
														assign node29248 = (inp[7]) ? 4'b0111 : node29249;
															assign node29249 = (inp[2]) ? 4'b0110 : node29250;
																assign node29250 = (inp[14]) ? 4'b0110 : 4'b0111;
													assign node29256 = (inp[8]) ? node29262 : node29257;
														assign node29257 = (inp[7]) ? 4'b0011 : node29258;
															assign node29258 = (inp[2]) ? 4'b0010 : 4'b0011;
														assign node29262 = (inp[7]) ? 4'b0010 : 4'b0011;
												assign node29265 = (inp[12]) ? node29273 : node29266;
													assign node29266 = (inp[8]) ? 4'b0010 : node29267;
														assign node29267 = (inp[7]) ? 4'b0011 : node29268;
															assign node29268 = (inp[14]) ? 4'b0010 : 4'b0011;
													assign node29273 = (inp[14]) ? node29283 : node29274;
														assign node29274 = (inp[7]) ? node29276 : 4'b0101;
															assign node29276 = (inp[2]) ? node29280 : node29277;
																assign node29277 = (inp[8]) ? 4'b0101 : 4'b0100;
																assign node29280 = (inp[8]) ? 4'b0100 : 4'b0101;
														assign node29283 = (inp[8]) ? node29287 : node29284;
															assign node29284 = (inp[7]) ? 4'b0101 : 4'b0100;
															assign node29287 = (inp[7]) ? 4'b0100 : 4'b0101;
											assign node29290 = (inp[14]) ? node29318 : node29291;
												assign node29291 = (inp[8]) ? node29309 : node29292;
													assign node29292 = (inp[2]) ? node29300 : node29293;
														assign node29293 = (inp[7]) ? node29295 : 4'b0001;
															assign node29295 = (inp[4]) ? node29297 : 4'b0000;
																assign node29297 = (inp[12]) ? 4'b0100 : 4'b0000;
														assign node29300 = (inp[7]) ? node29304 : node29301;
															assign node29301 = (inp[12]) ? 4'b0100 : 4'b0000;
															assign node29304 = (inp[12]) ? 4'b0101 : node29305;
																assign node29305 = (inp[4]) ? 4'b0001 : 4'b0101;
													assign node29309 = (inp[2]) ? node29315 : node29310;
														assign node29310 = (inp[4]) ? 4'b0101 : node29311;
															assign node29311 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node29315 = (inp[7]) ? 4'b0000 : 4'b0001;
												assign node29318 = (inp[8]) ? node29334 : node29319;
													assign node29319 = (inp[7]) ? node29327 : node29320;
														assign node29320 = (inp[2]) ? node29322 : 4'b0100;
															assign node29322 = (inp[4]) ? node29324 : 4'b0000;
																assign node29324 = (inp[12]) ? 4'b0100 : 4'b0000;
														assign node29327 = (inp[2]) ? 4'b0101 : node29328;
															assign node29328 = (inp[4]) ? 4'b0001 : node29329;
																assign node29329 = (inp[12]) ? 4'b0001 : 4'b0101;
													assign node29334 = (inp[7]) ? node29342 : node29335;
														assign node29335 = (inp[2]) ? node29337 : 4'b0101;
															assign node29337 = (inp[4]) ? 4'b0001 : node29338;
																assign node29338 = (inp[12]) ? 4'b0001 : 4'b0101;
														assign node29342 = (inp[2]) ? node29348 : node29343;
															assign node29343 = (inp[12]) ? 4'b0100 : node29344;
																assign node29344 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node29348 = (inp[12]) ? node29352 : node29349;
																assign node29349 = (inp[4]) ? 4'b0000 : 4'b0100;
																assign node29352 = (inp[4]) ? 4'b0100 : 4'b0000;
									assign node29355 = (inp[3]) ? node29467 : node29356;
										assign node29356 = (inp[4]) ? node29414 : node29357;
											assign node29357 = (inp[12]) ? node29389 : node29358;
												assign node29358 = (inp[5]) ? node29366 : node29359;
													assign node29359 = (inp[8]) ? 4'b0100 : node29360;
														assign node29360 = (inp[2]) ? node29362 : 4'b0101;
															assign node29362 = (inp[7]) ? 4'b0101 : 4'b0100;
													assign node29366 = (inp[2]) ? node29382 : node29367;
														assign node29367 = (inp[14]) ? node29375 : node29368;
															assign node29368 = (inp[7]) ? node29372 : node29369;
																assign node29369 = (inp[8]) ? 4'b0100 : 4'b0101;
																assign node29372 = (inp[8]) ? 4'b0101 : 4'b0100;
															assign node29375 = (inp[7]) ? node29379 : node29376;
																assign node29376 = (inp[8]) ? 4'b0101 : 4'b0100;
																assign node29379 = (inp[8]) ? 4'b0100 : 4'b0101;
														assign node29382 = (inp[7]) ? node29386 : node29383;
															assign node29383 = (inp[8]) ? 4'b0101 : 4'b0100;
															assign node29386 = (inp[8]) ? 4'b0100 : 4'b0101;
												assign node29389 = (inp[8]) ? node29403 : node29390;
													assign node29390 = (inp[5]) ? node29396 : node29391;
														assign node29391 = (inp[7]) ? node29393 : 4'b0000;
															assign node29393 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node29396 = (inp[2]) ? 4'b0000 : node29397;
															assign node29397 = (inp[14]) ? 4'b0001 : node29398;
																assign node29398 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node29403 = (inp[2]) ? node29411 : node29404;
														assign node29404 = (inp[7]) ? node29408 : node29405;
															assign node29405 = (inp[14]) ? 4'b0001 : 4'b0000;
															assign node29408 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node29411 = (inp[7]) ? 4'b0000 : 4'b0001;
											assign node29414 = (inp[12]) ? node29438 : node29415;
												assign node29415 = (inp[8]) ? node29429 : node29416;
													assign node29416 = (inp[5]) ? node29424 : node29417;
														assign node29417 = (inp[7]) ? node29421 : node29418;
															assign node29418 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node29421 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node29424 = (inp[2]) ? 4'b0000 : node29425;
															assign node29425 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node29429 = (inp[7]) ? node29433 : node29430;
														assign node29430 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node29433 = (inp[2]) ? 4'b0000 : node29434;
															assign node29434 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node29438 = (inp[5]) ? node29454 : node29439;
													assign node29439 = (inp[7]) ? node29445 : node29440;
														assign node29440 = (inp[8]) ? node29442 : 4'b0100;
															assign node29442 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node29445 = (inp[8]) ? node29451 : node29446;
															assign node29446 = (inp[14]) ? 4'b0101 : node29447;
																assign node29447 = (inp[2]) ? 4'b0101 : 4'b0100;
															assign node29451 = (inp[2]) ? 4'b0100 : 4'b0101;
													assign node29454 = (inp[14]) ? 4'b0111 : node29455;
														assign node29455 = (inp[7]) ? node29461 : node29456;
															assign node29456 = (inp[2]) ? node29458 : 4'b0111;
																assign node29458 = (inp[8]) ? 4'b0111 : 4'b0110;
															assign node29461 = (inp[8]) ? 4'b0110 : node29462;
																assign node29462 = (inp[2]) ? 4'b0111 : 4'b0110;
										assign node29467 = (inp[5]) ? node29529 : node29468;
											assign node29468 = (inp[12]) ? node29502 : node29469;
												assign node29469 = (inp[4]) ? node29487 : node29470;
													assign node29470 = (inp[8]) ? node29482 : node29471;
														assign node29471 = (inp[7]) ? node29477 : node29472;
															assign node29472 = (inp[14]) ? 4'b0100 : node29473;
																assign node29473 = (inp[2]) ? 4'b0100 : 4'b0101;
															assign node29477 = (inp[14]) ? 4'b0101 : node29478;
																assign node29478 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node29482 = (inp[7]) ? node29484 : 4'b0101;
															assign node29484 = (inp[14]) ? 4'b0100 : 4'b0101;
													assign node29487 = (inp[14]) ? node29495 : node29488;
														assign node29488 = (inp[8]) ? 4'b0000 : node29489;
															assign node29489 = (inp[2]) ? node29491 : 4'b0000;
																assign node29491 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node29495 = (inp[7]) ? node29499 : node29496;
															assign node29496 = (inp[8]) ? 4'b0001 : 4'b0000;
															assign node29499 = (inp[8]) ? 4'b0000 : 4'b0001;
												assign node29502 = (inp[4]) ? node29510 : node29503;
													assign node29503 = (inp[7]) ? node29505 : 4'b0000;
														assign node29505 = (inp[8]) ? 4'b0000 : node29506;
															assign node29506 = (inp[2]) ? 4'b0001 : 4'b0000;
													assign node29510 = (inp[14]) ? node29520 : node29511;
														assign node29511 = (inp[8]) ? 4'b0111 : node29512;
															assign node29512 = (inp[2]) ? node29516 : node29513;
																assign node29513 = (inp[7]) ? 4'b0110 : 4'b0111;
																assign node29516 = (inp[7]) ? 4'b0111 : 4'b0110;
														assign node29520 = (inp[2]) ? node29522 : 4'b0110;
															assign node29522 = (inp[7]) ? node29526 : node29523;
																assign node29523 = (inp[8]) ? 4'b0111 : 4'b0110;
																assign node29526 = (inp[8]) ? 4'b0110 : 4'b0111;
											assign node29529 = (inp[2]) ? node29571 : node29530;
												assign node29530 = (inp[8]) ? node29554 : node29531;
													assign node29531 = (inp[7]) ? node29541 : node29532;
														assign node29532 = (inp[14]) ? 4'b0010 : node29533;
															assign node29533 = (inp[4]) ? node29537 : node29534;
																assign node29534 = (inp[12]) ? 4'b0011 : 4'b0111;
																assign node29537 = (inp[12]) ? 4'b0111 : 4'b0011;
														assign node29541 = (inp[14]) ? node29549 : node29542;
															assign node29542 = (inp[4]) ? node29546 : node29543;
																assign node29543 = (inp[12]) ? 4'b0010 : 4'b0110;
																assign node29546 = (inp[12]) ? 4'b0110 : 4'b0010;
															assign node29549 = (inp[12]) ? 4'b0111 : node29550;
																assign node29550 = (inp[4]) ? 4'b0011 : 4'b0111;
													assign node29554 = (inp[7]) ? node29562 : node29555;
														assign node29555 = (inp[14]) ? 4'b0111 : node29556;
															assign node29556 = (inp[4]) ? node29558 : 4'b0010;
																assign node29558 = (inp[12]) ? 4'b0110 : 4'b0010;
														assign node29562 = (inp[14]) ? node29566 : node29563;
															assign node29563 = (inp[4]) ? 4'b0111 : 4'b0011;
															assign node29566 = (inp[12]) ? 4'b0010 : node29567;
																assign node29567 = (inp[4]) ? 4'b0010 : 4'b0110;
												assign node29571 = (inp[12]) ? node29591 : node29572;
													assign node29572 = (inp[4]) ? node29586 : node29573;
														assign node29573 = (inp[14]) ? node29581 : node29574;
															assign node29574 = (inp[8]) ? node29578 : node29575;
																assign node29575 = (inp[7]) ? 4'b0111 : 4'b0110;
																assign node29578 = (inp[7]) ? 4'b0110 : 4'b0111;
															assign node29581 = (inp[8]) ? node29583 : 4'b0110;
																assign node29583 = (inp[7]) ? 4'b0110 : 4'b0111;
														assign node29586 = (inp[7]) ? node29588 : 4'b0010;
															assign node29588 = (inp[8]) ? 4'b0010 : 4'b0011;
													assign node29591 = (inp[4]) ? node29593 : 4'b0011;
														assign node29593 = (inp[8]) ? node29597 : node29594;
															assign node29594 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node29597 = (inp[7]) ? 4'b0110 : 4'b0111;
								assign node29600 = (inp[15]) ? node29846 : node29601;
									assign node29601 = (inp[5]) ? node29735 : node29602;
										assign node29602 = (inp[3]) ? node29670 : node29603;
											assign node29603 = (inp[2]) ? node29645 : node29604;
												assign node29604 = (inp[14]) ? node29620 : node29605;
													assign node29605 = (inp[4]) ? node29613 : node29606;
														assign node29606 = (inp[7]) ? node29610 : node29607;
															assign node29607 = (inp[8]) ? 4'b0110 : 4'b0111;
															assign node29610 = (inp[8]) ? 4'b0111 : 4'b0110;
														assign node29613 = (inp[7]) ? node29617 : node29614;
															assign node29614 = (inp[8]) ? 4'b0010 : 4'b0011;
															assign node29617 = (inp[8]) ? 4'b0111 : 4'b0110;
													assign node29620 = (inp[12]) ? node29634 : node29621;
														assign node29621 = (inp[4]) ? node29627 : node29622;
															assign node29622 = (inp[8]) ? 4'b0011 : node29623;
																assign node29623 = (inp[7]) ? 4'b0011 : 4'b0010;
															assign node29627 = (inp[8]) ? node29631 : node29628;
																assign node29628 = (inp[7]) ? 4'b0111 : 4'b0110;
																assign node29631 = (inp[7]) ? 4'b0110 : 4'b0111;
														assign node29634 = (inp[4]) ? node29640 : node29635;
															assign node29635 = (inp[7]) ? 4'b0110 : node29636;
																assign node29636 = (inp[8]) ? 4'b0111 : 4'b0110;
															assign node29640 = (inp[7]) ? node29642 : 4'b0011;
																assign node29642 = (inp[8]) ? 4'b0010 : 4'b0011;
												assign node29645 = (inp[8]) ? node29655 : node29646;
													assign node29646 = (inp[7]) ? node29652 : node29647;
														assign node29647 = (inp[12]) ? node29649 : 4'b0110;
															assign node29649 = (inp[4]) ? 4'b0010 : 4'b0110;
														assign node29652 = (inp[14]) ? 4'b0111 : 4'b0011;
													assign node29655 = (inp[7]) ? node29663 : node29656;
														assign node29656 = (inp[12]) ? node29660 : node29657;
															assign node29657 = (inp[4]) ? 4'b0111 : 4'b0011;
															assign node29660 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node29663 = (inp[4]) ? node29667 : node29664;
															assign node29664 = (inp[12]) ? 4'b0110 : 4'b0010;
															assign node29667 = (inp[12]) ? 4'b0010 : 4'b0110;
											assign node29670 = (inp[4]) ? node29710 : node29671;
												assign node29671 = (inp[12]) ? node29697 : node29672;
													assign node29672 = (inp[14]) ? node29686 : node29673;
														assign node29673 = (inp[7]) ? node29681 : node29674;
															assign node29674 = (inp[2]) ? node29678 : node29675;
																assign node29675 = (inp[8]) ? 4'b0010 : 4'b0011;
																assign node29678 = (inp[8]) ? 4'b0011 : 4'b0010;
															assign node29681 = (inp[8]) ? node29683 : 4'b0010;
																assign node29683 = (inp[2]) ? 4'b0010 : 4'b0011;
														assign node29686 = (inp[2]) ? node29692 : node29687;
															assign node29687 = (inp[7]) ? node29689 : 4'b0010;
																assign node29689 = (inp[8]) ? 4'b0010 : 4'b0011;
															assign node29692 = (inp[8]) ? node29694 : 4'b0010;
																assign node29694 = (inp[7]) ? 4'b0010 : 4'b0011;
													assign node29697 = (inp[8]) ? node29705 : node29698;
														assign node29698 = (inp[2]) ? 4'b0101 : node29699;
															assign node29699 = (inp[14]) ? node29701 : 4'b0100;
																assign node29701 = (inp[7]) ? 4'b0101 : 4'b0100;
														assign node29705 = (inp[7]) ? node29707 : 4'b0101;
															assign node29707 = (inp[14]) ? 4'b0100 : 4'b0101;
												assign node29710 = (inp[12]) ? node29728 : node29711;
													assign node29711 = (inp[2]) ? node29723 : node29712;
														assign node29712 = (inp[7]) ? node29718 : node29713;
															assign node29713 = (inp[8]) ? 4'b0100 : node29714;
																assign node29714 = (inp[14]) ? 4'b0100 : 4'b0101;
															assign node29718 = (inp[8]) ? 4'b0101 : node29719;
																assign node29719 = (inp[14]) ? 4'b0101 : 4'b0100;
														assign node29723 = (inp[8]) ? node29725 : 4'b0101;
															assign node29725 = (inp[7]) ? 4'b0100 : 4'b0101;
													assign node29728 = (inp[8]) ? 4'b0000 : node29729;
														assign node29729 = (inp[14]) ? node29731 : 4'b0000;
															assign node29731 = (inp[7]) ? 4'b0001 : 4'b0000;
										assign node29735 = (inp[3]) ? node29791 : node29736;
											assign node29736 = (inp[4]) ? node29762 : node29737;
												assign node29737 = (inp[12]) ? node29755 : node29738;
													assign node29738 = (inp[14]) ? node29748 : node29739;
														assign node29739 = (inp[2]) ? node29741 : 4'b0010;
															assign node29741 = (inp[8]) ? node29745 : node29742;
																assign node29742 = (inp[7]) ? 4'b0011 : 4'b0010;
																assign node29745 = (inp[7]) ? 4'b0010 : 4'b0011;
														assign node29748 = (inp[2]) ? node29750 : 4'b0011;
															assign node29750 = (inp[7]) ? 4'b0010 : node29751;
																assign node29751 = (inp[8]) ? 4'b0011 : 4'b0010;
													assign node29755 = (inp[8]) ? node29759 : node29756;
														assign node29756 = (inp[7]) ? 4'b0101 : 4'b0100;
														assign node29759 = (inp[7]) ? 4'b0100 : 4'b0101;
												assign node29762 = (inp[12]) ? node29776 : node29763;
													assign node29763 = (inp[2]) ? node29769 : node29764;
														assign node29764 = (inp[14]) ? 4'b0100 : node29765;
															assign node29765 = (inp[8]) ? 4'b0101 : 4'b0100;
														assign node29769 = (inp[7]) ? node29773 : node29770;
															assign node29770 = (inp[8]) ? 4'b0101 : 4'b0100;
															assign node29773 = (inp[8]) ? 4'b0100 : 4'b0101;
													assign node29776 = (inp[14]) ? node29782 : node29777;
														assign node29777 = (inp[8]) ? 4'b0000 : node29778;
															assign node29778 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node29782 = (inp[2]) ? 4'b0001 : node29783;
															assign node29783 = (inp[8]) ? node29787 : node29784;
																assign node29784 = (inp[7]) ? 4'b0001 : 4'b0000;
																assign node29787 = (inp[7]) ? 4'b0000 : 4'b0001;
											assign node29791 = (inp[7]) ? node29817 : node29792;
												assign node29792 = (inp[8]) ? node29802 : node29793;
													assign node29793 = (inp[14]) ? node29795 : 4'b0000;
														assign node29795 = (inp[12]) ? node29799 : node29796;
															assign node29796 = (inp[4]) ? 4'b0100 : 4'b0000;
															assign node29799 = (inp[4]) ? 4'b0000 : 4'b0100;
													assign node29802 = (inp[14]) ? node29812 : node29803;
														assign node29803 = (inp[2]) ? node29809 : node29804;
															assign node29804 = (inp[12]) ? 4'b0100 : node29805;
																assign node29805 = (inp[4]) ? 4'b0100 : 4'b0000;
															assign node29809 = (inp[4]) ? 4'b0101 : 4'b0001;
														assign node29812 = (inp[12]) ? node29814 : 4'b0001;
															assign node29814 = (inp[4]) ? 4'b0001 : 4'b0101;
												assign node29817 = (inp[8]) ? node29837 : node29818;
													assign node29818 = (inp[14]) ? node29830 : node29819;
														assign node29819 = (inp[2]) ? node29825 : node29820;
															assign node29820 = (inp[12]) ? node29822 : 4'b0100;
																assign node29822 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node29825 = (inp[12]) ? node29827 : 4'b0001;
																assign node29827 = (inp[4]) ? 4'b0001 : 4'b0101;
														assign node29830 = (inp[12]) ? node29834 : node29831;
															assign node29831 = (inp[4]) ? 4'b0101 : 4'b0001;
															assign node29834 = (inp[4]) ? 4'b0001 : 4'b0101;
													assign node29837 = (inp[14]) ? node29841 : node29838;
														assign node29838 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node29841 = (inp[2]) ? node29843 : 4'b0000;
															assign node29843 = (inp[4]) ? 4'b0100 : 4'b0000;
									assign node29846 = (inp[3]) ? node29968 : node29847;
										assign node29847 = (inp[5]) ? node29909 : node29848;
											assign node29848 = (inp[8]) ? node29880 : node29849;
												assign node29849 = (inp[7]) ? node29863 : node29850;
													assign node29850 = (inp[2]) ? node29858 : node29851;
														assign node29851 = (inp[14]) ? node29853 : 4'b0001;
															assign node29853 = (inp[12]) ? node29855 : 4'b0100;
																assign node29855 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node29858 = (inp[4]) ? 4'b0100 : node29859;
															assign node29859 = (inp[12]) ? 4'b0100 : 4'b0000;
													assign node29863 = (inp[14]) ? node29873 : node29864;
														assign node29864 = (inp[2]) ? node29870 : node29865;
															assign node29865 = (inp[4]) ? node29867 : 4'b0000;
																assign node29867 = (inp[12]) ? 4'b0000 : 4'b0100;
															assign node29870 = (inp[12]) ? 4'b0101 : 4'b0001;
														assign node29873 = (inp[12]) ? node29877 : node29874;
															assign node29874 = (inp[4]) ? 4'b0101 : 4'b0001;
															assign node29877 = (inp[2]) ? 4'b0001 : 4'b0101;
												assign node29880 = (inp[7]) ? node29894 : node29881;
													assign node29881 = (inp[2]) ? node29889 : node29882;
														assign node29882 = (inp[14]) ? 4'b0001 : node29883;
															assign node29883 = (inp[12]) ? node29885 : 4'b0000;
																assign node29885 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node29889 = (inp[4]) ? node29891 : 4'b0001;
															assign node29891 = (inp[14]) ? 4'b0001 : 4'b0101;
													assign node29894 = (inp[14]) ? node29904 : node29895;
														assign node29895 = (inp[2]) ? node29901 : node29896;
															assign node29896 = (inp[12]) ? 4'b0001 : node29897;
																assign node29897 = (inp[4]) ? 4'b0101 : 4'b0001;
															assign node29901 = (inp[12]) ? 4'b0000 : 4'b0100;
														assign node29904 = (inp[12]) ? node29906 : 4'b0000;
															assign node29906 = (inp[4]) ? 4'b0000 : 4'b0100;
											assign node29909 = (inp[12]) ? node29939 : node29910;
												assign node29910 = (inp[4]) ? node29928 : node29911;
													assign node29911 = (inp[2]) ? node29923 : node29912;
														assign node29912 = (inp[7]) ? node29918 : node29913;
															assign node29913 = (inp[8]) ? node29915 : 4'b0001;
																assign node29915 = (inp[14]) ? 4'b0001 : 4'b0000;
															assign node29918 = (inp[8]) ? 4'b0000 : node29919;
																assign node29919 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node29923 = (inp[14]) ? node29925 : 4'b0001;
															assign node29925 = (inp[7]) ? 4'b0001 : 4'b0000;
													assign node29928 = (inp[7]) ? node29932 : node29929;
														assign node29929 = (inp[8]) ? 4'b0111 : 4'b0110;
														assign node29932 = (inp[8]) ? node29934 : 4'b0111;
															assign node29934 = (inp[2]) ? 4'b0110 : node29935;
																assign node29935 = (inp[14]) ? 4'b0110 : 4'b0111;
												assign node29939 = (inp[4]) ? node29959 : node29940;
													assign node29940 = (inp[14]) ? node29954 : node29941;
														assign node29941 = (inp[7]) ? node29947 : node29942;
															assign node29942 = (inp[2]) ? 4'b0111 : node29943;
																assign node29943 = (inp[8]) ? 4'b0110 : 4'b0111;
															assign node29947 = (inp[2]) ? node29951 : node29948;
																assign node29948 = (inp[8]) ? 4'b0111 : 4'b0110;
																assign node29951 = (inp[8]) ? 4'b0110 : 4'b0111;
														assign node29954 = (inp[2]) ? node29956 : 4'b0111;
															assign node29956 = (inp[8]) ? 4'b0111 : 4'b0110;
													assign node29959 = (inp[8]) ? node29961 : 4'b0010;
														assign node29961 = (inp[7]) ? 4'b0010 : node29962;
															assign node29962 = (inp[2]) ? 4'b0011 : node29963;
																assign node29963 = (inp[14]) ? 4'b0011 : 4'b0010;
										assign node29968 = (inp[4]) ? node30028 : node29969;
											assign node29969 = (inp[12]) ? node30007 : node29970;
												assign node29970 = (inp[5]) ? node29992 : node29971;
													assign node29971 = (inp[2]) ? node29983 : node29972;
														assign node29972 = (inp[7]) ? node29978 : node29973;
															assign node29973 = (inp[8]) ? node29975 : 4'b0000;
																assign node29975 = (inp[14]) ? 4'b0001 : 4'b0000;
															assign node29978 = (inp[8]) ? node29980 : 4'b0001;
																assign node29980 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node29983 = (inp[14]) ? node29987 : node29984;
															assign node29984 = (inp[7]) ? 4'b0000 : 4'b0001;
															assign node29987 = (inp[8]) ? 4'b0001 : node29988;
																assign node29988 = (inp[7]) ? 4'b0001 : 4'b0000;
													assign node29992 = (inp[8]) ? node30004 : node29993;
														assign node29993 = (inp[7]) ? node29999 : node29994;
															assign node29994 = (inp[14]) ? 4'b0010 : node29995;
																assign node29995 = (inp[2]) ? 4'b0010 : 4'b0011;
															assign node29999 = (inp[14]) ? 4'b0011 : node30000;
																assign node30000 = (inp[2]) ? 4'b0011 : 4'b0010;
														assign node30004 = (inp[7]) ? 4'b0010 : 4'b0011;
												assign node30007 = (inp[7]) ? node30019 : node30008;
													assign node30008 = (inp[8]) ? node30014 : node30009;
														assign node30009 = (inp[2]) ? 4'b0110 : node30010;
															assign node30010 = (inp[14]) ? 4'b0110 : 4'b0111;
														assign node30014 = (inp[2]) ? 4'b0111 : node30015;
															assign node30015 = (inp[14]) ? 4'b0111 : 4'b0110;
													assign node30019 = (inp[14]) ? 4'b0111 : node30020;
														assign node30020 = (inp[8]) ? node30024 : node30021;
															assign node30021 = (inp[2]) ? 4'b0111 : 4'b0110;
															assign node30024 = (inp[2]) ? 4'b0110 : 4'b0111;
											assign node30028 = (inp[12]) ? node30068 : node30029;
												assign node30029 = (inp[5]) ? node30049 : node30030;
													assign node30030 = (inp[2]) ? node30044 : node30031;
														assign node30031 = (inp[7]) ? node30039 : node30032;
															assign node30032 = (inp[8]) ? node30036 : node30033;
																assign node30033 = (inp[14]) ? 4'b0110 : 4'b0111;
																assign node30036 = (inp[14]) ? 4'b0111 : 4'b0110;
															assign node30039 = (inp[14]) ? 4'b0111 : node30040;
																assign node30040 = (inp[8]) ? 4'b0111 : 4'b0110;
														assign node30044 = (inp[8]) ? node30046 : 4'b0110;
															assign node30046 = (inp[7]) ? 4'b0110 : 4'b0111;
													assign node30049 = (inp[2]) ? node30055 : node30050;
														assign node30050 = (inp[7]) ? node30052 : 4'b0110;
															assign node30052 = (inp[8]) ? 4'b0110 : 4'b0111;
														assign node30055 = (inp[14]) ? node30063 : node30056;
															assign node30056 = (inp[8]) ? node30060 : node30057;
																assign node30057 = (inp[7]) ? 4'b0111 : 4'b0110;
																assign node30060 = (inp[7]) ? 4'b0110 : 4'b0111;
															assign node30063 = (inp[7]) ? 4'b0110 : node30064;
																assign node30064 = (inp[8]) ? 4'b0111 : 4'b0110;
												assign node30068 = (inp[5]) ? node30082 : node30069;
													assign node30069 = (inp[8]) ? node30075 : node30070;
														assign node30070 = (inp[7]) ? node30072 : 4'b0010;
															assign node30072 = (inp[14]) ? 4'b0011 : 4'b0010;
														assign node30075 = (inp[7]) ? node30079 : node30076;
															assign node30076 = (inp[14]) ? 4'b0011 : 4'b0010;
															assign node30079 = (inp[2]) ? 4'b0010 : 4'b0011;
													assign node30082 = (inp[14]) ? node30094 : node30083;
														assign node30083 = (inp[2]) ? node30089 : node30084;
															assign node30084 = (inp[8]) ? 4'b0011 : node30085;
																assign node30085 = (inp[7]) ? 4'b0010 : 4'b0011;
															assign node30089 = (inp[8]) ? 4'b0010 : node30090;
																assign node30090 = (inp[7]) ? 4'b0011 : 4'b0010;
														assign node30094 = (inp[7]) ? 4'b0011 : node30095;
															assign node30095 = (inp[8]) ? 4'b0011 : 4'b0010;
							assign node30099 = (inp[14]) ? node30687 : node30100;
								assign node30100 = (inp[9]) ? node30386 : node30101;
									assign node30101 = (inp[15]) ? node30249 : node30102;
										assign node30102 = (inp[3]) ? node30170 : node30103;
											assign node30103 = (inp[2]) ? node30141 : node30104;
												assign node30104 = (inp[5]) ? node30128 : node30105;
													assign node30105 = (inp[8]) ? node30119 : node30106;
														assign node30106 = (inp[7]) ? node30114 : node30107;
															assign node30107 = (inp[4]) ? node30111 : node30108;
																assign node30108 = (inp[12]) ? 4'b0001 : 4'b0101;
																assign node30111 = (inp[12]) ? 4'b0101 : 4'b0001;
															assign node30114 = (inp[12]) ? node30116 : 4'b0100;
																assign node30116 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node30119 = (inp[7]) ? 4'b0101 : node30120;
															assign node30120 = (inp[4]) ? node30124 : node30121;
																assign node30121 = (inp[12]) ? 4'b0000 : 4'b0100;
																assign node30124 = (inp[12]) ? 4'b0100 : 4'b0000;
													assign node30128 = (inp[12]) ? node30138 : node30129;
														assign node30129 = (inp[4]) ? 4'b0001 : node30130;
															assign node30130 = (inp[7]) ? node30134 : node30131;
																assign node30131 = (inp[8]) ? 4'b0100 : 4'b0101;
																assign node30134 = (inp[8]) ? 4'b0101 : 4'b0100;
														assign node30138 = (inp[7]) ? 4'b0111 : 4'b0110;
												assign node30141 = (inp[4]) ? node30153 : node30142;
													assign node30142 = (inp[12]) ? node30146 : node30143;
														assign node30143 = (inp[5]) ? 4'b0101 : 4'b0100;
														assign node30146 = (inp[8]) ? node30150 : node30147;
															assign node30147 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node30150 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node30153 = (inp[12]) ? node30163 : node30154;
														assign node30154 = (inp[5]) ? node30156 : 4'b0000;
															assign node30156 = (inp[8]) ? node30160 : node30157;
																assign node30157 = (inp[7]) ? 4'b0001 : 4'b0000;
																assign node30160 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node30163 = (inp[5]) ? 4'b0110 : node30164;
															assign node30164 = (inp[7]) ? node30166 : 4'b0101;
																assign node30166 = (inp[8]) ? 4'b0100 : 4'b0101;
											assign node30170 = (inp[5]) ? node30214 : node30171;
												assign node30171 = (inp[4]) ? node30193 : node30172;
													assign node30172 = (inp[12]) ? node30180 : node30173;
														assign node30173 = (inp[7]) ? 4'b0101 : node30174;
															assign node30174 = (inp[2]) ? 4'b0100 : node30175;
																assign node30175 = (inp[8]) ? 4'b0100 : 4'b0101;
														assign node30180 = (inp[7]) ? node30186 : node30181;
															assign node30181 = (inp[8]) ? node30183 : 4'b0001;
																assign node30183 = (inp[2]) ? 4'b0001 : 4'b0000;
															assign node30186 = (inp[8]) ? node30190 : node30187;
																assign node30187 = (inp[2]) ? 4'b0001 : 4'b0000;
																assign node30190 = (inp[2]) ? 4'b0000 : 4'b0001;
													assign node30193 = (inp[12]) ? node30205 : node30194;
														assign node30194 = (inp[2]) ? node30200 : node30195;
															assign node30195 = (inp[7]) ? 4'b0001 : node30196;
																assign node30196 = (inp[8]) ? 4'b0000 : 4'b0001;
															assign node30200 = (inp[7]) ? 4'b0000 : node30201;
																assign node30201 = (inp[8]) ? 4'b0001 : 4'b0000;
														assign node30205 = (inp[2]) ? node30207 : 4'b0110;
															assign node30207 = (inp[7]) ? node30211 : node30208;
																assign node30208 = (inp[8]) ? 4'b0111 : 4'b0110;
																assign node30211 = (inp[8]) ? 4'b0110 : 4'b0111;
												assign node30214 = (inp[2]) ? node30230 : node30215;
													assign node30215 = (inp[4]) ? node30223 : node30216;
														assign node30216 = (inp[12]) ? 4'b0011 : node30217;
															assign node30217 = (inp[7]) ? node30219 : 4'b0110;
																assign node30219 = (inp[8]) ? 4'b0111 : 4'b0110;
														assign node30223 = (inp[12]) ? 4'b0110 : node30224;
															assign node30224 = (inp[8]) ? node30226 : 4'b0010;
																assign node30226 = (inp[7]) ? 4'b0011 : 4'b0010;
													assign node30230 = (inp[4]) ? node30240 : node30231;
														assign node30231 = (inp[12]) ? node30233 : 4'b0111;
															assign node30233 = (inp[8]) ? node30237 : node30234;
																assign node30234 = (inp[7]) ? 4'b0011 : 4'b0010;
																assign node30237 = (inp[7]) ? 4'b0010 : 4'b0011;
														assign node30240 = (inp[12]) ? node30244 : node30241;
															assign node30241 = (inp[8]) ? 4'b0010 : 4'b0011;
															assign node30244 = (inp[7]) ? 4'b0111 : node30245;
																assign node30245 = (inp[8]) ? 4'b0111 : 4'b0110;
										assign node30249 = (inp[3]) ? node30317 : node30250;
											assign node30250 = (inp[4]) ? node30274 : node30251;
												assign node30251 = (inp[12]) ? node30261 : node30252;
													assign node30252 = (inp[7]) ? node30254 : 4'b0110;
														assign node30254 = (inp[5]) ? 4'b0111 : node30255;
															assign node30255 = (inp[8]) ? node30257 : 4'b0110;
																assign node30257 = (inp[2]) ? 4'b0110 : 4'b0111;
													assign node30261 = (inp[7]) ? node30269 : node30262;
														assign node30262 = (inp[2]) ? node30266 : node30263;
															assign node30263 = (inp[8]) ? 4'b0010 : 4'b0011;
															assign node30266 = (inp[8]) ? 4'b0011 : 4'b0010;
														assign node30269 = (inp[2]) ? node30271 : 4'b0010;
															assign node30271 = (inp[8]) ? 4'b0010 : 4'b0011;
												assign node30274 = (inp[12]) ? node30294 : node30275;
													assign node30275 = (inp[5]) ? node30283 : node30276;
														assign node30276 = (inp[8]) ? 4'b0011 : node30277;
															assign node30277 = (inp[7]) ? 4'b0011 : node30278;
																assign node30278 = (inp[2]) ? 4'b0010 : 4'b0011;
														assign node30283 = (inp[2]) ? node30289 : node30284;
															assign node30284 = (inp[8]) ? node30286 : 4'b0011;
																assign node30286 = (inp[7]) ? 4'b0011 : 4'b0010;
															assign node30289 = (inp[8]) ? node30291 : 4'b0010;
																assign node30291 = (inp[7]) ? 4'b0010 : 4'b0011;
													assign node30294 = (inp[5]) ? node30308 : node30295;
														assign node30295 = (inp[7]) ? node30301 : node30296;
															assign node30296 = (inp[2]) ? node30298 : 4'b0111;
																assign node30298 = (inp[8]) ? 4'b0111 : 4'b0110;
															assign node30301 = (inp[8]) ? node30305 : node30302;
																assign node30302 = (inp[2]) ? 4'b0111 : 4'b0110;
																assign node30305 = (inp[2]) ? 4'b0110 : 4'b0111;
														assign node30308 = (inp[8]) ? 4'b0101 : node30309;
															assign node30309 = (inp[2]) ? node30313 : node30310;
																assign node30310 = (inp[7]) ? 4'b0100 : 4'b0101;
																assign node30313 = (inp[7]) ? 4'b0101 : 4'b0100;
											assign node30317 = (inp[5]) ? node30349 : node30318;
												assign node30318 = (inp[12]) ? node30334 : node30319;
													assign node30319 = (inp[4]) ? node30327 : node30320;
														assign node30320 = (inp[2]) ? 4'b0111 : node30321;
															assign node30321 = (inp[8]) ? 4'b0110 : node30322;
																assign node30322 = (inp[7]) ? 4'b0110 : 4'b0111;
														assign node30327 = (inp[2]) ? node30329 : 4'b0011;
															assign node30329 = (inp[7]) ? node30331 : 4'b0010;
																assign node30331 = (inp[8]) ? 4'b0010 : 4'b0011;
													assign node30334 = (inp[4]) ? node30342 : node30335;
														assign node30335 = (inp[2]) ? node30337 : 4'b0011;
															assign node30337 = (inp[7]) ? 4'b0010 : node30338;
																assign node30338 = (inp[8]) ? 4'b0011 : 4'b0010;
														assign node30342 = (inp[7]) ? 4'b0100 : node30343;
															assign node30343 = (inp[8]) ? node30345 : 4'b0101;
																assign node30345 = (inp[2]) ? 4'b0101 : 4'b0100;
												assign node30349 = (inp[12]) ? node30369 : node30350;
													assign node30350 = (inp[4]) ? node30356 : node30351;
														assign node30351 = (inp[8]) ? 4'b0100 : node30352;
															assign node30352 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node30356 = (inp[8]) ? node30362 : node30357;
															assign node30357 = (inp[7]) ? 4'b0001 : node30358;
																assign node30358 = (inp[2]) ? 4'b0000 : 4'b0001;
															assign node30362 = (inp[2]) ? node30366 : node30363;
																assign node30363 = (inp[7]) ? 4'b0001 : 4'b0000;
																assign node30366 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node30369 = (inp[4]) ? node30377 : node30370;
														assign node30370 = (inp[2]) ? 4'b0001 : node30371;
															assign node30371 = (inp[7]) ? node30373 : 4'b0000;
																assign node30373 = (inp[8]) ? 4'b0001 : 4'b0000;
														assign node30377 = (inp[7]) ? node30379 : 4'b0100;
															assign node30379 = (inp[2]) ? node30383 : node30380;
																assign node30380 = (inp[8]) ? 4'b0101 : 4'b0100;
																assign node30383 = (inp[8]) ? 4'b0100 : 4'b0101;
									assign node30386 = (inp[15]) ? node30540 : node30387;
										assign node30387 = (inp[5]) ? node30465 : node30388;
											assign node30388 = (inp[3]) ? node30432 : node30389;
												assign node30389 = (inp[7]) ? node30409 : node30390;
													assign node30390 = (inp[4]) ? node30398 : node30391;
														assign node30391 = (inp[12]) ? 4'b0101 : node30392;
															assign node30392 = (inp[2]) ? node30394 : 4'b0001;
																assign node30394 = (inp[8]) ? 4'b0001 : 4'b0000;
														assign node30398 = (inp[12]) ? node30404 : node30399;
															assign node30399 = (inp[8]) ? node30401 : 4'b0101;
																assign node30401 = (inp[2]) ? 4'b0101 : 4'b0100;
															assign node30404 = (inp[8]) ? node30406 : 4'b0000;
																assign node30406 = (inp[2]) ? 4'b0001 : 4'b0000;
													assign node30409 = (inp[2]) ? node30423 : node30410;
														assign node30410 = (inp[8]) ? node30416 : node30411;
															assign node30411 = (inp[12]) ? 4'b0100 : node30412;
																assign node30412 = (inp[4]) ? 4'b0100 : 4'b0000;
															assign node30416 = (inp[12]) ? node30420 : node30417;
																assign node30417 = (inp[4]) ? 4'b0101 : 4'b0001;
																assign node30420 = (inp[4]) ? 4'b0001 : 4'b0101;
														assign node30423 = (inp[8]) ? node30425 : 4'b0101;
															assign node30425 = (inp[12]) ? node30429 : node30426;
																assign node30426 = (inp[4]) ? 4'b0100 : 4'b0000;
																assign node30429 = (inp[4]) ? 4'b0000 : 4'b0100;
												assign node30432 = (inp[4]) ? node30446 : node30433;
													assign node30433 = (inp[12]) ? node30441 : node30434;
														assign node30434 = (inp[8]) ? 4'b0001 : node30435;
															assign node30435 = (inp[2]) ? node30437 : 4'b0000;
																assign node30437 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node30441 = (inp[8]) ? node30443 : 4'b0111;
															assign node30443 = (inp[2]) ? 4'b0110 : 4'b0111;
													assign node30446 = (inp[12]) ? node30454 : node30447;
														assign node30447 = (inp[2]) ? node30449 : 4'b0111;
															assign node30449 = (inp[8]) ? node30451 : 4'b0111;
																assign node30451 = (inp[7]) ? 4'b0110 : 4'b0111;
														assign node30454 = (inp[7]) ? node30460 : node30455;
															assign node30455 = (inp[2]) ? 4'b0011 : node30456;
																assign node30456 = (inp[8]) ? 4'b0010 : 4'b0011;
															assign node30460 = (inp[2]) ? 4'b0010 : node30461;
																assign node30461 = (inp[8]) ? 4'b0011 : 4'b0010;
											assign node30465 = (inp[3]) ? node30503 : node30466;
												assign node30466 = (inp[4]) ? node30480 : node30467;
													assign node30467 = (inp[12]) ? node30471 : node30468;
														assign node30468 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node30471 = (inp[2]) ? 4'b0111 : node30472;
															assign node30472 = (inp[8]) ? node30476 : node30473;
																assign node30473 = (inp[7]) ? 4'b0110 : 4'b0111;
																assign node30476 = (inp[7]) ? 4'b0111 : 4'b0110;
													assign node30480 = (inp[12]) ? node30494 : node30481;
														assign node30481 = (inp[2]) ? node30487 : node30482;
															assign node30482 = (inp[7]) ? 4'b0111 : node30483;
																assign node30483 = (inp[8]) ? 4'b0110 : 4'b0111;
															assign node30487 = (inp[7]) ? node30491 : node30488;
																assign node30488 = (inp[8]) ? 4'b0111 : 4'b0110;
																assign node30491 = (inp[8]) ? 4'b0110 : 4'b0111;
														assign node30494 = (inp[2]) ? 4'b0011 : node30495;
															assign node30495 = (inp[7]) ? node30499 : node30496;
																assign node30496 = (inp[8]) ? 4'b0010 : 4'b0011;
																assign node30499 = (inp[8]) ? 4'b0011 : 4'b0010;
												assign node30503 = (inp[8]) ? node30525 : node30504;
													assign node30504 = (inp[4]) ? node30514 : node30505;
														assign node30505 = (inp[12]) ? 4'b0110 : node30506;
															assign node30506 = (inp[2]) ? node30510 : node30507;
																assign node30507 = (inp[7]) ? 4'b0010 : 4'b0011;
																assign node30510 = (inp[7]) ? 4'b0011 : 4'b0010;
														assign node30514 = (inp[12]) ? node30520 : node30515;
															assign node30515 = (inp[2]) ? node30517 : 4'b0110;
																assign node30517 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node30520 = (inp[2]) ? 4'b0010 : node30521;
																assign node30521 = (inp[7]) ? 4'b0010 : 4'b0011;
													assign node30525 = (inp[12]) ? node30535 : node30526;
														assign node30526 = (inp[4]) ? node30530 : node30527;
															assign node30527 = (inp[2]) ? 4'b0011 : 4'b0010;
															assign node30530 = (inp[2]) ? 4'b0111 : node30531;
																assign node30531 = (inp[7]) ? 4'b0111 : 4'b0110;
														assign node30535 = (inp[4]) ? node30537 : 4'b0111;
															assign node30537 = (inp[2]) ? 4'b0010 : 4'b0011;
										assign node30540 = (inp[3]) ? node30610 : node30541;
											assign node30541 = (inp[5]) ? node30573 : node30542;
												assign node30542 = (inp[4]) ? node30558 : node30543;
													assign node30543 = (inp[12]) ? node30551 : node30544;
														assign node30544 = (inp[2]) ? 4'b0011 : node30545;
															assign node30545 = (inp[7]) ? 4'b0010 : node30546;
																assign node30546 = (inp[8]) ? 4'b0010 : 4'b0011;
														assign node30551 = (inp[2]) ? 4'b0110 : node30552;
															assign node30552 = (inp[8]) ? 4'b0111 : node30553;
																assign node30553 = (inp[7]) ? 4'b0110 : 4'b0111;
													assign node30558 = (inp[12]) ? node30566 : node30559;
														assign node30559 = (inp[8]) ? node30561 : 4'b0111;
															assign node30561 = (inp[7]) ? node30563 : 4'b0111;
																assign node30563 = (inp[2]) ? 4'b0110 : 4'b0111;
														assign node30566 = (inp[2]) ? node30568 : 4'b0011;
															assign node30568 = (inp[8]) ? node30570 : 4'b0011;
																assign node30570 = (inp[7]) ? 4'b0010 : 4'b0011;
												assign node30573 = (inp[4]) ? node30591 : node30574;
													assign node30574 = (inp[12]) ? node30584 : node30575;
														assign node30575 = (inp[8]) ? 4'b0011 : node30576;
															assign node30576 = (inp[2]) ? node30580 : node30577;
																assign node30577 = (inp[7]) ? 4'b0010 : 4'b0011;
																assign node30580 = (inp[7]) ? 4'b0011 : 4'b0010;
														assign node30584 = (inp[7]) ? node30586 : 4'b0101;
															assign node30586 = (inp[2]) ? node30588 : 4'b0100;
																assign node30588 = (inp[8]) ? 4'b0100 : 4'b0101;
													assign node30591 = (inp[12]) ? node30603 : node30592;
														assign node30592 = (inp[8]) ? node30598 : node30593;
															assign node30593 = (inp[2]) ? 4'b0100 : node30594;
																assign node30594 = (inp[7]) ? 4'b0100 : 4'b0101;
															assign node30598 = (inp[7]) ? node30600 : 4'b0101;
																assign node30600 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node30603 = (inp[7]) ? node30605 : 4'b0000;
															assign node30605 = (inp[8]) ? node30607 : 4'b0001;
																assign node30607 = (inp[2]) ? 4'b0000 : 4'b0001;
											assign node30610 = (inp[12]) ? node30646 : node30611;
												assign node30611 = (inp[4]) ? node30629 : node30612;
													assign node30612 = (inp[5]) ? node30622 : node30613;
														assign node30613 = (inp[2]) ? node30615 : 4'b0011;
															assign node30615 = (inp[7]) ? node30619 : node30616;
																assign node30616 = (inp[8]) ? 4'b0011 : 4'b0010;
																assign node30619 = (inp[8]) ? 4'b0010 : 4'b0011;
														assign node30622 = (inp[2]) ? node30624 : 4'b0000;
															assign node30624 = (inp[7]) ? node30626 : 4'b0001;
																assign node30626 = (inp[8]) ? 4'b0000 : 4'b0001;
													assign node30629 = (inp[8]) ? node30639 : node30630;
														assign node30630 = (inp[5]) ? node30636 : node30631;
															assign node30631 = (inp[7]) ? node30633 : 4'b0100;
																assign node30633 = (inp[2]) ? 4'b0101 : 4'b0100;
															assign node30636 = (inp[7]) ? 4'b0100 : 4'b0101;
														assign node30639 = (inp[7]) ? node30643 : node30640;
															assign node30640 = (inp[2]) ? 4'b0101 : 4'b0100;
															assign node30643 = (inp[2]) ? 4'b0100 : 4'b0101;
												assign node30646 = (inp[4]) ? node30672 : node30647;
													assign node30647 = (inp[5]) ? node30663 : node30648;
														assign node30648 = (inp[8]) ? node30656 : node30649;
															assign node30649 = (inp[7]) ? node30653 : node30650;
																assign node30650 = (inp[2]) ? 4'b0100 : 4'b0101;
																assign node30653 = (inp[2]) ? 4'b0101 : 4'b0100;
															assign node30656 = (inp[7]) ? node30660 : node30657;
																assign node30657 = (inp[2]) ? 4'b0101 : 4'b0100;
																assign node30660 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node30663 = (inp[8]) ? 4'b0101 : node30664;
															assign node30664 = (inp[2]) ? node30668 : node30665;
																assign node30665 = (inp[7]) ? 4'b0100 : 4'b0101;
																assign node30668 = (inp[7]) ? 4'b0101 : 4'b0100;
													assign node30672 = (inp[2]) ? node30682 : node30673;
														assign node30673 = (inp[5]) ? 4'b0000 : node30674;
															assign node30674 = (inp[8]) ? node30678 : node30675;
																assign node30675 = (inp[7]) ? 4'b0000 : 4'b0001;
																assign node30678 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node30682 = (inp[7]) ? 4'b0001 : node30683;
															assign node30683 = (inp[5]) ? 4'b0001 : 4'b0000;
								assign node30687 = (inp[5]) ? node30917 : node30688;
									assign node30688 = (inp[15]) ? node30806 : node30689;
										assign node30689 = (inp[3]) ? node30763 : node30690;
											assign node30690 = (inp[12]) ? node30728 : node30691;
												assign node30691 = (inp[2]) ? node30713 : node30692;
													assign node30692 = (inp[9]) ? node30704 : node30693;
														assign node30693 = (inp[4]) ? node30699 : node30694;
															assign node30694 = (inp[7]) ? 4'b0100 : node30695;
																assign node30695 = (inp[8]) ? 4'b0101 : 4'b0100;
															assign node30699 = (inp[7]) ? node30701 : 4'b0001;
																assign node30701 = (inp[8]) ? 4'b0000 : 4'b0001;
														assign node30704 = (inp[4]) ? node30706 : 4'b0001;
															assign node30706 = (inp[7]) ? node30710 : node30707;
																assign node30707 = (inp[8]) ? 4'b0101 : 4'b0100;
																assign node30710 = (inp[8]) ? 4'b0100 : 4'b0101;
													assign node30713 = (inp[4]) ? node30717 : node30714;
														assign node30714 = (inp[9]) ? 4'b0001 : 4'b0101;
														assign node30717 = (inp[9]) ? node30723 : node30718;
															assign node30718 = (inp[7]) ? 4'b0001 : node30719;
																assign node30719 = (inp[8]) ? 4'b0001 : 4'b0000;
															assign node30723 = (inp[7]) ? node30725 : 4'b0101;
																assign node30725 = (inp[8]) ? 4'b0100 : 4'b0101;
												assign node30728 = (inp[4]) ? node30740 : node30729;
													assign node30729 = (inp[9]) ? node30735 : node30730;
														assign node30730 = (inp[7]) ? 4'b0000 : node30731;
															assign node30731 = (inp[8]) ? 4'b0001 : 4'b0000;
														assign node30735 = (inp[8]) ? node30737 : 4'b0100;
															assign node30737 = (inp[7]) ? 4'b0100 : 4'b0101;
													assign node30740 = (inp[9]) ? node30756 : node30741;
														assign node30741 = (inp[2]) ? node30749 : node30742;
															assign node30742 = (inp[7]) ? node30746 : node30743;
																assign node30743 = (inp[8]) ? 4'b0101 : 4'b0100;
																assign node30746 = (inp[8]) ? 4'b0100 : 4'b0101;
															assign node30749 = (inp[7]) ? node30753 : node30750;
																assign node30750 = (inp[8]) ? 4'b0101 : 4'b0100;
																assign node30753 = (inp[8]) ? 4'b0100 : 4'b0101;
														assign node30756 = (inp[7]) ? node30760 : node30757;
															assign node30757 = (inp[8]) ? 4'b0001 : 4'b0000;
															assign node30760 = (inp[8]) ? 4'b0000 : 4'b0001;
											assign node30763 = (inp[12]) ? node30789 : node30764;
												assign node30764 = (inp[9]) ? node30780 : node30765;
													assign node30765 = (inp[4]) ? node30771 : node30766;
														assign node30766 = (inp[7]) ? node30768 : 4'b0101;
															assign node30768 = (inp[8]) ? 4'b0100 : 4'b0101;
														assign node30771 = (inp[2]) ? 4'b0001 : node30772;
															assign node30772 = (inp[7]) ? node30776 : node30773;
																assign node30773 = (inp[8]) ? 4'b0001 : 4'b0000;
																assign node30776 = (inp[8]) ? 4'b0000 : 4'b0001;
													assign node30780 = (inp[4]) ? node30784 : node30781;
														assign node30781 = (inp[8]) ? 4'b0000 : 4'b0001;
														assign node30784 = (inp[7]) ? 4'b0110 : node30785;
															assign node30785 = (inp[8]) ? 4'b0111 : 4'b0110;
												assign node30789 = (inp[8]) ? node30801 : node30790;
													assign node30790 = (inp[7]) ? node30794 : node30791;
														assign node30791 = (inp[9]) ? 4'b0010 : 4'b0000;
														assign node30794 = (inp[4]) ? node30798 : node30795;
															assign node30795 = (inp[9]) ? 4'b0111 : 4'b0001;
															assign node30798 = (inp[9]) ? 4'b0011 : 4'b0111;
													assign node30801 = (inp[7]) ? node30803 : 4'b0111;
														assign node30803 = (inp[9]) ? 4'b0010 : 4'b0110;
										assign node30806 = (inp[3]) ? node30862 : node30807;
											assign node30807 = (inp[12]) ? node30829 : node30808;
												assign node30808 = (inp[4]) ? node30816 : node30809;
													assign node30809 = (inp[9]) ? 4'b0010 : node30810;
														assign node30810 = (inp[7]) ? 4'b0110 : node30811;
															assign node30811 = (inp[8]) ? 4'b0111 : 4'b0110;
													assign node30816 = (inp[9]) ? node30822 : node30817;
														assign node30817 = (inp[8]) ? node30819 : 4'b0010;
															assign node30819 = (inp[7]) ? 4'b0010 : 4'b0011;
														assign node30822 = (inp[8]) ? node30826 : node30823;
															assign node30823 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node30826 = (inp[2]) ? 4'b0111 : 4'b0110;
												assign node30829 = (inp[9]) ? node30851 : node30830;
													assign node30830 = (inp[4]) ? node30838 : node30831;
														assign node30831 = (inp[2]) ? 4'b0011 : node30832;
															assign node30832 = (inp[7]) ? node30834 : 4'b0010;
																assign node30834 = (inp[8]) ? 4'b0010 : 4'b0011;
														assign node30838 = (inp[2]) ? node30844 : node30839;
															assign node30839 = (inp[7]) ? node30841 : 4'b0110;
																assign node30841 = (inp[8]) ? 4'b0110 : 4'b0111;
															assign node30844 = (inp[8]) ? node30848 : node30845;
																assign node30845 = (inp[7]) ? 4'b0111 : 4'b0110;
																assign node30848 = (inp[7]) ? 4'b0110 : 4'b0111;
													assign node30851 = (inp[4]) ? node30855 : node30852;
														assign node30852 = (inp[2]) ? 4'b0110 : 4'b0111;
														assign node30855 = (inp[8]) ? node30859 : node30856;
															assign node30856 = (inp[7]) ? 4'b0011 : 4'b0010;
															assign node30859 = (inp[7]) ? 4'b0010 : 4'b0011;
											assign node30862 = (inp[9]) ? node30890 : node30863;
												assign node30863 = (inp[12]) ? node30877 : node30864;
													assign node30864 = (inp[4]) ? node30870 : node30865;
														assign node30865 = (inp[7]) ? node30867 : 4'b0111;
															assign node30867 = (inp[8]) ? 4'b0110 : 4'b0111;
														assign node30870 = (inp[7]) ? node30874 : node30871;
															assign node30871 = (inp[8]) ? 4'b0011 : 4'b0010;
															assign node30874 = (inp[8]) ? 4'b0010 : 4'b0011;
													assign node30877 = (inp[4]) ? node30885 : node30878;
														assign node30878 = (inp[7]) ? node30882 : node30879;
															assign node30879 = (inp[8]) ? 4'b0011 : 4'b0010;
															assign node30882 = (inp[8]) ? 4'b0010 : 4'b0011;
														assign node30885 = (inp[8]) ? node30887 : 4'b0101;
															assign node30887 = (inp[7]) ? 4'b0100 : 4'b0101;
												assign node30890 = (inp[12]) ? node30902 : node30891;
													assign node30891 = (inp[4]) ? node30897 : node30892;
														assign node30892 = (inp[8]) ? 4'b0010 : node30893;
															assign node30893 = (inp[7]) ? 4'b0011 : 4'b0010;
														assign node30897 = (inp[7]) ? node30899 : 4'b0100;
															assign node30899 = (inp[8]) ? 4'b0100 : 4'b0101;
													assign node30902 = (inp[4]) ? node30910 : node30903;
														assign node30903 = (inp[2]) ? node30905 : 4'b0101;
															assign node30905 = (inp[8]) ? node30907 : 4'b0101;
																assign node30907 = (inp[7]) ? 4'b0100 : 4'b0101;
														assign node30910 = (inp[2]) ? 4'b0000 : node30911;
															assign node30911 = (inp[7]) ? 4'b0001 : node30912;
																assign node30912 = (inp[8]) ? 4'b0001 : 4'b0000;
									assign node30917 = (inp[15]) ? node31051 : node30918;
										assign node30918 = (inp[3]) ? node30988 : node30919;
											assign node30919 = (inp[12]) ? node30953 : node30920;
												assign node30920 = (inp[9]) ? node30942 : node30921;
													assign node30921 = (inp[4]) ? node30929 : node30922;
														assign node30922 = (inp[7]) ? node30926 : node30923;
															assign node30923 = (inp[8]) ? 4'b0101 : 4'b0100;
															assign node30926 = (inp[8]) ? 4'b0100 : 4'b0101;
														assign node30929 = (inp[2]) ? node30935 : node30930;
															assign node30930 = (inp[7]) ? node30932 : 4'b0000;
																assign node30932 = (inp[8]) ? 4'b0000 : 4'b0001;
															assign node30935 = (inp[8]) ? node30939 : node30936;
																assign node30936 = (inp[7]) ? 4'b0001 : 4'b0000;
																assign node30939 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node30942 = (inp[4]) ? node30950 : node30943;
														assign node30943 = (inp[8]) ? node30947 : node30944;
															assign node30944 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node30947 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node30950 = (inp[2]) ? 4'b0111 : 4'b0110;
												assign node30953 = (inp[9]) ? node30969 : node30954;
													assign node30954 = (inp[4]) ? node30962 : node30955;
														assign node30955 = (inp[7]) ? node30959 : node30956;
															assign node30956 = (inp[8]) ? 4'b0001 : 4'b0000;
															assign node30959 = (inp[8]) ? 4'b0000 : 4'b0001;
														assign node30962 = (inp[2]) ? node30964 : 4'b0110;
															assign node30964 = (inp[7]) ? 4'b0111 : node30965;
																assign node30965 = (inp[8]) ? 4'b0111 : 4'b0110;
													assign node30969 = (inp[4]) ? node30983 : node30970;
														assign node30970 = (inp[2]) ? node30978 : node30971;
															assign node30971 = (inp[8]) ? node30975 : node30972;
																assign node30972 = (inp[7]) ? 4'b0111 : 4'b0110;
																assign node30975 = (inp[7]) ? 4'b0110 : 4'b0111;
															assign node30978 = (inp[7]) ? 4'b0111 : node30979;
																assign node30979 = (inp[8]) ? 4'b0111 : 4'b0110;
														assign node30983 = (inp[8]) ? node30985 : 4'b0011;
															assign node30985 = (inp[7]) ? 4'b0010 : 4'b0011;
											assign node30988 = (inp[9]) ? node31032 : node30989;
												assign node30989 = (inp[4]) ? node31005 : node30990;
													assign node30990 = (inp[12]) ? node30998 : node30991;
														assign node30991 = (inp[8]) ? node30995 : node30992;
															assign node30992 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node30995 = (inp[7]) ? 4'b0110 : 4'b0111;
														assign node30998 = (inp[7]) ? node31002 : node30999;
															assign node30999 = (inp[8]) ? 4'b0011 : 4'b0010;
															assign node31002 = (inp[8]) ? 4'b0010 : 4'b0011;
													assign node31005 = (inp[12]) ? node31021 : node31006;
														assign node31006 = (inp[2]) ? node31014 : node31007;
															assign node31007 = (inp[7]) ? node31011 : node31008;
																assign node31008 = (inp[8]) ? 4'b0011 : 4'b0010;
																assign node31011 = (inp[8]) ? 4'b0010 : 4'b0011;
															assign node31014 = (inp[8]) ? node31018 : node31015;
																assign node31015 = (inp[7]) ? 4'b0011 : 4'b0010;
																assign node31018 = (inp[7]) ? 4'b0010 : 4'b0011;
														assign node31021 = (inp[2]) ? node31027 : node31022;
															assign node31022 = (inp[7]) ? node31024 : 4'b0111;
																assign node31024 = (inp[8]) ? 4'b0110 : 4'b0111;
															assign node31027 = (inp[7]) ? 4'b0110 : node31028;
																assign node31028 = (inp[8]) ? 4'b0111 : 4'b0110;
												assign node31032 = (inp[12]) ? node31036 : node31033;
													assign node31033 = (inp[4]) ? 4'b0110 : 4'b0010;
													assign node31036 = (inp[4]) ? node31048 : node31037;
														assign node31037 = (inp[2]) ? node31043 : node31038;
															assign node31038 = (inp[7]) ? 4'b0111 : node31039;
																assign node31039 = (inp[8]) ? 4'b0111 : 4'b0110;
															assign node31043 = (inp[8]) ? node31045 : 4'b0110;
																assign node31045 = (inp[7]) ? 4'b0110 : 4'b0111;
														assign node31048 = (inp[7]) ? 4'b0010 : 4'b0011;
										assign node31051 = (inp[3]) ? node31129 : node31052;
											assign node31052 = (inp[12]) ? node31092 : node31053;
												assign node31053 = (inp[4]) ? node31077 : node31054;
													assign node31054 = (inp[9]) ? node31068 : node31055;
														assign node31055 = (inp[2]) ? node31063 : node31056;
															assign node31056 = (inp[8]) ? node31060 : node31057;
																assign node31057 = (inp[7]) ? 4'b0111 : 4'b0110;
																assign node31060 = (inp[7]) ? 4'b0110 : 4'b0111;
															assign node31063 = (inp[8]) ? node31065 : 4'b0110;
																assign node31065 = (inp[7]) ? 4'b0110 : 4'b0111;
														assign node31068 = (inp[2]) ? node31070 : 4'b0010;
															assign node31070 = (inp[8]) ? node31074 : node31071;
																assign node31071 = (inp[7]) ? 4'b0011 : 4'b0010;
																assign node31074 = (inp[7]) ? 4'b0010 : 4'b0011;
													assign node31077 = (inp[9]) ? node31083 : node31078;
														assign node31078 = (inp[7]) ? node31080 : 4'b0011;
															assign node31080 = (inp[8]) ? 4'b0010 : 4'b0011;
														assign node31083 = (inp[2]) ? node31085 : 4'b0100;
															assign node31085 = (inp[8]) ? node31089 : node31086;
																assign node31086 = (inp[7]) ? 4'b0101 : 4'b0100;
																assign node31089 = (inp[7]) ? 4'b0100 : 4'b0101;
												assign node31092 = (inp[4]) ? node31110 : node31093;
													assign node31093 = (inp[9]) ? node31099 : node31094;
														assign node31094 = (inp[8]) ? 4'b0010 : node31095;
															assign node31095 = (inp[7]) ? 4'b0011 : 4'b0010;
														assign node31099 = (inp[2]) ? node31105 : node31100;
															assign node31100 = (inp[8]) ? node31102 : 4'b0100;
																assign node31102 = (inp[7]) ? 4'b0100 : 4'b0101;
															assign node31105 = (inp[8]) ? node31107 : 4'b0101;
																assign node31107 = (inp[7]) ? 4'b0100 : 4'b0101;
													assign node31110 = (inp[9]) ? node31118 : node31111;
														assign node31111 = (inp[7]) ? node31115 : node31112;
															assign node31112 = (inp[8]) ? 4'b0101 : 4'b0100;
															assign node31115 = (inp[8]) ? 4'b0100 : 4'b0101;
														assign node31118 = (inp[2]) ? node31124 : node31119;
															assign node31119 = (inp[8]) ? node31121 : 4'b0001;
																assign node31121 = (inp[7]) ? 4'b0000 : 4'b0001;
															assign node31124 = (inp[8]) ? node31126 : 4'b0000;
																assign node31126 = (inp[7]) ? 4'b0000 : 4'b0001;
											assign node31129 = (inp[9]) ? node31165 : node31130;
												assign node31130 = (inp[8]) ? node31144 : node31131;
													assign node31131 = (inp[7]) ? node31137 : node31132;
														assign node31132 = (inp[4]) ? node31134 : 4'b0000;
															assign node31134 = (inp[12]) ? 4'b0100 : 4'b0000;
														assign node31137 = (inp[4]) ? node31141 : node31138;
															assign node31138 = (inp[2]) ? 4'b0101 : 4'b0001;
															assign node31141 = (inp[2]) ? 4'b0001 : 4'b0101;
													assign node31144 = (inp[7]) ? node31152 : node31145;
														assign node31145 = (inp[2]) ? 4'b0101 : node31146;
															assign node31146 = (inp[12]) ? 4'b0001 : node31147;
																assign node31147 = (inp[4]) ? 4'b0001 : 4'b0101;
														assign node31152 = (inp[2]) ? node31160 : node31153;
															assign node31153 = (inp[12]) ? node31157 : node31154;
																assign node31154 = (inp[4]) ? 4'b0000 : 4'b0100;
																assign node31157 = (inp[4]) ? 4'b0100 : 4'b0000;
															assign node31160 = (inp[12]) ? 4'b0000 : node31161;
																assign node31161 = (inp[4]) ? 4'b0000 : 4'b0100;
												assign node31165 = (inp[8]) ? node31179 : node31166;
													assign node31166 = (inp[7]) ? node31172 : node31167;
														assign node31167 = (inp[4]) ? 4'b0100 : node31168;
															assign node31168 = (inp[12]) ? 4'b0100 : 4'b0000;
														assign node31172 = (inp[12]) ? node31176 : node31173;
															assign node31173 = (inp[4]) ? 4'b0101 : 4'b0001;
															assign node31176 = (inp[4]) ? 4'b0001 : 4'b0101;
													assign node31179 = (inp[7]) ? node31187 : node31180;
														assign node31180 = (inp[12]) ? node31184 : node31181;
															assign node31181 = (inp[4]) ? 4'b0101 : 4'b0001;
															assign node31184 = (inp[2]) ? 4'b0001 : 4'b0101;
														assign node31187 = (inp[12]) ? node31189 : 4'b0100;
															assign node31189 = (inp[4]) ? 4'b0000 : 4'b0100;
		assign node31192 = (inp[11]) ? node47420 : node31193;
			assign node31193 = (inp[6]) ? node40135 : node31194;
				assign node31194 = (inp[1]) ? node35644 : node31195;
					assign node31195 = (inp[13]) ? node33403 : node31196;
						assign node31196 = (inp[2]) ? node32442 : node31197;
							assign node31197 = (inp[15]) ? node31815 : node31198;
								assign node31198 = (inp[5]) ? node31508 : node31199;
									assign node31199 = (inp[0]) ? node31373 : node31200;
										assign node31200 = (inp[3]) ? node31284 : node31201;
											assign node31201 = (inp[8]) ? node31241 : node31202;
												assign node31202 = (inp[9]) ? node31224 : node31203;
													assign node31203 = (inp[14]) ? node31213 : node31204;
														assign node31204 = (inp[7]) ? node31206 : 4'b1111;
															assign node31206 = (inp[4]) ? node31210 : node31207;
																assign node31207 = (inp[12]) ? 4'b1010 : 4'b1110;
																assign node31210 = (inp[12]) ? 4'b1110 : 4'b1010;
														assign node31213 = (inp[7]) ? node31217 : node31214;
															assign node31214 = (inp[4]) ? 4'b1110 : 4'b1010;
															assign node31217 = (inp[12]) ? node31221 : node31218;
																assign node31218 = (inp[4]) ? 4'b1011 : 4'b1111;
																assign node31221 = (inp[4]) ? 4'b1111 : 4'b1011;
													assign node31224 = (inp[7]) ? node31232 : node31225;
														assign node31225 = (inp[14]) ? node31227 : 4'b1011;
															assign node31227 = (inp[4]) ? node31229 : 4'b1110;
																assign node31229 = (inp[12]) ? 4'b1010 : 4'b1110;
														assign node31232 = (inp[14]) ? 4'b1011 : node31233;
															assign node31233 = (inp[12]) ? node31237 : node31234;
																assign node31234 = (inp[4]) ? 4'b1110 : 4'b1010;
																assign node31237 = (inp[4]) ? 4'b1010 : 4'b1110;
												assign node31241 = (inp[7]) ? node31265 : node31242;
													assign node31242 = (inp[14]) ? node31252 : node31243;
														assign node31243 = (inp[12]) ? 4'b1110 : node31244;
															assign node31244 = (inp[9]) ? node31248 : node31245;
																assign node31245 = (inp[4]) ? 4'b1010 : 4'b1110;
																assign node31248 = (inp[4]) ? 4'b1110 : 4'b1010;
														assign node31252 = (inp[4]) ? node31258 : node31253;
															assign node31253 = (inp[9]) ? node31255 : 4'b1111;
																assign node31255 = (inp[12]) ? 4'b1111 : 4'b1011;
															assign node31258 = (inp[12]) ? node31262 : node31259;
																assign node31259 = (inp[9]) ? 4'b1111 : 4'b1011;
																assign node31262 = (inp[9]) ? 4'b1011 : 4'b1111;
													assign node31265 = (inp[14]) ? node31279 : node31266;
														assign node31266 = (inp[12]) ? node31272 : node31267;
															assign node31267 = (inp[9]) ? node31269 : 4'b1111;
																assign node31269 = (inp[4]) ? 4'b1111 : 4'b1011;
															assign node31272 = (inp[9]) ? node31276 : node31273;
																assign node31273 = (inp[4]) ? 4'b1111 : 4'b1011;
																assign node31276 = (inp[4]) ? 4'b1011 : 4'b1111;
														assign node31279 = (inp[9]) ? 4'b1110 : node31280;
															assign node31280 = (inp[12]) ? 4'b1010 : 4'b1110;
											assign node31284 = (inp[4]) ? node31326 : node31285;
												assign node31285 = (inp[12]) ? node31311 : node31286;
													assign node31286 = (inp[9]) ? node31298 : node31287;
														assign node31287 = (inp[7]) ? node31293 : node31288;
															assign node31288 = (inp[8]) ? 4'b1111 : node31289;
																assign node31289 = (inp[14]) ? 4'b1110 : 4'b1111;
															assign node31293 = (inp[8]) ? 4'b1110 : node31294;
																assign node31294 = (inp[14]) ? 4'b1111 : 4'b1110;
														assign node31298 = (inp[7]) ? node31306 : node31299;
															assign node31299 = (inp[8]) ? node31303 : node31300;
																assign node31300 = (inp[14]) ? 4'b1010 : 4'b1011;
																assign node31303 = (inp[14]) ? 4'b1011 : 4'b1010;
															assign node31306 = (inp[8]) ? 4'b1010 : node31307;
																assign node31307 = (inp[14]) ? 4'b1011 : 4'b1010;
													assign node31311 = (inp[9]) ? node31319 : node31312;
														assign node31312 = (inp[14]) ? node31314 : 4'b1010;
															assign node31314 = (inp[7]) ? node31316 : 4'b1011;
																assign node31316 = (inp[8]) ? 4'b1010 : 4'b1011;
														assign node31319 = (inp[14]) ? 4'b1101 : node31320;
															assign node31320 = (inp[7]) ? node31322 : 4'b1100;
																assign node31322 = (inp[8]) ? 4'b1101 : 4'b1100;
												assign node31326 = (inp[9]) ? node31348 : node31327;
													assign node31327 = (inp[12]) ? node31341 : node31328;
														assign node31328 = (inp[8]) ? node31336 : node31329;
															assign node31329 = (inp[14]) ? node31333 : node31330;
																assign node31330 = (inp[7]) ? 4'b1010 : 4'b1011;
																assign node31333 = (inp[7]) ? 4'b1011 : 4'b1010;
															assign node31336 = (inp[14]) ? node31338 : 4'b1010;
																assign node31338 = (inp[7]) ? 4'b1010 : 4'b1011;
														assign node31341 = (inp[8]) ? node31343 : 4'b1100;
															assign node31343 = (inp[14]) ? node31345 : 4'b1101;
																assign node31345 = (inp[7]) ? 4'b1100 : 4'b1101;
													assign node31348 = (inp[12]) ? node31362 : node31349;
														assign node31349 = (inp[7]) ? node31357 : node31350;
															assign node31350 = (inp[14]) ? node31354 : node31351;
																assign node31351 = (inp[8]) ? 4'b1100 : 4'b1101;
																assign node31354 = (inp[8]) ? 4'b1101 : 4'b1100;
															assign node31357 = (inp[14]) ? node31359 : 4'b1100;
																assign node31359 = (inp[8]) ? 4'b1100 : 4'b1101;
														assign node31362 = (inp[7]) ? node31368 : node31363;
															assign node31363 = (inp[14]) ? node31365 : 4'b1001;
																assign node31365 = (inp[8]) ? 4'b1001 : 4'b1000;
															assign node31368 = (inp[14]) ? 4'b1000 : node31369;
																assign node31369 = (inp[8]) ? 4'b1001 : 4'b1000;
										assign node31373 = (inp[3]) ? node31437 : node31374;
											assign node31374 = (inp[12]) ? node31406 : node31375;
												assign node31375 = (inp[7]) ? node31391 : node31376;
													assign node31376 = (inp[4]) ? node31384 : node31377;
														assign node31377 = (inp[9]) ? node31379 : 4'b1100;
															assign node31379 = (inp[8]) ? 4'b1001 : node31380;
																assign node31380 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node31384 = (inp[9]) ? node31386 : 4'b1000;
															assign node31386 = (inp[14]) ? node31388 : 4'b1100;
																assign node31388 = (inp[8]) ? 4'b1101 : 4'b1100;
													assign node31391 = (inp[4]) ? node31399 : node31392;
														assign node31392 = (inp[14]) ? node31396 : node31393;
															assign node31393 = (inp[8]) ? 4'b1101 : 4'b1100;
															assign node31396 = (inp[8]) ? 4'b1100 : 4'b1101;
														assign node31399 = (inp[9]) ? node31401 : 4'b1000;
															assign node31401 = (inp[14]) ? 4'b1100 : node31402;
																assign node31402 = (inp[8]) ? 4'b1101 : 4'b1100;
												assign node31406 = (inp[14]) ? node31422 : node31407;
													assign node31407 = (inp[4]) ? node31419 : node31408;
														assign node31408 = (inp[9]) ? node31414 : node31409;
															assign node31409 = (inp[8]) ? node31411 : 4'b1001;
																assign node31411 = (inp[7]) ? 4'b1001 : 4'b1000;
															assign node31414 = (inp[7]) ? node31416 : 4'b1101;
																assign node31416 = (inp[8]) ? 4'b1101 : 4'b1100;
														assign node31419 = (inp[9]) ? 4'b1001 : 4'b1101;
													assign node31422 = (inp[4]) ? node31428 : node31423;
														assign node31423 = (inp[7]) ? 4'b1101 : node31424;
															assign node31424 = (inp[8]) ? 4'b1101 : 4'b1100;
														assign node31428 = (inp[9]) ? node31432 : node31429;
															assign node31429 = (inp[7]) ? 4'b1100 : 4'b1101;
															assign node31432 = (inp[8]) ? node31434 : 4'b1000;
																assign node31434 = (inp[7]) ? 4'b1000 : 4'b1001;
											assign node31437 = (inp[9]) ? node31467 : node31438;
												assign node31438 = (inp[4]) ? node31458 : node31439;
													assign node31439 = (inp[12]) ? node31449 : node31440;
														assign node31440 = (inp[7]) ? node31442 : 4'b1101;
															assign node31442 = (inp[14]) ? node31446 : node31443;
																assign node31443 = (inp[8]) ? 4'b1101 : 4'b1100;
																assign node31446 = (inp[8]) ? 4'b1100 : 4'b1101;
														assign node31449 = (inp[8]) ? node31451 : 4'b1000;
															assign node31451 = (inp[7]) ? node31455 : node31452;
																assign node31452 = (inp[14]) ? 4'b1001 : 4'b1000;
																assign node31455 = (inp[14]) ? 4'b1000 : 4'b1001;
													assign node31458 = (inp[12]) ? node31460 : 4'b1000;
														assign node31460 = (inp[14]) ? node31462 : 4'b1111;
															assign node31462 = (inp[8]) ? node31464 : 4'b1110;
																assign node31464 = (inp[7]) ? 4'b1110 : 4'b1111;
												assign node31467 = (inp[4]) ? node31487 : node31468;
													assign node31468 = (inp[12]) ? node31476 : node31469;
														assign node31469 = (inp[14]) ? 4'b1001 : node31470;
															assign node31470 = (inp[8]) ? node31472 : 4'b1001;
																assign node31472 = (inp[7]) ? 4'b1001 : 4'b1000;
														assign node31476 = (inp[7]) ? node31482 : node31477;
															assign node31477 = (inp[14]) ? 4'b1110 : node31478;
																assign node31478 = (inp[8]) ? 4'b1110 : 4'b1111;
															assign node31482 = (inp[14]) ? 4'b1111 : node31483;
																assign node31483 = (inp[8]) ? 4'b1111 : 4'b1110;
													assign node31487 = (inp[12]) ? node31501 : node31488;
														assign node31488 = (inp[7]) ? node31494 : node31489;
															assign node31489 = (inp[14]) ? node31491 : 4'b1111;
																assign node31491 = (inp[8]) ? 4'b1111 : 4'b1110;
															assign node31494 = (inp[8]) ? node31498 : node31495;
																assign node31495 = (inp[14]) ? 4'b1111 : 4'b1110;
																assign node31498 = (inp[14]) ? 4'b1110 : 4'b1111;
														assign node31501 = (inp[8]) ? 4'b1011 : node31502;
															assign node31502 = (inp[7]) ? node31504 : 4'b1010;
																assign node31504 = (inp[14]) ? 4'b1011 : 4'b1010;
									assign node31508 = (inp[0]) ? node31656 : node31509;
										assign node31509 = (inp[3]) ? node31577 : node31510;
											assign node31510 = (inp[9]) ? node31548 : node31511;
												assign node31511 = (inp[4]) ? node31531 : node31512;
													assign node31512 = (inp[12]) ? node31520 : node31513;
														assign node31513 = (inp[7]) ? 4'b1110 : node31514;
															assign node31514 = (inp[8]) ? node31516 : 4'b1110;
																assign node31516 = (inp[14]) ? 4'b1111 : 4'b1110;
														assign node31520 = (inp[8]) ? node31526 : node31521;
															assign node31521 = (inp[7]) ? node31523 : 4'b1011;
																assign node31523 = (inp[14]) ? 4'b1011 : 4'b1010;
															assign node31526 = (inp[14]) ? node31528 : 4'b1010;
																assign node31528 = (inp[7]) ? 4'b1010 : 4'b1011;
													assign node31531 = (inp[12]) ? node31545 : node31532;
														assign node31532 = (inp[14]) ? node31538 : node31533;
															assign node31533 = (inp[8]) ? node31535 : 4'b1011;
																assign node31535 = (inp[7]) ? 4'b1011 : 4'b1010;
															assign node31538 = (inp[8]) ? node31542 : node31539;
																assign node31539 = (inp[7]) ? 4'b1011 : 4'b1010;
																assign node31542 = (inp[7]) ? 4'b1010 : 4'b1011;
														assign node31545 = (inp[14]) ? 4'b1101 : 4'b1100;
												assign node31548 = (inp[4]) ? node31564 : node31549;
													assign node31549 = (inp[12]) ? node31553 : node31550;
														assign node31550 = (inp[8]) ? 4'b1010 : 4'b1011;
														assign node31553 = (inp[8]) ? node31559 : node31554;
															assign node31554 = (inp[7]) ? node31556 : 4'b1101;
																assign node31556 = (inp[14]) ? 4'b1101 : 4'b1100;
															assign node31559 = (inp[14]) ? 4'b1100 : node31560;
																assign node31560 = (inp[7]) ? 4'b1101 : 4'b1100;
													assign node31564 = (inp[12]) ? node31572 : node31565;
														assign node31565 = (inp[7]) ? 4'b1100 : node31566;
															assign node31566 = (inp[8]) ? 4'b1100 : node31567;
																assign node31567 = (inp[14]) ? 4'b1100 : 4'b1101;
														assign node31572 = (inp[14]) ? node31574 : 4'b1000;
															assign node31574 = (inp[7]) ? 4'b1001 : 4'b1000;
											assign node31577 = (inp[7]) ? node31611 : node31578;
												assign node31578 = (inp[9]) ? node31604 : node31579;
													assign node31579 = (inp[8]) ? node31593 : node31580;
														assign node31580 = (inp[14]) ? node31588 : node31581;
															assign node31581 = (inp[4]) ? node31585 : node31582;
																assign node31582 = (inp[12]) ? 4'b1001 : 4'b1101;
																assign node31585 = (inp[12]) ? 4'b1101 : 4'b1001;
															assign node31588 = (inp[4]) ? node31590 : 4'b1100;
																assign node31590 = (inp[12]) ? 4'b1100 : 4'b1000;
														assign node31593 = (inp[14]) ? node31599 : node31594;
															assign node31594 = (inp[12]) ? node31596 : 4'b1000;
																assign node31596 = (inp[4]) ? 4'b1100 : 4'b1000;
															assign node31599 = (inp[12]) ? 4'b1001 : node31600;
																assign node31600 = (inp[4]) ? 4'b1001 : 4'b1101;
													assign node31604 = (inp[14]) ? 4'b1101 : node31605;
														assign node31605 = (inp[8]) ? 4'b1000 : node31606;
															assign node31606 = (inp[12]) ? 4'b1001 : 4'b1101;
												assign node31611 = (inp[9]) ? node31635 : node31612;
													assign node31612 = (inp[8]) ? node31626 : node31613;
														assign node31613 = (inp[14]) ? node31621 : node31614;
															assign node31614 = (inp[4]) ? node31618 : node31615;
																assign node31615 = (inp[12]) ? 4'b1000 : 4'b1100;
																assign node31618 = (inp[12]) ? 4'b1100 : 4'b1000;
															assign node31621 = (inp[4]) ? 4'b1101 : node31622;
																assign node31622 = (inp[12]) ? 4'b1001 : 4'b1101;
														assign node31626 = (inp[14]) ? node31628 : 4'b1101;
															assign node31628 = (inp[12]) ? node31632 : node31629;
																assign node31629 = (inp[4]) ? 4'b1000 : 4'b1100;
																assign node31632 = (inp[4]) ? 4'b1100 : 4'b1000;
													assign node31635 = (inp[8]) ? node31643 : node31636;
														assign node31636 = (inp[14]) ? 4'b1001 : node31637;
															assign node31637 = (inp[4]) ? 4'b1000 : node31638;
																assign node31638 = (inp[12]) ? 4'b1100 : 4'b1000;
														assign node31643 = (inp[14]) ? node31651 : node31644;
															assign node31644 = (inp[4]) ? node31648 : node31645;
																assign node31645 = (inp[12]) ? 4'b1101 : 4'b1001;
																assign node31648 = (inp[12]) ? 4'b1001 : 4'b1101;
															assign node31651 = (inp[12]) ? 4'b1100 : node31652;
																assign node31652 = (inp[4]) ? 4'b1100 : 4'b1000;
										assign node31656 = (inp[3]) ? node31722 : node31657;
											assign node31657 = (inp[4]) ? node31685 : node31658;
												assign node31658 = (inp[9]) ? node31674 : node31659;
													assign node31659 = (inp[12]) ? node31663 : node31660;
														assign node31660 = (inp[8]) ? 4'b1101 : 4'b1100;
														assign node31663 = (inp[8]) ? node31669 : node31664;
															assign node31664 = (inp[14]) ? node31666 : 4'b1001;
																assign node31666 = (inp[7]) ? 4'b1001 : 4'b1000;
															assign node31669 = (inp[7]) ? 4'b1000 : node31670;
																assign node31670 = (inp[14]) ? 4'b1001 : 4'b1000;
													assign node31674 = (inp[12]) ? 4'b1110 : node31675;
														assign node31675 = (inp[8]) ? node31677 : 4'b1000;
															assign node31677 = (inp[7]) ? node31681 : node31678;
																assign node31678 = (inp[14]) ? 4'b1001 : 4'b1000;
																assign node31681 = (inp[14]) ? 4'b1000 : 4'b1001;
												assign node31685 = (inp[9]) ? node31703 : node31686;
													assign node31686 = (inp[12]) ? node31694 : node31687;
														assign node31687 = (inp[14]) ? node31689 : 4'b1000;
															assign node31689 = (inp[8]) ? 4'b1001 : node31690;
																assign node31690 = (inp[7]) ? 4'b1001 : 4'b1000;
														assign node31694 = (inp[14]) ? node31696 : 4'b1110;
															assign node31696 = (inp[8]) ? node31700 : node31697;
																assign node31697 = (inp[7]) ? 4'b1111 : 4'b1110;
																assign node31700 = (inp[7]) ? 4'b1110 : 4'b1111;
													assign node31703 = (inp[12]) ? node31713 : node31704;
														assign node31704 = (inp[8]) ? node31706 : 4'b1110;
															assign node31706 = (inp[14]) ? node31710 : node31707;
																assign node31707 = (inp[7]) ? 4'b1111 : 4'b1110;
																assign node31710 = (inp[7]) ? 4'b1110 : 4'b1111;
														assign node31713 = (inp[14]) ? node31715 : 4'b1010;
															assign node31715 = (inp[8]) ? node31719 : node31716;
																assign node31716 = (inp[7]) ? 4'b1011 : 4'b1010;
																assign node31719 = (inp[7]) ? 4'b1010 : 4'b1011;
											assign node31722 = (inp[9]) ? node31772 : node31723;
												assign node31723 = (inp[12]) ? node31743 : node31724;
													assign node31724 = (inp[4]) ? node31738 : node31725;
														assign node31725 = (inp[7]) ? node31731 : node31726;
															assign node31726 = (inp[14]) ? node31728 : 4'b1110;
																assign node31728 = (inp[8]) ? 4'b1111 : 4'b1110;
															assign node31731 = (inp[14]) ? node31735 : node31732;
																assign node31732 = (inp[8]) ? 4'b1111 : 4'b1110;
																assign node31735 = (inp[8]) ? 4'b1110 : 4'b1111;
														assign node31738 = (inp[14]) ? node31740 : 4'b1010;
															assign node31740 = (inp[8]) ? 4'b1010 : 4'b1011;
													assign node31743 = (inp[4]) ? node31757 : node31744;
														assign node31744 = (inp[14]) ? node31752 : node31745;
															assign node31745 = (inp[7]) ? node31749 : node31746;
																assign node31746 = (inp[8]) ? 4'b1010 : 4'b1011;
																assign node31749 = (inp[8]) ? 4'b1011 : 4'b1010;
															assign node31752 = (inp[8]) ? node31754 : 4'b1011;
																assign node31754 = (inp[7]) ? 4'b1010 : 4'b1011;
														assign node31757 = (inp[14]) ? node31765 : node31758;
															assign node31758 = (inp[7]) ? node31762 : node31759;
																assign node31759 = (inp[8]) ? 4'b1110 : 4'b1111;
																assign node31762 = (inp[8]) ? 4'b1111 : 4'b1110;
															assign node31765 = (inp[8]) ? node31769 : node31766;
																assign node31766 = (inp[7]) ? 4'b1111 : 4'b1110;
																assign node31769 = (inp[7]) ? 4'b1110 : 4'b1111;
												assign node31772 = (inp[4]) ? node31794 : node31773;
													assign node31773 = (inp[12]) ? node31783 : node31774;
														assign node31774 = (inp[8]) ? node31776 : 4'b1011;
															assign node31776 = (inp[14]) ? node31780 : node31777;
																assign node31777 = (inp[7]) ? 4'b1011 : 4'b1010;
																assign node31780 = (inp[7]) ? 4'b1010 : 4'b1011;
														assign node31783 = (inp[8]) ? node31789 : node31784;
															assign node31784 = (inp[14]) ? node31786 : 4'b1110;
																assign node31786 = (inp[7]) ? 4'b1111 : 4'b1110;
															assign node31789 = (inp[14]) ? node31791 : 4'b1111;
																assign node31791 = (inp[7]) ? 4'b1110 : 4'b1111;
													assign node31794 = (inp[12]) ? node31802 : node31795;
														assign node31795 = (inp[7]) ? 4'b1110 : node31796;
															assign node31796 = (inp[8]) ? node31798 : 4'b1111;
																assign node31798 = (inp[14]) ? 4'b1111 : 4'b1110;
														assign node31802 = (inp[8]) ? node31810 : node31803;
															assign node31803 = (inp[14]) ? node31807 : node31804;
																assign node31804 = (inp[7]) ? 4'b1010 : 4'b1011;
																assign node31807 = (inp[7]) ? 4'b1011 : 4'b1010;
															assign node31810 = (inp[14]) ? 4'b1010 : node31811;
																assign node31811 = (inp[7]) ? 4'b1011 : 4'b1010;
								assign node31815 = (inp[9]) ? node32135 : node31816;
									assign node31816 = (inp[0]) ? node31956 : node31817;
										assign node31817 = (inp[3]) ? node31881 : node31818;
											assign node31818 = (inp[4]) ? node31844 : node31819;
												assign node31819 = (inp[12]) ? node31829 : node31820;
													assign node31820 = (inp[14]) ? node31822 : 4'b1101;
														assign node31822 = (inp[8]) ? node31826 : node31823;
															assign node31823 = (inp[7]) ? 4'b1101 : 4'b1100;
															assign node31826 = (inp[7]) ? 4'b1100 : 4'b1101;
													assign node31829 = (inp[8]) ? node31837 : node31830;
														assign node31830 = (inp[7]) ? node31834 : node31831;
															assign node31831 = (inp[14]) ? 4'b1000 : 4'b1001;
															assign node31834 = (inp[14]) ? 4'b1001 : 4'b1000;
														assign node31837 = (inp[5]) ? 4'b1001 : node31838;
															assign node31838 = (inp[14]) ? 4'b1001 : node31839;
																assign node31839 = (inp[7]) ? 4'b1001 : 4'b1000;
												assign node31844 = (inp[12]) ? node31858 : node31845;
													assign node31845 = (inp[14]) ? node31851 : node31846;
														assign node31846 = (inp[8]) ? 4'b1000 : node31847;
															assign node31847 = (inp[7]) ? 4'b1000 : 4'b1001;
														assign node31851 = (inp[8]) ? node31855 : node31852;
															assign node31852 = (inp[7]) ? 4'b1001 : 4'b1000;
															assign node31855 = (inp[7]) ? 4'b1000 : 4'b1001;
													assign node31858 = (inp[5]) ? node31870 : node31859;
														assign node31859 = (inp[8]) ? node31865 : node31860;
															assign node31860 = (inp[14]) ? node31862 : 4'b1100;
																assign node31862 = (inp[7]) ? 4'b1101 : 4'b1100;
															assign node31865 = (inp[7]) ? node31867 : 4'b1101;
																assign node31867 = (inp[14]) ? 4'b1100 : 4'b1101;
														assign node31870 = (inp[7]) ? node31876 : node31871;
															assign node31871 = (inp[14]) ? node31873 : 4'b1111;
																assign node31873 = (inp[8]) ? 4'b1111 : 4'b1110;
															assign node31876 = (inp[8]) ? 4'b1110 : node31877;
																assign node31877 = (inp[14]) ? 4'b1111 : 4'b1110;
											assign node31881 = (inp[5]) ? node31919 : node31882;
												assign node31882 = (inp[4]) ? node31900 : node31883;
													assign node31883 = (inp[12]) ? node31891 : node31884;
														assign node31884 = (inp[14]) ? node31886 : 4'b1101;
															assign node31886 = (inp[8]) ? node31888 : 4'b1101;
																assign node31888 = (inp[7]) ? 4'b1100 : 4'b1101;
														assign node31891 = (inp[14]) ? node31893 : 4'b1001;
															assign node31893 = (inp[8]) ? node31897 : node31894;
																assign node31894 = (inp[7]) ? 4'b1001 : 4'b1000;
																assign node31897 = (inp[7]) ? 4'b1000 : 4'b1001;
													assign node31900 = (inp[12]) ? node31906 : node31901;
														assign node31901 = (inp[8]) ? 4'b1001 : node31902;
															assign node31902 = (inp[7]) ? 4'b1000 : 4'b1001;
														assign node31906 = (inp[8]) ? node31912 : node31907;
															assign node31907 = (inp[7]) ? node31909 : 4'b1111;
																assign node31909 = (inp[14]) ? 4'b1111 : 4'b1110;
															assign node31912 = (inp[7]) ? node31916 : node31913;
																assign node31913 = (inp[14]) ? 4'b1111 : 4'b1110;
																assign node31916 = (inp[14]) ? 4'b1110 : 4'b1111;
												assign node31919 = (inp[4]) ? node31939 : node31920;
													assign node31920 = (inp[12]) ? node31930 : node31921;
														assign node31921 = (inp[8]) ? node31923 : 4'b1110;
															assign node31923 = (inp[7]) ? node31927 : node31924;
																assign node31924 = (inp[14]) ? 4'b1111 : 4'b1110;
																assign node31927 = (inp[14]) ? 4'b1110 : 4'b1111;
														assign node31930 = (inp[14]) ? node31932 : 4'b1010;
															assign node31932 = (inp[7]) ? node31936 : node31933;
																assign node31933 = (inp[8]) ? 4'b1011 : 4'b1010;
																assign node31936 = (inp[8]) ? 4'b1010 : 4'b1011;
													assign node31939 = (inp[12]) ? node31945 : node31940;
														assign node31940 = (inp[7]) ? 4'b1011 : node31941;
															assign node31941 = (inp[14]) ? 4'b1010 : 4'b1011;
														assign node31945 = (inp[7]) ? node31951 : node31946;
															assign node31946 = (inp[8]) ? 4'b1111 : node31947;
																assign node31947 = (inp[14]) ? 4'b1110 : 4'b1111;
															assign node31951 = (inp[8]) ? 4'b1110 : node31952;
																assign node31952 = (inp[14]) ? 4'b1111 : 4'b1110;
										assign node31956 = (inp[5]) ? node32042 : node31957;
											assign node31957 = (inp[3]) ? node32001 : node31958;
												assign node31958 = (inp[7]) ? node31984 : node31959;
													assign node31959 = (inp[4]) ? node31971 : node31960;
														assign node31960 = (inp[12]) ? node31966 : node31961;
															assign node31961 = (inp[14]) ? node31963 : 4'b1111;
																assign node31963 = (inp[8]) ? 4'b1111 : 4'b1110;
															assign node31966 = (inp[14]) ? node31968 : 4'b1011;
																assign node31968 = (inp[8]) ? 4'b1011 : 4'b1010;
														assign node31971 = (inp[12]) ? node31979 : node31972;
															assign node31972 = (inp[14]) ? node31976 : node31973;
																assign node31973 = (inp[8]) ? 4'b1010 : 4'b1011;
																assign node31976 = (inp[8]) ? 4'b1011 : 4'b1010;
															assign node31979 = (inp[14]) ? 4'b1110 : node31980;
																assign node31980 = (inp[8]) ? 4'b1110 : 4'b1111;
													assign node31984 = (inp[4]) ? node31994 : node31985;
														assign node31985 = (inp[12]) ? node31989 : node31986;
															assign node31986 = (inp[8]) ? 4'b1110 : 4'b1111;
															assign node31989 = (inp[14]) ? node31991 : 4'b1010;
																assign node31991 = (inp[8]) ? 4'b1010 : 4'b1011;
														assign node31994 = (inp[12]) ? node31996 : 4'b1010;
															assign node31996 = (inp[14]) ? 4'b1111 : node31997;
																assign node31997 = (inp[8]) ? 4'b1111 : 4'b1110;
												assign node32001 = (inp[12]) ? node32025 : node32002;
													assign node32002 = (inp[4]) ? node32014 : node32003;
														assign node32003 = (inp[7]) ? node32009 : node32004;
															assign node32004 = (inp[14]) ? node32006 : 4'b1110;
																assign node32006 = (inp[8]) ? 4'b1111 : 4'b1110;
															assign node32009 = (inp[14]) ? 4'b1111 : node32010;
																assign node32010 = (inp[8]) ? 4'b1111 : 4'b1110;
														assign node32014 = (inp[14]) ? node32020 : node32015;
															assign node32015 = (inp[7]) ? node32017 : 4'b1011;
																assign node32017 = (inp[8]) ? 4'b1011 : 4'b1010;
															assign node32020 = (inp[7]) ? node32022 : 4'b1010;
																assign node32022 = (inp[8]) ? 4'b1010 : 4'b1011;
													assign node32025 = (inp[4]) ? node32033 : node32026;
														assign node32026 = (inp[14]) ? node32028 : 4'b1010;
															assign node32028 = (inp[8]) ? 4'b1010 : node32029;
																assign node32029 = (inp[7]) ? 4'b1011 : 4'b1010;
														assign node32033 = (inp[8]) ? node32035 : 4'b1100;
															assign node32035 = (inp[7]) ? node32039 : node32036;
																assign node32036 = (inp[14]) ? 4'b1101 : 4'b1100;
																assign node32039 = (inp[14]) ? 4'b1100 : 4'b1101;
											assign node32042 = (inp[3]) ? node32090 : node32043;
												assign node32043 = (inp[12]) ? node32065 : node32044;
													assign node32044 = (inp[4]) ? node32054 : node32045;
														assign node32045 = (inp[8]) ? 4'b1111 : node32046;
															assign node32046 = (inp[7]) ? node32050 : node32047;
																assign node32047 = (inp[14]) ? 4'b1110 : 4'b1111;
																assign node32050 = (inp[14]) ? 4'b1111 : 4'b1110;
														assign node32054 = (inp[7]) ? node32060 : node32055;
															assign node32055 = (inp[14]) ? 4'b1011 : node32056;
																assign node32056 = (inp[8]) ? 4'b1010 : 4'b1011;
															assign node32060 = (inp[14]) ? node32062 : 4'b1010;
																assign node32062 = (inp[8]) ? 4'b1010 : 4'b1011;
													assign node32065 = (inp[4]) ? node32077 : node32066;
														assign node32066 = (inp[7]) ? node32072 : node32067;
															assign node32067 = (inp[14]) ? 4'b1010 : node32068;
																assign node32068 = (inp[8]) ? 4'b1010 : 4'b1011;
															assign node32072 = (inp[8]) ? 4'b1011 : node32073;
																assign node32073 = (inp[14]) ? 4'b1011 : 4'b1010;
														assign node32077 = (inp[14]) ? node32083 : node32078;
															assign node32078 = (inp[7]) ? 4'b1101 : node32079;
																assign node32079 = (inp[8]) ? 4'b1100 : 4'b1101;
															assign node32083 = (inp[7]) ? node32087 : node32084;
																assign node32084 = (inp[8]) ? 4'b1101 : 4'b1100;
																assign node32087 = (inp[8]) ? 4'b1100 : 4'b1101;
												assign node32090 = (inp[8]) ? node32120 : node32091;
													assign node32091 = (inp[12]) ? node32107 : node32092;
														assign node32092 = (inp[4]) ? node32100 : node32093;
															assign node32093 = (inp[14]) ? node32097 : node32094;
																assign node32094 = (inp[7]) ? 4'b1100 : 4'b1101;
																assign node32097 = (inp[7]) ? 4'b1101 : 4'b1100;
															assign node32100 = (inp[7]) ? node32104 : node32101;
																assign node32101 = (inp[14]) ? 4'b1000 : 4'b1001;
																assign node32104 = (inp[14]) ? 4'b1001 : 4'b1000;
														assign node32107 = (inp[4]) ? node32113 : node32108;
															assign node32108 = (inp[14]) ? node32110 : 4'b1000;
																assign node32110 = (inp[7]) ? 4'b1001 : 4'b1000;
															assign node32113 = (inp[14]) ? node32117 : node32114;
																assign node32114 = (inp[7]) ? 4'b1100 : 4'b1101;
																assign node32117 = (inp[7]) ? 4'b1101 : 4'b1100;
													assign node32120 = (inp[7]) ? node32126 : node32121;
														assign node32121 = (inp[14]) ? node32123 : 4'b1000;
															assign node32123 = (inp[4]) ? 4'b1001 : 4'b1101;
														assign node32126 = (inp[14]) ? node32132 : node32127;
															assign node32127 = (inp[4]) ? 4'b1101 : node32128;
																assign node32128 = (inp[12]) ? 4'b1001 : 4'b1101;
															assign node32132 = (inp[4]) ? 4'b1100 : 4'b1000;
									assign node32135 = (inp[0]) ? node32299 : node32136;
										assign node32136 = (inp[3]) ? node32214 : node32137;
											assign node32137 = (inp[5]) ? node32173 : node32138;
												assign node32138 = (inp[7]) ? node32160 : node32139;
													assign node32139 = (inp[12]) ? node32151 : node32140;
														assign node32140 = (inp[4]) ? node32148 : node32141;
															assign node32141 = (inp[14]) ? node32145 : node32142;
																assign node32142 = (inp[8]) ? 4'b1000 : 4'b1001;
																assign node32145 = (inp[8]) ? 4'b1001 : 4'b1000;
															assign node32148 = (inp[14]) ? 4'b1101 : 4'b1100;
														assign node32151 = (inp[4]) ? node32157 : node32152;
															assign node32152 = (inp[8]) ? 4'b1100 : node32153;
																assign node32153 = (inp[14]) ? 4'b1100 : 4'b1101;
															assign node32157 = (inp[8]) ? 4'b1001 : 4'b1000;
													assign node32160 = (inp[4]) ? node32164 : node32161;
														assign node32161 = (inp[12]) ? 4'b1101 : 4'b1001;
														assign node32164 = (inp[12]) ? node32166 : 4'b1101;
															assign node32166 = (inp[14]) ? node32170 : node32167;
																assign node32167 = (inp[8]) ? 4'b1001 : 4'b1000;
																assign node32170 = (inp[8]) ? 4'b1000 : 4'b1001;
												assign node32173 = (inp[4]) ? node32193 : node32174;
													assign node32174 = (inp[12]) ? node32186 : node32175;
														assign node32175 = (inp[8]) ? node32181 : node32176;
															assign node32176 = (inp[14]) ? 4'b1000 : node32177;
																assign node32177 = (inp[7]) ? 4'b1000 : 4'b1001;
															assign node32181 = (inp[7]) ? 4'b1001 : node32182;
																assign node32182 = (inp[14]) ? 4'b1001 : 4'b1000;
														assign node32186 = (inp[7]) ? 4'b1110 : node32187;
															assign node32187 = (inp[8]) ? 4'b1111 : node32188;
																assign node32188 = (inp[14]) ? 4'b1110 : 4'b1111;
													assign node32193 = (inp[12]) ? node32205 : node32194;
														assign node32194 = (inp[8]) ? node32200 : node32195;
															assign node32195 = (inp[7]) ? node32197 : 4'b1111;
																assign node32197 = (inp[14]) ? 4'b1111 : 4'b1110;
															assign node32200 = (inp[14]) ? node32202 : 4'b1110;
																assign node32202 = (inp[7]) ? 4'b1110 : 4'b1111;
														assign node32205 = (inp[14]) ? 4'b1011 : node32206;
															assign node32206 = (inp[7]) ? node32210 : node32207;
																assign node32207 = (inp[8]) ? 4'b1010 : 4'b1011;
																assign node32210 = (inp[8]) ? 4'b1011 : 4'b1010;
											assign node32214 = (inp[5]) ? node32254 : node32215;
												assign node32215 = (inp[4]) ? node32227 : node32216;
													assign node32216 = (inp[12]) ? node32224 : node32217;
														assign node32217 = (inp[7]) ? node32219 : 4'b1001;
															assign node32219 = (inp[8]) ? node32221 : 4'b1000;
																assign node32221 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node32224 = (inp[7]) ? 4'b1111 : 4'b1110;
													assign node32227 = (inp[12]) ? node32239 : node32228;
														assign node32228 = (inp[8]) ? node32234 : node32229;
															assign node32229 = (inp[7]) ? node32231 : 4'b1110;
																assign node32231 = (inp[14]) ? 4'b1111 : 4'b1110;
															assign node32234 = (inp[7]) ? node32236 : 4'b1111;
																assign node32236 = (inp[14]) ? 4'b1110 : 4'b1111;
														assign node32239 = (inp[7]) ? node32247 : node32240;
															assign node32240 = (inp[8]) ? node32244 : node32241;
																assign node32241 = (inp[14]) ? 4'b1010 : 4'b1011;
																assign node32244 = (inp[14]) ? 4'b1011 : 4'b1010;
															assign node32247 = (inp[14]) ? node32251 : node32248;
																assign node32248 = (inp[8]) ? 4'b1011 : 4'b1010;
																assign node32251 = (inp[8]) ? 4'b1010 : 4'b1011;
												assign node32254 = (inp[14]) ? node32274 : node32255;
													assign node32255 = (inp[7]) ? node32265 : node32256;
														assign node32256 = (inp[8]) ? node32262 : node32257;
															assign node32257 = (inp[4]) ? node32259 : 4'b1111;
																assign node32259 = (inp[12]) ? 4'b1011 : 4'b1111;
															assign node32262 = (inp[12]) ? 4'b1110 : 4'b1010;
														assign node32265 = (inp[8]) ? 4'b1111 : node32266;
															assign node32266 = (inp[4]) ? node32270 : node32267;
																assign node32267 = (inp[12]) ? 4'b1110 : 4'b1010;
																assign node32270 = (inp[12]) ? 4'b1010 : 4'b1110;
													assign node32274 = (inp[8]) ? node32288 : node32275;
														assign node32275 = (inp[7]) ? node32281 : node32276;
															assign node32276 = (inp[12]) ? node32278 : 4'b1110;
																assign node32278 = (inp[4]) ? 4'b1010 : 4'b1110;
															assign node32281 = (inp[12]) ? node32285 : node32282;
																assign node32282 = (inp[4]) ? 4'b1111 : 4'b1011;
																assign node32285 = (inp[4]) ? 4'b1011 : 4'b1111;
														assign node32288 = (inp[7]) ? node32294 : node32289;
															assign node32289 = (inp[4]) ? 4'b1011 : node32290;
																assign node32290 = (inp[12]) ? 4'b1111 : 4'b1011;
															assign node32294 = (inp[12]) ? node32296 : 4'b1010;
																assign node32296 = (inp[4]) ? 4'b1010 : 4'b1110;
										assign node32299 = (inp[3]) ? node32385 : node32300;
											assign node32300 = (inp[5]) ? node32354 : node32301;
												assign node32301 = (inp[14]) ? node32331 : node32302;
													assign node32302 = (inp[12]) ? node32318 : node32303;
														assign node32303 = (inp[4]) ? node32311 : node32304;
															assign node32304 = (inp[7]) ? node32308 : node32305;
																assign node32305 = (inp[8]) ? 4'b1010 : 4'b1011;
																assign node32308 = (inp[8]) ? 4'b1011 : 4'b1010;
															assign node32311 = (inp[8]) ? node32315 : node32312;
																assign node32312 = (inp[7]) ? 4'b1110 : 4'b1111;
																assign node32315 = (inp[7]) ? 4'b1111 : 4'b1110;
														assign node32318 = (inp[4]) ? node32324 : node32319;
															assign node32319 = (inp[7]) ? node32321 : 4'b1111;
																assign node32321 = (inp[8]) ? 4'b1111 : 4'b1110;
															assign node32324 = (inp[8]) ? node32328 : node32325;
																assign node32325 = (inp[7]) ? 4'b1010 : 4'b1011;
																assign node32328 = (inp[7]) ? 4'b1011 : 4'b1010;
													assign node32331 = (inp[12]) ? node32343 : node32332;
														assign node32332 = (inp[4]) ? node32338 : node32333;
															assign node32333 = (inp[7]) ? 4'b1011 : node32334;
																assign node32334 = (inp[8]) ? 4'b1011 : 4'b1010;
															assign node32338 = (inp[7]) ? node32340 : 4'b1111;
																assign node32340 = (inp[8]) ? 4'b1110 : 4'b1111;
														assign node32343 = (inp[4]) ? node32349 : node32344;
															assign node32344 = (inp[7]) ? 4'b1111 : node32345;
																assign node32345 = (inp[8]) ? 4'b1111 : 4'b1110;
															assign node32349 = (inp[7]) ? node32351 : 4'b1011;
																assign node32351 = (inp[8]) ? 4'b1010 : 4'b1011;
												assign node32354 = (inp[12]) ? node32370 : node32355;
													assign node32355 = (inp[4]) ? node32365 : node32356;
														assign node32356 = (inp[8]) ? node32358 : 4'b1011;
															assign node32358 = (inp[7]) ? node32362 : node32359;
																assign node32359 = (inp[14]) ? 4'b1011 : 4'b1010;
																assign node32362 = (inp[14]) ? 4'b1010 : 4'b1011;
														assign node32365 = (inp[7]) ? node32367 : 4'b1100;
															assign node32367 = (inp[14]) ? 4'b1101 : 4'b1100;
													assign node32370 = (inp[4]) ? node32378 : node32371;
														assign node32371 = (inp[7]) ? node32373 : 4'b1101;
															assign node32373 = (inp[14]) ? 4'b1100 : node32374;
																assign node32374 = (inp[8]) ? 4'b1101 : 4'b1100;
														assign node32378 = (inp[8]) ? node32380 : 4'b1000;
															assign node32380 = (inp[14]) ? node32382 : 4'b1001;
																assign node32382 = (inp[7]) ? 4'b1000 : 4'b1001;
											assign node32385 = (inp[12]) ? node32415 : node32386;
												assign node32386 = (inp[4]) ? node32404 : node32387;
													assign node32387 = (inp[5]) ? node32397 : node32388;
														assign node32388 = (inp[7]) ? 4'b1011 : node32389;
															assign node32389 = (inp[8]) ? node32393 : node32390;
																assign node32390 = (inp[14]) ? 4'b1010 : 4'b1011;
																assign node32393 = (inp[14]) ? 4'b1011 : 4'b1010;
														assign node32397 = (inp[8]) ? 4'b1000 : node32398;
															assign node32398 = (inp[14]) ? node32400 : 4'b1001;
																assign node32400 = (inp[7]) ? 4'b1001 : 4'b1000;
													assign node32404 = (inp[8]) ? node32410 : node32405;
														assign node32405 = (inp[5]) ? 4'b1100 : node32406;
															assign node32406 = (inp[14]) ? 4'b1100 : 4'b1101;
														assign node32410 = (inp[7]) ? 4'b1101 : node32411;
															assign node32411 = (inp[14]) ? 4'b1101 : 4'b1100;
												assign node32415 = (inp[4]) ? node32423 : node32416;
													assign node32416 = (inp[14]) ? node32420 : node32417;
														assign node32417 = (inp[7]) ? 4'b1101 : 4'b1100;
														assign node32420 = (inp[7]) ? 4'b1100 : 4'b1101;
													assign node32423 = (inp[14]) ? node32433 : node32424;
														assign node32424 = (inp[5]) ? 4'b1001 : node32425;
															assign node32425 = (inp[8]) ? node32429 : node32426;
																assign node32426 = (inp[7]) ? 4'b1000 : 4'b1001;
																assign node32429 = (inp[7]) ? 4'b1001 : 4'b1000;
														assign node32433 = (inp[5]) ? node32437 : node32434;
															assign node32434 = (inp[7]) ? 4'b1001 : 4'b1000;
															assign node32437 = (inp[8]) ? node32439 : 4'b1000;
																assign node32439 = (inp[7]) ? 4'b1000 : 4'b1001;
							assign node32442 = (inp[3]) ? node32964 : node32443;
								assign node32443 = (inp[5]) ? node32739 : node32444;
									assign node32444 = (inp[8]) ? node32606 : node32445;
										assign node32445 = (inp[7]) ? node32537 : node32446;
											assign node32446 = (inp[0]) ? node32496 : node32447;
												assign node32447 = (inp[15]) ? node32469 : node32448;
													assign node32448 = (inp[9]) ? node32456 : node32449;
														assign node32449 = (inp[14]) ? node32451 : 4'b1010;
															assign node32451 = (inp[12]) ? 4'b1010 : node32452;
																assign node32452 = (inp[4]) ? 4'b1010 : 4'b1110;
														assign node32456 = (inp[14]) ? node32462 : node32457;
															assign node32457 = (inp[4]) ? node32459 : 4'b1110;
																assign node32459 = (inp[12]) ? 4'b1010 : 4'b1110;
															assign node32462 = (inp[12]) ? node32466 : node32463;
																assign node32463 = (inp[4]) ? 4'b1110 : 4'b1010;
																assign node32466 = (inp[4]) ? 4'b1010 : 4'b1110;
													assign node32469 = (inp[14]) ? node32483 : node32470;
														assign node32470 = (inp[12]) ? node32478 : node32471;
															assign node32471 = (inp[9]) ? node32475 : node32472;
																assign node32472 = (inp[4]) ? 4'b1000 : 4'b1100;
																assign node32475 = (inp[4]) ? 4'b1100 : 4'b1000;
															assign node32478 = (inp[9]) ? node32480 : 4'b1000;
																assign node32480 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node32483 = (inp[12]) ? node32489 : node32484;
															assign node32484 = (inp[9]) ? node32486 : 4'b1100;
																assign node32486 = (inp[4]) ? 4'b1100 : 4'b1000;
															assign node32489 = (inp[4]) ? node32493 : node32490;
																assign node32490 = (inp[9]) ? 4'b1100 : 4'b1000;
																assign node32493 = (inp[9]) ? 4'b1000 : 4'b1100;
												assign node32496 = (inp[15]) ? node32512 : node32497;
													assign node32497 = (inp[12]) ? 4'b1100 : node32498;
														assign node32498 = (inp[14]) ? node32506 : node32499;
															assign node32499 = (inp[9]) ? node32503 : node32500;
																assign node32500 = (inp[4]) ? 4'b1000 : 4'b1100;
																assign node32503 = (inp[4]) ? 4'b1100 : 4'b1000;
															assign node32506 = (inp[4]) ? node32508 : 4'b1000;
																assign node32508 = (inp[9]) ? 4'b1100 : 4'b1000;
													assign node32512 = (inp[14]) ? node32522 : node32513;
														assign node32513 = (inp[4]) ? 4'b1110 : node32514;
															assign node32514 = (inp[9]) ? node32518 : node32515;
																assign node32515 = (inp[12]) ? 4'b1010 : 4'b1110;
																assign node32518 = (inp[12]) ? 4'b1110 : 4'b1010;
														assign node32522 = (inp[9]) ? node32530 : node32523;
															assign node32523 = (inp[12]) ? node32527 : node32524;
																assign node32524 = (inp[4]) ? 4'b1010 : 4'b1110;
																assign node32527 = (inp[4]) ? 4'b1110 : 4'b1010;
															assign node32530 = (inp[12]) ? node32534 : node32531;
																assign node32531 = (inp[4]) ? 4'b1110 : 4'b1010;
																assign node32534 = (inp[4]) ? 4'b1010 : 4'b1110;
											assign node32537 = (inp[14]) ? node32569 : node32538;
												assign node32538 = (inp[9]) ? node32554 : node32539;
													assign node32539 = (inp[12]) ? node32545 : node32540;
														assign node32540 = (inp[4]) ? 4'b1011 : node32541;
															assign node32541 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node32545 = (inp[4]) ? node32547 : 4'b1011;
															assign node32547 = (inp[0]) ? node32551 : node32548;
																assign node32548 = (inp[15]) ? 4'b1101 : 4'b1111;
																assign node32551 = (inp[15]) ? 4'b1111 : 4'b1101;
													assign node32554 = (inp[0]) ? node32558 : node32555;
														assign node32555 = (inp[15]) ? 4'b1101 : 4'b1111;
														assign node32558 = (inp[15]) ? node32566 : node32559;
															assign node32559 = (inp[12]) ? node32563 : node32560;
																assign node32560 = (inp[4]) ? 4'b1101 : 4'b1001;
																assign node32563 = (inp[4]) ? 4'b1001 : 4'b1101;
															assign node32566 = (inp[4]) ? 4'b1011 : 4'b1111;
												assign node32569 = (inp[15]) ? node32587 : node32570;
													assign node32570 = (inp[0]) ? node32578 : node32571;
														assign node32571 = (inp[4]) ? 4'b1011 : node32572;
															assign node32572 = (inp[12]) ? 4'b1011 : node32573;
																assign node32573 = (inp[9]) ? 4'b1011 : 4'b1111;
														assign node32578 = (inp[9]) ? 4'b1001 : node32579;
															assign node32579 = (inp[12]) ? node32583 : node32580;
																assign node32580 = (inp[4]) ? 4'b1001 : 4'b1101;
																assign node32583 = (inp[4]) ? 4'b1101 : 4'b1001;
													assign node32587 = (inp[0]) ? node32599 : node32588;
														assign node32588 = (inp[4]) ? node32594 : node32589;
															assign node32589 = (inp[9]) ? 4'b1001 : node32590;
																assign node32590 = (inp[12]) ? 4'b1001 : 4'b1101;
															assign node32594 = (inp[12]) ? 4'b1101 : node32595;
																assign node32595 = (inp[9]) ? 4'b1101 : 4'b1001;
														assign node32599 = (inp[12]) ? 4'b1111 : node32600;
															assign node32600 = (inp[9]) ? node32602 : 4'b1011;
																assign node32602 = (inp[4]) ? 4'b1111 : 4'b1011;
										assign node32606 = (inp[7]) ? node32678 : node32607;
											assign node32607 = (inp[9]) ? node32653 : node32608;
												assign node32608 = (inp[14]) ? node32626 : node32609;
													assign node32609 = (inp[0]) ? node32617 : node32610;
														assign node32610 = (inp[15]) ? 4'b1001 : node32611;
															assign node32611 = (inp[4]) ? 4'b1011 : node32612;
																assign node32612 = (inp[12]) ? 4'b1011 : 4'b1111;
														assign node32617 = (inp[15]) ? node32623 : node32618;
															assign node32618 = (inp[12]) ? 4'b1001 : node32619;
																assign node32619 = (inp[4]) ? 4'b1001 : 4'b1101;
															assign node32623 = (inp[12]) ? 4'b1111 : 4'b1011;
													assign node32626 = (inp[0]) ? node32642 : node32627;
														assign node32627 = (inp[15]) ? node32635 : node32628;
															assign node32628 = (inp[4]) ? node32632 : node32629;
																assign node32629 = (inp[12]) ? 4'b1011 : 4'b1111;
																assign node32632 = (inp[12]) ? 4'b1111 : 4'b1011;
															assign node32635 = (inp[4]) ? node32639 : node32636;
																assign node32636 = (inp[12]) ? 4'b1001 : 4'b1101;
																assign node32639 = (inp[12]) ? 4'b1101 : 4'b1001;
														assign node32642 = (inp[15]) ? node32648 : node32643;
															assign node32643 = (inp[12]) ? 4'b1101 : node32644;
																assign node32644 = (inp[4]) ? 4'b1001 : 4'b1101;
															assign node32648 = (inp[12]) ? node32650 : 4'b1111;
																assign node32650 = (inp[4]) ? 4'b1111 : 4'b1011;
												assign node32653 = (inp[0]) ? node32667 : node32654;
													assign node32654 = (inp[15]) ? node32662 : node32655;
														assign node32655 = (inp[4]) ? node32659 : node32656;
															assign node32656 = (inp[12]) ? 4'b1111 : 4'b1011;
															assign node32659 = (inp[12]) ? 4'b1011 : 4'b1111;
														assign node32662 = (inp[12]) ? node32664 : 4'b1001;
															assign node32664 = (inp[4]) ? 4'b1001 : 4'b1101;
													assign node32667 = (inp[15]) ? node32671 : node32668;
														assign node32668 = (inp[12]) ? 4'b1001 : 4'b1101;
														assign node32671 = (inp[12]) ? node32675 : node32672;
															assign node32672 = (inp[4]) ? 4'b1111 : 4'b1011;
															assign node32675 = (inp[4]) ? 4'b1011 : 4'b1111;
											assign node32678 = (inp[0]) ? node32706 : node32679;
												assign node32679 = (inp[15]) ? node32697 : node32680;
													assign node32680 = (inp[12]) ? node32690 : node32681;
														assign node32681 = (inp[14]) ? 4'b1010 : node32682;
															assign node32682 = (inp[9]) ? node32686 : node32683;
																assign node32683 = (inp[4]) ? 4'b1010 : 4'b1110;
																assign node32686 = (inp[4]) ? 4'b1110 : 4'b1010;
														assign node32690 = (inp[4]) ? node32694 : node32691;
															assign node32691 = (inp[9]) ? 4'b1110 : 4'b1010;
															assign node32694 = (inp[9]) ? 4'b1010 : 4'b1110;
													assign node32697 = (inp[12]) ? 4'b1000 : node32698;
														assign node32698 = (inp[9]) ? node32702 : node32699;
															assign node32699 = (inp[4]) ? 4'b1000 : 4'b1100;
															assign node32702 = (inp[4]) ? 4'b1100 : 4'b1000;
												assign node32706 = (inp[15]) ? node32722 : node32707;
													assign node32707 = (inp[4]) ? node32715 : node32708;
														assign node32708 = (inp[14]) ? node32710 : 4'b1100;
															assign node32710 = (inp[12]) ? node32712 : 4'b1100;
																assign node32712 = (inp[9]) ? 4'b1100 : 4'b1000;
														assign node32715 = (inp[14]) ? node32717 : 4'b1000;
															assign node32717 = (inp[9]) ? 4'b1000 : node32718;
																assign node32718 = (inp[12]) ? 4'b1100 : 4'b1000;
													assign node32722 = (inp[12]) ? node32730 : node32723;
														assign node32723 = (inp[9]) ? node32727 : node32724;
															assign node32724 = (inp[4]) ? 4'b1010 : 4'b1110;
															assign node32727 = (inp[4]) ? 4'b1110 : 4'b1010;
														assign node32730 = (inp[14]) ? node32732 : 4'b1110;
															assign node32732 = (inp[9]) ? node32736 : node32733;
																assign node32733 = (inp[4]) ? 4'b1110 : 4'b1010;
																assign node32736 = (inp[4]) ? 4'b1010 : 4'b1110;
									assign node32739 = (inp[9]) ? node32857 : node32740;
										assign node32740 = (inp[8]) ? node32794 : node32741;
											assign node32741 = (inp[7]) ? node32767 : node32742;
												assign node32742 = (inp[0]) ? node32756 : node32743;
													assign node32743 = (inp[15]) ? node32751 : node32744;
														assign node32744 = (inp[4]) ? node32748 : node32745;
															assign node32745 = (inp[12]) ? 4'b1010 : 4'b1110;
															assign node32748 = (inp[12]) ? 4'b1100 : 4'b1010;
														assign node32751 = (inp[12]) ? node32753 : 4'b1000;
															assign node32753 = (inp[4]) ? 4'b1110 : 4'b1000;
													assign node32756 = (inp[15]) ? node32764 : node32757;
														assign node32757 = (inp[4]) ? node32761 : node32758;
															assign node32758 = (inp[12]) ? 4'b1000 : 4'b1100;
															assign node32761 = (inp[12]) ? 4'b1110 : 4'b1000;
														assign node32764 = (inp[4]) ? 4'b1010 : 4'b1110;
												assign node32767 = (inp[15]) ? node32779 : node32768;
													assign node32768 = (inp[0]) ? node32774 : node32769;
														assign node32769 = (inp[12]) ? 4'b1011 : node32770;
															assign node32770 = (inp[4]) ? 4'b1011 : 4'b1111;
														assign node32774 = (inp[4]) ? 4'b1111 : node32775;
															assign node32775 = (inp[12]) ? 4'b1001 : 4'b1101;
													assign node32779 = (inp[0]) ? node32785 : node32780;
														assign node32780 = (inp[12]) ? 4'b1111 : node32781;
															assign node32781 = (inp[4]) ? 4'b1001 : 4'b1101;
														assign node32785 = (inp[14]) ? node32787 : 4'b1011;
															assign node32787 = (inp[4]) ? node32791 : node32788;
																assign node32788 = (inp[12]) ? 4'b1011 : 4'b1111;
																assign node32791 = (inp[12]) ? 4'b1101 : 4'b1011;
											assign node32794 = (inp[7]) ? node32826 : node32795;
												assign node32795 = (inp[14]) ? node32809 : node32796;
													assign node32796 = (inp[0]) ? node32806 : node32797;
														assign node32797 = (inp[15]) ? node32801 : node32798;
															assign node32798 = (inp[12]) ? 4'b1011 : 4'b1111;
															assign node32801 = (inp[12]) ? 4'b1001 : node32802;
																assign node32802 = (inp[4]) ? 4'b1001 : 4'b1101;
														assign node32806 = (inp[15]) ? 4'b1011 : 4'b1001;
													assign node32809 = (inp[4]) ? node32817 : node32810;
														assign node32810 = (inp[12]) ? node32812 : 4'b1111;
															assign node32812 = (inp[15]) ? node32814 : 4'b1011;
																assign node32814 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node32817 = (inp[12]) ? node32819 : 4'b1001;
															assign node32819 = (inp[15]) ? node32823 : node32820;
																assign node32820 = (inp[0]) ? 4'b1111 : 4'b1101;
																assign node32823 = (inp[0]) ? 4'b1101 : 4'b1111;
												assign node32826 = (inp[15]) ? node32842 : node32827;
													assign node32827 = (inp[0]) ? node32833 : node32828;
														assign node32828 = (inp[12]) ? node32830 : 4'b1010;
															assign node32830 = (inp[4]) ? 4'b1100 : 4'b1010;
														assign node32833 = (inp[14]) ? node32839 : node32834;
															assign node32834 = (inp[12]) ? 4'b1000 : node32835;
																assign node32835 = (inp[4]) ? 4'b1000 : 4'b1100;
															assign node32839 = (inp[4]) ? 4'b1110 : 4'b1000;
													assign node32842 = (inp[0]) ? node32850 : node32843;
														assign node32843 = (inp[12]) ? node32847 : node32844;
															assign node32844 = (inp[4]) ? 4'b1000 : 4'b1100;
															assign node32847 = (inp[4]) ? 4'b1110 : 4'b1000;
														assign node32850 = (inp[4]) ? node32854 : node32851;
															assign node32851 = (inp[12]) ? 4'b1010 : 4'b1110;
															assign node32854 = (inp[12]) ? 4'b1100 : 4'b1010;
										assign node32857 = (inp[12]) ? node32917 : node32858;
											assign node32858 = (inp[4]) ? node32882 : node32859;
												assign node32859 = (inp[0]) ? node32869 : node32860;
													assign node32860 = (inp[15]) ? node32862 : 4'b1011;
														assign node32862 = (inp[8]) ? node32866 : node32863;
															assign node32863 = (inp[7]) ? 4'b1001 : 4'b1000;
															assign node32866 = (inp[7]) ? 4'b1000 : 4'b1001;
													assign node32869 = (inp[15]) ? node32877 : node32870;
														assign node32870 = (inp[7]) ? node32874 : node32871;
															assign node32871 = (inp[14]) ? 4'b1001 : 4'b1000;
															assign node32874 = (inp[8]) ? 4'b1000 : 4'b1001;
														assign node32877 = (inp[7]) ? 4'b1010 : node32878;
															assign node32878 = (inp[8]) ? 4'b1011 : 4'b1010;
												assign node32882 = (inp[8]) ? node32904 : node32883;
													assign node32883 = (inp[7]) ? node32891 : node32884;
														assign node32884 = (inp[14]) ? node32886 : 4'b1110;
															assign node32886 = (inp[15]) ? node32888 : 4'b1100;
																assign node32888 = (inp[0]) ? 4'b1100 : 4'b1110;
														assign node32891 = (inp[14]) ? node32897 : node32892;
															assign node32892 = (inp[0]) ? 4'b1101 : node32893;
																assign node32893 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node32897 = (inp[0]) ? node32901 : node32898;
																assign node32898 = (inp[15]) ? 4'b1111 : 4'b1101;
																assign node32901 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node32904 = (inp[7]) ? node32914 : node32905;
														assign node32905 = (inp[14]) ? 4'b1101 : node32906;
															assign node32906 = (inp[15]) ? node32910 : node32907;
																assign node32907 = (inp[0]) ? 4'b1111 : 4'b1101;
																assign node32910 = (inp[0]) ? 4'b1101 : 4'b1111;
														assign node32914 = (inp[14]) ? 4'b1110 : 4'b1100;
											assign node32917 = (inp[4]) ? node32941 : node32918;
												assign node32918 = (inp[8]) ? node32928 : node32919;
													assign node32919 = (inp[7]) ? node32921 : 4'b1100;
														assign node32921 = (inp[15]) ? node32925 : node32922;
															assign node32922 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node32925 = (inp[0]) ? 4'b1101 : 4'b1111;
													assign node32928 = (inp[7]) ? node32932 : node32929;
														assign node32929 = (inp[15]) ? 4'b1101 : 4'b1111;
														assign node32932 = (inp[14]) ? 4'b1110 : node32933;
															assign node32933 = (inp[15]) ? node32937 : node32934;
																assign node32934 = (inp[0]) ? 4'b1110 : 4'b1100;
																assign node32937 = (inp[0]) ? 4'b1100 : 4'b1110;
												assign node32941 = (inp[8]) ? node32953 : node32942;
													assign node32942 = (inp[7]) ? 4'b1001 : node32943;
														assign node32943 = (inp[14]) ? node32945 : 4'b1000;
															assign node32945 = (inp[0]) ? node32949 : node32946;
																assign node32946 = (inp[15]) ? 4'b1010 : 4'b1000;
																assign node32949 = (inp[15]) ? 4'b1000 : 4'b1010;
													assign node32953 = (inp[7]) ? node32957 : node32954;
														assign node32954 = (inp[15]) ? 4'b1001 : 4'b1011;
														assign node32957 = (inp[0]) ? node32961 : node32958;
															assign node32958 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node32961 = (inp[15]) ? 4'b1000 : 4'b1010;
								assign node32964 = (inp[9]) ? node33202 : node32965;
									assign node32965 = (inp[12]) ? node33107 : node32966;
										assign node32966 = (inp[4]) ? node33044 : node32967;
											assign node32967 = (inp[0]) ? node33003 : node32968;
												assign node32968 = (inp[5]) ? node32984 : node32969;
													assign node32969 = (inp[15]) ? node32977 : node32970;
														assign node32970 = (inp[7]) ? node32974 : node32971;
															assign node32971 = (inp[8]) ? 4'b1111 : 4'b1110;
															assign node32974 = (inp[8]) ? 4'b1110 : 4'b1111;
														assign node32977 = (inp[7]) ? node32981 : node32978;
															assign node32978 = (inp[8]) ? 4'b1101 : 4'b1100;
															assign node32981 = (inp[8]) ? 4'b1100 : 4'b1101;
													assign node32984 = (inp[15]) ? node32992 : node32985;
														assign node32985 = (inp[7]) ? node32989 : node32986;
															assign node32986 = (inp[8]) ? 4'b1101 : 4'b1100;
															assign node32989 = (inp[8]) ? 4'b1100 : 4'b1101;
														assign node32992 = (inp[14]) ? node32998 : node32993;
															assign node32993 = (inp[8]) ? 4'b1111 : node32994;
																assign node32994 = (inp[7]) ? 4'b1111 : 4'b1110;
															assign node32998 = (inp[7]) ? node33000 : 4'b1111;
																assign node33000 = (inp[8]) ? 4'b1110 : 4'b1111;
												assign node33003 = (inp[14]) ? node33021 : node33004;
													assign node33004 = (inp[7]) ? node33010 : node33005;
														assign node33005 = (inp[5]) ? node33007 : 4'b1100;
															assign node33007 = (inp[15]) ? 4'b1100 : 4'b1110;
														assign node33010 = (inp[8]) ? node33016 : node33011;
															assign node33011 = (inp[15]) ? node33013 : 4'b1111;
																assign node33013 = (inp[5]) ? 4'b1101 : 4'b1111;
															assign node33016 = (inp[5]) ? 4'b1110 : node33017;
																assign node33017 = (inp[15]) ? 4'b1110 : 4'b1100;
													assign node33021 = (inp[5]) ? node33031 : node33022;
														assign node33022 = (inp[15]) ? 4'b1110 : node33023;
															assign node33023 = (inp[7]) ? node33027 : node33024;
																assign node33024 = (inp[8]) ? 4'b1101 : 4'b1100;
																assign node33027 = (inp[8]) ? 4'b1100 : 4'b1101;
														assign node33031 = (inp[15]) ? node33037 : node33032;
															assign node33032 = (inp[8]) ? node33034 : 4'b1110;
																assign node33034 = (inp[7]) ? 4'b1110 : 4'b1111;
															assign node33037 = (inp[8]) ? node33041 : node33038;
																assign node33038 = (inp[7]) ? 4'b1101 : 4'b1100;
																assign node33041 = (inp[7]) ? 4'b1100 : 4'b1101;
											assign node33044 = (inp[7]) ? node33068 : node33045;
												assign node33045 = (inp[8]) ? node33059 : node33046;
													assign node33046 = (inp[15]) ? node33052 : node33047;
														assign node33047 = (inp[0]) ? node33049 : 4'b1010;
															assign node33049 = (inp[14]) ? 4'b1010 : 4'b1000;
														assign node33052 = (inp[0]) ? node33056 : node33053;
															assign node33053 = (inp[5]) ? 4'b1010 : 4'b1000;
															assign node33056 = (inp[5]) ? 4'b1000 : 4'b1010;
													assign node33059 = (inp[14]) ? 4'b1011 : node33060;
														assign node33060 = (inp[15]) ? 4'b1011 : node33061;
															assign node33061 = (inp[0]) ? node33063 : 4'b1001;
																assign node33063 = (inp[5]) ? 4'b1011 : 4'b1001;
												assign node33068 = (inp[8]) ? node33088 : node33069;
													assign node33069 = (inp[14]) ? node33083 : node33070;
														assign node33070 = (inp[5]) ? node33076 : node33071;
															assign node33071 = (inp[15]) ? 4'b1011 : node33072;
																assign node33072 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node33076 = (inp[15]) ? node33080 : node33077;
																assign node33077 = (inp[0]) ? 4'b1011 : 4'b1001;
																assign node33080 = (inp[0]) ? 4'b1001 : 4'b1011;
														assign node33083 = (inp[5]) ? 4'b1001 : node33084;
															assign node33084 = (inp[15]) ? 4'b1001 : 4'b1011;
													assign node33088 = (inp[0]) ? node33096 : node33089;
														assign node33089 = (inp[15]) ? node33093 : node33090;
															assign node33090 = (inp[5]) ? 4'b1000 : 4'b1010;
															assign node33093 = (inp[5]) ? 4'b1010 : 4'b1000;
														assign node33096 = (inp[14]) ? node33102 : node33097;
															assign node33097 = (inp[5]) ? node33099 : 4'b1000;
																assign node33099 = (inp[15]) ? 4'b1000 : 4'b1010;
															assign node33102 = (inp[15]) ? node33104 : 4'b1000;
																assign node33104 = (inp[5]) ? 4'b1000 : 4'b1010;
										assign node33107 = (inp[4]) ? node33173 : node33108;
											assign node33108 = (inp[8]) ? node33140 : node33109;
												assign node33109 = (inp[7]) ? node33125 : node33110;
													assign node33110 = (inp[15]) ? node33118 : node33111;
														assign node33111 = (inp[14]) ? 4'b1010 : node33112;
															assign node33112 = (inp[0]) ? node33114 : 4'b1000;
																assign node33114 = (inp[5]) ? 4'b1010 : 4'b1000;
														assign node33118 = (inp[14]) ? node33120 : 4'b1010;
															assign node33120 = (inp[0]) ? node33122 : 4'b1010;
																assign node33122 = (inp[5]) ? 4'b1000 : 4'b1010;
													assign node33125 = (inp[14]) ? 4'b1001 : node33126;
														assign node33126 = (inp[5]) ? node33132 : node33127;
															assign node33127 = (inp[15]) ? 4'b1001 : node33128;
																assign node33128 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node33132 = (inp[15]) ? node33136 : node33133;
																assign node33133 = (inp[0]) ? 4'b1011 : 4'b1001;
																assign node33136 = (inp[0]) ? 4'b1001 : 4'b1011;
												assign node33140 = (inp[7]) ? node33150 : node33141;
													assign node33141 = (inp[5]) ? node33145 : node33142;
														assign node33142 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node33145 = (inp[15]) ? 4'b1001 : node33146;
															assign node33146 = (inp[0]) ? 4'b1011 : 4'b1001;
													assign node33150 = (inp[15]) ? node33166 : node33151;
														assign node33151 = (inp[14]) ? node33159 : node33152;
															assign node33152 = (inp[0]) ? node33156 : node33153;
																assign node33153 = (inp[5]) ? 4'b1000 : 4'b1010;
																assign node33156 = (inp[5]) ? 4'b1010 : 4'b1000;
															assign node33159 = (inp[0]) ? node33163 : node33160;
																assign node33160 = (inp[5]) ? 4'b1000 : 4'b1010;
																assign node33163 = (inp[5]) ? 4'b1010 : 4'b1000;
														assign node33166 = (inp[0]) ? node33170 : node33167;
															assign node33167 = (inp[5]) ? 4'b1010 : 4'b1000;
															assign node33170 = (inp[5]) ? 4'b1000 : 4'b1010;
											assign node33173 = (inp[7]) ? node33189 : node33174;
												assign node33174 = (inp[8]) ? node33184 : node33175;
													assign node33175 = (inp[14]) ? node33177 : 4'b1100;
														assign node33177 = (inp[15]) ? node33181 : node33178;
															assign node33178 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node33181 = (inp[0]) ? 4'b1100 : 4'b1110;
													assign node33184 = (inp[15]) ? node33186 : 4'b1101;
														assign node33186 = (inp[0]) ? 4'b1101 : 4'b1111;
												assign node33189 = (inp[8]) ? node33195 : node33190;
													assign node33190 = (inp[0]) ? node33192 : 4'b1101;
														assign node33192 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node33195 = (inp[0]) ? node33199 : node33196;
														assign node33196 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node33199 = (inp[15]) ? 4'b1100 : 4'b1110;
									assign node33202 = (inp[15]) ? node33302 : node33203;
										assign node33203 = (inp[0]) ? node33261 : node33204;
											assign node33204 = (inp[12]) ? node33232 : node33205;
												assign node33205 = (inp[4]) ? node33223 : node33206;
													assign node33206 = (inp[5]) ? node33212 : node33207;
														assign node33207 = (inp[7]) ? 4'b1011 : node33208;
															assign node33208 = (inp[8]) ? 4'b1011 : 4'b1010;
														assign node33212 = (inp[14]) ? node33218 : node33213;
															assign node33213 = (inp[8]) ? node33215 : 4'b1000;
																assign node33215 = (inp[7]) ? 4'b1000 : 4'b1001;
															assign node33218 = (inp[7]) ? node33220 : 4'b1000;
																assign node33220 = (inp[8]) ? 4'b1000 : 4'b1001;
													assign node33223 = (inp[14]) ? 4'b1100 : node33224;
														assign node33224 = (inp[8]) ? node33228 : node33225;
															assign node33225 = (inp[7]) ? 4'b1101 : 4'b1100;
															assign node33228 = (inp[7]) ? 4'b1100 : 4'b1101;
												assign node33232 = (inp[4]) ? node33246 : node33233;
													assign node33233 = (inp[5]) ? node33241 : node33234;
														assign node33234 = (inp[7]) ? node33238 : node33235;
															assign node33235 = (inp[8]) ? 4'b1101 : 4'b1100;
															assign node33238 = (inp[8]) ? 4'b1100 : 4'b1101;
														assign node33241 = (inp[7]) ? node33243 : 4'b1101;
															assign node33243 = (inp[8]) ? 4'b1100 : 4'b1101;
													assign node33246 = (inp[14]) ? node33254 : node33247;
														assign node33247 = (inp[8]) ? node33251 : node33248;
															assign node33248 = (inp[7]) ? 4'b1001 : 4'b1000;
															assign node33251 = (inp[7]) ? 4'b1000 : 4'b1001;
														assign node33254 = (inp[7]) ? node33258 : node33255;
															assign node33255 = (inp[8]) ? 4'b1001 : 4'b1000;
															assign node33258 = (inp[8]) ? 4'b1000 : 4'b1001;
											assign node33261 = (inp[12]) ? node33285 : node33262;
												assign node33262 = (inp[4]) ? node33278 : node33263;
													assign node33263 = (inp[5]) ? node33271 : node33264;
														assign node33264 = (inp[7]) ? node33268 : node33265;
															assign node33265 = (inp[8]) ? 4'b1001 : 4'b1000;
															assign node33268 = (inp[8]) ? 4'b1000 : 4'b1001;
														assign node33271 = (inp[14]) ? node33275 : node33272;
															assign node33272 = (inp[7]) ? 4'b1010 : 4'b1011;
															assign node33275 = (inp[7]) ? 4'b1011 : 4'b1010;
													assign node33278 = (inp[14]) ? 4'b1111 : node33279;
														assign node33279 = (inp[8]) ? node33281 : 4'b1110;
															assign node33281 = (inp[7]) ? 4'b1110 : 4'b1111;
												assign node33285 = (inp[4]) ? node33297 : node33286;
													assign node33286 = (inp[5]) ? node33290 : node33287;
														assign node33287 = (inp[14]) ? 4'b1110 : 4'b1111;
														assign node33290 = (inp[7]) ? node33294 : node33291;
															assign node33291 = (inp[8]) ? 4'b1111 : 4'b1110;
															assign node33294 = (inp[8]) ? 4'b1110 : 4'b1111;
													assign node33297 = (inp[7]) ? node33299 : 4'b1011;
														assign node33299 = (inp[8]) ? 4'b1010 : 4'b1011;
										assign node33302 = (inp[0]) ? node33346 : node33303;
											assign node33303 = (inp[4]) ? node33333 : node33304;
												assign node33304 = (inp[12]) ? node33318 : node33305;
													assign node33305 = (inp[5]) ? node33313 : node33306;
														assign node33306 = (inp[8]) ? node33310 : node33307;
															assign node33307 = (inp[7]) ? 4'b1001 : 4'b1000;
															assign node33310 = (inp[7]) ? 4'b1000 : 4'b1001;
														assign node33313 = (inp[7]) ? 4'b1010 : node33314;
															assign node33314 = (inp[8]) ? 4'b1011 : 4'b1010;
													assign node33318 = (inp[5]) ? node33320 : 4'b1110;
														assign node33320 = (inp[14]) ? node33328 : node33321;
															assign node33321 = (inp[7]) ? node33325 : node33322;
																assign node33322 = (inp[8]) ? 4'b1111 : 4'b1110;
																assign node33325 = (inp[8]) ? 4'b1110 : 4'b1111;
															assign node33328 = (inp[8]) ? 4'b1110 : node33329;
																assign node33329 = (inp[7]) ? 4'b1111 : 4'b1110;
												assign node33333 = (inp[12]) ? node33341 : node33334;
													assign node33334 = (inp[7]) ? node33338 : node33335;
														assign node33335 = (inp[8]) ? 4'b1111 : 4'b1110;
														assign node33338 = (inp[8]) ? 4'b1110 : 4'b1111;
													assign node33341 = (inp[7]) ? 4'b1011 : node33342;
														assign node33342 = (inp[8]) ? 4'b1011 : 4'b1010;
											assign node33346 = (inp[5]) ? node33374 : node33347;
												assign node33347 = (inp[12]) ? node33361 : node33348;
													assign node33348 = (inp[4]) ? node33354 : node33349;
														assign node33349 = (inp[8]) ? node33351 : 4'b1011;
															assign node33351 = (inp[7]) ? 4'b1010 : 4'b1011;
														assign node33354 = (inp[7]) ? node33358 : node33355;
															assign node33355 = (inp[8]) ? 4'b1101 : 4'b1100;
															assign node33358 = (inp[8]) ? 4'b1100 : 4'b1101;
													assign node33361 = (inp[4]) ? node33369 : node33362;
														assign node33362 = (inp[8]) ? node33366 : node33363;
															assign node33363 = (inp[7]) ? 4'b1101 : 4'b1100;
															assign node33366 = (inp[7]) ? 4'b1100 : 4'b1101;
														assign node33369 = (inp[8]) ? 4'b1001 : node33370;
															assign node33370 = (inp[14]) ? 4'b1001 : 4'b1000;
												assign node33374 = (inp[8]) ? node33392 : node33375;
													assign node33375 = (inp[7]) ? node33383 : node33376;
														assign node33376 = (inp[12]) ? node33380 : node33377;
															assign node33377 = (inp[4]) ? 4'b1100 : 4'b1000;
															assign node33380 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node33383 = (inp[14]) ? 4'b1001 : node33384;
															assign node33384 = (inp[4]) ? node33388 : node33385;
																assign node33385 = (inp[12]) ? 4'b1101 : 4'b1001;
																assign node33388 = (inp[12]) ? 4'b1001 : 4'b1101;
													assign node33392 = (inp[7]) ? node33398 : node33393;
														assign node33393 = (inp[14]) ? node33395 : 4'b1101;
															assign node33395 = (inp[4]) ? 4'b1101 : 4'b1001;
														assign node33398 = (inp[4]) ? node33400 : 4'b1100;
															assign node33400 = (inp[12]) ? 4'b1000 : 4'b1100;
						assign node33403 = (inp[7]) ? node34551 : node33404;
							assign node33404 = (inp[8]) ? node33986 : node33405;
								assign node33405 = (inp[14]) ? node33699 : node33406;
									assign node33406 = (inp[2]) ? node33568 : node33407;
										assign node33407 = (inp[9]) ? node33497 : node33408;
											assign node33408 = (inp[0]) ? node33446 : node33409;
												assign node33409 = (inp[3]) ? node33429 : node33410;
													assign node33410 = (inp[15]) ? node33422 : node33411;
														assign node33411 = (inp[5]) ? node33417 : node33412;
															assign node33412 = (inp[12]) ? 4'b1111 : node33413;
																assign node33413 = (inp[4]) ? 4'b1011 : 4'b1111;
															assign node33417 = (inp[4]) ? node33419 : 4'b1011;
																assign node33419 = (inp[12]) ? 4'b1101 : 4'b1011;
														assign node33422 = (inp[5]) ? node33424 : 4'b1001;
															assign node33424 = (inp[4]) ? 4'b1111 : node33425;
																assign node33425 = (inp[12]) ? 4'b1001 : 4'b1101;
													assign node33429 = (inp[15]) ? node33441 : node33430;
														assign node33430 = (inp[5]) ? node33436 : node33431;
															assign node33431 = (inp[12]) ? 4'b1101 : node33432;
																assign node33432 = (inp[4]) ? 4'b1011 : 4'b1111;
															assign node33436 = (inp[12]) ? node33438 : 4'b1101;
																assign node33438 = (inp[4]) ? 4'b1101 : 4'b1001;
														assign node33441 = (inp[5]) ? node33443 : 4'b1101;
															assign node33443 = (inp[4]) ? 4'b1111 : 4'b1011;
												assign node33446 = (inp[15]) ? node33474 : node33447;
													assign node33447 = (inp[3]) ? node33461 : node33448;
														assign node33448 = (inp[5]) ? node33456 : node33449;
															assign node33449 = (inp[4]) ? node33453 : node33450;
																assign node33450 = (inp[12]) ? 4'b1001 : 4'b1101;
																assign node33453 = (inp[12]) ? 4'b1101 : 4'b1001;
															assign node33456 = (inp[4]) ? 4'b1001 : node33457;
																assign node33457 = (inp[12]) ? 4'b1001 : 4'b1101;
														assign node33461 = (inp[5]) ? node33467 : node33462;
															assign node33462 = (inp[4]) ? 4'b1001 : node33463;
																assign node33463 = (inp[12]) ? 4'b1001 : 4'b1101;
															assign node33467 = (inp[4]) ? node33471 : node33468;
																assign node33468 = (inp[12]) ? 4'b1011 : 4'b1111;
																assign node33471 = (inp[12]) ? 4'b1111 : 4'b1011;
													assign node33474 = (inp[3]) ? node33482 : node33475;
														assign node33475 = (inp[12]) ? node33479 : node33476;
															assign node33476 = (inp[4]) ? 4'b1011 : 4'b1111;
															assign node33479 = (inp[4]) ? 4'b1101 : 4'b1011;
														assign node33482 = (inp[5]) ? node33490 : node33483;
															assign node33483 = (inp[4]) ? node33487 : node33484;
																assign node33484 = (inp[12]) ? 4'b1011 : 4'b1111;
																assign node33487 = (inp[12]) ? 4'b1101 : 4'b1011;
															assign node33490 = (inp[12]) ? node33494 : node33491;
																assign node33491 = (inp[4]) ? 4'b1001 : 4'b1101;
																assign node33494 = (inp[4]) ? 4'b1101 : 4'b1001;
											assign node33497 = (inp[12]) ? node33537 : node33498;
												assign node33498 = (inp[4]) ? node33522 : node33499;
													assign node33499 = (inp[3]) ? node33507 : node33500;
														assign node33500 = (inp[15]) ? node33504 : node33501;
															assign node33501 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node33504 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node33507 = (inp[15]) ? node33515 : node33508;
															assign node33508 = (inp[0]) ? node33512 : node33509;
																assign node33509 = (inp[5]) ? 4'b1001 : 4'b1011;
																assign node33512 = (inp[5]) ? 4'b1011 : 4'b1001;
															assign node33515 = (inp[0]) ? node33519 : node33516;
																assign node33516 = (inp[5]) ? 4'b1011 : 4'b1001;
																assign node33519 = (inp[5]) ? 4'b1001 : 4'b1011;
													assign node33522 = (inp[0]) ? node33528 : node33523;
														assign node33523 = (inp[15]) ? 4'b1111 : node33524;
															assign node33524 = (inp[5]) ? 4'b1101 : 4'b1111;
														assign node33528 = (inp[15]) ? node33534 : node33529;
															assign node33529 = (inp[3]) ? 4'b1111 : node33530;
																assign node33530 = (inp[5]) ? 4'b1111 : 4'b1101;
															assign node33534 = (inp[3]) ? 4'b1101 : 4'b1111;
												assign node33537 = (inp[4]) ? node33553 : node33538;
													assign node33538 = (inp[0]) ? node33548 : node33539;
														assign node33539 = (inp[15]) ? node33545 : node33540;
															assign node33540 = (inp[5]) ? 4'b1101 : node33541;
																assign node33541 = (inp[3]) ? 4'b1101 : 4'b1111;
															assign node33545 = (inp[3]) ? 4'b1111 : 4'b1101;
														assign node33548 = (inp[15]) ? node33550 : 4'b1111;
															assign node33550 = (inp[3]) ? 4'b1101 : 4'b1111;
													assign node33553 = (inp[15]) ? node33563 : node33554;
														assign node33554 = (inp[0]) ? node33558 : node33555;
															assign node33555 = (inp[5]) ? 4'b1001 : 4'b1011;
															assign node33558 = (inp[3]) ? 4'b1011 : node33559;
																assign node33559 = (inp[5]) ? 4'b1011 : 4'b1001;
														assign node33563 = (inp[0]) ? 4'b1001 : node33564;
															assign node33564 = (inp[5]) ? 4'b1011 : 4'b1001;
										assign node33568 = (inp[12]) ? node33630 : node33569;
											assign node33569 = (inp[3]) ? node33591 : node33570;
												assign node33570 = (inp[9]) ? node33582 : node33571;
													assign node33571 = (inp[4]) ? 4'b1010 : node33572;
														assign node33572 = (inp[5]) ? node33574 : 4'b1100;
															assign node33574 = (inp[0]) ? node33578 : node33575;
																assign node33575 = (inp[15]) ? 4'b1100 : 4'b1110;
																assign node33578 = (inp[15]) ? 4'b1110 : 4'b1100;
													assign node33582 = (inp[4]) ? node33584 : 4'b1010;
														assign node33584 = (inp[15]) ? 4'b1110 : node33585;
															assign node33585 = (inp[5]) ? node33587 : 4'b1110;
																assign node33587 = (inp[0]) ? 4'b1110 : 4'b1100;
												assign node33591 = (inp[5]) ? node33611 : node33592;
													assign node33592 = (inp[9]) ? node33600 : node33593;
														assign node33593 = (inp[4]) ? node33595 : 4'b1110;
															assign node33595 = (inp[15]) ? 4'b1000 : node33596;
																assign node33596 = (inp[0]) ? 4'b1000 : 4'b1010;
														assign node33600 = (inp[4]) ? node33606 : node33601;
															assign node33601 = (inp[15]) ? node33603 : 4'b1000;
																assign node33603 = (inp[0]) ? 4'b1010 : 4'b1000;
															assign node33606 = (inp[15]) ? 4'b1100 : node33607;
																assign node33607 = (inp[0]) ? 4'b1110 : 4'b1100;
													assign node33611 = (inp[0]) ? node33621 : node33612;
														assign node33612 = (inp[15]) ? node33614 : 4'b1000;
															assign node33614 = (inp[9]) ? node33618 : node33615;
																assign node33615 = (inp[4]) ? 4'b1010 : 4'b1110;
																assign node33618 = (inp[4]) ? 4'b1110 : 4'b1010;
														assign node33621 = (inp[15]) ? node33627 : node33622;
															assign node33622 = (inp[4]) ? node33624 : 4'b1110;
																assign node33624 = (inp[9]) ? 4'b1110 : 4'b1010;
															assign node33627 = (inp[4]) ? 4'b1000 : 4'b1100;
											assign node33630 = (inp[9]) ? node33664 : node33631;
												assign node33631 = (inp[4]) ? node33649 : node33632;
													assign node33632 = (inp[15]) ? node33638 : node33633;
														assign node33633 = (inp[0]) ? 4'b1000 : node33634;
															assign node33634 = (inp[3]) ? 4'b1000 : 4'b1010;
														assign node33638 = (inp[0]) ? node33644 : node33639;
															assign node33639 = (inp[5]) ? node33641 : 4'b1000;
																assign node33641 = (inp[3]) ? 4'b1010 : 4'b1000;
															assign node33644 = (inp[3]) ? node33646 : 4'b1010;
																assign node33646 = (inp[5]) ? 4'b1000 : 4'b1010;
													assign node33649 = (inp[15]) ? node33653 : node33650;
														assign node33650 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node33653 = (inp[0]) ? node33659 : node33654;
															assign node33654 = (inp[5]) ? 4'b1110 : node33655;
																assign node33655 = (inp[3]) ? 4'b1110 : 4'b1100;
															assign node33659 = (inp[5]) ? 4'b1100 : node33660;
																assign node33660 = (inp[3]) ? 4'b1100 : 4'b1110;
												assign node33664 = (inp[4]) ? node33682 : node33665;
													assign node33665 = (inp[5]) ? node33675 : node33666;
														assign node33666 = (inp[3]) ? 4'b1100 : node33667;
															assign node33667 = (inp[0]) ? node33671 : node33668;
																assign node33668 = (inp[15]) ? 4'b1100 : 4'b1110;
																assign node33671 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node33675 = (inp[15]) ? node33679 : node33676;
															assign node33676 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node33679 = (inp[3]) ? 4'b1110 : 4'b1100;
													assign node33682 = (inp[15]) ? node33688 : node33683;
														assign node33683 = (inp[0]) ? 4'b1010 : node33684;
															assign node33684 = (inp[5]) ? 4'b1000 : 4'b1010;
														assign node33688 = (inp[0]) ? node33694 : node33689;
															assign node33689 = (inp[3]) ? 4'b1010 : node33690;
																assign node33690 = (inp[5]) ? 4'b1010 : 4'b1000;
															assign node33694 = (inp[3]) ? 4'b1000 : node33695;
																assign node33695 = (inp[5]) ? 4'b1000 : 4'b1010;
									assign node33699 = (inp[3]) ? node33813 : node33700;
										assign node33700 = (inp[9]) ? node33744 : node33701;
											assign node33701 = (inp[0]) ? node33715 : node33702;
												assign node33702 = (inp[15]) ? node33708 : node33703;
													assign node33703 = (inp[4]) ? 4'b1010 : node33704;
														assign node33704 = (inp[12]) ? 4'b1010 : 4'b1110;
													assign node33708 = (inp[4]) ? node33712 : node33709;
														assign node33709 = (inp[12]) ? 4'b1000 : 4'b1100;
														assign node33712 = (inp[12]) ? 4'b1100 : 4'b1000;
												assign node33715 = (inp[15]) ? node33727 : node33716;
													assign node33716 = (inp[2]) ? node33722 : node33717;
														assign node33717 = (inp[12]) ? node33719 : 4'b1000;
															assign node33719 = (inp[5]) ? 4'b1110 : 4'b1000;
														assign node33722 = (inp[12]) ? node33724 : 4'b1100;
															assign node33724 = (inp[4]) ? 4'b1100 : 4'b1000;
													assign node33727 = (inp[2]) ? node33735 : node33728;
														assign node33728 = (inp[12]) ? node33732 : node33729;
															assign node33729 = (inp[4]) ? 4'b1010 : 4'b1110;
															assign node33732 = (inp[4]) ? 4'b1110 : 4'b1010;
														assign node33735 = (inp[4]) ? node33739 : node33736;
															assign node33736 = (inp[12]) ? 4'b1010 : 4'b1110;
															assign node33739 = (inp[12]) ? node33741 : 4'b1010;
																assign node33741 = (inp[5]) ? 4'b1100 : 4'b1110;
											assign node33744 = (inp[15]) ? node33784 : node33745;
												assign node33745 = (inp[0]) ? node33761 : node33746;
													assign node33746 = (inp[5]) ? node33754 : node33747;
														assign node33747 = (inp[12]) ? node33751 : node33748;
															assign node33748 = (inp[4]) ? 4'b1110 : 4'b1010;
															assign node33751 = (inp[4]) ? 4'b1010 : 4'b1110;
														assign node33754 = (inp[4]) ? node33758 : node33755;
															assign node33755 = (inp[12]) ? 4'b1100 : 4'b1010;
															assign node33758 = (inp[12]) ? 4'b1000 : 4'b1100;
													assign node33761 = (inp[5]) ? node33777 : node33762;
														assign node33762 = (inp[2]) ? node33770 : node33763;
															assign node33763 = (inp[12]) ? node33767 : node33764;
																assign node33764 = (inp[4]) ? 4'b1100 : 4'b1000;
																assign node33767 = (inp[4]) ? 4'b1000 : 4'b1100;
															assign node33770 = (inp[12]) ? node33774 : node33771;
																assign node33771 = (inp[4]) ? 4'b1100 : 4'b1000;
																assign node33774 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node33777 = (inp[4]) ? node33781 : node33778;
															assign node33778 = (inp[12]) ? 4'b1110 : 4'b1000;
															assign node33781 = (inp[12]) ? 4'b1010 : 4'b1110;
												assign node33784 = (inp[0]) ? node33800 : node33785;
													assign node33785 = (inp[5]) ? node33795 : node33786;
														assign node33786 = (inp[2]) ? 4'b1000 : node33787;
															assign node33787 = (inp[12]) ? node33791 : node33788;
																assign node33788 = (inp[4]) ? 4'b1100 : 4'b1000;
																assign node33791 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node33795 = (inp[4]) ? node33797 : 4'b1000;
															assign node33797 = (inp[12]) ? 4'b1010 : 4'b1110;
													assign node33800 = (inp[5]) ? node33806 : node33801;
														assign node33801 = (inp[12]) ? 4'b1010 : node33802;
															assign node33802 = (inp[4]) ? 4'b1110 : 4'b1010;
														assign node33806 = (inp[12]) ? node33810 : node33807;
															assign node33807 = (inp[2]) ? 4'b1100 : 4'b1010;
															assign node33810 = (inp[4]) ? 4'b1000 : 4'b1100;
										assign node33813 = (inp[2]) ? node33901 : node33814;
											assign node33814 = (inp[12]) ? node33860 : node33815;
												assign node33815 = (inp[15]) ? node33843 : node33816;
													assign node33816 = (inp[5]) ? node33830 : node33817;
														assign node33817 = (inp[0]) ? node33825 : node33818;
															assign node33818 = (inp[9]) ? node33822 : node33819;
																assign node33819 = (inp[4]) ? 4'b1010 : 4'b1110;
																assign node33822 = (inp[4]) ? 4'b1100 : 4'b1010;
															assign node33825 = (inp[4]) ? 4'b1000 : node33826;
																assign node33826 = (inp[9]) ? 4'b1000 : 4'b1100;
														assign node33830 = (inp[0]) ? node33836 : node33831;
															assign node33831 = (inp[4]) ? node33833 : 4'b1000;
																assign node33833 = (inp[9]) ? 4'b1100 : 4'b1000;
															assign node33836 = (inp[4]) ? node33840 : node33837;
																assign node33837 = (inp[9]) ? 4'b1010 : 4'b1110;
																assign node33840 = (inp[9]) ? 4'b1110 : 4'b1010;
													assign node33843 = (inp[4]) ? node33851 : node33844;
														assign node33844 = (inp[9]) ? node33846 : 4'b1100;
															assign node33846 = (inp[0]) ? node33848 : 4'b1000;
																assign node33848 = (inp[5]) ? 4'b1000 : 4'b1010;
														assign node33851 = (inp[9]) ? node33857 : node33852;
															assign node33852 = (inp[5]) ? node33854 : 4'b1010;
																assign node33854 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node33857 = (inp[5]) ? 4'b1110 : 4'b1100;
												assign node33860 = (inp[15]) ? node33878 : node33861;
													assign node33861 = (inp[0]) ? node33869 : node33862;
														assign node33862 = (inp[5]) ? node33864 : 4'b1000;
															assign node33864 = (inp[9]) ? 4'b1100 : node33865;
																assign node33865 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node33869 = (inp[4]) ? node33875 : node33870;
															assign node33870 = (inp[9]) ? 4'b1110 : node33871;
																assign node33871 = (inp[5]) ? 4'b1010 : 4'b1000;
															assign node33875 = (inp[9]) ? 4'b1010 : 4'b1110;
													assign node33878 = (inp[0]) ? node33892 : node33879;
														assign node33879 = (inp[5]) ? node33885 : node33880;
															assign node33880 = (inp[4]) ? 4'b1110 : node33881;
																assign node33881 = (inp[9]) ? 4'b1110 : 4'b1000;
															assign node33885 = (inp[9]) ? node33889 : node33886;
																assign node33886 = (inp[4]) ? 4'b1110 : 4'b1010;
																assign node33889 = (inp[4]) ? 4'b1010 : 4'b1110;
														assign node33892 = (inp[4]) ? node33898 : node33893;
															assign node33893 = (inp[9]) ? 4'b1100 : node33894;
																assign node33894 = (inp[5]) ? 4'b1000 : 4'b1010;
															assign node33898 = (inp[9]) ? 4'b1000 : 4'b1100;
											assign node33901 = (inp[12]) ? node33945 : node33902;
												assign node33902 = (inp[5]) ? node33918 : node33903;
													assign node33903 = (inp[9]) ? node33915 : node33904;
														assign node33904 = (inp[4]) ? node33910 : node33905;
															assign node33905 = (inp[15]) ? 4'b1110 : node33906;
																assign node33906 = (inp[0]) ? 4'b1100 : 4'b1110;
															assign node33910 = (inp[15]) ? node33912 : 4'b1010;
																assign node33912 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node33915 = (inp[4]) ? 4'b1110 : 4'b1010;
													assign node33918 = (inp[4]) ? node33930 : node33919;
														assign node33919 = (inp[9]) ? node33925 : node33920;
															assign node33920 = (inp[15]) ? 4'b1110 : node33921;
																assign node33921 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node33925 = (inp[15]) ? node33927 : 4'b1010;
																assign node33927 = (inp[0]) ? 4'b1000 : 4'b1010;
														assign node33930 = (inp[9]) ? node33938 : node33931;
															assign node33931 = (inp[0]) ? node33935 : node33932;
																assign node33932 = (inp[15]) ? 4'b1010 : 4'b1000;
																assign node33935 = (inp[15]) ? 4'b1000 : 4'b1010;
															assign node33938 = (inp[15]) ? node33942 : node33939;
																assign node33939 = (inp[0]) ? 4'b1110 : 4'b1100;
																assign node33942 = (inp[0]) ? 4'b1100 : 4'b1110;
												assign node33945 = (inp[5]) ? node33963 : node33946;
													assign node33946 = (inp[15]) ? node33956 : node33947;
														assign node33947 = (inp[0]) ? 4'b1010 : node33948;
															assign node33948 = (inp[9]) ? node33952 : node33949;
																assign node33949 = (inp[4]) ? 4'b1100 : 4'b1010;
																assign node33952 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node33956 = (inp[0]) ? 4'b1100 : node33957;
															assign node33957 = (inp[4]) ? node33959 : 4'b1110;
																assign node33959 = (inp[9]) ? 4'b1010 : 4'b1110;
													assign node33963 = (inp[9]) ? node33975 : node33964;
														assign node33964 = (inp[4]) ? node33972 : node33965;
															assign node33965 = (inp[0]) ? node33969 : node33966;
																assign node33966 = (inp[15]) ? 4'b1010 : 4'b1000;
																assign node33969 = (inp[15]) ? 4'b1000 : 4'b1010;
															assign node33972 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node33975 = (inp[4]) ? node33983 : node33976;
															assign node33976 = (inp[0]) ? node33980 : node33977;
																assign node33977 = (inp[15]) ? 4'b1110 : 4'b1100;
																assign node33980 = (inp[15]) ? 4'b1100 : 4'b1110;
															assign node33983 = (inp[15]) ? 4'b1000 : 4'b1010;
								assign node33986 = (inp[14]) ? node34296 : node33987;
									assign node33987 = (inp[2]) ? node34141 : node33988;
										assign node33988 = (inp[9]) ? node34064 : node33989;
											assign node33989 = (inp[3]) ? node34029 : node33990;
												assign node33990 = (inp[12]) ? node34010 : node33991;
													assign node33991 = (inp[4]) ? node33999 : node33992;
														assign node33992 = (inp[0]) ? node33996 : node33993;
															assign node33993 = (inp[15]) ? 4'b1100 : 4'b1110;
															assign node33996 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node33999 = (inp[5]) ? node34005 : node34000;
															assign node34000 = (inp[15]) ? 4'b1010 : node34001;
																assign node34001 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node34005 = (inp[15]) ? 4'b1000 : node34006;
																assign node34006 = (inp[0]) ? 4'b1000 : 4'b1010;
													assign node34010 = (inp[4]) ? node34020 : node34011;
														assign node34011 = (inp[5]) ? 4'b1010 : node34012;
															assign node34012 = (inp[15]) ? node34016 : node34013;
																assign node34013 = (inp[0]) ? 4'b1000 : 4'b1010;
																assign node34016 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node34020 = (inp[15]) ? 4'b1110 : node34021;
															assign node34021 = (inp[5]) ? node34025 : node34022;
																assign node34022 = (inp[0]) ? 4'b1100 : 4'b1110;
																assign node34025 = (inp[0]) ? 4'b1110 : 4'b1100;
												assign node34029 = (inp[15]) ? node34047 : node34030;
													assign node34030 = (inp[4]) ? node34040 : node34031;
														assign node34031 = (inp[12]) ? node34035 : node34032;
															assign node34032 = (inp[5]) ? 4'b1110 : 4'b1100;
															assign node34035 = (inp[5]) ? 4'b1000 : node34036;
																assign node34036 = (inp[0]) ? 4'b1000 : 4'b1010;
														assign node34040 = (inp[12]) ? 4'b1100 : node34041;
															assign node34041 = (inp[0]) ? node34043 : 4'b1000;
																assign node34043 = (inp[5]) ? 4'b1010 : 4'b1000;
													assign node34047 = (inp[4]) ? node34053 : node34048;
														assign node34048 = (inp[12]) ? 4'b1000 : node34049;
															assign node34049 = (inp[5]) ? 4'b1100 : 4'b1110;
														assign node34053 = (inp[12]) ? node34061 : node34054;
															assign node34054 = (inp[5]) ? node34058 : node34055;
																assign node34055 = (inp[0]) ? 4'b1010 : 4'b1000;
																assign node34058 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node34061 = (inp[0]) ? 4'b1100 : 4'b1110;
											assign node34064 = (inp[15]) ? node34100 : node34065;
												assign node34065 = (inp[0]) ? node34085 : node34066;
													assign node34066 = (inp[3]) ? node34078 : node34067;
														assign node34067 = (inp[5]) ? node34073 : node34068;
															assign node34068 = (inp[12]) ? node34070 : 4'b1010;
																assign node34070 = (inp[4]) ? 4'b1010 : 4'b1110;
															assign node34073 = (inp[12]) ? 4'b1100 : node34074;
																assign node34074 = (inp[4]) ? 4'b1100 : 4'b1010;
														assign node34078 = (inp[4]) ? 4'b1100 : node34079;
															assign node34079 = (inp[12]) ? 4'b1100 : node34080;
																assign node34080 = (inp[5]) ? 4'b1000 : 4'b1010;
													assign node34085 = (inp[5]) ? node34093 : node34086;
														assign node34086 = (inp[4]) ? node34090 : node34087;
															assign node34087 = (inp[3]) ? 4'b1000 : 4'b1100;
															assign node34090 = (inp[12]) ? 4'b1010 : 4'b1110;
														assign node34093 = (inp[4]) ? node34097 : node34094;
															assign node34094 = (inp[12]) ? 4'b1110 : 4'b1010;
															assign node34097 = (inp[12]) ? 4'b1010 : 4'b1110;
												assign node34100 = (inp[0]) ? node34124 : node34101;
													assign node34101 = (inp[3]) ? node34111 : node34102;
														assign node34102 = (inp[12]) ? node34106 : node34103;
															assign node34103 = (inp[4]) ? 4'b1100 : 4'b1000;
															assign node34106 = (inp[5]) ? node34108 : 4'b1100;
																assign node34108 = (inp[4]) ? 4'b1010 : 4'b1110;
														assign node34111 = (inp[5]) ? node34119 : node34112;
															assign node34112 = (inp[4]) ? node34116 : node34113;
																assign node34113 = (inp[12]) ? 4'b1110 : 4'b1000;
																assign node34116 = (inp[12]) ? 4'b1010 : 4'b1110;
															assign node34119 = (inp[12]) ? 4'b1110 : node34120;
																assign node34120 = (inp[4]) ? 4'b1110 : 4'b1010;
													assign node34124 = (inp[5]) ? node34136 : node34125;
														assign node34125 = (inp[3]) ? node34133 : node34126;
															assign node34126 = (inp[12]) ? node34130 : node34127;
																assign node34127 = (inp[4]) ? 4'b1110 : 4'b1010;
																assign node34130 = (inp[4]) ? 4'b1010 : 4'b1110;
															assign node34133 = (inp[4]) ? 4'b1000 : 4'b1010;
														assign node34136 = (inp[12]) ? 4'b1000 : node34137;
															assign node34137 = (inp[4]) ? 4'b1100 : 4'b1000;
										assign node34141 = (inp[5]) ? node34223 : node34142;
											assign node34142 = (inp[12]) ? node34184 : node34143;
												assign node34143 = (inp[3]) ? node34165 : node34144;
													assign node34144 = (inp[9]) ? node34154 : node34145;
														assign node34145 = (inp[4]) ? node34151 : node34146;
															assign node34146 = (inp[15]) ? node34148 : 4'b0101;
																assign node34148 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node34151 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node34154 = (inp[4]) ? node34160 : node34155;
															assign node34155 = (inp[0]) ? 4'b0001 : node34156;
																assign node34156 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node34160 = (inp[15]) ? 4'b0101 : node34161;
																assign node34161 = (inp[0]) ? 4'b0101 : 4'b0111;
													assign node34165 = (inp[15]) ? node34175 : node34166;
														assign node34166 = (inp[0]) ? node34172 : node34167;
															assign node34167 = (inp[4]) ? node34169 : 4'b0011;
																assign node34169 = (inp[9]) ? 4'b0101 : 4'b0011;
															assign node34172 = (inp[4]) ? 4'b0001 : 4'b0101;
														assign node34175 = (inp[0]) ? node34181 : node34176;
															assign node34176 = (inp[9]) ? 4'b0001 : node34177;
																assign node34177 = (inp[4]) ? 4'b0001 : 4'b0101;
															assign node34181 = (inp[9]) ? 4'b0101 : 4'b0011;
												assign node34184 = (inp[4]) ? node34202 : node34185;
													assign node34185 = (inp[9]) ? node34193 : node34186;
														assign node34186 = (inp[0]) ? node34190 : node34187;
															assign node34187 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node34190 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node34193 = (inp[0]) ? 4'b0111 : node34194;
															assign node34194 = (inp[15]) ? node34198 : node34195;
																assign node34195 = (inp[3]) ? 4'b0101 : 4'b0111;
																assign node34198 = (inp[3]) ? 4'b0111 : 4'b0101;
													assign node34202 = (inp[9]) ? node34216 : node34203;
														assign node34203 = (inp[15]) ? node34209 : node34204;
															assign node34204 = (inp[3]) ? node34206 : 4'b0101;
																assign node34206 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node34209 = (inp[3]) ? node34213 : node34210;
																assign node34210 = (inp[0]) ? 4'b0111 : 4'b0101;
																assign node34213 = (inp[0]) ? 4'b0101 : 4'b0111;
														assign node34216 = (inp[0]) ? 4'b0011 : node34217;
															assign node34217 = (inp[15]) ? node34219 : 4'b0001;
																assign node34219 = (inp[3]) ? 4'b0011 : 4'b0001;
											assign node34223 = (inp[3]) ? node34259 : node34224;
												assign node34224 = (inp[4]) ? node34244 : node34225;
													assign node34225 = (inp[0]) ? node34233 : node34226;
														assign node34226 = (inp[15]) ? node34230 : node34227;
															assign node34227 = (inp[9]) ? 4'b0101 : 4'b0111;
															assign node34230 = (inp[9]) ? 4'b0111 : 4'b0101;
														assign node34233 = (inp[15]) ? node34237 : node34234;
															assign node34234 = (inp[12]) ? 4'b0111 : 4'b0101;
															assign node34237 = (inp[9]) ? node34241 : node34238;
																assign node34238 = (inp[12]) ? 4'b0011 : 4'b0111;
																assign node34241 = (inp[12]) ? 4'b0101 : 4'b0011;
													assign node34244 = (inp[15]) ? node34256 : node34245;
														assign node34245 = (inp[0]) ? node34249 : node34246;
															assign node34246 = (inp[12]) ? 4'b0001 : 4'b0011;
															assign node34249 = (inp[12]) ? node34253 : node34250;
																assign node34250 = (inp[9]) ? 4'b0111 : 4'b0001;
																assign node34253 = (inp[9]) ? 4'b0011 : 4'b0111;
														assign node34256 = (inp[12]) ? 4'b0101 : 4'b0111;
												assign node34259 = (inp[0]) ? node34281 : node34260;
													assign node34260 = (inp[15]) ? node34274 : node34261;
														assign node34261 = (inp[4]) ? node34269 : node34262;
															assign node34262 = (inp[12]) ? node34266 : node34263;
																assign node34263 = (inp[9]) ? 4'b0001 : 4'b0101;
																assign node34266 = (inp[9]) ? 4'b0101 : 4'b0001;
															assign node34269 = (inp[9]) ? 4'b0101 : node34270;
																assign node34270 = (inp[12]) ? 4'b0101 : 4'b0001;
														assign node34274 = (inp[12]) ? node34276 : 4'b0111;
															assign node34276 = (inp[9]) ? 4'b0111 : node34277;
																assign node34277 = (inp[4]) ? 4'b0111 : 4'b0011;
													assign node34281 = (inp[15]) ? node34289 : node34282;
														assign node34282 = (inp[9]) ? node34284 : 4'b0111;
															assign node34284 = (inp[12]) ? 4'b0011 : node34285;
																assign node34285 = (inp[4]) ? 4'b0111 : 4'b0011;
														assign node34289 = (inp[9]) ? node34291 : 4'b0001;
															assign node34291 = (inp[4]) ? 4'b0001 : node34292;
																assign node34292 = (inp[12]) ? 4'b0101 : 4'b0001;
									assign node34296 = (inp[0]) ? node34406 : node34297;
										assign node34297 = (inp[12]) ? node34353 : node34298;
											assign node34298 = (inp[15]) ? node34330 : node34299;
												assign node34299 = (inp[3]) ? node34315 : node34300;
													assign node34300 = (inp[5]) ? node34308 : node34301;
														assign node34301 = (inp[9]) ? node34305 : node34302;
															assign node34302 = (inp[4]) ? 4'b0011 : 4'b0111;
															assign node34305 = (inp[4]) ? 4'b0111 : 4'b0011;
														assign node34308 = (inp[4]) ? node34312 : node34309;
															assign node34309 = (inp[9]) ? 4'b0011 : 4'b0111;
															assign node34312 = (inp[9]) ? 4'b0101 : 4'b0011;
													assign node34315 = (inp[5]) ? node34323 : node34316;
														assign node34316 = (inp[9]) ? node34320 : node34317;
															assign node34317 = (inp[4]) ? 4'b0011 : 4'b0111;
															assign node34320 = (inp[4]) ? 4'b0101 : 4'b0011;
														assign node34323 = (inp[4]) ? node34327 : node34324;
															assign node34324 = (inp[9]) ? 4'b0001 : 4'b0101;
															assign node34327 = (inp[9]) ? 4'b0101 : 4'b0001;
												assign node34330 = (inp[3]) ? node34340 : node34331;
													assign node34331 = (inp[9]) ? node34335 : node34332;
														assign node34332 = (inp[4]) ? 4'b0001 : 4'b0101;
														assign node34335 = (inp[4]) ? node34337 : 4'b0001;
															assign node34337 = (inp[5]) ? 4'b0111 : 4'b0101;
													assign node34340 = (inp[5]) ? node34346 : node34341;
														assign node34341 = (inp[4]) ? node34343 : 4'b0001;
															assign node34343 = (inp[9]) ? 4'b0111 : 4'b0001;
														assign node34346 = (inp[4]) ? node34350 : node34347;
															assign node34347 = (inp[9]) ? 4'b0011 : 4'b0111;
															assign node34350 = (inp[9]) ? 4'b0111 : 4'b0011;
											assign node34353 = (inp[15]) ? node34373 : node34354;
												assign node34354 = (inp[5]) ? node34364 : node34355;
													assign node34355 = (inp[9]) ? node34357 : 4'b0011;
														assign node34357 = (inp[4]) ? node34361 : node34358;
															assign node34358 = (inp[3]) ? 4'b0101 : 4'b0111;
															assign node34361 = (inp[3]) ? 4'b0001 : 4'b0011;
													assign node34364 = (inp[9]) ? node34370 : node34365;
														assign node34365 = (inp[4]) ? 4'b0101 : node34366;
															assign node34366 = (inp[2]) ? 4'b0001 : 4'b0011;
														assign node34370 = (inp[4]) ? 4'b0001 : 4'b0101;
												assign node34373 = (inp[5]) ? node34389 : node34374;
													assign node34374 = (inp[3]) ? node34382 : node34375;
														assign node34375 = (inp[2]) ? 4'b0101 : node34376;
															assign node34376 = (inp[4]) ? node34378 : 4'b0001;
																assign node34378 = (inp[9]) ? 4'b0001 : 4'b0101;
														assign node34382 = (inp[9]) ? node34386 : node34383;
															assign node34383 = (inp[4]) ? 4'b0111 : 4'b0001;
															assign node34386 = (inp[4]) ? 4'b0011 : 4'b0111;
													assign node34389 = (inp[3]) ? node34399 : node34390;
														assign node34390 = (inp[2]) ? 4'b0111 : node34391;
															assign node34391 = (inp[4]) ? node34395 : node34392;
																assign node34392 = (inp[9]) ? 4'b0111 : 4'b0001;
																assign node34395 = (inp[9]) ? 4'b0011 : 4'b0111;
														assign node34399 = (inp[2]) ? node34401 : 4'b0011;
															assign node34401 = (inp[4]) ? node34403 : 4'b0011;
																assign node34403 = (inp[9]) ? 4'b0011 : 4'b0111;
										assign node34406 = (inp[2]) ? node34474 : node34407;
											assign node34407 = (inp[15]) ? node34445 : node34408;
												assign node34408 = (inp[5]) ? node34428 : node34409;
													assign node34409 = (inp[4]) ? node34419 : node34410;
														assign node34410 = (inp[3]) ? 4'b0001 : node34411;
															assign node34411 = (inp[9]) ? node34415 : node34412;
																assign node34412 = (inp[12]) ? 4'b0001 : 4'b0101;
																assign node34415 = (inp[12]) ? 4'b0101 : 4'b0001;
														assign node34419 = (inp[3]) ? 4'b0111 : node34420;
															assign node34420 = (inp[9]) ? node34424 : node34421;
																assign node34421 = (inp[12]) ? 4'b0101 : 4'b0001;
																assign node34424 = (inp[12]) ? 4'b0001 : 4'b0101;
													assign node34428 = (inp[3]) ? 4'b0111 : node34429;
														assign node34429 = (inp[9]) ? node34437 : node34430;
															assign node34430 = (inp[4]) ? node34434 : node34431;
																assign node34431 = (inp[12]) ? 4'b0001 : 4'b0101;
																assign node34434 = (inp[12]) ? 4'b0111 : 4'b0001;
															assign node34437 = (inp[12]) ? node34441 : node34438;
																assign node34438 = (inp[4]) ? 4'b0111 : 4'b0001;
																assign node34441 = (inp[4]) ? 4'b0011 : 4'b0111;
												assign node34445 = (inp[5]) ? node34463 : node34446;
													assign node34446 = (inp[3]) ? node34454 : node34447;
														assign node34447 = (inp[4]) ? node34449 : 4'b0111;
															assign node34449 = (inp[12]) ? 4'b0011 : node34450;
																assign node34450 = (inp[9]) ? 4'b0111 : 4'b0011;
														assign node34454 = (inp[12]) ? 4'b0101 : node34455;
															assign node34455 = (inp[4]) ? node34459 : node34456;
																assign node34456 = (inp[9]) ? 4'b0011 : 4'b0111;
																assign node34459 = (inp[9]) ? 4'b0101 : 4'b0011;
													assign node34463 = (inp[12]) ? node34469 : node34464;
														assign node34464 = (inp[4]) ? 4'b0101 : node34465;
															assign node34465 = (inp[3]) ? 4'b0101 : 4'b0111;
														assign node34469 = (inp[4]) ? 4'b0101 : node34470;
															assign node34470 = (inp[9]) ? 4'b0101 : 4'b0001;
											assign node34474 = (inp[5]) ? node34514 : node34475;
												assign node34475 = (inp[15]) ? node34489 : node34476;
													assign node34476 = (inp[3]) ? node34484 : node34477;
														assign node34477 = (inp[4]) ? node34479 : 4'b0101;
															assign node34479 = (inp[12]) ? 4'b0001 : node34480;
																assign node34480 = (inp[9]) ? 4'b0101 : 4'b0001;
														assign node34484 = (inp[4]) ? node34486 : 4'b0001;
															assign node34486 = (inp[12]) ? 4'b0011 : 4'b0111;
													assign node34489 = (inp[3]) ? node34503 : node34490;
														assign node34490 = (inp[9]) ? node34496 : node34491;
															assign node34491 = (inp[12]) ? 4'b0011 : node34492;
																assign node34492 = (inp[4]) ? 4'b0011 : 4'b0111;
															assign node34496 = (inp[4]) ? node34500 : node34497;
																assign node34497 = (inp[12]) ? 4'b0111 : 4'b0011;
																assign node34500 = (inp[12]) ? 4'b0011 : 4'b0111;
														assign node34503 = (inp[12]) ? node34509 : node34504;
															assign node34504 = (inp[4]) ? node34506 : 4'b0011;
																assign node34506 = (inp[9]) ? 4'b0101 : 4'b0011;
															assign node34509 = (inp[9]) ? node34511 : 4'b0101;
																assign node34511 = (inp[4]) ? 4'b0001 : 4'b0101;
												assign node34514 = (inp[15]) ? node34530 : node34515;
													assign node34515 = (inp[3]) ? node34523 : node34516;
														assign node34516 = (inp[12]) ? 4'b0111 : node34517;
															assign node34517 = (inp[9]) ? 4'b0001 : node34518;
																assign node34518 = (inp[4]) ? 4'b0001 : 4'b0101;
														assign node34523 = (inp[4]) ? 4'b0011 : node34524;
															assign node34524 = (inp[12]) ? 4'b0011 : node34525;
																assign node34525 = (inp[9]) ? 4'b0011 : 4'b0111;
													assign node34530 = (inp[3]) ? node34542 : node34531;
														assign node34531 = (inp[4]) ? node34537 : node34532;
															assign node34532 = (inp[12]) ? node34534 : 4'b0011;
																assign node34534 = (inp[9]) ? 4'b0101 : 4'b0011;
															assign node34537 = (inp[9]) ? node34539 : 4'b0101;
																assign node34539 = (inp[12]) ? 4'b0001 : 4'b0101;
														assign node34542 = (inp[12]) ? 4'b0001 : node34543;
															assign node34543 = (inp[9]) ? node34547 : node34544;
																assign node34544 = (inp[4]) ? 4'b0001 : 4'b0101;
																assign node34547 = (inp[4]) ? 4'b0101 : 4'b0001;
							assign node34551 = (inp[8]) ? node35051 : node34552;
								assign node34552 = (inp[2]) ? node34814 : node34553;
									assign node34553 = (inp[14]) ? node34683 : node34554;
										assign node34554 = (inp[12]) ? node34622 : node34555;
											assign node34555 = (inp[5]) ? node34593 : node34556;
												assign node34556 = (inp[9]) ? node34572 : node34557;
													assign node34557 = (inp[4]) ? node34565 : node34558;
														assign node34558 = (inp[0]) ? node34562 : node34559;
															assign node34559 = (inp[15]) ? 4'b1100 : 4'b1110;
															assign node34562 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node34565 = (inp[3]) ? node34567 : 4'b1000;
															assign node34567 = (inp[0]) ? 4'b1010 : node34568;
																assign node34568 = (inp[15]) ? 4'b1000 : 4'b1010;
													assign node34572 = (inp[4]) ? node34580 : node34573;
														assign node34573 = (inp[0]) ? node34577 : node34574;
															assign node34574 = (inp[15]) ? 4'b1000 : 4'b1010;
															assign node34577 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node34580 = (inp[0]) ? node34586 : node34581;
															assign node34581 = (inp[15]) ? 4'b1100 : node34582;
																assign node34582 = (inp[3]) ? 4'b1100 : 4'b1110;
															assign node34586 = (inp[3]) ? node34590 : node34587;
																assign node34587 = (inp[15]) ? 4'b1110 : 4'b1100;
																assign node34590 = (inp[15]) ? 4'b1100 : 4'b1110;
												assign node34593 = (inp[9]) ? node34607 : node34594;
													assign node34594 = (inp[4]) ? node34598 : node34595;
														assign node34595 = (inp[15]) ? 4'b1100 : 4'b1110;
														assign node34598 = (inp[15]) ? 4'b1010 : node34599;
															assign node34599 = (inp[0]) ? node34603 : node34600;
																assign node34600 = (inp[3]) ? 4'b1000 : 4'b1010;
																assign node34603 = (inp[3]) ? 4'b1010 : 4'b1000;
													assign node34607 = (inp[4]) ? node34613 : node34608;
														assign node34608 = (inp[0]) ? node34610 : 4'b1010;
															assign node34610 = (inp[3]) ? 4'b1010 : 4'b1000;
														assign node34613 = (inp[3]) ? 4'b1110 : node34614;
															assign node34614 = (inp[0]) ? node34618 : node34615;
																assign node34615 = (inp[15]) ? 4'b1110 : 4'b1100;
																assign node34618 = (inp[15]) ? 4'b1100 : 4'b1110;
											assign node34622 = (inp[4]) ? node34652 : node34623;
												assign node34623 = (inp[9]) ? node34643 : node34624;
													assign node34624 = (inp[5]) ? node34630 : node34625;
														assign node34625 = (inp[15]) ? node34627 : 4'b1000;
															assign node34627 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node34630 = (inp[0]) ? node34638 : node34631;
															assign node34631 = (inp[3]) ? node34635 : node34632;
																assign node34632 = (inp[15]) ? 4'b1000 : 4'b1010;
																assign node34635 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node34638 = (inp[15]) ? node34640 : 4'b1010;
																assign node34640 = (inp[3]) ? 4'b1000 : 4'b1010;
													assign node34643 = (inp[5]) ? node34647 : node34644;
														assign node34644 = (inp[3]) ? 4'b1100 : 4'b1110;
														assign node34647 = (inp[3]) ? node34649 : 4'b1100;
															assign node34649 = (inp[0]) ? 4'b1110 : 4'b1100;
												assign node34652 = (inp[9]) ? node34672 : node34653;
													assign node34653 = (inp[5]) ? node34663 : node34654;
														assign node34654 = (inp[0]) ? node34656 : 4'b1110;
															assign node34656 = (inp[3]) ? node34660 : node34657;
																assign node34657 = (inp[15]) ? 4'b1110 : 4'b1100;
																assign node34660 = (inp[15]) ? 4'b1100 : 4'b1110;
														assign node34663 = (inp[3]) ? node34665 : 4'b1100;
															assign node34665 = (inp[15]) ? node34669 : node34666;
																assign node34666 = (inp[0]) ? 4'b1110 : 4'b1100;
																assign node34669 = (inp[0]) ? 4'b1100 : 4'b1110;
													assign node34672 = (inp[0]) ? node34678 : node34673;
														assign node34673 = (inp[15]) ? 4'b1010 : node34674;
															assign node34674 = (inp[3]) ? 4'b1000 : 4'b1010;
														assign node34678 = (inp[3]) ? node34680 : 4'b1000;
															assign node34680 = (inp[15]) ? 4'b1000 : 4'b1010;
										assign node34683 = (inp[9]) ? node34755 : node34684;
											assign node34684 = (inp[15]) ? node34712 : node34685;
												assign node34685 = (inp[0]) ? node34699 : node34686;
													assign node34686 = (inp[3]) ? node34696 : node34687;
														assign node34687 = (inp[4]) ? node34691 : node34688;
															assign node34688 = (inp[12]) ? 4'b0011 : 4'b0111;
															assign node34691 = (inp[12]) ? node34693 : 4'b0011;
																assign node34693 = (inp[5]) ? 4'b0101 : 4'b0111;
														assign node34696 = (inp[5]) ? 4'b0101 : 4'b0111;
													assign node34699 = (inp[5]) ? node34709 : node34700;
														assign node34700 = (inp[4]) ? node34704 : node34701;
															assign node34701 = (inp[12]) ? 4'b0001 : 4'b0101;
															assign node34704 = (inp[12]) ? node34706 : 4'b0001;
																assign node34706 = (inp[3]) ? 4'b0111 : 4'b0101;
														assign node34709 = (inp[3]) ? 4'b0111 : 4'b0101;
												assign node34712 = (inp[0]) ? node34728 : node34713;
													assign node34713 = (inp[3]) ? node34721 : node34714;
														assign node34714 = (inp[12]) ? node34718 : node34715;
															assign node34715 = (inp[4]) ? 4'b0001 : 4'b0101;
															assign node34718 = (inp[4]) ? 4'b0111 : 4'b0001;
														assign node34721 = (inp[4]) ? node34725 : node34722;
															assign node34722 = (inp[5]) ? 4'b0011 : 4'b0001;
															assign node34725 = (inp[12]) ? 4'b0111 : 4'b0011;
													assign node34728 = (inp[3]) ? node34742 : node34729;
														assign node34729 = (inp[5]) ? node34737 : node34730;
															assign node34730 = (inp[12]) ? node34734 : node34731;
																assign node34731 = (inp[4]) ? 4'b0011 : 4'b0111;
																assign node34734 = (inp[4]) ? 4'b0111 : 4'b0011;
															assign node34737 = (inp[4]) ? 4'b0011 : node34738;
																assign node34738 = (inp[12]) ? 4'b0011 : 4'b0111;
														assign node34742 = (inp[5]) ? node34750 : node34743;
															assign node34743 = (inp[4]) ? node34747 : node34744;
																assign node34744 = (inp[12]) ? 4'b0011 : 4'b0111;
																assign node34747 = (inp[12]) ? 4'b0101 : 4'b0011;
															assign node34750 = (inp[4]) ? 4'b0101 : node34751;
																assign node34751 = (inp[12]) ? 4'b0001 : 4'b0101;
											assign node34755 = (inp[15]) ? node34781 : node34756;
												assign node34756 = (inp[4]) ? node34768 : node34757;
													assign node34757 = (inp[12]) ? node34761 : node34758;
														assign node34758 = (inp[0]) ? 4'b0001 : 4'b0011;
														assign node34761 = (inp[0]) ? node34763 : 4'b0101;
															assign node34763 = (inp[5]) ? 4'b0111 : node34764;
																assign node34764 = (inp[3]) ? 4'b0111 : 4'b0101;
													assign node34768 = (inp[12]) ? node34772 : node34769;
														assign node34769 = (inp[5]) ? 4'b0111 : 4'b0101;
														assign node34772 = (inp[0]) ? node34778 : node34773;
															assign node34773 = (inp[3]) ? 4'b0001 : node34774;
																assign node34774 = (inp[5]) ? 4'b0001 : 4'b0011;
															assign node34778 = (inp[5]) ? 4'b0011 : 4'b0001;
												assign node34781 = (inp[0]) ? node34799 : node34782;
													assign node34782 = (inp[3]) ? node34790 : node34783;
														assign node34783 = (inp[5]) ? 4'b0011 : node34784;
															assign node34784 = (inp[4]) ? 4'b0001 : node34785;
																assign node34785 = (inp[12]) ? 4'b0101 : 4'b0001;
														assign node34790 = (inp[5]) ? node34792 : 4'b0111;
															assign node34792 = (inp[12]) ? node34796 : node34793;
																assign node34793 = (inp[4]) ? 4'b0111 : 4'b0011;
																assign node34796 = (inp[4]) ? 4'b0011 : 4'b0111;
													assign node34799 = (inp[4]) ? node34807 : node34800;
														assign node34800 = (inp[12]) ? node34802 : 4'b0011;
															assign node34802 = (inp[3]) ? 4'b0101 : node34803;
																assign node34803 = (inp[5]) ? 4'b0101 : 4'b0111;
														assign node34807 = (inp[12]) ? 4'b0001 : node34808;
															assign node34808 = (inp[3]) ? 4'b0101 : node34809;
																assign node34809 = (inp[5]) ? 4'b0101 : 4'b0111;
									assign node34814 = (inp[15]) ? node34920 : node34815;
										assign node34815 = (inp[12]) ? node34871 : node34816;
											assign node34816 = (inp[0]) ? node34842 : node34817;
												assign node34817 = (inp[5]) ? node34827 : node34818;
													assign node34818 = (inp[4]) ? node34822 : node34819;
														assign node34819 = (inp[9]) ? 4'b0011 : 4'b0111;
														assign node34822 = (inp[9]) ? node34824 : 4'b0011;
															assign node34824 = (inp[3]) ? 4'b0101 : 4'b0111;
													assign node34827 = (inp[3]) ? node34835 : node34828;
														assign node34828 = (inp[9]) ? node34832 : node34829;
															assign node34829 = (inp[4]) ? 4'b0011 : 4'b0111;
															assign node34832 = (inp[4]) ? 4'b0101 : 4'b0011;
														assign node34835 = (inp[9]) ? node34839 : node34836;
															assign node34836 = (inp[4]) ? 4'b0001 : 4'b0101;
															assign node34839 = (inp[4]) ? 4'b0101 : 4'b0001;
												assign node34842 = (inp[5]) ? node34862 : node34843;
													assign node34843 = (inp[14]) ? node34855 : node34844;
														assign node34844 = (inp[3]) ? node34850 : node34845;
															assign node34845 = (inp[9]) ? node34847 : 4'b0101;
																assign node34847 = (inp[4]) ? 4'b0101 : 4'b0001;
															assign node34850 = (inp[9]) ? 4'b0111 : node34851;
																assign node34851 = (inp[4]) ? 4'b0001 : 4'b0101;
														assign node34855 = (inp[4]) ? node34859 : node34856;
															assign node34856 = (inp[9]) ? 4'b0001 : 4'b0101;
															assign node34859 = (inp[9]) ? 4'b0101 : 4'b0001;
													assign node34862 = (inp[4]) ? 4'b0111 : node34863;
														assign node34863 = (inp[3]) ? node34867 : node34864;
															assign node34864 = (inp[9]) ? 4'b0001 : 4'b0101;
															assign node34867 = (inp[9]) ? 4'b0011 : 4'b0111;
											assign node34871 = (inp[0]) ? node34897 : node34872;
												assign node34872 = (inp[5]) ? node34888 : node34873;
													assign node34873 = (inp[3]) ? node34881 : node34874;
														assign node34874 = (inp[4]) ? node34878 : node34875;
															assign node34875 = (inp[9]) ? 4'b0111 : 4'b0011;
															assign node34878 = (inp[9]) ? 4'b0011 : 4'b0111;
														assign node34881 = (inp[4]) ? node34885 : node34882;
															assign node34882 = (inp[9]) ? 4'b0101 : 4'b0011;
															assign node34885 = (inp[9]) ? 4'b0001 : 4'b0101;
													assign node34888 = (inp[4]) ? node34894 : node34889;
														assign node34889 = (inp[9]) ? 4'b0101 : node34890;
															assign node34890 = (inp[3]) ? 4'b0001 : 4'b0011;
														assign node34894 = (inp[9]) ? 4'b0001 : 4'b0101;
												assign node34897 = (inp[3]) ? node34911 : node34898;
													assign node34898 = (inp[5]) ? node34904 : node34899;
														assign node34899 = (inp[4]) ? 4'b0001 : node34900;
															assign node34900 = (inp[9]) ? 4'b0101 : 4'b0001;
														assign node34904 = (inp[4]) ? node34908 : node34905;
															assign node34905 = (inp[9]) ? 4'b0111 : 4'b0001;
															assign node34908 = (inp[9]) ? 4'b0011 : 4'b0111;
													assign node34911 = (inp[9]) ? node34917 : node34912;
														assign node34912 = (inp[4]) ? 4'b0111 : node34913;
															assign node34913 = (inp[5]) ? 4'b0011 : 4'b0001;
														assign node34917 = (inp[4]) ? 4'b0011 : 4'b0111;
										assign node34920 = (inp[5]) ? node34988 : node34921;
											assign node34921 = (inp[0]) ? node34959 : node34922;
												assign node34922 = (inp[3]) ? node34944 : node34923;
													assign node34923 = (inp[14]) ? node34935 : node34924;
														assign node34924 = (inp[12]) ? node34930 : node34925;
															assign node34925 = (inp[9]) ? 4'b0001 : node34926;
																assign node34926 = (inp[4]) ? 4'b0001 : 4'b0101;
															assign node34930 = (inp[9]) ? 4'b0101 : node34931;
																assign node34931 = (inp[4]) ? 4'b0101 : 4'b0001;
														assign node34935 = (inp[12]) ? node34937 : 4'b0101;
															assign node34937 = (inp[4]) ? node34941 : node34938;
																assign node34938 = (inp[9]) ? 4'b0101 : 4'b0001;
																assign node34941 = (inp[9]) ? 4'b0001 : 4'b0101;
													assign node34944 = (inp[12]) ? node34952 : node34945;
														assign node34945 = (inp[4]) ? node34949 : node34946;
															assign node34946 = (inp[9]) ? 4'b0001 : 4'b0101;
															assign node34949 = (inp[9]) ? 4'b0111 : 4'b0001;
														assign node34952 = (inp[9]) ? node34956 : node34953;
															assign node34953 = (inp[4]) ? 4'b0111 : 4'b0001;
															assign node34956 = (inp[4]) ? 4'b0011 : 4'b0111;
												assign node34959 = (inp[3]) ? node34973 : node34960;
													assign node34960 = (inp[12]) ? node34968 : node34961;
														assign node34961 = (inp[9]) ? node34965 : node34962;
															assign node34962 = (inp[4]) ? 4'b0011 : 4'b0111;
															assign node34965 = (inp[4]) ? 4'b0111 : 4'b0011;
														assign node34968 = (inp[9]) ? node34970 : 4'b0011;
															assign node34970 = (inp[4]) ? 4'b0011 : 4'b0111;
													assign node34973 = (inp[4]) ? node34981 : node34974;
														assign node34974 = (inp[9]) ? node34978 : node34975;
															assign node34975 = (inp[12]) ? 4'b0011 : 4'b0111;
															assign node34978 = (inp[12]) ? 4'b0101 : 4'b0011;
														assign node34981 = (inp[12]) ? node34985 : node34982;
															assign node34982 = (inp[9]) ? 4'b0101 : 4'b0011;
															assign node34985 = (inp[9]) ? 4'b0001 : 4'b0101;
											assign node34988 = (inp[0]) ? node35020 : node34989;
												assign node34989 = (inp[3]) ? node35005 : node34990;
													assign node34990 = (inp[9]) ? node34998 : node34991;
														assign node34991 = (inp[12]) ? node34995 : node34992;
															assign node34992 = (inp[4]) ? 4'b0001 : 4'b0101;
															assign node34995 = (inp[4]) ? 4'b0111 : 4'b0001;
														assign node34998 = (inp[4]) ? node35002 : node34999;
															assign node34999 = (inp[12]) ? 4'b0111 : 4'b0001;
															assign node35002 = (inp[12]) ? 4'b0011 : 4'b0111;
													assign node35005 = (inp[9]) ? node35013 : node35006;
														assign node35006 = (inp[12]) ? node35010 : node35007;
															assign node35007 = (inp[4]) ? 4'b0011 : 4'b0111;
															assign node35010 = (inp[4]) ? 4'b0111 : 4'b0011;
														assign node35013 = (inp[12]) ? node35017 : node35014;
															assign node35014 = (inp[4]) ? 4'b0111 : 4'b0011;
															assign node35017 = (inp[4]) ? 4'b0011 : 4'b0111;
												assign node35020 = (inp[3]) ? node35032 : node35021;
													assign node35021 = (inp[9]) ? node35027 : node35022;
														assign node35022 = (inp[12]) ? 4'b0011 : node35023;
															assign node35023 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node35027 = (inp[14]) ? 4'b0011 : node35028;
															assign node35028 = (inp[4]) ? 4'b0001 : 4'b0101;
													assign node35032 = (inp[12]) ? node35038 : node35033;
														assign node35033 = (inp[4]) ? 4'b0101 : node35034;
															assign node35034 = (inp[9]) ? 4'b0001 : 4'b0101;
														assign node35038 = (inp[14]) ? node35046 : node35039;
															assign node35039 = (inp[4]) ? node35043 : node35040;
																assign node35040 = (inp[9]) ? 4'b0101 : 4'b0001;
																assign node35043 = (inp[9]) ? 4'b0001 : 4'b0101;
															assign node35046 = (inp[4]) ? node35048 : 4'b0001;
																assign node35048 = (inp[9]) ? 4'b0001 : 4'b0101;
								assign node35051 = (inp[2]) ? node35317 : node35052;
									assign node35052 = (inp[14]) ? node35182 : node35053;
										assign node35053 = (inp[3]) ? node35123 : node35054;
											assign node35054 = (inp[4]) ? node35092 : node35055;
												assign node35055 = (inp[5]) ? node35077 : node35056;
													assign node35056 = (inp[9]) ? node35064 : node35057;
														assign node35057 = (inp[12]) ? node35059 : 4'b0101;
															assign node35059 = (inp[15]) ? node35061 : 4'b0001;
																assign node35061 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node35064 = (inp[12]) ? node35070 : node35065;
															assign node35065 = (inp[0]) ? 4'b0001 : node35066;
																assign node35066 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node35070 = (inp[0]) ? node35074 : node35071;
																assign node35071 = (inp[15]) ? 4'b0101 : 4'b0111;
																assign node35074 = (inp[15]) ? 4'b0111 : 4'b0101;
													assign node35077 = (inp[15]) ? node35087 : node35078;
														assign node35078 = (inp[0]) ? node35084 : node35079;
															assign node35079 = (inp[12]) ? 4'b0101 : node35080;
																assign node35080 = (inp[9]) ? 4'b0011 : 4'b0111;
															assign node35084 = (inp[9]) ? 4'b0111 : 4'b0101;
														assign node35087 = (inp[12]) ? 4'b0101 : node35088;
															assign node35088 = (inp[0]) ? 4'b0111 : 4'b0101;
												assign node35092 = (inp[15]) ? node35106 : node35093;
													assign node35093 = (inp[9]) ? node35097 : node35094;
														assign node35094 = (inp[12]) ? 4'b0101 : 4'b0001;
														assign node35097 = (inp[12]) ? node35103 : node35098;
															assign node35098 = (inp[5]) ? node35100 : 4'b0101;
																assign node35100 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node35103 = (inp[0]) ? 4'b0001 : 4'b0011;
													assign node35106 = (inp[0]) ? node35114 : node35107;
														assign node35107 = (inp[12]) ? node35111 : node35108;
															assign node35108 = (inp[9]) ? 4'b0101 : 4'b0001;
															assign node35111 = (inp[9]) ? 4'b0011 : 4'b0111;
														assign node35114 = (inp[5]) ? 4'b0001 : node35115;
															assign node35115 = (inp[9]) ? node35119 : node35116;
																assign node35116 = (inp[12]) ? 4'b0111 : 4'b0011;
																assign node35119 = (inp[12]) ? 4'b0011 : 4'b0111;
											assign node35123 = (inp[9]) ? node35151 : node35124;
												assign node35124 = (inp[5]) ? node35140 : node35125;
													assign node35125 = (inp[0]) ? node35127 : 4'b0001;
														assign node35127 = (inp[15]) ? node35135 : node35128;
															assign node35128 = (inp[12]) ? node35132 : node35129;
																assign node35129 = (inp[4]) ? 4'b0001 : 4'b0101;
																assign node35132 = (inp[4]) ? 4'b0111 : 4'b0001;
															assign node35135 = (inp[12]) ? 4'b0011 : node35136;
																assign node35136 = (inp[4]) ? 4'b0011 : 4'b0111;
													assign node35140 = (inp[4]) ? node35144 : node35141;
														assign node35141 = (inp[12]) ? 4'b0011 : 4'b0111;
														assign node35144 = (inp[12]) ? node35146 : 4'b0011;
															assign node35146 = (inp[15]) ? 4'b0111 : node35147;
																assign node35147 = (inp[0]) ? 4'b0111 : 4'b0101;
												assign node35151 = (inp[15]) ? node35169 : node35152;
													assign node35152 = (inp[5]) ? node35162 : node35153;
														assign node35153 = (inp[0]) ? node35155 : 4'b0011;
															assign node35155 = (inp[12]) ? node35159 : node35156;
																assign node35156 = (inp[4]) ? 4'b0111 : 4'b0001;
																assign node35159 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node35162 = (inp[0]) ? 4'b0011 : node35163;
															assign node35163 = (inp[4]) ? 4'b0001 : node35164;
																assign node35164 = (inp[12]) ? 4'b0101 : 4'b0001;
													assign node35169 = (inp[0]) ? node35175 : node35170;
														assign node35170 = (inp[4]) ? node35172 : 4'b0001;
															assign node35172 = (inp[12]) ? 4'b0011 : 4'b0111;
														assign node35175 = (inp[12]) ? node35179 : node35176;
															assign node35176 = (inp[4]) ? 4'b0101 : 4'b0001;
															assign node35179 = (inp[4]) ? 4'b0001 : 4'b0101;
										assign node35182 = (inp[15]) ? node35246 : node35183;
											assign node35183 = (inp[9]) ? node35215 : node35184;
												assign node35184 = (inp[3]) ? node35200 : node35185;
													assign node35185 = (inp[0]) ? node35195 : node35186;
														assign node35186 = (inp[4]) ? node35190 : node35187;
															assign node35187 = (inp[12]) ? 4'b0010 : 4'b0110;
															assign node35190 = (inp[12]) ? node35192 : 4'b0010;
																assign node35192 = (inp[5]) ? 4'b0100 : 4'b0110;
														assign node35195 = (inp[12]) ? 4'b0110 : node35196;
															assign node35196 = (inp[5]) ? 4'b0000 : 4'b0100;
													assign node35200 = (inp[0]) ? node35208 : node35201;
														assign node35201 = (inp[12]) ? node35205 : node35202;
															assign node35202 = (inp[4]) ? 4'b0010 : 4'b0110;
															assign node35205 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node35208 = (inp[5]) ? 4'b0010 : node35209;
															assign node35209 = (inp[12]) ? 4'b0000 : node35210;
																assign node35210 = (inp[4]) ? 4'b0000 : 4'b0100;
												assign node35215 = (inp[5]) ? node35239 : node35216;
													assign node35216 = (inp[0]) ? node35228 : node35217;
														assign node35217 = (inp[3]) ? node35223 : node35218;
															assign node35218 = (inp[4]) ? 4'b0010 : node35219;
																assign node35219 = (inp[12]) ? 4'b0110 : 4'b0010;
															assign node35223 = (inp[12]) ? node35225 : 4'b0100;
																assign node35225 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node35228 = (inp[3]) ? node35234 : node35229;
															assign node35229 = (inp[12]) ? 4'b0100 : node35230;
																assign node35230 = (inp[4]) ? 4'b0100 : 4'b0000;
															assign node35234 = (inp[12]) ? 4'b0110 : node35235;
																assign node35235 = (inp[4]) ? 4'b0110 : 4'b0000;
													assign node35239 = (inp[0]) ? node35241 : 4'b0100;
														assign node35241 = (inp[4]) ? 4'b0110 : node35242;
															assign node35242 = (inp[12]) ? 4'b0110 : 4'b0010;
											assign node35246 = (inp[4]) ? node35284 : node35247;
												assign node35247 = (inp[5]) ? node35265 : node35248;
													assign node35248 = (inp[0]) ? node35256 : node35249;
														assign node35249 = (inp[3]) ? 4'b0000 : node35250;
															assign node35250 = (inp[9]) ? 4'b0000 : node35251;
																assign node35251 = (inp[12]) ? 4'b0000 : 4'b0100;
														assign node35256 = (inp[12]) ? node35260 : node35257;
															assign node35257 = (inp[3]) ? 4'b0110 : 4'b0010;
															assign node35260 = (inp[9]) ? node35262 : 4'b0010;
																assign node35262 = (inp[3]) ? 4'b0100 : 4'b0110;
													assign node35265 = (inp[0]) ? node35277 : node35266;
														assign node35266 = (inp[3]) ? node35270 : node35267;
															assign node35267 = (inp[9]) ? 4'b0110 : 4'b0100;
															assign node35270 = (inp[12]) ? node35274 : node35271;
																assign node35271 = (inp[9]) ? 4'b0010 : 4'b0110;
																assign node35274 = (inp[9]) ? 4'b0110 : 4'b0010;
														assign node35277 = (inp[12]) ? node35281 : node35278;
															assign node35278 = (inp[3]) ? 4'b0100 : 4'b0010;
															assign node35281 = (inp[9]) ? 4'b0100 : 4'b0000;
												assign node35284 = (inp[0]) ? node35300 : node35285;
													assign node35285 = (inp[3]) ? node35293 : node35286;
														assign node35286 = (inp[9]) ? node35290 : node35287;
															assign node35287 = (inp[12]) ? 4'b0100 : 4'b0000;
															assign node35290 = (inp[12]) ? 4'b0000 : 4'b0100;
														assign node35293 = (inp[12]) ? node35297 : node35294;
															assign node35294 = (inp[9]) ? 4'b0110 : 4'b0000;
															assign node35297 = (inp[9]) ? 4'b0010 : 4'b0110;
													assign node35300 = (inp[3]) ? node35310 : node35301;
														assign node35301 = (inp[5]) ? node35307 : node35302;
															assign node35302 = (inp[12]) ? node35304 : 4'b0010;
																assign node35304 = (inp[9]) ? 4'b0010 : 4'b0110;
															assign node35307 = (inp[12]) ? 4'b0000 : 4'b0010;
														assign node35310 = (inp[12]) ? node35314 : node35311;
															assign node35311 = (inp[5]) ? 4'b0000 : 4'b0010;
															assign node35314 = (inp[9]) ? 4'b0000 : 4'b0100;
									assign node35317 = (inp[14]) ? node35471 : node35318;
										assign node35318 = (inp[3]) ? node35408 : node35319;
											assign node35319 = (inp[5]) ? node35365 : node35320;
												assign node35320 = (inp[9]) ? node35348 : node35321;
													assign node35321 = (inp[0]) ? node35337 : node35322;
														assign node35322 = (inp[15]) ? node35330 : node35323;
															assign node35323 = (inp[12]) ? node35327 : node35324;
																assign node35324 = (inp[4]) ? 4'b0010 : 4'b0110;
																assign node35327 = (inp[4]) ? 4'b0110 : 4'b0010;
															assign node35330 = (inp[4]) ? node35334 : node35331;
																assign node35331 = (inp[12]) ? 4'b0000 : 4'b0100;
																assign node35334 = (inp[12]) ? 4'b0100 : 4'b0000;
														assign node35337 = (inp[15]) ? node35343 : node35338;
															assign node35338 = (inp[4]) ? node35340 : 4'b0100;
																assign node35340 = (inp[12]) ? 4'b0100 : 4'b0000;
															assign node35343 = (inp[4]) ? node35345 : 4'b0110;
																assign node35345 = (inp[12]) ? 4'b0110 : 4'b0010;
													assign node35348 = (inp[0]) ? node35358 : node35349;
														assign node35349 = (inp[15]) ? node35351 : 4'b0110;
															assign node35351 = (inp[12]) ? node35355 : node35352;
																assign node35352 = (inp[4]) ? 4'b0100 : 4'b0000;
																assign node35355 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node35358 = (inp[15]) ? 4'b0110 : node35359;
															assign node35359 = (inp[4]) ? node35361 : 4'b0100;
																assign node35361 = (inp[12]) ? 4'b0000 : 4'b0100;
												assign node35365 = (inp[12]) ? node35385 : node35366;
													assign node35366 = (inp[15]) ? node35376 : node35367;
														assign node35367 = (inp[0]) ? node35373 : node35368;
															assign node35368 = (inp[9]) ? 4'b0010 : node35369;
																assign node35369 = (inp[4]) ? 4'b0010 : 4'b0110;
															assign node35373 = (inp[4]) ? 4'b0110 : 4'b0100;
														assign node35376 = (inp[0]) ? node35378 : 4'b0100;
															assign node35378 = (inp[4]) ? node35382 : node35379;
																assign node35379 = (inp[9]) ? 4'b0010 : 4'b0110;
																assign node35382 = (inp[9]) ? 4'b0100 : 4'b0010;
													assign node35385 = (inp[15]) ? node35397 : node35386;
														assign node35386 = (inp[0]) ? node35394 : node35387;
															assign node35387 = (inp[4]) ? node35391 : node35388;
																assign node35388 = (inp[9]) ? 4'b0100 : 4'b0010;
																assign node35391 = (inp[9]) ? 4'b0000 : 4'b0100;
															assign node35394 = (inp[4]) ? 4'b0010 : 4'b0000;
														assign node35397 = (inp[4]) ? node35405 : node35398;
															assign node35398 = (inp[9]) ? node35402 : node35399;
																assign node35399 = (inp[0]) ? 4'b0010 : 4'b0000;
																assign node35402 = (inp[0]) ? 4'b0100 : 4'b0110;
															assign node35405 = (inp[9]) ? 4'b0010 : 4'b0110;
											assign node35408 = (inp[0]) ? node35432 : node35409;
												assign node35409 = (inp[15]) ? node35419 : node35410;
													assign node35410 = (inp[5]) ? node35414 : node35411;
														assign node35411 = (inp[9]) ? 4'b0010 : 4'b0110;
														assign node35414 = (inp[9]) ? node35416 : 4'b0100;
															assign node35416 = (inp[4]) ? 4'b0000 : 4'b0100;
													assign node35419 = (inp[4]) ? node35427 : node35420;
														assign node35420 = (inp[12]) ? node35424 : node35421;
															assign node35421 = (inp[9]) ? 4'b0000 : 4'b0100;
															assign node35424 = (inp[5]) ? 4'b0010 : 4'b0110;
														assign node35427 = (inp[12]) ? node35429 : 4'b0110;
															assign node35429 = (inp[9]) ? 4'b0010 : 4'b0110;
												assign node35432 = (inp[15]) ? node35454 : node35433;
													assign node35433 = (inp[5]) ? node35441 : node35434;
														assign node35434 = (inp[4]) ? node35436 : 4'b0000;
															assign node35436 = (inp[9]) ? node35438 : 4'b0110;
																assign node35438 = (inp[12]) ? 4'b0010 : 4'b0110;
														assign node35441 = (inp[4]) ? node35447 : node35442;
															assign node35442 = (inp[9]) ? node35444 : 4'b0110;
																assign node35444 = (inp[12]) ? 4'b0110 : 4'b0010;
															assign node35447 = (inp[9]) ? node35451 : node35448;
																assign node35448 = (inp[12]) ? 4'b0110 : 4'b0010;
																assign node35451 = (inp[12]) ? 4'b0010 : 4'b0110;
													assign node35454 = (inp[5]) ? node35462 : node35455;
														assign node35455 = (inp[9]) ? 4'b0000 : node35456;
															assign node35456 = (inp[12]) ? 4'b0010 : node35457;
																assign node35457 = (inp[4]) ? 4'b0010 : 4'b0110;
														assign node35462 = (inp[12]) ? 4'b0000 : node35463;
															assign node35463 = (inp[9]) ? node35467 : node35464;
																assign node35464 = (inp[4]) ? 4'b0000 : 4'b0100;
																assign node35467 = (inp[4]) ? 4'b0100 : 4'b0000;
										assign node35471 = (inp[3]) ? node35563 : node35472;
											assign node35472 = (inp[5]) ? node35524 : node35473;
												assign node35473 = (inp[9]) ? node35501 : node35474;
													assign node35474 = (inp[12]) ? node35488 : node35475;
														assign node35475 = (inp[4]) ? node35481 : node35476;
															assign node35476 = (inp[0]) ? 4'b0110 : node35477;
																assign node35477 = (inp[15]) ? 4'b0100 : 4'b0110;
															assign node35481 = (inp[15]) ? node35485 : node35482;
																assign node35482 = (inp[0]) ? 4'b0000 : 4'b0010;
																assign node35485 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node35488 = (inp[4]) ? node35494 : node35489;
															assign node35489 = (inp[15]) ? node35491 : 4'b0000;
																assign node35491 = (inp[0]) ? 4'b0010 : 4'b0000;
															assign node35494 = (inp[0]) ? node35498 : node35495;
																assign node35495 = (inp[15]) ? 4'b0100 : 4'b0110;
																assign node35498 = (inp[15]) ? 4'b0110 : 4'b0100;
													assign node35501 = (inp[12]) ? node35511 : node35502;
														assign node35502 = (inp[4]) ? 4'b0100 : node35503;
															assign node35503 = (inp[0]) ? node35507 : node35504;
																assign node35504 = (inp[15]) ? 4'b0000 : 4'b0010;
																assign node35507 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node35511 = (inp[4]) ? node35517 : node35512;
															assign node35512 = (inp[15]) ? 4'b0110 : node35513;
																assign node35513 = (inp[0]) ? 4'b0100 : 4'b0110;
															assign node35517 = (inp[0]) ? node35521 : node35518;
																assign node35518 = (inp[15]) ? 4'b0000 : 4'b0010;
																assign node35521 = (inp[15]) ? 4'b0010 : 4'b0000;
												assign node35524 = (inp[15]) ? node35546 : node35525;
													assign node35525 = (inp[12]) ? node35539 : node35526;
														assign node35526 = (inp[0]) ? node35534 : node35527;
															assign node35527 = (inp[4]) ? node35531 : node35528;
																assign node35528 = (inp[9]) ? 4'b0010 : 4'b0110;
																assign node35531 = (inp[9]) ? 4'b0100 : 4'b0010;
															assign node35534 = (inp[9]) ? 4'b0110 : node35535;
																assign node35535 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node35539 = (inp[0]) ? node35541 : 4'b0100;
															assign node35541 = (inp[4]) ? node35543 : 4'b0000;
																assign node35543 = (inp[9]) ? 4'b0010 : 4'b0110;
													assign node35546 = (inp[12]) ? node35558 : node35547;
														assign node35547 = (inp[0]) ? node35551 : node35548;
															assign node35548 = (inp[4]) ? 4'b0110 : 4'b0100;
															assign node35551 = (inp[9]) ? node35555 : node35552;
																assign node35552 = (inp[4]) ? 4'b0010 : 4'b0110;
																assign node35555 = (inp[4]) ? 4'b0100 : 4'b0010;
														assign node35558 = (inp[4]) ? 4'b0010 : node35559;
															assign node35559 = (inp[9]) ? 4'b0100 : 4'b0010;
											assign node35563 = (inp[5]) ? node35607 : node35564;
												assign node35564 = (inp[4]) ? node35582 : node35565;
													assign node35565 = (inp[12]) ? node35573 : node35566;
														assign node35566 = (inp[9]) ? node35568 : 4'b0110;
															assign node35568 = (inp[0]) ? 4'b0000 : node35569;
																assign node35569 = (inp[15]) ? 4'b0000 : 4'b0010;
														assign node35573 = (inp[9]) ? 4'b0110 : node35574;
															assign node35574 = (inp[15]) ? node35578 : node35575;
																assign node35575 = (inp[0]) ? 4'b0000 : 4'b0010;
																assign node35578 = (inp[0]) ? 4'b0010 : 4'b0000;
													assign node35582 = (inp[9]) ? node35596 : node35583;
														assign node35583 = (inp[12]) ? node35589 : node35584;
															assign node35584 = (inp[15]) ? node35586 : 4'b0000;
																assign node35586 = (inp[0]) ? 4'b0010 : 4'b0000;
															assign node35589 = (inp[0]) ? node35593 : node35590;
																assign node35590 = (inp[15]) ? 4'b0110 : 4'b0100;
																assign node35593 = (inp[15]) ? 4'b0100 : 4'b0110;
														assign node35596 = (inp[12]) ? node35600 : node35597;
															assign node35597 = (inp[0]) ? 4'b0100 : 4'b0110;
															assign node35600 = (inp[15]) ? node35604 : node35601;
																assign node35601 = (inp[0]) ? 4'b0010 : 4'b0000;
																assign node35604 = (inp[0]) ? 4'b0000 : 4'b0010;
												assign node35607 = (inp[4]) ? node35621 : node35608;
													assign node35608 = (inp[9]) ? node35612 : node35609;
														assign node35609 = (inp[12]) ? 4'b0000 : 4'b0100;
														assign node35612 = (inp[12]) ? 4'b0100 : node35613;
															assign node35613 = (inp[15]) ? node35617 : node35614;
																assign node35614 = (inp[0]) ? 4'b0010 : 4'b0000;
																assign node35617 = (inp[0]) ? 4'b0000 : 4'b0010;
													assign node35621 = (inp[12]) ? node35633 : node35622;
														assign node35622 = (inp[9]) ? node35628 : node35623;
															assign node35623 = (inp[15]) ? 4'b0000 : node35624;
																assign node35624 = (inp[0]) ? 4'b0010 : 4'b0000;
															assign node35628 = (inp[15]) ? 4'b0100 : node35629;
																assign node35629 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node35633 = (inp[9]) ? node35637 : node35634;
															assign node35634 = (inp[15]) ? 4'b0110 : 4'b0100;
															assign node35637 = (inp[0]) ? node35641 : node35638;
																assign node35638 = (inp[15]) ? 4'b0010 : 4'b0000;
																assign node35641 = (inp[15]) ? 4'b0000 : 4'b0010;
					assign node35644 = (inp[13]) ? node37870 : node35645;
						assign node35645 = (inp[8]) ? node36801 : node35646;
							assign node35646 = (inp[7]) ? node36230 : node35647;
								assign node35647 = (inp[2]) ? node35937 : node35648;
									assign node35648 = (inp[14]) ? node35794 : node35649;
										assign node35649 = (inp[15]) ? node35717 : node35650;
											assign node35650 = (inp[9]) ? node35684 : node35651;
												assign node35651 = (inp[5]) ? node35663 : node35652;
													assign node35652 = (inp[0]) ? node35658 : node35653;
														assign node35653 = (inp[12]) ? node35655 : 4'b1011;
															assign node35655 = (inp[4]) ? 4'b1101 : 4'b1011;
														assign node35658 = (inp[3]) ? node35660 : 4'b1001;
															assign node35660 = (inp[4]) ? 4'b1001 : 4'b1101;
													assign node35663 = (inp[3]) ? node35677 : node35664;
														assign node35664 = (inp[0]) ? node35670 : node35665;
															assign node35665 = (inp[12]) ? 4'b1101 : node35666;
																assign node35666 = (inp[4]) ? 4'b1011 : 4'b1111;
															assign node35670 = (inp[4]) ? node35674 : node35671;
																assign node35671 = (inp[12]) ? 4'b1001 : 4'b1101;
																assign node35674 = (inp[12]) ? 4'b1111 : 4'b1001;
														assign node35677 = (inp[0]) ? node35679 : 4'b1001;
															assign node35679 = (inp[12]) ? 4'b1011 : node35680;
																assign node35680 = (inp[4]) ? 4'b1011 : 4'b1111;
												assign node35684 = (inp[0]) ? node35700 : node35685;
													assign node35685 = (inp[3]) ? node35693 : node35686;
														assign node35686 = (inp[12]) ? 4'b1011 : node35687;
															assign node35687 = (inp[4]) ? node35689 : 4'b1011;
																assign node35689 = (inp[5]) ? 4'b1101 : 4'b1111;
														assign node35693 = (inp[5]) ? node35695 : 4'b1101;
															assign node35695 = (inp[4]) ? node35697 : 4'b1001;
																assign node35697 = (inp[12]) ? 4'b1001 : 4'b1101;
													assign node35700 = (inp[3]) ? node35710 : node35701;
														assign node35701 = (inp[5]) ? node35703 : 4'b1001;
															assign node35703 = (inp[4]) ? node35707 : node35704;
																assign node35704 = (inp[12]) ? 4'b1111 : 4'b1001;
																assign node35707 = (inp[12]) ? 4'b1011 : 4'b1111;
														assign node35710 = (inp[4]) ? node35714 : node35711;
															assign node35711 = (inp[12]) ? 4'b1111 : 4'b1011;
															assign node35714 = (inp[12]) ? 4'b1011 : 4'b1111;
											assign node35717 = (inp[4]) ? node35763 : node35718;
												assign node35718 = (inp[0]) ? node35742 : node35719;
													assign node35719 = (inp[5]) ? node35731 : node35720;
														assign node35720 = (inp[3]) ? node35726 : node35721;
															assign node35721 = (inp[9]) ? 4'b1101 : node35722;
																assign node35722 = (inp[12]) ? 4'b1001 : 4'b1101;
															assign node35726 = (inp[12]) ? 4'b1001 : node35727;
																assign node35727 = (inp[9]) ? 4'b1001 : 4'b1101;
														assign node35731 = (inp[3]) ? node35739 : node35732;
															assign node35732 = (inp[9]) ? node35736 : node35733;
																assign node35733 = (inp[12]) ? 4'b1001 : 4'b1101;
																assign node35736 = (inp[12]) ? 4'b1111 : 4'b1001;
															assign node35739 = (inp[12]) ? 4'b1111 : 4'b1011;
													assign node35742 = (inp[5]) ? node35752 : node35743;
														assign node35743 = (inp[3]) ? node35749 : node35744;
															assign node35744 = (inp[9]) ? 4'b1111 : node35745;
																assign node35745 = (inp[12]) ? 4'b1011 : 4'b1111;
															assign node35749 = (inp[12]) ? 4'b1101 : 4'b1011;
														assign node35752 = (inp[3]) ? node35756 : node35753;
															assign node35753 = (inp[9]) ? 4'b1101 : 4'b1011;
															assign node35756 = (inp[12]) ? node35760 : node35757;
																assign node35757 = (inp[9]) ? 4'b1001 : 4'b1101;
																assign node35760 = (inp[9]) ? 4'b1101 : 4'b1001;
												assign node35763 = (inp[0]) ? node35779 : node35764;
													assign node35764 = (inp[5]) ? node35772 : node35765;
														assign node35765 = (inp[3]) ? 4'b1111 : node35766;
															assign node35766 = (inp[12]) ? node35768 : 4'b1001;
																assign node35768 = (inp[9]) ? 4'b1001 : 4'b1101;
														assign node35772 = (inp[12]) ? node35776 : node35773;
															assign node35773 = (inp[3]) ? 4'b1011 : 4'b1111;
															assign node35776 = (inp[9]) ? 4'b1011 : 4'b1111;
													assign node35779 = (inp[5]) ? node35787 : node35780;
														assign node35780 = (inp[9]) ? node35784 : node35781;
															assign node35781 = (inp[3]) ? 4'b1011 : 4'b1111;
															assign node35784 = (inp[12]) ? 4'b1001 : 4'b1101;
														assign node35787 = (inp[9]) ? node35791 : node35788;
															assign node35788 = (inp[12]) ? 4'b1101 : 4'b1001;
															assign node35791 = (inp[12]) ? 4'b1001 : 4'b1101;
										assign node35794 = (inp[5]) ? node35866 : node35795;
											assign node35795 = (inp[4]) ? node35829 : node35796;
												assign node35796 = (inp[15]) ? node35806 : node35797;
													assign node35797 = (inp[0]) ? node35801 : node35798;
														assign node35798 = (inp[9]) ? 4'b1010 : 4'b1110;
														assign node35801 = (inp[12]) ? 4'b1000 : node35802;
															assign node35802 = (inp[9]) ? 4'b1000 : 4'b1100;
													assign node35806 = (inp[0]) ? node35816 : node35807;
														assign node35807 = (inp[9]) ? node35811 : node35808;
															assign node35808 = (inp[12]) ? 4'b1000 : 4'b1100;
															assign node35811 = (inp[12]) ? node35813 : 4'b1000;
																assign node35813 = (inp[3]) ? 4'b1110 : 4'b1100;
														assign node35816 = (inp[3]) ? node35824 : node35817;
															assign node35817 = (inp[9]) ? node35821 : node35818;
																assign node35818 = (inp[12]) ? 4'b1010 : 4'b1110;
																assign node35821 = (inp[12]) ? 4'b1110 : 4'b1010;
															assign node35824 = (inp[9]) ? 4'b1010 : node35825;
																assign node35825 = (inp[12]) ? 4'b1010 : 4'b1110;
												assign node35829 = (inp[15]) ? node35843 : node35830;
													assign node35830 = (inp[0]) ? node35840 : node35831;
														assign node35831 = (inp[3]) ? 4'b1010 : node35832;
															assign node35832 = (inp[12]) ? node35836 : node35833;
																assign node35833 = (inp[9]) ? 4'b1110 : 4'b1010;
																assign node35836 = (inp[9]) ? 4'b1010 : 4'b1110;
														assign node35840 = (inp[3]) ? 4'b1110 : 4'b1100;
													assign node35843 = (inp[0]) ? node35857 : node35844;
														assign node35844 = (inp[3]) ? node35850 : node35845;
															assign node35845 = (inp[9]) ? node35847 : 4'b1100;
																assign node35847 = (inp[12]) ? 4'b1000 : 4'b1100;
															assign node35850 = (inp[9]) ? node35854 : node35851;
																assign node35851 = (inp[12]) ? 4'b1110 : 4'b1000;
																assign node35854 = (inp[12]) ? 4'b1010 : 4'b1110;
														assign node35857 = (inp[3]) ? node35863 : node35858;
															assign node35858 = (inp[9]) ? 4'b1010 : node35859;
																assign node35859 = (inp[12]) ? 4'b1110 : 4'b1010;
															assign node35863 = (inp[9]) ? 4'b1100 : 4'b1010;
											assign node35866 = (inp[0]) ? node35904 : node35867;
												assign node35867 = (inp[15]) ? node35885 : node35868;
													assign node35868 = (inp[12]) ? node35880 : node35869;
														assign node35869 = (inp[3]) ? node35873 : node35870;
															assign node35870 = (inp[9]) ? 4'b1010 : 4'b1110;
															assign node35873 = (inp[4]) ? node35877 : node35874;
																assign node35874 = (inp[9]) ? 4'b1000 : 4'b1100;
																assign node35877 = (inp[9]) ? 4'b1100 : 4'b1000;
														assign node35880 = (inp[4]) ? node35882 : 4'b1100;
															assign node35882 = (inp[9]) ? 4'b1000 : 4'b1100;
													assign node35885 = (inp[3]) ? node35895 : node35886;
														assign node35886 = (inp[9]) ? node35892 : node35887;
															assign node35887 = (inp[4]) ? 4'b1000 : node35888;
																assign node35888 = (inp[12]) ? 4'b1000 : 4'b1100;
															assign node35892 = (inp[12]) ? 4'b1010 : 4'b1110;
														assign node35895 = (inp[9]) ? 4'b1110 : node35896;
															assign node35896 = (inp[12]) ? node35900 : node35897;
																assign node35897 = (inp[4]) ? 4'b1010 : 4'b1110;
																assign node35900 = (inp[4]) ? 4'b1110 : 4'b1010;
												assign node35904 = (inp[15]) ? node35922 : node35905;
													assign node35905 = (inp[12]) ? node35917 : node35906;
														assign node35906 = (inp[3]) ? node35912 : node35907;
															assign node35907 = (inp[9]) ? node35909 : 4'b1000;
																assign node35909 = (inp[4]) ? 4'b1110 : 4'b1000;
															assign node35912 = (inp[9]) ? node35914 : 4'b1010;
																assign node35914 = (inp[4]) ? 4'b1110 : 4'b1010;
														assign node35917 = (inp[9]) ? node35919 : 4'b1110;
															assign node35919 = (inp[4]) ? 4'b1010 : 4'b1110;
													assign node35922 = (inp[4]) ? 4'b1100 : node35923;
														assign node35923 = (inp[3]) ? node35931 : node35924;
															assign node35924 = (inp[12]) ? node35928 : node35925;
																assign node35925 = (inp[9]) ? 4'b1010 : 4'b1110;
																assign node35928 = (inp[9]) ? 4'b1100 : 4'b1010;
															assign node35931 = (inp[12]) ? node35933 : 4'b1100;
																assign node35933 = (inp[9]) ? 4'b1100 : 4'b1000;
									assign node35937 = (inp[14]) ? node36095 : node35938;
										assign node35938 = (inp[9]) ? node36024 : node35939;
											assign node35939 = (inp[5]) ? node35987 : node35940;
												assign node35940 = (inp[4]) ? node35966 : node35941;
													assign node35941 = (inp[12]) ? node35951 : node35942;
														assign node35942 = (inp[3]) ? node35944 : 4'b1100;
															assign node35944 = (inp[0]) ? node35948 : node35945;
																assign node35945 = (inp[15]) ? 4'b1100 : 4'b1110;
																assign node35948 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node35951 = (inp[3]) ? node35959 : node35952;
															assign node35952 = (inp[15]) ? node35956 : node35953;
																assign node35953 = (inp[0]) ? 4'b1000 : 4'b1010;
																assign node35956 = (inp[0]) ? 4'b1010 : 4'b1000;
															assign node35959 = (inp[0]) ? node35963 : node35960;
																assign node35960 = (inp[15]) ? 4'b1000 : 4'b1010;
																assign node35963 = (inp[15]) ? 4'b1010 : 4'b1000;
													assign node35966 = (inp[12]) ? node35974 : node35967;
														assign node35967 = (inp[0]) ? node35971 : node35968;
															assign node35968 = (inp[15]) ? 4'b1000 : 4'b1010;
															assign node35971 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node35974 = (inp[3]) ? node35982 : node35975;
															assign node35975 = (inp[0]) ? node35979 : node35976;
																assign node35976 = (inp[15]) ? 4'b1100 : 4'b1110;
																assign node35979 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node35982 = (inp[15]) ? node35984 : 4'b1110;
																assign node35984 = (inp[0]) ? 4'b1100 : 4'b1110;
												assign node35987 = (inp[4]) ? node36009 : node35988;
													assign node35988 = (inp[12]) ? node36002 : node35989;
														assign node35989 = (inp[15]) ? node35997 : node35990;
															assign node35990 = (inp[0]) ? node35994 : node35991;
																assign node35991 = (inp[3]) ? 4'b1100 : 4'b1110;
																assign node35994 = (inp[3]) ? 4'b1110 : 4'b1100;
															assign node35997 = (inp[3]) ? node35999 : 4'b1100;
																assign node35999 = (inp[0]) ? 4'b1100 : 4'b1110;
														assign node36002 = (inp[15]) ? node36004 : 4'b1000;
															assign node36004 = (inp[3]) ? 4'b1010 : node36005;
																assign node36005 = (inp[0]) ? 4'b1010 : 4'b1000;
													assign node36009 = (inp[12]) ? node36017 : node36010;
														assign node36010 = (inp[15]) ? 4'b1000 : node36011;
															assign node36011 = (inp[3]) ? node36013 : 4'b1010;
																assign node36013 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node36017 = (inp[15]) ? node36021 : node36018;
															assign node36018 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node36021 = (inp[0]) ? 4'b1100 : 4'b1110;
											assign node36024 = (inp[0]) ? node36058 : node36025;
												assign node36025 = (inp[15]) ? node36045 : node36026;
													assign node36026 = (inp[5]) ? node36040 : node36027;
														assign node36027 = (inp[3]) ? node36035 : node36028;
															assign node36028 = (inp[4]) ? node36032 : node36029;
																assign node36029 = (inp[12]) ? 4'b1110 : 4'b1010;
																assign node36032 = (inp[12]) ? 4'b1010 : 4'b1110;
															assign node36035 = (inp[12]) ? node36037 : 4'b1010;
																assign node36037 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node36040 = (inp[12]) ? node36042 : 4'b1100;
															assign node36042 = (inp[4]) ? 4'b1000 : 4'b1100;
													assign node36045 = (inp[5]) ? node36053 : node36046;
														assign node36046 = (inp[3]) ? node36048 : 4'b1000;
															assign node36048 = (inp[4]) ? node36050 : 4'b1110;
																assign node36050 = (inp[12]) ? 4'b1010 : 4'b1110;
														assign node36053 = (inp[4]) ? node36055 : 4'b1110;
															assign node36055 = (inp[12]) ? 4'b1010 : 4'b1110;
												assign node36058 = (inp[15]) ? node36080 : node36059;
													assign node36059 = (inp[3]) ? node36069 : node36060;
														assign node36060 = (inp[4]) ? node36064 : node36061;
															assign node36061 = (inp[12]) ? 4'b1100 : 4'b1000;
															assign node36064 = (inp[5]) ? node36066 : 4'b1100;
																assign node36066 = (inp[12]) ? 4'b1010 : 4'b1110;
														assign node36069 = (inp[5]) ? node36075 : node36070;
															assign node36070 = (inp[4]) ? node36072 : 4'b1110;
																assign node36072 = (inp[12]) ? 4'b1010 : 4'b1110;
															assign node36075 = (inp[12]) ? 4'b1110 : node36076;
																assign node36076 = (inp[4]) ? 4'b1110 : 4'b1010;
													assign node36080 = (inp[3]) ? node36090 : node36081;
														assign node36081 = (inp[5]) ? node36085 : node36082;
															assign node36082 = (inp[12]) ? 4'b1010 : 4'b1110;
															assign node36085 = (inp[4]) ? node36087 : 4'b1010;
																assign node36087 = (inp[12]) ? 4'b1000 : 4'b1100;
														assign node36090 = (inp[12]) ? node36092 : 4'b1100;
															assign node36092 = (inp[4]) ? 4'b1000 : 4'b1100;
										assign node36095 = (inp[12]) ? node36159 : node36096;
											assign node36096 = (inp[9]) ? node36136 : node36097;
												assign node36097 = (inp[4]) ? node36117 : node36098;
													assign node36098 = (inp[3]) ? node36112 : node36099;
														assign node36099 = (inp[5]) ? node36105 : node36100;
															assign node36100 = (inp[15]) ? 4'b1110 : node36101;
																assign node36101 = (inp[0]) ? 4'b1100 : 4'b1110;
															assign node36105 = (inp[15]) ? node36109 : node36106;
																assign node36106 = (inp[0]) ? 4'b1100 : 4'b1110;
																assign node36109 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node36112 = (inp[5]) ? 4'b1110 : node36113;
															assign node36113 = (inp[15]) ? 4'b1100 : 4'b1110;
													assign node36117 = (inp[0]) ? node36127 : node36118;
														assign node36118 = (inp[15]) ? node36122 : node36119;
															assign node36119 = (inp[3]) ? 4'b1000 : 4'b1010;
															assign node36122 = (inp[5]) ? node36124 : 4'b1000;
																assign node36124 = (inp[3]) ? 4'b1010 : 4'b1000;
														assign node36127 = (inp[15]) ? node36131 : node36128;
															assign node36128 = (inp[3]) ? 4'b1010 : 4'b1000;
															assign node36131 = (inp[3]) ? node36133 : 4'b1010;
																assign node36133 = (inp[5]) ? 4'b1000 : 4'b1010;
												assign node36136 = (inp[4]) ? node36144 : node36137;
													assign node36137 = (inp[15]) ? 4'b1000 : node36138;
														assign node36138 = (inp[0]) ? node36140 : 4'b1010;
															assign node36140 = (inp[5]) ? 4'b1010 : 4'b1000;
													assign node36144 = (inp[15]) ? node36148 : node36145;
														assign node36145 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node36148 = (inp[0]) ? node36154 : node36149;
															assign node36149 = (inp[3]) ? 4'b1110 : node36150;
																assign node36150 = (inp[5]) ? 4'b1110 : 4'b1100;
															assign node36154 = (inp[5]) ? 4'b1100 : node36155;
																assign node36155 = (inp[3]) ? 4'b1100 : 4'b1110;
											assign node36159 = (inp[5]) ? node36197 : node36160;
												assign node36160 = (inp[0]) ? node36174 : node36161;
													assign node36161 = (inp[9]) ? node36171 : node36162;
														assign node36162 = (inp[4]) ? node36164 : 4'b1010;
															assign node36164 = (inp[15]) ? node36168 : node36165;
																assign node36165 = (inp[3]) ? 4'b1100 : 4'b1110;
																assign node36168 = (inp[3]) ? 4'b1110 : 4'b1100;
														assign node36171 = (inp[4]) ? 4'b1010 : 4'b1110;
													assign node36174 = (inp[15]) ? node36188 : node36175;
														assign node36175 = (inp[3]) ? node36181 : node36176;
															assign node36176 = (inp[9]) ? node36178 : 4'b1000;
																assign node36178 = (inp[4]) ? 4'b1000 : 4'b1100;
															assign node36181 = (inp[4]) ? node36185 : node36182;
																assign node36182 = (inp[9]) ? 4'b1110 : 4'b1000;
																assign node36185 = (inp[9]) ? 4'b1010 : 4'b1110;
														assign node36188 = (inp[3]) ? node36194 : node36189;
															assign node36189 = (inp[4]) ? 4'b1110 : node36190;
																assign node36190 = (inp[9]) ? 4'b1110 : 4'b1010;
															assign node36194 = (inp[9]) ? 4'b1000 : 4'b1100;
												assign node36197 = (inp[15]) ? node36213 : node36198;
													assign node36198 = (inp[0]) ? node36204 : node36199;
														assign node36199 = (inp[4]) ? node36201 : 4'b1010;
															assign node36201 = (inp[9]) ? 4'b1000 : 4'b1100;
														assign node36204 = (inp[3]) ? node36206 : 4'b1110;
															assign node36206 = (inp[9]) ? node36210 : node36207;
																assign node36207 = (inp[4]) ? 4'b1110 : 4'b1010;
																assign node36210 = (inp[4]) ? 4'b1010 : 4'b1110;
													assign node36213 = (inp[0]) ? node36223 : node36214;
														assign node36214 = (inp[9]) ? node36220 : node36215;
															assign node36215 = (inp[3]) ? node36217 : 4'b1000;
																assign node36217 = (inp[4]) ? 4'b1110 : 4'b1010;
															assign node36220 = (inp[4]) ? 4'b1010 : 4'b1110;
														assign node36223 = (inp[9]) ? node36227 : node36224;
															assign node36224 = (inp[3]) ? 4'b1000 : 4'b1010;
															assign node36227 = (inp[4]) ? 4'b1000 : 4'b1100;
								assign node36230 = (inp[2]) ? node36532 : node36231;
									assign node36231 = (inp[14]) ? node36383 : node36232;
										assign node36232 = (inp[15]) ? node36306 : node36233;
											assign node36233 = (inp[12]) ? node36271 : node36234;
												assign node36234 = (inp[3]) ? node36250 : node36235;
													assign node36235 = (inp[0]) ? node36245 : node36236;
														assign node36236 = (inp[5]) ? node36238 : 4'b1010;
															assign node36238 = (inp[9]) ? node36242 : node36239;
																assign node36239 = (inp[4]) ? 4'b1010 : 4'b1110;
																assign node36242 = (inp[4]) ? 4'b1100 : 4'b1010;
														assign node36245 = (inp[4]) ? node36247 : 4'b1000;
															assign node36247 = (inp[9]) ? 4'b1110 : 4'b1000;
													assign node36250 = (inp[9]) ? node36262 : node36251;
														assign node36251 = (inp[4]) ? node36257 : node36252;
															assign node36252 = (inp[5]) ? 4'b1100 : node36253;
																assign node36253 = (inp[0]) ? 4'b1100 : 4'b1110;
															assign node36257 = (inp[0]) ? node36259 : 4'b1000;
																assign node36259 = (inp[5]) ? 4'b1010 : 4'b1000;
														assign node36262 = (inp[4]) ? node36268 : node36263;
															assign node36263 = (inp[0]) ? 4'b1010 : node36264;
																assign node36264 = (inp[5]) ? 4'b1000 : 4'b1010;
															assign node36268 = (inp[0]) ? 4'b1110 : 4'b1100;
												assign node36271 = (inp[0]) ? node36287 : node36272;
													assign node36272 = (inp[5]) ? node36282 : node36273;
														assign node36273 = (inp[3]) ? 4'b1100 : node36274;
															assign node36274 = (inp[9]) ? node36278 : node36275;
																assign node36275 = (inp[4]) ? 4'b1110 : 4'b1010;
																assign node36278 = (inp[4]) ? 4'b1010 : 4'b1110;
														assign node36282 = (inp[3]) ? node36284 : 4'b1100;
															assign node36284 = (inp[4]) ? 4'b1100 : 4'b1000;
													assign node36287 = (inp[5]) ? node36301 : node36288;
														assign node36288 = (inp[3]) ? node36294 : node36289;
															assign node36289 = (inp[9]) ? node36291 : 4'b1100;
																assign node36291 = (inp[4]) ? 4'b1000 : 4'b1100;
															assign node36294 = (inp[9]) ? node36298 : node36295;
																assign node36295 = (inp[4]) ? 4'b1110 : 4'b1000;
																assign node36298 = (inp[4]) ? 4'b1010 : 4'b1110;
														assign node36301 = (inp[3]) ? 4'b1010 : node36302;
															assign node36302 = (inp[9]) ? 4'b1010 : 4'b1110;
											assign node36306 = (inp[5]) ? node36340 : node36307;
												assign node36307 = (inp[0]) ? node36325 : node36308;
													assign node36308 = (inp[3]) ? node36318 : node36309;
														assign node36309 = (inp[4]) ? 4'b1100 : node36310;
															assign node36310 = (inp[12]) ? node36314 : node36311;
																assign node36311 = (inp[9]) ? 4'b1000 : 4'b1100;
																assign node36314 = (inp[9]) ? 4'b1100 : 4'b1000;
														assign node36318 = (inp[4]) ? 4'b1110 : node36319;
															assign node36319 = (inp[9]) ? 4'b1110 : node36320;
																assign node36320 = (inp[12]) ? 4'b1000 : 4'b1100;
													assign node36325 = (inp[3]) ? node36333 : node36326;
														assign node36326 = (inp[12]) ? 4'b1110 : node36327;
															assign node36327 = (inp[9]) ? 4'b1010 : node36328;
																assign node36328 = (inp[4]) ? 4'b1010 : 4'b1110;
														assign node36333 = (inp[4]) ? 4'b1100 : node36334;
															assign node36334 = (inp[9]) ? 4'b1100 : node36335;
																assign node36335 = (inp[12]) ? 4'b1010 : 4'b1110;
												assign node36340 = (inp[0]) ? node36354 : node36341;
													assign node36341 = (inp[3]) ? node36345 : node36342;
														assign node36342 = (inp[9]) ? 4'b1110 : 4'b1000;
														assign node36345 = (inp[12]) ? 4'b1010 : node36346;
															assign node36346 = (inp[9]) ? node36350 : node36347;
																assign node36347 = (inp[4]) ? 4'b1010 : 4'b1110;
																assign node36350 = (inp[4]) ? 4'b1110 : 4'b1010;
													assign node36354 = (inp[3]) ? node36368 : node36355;
														assign node36355 = (inp[9]) ? node36363 : node36356;
															assign node36356 = (inp[12]) ? node36360 : node36357;
																assign node36357 = (inp[4]) ? 4'b1010 : 4'b1110;
																assign node36360 = (inp[4]) ? 4'b1100 : 4'b1010;
															assign node36363 = (inp[4]) ? node36365 : 4'b1100;
																assign node36365 = (inp[12]) ? 4'b1000 : 4'b1100;
														assign node36368 = (inp[12]) ? node36376 : node36369;
															assign node36369 = (inp[4]) ? node36373 : node36370;
																assign node36370 = (inp[9]) ? 4'b1000 : 4'b1100;
																assign node36373 = (inp[9]) ? 4'b1100 : 4'b1000;
															assign node36376 = (inp[4]) ? node36380 : node36377;
																assign node36377 = (inp[9]) ? 4'b1100 : 4'b1000;
																assign node36380 = (inp[9]) ? 4'b1000 : 4'b1100;
										assign node36383 = (inp[5]) ? node36451 : node36384;
											assign node36384 = (inp[4]) ? node36418 : node36385;
												assign node36385 = (inp[0]) ? node36403 : node36386;
													assign node36386 = (inp[15]) ? node36396 : node36387;
														assign node36387 = (inp[9]) ? node36391 : node36388;
															assign node36388 = (inp[12]) ? 4'b0011 : 4'b0111;
															assign node36391 = (inp[3]) ? 4'b0101 : node36392;
																assign node36392 = (inp[12]) ? 4'b0111 : 4'b0011;
														assign node36396 = (inp[12]) ? node36400 : node36397;
															assign node36397 = (inp[9]) ? 4'b0001 : 4'b0101;
															assign node36400 = (inp[3]) ? 4'b0111 : 4'b0101;
													assign node36403 = (inp[15]) ? node36411 : node36404;
														assign node36404 = (inp[12]) ? node36408 : node36405;
															assign node36405 = (inp[9]) ? 4'b0001 : 4'b0101;
															assign node36408 = (inp[9]) ? 4'b0111 : 4'b0001;
														assign node36411 = (inp[9]) ? node36415 : node36412;
															assign node36412 = (inp[12]) ? 4'b0011 : 4'b0111;
															assign node36415 = (inp[12]) ? 4'b0111 : 4'b0011;
												assign node36418 = (inp[15]) ? node36430 : node36419;
													assign node36419 = (inp[12]) ? node36421 : 4'b0011;
														assign node36421 = (inp[9]) ? node36423 : 4'b0101;
															assign node36423 = (inp[3]) ? node36427 : node36424;
																assign node36424 = (inp[0]) ? 4'b0001 : 4'b0011;
																assign node36427 = (inp[0]) ? 4'b0011 : 4'b0001;
													assign node36430 = (inp[0]) ? node36444 : node36431;
														assign node36431 = (inp[3]) ? node36437 : node36432;
															assign node36432 = (inp[12]) ? 4'b0101 : node36433;
																assign node36433 = (inp[9]) ? 4'b0101 : 4'b0001;
															assign node36437 = (inp[12]) ? node36441 : node36438;
																assign node36438 = (inp[9]) ? 4'b0111 : 4'b0001;
																assign node36441 = (inp[9]) ? 4'b0011 : 4'b0111;
														assign node36444 = (inp[3]) ? 4'b0001 : node36445;
															assign node36445 = (inp[9]) ? node36447 : 4'b0011;
																assign node36447 = (inp[12]) ? 4'b0011 : 4'b0111;
											assign node36451 = (inp[3]) ? node36493 : node36452;
												assign node36452 = (inp[15]) ? node36474 : node36453;
													assign node36453 = (inp[0]) ? node36465 : node36454;
														assign node36454 = (inp[12]) ? node36458 : node36455;
															assign node36455 = (inp[9]) ? 4'b0011 : 4'b0111;
															assign node36458 = (inp[4]) ? node36462 : node36459;
																assign node36459 = (inp[9]) ? 4'b0101 : 4'b0011;
																assign node36462 = (inp[9]) ? 4'b0001 : 4'b0101;
														assign node36465 = (inp[4]) ? node36471 : node36466;
															assign node36466 = (inp[9]) ? 4'b0001 : node36467;
																assign node36467 = (inp[12]) ? 4'b0001 : 4'b0101;
															assign node36471 = (inp[9]) ? 4'b0111 : 4'b0001;
													assign node36474 = (inp[12]) ? node36484 : node36475;
														assign node36475 = (inp[0]) ? node36479 : node36476;
															assign node36476 = (inp[4]) ? 4'b0001 : 4'b0101;
															assign node36479 = (inp[9]) ? node36481 : 4'b0011;
																assign node36481 = (inp[4]) ? 4'b0101 : 4'b0011;
														assign node36484 = (inp[0]) ? 4'b0011 : node36485;
															assign node36485 = (inp[4]) ? node36489 : node36486;
																assign node36486 = (inp[9]) ? 4'b0111 : 4'b0001;
																assign node36489 = (inp[9]) ? 4'b0011 : 4'b0111;
												assign node36493 = (inp[0]) ? node36515 : node36494;
													assign node36494 = (inp[15]) ? node36508 : node36495;
														assign node36495 = (inp[12]) ? node36503 : node36496;
															assign node36496 = (inp[4]) ? node36500 : node36497;
																assign node36497 = (inp[9]) ? 4'b0001 : 4'b0101;
																assign node36500 = (inp[9]) ? 4'b0101 : 4'b0001;
															assign node36503 = (inp[9]) ? node36505 : 4'b0001;
																assign node36505 = (inp[4]) ? 4'b0001 : 4'b0101;
														assign node36508 = (inp[12]) ? node36512 : node36509;
															assign node36509 = (inp[4]) ? 4'b0111 : 4'b0011;
															assign node36512 = (inp[4]) ? 4'b0011 : 4'b0111;
													assign node36515 = (inp[15]) ? node36525 : node36516;
														assign node36516 = (inp[9]) ? 4'b0111 : node36517;
															assign node36517 = (inp[12]) ? node36521 : node36518;
																assign node36518 = (inp[4]) ? 4'b0011 : 4'b0111;
																assign node36521 = (inp[4]) ? 4'b0111 : 4'b0011;
														assign node36525 = (inp[12]) ? node36527 : 4'b0101;
															assign node36527 = (inp[9]) ? 4'b0101 : node36528;
																assign node36528 = (inp[4]) ? 4'b0101 : 4'b0001;
									assign node36532 = (inp[5]) ? node36680 : node36533;
										assign node36533 = (inp[4]) ? node36585 : node36534;
											assign node36534 = (inp[12]) ? node36556 : node36535;
												assign node36535 = (inp[9]) ? node36549 : node36536;
													assign node36536 = (inp[3]) ? node36542 : node36537;
														assign node36537 = (inp[15]) ? 4'b0111 : node36538;
															assign node36538 = (inp[0]) ? 4'b0101 : 4'b0111;
														assign node36542 = (inp[15]) ? node36546 : node36543;
															assign node36543 = (inp[0]) ? 4'b0101 : 4'b0111;
															assign node36546 = (inp[0]) ? 4'b0111 : 4'b0101;
													assign node36549 = (inp[0]) ? node36553 : node36550;
														assign node36550 = (inp[15]) ? 4'b0001 : 4'b0011;
														assign node36553 = (inp[15]) ? 4'b0011 : 4'b0001;
												assign node36556 = (inp[9]) ? node36562 : node36557;
													assign node36557 = (inp[3]) ? node36559 : 4'b0001;
														assign node36559 = (inp[0]) ? 4'b0001 : 4'b0011;
													assign node36562 = (inp[0]) ? node36576 : node36563;
														assign node36563 = (inp[14]) ? node36569 : node36564;
															assign node36564 = (inp[3]) ? node36566 : 4'b0111;
																assign node36566 = (inp[15]) ? 4'b0111 : 4'b0101;
															assign node36569 = (inp[3]) ? node36573 : node36570;
																assign node36570 = (inp[15]) ? 4'b0101 : 4'b0111;
																assign node36573 = (inp[15]) ? 4'b0111 : 4'b0101;
														assign node36576 = (inp[14]) ? node36582 : node36577;
															assign node36577 = (inp[15]) ? 4'b0101 : node36578;
																assign node36578 = (inp[3]) ? 4'b0111 : 4'b0101;
															assign node36582 = (inp[15]) ? 4'b0111 : 4'b0101;
											assign node36585 = (inp[3]) ? node36643 : node36586;
												assign node36586 = (inp[14]) ? node36618 : node36587;
													assign node36587 = (inp[15]) ? node36603 : node36588;
														assign node36588 = (inp[0]) ? node36596 : node36589;
															assign node36589 = (inp[9]) ? node36593 : node36590;
																assign node36590 = (inp[12]) ? 4'b0111 : 4'b0011;
																assign node36593 = (inp[12]) ? 4'b0011 : 4'b0111;
															assign node36596 = (inp[12]) ? node36600 : node36597;
																assign node36597 = (inp[9]) ? 4'b0101 : 4'b0001;
																assign node36600 = (inp[9]) ? 4'b0001 : 4'b0101;
														assign node36603 = (inp[0]) ? node36611 : node36604;
															assign node36604 = (inp[9]) ? node36608 : node36605;
																assign node36605 = (inp[12]) ? 4'b0101 : 4'b0001;
																assign node36608 = (inp[12]) ? 4'b0001 : 4'b0101;
															assign node36611 = (inp[12]) ? node36615 : node36612;
																assign node36612 = (inp[9]) ? 4'b0111 : 4'b0011;
																assign node36615 = (inp[9]) ? 4'b0011 : 4'b0111;
													assign node36618 = (inp[12]) ? node36632 : node36619;
														assign node36619 = (inp[9]) ? node36625 : node36620;
															assign node36620 = (inp[15]) ? 4'b0001 : node36621;
																assign node36621 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node36625 = (inp[0]) ? node36629 : node36626;
																assign node36626 = (inp[15]) ? 4'b0101 : 4'b0111;
																assign node36629 = (inp[15]) ? 4'b0111 : 4'b0101;
														assign node36632 = (inp[9]) ? node36638 : node36633;
															assign node36633 = (inp[0]) ? 4'b0101 : node36634;
																assign node36634 = (inp[15]) ? 4'b0101 : 4'b0111;
															assign node36638 = (inp[0]) ? node36640 : 4'b0001;
																assign node36640 = (inp[15]) ? 4'b0011 : 4'b0001;
												assign node36643 = (inp[14]) ? node36659 : node36644;
													assign node36644 = (inp[9]) ? node36652 : node36645;
														assign node36645 = (inp[12]) ? node36649 : node36646;
															assign node36646 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node36649 = (inp[15]) ? 4'b0101 : 4'b0111;
														assign node36652 = (inp[12]) ? node36654 : 4'b0101;
															assign node36654 = (inp[0]) ? 4'b0001 : node36655;
																assign node36655 = (inp[15]) ? 4'b0011 : 4'b0001;
													assign node36659 = (inp[9]) ? node36667 : node36660;
														assign node36660 = (inp[12]) ? 4'b0111 : node36661;
															assign node36661 = (inp[15]) ? 4'b0011 : node36662;
																assign node36662 = (inp[0]) ? 4'b0001 : 4'b0011;
														assign node36667 = (inp[12]) ? node36675 : node36668;
															assign node36668 = (inp[0]) ? node36672 : node36669;
																assign node36669 = (inp[15]) ? 4'b0111 : 4'b0101;
																assign node36672 = (inp[15]) ? 4'b0101 : 4'b0111;
															assign node36675 = (inp[15]) ? 4'b0011 : node36676;
																assign node36676 = (inp[0]) ? 4'b0011 : 4'b0001;
										assign node36680 = (inp[12]) ? node36748 : node36681;
											assign node36681 = (inp[0]) ? node36717 : node36682;
												assign node36682 = (inp[15]) ? node36700 : node36683;
													assign node36683 = (inp[3]) ? node36693 : node36684;
														assign node36684 = (inp[14]) ? node36686 : 4'b0101;
															assign node36686 = (inp[9]) ? node36690 : node36687;
																assign node36687 = (inp[4]) ? 4'b0011 : 4'b0111;
																assign node36690 = (inp[4]) ? 4'b0101 : 4'b0011;
														assign node36693 = (inp[4]) ? node36697 : node36694;
															assign node36694 = (inp[9]) ? 4'b0001 : 4'b0101;
															assign node36697 = (inp[9]) ? 4'b0101 : 4'b0001;
													assign node36700 = (inp[3]) ? node36708 : node36701;
														assign node36701 = (inp[4]) ? node36705 : node36702;
															assign node36702 = (inp[9]) ? 4'b0001 : 4'b0101;
															assign node36705 = (inp[9]) ? 4'b0111 : 4'b0001;
														assign node36708 = (inp[14]) ? 4'b0111 : node36709;
															assign node36709 = (inp[9]) ? node36713 : node36710;
																assign node36710 = (inp[4]) ? 4'b0011 : 4'b0111;
																assign node36713 = (inp[4]) ? 4'b0111 : 4'b0011;
												assign node36717 = (inp[15]) ? node36731 : node36718;
													assign node36718 = (inp[3]) ? node36724 : node36719;
														assign node36719 = (inp[9]) ? node36721 : 4'b0001;
															assign node36721 = (inp[4]) ? 4'b0111 : 4'b0001;
														assign node36724 = (inp[4]) ? node36728 : node36725;
															assign node36725 = (inp[9]) ? 4'b0011 : 4'b0111;
															assign node36728 = (inp[9]) ? 4'b0111 : 4'b0011;
													assign node36731 = (inp[3]) ? node36739 : node36732;
														assign node36732 = (inp[9]) ? node36736 : node36733;
															assign node36733 = (inp[4]) ? 4'b0011 : 4'b0111;
															assign node36736 = (inp[4]) ? 4'b0101 : 4'b0011;
														assign node36739 = (inp[14]) ? 4'b0001 : node36740;
															assign node36740 = (inp[4]) ? node36744 : node36741;
																assign node36741 = (inp[9]) ? 4'b0001 : 4'b0101;
																assign node36744 = (inp[9]) ? 4'b0101 : 4'b0001;
											assign node36748 = (inp[14]) ? node36774 : node36749;
												assign node36749 = (inp[4]) ? node36763 : node36750;
													assign node36750 = (inp[9]) ? node36760 : node36751;
														assign node36751 = (inp[0]) ? node36753 : 4'b0011;
															assign node36753 = (inp[15]) ? node36757 : node36754;
																assign node36754 = (inp[3]) ? 4'b0011 : 4'b0001;
																assign node36757 = (inp[3]) ? 4'b0001 : 4'b0011;
														assign node36760 = (inp[3]) ? 4'b0111 : 4'b0101;
													assign node36763 = (inp[9]) ? node36771 : node36764;
														assign node36764 = (inp[0]) ? node36768 : node36765;
															assign node36765 = (inp[15]) ? 4'b0111 : 4'b0101;
															assign node36768 = (inp[15]) ? 4'b0101 : 4'b0111;
														assign node36771 = (inp[3]) ? 4'b0001 : 4'b0011;
												assign node36774 = (inp[0]) ? node36792 : node36775;
													assign node36775 = (inp[15]) ? node36785 : node36776;
														assign node36776 = (inp[3]) ? 4'b0101 : node36777;
															assign node36777 = (inp[4]) ? node36781 : node36778;
																assign node36778 = (inp[9]) ? 4'b0101 : 4'b0011;
																assign node36781 = (inp[9]) ? 4'b0001 : 4'b0101;
														assign node36785 = (inp[9]) ? node36789 : node36786;
															assign node36786 = (inp[4]) ? 4'b0111 : 4'b0001;
															assign node36789 = (inp[4]) ? 4'b0011 : 4'b0111;
													assign node36792 = (inp[15]) ? 4'b0101 : node36793;
														assign node36793 = (inp[9]) ? node36797 : node36794;
															assign node36794 = (inp[4]) ? 4'b0111 : 4'b0011;
															assign node36797 = (inp[4]) ? 4'b0011 : 4'b0111;
							assign node36801 = (inp[7]) ? node37345 : node36802;
								assign node36802 = (inp[2]) ? node37092 : node36803;
									assign node36803 = (inp[14]) ? node36951 : node36804;
										assign node36804 = (inp[0]) ? node36886 : node36805;
											assign node36805 = (inp[4]) ? node36845 : node36806;
												assign node36806 = (inp[15]) ? node36822 : node36807;
													assign node36807 = (inp[3]) ? node36817 : node36808;
														assign node36808 = (inp[9]) ? node36812 : node36809;
															assign node36809 = (inp[12]) ? 4'b1010 : 4'b1110;
															assign node36812 = (inp[12]) ? node36814 : 4'b1010;
																assign node36814 = (inp[5]) ? 4'b1100 : 4'b1110;
														assign node36817 = (inp[12]) ? 4'b1100 : node36818;
															assign node36818 = (inp[9]) ? 4'b1000 : 4'b1100;
													assign node36822 = (inp[5]) ? node36832 : node36823;
														assign node36823 = (inp[12]) ? node36827 : node36824;
															assign node36824 = (inp[9]) ? 4'b1000 : 4'b1100;
															assign node36827 = (inp[9]) ? node36829 : 4'b1000;
																assign node36829 = (inp[3]) ? 4'b1110 : 4'b1100;
														assign node36832 = (inp[3]) ? node36840 : node36833;
															assign node36833 = (inp[9]) ? node36837 : node36834;
																assign node36834 = (inp[12]) ? 4'b1000 : 4'b1100;
																assign node36837 = (inp[12]) ? 4'b1110 : 4'b1000;
															assign node36840 = (inp[9]) ? 4'b1110 : node36841;
																assign node36841 = (inp[12]) ? 4'b1010 : 4'b1110;
												assign node36845 = (inp[15]) ? node36865 : node36846;
													assign node36846 = (inp[5]) ? node36860 : node36847;
														assign node36847 = (inp[3]) ? node36853 : node36848;
															assign node36848 = (inp[9]) ? node36850 : 4'b1110;
																assign node36850 = (inp[12]) ? 4'b1010 : 4'b1110;
															assign node36853 = (inp[9]) ? node36857 : node36854;
																assign node36854 = (inp[12]) ? 4'b1100 : 4'b1010;
																assign node36857 = (inp[12]) ? 4'b1000 : 4'b1100;
														assign node36860 = (inp[9]) ? 4'b1000 : node36861;
															assign node36861 = (inp[12]) ? 4'b1100 : 4'b1000;
													assign node36865 = (inp[3]) ? node36877 : node36866;
														assign node36866 = (inp[5]) ? node36872 : node36867;
															assign node36867 = (inp[12]) ? node36869 : 4'b1100;
																assign node36869 = (inp[9]) ? 4'b1000 : 4'b1100;
															assign node36872 = (inp[9]) ? 4'b1110 : node36873;
																assign node36873 = (inp[12]) ? 4'b1110 : 4'b1000;
														assign node36877 = (inp[9]) ? node36883 : node36878;
															assign node36878 = (inp[12]) ? 4'b1110 : node36879;
																assign node36879 = (inp[5]) ? 4'b1010 : 4'b1000;
															assign node36883 = (inp[12]) ? 4'b1010 : 4'b1110;
											assign node36886 = (inp[4]) ? node36920 : node36887;
												assign node36887 = (inp[15]) ? node36901 : node36888;
													assign node36888 = (inp[3]) ? node36894 : node36889;
														assign node36889 = (inp[12]) ? 4'b1000 : node36890;
															assign node36890 = (inp[9]) ? 4'b1000 : 4'b1100;
														assign node36894 = (inp[5]) ? node36896 : 4'b1000;
															assign node36896 = (inp[9]) ? node36898 : 4'b1010;
																assign node36898 = (inp[12]) ? 4'b1110 : 4'b1010;
													assign node36901 = (inp[5]) ? node36913 : node36902;
														assign node36902 = (inp[3]) ? node36908 : node36903;
															assign node36903 = (inp[9]) ? node36905 : 4'b1010;
																assign node36905 = (inp[12]) ? 4'b1110 : 4'b1010;
															assign node36908 = (inp[9]) ? 4'b1100 : node36909;
																assign node36909 = (inp[12]) ? 4'b1010 : 4'b1110;
														assign node36913 = (inp[12]) ? 4'b1100 : node36914;
															assign node36914 = (inp[3]) ? node36916 : 4'b1010;
																assign node36916 = (inp[9]) ? 4'b1000 : 4'b1100;
												assign node36920 = (inp[9]) ? node36936 : node36921;
													assign node36921 = (inp[12]) ? node36931 : node36922;
														assign node36922 = (inp[3]) ? node36926 : node36923;
															assign node36923 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node36926 = (inp[15]) ? 4'b1000 : node36927;
																assign node36927 = (inp[5]) ? 4'b1010 : 4'b1000;
														assign node36931 = (inp[15]) ? node36933 : 4'b1110;
															assign node36933 = (inp[5]) ? 4'b1100 : 4'b1110;
													assign node36936 = (inp[12]) ? node36946 : node36937;
														assign node36937 = (inp[3]) ? 4'b1100 : node36938;
															assign node36938 = (inp[5]) ? node36942 : node36939;
																assign node36939 = (inp[15]) ? 4'b1110 : 4'b1100;
																assign node36942 = (inp[15]) ? 4'b1100 : 4'b1110;
														assign node36946 = (inp[15]) ? 4'b1000 : node36947;
															assign node36947 = (inp[3]) ? 4'b1010 : 4'b1000;
										assign node36951 = (inp[12]) ? node37013 : node36952;
											assign node36952 = (inp[5]) ? node36976 : node36953;
												assign node36953 = (inp[15]) ? node36963 : node36954;
													assign node36954 = (inp[0]) ? node36956 : 4'b0011;
														assign node36956 = (inp[3]) ? 4'b0001 : node36957;
															assign node36957 = (inp[9]) ? node36959 : 4'b0001;
																assign node36959 = (inp[4]) ? 4'b0101 : 4'b0001;
													assign node36963 = (inp[0]) ? node36969 : node36964;
														assign node36964 = (inp[4]) ? 4'b0001 : node36965;
															assign node36965 = (inp[9]) ? 4'b0001 : 4'b0101;
														assign node36969 = (inp[4]) ? node36973 : node36970;
															assign node36970 = (inp[9]) ? 4'b0011 : 4'b0111;
															assign node36973 = (inp[9]) ? 4'b0111 : 4'b0011;
												assign node36976 = (inp[3]) ? node37000 : node36977;
													assign node36977 = (inp[4]) ? node36993 : node36978;
														assign node36978 = (inp[9]) ? node36986 : node36979;
															assign node36979 = (inp[15]) ? node36983 : node36980;
																assign node36980 = (inp[0]) ? 4'b0101 : 4'b0111;
																assign node36983 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node36986 = (inp[15]) ? node36990 : node36987;
																assign node36987 = (inp[0]) ? 4'b0001 : 4'b0011;
																assign node36990 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node36993 = (inp[9]) ? node36995 : 4'b0001;
															assign node36995 = (inp[15]) ? 4'b0101 : node36996;
																assign node36996 = (inp[0]) ? 4'b0111 : 4'b0101;
													assign node37000 = (inp[9]) ? node37010 : node37001;
														assign node37001 = (inp[4]) ? node37003 : 4'b0101;
															assign node37003 = (inp[0]) ? node37007 : node37004;
																assign node37004 = (inp[15]) ? 4'b0011 : 4'b0001;
																assign node37007 = (inp[15]) ? 4'b0001 : 4'b0011;
														assign node37010 = (inp[4]) ? 4'b0101 : 4'b0001;
											assign node37013 = (inp[15]) ? node37051 : node37014;
												assign node37014 = (inp[0]) ? node37034 : node37015;
													assign node37015 = (inp[3]) ? node37027 : node37016;
														assign node37016 = (inp[5]) ? node37022 : node37017;
															assign node37017 = (inp[4]) ? node37019 : 4'b0111;
																assign node37019 = (inp[9]) ? 4'b0011 : 4'b0111;
															assign node37022 = (inp[9]) ? 4'b0101 : node37023;
																assign node37023 = (inp[4]) ? 4'b0101 : 4'b0011;
														assign node37027 = (inp[4]) ? node37031 : node37028;
															assign node37028 = (inp[9]) ? 4'b0101 : 4'b0011;
															assign node37031 = (inp[9]) ? 4'b0001 : 4'b0101;
													assign node37034 = (inp[3]) ? node37046 : node37035;
														assign node37035 = (inp[5]) ? node37043 : node37036;
															assign node37036 = (inp[9]) ? node37040 : node37037;
																assign node37037 = (inp[4]) ? 4'b0101 : 4'b0001;
																assign node37040 = (inp[4]) ? 4'b0001 : 4'b0101;
															assign node37043 = (inp[9]) ? 4'b0111 : 4'b0001;
														assign node37046 = (inp[4]) ? node37048 : 4'b0001;
															assign node37048 = (inp[9]) ? 4'b0011 : 4'b0111;
												assign node37051 = (inp[0]) ? node37081 : node37052;
													assign node37052 = (inp[5]) ? node37066 : node37053;
														assign node37053 = (inp[3]) ? node37059 : node37054;
															assign node37054 = (inp[9]) ? 4'b0001 : node37055;
																assign node37055 = (inp[4]) ? 4'b0101 : 4'b0001;
															assign node37059 = (inp[9]) ? node37063 : node37060;
																assign node37060 = (inp[4]) ? 4'b0111 : 4'b0001;
																assign node37063 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node37066 = (inp[3]) ? node37074 : node37067;
															assign node37067 = (inp[9]) ? node37071 : node37068;
																assign node37068 = (inp[4]) ? 4'b0111 : 4'b0001;
																assign node37071 = (inp[4]) ? 4'b0011 : 4'b0111;
															assign node37074 = (inp[9]) ? node37078 : node37075;
																assign node37075 = (inp[4]) ? 4'b0111 : 4'b0011;
																assign node37078 = (inp[4]) ? 4'b0011 : 4'b0111;
													assign node37081 = (inp[9]) ? node37089 : node37082;
														assign node37082 = (inp[4]) ? node37084 : 4'b0011;
															assign node37084 = (inp[3]) ? 4'b0101 : node37085;
																assign node37085 = (inp[5]) ? 4'b0101 : 4'b0111;
														assign node37089 = (inp[4]) ? 4'b0001 : 4'b0101;
									assign node37092 = (inp[9]) ? node37194 : node37093;
										assign node37093 = (inp[15]) ? node37145 : node37094;
											assign node37094 = (inp[0]) ? node37124 : node37095;
												assign node37095 = (inp[3]) ? node37111 : node37096;
													assign node37096 = (inp[5]) ? node37104 : node37097;
														assign node37097 = (inp[14]) ? node37099 : 4'b0111;
															assign node37099 = (inp[4]) ? node37101 : 4'b0011;
																assign node37101 = (inp[12]) ? 4'b0111 : 4'b0011;
														assign node37104 = (inp[4]) ? node37108 : node37105;
															assign node37105 = (inp[12]) ? 4'b0011 : 4'b0111;
															assign node37108 = (inp[12]) ? 4'b0101 : 4'b0011;
													assign node37111 = (inp[5]) ? node37117 : node37112;
														assign node37112 = (inp[4]) ? 4'b0101 : node37113;
															assign node37113 = (inp[12]) ? 4'b0011 : 4'b0111;
														assign node37117 = (inp[4]) ? node37121 : node37118;
															assign node37118 = (inp[12]) ? 4'b0001 : 4'b0101;
															assign node37121 = (inp[12]) ? 4'b0101 : 4'b0001;
												assign node37124 = (inp[3]) ? node37132 : node37125;
													assign node37125 = (inp[4]) ? node37129 : node37126;
														assign node37126 = (inp[12]) ? 4'b0001 : 4'b0101;
														assign node37129 = (inp[12]) ? 4'b0101 : 4'b0001;
													assign node37132 = (inp[5]) ? node37140 : node37133;
														assign node37133 = (inp[4]) ? node37137 : node37134;
															assign node37134 = (inp[12]) ? 4'b0001 : 4'b0101;
															assign node37137 = (inp[12]) ? 4'b0111 : 4'b0001;
														assign node37140 = (inp[4]) ? 4'b0111 : node37141;
															assign node37141 = (inp[12]) ? 4'b0011 : 4'b0111;
											assign node37145 = (inp[0]) ? node37175 : node37146;
												assign node37146 = (inp[5]) ? node37162 : node37147;
													assign node37147 = (inp[14]) ? node37155 : node37148;
														assign node37148 = (inp[12]) ? node37152 : node37149;
															assign node37149 = (inp[4]) ? 4'b0001 : 4'b0101;
															assign node37152 = (inp[4]) ? 4'b0101 : 4'b0001;
														assign node37155 = (inp[12]) ? node37159 : node37156;
															assign node37156 = (inp[4]) ? 4'b0001 : 4'b0101;
															assign node37159 = (inp[3]) ? 4'b0111 : 4'b0101;
													assign node37162 = (inp[3]) ? node37168 : node37163;
														assign node37163 = (inp[4]) ? 4'b0111 : node37164;
															assign node37164 = (inp[12]) ? 4'b0001 : 4'b0101;
														assign node37168 = (inp[4]) ? node37172 : node37169;
															assign node37169 = (inp[12]) ? 4'b0011 : 4'b0111;
															assign node37172 = (inp[12]) ? 4'b0111 : 4'b0011;
												assign node37175 = (inp[5]) ? node37185 : node37176;
													assign node37176 = (inp[12]) ? node37180 : node37177;
														assign node37177 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node37180 = (inp[4]) ? node37182 : 4'b0011;
															assign node37182 = (inp[3]) ? 4'b0101 : 4'b0111;
													assign node37185 = (inp[3]) ? 4'b0101 : node37186;
														assign node37186 = (inp[4]) ? node37190 : node37187;
															assign node37187 = (inp[12]) ? 4'b0011 : 4'b0111;
															assign node37190 = (inp[12]) ? 4'b0101 : 4'b0011;
										assign node37194 = (inp[14]) ? node37262 : node37195;
											assign node37195 = (inp[15]) ? node37233 : node37196;
												assign node37196 = (inp[0]) ? node37218 : node37197;
													assign node37197 = (inp[3]) ? node37207 : node37198;
														assign node37198 = (inp[5]) ? node37204 : node37199;
															assign node37199 = (inp[12]) ? node37201 : 4'b0111;
																assign node37201 = (inp[4]) ? 4'b0011 : 4'b0111;
															assign node37204 = (inp[12]) ? 4'b0101 : 4'b0011;
														assign node37207 = (inp[5]) ? node37211 : node37208;
															assign node37208 = (inp[12]) ? 4'b0001 : 4'b0011;
															assign node37211 = (inp[4]) ? node37215 : node37212;
																assign node37212 = (inp[12]) ? 4'b0101 : 4'b0001;
																assign node37215 = (inp[12]) ? 4'b0001 : 4'b0101;
													assign node37218 = (inp[5]) ? node37226 : node37219;
														assign node37219 = (inp[3]) ? 4'b0111 : node37220;
															assign node37220 = (inp[4]) ? 4'b0001 : node37221;
																assign node37221 = (inp[12]) ? 4'b0101 : 4'b0001;
														assign node37226 = (inp[4]) ? node37230 : node37227;
															assign node37227 = (inp[12]) ? 4'b0111 : 4'b0011;
															assign node37230 = (inp[12]) ? 4'b0011 : 4'b0111;
												assign node37233 = (inp[0]) ? node37251 : node37234;
													assign node37234 = (inp[12]) ? node37244 : node37235;
														assign node37235 = (inp[4]) ? node37241 : node37236;
															assign node37236 = (inp[3]) ? node37238 : 4'b0001;
																assign node37238 = (inp[5]) ? 4'b0011 : 4'b0001;
															assign node37241 = (inp[5]) ? 4'b0111 : 4'b0101;
														assign node37244 = (inp[4]) ? node37246 : 4'b0111;
															assign node37246 = (inp[3]) ? 4'b0011 : node37247;
																assign node37247 = (inp[5]) ? 4'b0011 : 4'b0001;
													assign node37251 = (inp[5]) ? node37253 : 4'b0011;
														assign node37253 = (inp[4]) ? node37259 : node37254;
															assign node37254 = (inp[12]) ? 4'b0101 : node37255;
																assign node37255 = (inp[3]) ? 4'b0001 : 4'b0011;
															assign node37259 = (inp[12]) ? 4'b0001 : 4'b0101;
											assign node37262 = (inp[5]) ? node37294 : node37263;
												assign node37263 = (inp[12]) ? node37273 : node37264;
													assign node37264 = (inp[4]) ? 4'b0101 : node37265;
														assign node37265 = (inp[15]) ? node37269 : node37266;
															assign node37266 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node37269 = (inp[0]) ? 4'b0011 : 4'b0001;
													assign node37273 = (inp[4]) ? node37285 : node37274;
														assign node37274 = (inp[3]) ? node37280 : node37275;
															assign node37275 = (inp[15]) ? 4'b0101 : node37276;
																assign node37276 = (inp[0]) ? 4'b0101 : 4'b0111;
															assign node37280 = (inp[0]) ? 4'b0111 : node37281;
																assign node37281 = (inp[15]) ? 4'b0111 : 4'b0101;
														assign node37285 = (inp[3]) ? node37287 : 4'b0001;
															assign node37287 = (inp[15]) ? node37291 : node37288;
																assign node37288 = (inp[0]) ? 4'b0011 : 4'b0001;
																assign node37291 = (inp[0]) ? 4'b0001 : 4'b0011;
												assign node37294 = (inp[3]) ? node37324 : node37295;
													assign node37295 = (inp[4]) ? node37311 : node37296;
														assign node37296 = (inp[12]) ? node37304 : node37297;
															assign node37297 = (inp[0]) ? node37301 : node37298;
																assign node37298 = (inp[15]) ? 4'b0001 : 4'b0011;
																assign node37301 = (inp[15]) ? 4'b0011 : 4'b0001;
															assign node37304 = (inp[15]) ? node37308 : node37305;
																assign node37305 = (inp[0]) ? 4'b0111 : 4'b0101;
																assign node37308 = (inp[0]) ? 4'b0101 : 4'b0111;
														assign node37311 = (inp[12]) ? node37317 : node37312;
															assign node37312 = (inp[15]) ? node37314 : 4'b0111;
																assign node37314 = (inp[0]) ? 4'b0101 : 4'b0111;
															assign node37317 = (inp[15]) ? node37321 : node37318;
																assign node37318 = (inp[0]) ? 4'b0011 : 4'b0001;
																assign node37321 = (inp[0]) ? 4'b0001 : 4'b0011;
													assign node37324 = (inp[15]) ? node37332 : node37325;
														assign node37325 = (inp[0]) ? 4'b0011 : node37326;
															assign node37326 = (inp[12]) ? node37328 : 4'b0001;
																assign node37328 = (inp[4]) ? 4'b0001 : 4'b0101;
														assign node37332 = (inp[0]) ? node37340 : node37333;
															assign node37333 = (inp[4]) ? node37337 : node37334;
																assign node37334 = (inp[12]) ? 4'b0111 : 4'b0011;
																assign node37337 = (inp[12]) ? 4'b0011 : 4'b0111;
															assign node37340 = (inp[12]) ? 4'b0001 : node37341;
																assign node37341 = (inp[4]) ? 4'b0101 : 4'b0001;
								assign node37345 = (inp[14]) ? node37605 : node37346;
									assign node37346 = (inp[2]) ? node37490 : node37347;
										assign node37347 = (inp[15]) ? node37423 : node37348;
											assign node37348 = (inp[9]) ? node37398 : node37349;
												assign node37349 = (inp[0]) ? node37369 : node37350;
													assign node37350 = (inp[3]) ? node37360 : node37351;
														assign node37351 = (inp[4]) ? node37355 : node37352;
															assign node37352 = (inp[12]) ? 4'b0011 : 4'b0111;
															assign node37355 = (inp[12]) ? node37357 : 4'b0011;
																assign node37357 = (inp[5]) ? 4'b0101 : 4'b0111;
														assign node37360 = (inp[5]) ? node37366 : node37361;
															assign node37361 = (inp[12]) ? 4'b0101 : node37362;
																assign node37362 = (inp[4]) ? 4'b0011 : 4'b0111;
															assign node37366 = (inp[4]) ? 4'b0001 : 4'b0101;
													assign node37369 = (inp[3]) ? node37385 : node37370;
														assign node37370 = (inp[5]) ? node37378 : node37371;
															assign node37371 = (inp[4]) ? node37375 : node37372;
																assign node37372 = (inp[12]) ? 4'b0001 : 4'b0101;
																assign node37375 = (inp[12]) ? 4'b0101 : 4'b0001;
															assign node37378 = (inp[4]) ? node37382 : node37379;
																assign node37379 = (inp[12]) ? 4'b0001 : 4'b0101;
																assign node37382 = (inp[12]) ? 4'b0111 : 4'b0001;
														assign node37385 = (inp[5]) ? node37393 : node37386;
															assign node37386 = (inp[12]) ? node37390 : node37387;
																assign node37387 = (inp[4]) ? 4'b0001 : 4'b0101;
																assign node37390 = (inp[4]) ? 4'b0111 : 4'b0001;
															assign node37393 = (inp[4]) ? node37395 : 4'b0111;
																assign node37395 = (inp[12]) ? 4'b0111 : 4'b0011;
												assign node37398 = (inp[0]) ? node37412 : node37399;
													assign node37399 = (inp[3]) ? node37405 : node37400;
														assign node37400 = (inp[12]) ? node37402 : 4'b0011;
															assign node37402 = (inp[4]) ? 4'b0001 : 4'b0101;
														assign node37405 = (inp[12]) ? node37409 : node37406;
															assign node37406 = (inp[4]) ? 4'b0101 : 4'b0001;
															assign node37409 = (inp[4]) ? 4'b0001 : 4'b0101;
													assign node37412 = (inp[4]) ? node37418 : node37413;
														assign node37413 = (inp[12]) ? node37415 : 4'b0001;
															assign node37415 = (inp[3]) ? 4'b0111 : 4'b0101;
														assign node37418 = (inp[12]) ? node37420 : 4'b0111;
															assign node37420 = (inp[5]) ? 4'b0011 : 4'b0001;
											assign node37423 = (inp[0]) ? node37463 : node37424;
												assign node37424 = (inp[3]) ? node37446 : node37425;
													assign node37425 = (inp[5]) ? node37435 : node37426;
														assign node37426 = (inp[12]) ? node37428 : 4'b0101;
															assign node37428 = (inp[4]) ? node37432 : node37429;
																assign node37429 = (inp[9]) ? 4'b0101 : 4'b0001;
																assign node37432 = (inp[9]) ? 4'b0001 : 4'b0101;
														assign node37435 = (inp[4]) ? node37439 : node37436;
															assign node37436 = (inp[12]) ? 4'b0001 : 4'b0101;
															assign node37439 = (inp[12]) ? node37443 : node37440;
																assign node37440 = (inp[9]) ? 4'b0111 : 4'b0001;
																assign node37443 = (inp[9]) ? 4'b0011 : 4'b0111;
													assign node37446 = (inp[12]) ? node37456 : node37447;
														assign node37447 = (inp[4]) ? node37453 : node37448;
															assign node37448 = (inp[5]) ? 4'b0011 : node37449;
																assign node37449 = (inp[9]) ? 4'b0001 : 4'b0101;
															assign node37453 = (inp[9]) ? 4'b0111 : 4'b0011;
														assign node37456 = (inp[9]) ? node37460 : node37457;
															assign node37457 = (inp[4]) ? 4'b0111 : 4'b0011;
															assign node37460 = (inp[4]) ? 4'b0011 : 4'b0111;
												assign node37463 = (inp[5]) ? node37483 : node37464;
													assign node37464 = (inp[3]) ? node37476 : node37465;
														assign node37465 = (inp[12]) ? node37471 : node37466;
															assign node37466 = (inp[4]) ? node37468 : 4'b0111;
																assign node37468 = (inp[9]) ? 4'b0111 : 4'b0011;
															assign node37471 = (inp[9]) ? 4'b0011 : node37472;
																assign node37472 = (inp[4]) ? 4'b0111 : 4'b0011;
														assign node37476 = (inp[9]) ? node37478 : 4'b0011;
															assign node37478 = (inp[4]) ? node37480 : 4'b0011;
																assign node37480 = (inp[12]) ? 4'b0001 : 4'b0101;
													assign node37483 = (inp[3]) ? 4'b0101 : node37484;
														assign node37484 = (inp[4]) ? node37486 : 4'b0011;
															assign node37486 = (inp[12]) ? 4'b0101 : 4'b0011;
										assign node37490 = (inp[12]) ? node37550 : node37491;
											assign node37491 = (inp[5]) ? node37523 : node37492;
												assign node37492 = (inp[4]) ? node37504 : node37493;
													assign node37493 = (inp[9]) ? node37501 : node37494;
														assign node37494 = (inp[3]) ? 4'b0100 : node37495;
															assign node37495 = (inp[15]) ? node37497 : 4'b0100;
																assign node37497 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node37501 = (inp[15]) ? 4'b0010 : 4'b0000;
													assign node37504 = (inp[9]) ? node37512 : node37505;
														assign node37505 = (inp[15]) ? node37509 : node37506;
															assign node37506 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node37509 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node37512 = (inp[0]) ? node37518 : node37513;
															assign node37513 = (inp[15]) ? node37515 : 4'b0110;
																assign node37515 = (inp[3]) ? 4'b0110 : 4'b0100;
															assign node37518 = (inp[15]) ? 4'b0100 : node37519;
																assign node37519 = (inp[3]) ? 4'b0110 : 4'b0100;
												assign node37523 = (inp[4]) ? node37543 : node37524;
													assign node37524 = (inp[9]) ? node37534 : node37525;
														assign node37525 = (inp[3]) ? node37527 : 4'b0100;
															assign node37527 = (inp[0]) ? node37531 : node37528;
																assign node37528 = (inp[15]) ? 4'b0110 : 4'b0100;
																assign node37531 = (inp[15]) ? 4'b0100 : 4'b0110;
														assign node37534 = (inp[15]) ? 4'b0010 : node37535;
															assign node37535 = (inp[0]) ? node37539 : node37536;
																assign node37536 = (inp[3]) ? 4'b0000 : 4'b0010;
																assign node37539 = (inp[3]) ? 4'b0010 : 4'b0000;
													assign node37543 = (inp[9]) ? node37545 : 4'b0010;
														assign node37545 = (inp[3]) ? 4'b0110 : node37546;
															assign node37546 = (inp[0]) ? 4'b0110 : 4'b0100;
											assign node37550 = (inp[0]) ? node37578 : node37551;
												assign node37551 = (inp[15]) ? node37563 : node37552;
													assign node37552 = (inp[9]) ? node37558 : node37553;
														assign node37553 = (inp[4]) ? node37555 : 4'b0010;
															assign node37555 = (inp[5]) ? 4'b0100 : 4'b0110;
														assign node37558 = (inp[4]) ? node37560 : 4'b0100;
															assign node37560 = (inp[5]) ? 4'b0000 : 4'b0010;
													assign node37563 = (inp[3]) ? node37573 : node37564;
														assign node37564 = (inp[5]) ? 4'b0000 : node37565;
															assign node37565 = (inp[4]) ? node37569 : node37566;
																assign node37566 = (inp[9]) ? 4'b0100 : 4'b0000;
																assign node37569 = (inp[9]) ? 4'b0000 : 4'b0100;
														assign node37573 = (inp[9]) ? node37575 : 4'b0000;
															assign node37575 = (inp[5]) ? 4'b0010 : 4'b0110;
												assign node37578 = (inp[9]) ? node37590 : node37579;
													assign node37579 = (inp[4]) ? node37583 : node37580;
														assign node37580 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node37583 = (inp[3]) ? 4'b0110 : node37584;
															assign node37584 = (inp[5]) ? 4'b0100 : node37585;
																assign node37585 = (inp[15]) ? 4'b0110 : 4'b0100;
													assign node37590 = (inp[4]) ? node37598 : node37591;
														assign node37591 = (inp[15]) ? node37593 : 4'b0110;
															assign node37593 = (inp[3]) ? 4'b0100 : node37594;
																assign node37594 = (inp[5]) ? 4'b0100 : 4'b0110;
														assign node37598 = (inp[5]) ? 4'b0010 : node37599;
															assign node37599 = (inp[3]) ? 4'b0000 : node37600;
																assign node37600 = (inp[15]) ? 4'b0010 : 4'b0000;
									assign node37605 = (inp[3]) ? node37767 : node37606;
										assign node37606 = (inp[5]) ? node37698 : node37607;
											assign node37607 = (inp[2]) ? node37655 : node37608;
												assign node37608 = (inp[0]) ? node37630 : node37609;
													assign node37609 = (inp[15]) ? node37625 : node37610;
														assign node37610 = (inp[9]) ? node37618 : node37611;
															assign node37611 = (inp[4]) ? node37615 : node37612;
																assign node37612 = (inp[12]) ? 4'b0010 : 4'b0110;
																assign node37615 = (inp[12]) ? 4'b0110 : 4'b0010;
															assign node37618 = (inp[4]) ? node37622 : node37619;
																assign node37619 = (inp[12]) ? 4'b0110 : 4'b0010;
																assign node37622 = (inp[12]) ? 4'b0010 : 4'b0110;
														assign node37625 = (inp[12]) ? node37627 : 4'b0100;
															assign node37627 = (inp[4]) ? 4'b0100 : 4'b0000;
													assign node37630 = (inp[15]) ? node37642 : node37631;
														assign node37631 = (inp[9]) ? node37637 : node37632;
															assign node37632 = (inp[4]) ? 4'b0000 : node37633;
																assign node37633 = (inp[12]) ? 4'b0000 : 4'b0100;
															assign node37637 = (inp[12]) ? 4'b0100 : node37638;
																assign node37638 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node37642 = (inp[9]) ? node37650 : node37643;
															assign node37643 = (inp[4]) ? node37647 : node37644;
																assign node37644 = (inp[12]) ? 4'b0010 : 4'b0110;
																assign node37647 = (inp[12]) ? 4'b0110 : 4'b0010;
															assign node37650 = (inp[12]) ? 4'b0010 : node37651;
																assign node37651 = (inp[4]) ? 4'b0110 : 4'b0010;
												assign node37655 = (inp[12]) ? node37679 : node37656;
													assign node37656 = (inp[9]) ? node37666 : node37657;
														assign node37657 = (inp[4]) ? node37661 : node37658;
															assign node37658 = (inp[0]) ? 4'b0100 : 4'b0110;
															assign node37661 = (inp[0]) ? 4'b0010 : node37662;
																assign node37662 = (inp[15]) ? 4'b0000 : 4'b0010;
														assign node37666 = (inp[4]) ? node37674 : node37667;
															assign node37667 = (inp[0]) ? node37671 : node37668;
																assign node37668 = (inp[15]) ? 4'b0000 : 4'b0010;
																assign node37671 = (inp[15]) ? 4'b0010 : 4'b0000;
															assign node37674 = (inp[15]) ? node37676 : 4'b0100;
																assign node37676 = (inp[0]) ? 4'b0110 : 4'b0100;
													assign node37679 = (inp[15]) ? node37691 : node37680;
														assign node37680 = (inp[0]) ? node37688 : node37681;
															assign node37681 = (inp[4]) ? node37685 : node37682;
																assign node37682 = (inp[9]) ? 4'b0110 : 4'b0010;
																assign node37685 = (inp[9]) ? 4'b0010 : 4'b0110;
															assign node37688 = (inp[9]) ? 4'b0000 : 4'b0100;
														assign node37691 = (inp[0]) ? 4'b0110 : node37692;
															assign node37692 = (inp[9]) ? node37694 : 4'b0100;
																assign node37694 = (inp[4]) ? 4'b0000 : 4'b0100;
											assign node37698 = (inp[4]) ? node37724 : node37699;
												assign node37699 = (inp[9]) ? node37713 : node37700;
													assign node37700 = (inp[12]) ? node37708 : node37701;
														assign node37701 = (inp[15]) ? node37705 : node37702;
															assign node37702 = (inp[0]) ? 4'b0100 : 4'b0110;
															assign node37705 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node37708 = (inp[2]) ? node37710 : 4'b0000;
															assign node37710 = (inp[0]) ? 4'b0010 : 4'b0000;
													assign node37713 = (inp[12]) ? node37721 : node37714;
														assign node37714 = (inp[15]) ? node37718 : node37715;
															assign node37715 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node37718 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node37721 = (inp[0]) ? 4'b0100 : 4'b0110;
												assign node37724 = (inp[2]) ? node37744 : node37725;
													assign node37725 = (inp[0]) ? node37737 : node37726;
														assign node37726 = (inp[9]) ? node37732 : node37727;
															assign node37727 = (inp[12]) ? 4'b0110 : node37728;
																assign node37728 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node37732 = (inp[12]) ? 4'b0000 : node37733;
																assign node37733 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node37737 = (inp[9]) ? 4'b0010 : node37738;
															assign node37738 = (inp[12]) ? node37740 : 4'b0010;
																assign node37740 = (inp[15]) ? 4'b0100 : 4'b0110;
													assign node37744 = (inp[9]) ? node37754 : node37745;
														assign node37745 = (inp[12]) ? node37747 : 4'b0000;
															assign node37747 = (inp[15]) ? node37751 : node37748;
																assign node37748 = (inp[0]) ? 4'b0110 : 4'b0100;
																assign node37751 = (inp[0]) ? 4'b0100 : 4'b0110;
														assign node37754 = (inp[12]) ? node37762 : node37755;
															assign node37755 = (inp[0]) ? node37759 : node37756;
																assign node37756 = (inp[15]) ? 4'b0110 : 4'b0100;
																assign node37759 = (inp[15]) ? 4'b0100 : 4'b0110;
															assign node37762 = (inp[15]) ? 4'b0000 : node37763;
																assign node37763 = (inp[0]) ? 4'b0010 : 4'b0000;
										assign node37767 = (inp[0]) ? node37815 : node37768;
											assign node37768 = (inp[15]) ? node37788 : node37769;
												assign node37769 = (inp[9]) ? node37781 : node37770;
													assign node37770 = (inp[5]) ? node37778 : node37771;
														assign node37771 = (inp[4]) ? node37775 : node37772;
															assign node37772 = (inp[12]) ? 4'b0010 : 4'b0110;
															assign node37775 = (inp[12]) ? 4'b0100 : 4'b0010;
														assign node37778 = (inp[12]) ? 4'b0000 : 4'b0100;
													assign node37781 = (inp[12]) ? node37785 : node37782;
														assign node37782 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node37785 = (inp[4]) ? 4'b0000 : 4'b0100;
												assign node37788 = (inp[5]) ? node37804 : node37789;
													assign node37789 = (inp[9]) ? node37797 : node37790;
														assign node37790 = (inp[4]) ? node37794 : node37791;
															assign node37791 = (inp[12]) ? 4'b0000 : 4'b0100;
															assign node37794 = (inp[2]) ? 4'b0110 : 4'b0000;
														assign node37797 = (inp[12]) ? node37801 : node37798;
															assign node37798 = (inp[4]) ? 4'b0110 : 4'b0000;
															assign node37801 = (inp[4]) ? 4'b0010 : 4'b0110;
													assign node37804 = (inp[12]) ? node37812 : node37805;
														assign node37805 = (inp[4]) ? node37809 : node37806;
															assign node37806 = (inp[9]) ? 4'b0010 : 4'b0110;
															assign node37809 = (inp[9]) ? 4'b0110 : 4'b0010;
														assign node37812 = (inp[2]) ? 4'b0010 : 4'b0110;
											assign node37815 = (inp[15]) ? node37843 : node37816;
												assign node37816 = (inp[5]) ? node37830 : node37817;
													assign node37817 = (inp[9]) ? node37823 : node37818;
														assign node37818 = (inp[4]) ? 4'b0000 : node37819;
															assign node37819 = (inp[12]) ? 4'b0000 : 4'b0100;
														assign node37823 = (inp[12]) ? node37827 : node37824;
															assign node37824 = (inp[4]) ? 4'b0110 : 4'b0000;
															assign node37827 = (inp[4]) ? 4'b0010 : 4'b0110;
													assign node37830 = (inp[4]) ? 4'b0010 : node37831;
														assign node37831 = (inp[2]) ? node37837 : node37832;
															assign node37832 = (inp[12]) ? 4'b0010 : node37833;
																assign node37833 = (inp[9]) ? 4'b0010 : 4'b0110;
															assign node37837 = (inp[9]) ? 4'b0110 : node37838;
																assign node37838 = (inp[12]) ? 4'b0010 : 4'b0110;
												assign node37843 = (inp[5]) ? node37857 : node37844;
													assign node37844 = (inp[4]) ? node37850 : node37845;
														assign node37845 = (inp[9]) ? 4'b0010 : node37846;
															assign node37846 = (inp[12]) ? 4'b0010 : 4'b0110;
														assign node37850 = (inp[12]) ? node37854 : node37851;
															assign node37851 = (inp[9]) ? 4'b0100 : 4'b0010;
															assign node37854 = (inp[9]) ? 4'b0000 : 4'b0100;
													assign node37857 = (inp[12]) ? node37865 : node37858;
														assign node37858 = (inp[2]) ? 4'b0100 : node37859;
															assign node37859 = (inp[4]) ? 4'b0000 : node37860;
																assign node37860 = (inp[9]) ? 4'b0000 : 4'b0100;
														assign node37865 = (inp[9]) ? 4'b0000 : node37866;
															assign node37866 = (inp[4]) ? 4'b0100 : 4'b0000;
						assign node37870 = (inp[5]) ? node38976 : node37871;
							assign node37871 = (inp[14]) ? node38453 : node37872;
								assign node37872 = (inp[8]) ? node38174 : node37873;
									assign node37873 = (inp[9]) ? node37997 : node37874;
										assign node37874 = (inp[0]) ? node37934 : node37875;
											assign node37875 = (inp[15]) ? node37897 : node37876;
												assign node37876 = (inp[2]) ? node37890 : node37877;
													assign node37877 = (inp[7]) ? node37885 : node37878;
														assign node37878 = (inp[12]) ? node37882 : node37879;
															assign node37879 = (inp[4]) ? 4'b0011 : 4'b0111;
															assign node37882 = (inp[4]) ? 4'b0101 : 4'b0011;
														assign node37885 = (inp[12]) ? 4'b0010 : node37886;
															assign node37886 = (inp[4]) ? 4'b0010 : 4'b0110;
													assign node37890 = (inp[7]) ? node37892 : 4'b0010;
														assign node37892 = (inp[4]) ? node37894 : 4'b0011;
															assign node37894 = (inp[12]) ? 4'b0111 : 4'b0011;
												assign node37897 = (inp[3]) ? node37919 : node37898;
													assign node37898 = (inp[7]) ? node37910 : node37899;
														assign node37899 = (inp[2]) ? node37903 : node37900;
															assign node37900 = (inp[4]) ? 4'b0101 : 4'b0001;
															assign node37903 = (inp[4]) ? node37907 : node37904;
																assign node37904 = (inp[12]) ? 4'b0000 : 4'b0100;
																assign node37907 = (inp[12]) ? 4'b0100 : 4'b0000;
														assign node37910 = (inp[2]) ? node37914 : node37911;
															assign node37911 = (inp[12]) ? 4'b0000 : 4'b0100;
															assign node37914 = (inp[4]) ? node37916 : 4'b0101;
																assign node37916 = (inp[12]) ? 4'b0101 : 4'b0001;
													assign node37919 = (inp[12]) ? node37925 : node37920;
														assign node37920 = (inp[7]) ? node37922 : 4'b0000;
															assign node37922 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node37925 = (inp[4]) ? node37927 : 4'b0001;
															assign node37927 = (inp[7]) ? node37931 : node37928;
																assign node37928 = (inp[2]) ? 4'b0110 : 4'b0111;
																assign node37931 = (inp[2]) ? 4'b0111 : 4'b0110;
											assign node37934 = (inp[15]) ? node37962 : node37935;
												assign node37935 = (inp[3]) ? node37945 : node37936;
													assign node37936 = (inp[2]) ? node37942 : node37937;
														assign node37937 = (inp[4]) ? 4'b0001 : node37938;
															assign node37938 = (inp[12]) ? 4'b0001 : 4'b0101;
														assign node37942 = (inp[12]) ? 4'b0101 : 4'b0001;
													assign node37945 = (inp[12]) ? node37953 : node37946;
														assign node37946 = (inp[4]) ? node37948 : 4'b0101;
															assign node37948 = (inp[2]) ? node37950 : 4'b0001;
																assign node37950 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node37953 = (inp[4]) ? node37959 : node37954;
															assign node37954 = (inp[2]) ? 4'b0000 : node37955;
																assign node37955 = (inp[7]) ? 4'b0000 : 4'b0001;
															assign node37959 = (inp[2]) ? 4'b0110 : 4'b0111;
												assign node37962 = (inp[3]) ? node37984 : node37963;
													assign node37963 = (inp[12]) ? node37971 : node37964;
														assign node37964 = (inp[4]) ? node37966 : 4'b0110;
															assign node37966 = (inp[7]) ? node37968 : 4'b0011;
																assign node37968 = (inp[2]) ? 4'b0011 : 4'b0010;
														assign node37971 = (inp[4]) ? node37977 : node37972;
															assign node37972 = (inp[2]) ? 4'b0011 : node37973;
																assign node37973 = (inp[7]) ? 4'b0010 : 4'b0011;
															assign node37977 = (inp[7]) ? node37981 : node37978;
																assign node37978 = (inp[2]) ? 4'b0110 : 4'b0111;
																assign node37981 = (inp[2]) ? 4'b0111 : 4'b0110;
													assign node37984 = (inp[12]) ? node37992 : node37985;
														assign node37985 = (inp[4]) ? node37987 : 4'b0111;
															assign node37987 = (inp[2]) ? 4'b0011 : node37988;
																assign node37988 = (inp[7]) ? 4'b0010 : 4'b0011;
														assign node37992 = (inp[4]) ? 4'b0101 : node37993;
															assign node37993 = (inp[7]) ? 4'b0010 : 4'b0011;
										assign node37997 = (inp[15]) ? node38093 : node37998;
											assign node37998 = (inp[0]) ? node38040 : node37999;
												assign node37999 = (inp[3]) ? node38019 : node38000;
													assign node38000 = (inp[7]) ? node38010 : node38001;
														assign node38001 = (inp[2]) ? node38005 : node38002;
															assign node38002 = (inp[4]) ? 4'b0011 : 4'b0111;
															assign node38005 = (inp[4]) ? node38007 : 4'b0010;
																assign node38007 = (inp[12]) ? 4'b0010 : 4'b0110;
														assign node38010 = (inp[2]) ? node38012 : 4'b0010;
															assign node38012 = (inp[12]) ? node38016 : node38013;
																assign node38013 = (inp[4]) ? 4'b0111 : 4'b0011;
																assign node38016 = (inp[4]) ? 4'b0011 : 4'b0111;
													assign node38019 = (inp[12]) ? node38029 : node38020;
														assign node38020 = (inp[4]) ? node38026 : node38021;
															assign node38021 = (inp[7]) ? 4'b0010 : node38022;
																assign node38022 = (inp[2]) ? 4'b0010 : 4'b0011;
															assign node38026 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node38029 = (inp[4]) ? node38037 : node38030;
															assign node38030 = (inp[2]) ? node38034 : node38031;
																assign node38031 = (inp[7]) ? 4'b0100 : 4'b0101;
																assign node38034 = (inp[7]) ? 4'b0101 : 4'b0100;
															assign node38037 = (inp[7]) ? 4'b0000 : 4'b0001;
												assign node38040 = (inp[3]) ? node38064 : node38041;
													assign node38041 = (inp[7]) ? node38053 : node38042;
														assign node38042 = (inp[2]) ? node38050 : node38043;
															assign node38043 = (inp[4]) ? node38047 : node38044;
																assign node38044 = (inp[12]) ? 4'b0101 : 4'b0001;
																assign node38047 = (inp[12]) ? 4'b0001 : 4'b0101;
															assign node38050 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node38053 = (inp[2]) ? node38061 : node38054;
															assign node38054 = (inp[12]) ? node38058 : node38055;
																assign node38055 = (inp[4]) ? 4'b0100 : 4'b0000;
																assign node38058 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node38061 = (inp[12]) ? 4'b0101 : 4'b0001;
													assign node38064 = (inp[4]) ? node38080 : node38065;
														assign node38065 = (inp[12]) ? node38073 : node38066;
															assign node38066 = (inp[7]) ? node38070 : node38067;
																assign node38067 = (inp[2]) ? 4'b0000 : 4'b0001;
																assign node38070 = (inp[2]) ? 4'b0001 : 4'b0000;
															assign node38073 = (inp[2]) ? node38077 : node38074;
																assign node38074 = (inp[7]) ? 4'b0110 : 4'b0111;
																assign node38077 = (inp[7]) ? 4'b0111 : 4'b0110;
														assign node38080 = (inp[12]) ? node38088 : node38081;
															assign node38081 = (inp[7]) ? node38085 : node38082;
																assign node38082 = (inp[2]) ? 4'b0110 : 4'b0111;
																assign node38085 = (inp[2]) ? 4'b0111 : 4'b0110;
															assign node38088 = (inp[2]) ? 4'b0010 : node38089;
																assign node38089 = (inp[7]) ? 4'b0010 : 4'b0011;
											assign node38093 = (inp[0]) ? node38129 : node38094;
												assign node38094 = (inp[3]) ? node38108 : node38095;
													assign node38095 = (inp[4]) ? node38103 : node38096;
														assign node38096 = (inp[12]) ? 4'b0100 : node38097;
															assign node38097 = (inp[7]) ? 4'b0000 : node38098;
																assign node38098 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node38103 = (inp[12]) ? node38105 : 4'b0101;
															assign node38105 = (inp[2]) ? 4'b0000 : 4'b0001;
													assign node38108 = (inp[4]) ? node38118 : node38109;
														assign node38109 = (inp[12]) ? node38115 : node38110;
															assign node38110 = (inp[7]) ? node38112 : 4'b0001;
																assign node38112 = (inp[2]) ? 4'b0001 : 4'b0000;
															assign node38115 = (inp[2]) ? 4'b0111 : 4'b0110;
														assign node38118 = (inp[12]) ? node38124 : node38119;
															assign node38119 = (inp[2]) ? 4'b0110 : node38120;
																assign node38120 = (inp[7]) ? 4'b0110 : 4'b0111;
															assign node38124 = (inp[7]) ? 4'b0010 : node38125;
																assign node38125 = (inp[2]) ? 4'b0010 : 4'b0011;
												assign node38129 = (inp[3]) ? node38157 : node38130;
													assign node38130 = (inp[2]) ? node38142 : node38131;
														assign node38131 = (inp[7]) ? node38137 : node38132;
															assign node38132 = (inp[12]) ? 4'b0011 : node38133;
																assign node38133 = (inp[4]) ? 4'b0111 : 4'b0011;
															assign node38137 = (inp[4]) ? 4'b0010 : node38138;
																assign node38138 = (inp[12]) ? 4'b0110 : 4'b0010;
														assign node38142 = (inp[7]) ? node38150 : node38143;
															assign node38143 = (inp[4]) ? node38147 : node38144;
																assign node38144 = (inp[12]) ? 4'b0110 : 4'b0010;
																assign node38147 = (inp[12]) ? 4'b0010 : 4'b0110;
															assign node38150 = (inp[4]) ? node38154 : node38151;
																assign node38151 = (inp[12]) ? 4'b0111 : 4'b0011;
																assign node38154 = (inp[12]) ? 4'b0011 : 4'b0111;
													assign node38157 = (inp[4]) ? node38165 : node38158;
														assign node38158 = (inp[12]) ? 4'b0100 : node38159;
															assign node38159 = (inp[2]) ? 4'b0010 : node38160;
																assign node38160 = (inp[7]) ? 4'b0010 : 4'b0011;
														assign node38165 = (inp[12]) ? node38167 : 4'b0100;
															assign node38167 = (inp[2]) ? node38171 : node38168;
																assign node38168 = (inp[7]) ? 4'b0000 : 4'b0001;
																assign node38171 = (inp[7]) ? 4'b0001 : 4'b0000;
									assign node38174 = (inp[3]) ? node38312 : node38175;
										assign node38175 = (inp[7]) ? node38251 : node38176;
											assign node38176 = (inp[2]) ? node38220 : node38177;
												assign node38177 = (inp[9]) ? node38199 : node38178;
													assign node38178 = (inp[0]) ? node38186 : node38179;
														assign node38179 = (inp[15]) ? 4'b0100 : node38180;
															assign node38180 = (inp[12]) ? 4'b0110 : node38181;
																assign node38181 = (inp[4]) ? 4'b0010 : 4'b0110;
														assign node38186 = (inp[15]) ? node38194 : node38187;
															assign node38187 = (inp[4]) ? node38191 : node38188;
																assign node38188 = (inp[12]) ? 4'b0000 : 4'b0100;
																assign node38191 = (inp[12]) ? 4'b0100 : 4'b0000;
															assign node38194 = (inp[4]) ? node38196 : 4'b0010;
																assign node38196 = (inp[12]) ? 4'b0110 : 4'b0010;
													assign node38199 = (inp[15]) ? node38207 : node38200;
														assign node38200 = (inp[0]) ? node38202 : 4'b0010;
															assign node38202 = (inp[4]) ? 4'b0000 : node38203;
																assign node38203 = (inp[12]) ? 4'b0100 : 4'b0000;
														assign node38207 = (inp[0]) ? node38215 : node38208;
															assign node38208 = (inp[4]) ? node38212 : node38209;
																assign node38209 = (inp[12]) ? 4'b0100 : 4'b0000;
																assign node38212 = (inp[12]) ? 4'b0000 : 4'b0100;
															assign node38215 = (inp[12]) ? node38217 : 4'b0010;
																assign node38217 = (inp[4]) ? 4'b0010 : 4'b0110;
												assign node38220 = (inp[4]) ? node38234 : node38221;
													assign node38221 = (inp[15]) ? node38229 : node38222;
														assign node38222 = (inp[0]) ? 4'b0101 : node38223;
															assign node38223 = (inp[9]) ? 4'b0111 : node38224;
																assign node38224 = (inp[12]) ? 4'b0011 : 4'b0111;
														assign node38229 = (inp[0]) ? node38231 : 4'b0001;
															assign node38231 = (inp[9]) ? 4'b0011 : 4'b0111;
													assign node38234 = (inp[15]) ? node38238 : node38235;
														assign node38235 = (inp[0]) ? 4'b0001 : 4'b0011;
														assign node38238 = (inp[0]) ? node38244 : node38239;
															assign node38239 = (inp[9]) ? 4'b0101 : node38240;
																assign node38240 = (inp[12]) ? 4'b0101 : 4'b0001;
															assign node38244 = (inp[12]) ? node38248 : node38245;
																assign node38245 = (inp[9]) ? 4'b0111 : 4'b0011;
																assign node38248 = (inp[9]) ? 4'b0011 : 4'b0111;
											assign node38251 = (inp[2]) ? node38277 : node38252;
												assign node38252 = (inp[12]) ? node38262 : node38253;
													assign node38253 = (inp[4]) ? node38257 : node38254;
														assign node38254 = (inp[0]) ? 4'b0101 : 4'b0001;
														assign node38257 = (inp[0]) ? node38259 : 4'b0001;
															assign node38259 = (inp[15]) ? 4'b0011 : 4'b0001;
													assign node38262 = (inp[9]) ? node38272 : node38263;
														assign node38263 = (inp[4]) ? node38267 : node38264;
															assign node38264 = (inp[15]) ? 4'b0011 : 4'b0001;
															assign node38267 = (inp[0]) ? node38269 : 4'b0111;
																assign node38269 = (inp[15]) ? 4'b0111 : 4'b0101;
														assign node38272 = (inp[4]) ? 4'b0001 : node38273;
															assign node38273 = (inp[15]) ? 4'b0101 : 4'b0111;
												assign node38277 = (inp[4]) ? node38293 : node38278;
													assign node38278 = (inp[12]) ? node38282 : node38279;
														assign node38279 = (inp[9]) ? 4'b0000 : 4'b0100;
														assign node38282 = (inp[9]) ? node38290 : node38283;
															assign node38283 = (inp[15]) ? node38287 : node38284;
																assign node38284 = (inp[0]) ? 4'b0000 : 4'b0010;
																assign node38287 = (inp[0]) ? 4'b0010 : 4'b0000;
															assign node38290 = (inp[15]) ? 4'b0110 : 4'b0100;
													assign node38293 = (inp[15]) ? node38305 : node38294;
														assign node38294 = (inp[0]) ? node38300 : node38295;
															assign node38295 = (inp[9]) ? 4'b0110 : node38296;
																assign node38296 = (inp[12]) ? 4'b0110 : 4'b0010;
															assign node38300 = (inp[12]) ? node38302 : 4'b0100;
																assign node38302 = (inp[9]) ? 4'b0000 : 4'b0100;
														assign node38305 = (inp[9]) ? node38309 : node38306;
															assign node38306 = (inp[12]) ? 4'b0100 : 4'b0000;
															assign node38309 = (inp[12]) ? 4'b0000 : 4'b0100;
										assign node38312 = (inp[2]) ? node38382 : node38313;
											assign node38313 = (inp[7]) ? node38341 : node38314;
												assign node38314 = (inp[12]) ? node38330 : node38315;
													assign node38315 = (inp[9]) ? node38323 : node38316;
														assign node38316 = (inp[4]) ? 4'b0010 : node38317;
															assign node38317 = (inp[0]) ? node38319 : 4'b0100;
																assign node38319 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node38323 = (inp[4]) ? node38325 : 4'b0000;
															assign node38325 = (inp[15]) ? 4'b0100 : node38326;
																assign node38326 = (inp[0]) ? 4'b0110 : 4'b0100;
													assign node38330 = (inp[15]) ? 4'b0010 : node38331;
														assign node38331 = (inp[4]) ? node38337 : node38332;
															assign node38332 = (inp[9]) ? 4'b0110 : node38333;
																assign node38333 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node38337 = (inp[9]) ? 4'b0000 : 4'b0100;
												assign node38341 = (inp[9]) ? node38365 : node38342;
													assign node38342 = (inp[0]) ? node38350 : node38343;
														assign node38343 = (inp[15]) ? node38345 : 4'b0111;
															assign node38345 = (inp[12]) ? 4'b0111 : node38346;
																assign node38346 = (inp[4]) ? 4'b0001 : 4'b0101;
														assign node38350 = (inp[15]) ? node38358 : node38351;
															assign node38351 = (inp[12]) ? node38355 : node38352;
																assign node38352 = (inp[4]) ? 4'b0001 : 4'b0101;
																assign node38355 = (inp[4]) ? 4'b0111 : 4'b0001;
															assign node38358 = (inp[4]) ? node38362 : node38359;
																assign node38359 = (inp[12]) ? 4'b0011 : 4'b0111;
																assign node38362 = (inp[12]) ? 4'b0101 : 4'b0011;
													assign node38365 = (inp[4]) ? node38373 : node38366;
														assign node38366 = (inp[12]) ? node38368 : 4'b0011;
															assign node38368 = (inp[0]) ? 4'b0111 : node38369;
																assign node38369 = (inp[15]) ? 4'b0111 : 4'b0101;
														assign node38373 = (inp[12]) ? 4'b0011 : node38374;
															assign node38374 = (inp[0]) ? node38378 : node38375;
																assign node38375 = (inp[15]) ? 4'b0111 : 4'b0101;
																assign node38378 = (inp[15]) ? 4'b0101 : 4'b0111;
											assign node38382 = (inp[7]) ? node38408 : node38383;
												assign node38383 = (inp[12]) ? node38401 : node38384;
													assign node38384 = (inp[0]) ? node38394 : node38385;
														assign node38385 = (inp[15]) ? node38391 : node38386;
															assign node38386 = (inp[4]) ? 4'b0011 : node38387;
																assign node38387 = (inp[9]) ? 4'b0011 : 4'b0111;
															assign node38391 = (inp[4]) ? 4'b0111 : 4'b0001;
														assign node38394 = (inp[15]) ? node38396 : 4'b0001;
															assign node38396 = (inp[4]) ? 4'b0011 : node38397;
																assign node38397 = (inp[9]) ? 4'b0011 : 4'b0111;
													assign node38401 = (inp[9]) ? node38405 : node38402;
														assign node38402 = (inp[4]) ? 4'b0111 : 4'b0011;
														assign node38405 = (inp[0]) ? 4'b0111 : 4'b0101;
												assign node38408 = (inp[0]) ? node38432 : node38409;
													assign node38409 = (inp[9]) ? node38421 : node38410;
														assign node38410 = (inp[4]) ? node38416 : node38411;
															assign node38411 = (inp[15]) ? 4'b0000 : node38412;
																assign node38412 = (inp[12]) ? 4'b0010 : 4'b0110;
															assign node38416 = (inp[12]) ? node38418 : 4'b0000;
																assign node38418 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node38421 = (inp[15]) ? node38425 : node38422;
															assign node38422 = (inp[12]) ? 4'b0000 : 4'b0010;
															assign node38425 = (inp[12]) ? node38429 : node38426;
																assign node38426 = (inp[4]) ? 4'b0110 : 4'b0000;
																assign node38429 = (inp[4]) ? 4'b0010 : 4'b0110;
													assign node38432 = (inp[4]) ? node38444 : node38433;
														assign node38433 = (inp[12]) ? node38439 : node38434;
															assign node38434 = (inp[9]) ? 4'b0010 : node38435;
																assign node38435 = (inp[15]) ? 4'b0110 : 4'b0100;
															assign node38439 = (inp[9]) ? node38441 : 4'b0000;
																assign node38441 = (inp[15]) ? 4'b0100 : 4'b0110;
														assign node38444 = (inp[9]) ? node38450 : node38445;
															assign node38445 = (inp[12]) ? 4'b0110 : node38446;
																assign node38446 = (inp[15]) ? 4'b0010 : 4'b0000;
															assign node38450 = (inp[12]) ? 4'b0000 : 4'b0100;
								assign node38453 = (inp[0]) ? node38723 : node38454;
									assign node38454 = (inp[15]) ? node38588 : node38455;
										assign node38455 = (inp[3]) ? node38521 : node38456;
											assign node38456 = (inp[12]) ? node38494 : node38457;
												assign node38457 = (inp[7]) ? node38477 : node38458;
													assign node38458 = (inp[8]) ? node38470 : node38459;
														assign node38459 = (inp[2]) ? node38465 : node38460;
															assign node38460 = (inp[4]) ? 4'b0110 : node38461;
																assign node38461 = (inp[9]) ? 4'b0010 : 4'b0110;
															assign node38465 = (inp[9]) ? node38467 : 4'b0010;
																assign node38467 = (inp[4]) ? 4'b0110 : 4'b0010;
														assign node38470 = (inp[9]) ? node38474 : node38471;
															assign node38471 = (inp[4]) ? 4'b0011 : 4'b0111;
															assign node38474 = (inp[4]) ? 4'b0111 : 4'b0011;
													assign node38477 = (inp[8]) ? node38485 : node38478;
														assign node38478 = (inp[2]) ? node38480 : 4'b0011;
															assign node38480 = (inp[9]) ? node38482 : 4'b0011;
																assign node38482 = (inp[4]) ? 4'b0111 : 4'b0011;
														assign node38485 = (inp[2]) ? 4'b0010 : node38486;
															assign node38486 = (inp[9]) ? node38490 : node38487;
																assign node38487 = (inp[4]) ? 4'b0010 : 4'b0110;
																assign node38490 = (inp[4]) ? 4'b0110 : 4'b0010;
												assign node38494 = (inp[8]) ? node38506 : node38495;
													assign node38495 = (inp[7]) ? node38501 : node38496;
														assign node38496 = (inp[4]) ? node38498 : 4'b0110;
															assign node38498 = (inp[9]) ? 4'b0010 : 4'b0110;
														assign node38501 = (inp[9]) ? node38503 : 4'b0011;
															assign node38503 = (inp[4]) ? 4'b0011 : 4'b0111;
													assign node38506 = (inp[7]) ? node38516 : node38507;
														assign node38507 = (inp[2]) ? 4'b0111 : node38508;
															assign node38508 = (inp[4]) ? node38512 : node38509;
																assign node38509 = (inp[9]) ? 4'b0111 : 4'b0011;
																assign node38512 = (inp[9]) ? 4'b0011 : 4'b0111;
														assign node38516 = (inp[4]) ? 4'b0110 : node38517;
															assign node38517 = (inp[9]) ? 4'b0110 : 4'b0010;
											assign node38521 = (inp[12]) ? node38553 : node38522;
												assign node38522 = (inp[4]) ? node38542 : node38523;
													assign node38523 = (inp[9]) ? node38535 : node38524;
														assign node38524 = (inp[2]) ? node38530 : node38525;
															assign node38525 = (inp[8]) ? node38527 : 4'b0110;
																assign node38527 = (inp[7]) ? 4'b0110 : 4'b0111;
															assign node38530 = (inp[7]) ? 4'b0111 : node38531;
																assign node38531 = (inp[8]) ? 4'b0111 : 4'b0110;
														assign node38535 = (inp[2]) ? 4'b0011 : node38536;
															assign node38536 = (inp[7]) ? node38538 : 4'b0010;
																assign node38538 = (inp[8]) ? 4'b0010 : 4'b0011;
													assign node38542 = (inp[9]) ? node38548 : node38543;
														assign node38543 = (inp[7]) ? 4'b0011 : node38544;
															assign node38544 = (inp[8]) ? 4'b0011 : 4'b0010;
														assign node38548 = (inp[7]) ? 4'b0101 : node38549;
															assign node38549 = (inp[8]) ? 4'b0101 : 4'b0100;
												assign node38553 = (inp[9]) ? node38567 : node38554;
													assign node38554 = (inp[4]) ? node38560 : node38555;
														assign node38555 = (inp[8]) ? 4'b0011 : node38556;
															assign node38556 = (inp[7]) ? 4'b0011 : 4'b0010;
														assign node38560 = (inp[2]) ? 4'b0101 : node38561;
															assign node38561 = (inp[8]) ? node38563 : 4'b0100;
																assign node38563 = (inp[7]) ? 4'b0100 : 4'b0101;
													assign node38567 = (inp[4]) ? node38579 : node38568;
														assign node38568 = (inp[2]) ? node38574 : node38569;
															assign node38569 = (inp[7]) ? node38571 : 4'b0101;
																assign node38571 = (inp[8]) ? 4'b0100 : 4'b0101;
															assign node38574 = (inp[7]) ? node38576 : 4'b0100;
																assign node38576 = (inp[8]) ? 4'b0100 : 4'b0101;
														assign node38579 = (inp[2]) ? node38581 : 4'b0001;
															assign node38581 = (inp[7]) ? node38585 : node38582;
																assign node38582 = (inp[8]) ? 4'b0001 : 4'b0000;
																assign node38585 = (inp[8]) ? 4'b0000 : 4'b0001;
										assign node38588 = (inp[3]) ? node38662 : node38589;
											assign node38589 = (inp[2]) ? node38627 : node38590;
												assign node38590 = (inp[9]) ? node38612 : node38591;
													assign node38591 = (inp[7]) ? node38603 : node38592;
														assign node38592 = (inp[8]) ? node38598 : node38593;
															assign node38593 = (inp[12]) ? 4'b0100 : node38594;
																assign node38594 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node38598 = (inp[4]) ? node38600 : 4'b0101;
																assign node38600 = (inp[12]) ? 4'b0101 : 4'b0001;
														assign node38603 = (inp[8]) ? node38605 : 4'b0101;
															assign node38605 = (inp[4]) ? node38609 : node38606;
																assign node38606 = (inp[12]) ? 4'b0000 : 4'b0100;
																assign node38609 = (inp[12]) ? 4'b0100 : 4'b0000;
													assign node38612 = (inp[7]) ? node38618 : node38613;
														assign node38613 = (inp[8]) ? 4'b0101 : node38614;
															assign node38614 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node38618 = (inp[8]) ? 4'b0000 : node38619;
															assign node38619 = (inp[12]) ? node38623 : node38620;
																assign node38620 = (inp[4]) ? 4'b0101 : 4'b0001;
																assign node38623 = (inp[4]) ? 4'b0001 : 4'b0101;
												assign node38627 = (inp[12]) ? node38641 : node38628;
													assign node38628 = (inp[9]) ? node38638 : node38629;
														assign node38629 = (inp[4]) ? node38633 : node38630;
															assign node38630 = (inp[8]) ? 4'b0101 : 4'b0100;
															assign node38633 = (inp[7]) ? node38635 : 4'b0001;
																assign node38635 = (inp[8]) ? 4'b0000 : 4'b0001;
														assign node38638 = (inp[4]) ? 4'b0101 : 4'b0001;
													assign node38641 = (inp[8]) ? node38649 : node38642;
														assign node38642 = (inp[7]) ? 4'b0001 : node38643;
															assign node38643 = (inp[4]) ? 4'b0000 : node38644;
																assign node38644 = (inp[9]) ? 4'b0100 : 4'b0000;
														assign node38649 = (inp[7]) ? node38655 : node38650;
															assign node38650 = (inp[9]) ? node38652 : 4'b0001;
																assign node38652 = (inp[4]) ? 4'b0001 : 4'b0101;
															assign node38655 = (inp[9]) ? node38659 : node38656;
																assign node38656 = (inp[4]) ? 4'b0100 : 4'b0000;
																assign node38659 = (inp[4]) ? 4'b0000 : 4'b0100;
											assign node38662 = (inp[4]) ? node38696 : node38663;
												assign node38663 = (inp[9]) ? node38685 : node38664;
													assign node38664 = (inp[12]) ? node38672 : node38665;
														assign node38665 = (inp[7]) ? node38669 : node38666;
															assign node38666 = (inp[8]) ? 4'b0101 : 4'b0100;
															assign node38669 = (inp[8]) ? 4'b0100 : 4'b0101;
														assign node38672 = (inp[2]) ? node38680 : node38673;
															assign node38673 = (inp[8]) ? node38677 : node38674;
																assign node38674 = (inp[7]) ? 4'b0001 : 4'b0000;
																assign node38677 = (inp[7]) ? 4'b0000 : 4'b0001;
															assign node38680 = (inp[8]) ? node38682 : 4'b0000;
																assign node38682 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node38685 = (inp[12]) ? node38691 : node38686;
														assign node38686 = (inp[7]) ? 4'b0001 : node38687;
															assign node38687 = (inp[8]) ? 4'b0001 : 4'b0000;
														assign node38691 = (inp[8]) ? node38693 : 4'b0110;
															assign node38693 = (inp[7]) ? 4'b0110 : 4'b0111;
												assign node38696 = (inp[9]) ? node38708 : node38697;
													assign node38697 = (inp[12]) ? node38701 : node38698;
														assign node38698 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node38701 = (inp[2]) ? 4'b0111 : node38702;
															assign node38702 = (inp[8]) ? 4'b0110 : node38703;
																assign node38703 = (inp[7]) ? 4'b0111 : 4'b0110;
													assign node38708 = (inp[12]) ? node38718 : node38709;
														assign node38709 = (inp[2]) ? node38711 : 4'b0110;
															assign node38711 = (inp[8]) ? node38715 : node38712;
																assign node38712 = (inp[7]) ? 4'b0111 : 4'b0110;
																assign node38715 = (inp[7]) ? 4'b0110 : 4'b0111;
														assign node38718 = (inp[7]) ? node38720 : 4'b0011;
															assign node38720 = (inp[8]) ? 4'b0010 : 4'b0011;
									assign node38723 = (inp[15]) ? node38843 : node38724;
										assign node38724 = (inp[3]) ? node38784 : node38725;
											assign node38725 = (inp[7]) ? node38751 : node38726;
												assign node38726 = (inp[8]) ? node38740 : node38727;
													assign node38727 = (inp[4]) ? node38733 : node38728;
														assign node38728 = (inp[12]) ? node38730 : 4'b0100;
															assign node38730 = (inp[9]) ? 4'b0100 : 4'b0000;
														assign node38733 = (inp[12]) ? node38737 : node38734;
															assign node38734 = (inp[9]) ? 4'b0100 : 4'b0000;
															assign node38737 = (inp[9]) ? 4'b0000 : 4'b0100;
													assign node38740 = (inp[12]) ? node38746 : node38741;
														assign node38741 = (inp[2]) ? 4'b0101 : node38742;
															assign node38742 = (inp[9]) ? 4'b0001 : 4'b0101;
														assign node38746 = (inp[9]) ? node38748 : 4'b0001;
															assign node38748 = (inp[4]) ? 4'b0001 : 4'b0101;
												assign node38751 = (inp[8]) ? node38773 : node38752;
													assign node38752 = (inp[9]) ? node38764 : node38753;
														assign node38753 = (inp[2]) ? node38759 : node38754;
															assign node38754 = (inp[12]) ? node38756 : 4'b0001;
																assign node38756 = (inp[4]) ? 4'b0101 : 4'b0001;
															assign node38759 = (inp[12]) ? node38761 : 4'b0101;
																assign node38761 = (inp[4]) ? 4'b0101 : 4'b0001;
														assign node38764 = (inp[2]) ? 4'b0001 : node38765;
															assign node38765 = (inp[12]) ? node38769 : node38766;
																assign node38766 = (inp[4]) ? 4'b0101 : 4'b0001;
																assign node38769 = (inp[4]) ? 4'b0001 : 4'b0101;
													assign node38773 = (inp[9]) ? node38779 : node38774;
														assign node38774 = (inp[12]) ? 4'b0000 : node38775;
															assign node38775 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node38779 = (inp[12]) ? 4'b0100 : node38780;
															assign node38780 = (inp[4]) ? 4'b0100 : 4'b0000;
											assign node38784 = (inp[12]) ? node38816 : node38785;
												assign node38785 = (inp[4]) ? node38797 : node38786;
													assign node38786 = (inp[9]) ? node38792 : node38787;
														assign node38787 = (inp[8]) ? 4'b0100 : node38788;
															assign node38788 = (inp[7]) ? 4'b0101 : 4'b0100;
														assign node38792 = (inp[8]) ? 4'b0000 : node38793;
															assign node38793 = (inp[7]) ? 4'b0001 : 4'b0000;
													assign node38797 = (inp[9]) ? node38811 : node38798;
														assign node38798 = (inp[2]) ? node38806 : node38799;
															assign node38799 = (inp[8]) ? node38803 : node38800;
																assign node38800 = (inp[7]) ? 4'b0001 : 4'b0000;
																assign node38803 = (inp[7]) ? 4'b0000 : 4'b0001;
															assign node38806 = (inp[7]) ? 4'b0001 : node38807;
																assign node38807 = (inp[8]) ? 4'b0001 : 4'b0000;
														assign node38811 = (inp[8]) ? node38813 : 4'b0111;
															assign node38813 = (inp[7]) ? 4'b0110 : 4'b0111;
												assign node38816 = (inp[9]) ? node38828 : node38817;
													assign node38817 = (inp[4]) ? node38821 : node38818;
														assign node38818 = (inp[8]) ? 4'b0001 : 4'b0000;
														assign node38821 = (inp[2]) ? node38823 : 4'b0111;
															assign node38823 = (inp[7]) ? node38825 : 4'b0110;
																assign node38825 = (inp[8]) ? 4'b0110 : 4'b0111;
													assign node38828 = (inp[4]) ? node38838 : node38829;
														assign node38829 = (inp[2]) ? 4'b0110 : node38830;
															assign node38830 = (inp[8]) ? node38834 : node38831;
																assign node38831 = (inp[7]) ? 4'b0111 : 4'b0110;
																assign node38834 = (inp[7]) ? 4'b0110 : 4'b0111;
														assign node38838 = (inp[8]) ? node38840 : 4'b0010;
															assign node38840 = (inp[7]) ? 4'b0010 : 4'b0011;
										assign node38843 = (inp[3]) ? node38901 : node38844;
											assign node38844 = (inp[4]) ? node38870 : node38845;
												assign node38845 = (inp[12]) ? node38855 : node38846;
													assign node38846 = (inp[9]) ? node38850 : node38847;
														assign node38847 = (inp[7]) ? 4'b0110 : 4'b0111;
														assign node38850 = (inp[7]) ? node38852 : 4'b0010;
															assign node38852 = (inp[8]) ? 4'b0010 : 4'b0011;
													assign node38855 = (inp[9]) ? node38867 : node38856;
														assign node38856 = (inp[2]) ? node38862 : node38857;
															assign node38857 = (inp[7]) ? node38859 : 4'b0011;
																assign node38859 = (inp[8]) ? 4'b0010 : 4'b0011;
															assign node38862 = (inp[7]) ? 4'b0010 : node38863;
																assign node38863 = (inp[8]) ? 4'b0011 : 4'b0010;
														assign node38867 = (inp[7]) ? 4'b0111 : 4'b0110;
												assign node38870 = (inp[7]) ? node38892 : node38871;
													assign node38871 = (inp[8]) ? node38885 : node38872;
														assign node38872 = (inp[2]) ? node38880 : node38873;
															assign node38873 = (inp[12]) ? node38877 : node38874;
																assign node38874 = (inp[9]) ? 4'b0110 : 4'b0010;
																assign node38877 = (inp[9]) ? 4'b0010 : 4'b0110;
															assign node38880 = (inp[9]) ? 4'b0010 : node38881;
																assign node38881 = (inp[12]) ? 4'b0110 : 4'b0010;
														assign node38885 = (inp[9]) ? node38889 : node38886;
															assign node38886 = (inp[12]) ? 4'b0111 : 4'b0011;
															assign node38889 = (inp[12]) ? 4'b0011 : 4'b0111;
													assign node38892 = (inp[8]) ? node38898 : node38893;
														assign node38893 = (inp[9]) ? node38895 : 4'b0111;
															assign node38895 = (inp[12]) ? 4'b0011 : 4'b0111;
														assign node38898 = (inp[2]) ? 4'b0110 : 4'b0010;
											assign node38901 = (inp[4]) ? node38943 : node38902;
												assign node38902 = (inp[12]) ? node38928 : node38903;
													assign node38903 = (inp[9]) ? node38917 : node38904;
														assign node38904 = (inp[2]) ? node38910 : node38905;
															assign node38905 = (inp[7]) ? node38907 : 4'b0111;
																assign node38907 = (inp[8]) ? 4'b0110 : 4'b0111;
															assign node38910 = (inp[7]) ? node38914 : node38911;
																assign node38911 = (inp[8]) ? 4'b0111 : 4'b0110;
																assign node38914 = (inp[8]) ? 4'b0110 : 4'b0111;
														assign node38917 = (inp[2]) ? node38923 : node38918;
															assign node38918 = (inp[8]) ? node38920 : 4'b0011;
																assign node38920 = (inp[7]) ? 4'b0010 : 4'b0011;
															assign node38923 = (inp[8]) ? node38925 : 4'b0010;
																assign node38925 = (inp[7]) ? 4'b0010 : 4'b0011;
													assign node38928 = (inp[9]) ? node38938 : node38929;
														assign node38929 = (inp[2]) ? 4'b0011 : node38930;
															assign node38930 = (inp[8]) ? node38934 : node38931;
																assign node38931 = (inp[7]) ? 4'b0011 : 4'b0010;
																assign node38934 = (inp[7]) ? 4'b0010 : 4'b0011;
														assign node38938 = (inp[8]) ? node38940 : 4'b0101;
															assign node38940 = (inp[7]) ? 4'b0100 : 4'b0101;
												assign node38943 = (inp[9]) ? node38955 : node38944;
													assign node38944 = (inp[12]) ? node38950 : node38945;
														assign node38945 = (inp[8]) ? node38947 : 4'b0011;
															assign node38947 = (inp[7]) ? 4'b0010 : 4'b0011;
														assign node38950 = (inp[2]) ? 4'b0100 : node38951;
															assign node38951 = (inp[7]) ? 4'b0101 : 4'b0100;
													assign node38955 = (inp[12]) ? node38963 : node38956;
														assign node38956 = (inp[8]) ? node38960 : node38957;
															assign node38957 = (inp[7]) ? 4'b0101 : 4'b0100;
															assign node38960 = (inp[7]) ? 4'b0100 : 4'b0101;
														assign node38963 = (inp[2]) ? node38971 : node38964;
															assign node38964 = (inp[7]) ? node38968 : node38965;
																assign node38965 = (inp[8]) ? 4'b0001 : 4'b0000;
																assign node38968 = (inp[8]) ? 4'b0000 : 4'b0001;
															assign node38971 = (inp[7]) ? node38973 : 4'b0001;
																assign node38973 = (inp[8]) ? 4'b0000 : 4'b0001;
							assign node38976 = (inp[2]) ? node39596 : node38977;
								assign node38977 = (inp[0]) ? node39279 : node38978;
									assign node38978 = (inp[15]) ? node39136 : node38979;
										assign node38979 = (inp[3]) ? node39043 : node38980;
											assign node38980 = (inp[12]) ? node39008 : node38981;
												assign node38981 = (inp[4]) ? node38999 : node38982;
													assign node38982 = (inp[9]) ? node38992 : node38983;
														assign node38983 = (inp[8]) ? 4'b0110 : node38984;
															assign node38984 = (inp[14]) ? node38988 : node38985;
																assign node38985 = (inp[7]) ? 4'b0110 : 4'b0111;
																assign node38988 = (inp[7]) ? 4'b0111 : 4'b0110;
														assign node38992 = (inp[14]) ? 4'b0010 : node38993;
															assign node38993 = (inp[7]) ? node38995 : 4'b0011;
																assign node38995 = (inp[8]) ? 4'b0011 : 4'b0010;
													assign node38999 = (inp[9]) ? node39001 : 4'b0011;
														assign node39001 = (inp[8]) ? node39003 : 4'b0100;
															assign node39003 = (inp[14]) ? node39005 : 4'b0101;
																assign node39005 = (inp[7]) ? 4'b0100 : 4'b0101;
												assign node39008 = (inp[4]) ? node39028 : node39009;
													assign node39009 = (inp[9]) ? node39015 : node39010;
														assign node39010 = (inp[7]) ? 4'b0011 : node39011;
															assign node39011 = (inp[8]) ? 4'b0011 : 4'b0010;
														assign node39015 = (inp[7]) ? node39023 : node39016;
															assign node39016 = (inp[8]) ? node39020 : node39017;
																assign node39017 = (inp[14]) ? 4'b0100 : 4'b0101;
																assign node39020 = (inp[14]) ? 4'b0101 : 4'b0100;
															assign node39023 = (inp[14]) ? node39025 : 4'b0100;
																assign node39025 = (inp[8]) ? 4'b0100 : 4'b0101;
													assign node39028 = (inp[9]) ? node39034 : node39029;
														assign node39029 = (inp[8]) ? node39031 : 4'b0100;
															assign node39031 = (inp[7]) ? 4'b0101 : 4'b0100;
														assign node39034 = (inp[14]) ? 4'b0001 : node39035;
															assign node39035 = (inp[8]) ? node39039 : node39036;
																assign node39036 = (inp[7]) ? 4'b0000 : 4'b0001;
																assign node39039 = (inp[7]) ? 4'b0001 : 4'b0000;
											assign node39043 = (inp[7]) ? node39087 : node39044;
												assign node39044 = (inp[9]) ? node39064 : node39045;
													assign node39045 = (inp[8]) ? node39053 : node39046;
														assign node39046 = (inp[14]) ? 4'b0000 : node39047;
															assign node39047 = (inp[4]) ? node39049 : 4'b0001;
																assign node39049 = (inp[12]) ? 4'b0101 : 4'b0001;
														assign node39053 = (inp[14]) ? node39059 : node39054;
															assign node39054 = (inp[4]) ? 4'b0100 : node39055;
																assign node39055 = (inp[12]) ? 4'b0000 : 4'b0100;
															assign node39059 = (inp[4]) ? 4'b0001 : node39060;
																assign node39060 = (inp[12]) ? 4'b0001 : 4'b0101;
													assign node39064 = (inp[14]) ? node39074 : node39065;
														assign node39065 = (inp[8]) ? 4'b0000 : node39066;
															assign node39066 = (inp[4]) ? node39070 : node39067;
																assign node39067 = (inp[12]) ? 4'b0101 : 4'b0001;
																assign node39070 = (inp[12]) ? 4'b0001 : 4'b0101;
														assign node39074 = (inp[8]) ? node39082 : node39075;
															assign node39075 = (inp[12]) ? node39079 : node39076;
																assign node39076 = (inp[4]) ? 4'b0100 : 4'b0000;
																assign node39079 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node39082 = (inp[12]) ? node39084 : 4'b0101;
																assign node39084 = (inp[4]) ? 4'b0001 : 4'b0101;
												assign node39087 = (inp[8]) ? node39111 : node39088;
													assign node39088 = (inp[14]) ? node39104 : node39089;
														assign node39089 = (inp[4]) ? node39097 : node39090;
															assign node39090 = (inp[9]) ? node39094 : node39091;
																assign node39091 = (inp[12]) ? 4'b0000 : 4'b0100;
																assign node39094 = (inp[12]) ? 4'b0100 : 4'b0000;
															assign node39097 = (inp[12]) ? node39101 : node39098;
																assign node39098 = (inp[9]) ? 4'b0100 : 4'b0000;
																assign node39101 = (inp[9]) ? 4'b0000 : 4'b0100;
														assign node39104 = (inp[12]) ? node39106 : 4'b0101;
															assign node39106 = (inp[9]) ? 4'b0001 : node39107;
																assign node39107 = (inp[4]) ? 4'b0101 : 4'b0001;
													assign node39111 = (inp[14]) ? node39127 : node39112;
														assign node39112 = (inp[9]) ? node39120 : node39113;
															assign node39113 = (inp[4]) ? node39117 : node39114;
																assign node39114 = (inp[12]) ? 4'b0001 : 4'b0101;
																assign node39117 = (inp[12]) ? 4'b0101 : 4'b0001;
															assign node39120 = (inp[12]) ? node39124 : node39121;
																assign node39121 = (inp[4]) ? 4'b0101 : 4'b0001;
																assign node39124 = (inp[4]) ? 4'b0001 : 4'b0101;
														assign node39127 = (inp[9]) ? node39129 : 4'b0100;
															assign node39129 = (inp[12]) ? node39133 : node39130;
																assign node39130 = (inp[4]) ? 4'b0100 : 4'b0000;
																assign node39133 = (inp[4]) ? 4'b0000 : 4'b0100;
										assign node39136 = (inp[3]) ? node39206 : node39137;
											assign node39137 = (inp[4]) ? node39175 : node39138;
												assign node39138 = (inp[9]) ? node39160 : node39139;
													assign node39139 = (inp[12]) ? node39147 : node39140;
														assign node39140 = (inp[7]) ? node39142 : 4'b0101;
															assign node39142 = (inp[8]) ? node39144 : 4'b0100;
																assign node39144 = (inp[14]) ? 4'b0100 : 4'b0101;
														assign node39147 = (inp[8]) ? node39155 : node39148;
															assign node39148 = (inp[14]) ? node39152 : node39149;
																assign node39149 = (inp[7]) ? 4'b0000 : 4'b0001;
																assign node39152 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node39155 = (inp[14]) ? node39157 : 4'b0000;
																assign node39157 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node39160 = (inp[12]) ? node39168 : node39161;
														assign node39161 = (inp[14]) ? node39163 : 4'b0001;
															assign node39163 = (inp[8]) ? node39165 : 4'b0000;
																assign node39165 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node39168 = (inp[7]) ? 4'b0111 : node39169;
															assign node39169 = (inp[8]) ? 4'b0110 : node39170;
																assign node39170 = (inp[14]) ? 4'b0110 : 4'b0111;
												assign node39175 = (inp[9]) ? node39189 : node39176;
													assign node39176 = (inp[12]) ? node39184 : node39177;
														assign node39177 = (inp[14]) ? 4'b0000 : node39178;
															assign node39178 = (inp[7]) ? node39180 : 4'b0000;
																assign node39180 = (inp[8]) ? 4'b0001 : 4'b0000;
														assign node39184 = (inp[14]) ? 4'b0110 : node39185;
															assign node39185 = (inp[7]) ? 4'b0111 : 4'b0110;
													assign node39189 = (inp[12]) ? node39197 : node39190;
														assign node39190 = (inp[8]) ? node39192 : 4'b0111;
															assign node39192 = (inp[7]) ? 4'b0110 : node39193;
																assign node39193 = (inp[14]) ? 4'b0111 : 4'b0110;
														assign node39197 = (inp[14]) ? 4'b0010 : node39198;
															assign node39198 = (inp[8]) ? node39202 : node39199;
																assign node39199 = (inp[7]) ? 4'b0010 : 4'b0011;
																assign node39202 = (inp[7]) ? 4'b0011 : 4'b0010;
											assign node39206 = (inp[12]) ? node39236 : node39207;
												assign node39207 = (inp[4]) ? node39219 : node39208;
													assign node39208 = (inp[9]) ? node39214 : node39209;
														assign node39209 = (inp[14]) ? 4'b0111 : node39210;
															assign node39210 = (inp[8]) ? 4'b0110 : 4'b0111;
														assign node39214 = (inp[8]) ? node39216 : 4'b0011;
															assign node39216 = (inp[14]) ? 4'b0011 : 4'b0010;
													assign node39219 = (inp[9]) ? node39221 : 4'b0011;
														assign node39221 = (inp[14]) ? node39229 : node39222;
															assign node39222 = (inp[8]) ? node39226 : node39223;
																assign node39223 = (inp[7]) ? 4'b0110 : 4'b0111;
																assign node39226 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node39229 = (inp[8]) ? node39233 : node39230;
																assign node39230 = (inp[7]) ? 4'b0111 : 4'b0110;
																assign node39233 = (inp[7]) ? 4'b0110 : 4'b0111;
												assign node39236 = (inp[4]) ? node39256 : node39237;
													assign node39237 = (inp[9]) ? node39251 : node39238;
														assign node39238 = (inp[8]) ? node39246 : node39239;
															assign node39239 = (inp[14]) ? node39243 : node39240;
																assign node39240 = (inp[7]) ? 4'b0010 : 4'b0011;
																assign node39243 = (inp[7]) ? 4'b0011 : 4'b0010;
															assign node39246 = (inp[7]) ? node39248 : 4'b0011;
																assign node39248 = (inp[14]) ? 4'b0010 : 4'b0011;
														assign node39251 = (inp[7]) ? node39253 : 4'b0111;
															assign node39253 = (inp[8]) ? 4'b0111 : 4'b0110;
													assign node39256 = (inp[9]) ? node39268 : node39257;
														assign node39257 = (inp[7]) ? node39263 : node39258;
															assign node39258 = (inp[14]) ? 4'b0110 : node39259;
																assign node39259 = (inp[8]) ? 4'b0110 : 4'b0111;
															assign node39263 = (inp[8]) ? node39265 : 4'b0111;
																assign node39265 = (inp[14]) ? 4'b0110 : 4'b0111;
														assign node39268 = (inp[7]) ? node39274 : node39269;
															assign node39269 = (inp[14]) ? 4'b0011 : node39270;
																assign node39270 = (inp[8]) ? 4'b0010 : 4'b0011;
															assign node39274 = (inp[14]) ? node39276 : 4'b0010;
																assign node39276 = (inp[8]) ? 4'b0010 : 4'b0011;
									assign node39279 = (inp[15]) ? node39447 : node39280;
										assign node39280 = (inp[3]) ? node39362 : node39281;
											assign node39281 = (inp[12]) ? node39323 : node39282;
												assign node39282 = (inp[4]) ? node39306 : node39283;
													assign node39283 = (inp[9]) ? node39295 : node39284;
														assign node39284 = (inp[8]) ? node39290 : node39285;
															assign node39285 = (inp[14]) ? node39287 : 4'b0100;
																assign node39287 = (inp[7]) ? 4'b0101 : 4'b0100;
															assign node39290 = (inp[7]) ? 4'b0101 : node39291;
																assign node39291 = (inp[14]) ? 4'b0101 : 4'b0100;
														assign node39295 = (inp[14]) ? node39301 : node39296;
															assign node39296 = (inp[8]) ? node39298 : 4'b0000;
																assign node39298 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node39301 = (inp[8]) ? 4'b0001 : node39302;
																assign node39302 = (inp[7]) ? 4'b0001 : 4'b0000;
													assign node39306 = (inp[9]) ? node39316 : node39307;
														assign node39307 = (inp[7]) ? 4'b0000 : node39308;
															assign node39308 = (inp[14]) ? node39312 : node39309;
																assign node39309 = (inp[8]) ? 4'b0000 : 4'b0001;
																assign node39312 = (inp[8]) ? 4'b0001 : 4'b0000;
														assign node39316 = (inp[7]) ? 4'b0110 : node39317;
															assign node39317 = (inp[8]) ? 4'b0111 : node39318;
																assign node39318 = (inp[14]) ? 4'b0110 : 4'b0111;
												assign node39323 = (inp[4]) ? node39343 : node39324;
													assign node39324 = (inp[9]) ? node39336 : node39325;
														assign node39325 = (inp[8]) ? node39331 : node39326;
															assign node39326 = (inp[14]) ? node39328 : 4'b0000;
																assign node39328 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node39331 = (inp[14]) ? 4'b0001 : node39332;
																assign node39332 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node39336 = (inp[14]) ? 4'b0110 : node39337;
															assign node39337 = (inp[7]) ? node39339 : 4'b0110;
																assign node39339 = (inp[8]) ? 4'b0111 : 4'b0110;
													assign node39343 = (inp[9]) ? node39355 : node39344;
														assign node39344 = (inp[8]) ? node39350 : node39345;
															assign node39345 = (inp[7]) ? node39347 : 4'b0110;
																assign node39347 = (inp[14]) ? 4'b0111 : 4'b0110;
															assign node39350 = (inp[14]) ? node39352 : 4'b0111;
																assign node39352 = (inp[7]) ? 4'b0110 : 4'b0111;
														assign node39355 = (inp[8]) ? 4'b0011 : node39356;
															assign node39356 = (inp[14]) ? 4'b0010 : node39357;
																assign node39357 = (inp[7]) ? 4'b0010 : 4'b0011;
											assign node39362 = (inp[9]) ? node39406 : node39363;
												assign node39363 = (inp[7]) ? node39387 : node39364;
													assign node39364 = (inp[4]) ? node39376 : node39365;
														assign node39365 = (inp[12]) ? node39369 : node39366;
															assign node39366 = (inp[8]) ? 4'b0110 : 4'b0111;
															assign node39369 = (inp[8]) ? node39373 : node39370;
																assign node39370 = (inp[14]) ? 4'b0010 : 4'b0011;
																assign node39373 = (inp[14]) ? 4'b0011 : 4'b0010;
														assign node39376 = (inp[12]) ? node39382 : node39377;
															assign node39377 = (inp[8]) ? 4'b0010 : node39378;
																assign node39378 = (inp[14]) ? 4'b0010 : 4'b0011;
															assign node39382 = (inp[8]) ? node39384 : 4'b0110;
																assign node39384 = (inp[14]) ? 4'b0111 : 4'b0110;
													assign node39387 = (inp[14]) ? node39397 : node39388;
														assign node39388 = (inp[8]) ? node39394 : node39389;
															assign node39389 = (inp[12]) ? 4'b0110 : node39390;
																assign node39390 = (inp[4]) ? 4'b0010 : 4'b0110;
															assign node39394 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node39397 = (inp[8]) ? 4'b0110 : node39398;
															assign node39398 = (inp[12]) ? node39402 : node39399;
																assign node39399 = (inp[4]) ? 4'b0011 : 4'b0111;
																assign node39402 = (inp[4]) ? 4'b0111 : 4'b0011;
												assign node39406 = (inp[12]) ? node39428 : node39407;
													assign node39407 = (inp[4]) ? node39415 : node39408;
														assign node39408 = (inp[14]) ? 4'b0010 : node39409;
															assign node39409 = (inp[7]) ? 4'b0010 : node39410;
																assign node39410 = (inp[8]) ? 4'b0010 : 4'b0011;
														assign node39415 = (inp[8]) ? node39423 : node39416;
															assign node39416 = (inp[14]) ? node39420 : node39417;
																assign node39417 = (inp[7]) ? 4'b0110 : 4'b0111;
																assign node39420 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node39423 = (inp[7]) ? node39425 : 4'b0110;
																assign node39425 = (inp[14]) ? 4'b0110 : 4'b0111;
													assign node39428 = (inp[4]) ? node39442 : node39429;
														assign node39429 = (inp[7]) ? node39435 : node39430;
															assign node39430 = (inp[14]) ? node39432 : 4'b0111;
																assign node39432 = (inp[8]) ? 4'b0111 : 4'b0110;
															assign node39435 = (inp[8]) ? node39439 : node39436;
																assign node39436 = (inp[14]) ? 4'b0111 : 4'b0110;
																assign node39439 = (inp[14]) ? 4'b0110 : 4'b0111;
														assign node39442 = (inp[8]) ? node39444 : 4'b0011;
															assign node39444 = (inp[14]) ? 4'b0010 : 4'b0011;
										assign node39447 = (inp[3]) ? node39523 : node39448;
											assign node39448 = (inp[12]) ? node39486 : node39449;
												assign node39449 = (inp[4]) ? node39469 : node39450;
													assign node39450 = (inp[9]) ? node39458 : node39451;
														assign node39451 = (inp[8]) ? node39453 : 4'b0110;
															assign node39453 = (inp[7]) ? 4'b0110 : node39454;
																assign node39454 = (inp[14]) ? 4'b0111 : 4'b0110;
														assign node39458 = (inp[14]) ? node39464 : node39459;
															assign node39459 = (inp[7]) ? 4'b0010 : node39460;
																assign node39460 = (inp[8]) ? 4'b0010 : 4'b0011;
															assign node39464 = (inp[7]) ? 4'b0011 : node39465;
																assign node39465 = (inp[8]) ? 4'b0011 : 4'b0010;
													assign node39469 = (inp[9]) ? node39479 : node39470;
														assign node39470 = (inp[14]) ? 4'b0011 : node39471;
															assign node39471 = (inp[8]) ? node39475 : node39472;
																assign node39472 = (inp[7]) ? 4'b0010 : 4'b0011;
																assign node39475 = (inp[7]) ? 4'b0011 : 4'b0010;
														assign node39479 = (inp[8]) ? 4'b0100 : node39480;
															assign node39480 = (inp[7]) ? 4'b0101 : node39481;
																assign node39481 = (inp[14]) ? 4'b0100 : 4'b0101;
												assign node39486 = (inp[9]) ? node39506 : node39487;
													assign node39487 = (inp[4]) ? node39495 : node39488;
														assign node39488 = (inp[7]) ? node39490 : 4'b0010;
															assign node39490 = (inp[8]) ? node39492 : 4'b0011;
																assign node39492 = (inp[14]) ? 4'b0010 : 4'b0011;
														assign node39495 = (inp[14]) ? node39501 : node39496;
															assign node39496 = (inp[8]) ? 4'b0100 : node39497;
																assign node39497 = (inp[7]) ? 4'b0100 : 4'b0101;
															assign node39501 = (inp[8]) ? 4'b0101 : node39502;
																assign node39502 = (inp[7]) ? 4'b0101 : 4'b0100;
													assign node39506 = (inp[4]) ? node39520 : node39507;
														assign node39507 = (inp[7]) ? node39513 : node39508;
															assign node39508 = (inp[8]) ? node39510 : 4'b0101;
																assign node39510 = (inp[14]) ? 4'b0101 : 4'b0100;
															assign node39513 = (inp[8]) ? node39517 : node39514;
																assign node39514 = (inp[14]) ? 4'b0101 : 4'b0100;
																assign node39517 = (inp[14]) ? 4'b0100 : 4'b0101;
														assign node39520 = (inp[14]) ? 4'b0000 : 4'b0001;
											assign node39523 = (inp[9]) ? node39559 : node39524;
												assign node39524 = (inp[12]) ? node39542 : node39525;
													assign node39525 = (inp[4]) ? node39535 : node39526;
														assign node39526 = (inp[7]) ? 4'b0101 : node39527;
															assign node39527 = (inp[8]) ? node39531 : node39528;
																assign node39528 = (inp[14]) ? 4'b0100 : 4'b0101;
																assign node39531 = (inp[14]) ? 4'b0101 : 4'b0100;
														assign node39535 = (inp[14]) ? 4'b0001 : node39536;
															assign node39536 = (inp[8]) ? 4'b0001 : node39537;
																assign node39537 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node39542 = (inp[4]) ? node39546 : node39543;
														assign node39543 = (inp[8]) ? 4'b0001 : 4'b0000;
														assign node39546 = (inp[7]) ? node39552 : node39547;
															assign node39547 = (inp[8]) ? 4'b0100 : node39548;
																assign node39548 = (inp[14]) ? 4'b0100 : 4'b0101;
															assign node39552 = (inp[8]) ? node39556 : node39553;
																assign node39553 = (inp[14]) ? 4'b0101 : 4'b0100;
																assign node39556 = (inp[14]) ? 4'b0100 : 4'b0101;
												assign node39559 = (inp[8]) ? node39573 : node39560;
													assign node39560 = (inp[7]) ? node39568 : node39561;
														assign node39561 = (inp[14]) ? node39563 : 4'b0001;
															assign node39563 = (inp[4]) ? 4'b0000 : node39564;
																assign node39564 = (inp[12]) ? 4'b0100 : 4'b0000;
														assign node39568 = (inp[14]) ? 4'b0001 : node39569;
															assign node39569 = (inp[12]) ? 4'b0000 : 4'b0100;
													assign node39573 = (inp[14]) ? node39583 : node39574;
														assign node39574 = (inp[7]) ? 4'b0101 : node39575;
															assign node39575 = (inp[12]) ? node39579 : node39576;
																assign node39576 = (inp[4]) ? 4'b0100 : 4'b0000;
																assign node39579 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node39583 = (inp[7]) ? node39591 : node39584;
															assign node39584 = (inp[12]) ? node39588 : node39585;
																assign node39585 = (inp[4]) ? 4'b0101 : 4'b0001;
																assign node39588 = (inp[4]) ? 4'b0001 : 4'b0101;
															assign node39591 = (inp[12]) ? node39593 : 4'b0000;
																assign node39593 = (inp[4]) ? 4'b0000 : 4'b0100;
								assign node39596 = (inp[15]) ? node39878 : node39597;
									assign node39597 = (inp[0]) ? node39749 : node39598;
										assign node39598 = (inp[3]) ? node39656 : node39599;
											assign node39599 = (inp[9]) ? node39631 : node39600;
												assign node39600 = (inp[12]) ? node39620 : node39601;
													assign node39601 = (inp[4]) ? node39607 : node39602;
														assign node39602 = (inp[8]) ? 4'b0111 : node39603;
															assign node39603 = (inp[7]) ? 4'b0111 : 4'b0110;
														assign node39607 = (inp[14]) ? node39615 : node39608;
															assign node39608 = (inp[8]) ? node39612 : node39609;
																assign node39609 = (inp[7]) ? 4'b0011 : 4'b0010;
																assign node39612 = (inp[7]) ? 4'b0010 : 4'b0011;
															assign node39615 = (inp[7]) ? 4'b0011 : node39616;
																assign node39616 = (inp[8]) ? 4'b0011 : 4'b0010;
													assign node39620 = (inp[4]) ? node39626 : node39621;
														assign node39621 = (inp[7]) ? 4'b0010 : node39622;
															assign node39622 = (inp[8]) ? 4'b0011 : 4'b0010;
														assign node39626 = (inp[7]) ? node39628 : 4'b0101;
															assign node39628 = (inp[8]) ? 4'b0100 : 4'b0101;
												assign node39631 = (inp[4]) ? node39643 : node39632;
													assign node39632 = (inp[12]) ? node39638 : node39633;
														assign node39633 = (inp[7]) ? 4'b0011 : node39634;
															assign node39634 = (inp[8]) ? 4'b0011 : 4'b0010;
														assign node39638 = (inp[7]) ? 4'b0100 : node39639;
															assign node39639 = (inp[8]) ? 4'b0101 : 4'b0100;
													assign node39643 = (inp[12]) ? node39651 : node39644;
														assign node39644 = (inp[8]) ? node39648 : node39645;
															assign node39645 = (inp[7]) ? 4'b0101 : 4'b0100;
															assign node39648 = (inp[7]) ? 4'b0100 : 4'b0101;
														assign node39651 = (inp[7]) ? node39653 : 4'b0001;
															assign node39653 = (inp[8]) ? 4'b0000 : 4'b0001;
											assign node39656 = (inp[14]) ? node39706 : node39657;
												assign node39657 = (inp[12]) ? node39679 : node39658;
													assign node39658 = (inp[4]) ? node39666 : node39659;
														assign node39659 = (inp[9]) ? 4'b0000 : node39660;
															assign node39660 = (inp[8]) ? node39662 : 4'b0100;
																assign node39662 = (inp[7]) ? 4'b0100 : 4'b0101;
														assign node39666 = (inp[9]) ? node39674 : node39667;
															assign node39667 = (inp[8]) ? node39671 : node39668;
																assign node39668 = (inp[7]) ? 4'b0001 : 4'b0000;
																assign node39671 = (inp[7]) ? 4'b0000 : 4'b0001;
															assign node39674 = (inp[8]) ? 4'b0100 : node39675;
																assign node39675 = (inp[7]) ? 4'b0101 : 4'b0100;
													assign node39679 = (inp[4]) ? node39693 : node39680;
														assign node39680 = (inp[9]) ? node39688 : node39681;
															assign node39681 = (inp[7]) ? node39685 : node39682;
																assign node39682 = (inp[8]) ? 4'b0001 : 4'b0000;
																assign node39685 = (inp[8]) ? 4'b0000 : 4'b0001;
															assign node39688 = (inp[7]) ? node39690 : 4'b0101;
																assign node39690 = (inp[8]) ? 4'b0100 : 4'b0101;
														assign node39693 = (inp[9]) ? node39699 : node39694;
															assign node39694 = (inp[8]) ? 4'b0101 : node39695;
																assign node39695 = (inp[7]) ? 4'b0101 : 4'b0100;
															assign node39699 = (inp[7]) ? node39703 : node39700;
																assign node39700 = (inp[8]) ? 4'b0001 : 4'b0000;
																assign node39703 = (inp[8]) ? 4'b0000 : 4'b0001;
												assign node39706 = (inp[9]) ? node39722 : node39707;
													assign node39707 = (inp[4]) ? node39715 : node39708;
														assign node39708 = (inp[12]) ? 4'b0000 : node39709;
															assign node39709 = (inp[8]) ? node39711 : 4'b0101;
																assign node39711 = (inp[7]) ? 4'b0100 : 4'b0101;
														assign node39715 = (inp[12]) ? node39717 : 4'b0001;
															assign node39717 = (inp[8]) ? node39719 : 4'b0101;
																assign node39719 = (inp[7]) ? 4'b0100 : 4'b0101;
													assign node39722 = (inp[12]) ? node39736 : node39723;
														assign node39723 = (inp[4]) ? node39731 : node39724;
															assign node39724 = (inp[7]) ? node39728 : node39725;
																assign node39725 = (inp[8]) ? 4'b0001 : 4'b0000;
																assign node39728 = (inp[8]) ? 4'b0000 : 4'b0001;
															assign node39731 = (inp[7]) ? node39733 : 4'b0101;
																assign node39733 = (inp[8]) ? 4'b0100 : 4'b0101;
														assign node39736 = (inp[4]) ? node39742 : node39737;
															assign node39737 = (inp[8]) ? 4'b0101 : node39738;
																assign node39738 = (inp[7]) ? 4'b0101 : 4'b0100;
															assign node39742 = (inp[8]) ? node39746 : node39743;
																assign node39743 = (inp[7]) ? 4'b0001 : 4'b0000;
																assign node39746 = (inp[7]) ? 4'b0000 : 4'b0001;
										assign node39749 = (inp[3]) ? node39805 : node39750;
											assign node39750 = (inp[9]) ? node39772 : node39751;
												assign node39751 = (inp[12]) ? node39761 : node39752;
													assign node39752 = (inp[4]) ? node39754 : 4'b0101;
														assign node39754 = (inp[8]) ? node39758 : node39755;
															assign node39755 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node39758 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node39761 = (inp[4]) ? node39767 : node39762;
														assign node39762 = (inp[14]) ? 4'b0000 : node39763;
															assign node39763 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node39767 = (inp[14]) ? node39769 : 4'b0110;
															assign node39769 = (inp[7]) ? 4'b0110 : 4'b0111;
												assign node39772 = (inp[12]) ? node39788 : node39773;
													assign node39773 = (inp[4]) ? node39781 : node39774;
														assign node39774 = (inp[14]) ? 4'b0001 : node39775;
															assign node39775 = (inp[8]) ? node39777 : 4'b0000;
																assign node39777 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node39781 = (inp[14]) ? 4'b0110 : node39782;
															assign node39782 = (inp[8]) ? 4'b0111 : node39783;
																assign node39783 = (inp[7]) ? 4'b0111 : 4'b0110;
													assign node39788 = (inp[4]) ? node39796 : node39789;
														assign node39789 = (inp[8]) ? node39793 : node39790;
															assign node39790 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node39793 = (inp[7]) ? 4'b0110 : 4'b0111;
														assign node39796 = (inp[14]) ? 4'b0010 : node39797;
															assign node39797 = (inp[8]) ? node39801 : node39798;
																assign node39798 = (inp[7]) ? 4'b0011 : 4'b0010;
																assign node39801 = (inp[7]) ? 4'b0010 : 4'b0011;
											assign node39805 = (inp[14]) ? node39841 : node39806;
												assign node39806 = (inp[9]) ? node39818 : node39807;
													assign node39807 = (inp[12]) ? node39811 : node39808;
														assign node39808 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node39811 = (inp[4]) ? node39813 : 4'b0011;
															assign node39813 = (inp[7]) ? node39815 : 4'b0111;
																assign node39815 = (inp[8]) ? 4'b0110 : 4'b0111;
													assign node39818 = (inp[4]) ? node39830 : node39819;
														assign node39819 = (inp[12]) ? node39825 : node39820;
															assign node39820 = (inp[7]) ? 4'b0011 : node39821;
																assign node39821 = (inp[8]) ? 4'b0011 : 4'b0010;
															assign node39825 = (inp[7]) ? node39827 : 4'b0111;
																assign node39827 = (inp[8]) ? 4'b0110 : 4'b0111;
														assign node39830 = (inp[12]) ? node39836 : node39831;
															assign node39831 = (inp[8]) ? 4'b0111 : node39832;
																assign node39832 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node39836 = (inp[7]) ? node39838 : 4'b0011;
																assign node39838 = (inp[8]) ? 4'b0010 : 4'b0011;
												assign node39841 = (inp[7]) ? node39865 : node39842;
													assign node39842 = (inp[8]) ? node39854 : node39843;
														assign node39843 = (inp[9]) ? node39849 : node39844;
															assign node39844 = (inp[12]) ? node39846 : 4'b0110;
																assign node39846 = (inp[4]) ? 4'b0110 : 4'b0010;
															assign node39849 = (inp[4]) ? node39851 : 4'b0010;
																assign node39851 = (inp[12]) ? 4'b0010 : 4'b0110;
														assign node39854 = (inp[4]) ? node39860 : node39855;
															assign node39855 = (inp[12]) ? node39857 : 4'b0111;
																assign node39857 = (inp[9]) ? 4'b0111 : 4'b0011;
															assign node39860 = (inp[12]) ? 4'b0011 : node39861;
																assign node39861 = (inp[9]) ? 4'b0111 : 4'b0011;
													assign node39865 = (inp[8]) ? node39875 : node39866;
														assign node39866 = (inp[9]) ? node39868 : 4'b0011;
															assign node39868 = (inp[12]) ? node39872 : node39869;
																assign node39869 = (inp[4]) ? 4'b0111 : 4'b0011;
																assign node39872 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node39875 = (inp[9]) ? 4'b0010 : 4'b0110;
									assign node39878 = (inp[0]) ? node40012 : node39879;
										assign node39879 = (inp[3]) ? node39947 : node39880;
											assign node39880 = (inp[4]) ? node39914 : node39881;
												assign node39881 = (inp[9]) ? node39903 : node39882;
													assign node39882 = (inp[12]) ? node39892 : node39883;
														assign node39883 = (inp[14]) ? node39885 : 4'b0101;
															assign node39885 = (inp[7]) ? node39889 : node39886;
																assign node39886 = (inp[8]) ? 4'b0101 : 4'b0100;
																assign node39889 = (inp[8]) ? 4'b0100 : 4'b0101;
														assign node39892 = (inp[14]) ? node39898 : node39893;
															assign node39893 = (inp[7]) ? 4'b0001 : node39894;
																assign node39894 = (inp[8]) ? 4'b0001 : 4'b0000;
															assign node39898 = (inp[8]) ? node39900 : 4'b0001;
																assign node39900 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node39903 = (inp[12]) ? node39909 : node39904;
														assign node39904 = (inp[7]) ? 4'b0001 : node39905;
															assign node39905 = (inp[8]) ? 4'b0001 : 4'b0000;
														assign node39909 = (inp[14]) ? node39911 : 4'b0110;
															assign node39911 = (inp[7]) ? 4'b0110 : 4'b0111;
												assign node39914 = (inp[9]) ? node39932 : node39915;
													assign node39915 = (inp[12]) ? node39919 : node39916;
														assign node39916 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node39919 = (inp[14]) ? node39927 : node39920;
															assign node39920 = (inp[7]) ? node39924 : node39921;
																assign node39921 = (inp[8]) ? 4'b0111 : 4'b0110;
																assign node39924 = (inp[8]) ? 4'b0110 : 4'b0111;
															assign node39927 = (inp[7]) ? node39929 : 4'b0110;
																assign node39929 = (inp[8]) ? 4'b0110 : 4'b0111;
													assign node39932 = (inp[12]) ? node39940 : node39933;
														assign node39933 = (inp[8]) ? node39937 : node39934;
															assign node39934 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node39937 = (inp[7]) ? 4'b0110 : 4'b0111;
														assign node39940 = (inp[8]) ? node39944 : node39941;
															assign node39941 = (inp[7]) ? 4'b0011 : 4'b0010;
															assign node39944 = (inp[7]) ? 4'b0010 : 4'b0011;
											assign node39947 = (inp[4]) ? node39987 : node39948;
												assign node39948 = (inp[14]) ? node39966 : node39949;
													assign node39949 = (inp[9]) ? node39959 : node39950;
														assign node39950 = (inp[12]) ? node39952 : 4'b0111;
															assign node39952 = (inp[8]) ? node39956 : node39953;
																assign node39953 = (inp[7]) ? 4'b0011 : 4'b0010;
																assign node39956 = (inp[7]) ? 4'b0010 : 4'b0011;
														assign node39959 = (inp[12]) ? 4'b0111 : node39960;
															assign node39960 = (inp[8]) ? node39962 : 4'b0011;
																assign node39962 = (inp[7]) ? 4'b0010 : 4'b0011;
													assign node39966 = (inp[8]) ? node39976 : node39967;
														assign node39967 = (inp[7]) ? 4'b0011 : node39968;
															assign node39968 = (inp[9]) ? node39972 : node39969;
																assign node39969 = (inp[12]) ? 4'b0010 : 4'b0110;
																assign node39972 = (inp[12]) ? 4'b0110 : 4'b0010;
														assign node39976 = (inp[7]) ? node39982 : node39977;
															assign node39977 = (inp[9]) ? 4'b0111 : node39978;
																assign node39978 = (inp[12]) ? 4'b0011 : 4'b0111;
															assign node39982 = (inp[12]) ? 4'b0110 : node39983;
																assign node39983 = (inp[9]) ? 4'b0010 : 4'b0110;
												assign node39987 = (inp[7]) ? node40001 : node39988;
													assign node39988 = (inp[8]) ? node39994 : node39989;
														assign node39989 = (inp[9]) ? node39991 : 4'b0110;
															assign node39991 = (inp[12]) ? 4'b0010 : 4'b0110;
														assign node39994 = (inp[12]) ? node39998 : node39995;
															assign node39995 = (inp[9]) ? 4'b0111 : 4'b0011;
															assign node39998 = (inp[9]) ? 4'b0011 : 4'b0111;
													assign node40001 = (inp[8]) ? node40005 : node40002;
														assign node40002 = (inp[9]) ? 4'b0011 : 4'b0111;
														assign node40005 = (inp[9]) ? node40009 : node40006;
															assign node40006 = (inp[12]) ? 4'b0110 : 4'b0010;
															assign node40009 = (inp[12]) ? 4'b0010 : 4'b0110;
										assign node40012 = (inp[3]) ? node40074 : node40013;
											assign node40013 = (inp[4]) ? node40045 : node40014;
												assign node40014 = (inp[12]) ? node40030 : node40015;
													assign node40015 = (inp[9]) ? node40023 : node40016;
														assign node40016 = (inp[7]) ? node40020 : node40017;
															assign node40017 = (inp[8]) ? 4'b0111 : 4'b0110;
															assign node40020 = (inp[8]) ? 4'b0110 : 4'b0111;
														assign node40023 = (inp[8]) ? node40027 : node40024;
															assign node40024 = (inp[7]) ? 4'b0011 : 4'b0010;
															assign node40027 = (inp[7]) ? 4'b0010 : 4'b0011;
													assign node40030 = (inp[9]) ? 4'b0101 : node40031;
														assign node40031 = (inp[14]) ? node40037 : node40032;
															assign node40032 = (inp[8]) ? 4'b0011 : node40033;
																assign node40033 = (inp[7]) ? 4'b0011 : 4'b0010;
															assign node40037 = (inp[7]) ? node40041 : node40038;
																assign node40038 = (inp[8]) ? 4'b0011 : 4'b0010;
																assign node40041 = (inp[8]) ? 4'b0010 : 4'b0011;
												assign node40045 = (inp[9]) ? node40063 : node40046;
													assign node40046 = (inp[12]) ? node40058 : node40047;
														assign node40047 = (inp[14]) ? node40053 : node40048;
															assign node40048 = (inp[8]) ? 4'b0011 : node40049;
																assign node40049 = (inp[7]) ? 4'b0011 : 4'b0010;
															assign node40053 = (inp[7]) ? 4'b0010 : node40054;
																assign node40054 = (inp[8]) ? 4'b0011 : 4'b0010;
														assign node40058 = (inp[8]) ? node40060 : 4'b0100;
															assign node40060 = (inp[7]) ? 4'b0100 : 4'b0101;
													assign node40063 = (inp[12]) ? node40071 : node40064;
														assign node40064 = (inp[7]) ? node40068 : node40065;
															assign node40065 = (inp[8]) ? 4'b0101 : 4'b0100;
															assign node40068 = (inp[8]) ? 4'b0100 : 4'b0101;
														assign node40071 = (inp[8]) ? 4'b0001 : 4'b0000;
											assign node40074 = (inp[4]) ? node40100 : node40075;
												assign node40075 = (inp[7]) ? node40091 : node40076;
													assign node40076 = (inp[8]) ? node40086 : node40077;
														assign node40077 = (inp[14]) ? node40079 : 4'b0000;
															assign node40079 = (inp[12]) ? node40083 : node40080;
																assign node40080 = (inp[9]) ? 4'b0000 : 4'b0100;
																assign node40083 = (inp[9]) ? 4'b0100 : 4'b0000;
														assign node40086 = (inp[9]) ? node40088 : 4'b0101;
															assign node40088 = (inp[12]) ? 4'b0101 : 4'b0001;
													assign node40091 = (inp[8]) ? node40093 : 4'b0001;
														assign node40093 = (inp[12]) ? node40097 : node40094;
															assign node40094 = (inp[9]) ? 4'b0000 : 4'b0100;
															assign node40097 = (inp[9]) ? 4'b0100 : 4'b0000;
												assign node40100 = (inp[8]) ? node40120 : node40101;
													assign node40101 = (inp[7]) ? node40107 : node40102;
														assign node40102 = (inp[12]) ? node40104 : 4'b0100;
															assign node40104 = (inp[9]) ? 4'b0000 : 4'b0100;
														assign node40107 = (inp[14]) ? node40113 : node40108;
															assign node40108 = (inp[9]) ? 4'b0101 : node40109;
																assign node40109 = (inp[12]) ? 4'b0101 : 4'b0001;
															assign node40113 = (inp[9]) ? node40117 : node40114;
																assign node40114 = (inp[12]) ? 4'b0101 : 4'b0001;
																assign node40117 = (inp[12]) ? 4'b0001 : 4'b0101;
													assign node40120 = (inp[7]) ? node40126 : node40121;
														assign node40121 = (inp[14]) ? 4'b0001 : node40122;
															assign node40122 = (inp[9]) ? 4'b0001 : 4'b0101;
														assign node40126 = (inp[14]) ? 4'b0100 : node40127;
															assign node40127 = (inp[12]) ? node40131 : node40128;
																assign node40128 = (inp[9]) ? 4'b0100 : 4'b0000;
																assign node40131 = (inp[9]) ? 4'b0000 : 4'b0100;
				assign node40135 = (inp[13]) ? node43991 : node40136;
					assign node40136 = (inp[1]) ? node42406 : node40137;
						assign node40137 = (inp[2]) ? node41405 : node40138;
							assign node40138 = (inp[3]) ? node40782 : node40139;
								assign node40139 = (inp[4]) ? node40457 : node40140;
									assign node40140 = (inp[5]) ? node40306 : node40141;
										assign node40141 = (inp[7]) ? node40223 : node40142;
											assign node40142 = (inp[15]) ? node40178 : node40143;
												assign node40143 = (inp[0]) ? node40155 : node40144;
													assign node40144 = (inp[14]) ? node40148 : node40145;
														assign node40145 = (inp[8]) ? 4'b0110 : 4'b0111;
														assign node40148 = (inp[8]) ? 4'b0111 : node40149;
															assign node40149 = (inp[12]) ? 4'b0110 : node40150;
																assign node40150 = (inp[9]) ? 4'b0010 : 4'b0110;
													assign node40155 = (inp[12]) ? node40165 : node40156;
														assign node40156 = (inp[9]) ? 4'b0001 : node40157;
															assign node40157 = (inp[14]) ? node40161 : node40158;
																assign node40158 = (inp[8]) ? 4'b0100 : 4'b0101;
																assign node40161 = (inp[8]) ? 4'b0101 : 4'b0100;
														assign node40165 = (inp[9]) ? node40171 : node40166;
															assign node40166 = (inp[14]) ? node40168 : 4'b0001;
																assign node40168 = (inp[8]) ? 4'b0001 : 4'b0000;
															assign node40171 = (inp[8]) ? node40175 : node40172;
																assign node40172 = (inp[14]) ? 4'b0100 : 4'b0101;
																assign node40175 = (inp[14]) ? 4'b0101 : 4'b0100;
												assign node40178 = (inp[0]) ? node40200 : node40179;
													assign node40179 = (inp[14]) ? node40193 : node40180;
														assign node40180 = (inp[8]) ? node40186 : node40181;
															assign node40181 = (inp[9]) ? 4'b0001 : node40182;
																assign node40182 = (inp[12]) ? 4'b0001 : 4'b0101;
															assign node40186 = (inp[12]) ? node40190 : node40187;
																assign node40187 = (inp[9]) ? 4'b0000 : 4'b0100;
																assign node40190 = (inp[9]) ? 4'b0100 : 4'b0000;
														assign node40193 = (inp[8]) ? node40195 : 4'b0100;
															assign node40195 = (inp[9]) ? 4'b0101 : node40196;
																assign node40196 = (inp[12]) ? 4'b0001 : 4'b0101;
													assign node40200 = (inp[9]) ? node40212 : node40201;
														assign node40201 = (inp[12]) ? node40209 : node40202;
															assign node40202 = (inp[8]) ? node40206 : node40203;
																assign node40203 = (inp[14]) ? 4'b0110 : 4'b0111;
																assign node40206 = (inp[14]) ? 4'b0111 : 4'b0110;
															assign node40209 = (inp[8]) ? 4'b0011 : 4'b0010;
														assign node40212 = (inp[12]) ? node40220 : node40213;
															assign node40213 = (inp[8]) ? node40217 : node40214;
																assign node40214 = (inp[14]) ? 4'b0010 : 4'b0011;
																assign node40217 = (inp[14]) ? 4'b0011 : 4'b0010;
															assign node40220 = (inp[14]) ? 4'b0110 : 4'b0111;
											assign node40223 = (inp[15]) ? node40265 : node40224;
												assign node40224 = (inp[0]) ? node40248 : node40225;
													assign node40225 = (inp[8]) ? node40239 : node40226;
														assign node40226 = (inp[14]) ? node40232 : node40227;
															assign node40227 = (inp[9]) ? node40229 : 4'b0110;
																assign node40229 = (inp[12]) ? 4'b0110 : 4'b0010;
															assign node40232 = (inp[9]) ? node40236 : node40233;
																assign node40233 = (inp[12]) ? 4'b0011 : 4'b0111;
																assign node40236 = (inp[12]) ? 4'b0111 : 4'b0011;
														assign node40239 = (inp[14]) ? node40245 : node40240;
															assign node40240 = (inp[9]) ? node40242 : 4'b0011;
																assign node40242 = (inp[12]) ? 4'b0111 : 4'b0011;
															assign node40245 = (inp[12]) ? 4'b0010 : 4'b0110;
													assign node40248 = (inp[8]) ? node40260 : node40249;
														assign node40249 = (inp[14]) ? node40257 : node40250;
															assign node40250 = (inp[9]) ? node40254 : node40251;
																assign node40251 = (inp[12]) ? 4'b0000 : 4'b0100;
																assign node40254 = (inp[12]) ? 4'b0100 : 4'b0000;
															assign node40257 = (inp[9]) ? 4'b0101 : 4'b0001;
														assign node40260 = (inp[14]) ? 4'b0100 : node40261;
															assign node40261 = (inp[9]) ? 4'b0001 : 4'b0101;
												assign node40265 = (inp[0]) ? node40287 : node40266;
													assign node40266 = (inp[8]) ? node40278 : node40267;
														assign node40267 = (inp[14]) ? node40273 : node40268;
															assign node40268 = (inp[12]) ? 4'b0000 : node40269;
																assign node40269 = (inp[9]) ? 4'b0000 : 4'b0100;
															assign node40273 = (inp[12]) ? node40275 : 4'b0101;
																assign node40275 = (inp[9]) ? 4'b0101 : 4'b0001;
														assign node40278 = (inp[14]) ? node40280 : 4'b0101;
															assign node40280 = (inp[12]) ? node40284 : node40281;
																assign node40281 = (inp[9]) ? 4'b0000 : 4'b0100;
																assign node40284 = (inp[9]) ? 4'b0100 : 4'b0000;
													assign node40287 = (inp[12]) ? node40295 : node40288;
														assign node40288 = (inp[9]) ? 4'b0010 : node40289;
															assign node40289 = (inp[14]) ? 4'b0110 : node40290;
																assign node40290 = (inp[8]) ? 4'b0111 : 4'b0110;
														assign node40295 = (inp[9]) ? node40301 : node40296;
															assign node40296 = (inp[8]) ? 4'b0010 : node40297;
																assign node40297 = (inp[14]) ? 4'b0011 : 4'b0010;
															assign node40301 = (inp[8]) ? 4'b0110 : node40302;
																assign node40302 = (inp[14]) ? 4'b0111 : 4'b0110;
										assign node40306 = (inp[12]) ? node40384 : node40307;
											assign node40307 = (inp[9]) ? node40345 : node40308;
												assign node40308 = (inp[7]) ? node40326 : node40309;
													assign node40309 = (inp[0]) ? node40319 : node40310;
														assign node40310 = (inp[15]) ? node40316 : node40311;
															assign node40311 = (inp[8]) ? node40313 : 4'b0111;
																assign node40313 = (inp[14]) ? 4'b0111 : 4'b0110;
															assign node40316 = (inp[8]) ? 4'b0101 : 4'b0100;
														assign node40319 = (inp[15]) ? 4'b0111 : node40320;
															assign node40320 = (inp[14]) ? 4'b0101 : node40321;
																assign node40321 = (inp[8]) ? 4'b0100 : 4'b0101;
													assign node40326 = (inp[14]) ? node40338 : node40327;
														assign node40327 = (inp[8]) ? node40333 : node40328;
															assign node40328 = (inp[0]) ? 4'b0110 : node40329;
																assign node40329 = (inp[15]) ? 4'b0100 : 4'b0110;
															assign node40333 = (inp[0]) ? 4'b0101 : node40334;
																assign node40334 = (inp[15]) ? 4'b0101 : 4'b0111;
														assign node40338 = (inp[8]) ? node40340 : 4'b0111;
															assign node40340 = (inp[15]) ? 4'b0110 : node40341;
																assign node40341 = (inp[0]) ? 4'b0100 : 4'b0110;
												assign node40345 = (inp[14]) ? node40363 : node40346;
													assign node40346 = (inp[7]) ? node40354 : node40347;
														assign node40347 = (inp[8]) ? 4'b0010 : node40348;
															assign node40348 = (inp[15]) ? node40350 : 4'b0011;
																assign node40350 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node40354 = (inp[8]) ? node40358 : node40355;
															assign node40355 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node40358 = (inp[0]) ? 4'b0001 : node40359;
																assign node40359 = (inp[15]) ? 4'b0001 : 4'b0011;
													assign node40363 = (inp[15]) ? node40375 : node40364;
														assign node40364 = (inp[0]) ? node40368 : node40365;
															assign node40365 = (inp[7]) ? 4'b0011 : 4'b0010;
															assign node40368 = (inp[8]) ? node40372 : node40369;
																assign node40369 = (inp[7]) ? 4'b0001 : 4'b0000;
																assign node40372 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node40375 = (inp[0]) ? node40377 : 4'b0000;
															assign node40377 = (inp[7]) ? node40381 : node40378;
																assign node40378 = (inp[8]) ? 4'b0011 : 4'b0010;
																assign node40381 = (inp[8]) ? 4'b0010 : 4'b0011;
											assign node40384 = (inp[9]) ? node40416 : node40385;
												assign node40385 = (inp[7]) ? node40403 : node40386;
													assign node40386 = (inp[15]) ? node40396 : node40387;
														assign node40387 = (inp[0]) ? node40391 : node40388;
															assign node40388 = (inp[14]) ? 4'b0011 : 4'b0010;
															assign node40391 = (inp[14]) ? 4'b0000 : node40392;
																assign node40392 = (inp[8]) ? 4'b0000 : 4'b0001;
														assign node40396 = (inp[0]) ? node40398 : 4'b0000;
															assign node40398 = (inp[14]) ? node40400 : 4'b0011;
																assign node40400 = (inp[8]) ? 4'b0011 : 4'b0010;
													assign node40403 = (inp[15]) ? node40413 : node40404;
														assign node40404 = (inp[0]) ? 4'b0001 : node40405;
															assign node40405 = (inp[14]) ? node40409 : node40406;
																assign node40406 = (inp[8]) ? 4'b0011 : 4'b0010;
																assign node40409 = (inp[8]) ? 4'b0010 : 4'b0011;
														assign node40413 = (inp[0]) ? 4'b0010 : 4'b0001;
												assign node40416 = (inp[14]) ? node40442 : node40417;
													assign node40417 = (inp[8]) ? node40431 : node40418;
														assign node40418 = (inp[7]) ? node40424 : node40419;
															assign node40419 = (inp[0]) ? 4'b0101 : node40420;
																assign node40420 = (inp[15]) ? 4'b0111 : 4'b0101;
															assign node40424 = (inp[0]) ? node40428 : node40425;
																assign node40425 = (inp[15]) ? 4'b0110 : 4'b0100;
																assign node40428 = (inp[15]) ? 4'b0100 : 4'b0110;
														assign node40431 = (inp[7]) ? node40435 : node40432;
															assign node40432 = (inp[15]) ? 4'b0100 : 4'b0110;
															assign node40435 = (inp[0]) ? node40439 : node40436;
																assign node40436 = (inp[15]) ? 4'b0111 : 4'b0101;
																assign node40439 = (inp[15]) ? 4'b0101 : 4'b0111;
													assign node40442 = (inp[0]) ? node40454 : node40443;
														assign node40443 = (inp[15]) ? node40449 : node40444;
															assign node40444 = (inp[8]) ? 4'b0101 : node40445;
																assign node40445 = (inp[7]) ? 4'b0101 : 4'b0100;
															assign node40449 = (inp[8]) ? node40451 : 4'b0111;
																assign node40451 = (inp[7]) ? 4'b0110 : 4'b0111;
														assign node40454 = (inp[15]) ? 4'b0101 : 4'b0111;
									assign node40457 = (inp[15]) ? node40621 : node40458;
										assign node40458 = (inp[0]) ? node40538 : node40459;
											assign node40459 = (inp[5]) ? node40499 : node40460;
												assign node40460 = (inp[7]) ? node40480 : node40461;
													assign node40461 = (inp[12]) ? node40469 : node40462;
														assign node40462 = (inp[8]) ? node40466 : node40463;
															assign node40463 = (inp[14]) ? 4'b0010 : 4'b0011;
															assign node40466 = (inp[14]) ? 4'b0011 : 4'b0010;
														assign node40469 = (inp[9]) ? node40475 : node40470;
															assign node40470 = (inp[8]) ? 4'b0110 : node40471;
																assign node40471 = (inp[14]) ? 4'b0110 : 4'b0111;
															assign node40475 = (inp[8]) ? node40477 : 4'b0010;
																assign node40477 = (inp[14]) ? 4'b0011 : 4'b0010;
													assign node40480 = (inp[12]) ? node40492 : node40481;
														assign node40481 = (inp[9]) ? node40485 : node40482;
															assign node40482 = (inp[14]) ? 4'b0011 : 4'b0010;
															assign node40485 = (inp[14]) ? node40489 : node40486;
																assign node40486 = (inp[8]) ? 4'b0111 : 4'b0110;
																assign node40489 = (inp[8]) ? 4'b0110 : 4'b0111;
														assign node40492 = (inp[9]) ? node40494 : 4'b0111;
															assign node40494 = (inp[14]) ? 4'b0011 : node40495;
																assign node40495 = (inp[8]) ? 4'b0011 : 4'b0010;
												assign node40499 = (inp[9]) ? node40519 : node40500;
													assign node40500 = (inp[12]) ? node40510 : node40501;
														assign node40501 = (inp[7]) ? 4'b0010 : node40502;
															assign node40502 = (inp[8]) ? node40506 : node40503;
																assign node40503 = (inp[14]) ? 4'b0010 : 4'b0011;
																assign node40506 = (inp[14]) ? 4'b0011 : 4'b0010;
														assign node40510 = (inp[14]) ? node40512 : 4'b0100;
															assign node40512 = (inp[8]) ? node40516 : node40513;
																assign node40513 = (inp[7]) ? 4'b0101 : 4'b0100;
																assign node40516 = (inp[7]) ? 4'b0100 : 4'b0101;
													assign node40519 = (inp[12]) ? node40529 : node40520;
														assign node40520 = (inp[7]) ? node40522 : 4'b0100;
															assign node40522 = (inp[14]) ? node40526 : node40523;
																assign node40523 = (inp[8]) ? 4'b0101 : 4'b0100;
																assign node40526 = (inp[8]) ? 4'b0100 : 4'b0101;
														assign node40529 = (inp[7]) ? 4'b0001 : node40530;
															assign node40530 = (inp[14]) ? node40534 : node40531;
																assign node40531 = (inp[8]) ? 4'b0000 : 4'b0001;
																assign node40534 = (inp[8]) ? 4'b0001 : 4'b0000;
											assign node40538 = (inp[5]) ? node40580 : node40539;
												assign node40539 = (inp[12]) ? node40557 : node40540;
													assign node40540 = (inp[9]) ? node40550 : node40541;
														assign node40541 = (inp[8]) ? 4'b0000 : node40542;
															assign node40542 = (inp[7]) ? node40546 : node40543;
																assign node40543 = (inp[14]) ? 4'b0000 : 4'b0001;
																assign node40546 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node40550 = (inp[14]) ? node40552 : 4'b0100;
															assign node40552 = (inp[7]) ? node40554 : 4'b0100;
																assign node40554 = (inp[8]) ? 4'b0100 : 4'b0101;
													assign node40557 = (inp[9]) ? node40569 : node40558;
														assign node40558 = (inp[7]) ? node40564 : node40559;
															assign node40559 = (inp[14]) ? 4'b0100 : node40560;
																assign node40560 = (inp[8]) ? 4'b0100 : 4'b0101;
															assign node40564 = (inp[8]) ? node40566 : 4'b0101;
																assign node40566 = (inp[14]) ? 4'b0100 : 4'b0101;
														assign node40569 = (inp[14]) ? node40575 : node40570;
															assign node40570 = (inp[8]) ? node40572 : 4'b0001;
																assign node40572 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node40575 = (inp[8]) ? node40577 : 4'b0000;
																assign node40577 = (inp[7]) ? 4'b0000 : 4'b0001;
												assign node40580 = (inp[12]) ? node40600 : node40581;
													assign node40581 = (inp[9]) ? node40593 : node40582;
														assign node40582 = (inp[14]) ? node40588 : node40583;
															assign node40583 = (inp[8]) ? node40585 : 4'b0001;
																assign node40585 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node40588 = (inp[8]) ? node40590 : 4'b0000;
																assign node40590 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node40593 = (inp[14]) ? node40597 : node40594;
															assign node40594 = (inp[8]) ? 4'b0110 : 4'b0111;
															assign node40597 = (inp[8]) ? 4'b0111 : 4'b0110;
													assign node40600 = (inp[9]) ? node40608 : node40601;
														assign node40601 = (inp[7]) ? 4'b0111 : node40602;
															assign node40602 = (inp[14]) ? 4'b0111 : node40603;
																assign node40603 = (inp[8]) ? 4'b0110 : 4'b0111;
														assign node40608 = (inp[14]) ? node40614 : node40609;
															assign node40609 = (inp[7]) ? node40611 : 4'b0011;
																assign node40611 = (inp[8]) ? 4'b0011 : 4'b0010;
															assign node40614 = (inp[8]) ? node40618 : node40615;
																assign node40615 = (inp[7]) ? 4'b0011 : 4'b0010;
																assign node40618 = (inp[7]) ? 4'b0010 : 4'b0011;
										assign node40621 = (inp[0]) ? node40701 : node40622;
											assign node40622 = (inp[5]) ? node40666 : node40623;
												assign node40623 = (inp[14]) ? node40649 : node40624;
													assign node40624 = (inp[8]) ? node40636 : node40625;
														assign node40625 = (inp[7]) ? node40631 : node40626;
															assign node40626 = (inp[12]) ? 4'b0101 : node40627;
																assign node40627 = (inp[9]) ? 4'b0101 : 4'b0001;
															assign node40631 = (inp[9]) ? 4'b0100 : node40632;
																assign node40632 = (inp[12]) ? 4'b0100 : 4'b0000;
														assign node40636 = (inp[7]) ? node40644 : node40637;
															assign node40637 = (inp[9]) ? node40641 : node40638;
																assign node40638 = (inp[12]) ? 4'b0100 : 4'b0000;
																assign node40641 = (inp[12]) ? 4'b0000 : 4'b0100;
															assign node40644 = (inp[12]) ? 4'b0001 : node40645;
																assign node40645 = (inp[9]) ? 4'b0101 : 4'b0001;
													assign node40649 = (inp[7]) ? node40659 : node40650;
														assign node40650 = (inp[8]) ? node40654 : node40651;
															assign node40651 = (inp[12]) ? 4'b0100 : 4'b0000;
															assign node40654 = (inp[12]) ? node40656 : 4'b0001;
																assign node40656 = (inp[9]) ? 4'b0001 : 4'b0101;
														assign node40659 = (inp[8]) ? 4'b0000 : node40660;
															assign node40660 = (inp[12]) ? 4'b0001 : node40661;
																assign node40661 = (inp[9]) ? 4'b0101 : 4'b0001;
												assign node40666 = (inp[12]) ? node40680 : node40667;
													assign node40667 = (inp[9]) ? node40673 : node40668;
														assign node40668 = (inp[7]) ? node40670 : 4'b0001;
															assign node40670 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node40673 = (inp[8]) ? 4'b0111 : node40674;
															assign node40674 = (inp[7]) ? 4'b0110 : node40675;
																assign node40675 = (inp[14]) ? 4'b0110 : 4'b0111;
													assign node40680 = (inp[9]) ? node40694 : node40681;
														assign node40681 = (inp[14]) ? node40687 : node40682;
															assign node40682 = (inp[7]) ? 4'b0110 : node40683;
																assign node40683 = (inp[8]) ? 4'b0110 : 4'b0111;
															assign node40687 = (inp[7]) ? node40691 : node40688;
																assign node40688 = (inp[8]) ? 4'b0111 : 4'b0110;
																assign node40691 = (inp[8]) ? 4'b0110 : 4'b0111;
														assign node40694 = (inp[8]) ? 4'b0010 : node40695;
															assign node40695 = (inp[7]) ? node40697 : 4'b0011;
																assign node40697 = (inp[14]) ? 4'b0011 : 4'b0010;
											assign node40701 = (inp[5]) ? node40743 : node40702;
												assign node40702 = (inp[7]) ? node40726 : node40703;
													assign node40703 = (inp[9]) ? node40713 : node40704;
														assign node40704 = (inp[12]) ? node40710 : node40705;
															assign node40705 = (inp[8]) ? node40707 : 4'b0010;
																assign node40707 = (inp[14]) ? 4'b0011 : 4'b0010;
															assign node40710 = (inp[8]) ? 4'b0110 : 4'b0111;
														assign node40713 = (inp[12]) ? node40719 : node40714;
															assign node40714 = (inp[8]) ? 4'b0111 : node40715;
																assign node40715 = (inp[14]) ? 4'b0110 : 4'b0111;
															assign node40719 = (inp[8]) ? node40723 : node40720;
																assign node40720 = (inp[14]) ? 4'b0010 : 4'b0011;
																assign node40723 = (inp[14]) ? 4'b0011 : 4'b0010;
													assign node40726 = (inp[9]) ? node40736 : node40727;
														assign node40727 = (inp[12]) ? node40731 : node40728;
															assign node40728 = (inp[14]) ? 4'b0011 : 4'b0010;
															assign node40731 = (inp[14]) ? 4'b0111 : node40732;
																assign node40732 = (inp[8]) ? 4'b0111 : 4'b0110;
														assign node40736 = (inp[12]) ? 4'b0010 : node40737;
															assign node40737 = (inp[14]) ? 4'b0110 : node40738;
																assign node40738 = (inp[8]) ? 4'b0111 : 4'b0110;
												assign node40743 = (inp[9]) ? node40759 : node40744;
													assign node40744 = (inp[12]) ? node40752 : node40745;
														assign node40745 = (inp[14]) ? 4'b0011 : node40746;
															assign node40746 = (inp[8]) ? node40748 : 4'b0010;
																assign node40748 = (inp[7]) ? 4'b0011 : 4'b0010;
														assign node40752 = (inp[14]) ? node40754 : 4'b0100;
															assign node40754 = (inp[7]) ? node40756 : 4'b0101;
																assign node40756 = (inp[8]) ? 4'b0100 : 4'b0101;
													assign node40759 = (inp[12]) ? node40773 : node40760;
														assign node40760 = (inp[7]) ? node40768 : node40761;
															assign node40761 = (inp[14]) ? node40765 : node40762;
																assign node40762 = (inp[8]) ? 4'b0100 : 4'b0101;
																assign node40765 = (inp[8]) ? 4'b0101 : 4'b0100;
															assign node40768 = (inp[14]) ? node40770 : 4'b0100;
																assign node40770 = (inp[8]) ? 4'b0100 : 4'b0101;
														assign node40773 = (inp[8]) ? 4'b0001 : node40774;
															assign node40774 = (inp[14]) ? node40778 : node40775;
																assign node40775 = (inp[7]) ? 4'b0000 : 4'b0001;
																assign node40778 = (inp[7]) ? 4'b0001 : 4'b0000;
								assign node40782 = (inp[0]) ? node41100 : node40783;
									assign node40783 = (inp[15]) ? node40963 : node40784;
										assign node40784 = (inp[5]) ? node40868 : node40785;
											assign node40785 = (inp[12]) ? node40825 : node40786;
												assign node40786 = (inp[9]) ? node40806 : node40787;
													assign node40787 = (inp[4]) ? node40793 : node40788;
														assign node40788 = (inp[8]) ? node40790 : 4'b0111;
															assign node40790 = (inp[14]) ? 4'b0111 : 4'b0110;
														assign node40793 = (inp[7]) ? node40801 : node40794;
															assign node40794 = (inp[14]) ? node40798 : node40795;
																assign node40795 = (inp[8]) ? 4'b0010 : 4'b0011;
																assign node40798 = (inp[8]) ? 4'b0011 : 4'b0010;
															assign node40801 = (inp[8]) ? 4'b0011 : node40802;
																assign node40802 = (inp[14]) ? 4'b0011 : 4'b0010;
													assign node40806 = (inp[4]) ? node40816 : node40807;
														assign node40807 = (inp[7]) ? 4'b0010 : node40808;
															assign node40808 = (inp[14]) ? node40812 : node40809;
																assign node40809 = (inp[8]) ? 4'b0010 : 4'b0011;
																assign node40812 = (inp[8]) ? 4'b0011 : 4'b0010;
														assign node40816 = (inp[7]) ? 4'b0100 : node40817;
															assign node40817 = (inp[14]) ? node40821 : node40818;
																assign node40818 = (inp[8]) ? 4'b0100 : 4'b0101;
																assign node40821 = (inp[8]) ? 4'b0101 : 4'b0100;
												assign node40825 = (inp[9]) ? node40845 : node40826;
													assign node40826 = (inp[4]) ? node40834 : node40827;
														assign node40827 = (inp[7]) ? node40829 : 4'b0011;
															assign node40829 = (inp[8]) ? node40831 : 4'b0010;
																assign node40831 = (inp[14]) ? 4'b0010 : 4'b0011;
														assign node40834 = (inp[7]) ? node40840 : node40835;
															assign node40835 = (inp[14]) ? node40837 : 4'b0100;
																assign node40837 = (inp[8]) ? 4'b0101 : 4'b0100;
															assign node40840 = (inp[8]) ? node40842 : 4'b0101;
																assign node40842 = (inp[14]) ? 4'b0100 : 4'b0101;
													assign node40845 = (inp[4]) ? node40859 : node40846;
														assign node40846 = (inp[7]) ? node40854 : node40847;
															assign node40847 = (inp[8]) ? node40851 : node40848;
																assign node40848 = (inp[14]) ? 4'b0100 : 4'b0101;
																assign node40851 = (inp[14]) ? 4'b0101 : 4'b0100;
															assign node40854 = (inp[14]) ? node40856 : 4'b0101;
																assign node40856 = (inp[8]) ? 4'b0100 : 4'b0101;
														assign node40859 = (inp[14]) ? 4'b0001 : node40860;
															assign node40860 = (inp[8]) ? node40864 : node40861;
																assign node40861 = (inp[7]) ? 4'b0000 : 4'b0001;
																assign node40864 = (inp[7]) ? 4'b0001 : 4'b0000;
											assign node40868 = (inp[12]) ? node40926 : node40869;
												assign node40869 = (inp[14]) ? node40899 : node40870;
													assign node40870 = (inp[9]) ? node40884 : node40871;
														assign node40871 = (inp[4]) ? node40879 : node40872;
															assign node40872 = (inp[8]) ? node40876 : node40873;
																assign node40873 = (inp[7]) ? 4'b0100 : 4'b0101;
																assign node40876 = (inp[7]) ? 4'b0101 : 4'b0100;
															assign node40879 = (inp[7]) ? 4'b0000 : node40880;
																assign node40880 = (inp[8]) ? 4'b0000 : 4'b0001;
														assign node40884 = (inp[4]) ? node40892 : node40885;
															assign node40885 = (inp[7]) ? node40889 : node40886;
																assign node40886 = (inp[8]) ? 4'b0000 : 4'b0001;
																assign node40889 = (inp[8]) ? 4'b0001 : 4'b0000;
															assign node40892 = (inp[7]) ? node40896 : node40893;
																assign node40893 = (inp[8]) ? 4'b0100 : 4'b0101;
																assign node40896 = (inp[8]) ? 4'b0101 : 4'b0100;
													assign node40899 = (inp[7]) ? node40913 : node40900;
														assign node40900 = (inp[8]) ? node40906 : node40901;
															assign node40901 = (inp[9]) ? 4'b0100 : node40902;
																assign node40902 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node40906 = (inp[4]) ? node40910 : node40907;
																assign node40907 = (inp[9]) ? 4'b0001 : 4'b0101;
																assign node40910 = (inp[9]) ? 4'b0101 : 4'b0001;
														assign node40913 = (inp[8]) ? node40921 : node40914;
															assign node40914 = (inp[4]) ? node40918 : node40915;
																assign node40915 = (inp[9]) ? 4'b0001 : 4'b0101;
																assign node40918 = (inp[9]) ? 4'b0101 : 4'b0001;
															assign node40921 = (inp[4]) ? 4'b0100 : node40922;
																assign node40922 = (inp[9]) ? 4'b0000 : 4'b0100;
												assign node40926 = (inp[9]) ? node40950 : node40927;
													assign node40927 = (inp[4]) ? node40939 : node40928;
														assign node40928 = (inp[8]) ? node40934 : node40929;
															assign node40929 = (inp[14]) ? 4'b0000 : node40930;
																assign node40930 = (inp[7]) ? 4'b0000 : 4'b0001;
															assign node40934 = (inp[14]) ? 4'b0001 : node40935;
																assign node40935 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node40939 = (inp[14]) ? node40945 : node40940;
															assign node40940 = (inp[7]) ? 4'b0100 : node40941;
																assign node40941 = (inp[8]) ? 4'b0100 : 4'b0101;
															assign node40945 = (inp[7]) ? 4'b0101 : node40946;
																assign node40946 = (inp[8]) ? 4'b0101 : 4'b0100;
													assign node40950 = (inp[4]) ? node40956 : node40951;
														assign node40951 = (inp[8]) ? 4'b0100 : node40952;
															assign node40952 = (inp[7]) ? 4'b0101 : 4'b0100;
														assign node40956 = (inp[7]) ? 4'b0000 : node40957;
															assign node40957 = (inp[14]) ? node40959 : 4'b0001;
																assign node40959 = (inp[8]) ? 4'b0001 : 4'b0000;
										assign node40963 = (inp[5]) ? node41039 : node40964;
											assign node40964 = (inp[12]) ? node41000 : node40965;
												assign node40965 = (inp[4]) ? node40985 : node40966;
													assign node40966 = (inp[9]) ? node40976 : node40967;
														assign node40967 = (inp[14]) ? node40969 : 4'b0100;
															assign node40969 = (inp[7]) ? node40973 : node40970;
																assign node40970 = (inp[8]) ? 4'b0101 : 4'b0100;
																assign node40973 = (inp[8]) ? 4'b0100 : 4'b0101;
														assign node40976 = (inp[14]) ? node40978 : 4'b0000;
															assign node40978 = (inp[7]) ? node40982 : node40979;
																assign node40979 = (inp[8]) ? 4'b0001 : 4'b0000;
																assign node40982 = (inp[8]) ? 4'b0000 : 4'b0001;
													assign node40985 = (inp[9]) ? 4'b0110 : node40986;
														assign node40986 = (inp[14]) ? node40992 : node40987;
															assign node40987 = (inp[7]) ? node40989 : 4'b0000;
																assign node40989 = (inp[8]) ? 4'b0001 : 4'b0000;
															assign node40992 = (inp[8]) ? node40996 : node40993;
																assign node40993 = (inp[7]) ? 4'b0001 : 4'b0000;
																assign node40996 = (inp[7]) ? 4'b0000 : 4'b0001;
												assign node41000 = (inp[4]) ? node41020 : node41001;
													assign node41001 = (inp[9]) ? node41011 : node41002;
														assign node41002 = (inp[14]) ? node41004 : 4'b0001;
															assign node41004 = (inp[8]) ? node41008 : node41005;
																assign node41005 = (inp[7]) ? 4'b0001 : 4'b0000;
																assign node41008 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node41011 = (inp[7]) ? 4'b0110 : node41012;
															assign node41012 = (inp[14]) ? node41016 : node41013;
																assign node41013 = (inp[8]) ? 4'b0110 : 4'b0111;
																assign node41016 = (inp[8]) ? 4'b0111 : 4'b0110;
													assign node41020 = (inp[9]) ? node41034 : node41021;
														assign node41021 = (inp[8]) ? node41029 : node41022;
															assign node41022 = (inp[14]) ? node41026 : node41023;
																assign node41023 = (inp[7]) ? 4'b0110 : 4'b0111;
																assign node41026 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node41029 = (inp[14]) ? 4'b0110 : node41030;
																assign node41030 = (inp[7]) ? 4'b0111 : 4'b0110;
														assign node41034 = (inp[14]) ? 4'b0010 : node41035;
															assign node41035 = (inp[7]) ? 4'b0011 : 4'b0010;
											assign node41039 = (inp[12]) ? node41071 : node41040;
												assign node41040 = (inp[8]) ? node41062 : node41041;
													assign node41041 = (inp[7]) ? node41049 : node41042;
														assign node41042 = (inp[14]) ? 4'b0110 : node41043;
															assign node41043 = (inp[9]) ? node41045 : 4'b0011;
																assign node41045 = (inp[4]) ? 4'b0111 : 4'b0011;
														assign node41049 = (inp[14]) ? node41057 : node41050;
															assign node41050 = (inp[9]) ? node41054 : node41051;
																assign node41051 = (inp[4]) ? 4'b0010 : 4'b0110;
																assign node41054 = (inp[4]) ? 4'b0110 : 4'b0010;
															assign node41057 = (inp[9]) ? 4'b0011 : node41058;
																assign node41058 = (inp[4]) ? 4'b0011 : 4'b0111;
													assign node41062 = (inp[14]) ? node41066 : node41063;
														assign node41063 = (inp[7]) ? 4'b0011 : 4'b0010;
														assign node41066 = (inp[9]) ? 4'b0010 : node41067;
															assign node41067 = (inp[4]) ? 4'b0010 : 4'b0110;
												assign node41071 = (inp[4]) ? node41083 : node41072;
													assign node41072 = (inp[9]) ? node41078 : node41073;
														assign node41073 = (inp[7]) ? node41075 : 4'b0010;
															assign node41075 = (inp[14]) ? 4'b0010 : 4'b0011;
														assign node41078 = (inp[14]) ? node41080 : 4'b0110;
															assign node41080 = (inp[8]) ? 4'b0111 : 4'b0110;
													assign node41083 = (inp[9]) ? node41095 : node41084;
														assign node41084 = (inp[8]) ? node41090 : node41085;
															assign node41085 = (inp[14]) ? node41087 : 4'b0110;
																assign node41087 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node41090 = (inp[14]) ? 4'b0111 : node41091;
																assign node41091 = (inp[7]) ? 4'b0111 : 4'b0110;
														assign node41095 = (inp[7]) ? node41097 : 4'b0011;
															assign node41097 = (inp[14]) ? 4'b0011 : 4'b0010;
									assign node41100 = (inp[15]) ? node41260 : node41101;
										assign node41101 = (inp[5]) ? node41175 : node41102;
											assign node41102 = (inp[9]) ? node41144 : node41103;
												assign node41103 = (inp[12]) ? node41123 : node41104;
													assign node41104 = (inp[4]) ? node41114 : node41105;
														assign node41105 = (inp[7]) ? 4'b0101 : node41106;
															assign node41106 = (inp[8]) ? node41110 : node41107;
																assign node41107 = (inp[14]) ? 4'b0100 : 4'b0101;
																assign node41110 = (inp[14]) ? 4'b0101 : 4'b0100;
														assign node41114 = (inp[14]) ? node41116 : 4'b0001;
															assign node41116 = (inp[7]) ? node41120 : node41117;
																assign node41117 = (inp[8]) ? 4'b0001 : 4'b0000;
																assign node41120 = (inp[8]) ? 4'b0000 : 4'b0001;
													assign node41123 = (inp[4]) ? node41133 : node41124;
														assign node41124 = (inp[8]) ? node41126 : 4'b0001;
															assign node41126 = (inp[7]) ? node41130 : node41127;
																assign node41127 = (inp[14]) ? 4'b0001 : 4'b0000;
																assign node41130 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node41133 = (inp[14]) ? node41139 : node41134;
															assign node41134 = (inp[7]) ? 4'b0111 : node41135;
																assign node41135 = (inp[8]) ? 4'b0110 : 4'b0111;
															assign node41139 = (inp[7]) ? node41141 : 4'b0110;
																assign node41141 = (inp[8]) ? 4'b0110 : 4'b0111;
												assign node41144 = (inp[4]) ? node41160 : node41145;
													assign node41145 = (inp[12]) ? node41153 : node41146;
														assign node41146 = (inp[14]) ? node41148 : 4'b0000;
															assign node41148 = (inp[8]) ? 4'b0000 : node41149;
																assign node41149 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node41153 = (inp[14]) ? node41155 : 4'b0110;
															assign node41155 = (inp[7]) ? node41157 : 4'b0111;
																assign node41157 = (inp[8]) ? 4'b0110 : 4'b0111;
													assign node41160 = (inp[12]) ? 4'b0010 : node41161;
														assign node41161 = (inp[14]) ? node41167 : node41162;
															assign node41162 = (inp[7]) ? 4'b0111 : node41163;
																assign node41163 = (inp[8]) ? 4'b0110 : 4'b0111;
															assign node41167 = (inp[8]) ? node41171 : node41168;
																assign node41168 = (inp[7]) ? 4'b0111 : 4'b0110;
																assign node41171 = (inp[7]) ? 4'b0110 : 4'b0111;
											assign node41175 = (inp[9]) ? node41221 : node41176;
												assign node41176 = (inp[7]) ? node41196 : node41177;
													assign node41177 = (inp[4]) ? node41183 : node41178;
														assign node41178 = (inp[12]) ? node41180 : 4'b0110;
															assign node41180 = (inp[14]) ? 4'b0011 : 4'b0010;
														assign node41183 = (inp[12]) ? node41189 : node41184;
															assign node41184 = (inp[14]) ? node41186 : 4'b0011;
																assign node41186 = (inp[8]) ? 4'b0011 : 4'b0010;
															assign node41189 = (inp[8]) ? node41193 : node41190;
																assign node41190 = (inp[14]) ? 4'b0110 : 4'b0111;
																assign node41193 = (inp[14]) ? 4'b0111 : 4'b0110;
													assign node41196 = (inp[4]) ? node41210 : node41197;
														assign node41197 = (inp[12]) ? node41203 : node41198;
															assign node41198 = (inp[14]) ? node41200 : 4'b0111;
																assign node41200 = (inp[8]) ? 4'b0110 : 4'b0111;
															assign node41203 = (inp[14]) ? node41207 : node41204;
																assign node41204 = (inp[8]) ? 4'b0011 : 4'b0010;
																assign node41207 = (inp[8]) ? 4'b0010 : 4'b0011;
														assign node41210 = (inp[12]) ? node41216 : node41211;
															assign node41211 = (inp[14]) ? 4'b0011 : node41212;
																assign node41212 = (inp[8]) ? 4'b0011 : 4'b0010;
															assign node41216 = (inp[8]) ? 4'b0111 : node41217;
																assign node41217 = (inp[14]) ? 4'b0111 : 4'b0110;
												assign node41221 = (inp[14]) ? node41243 : node41222;
													assign node41222 = (inp[4]) ? node41230 : node41223;
														assign node41223 = (inp[12]) ? node41225 : 4'b0011;
															assign node41225 = (inp[7]) ? node41227 : 4'b0111;
																assign node41227 = (inp[8]) ? 4'b0111 : 4'b0110;
														assign node41230 = (inp[12]) ? node41238 : node41231;
															assign node41231 = (inp[7]) ? node41235 : node41232;
																assign node41232 = (inp[8]) ? 4'b0110 : 4'b0111;
																assign node41235 = (inp[8]) ? 4'b0111 : 4'b0110;
															assign node41238 = (inp[7]) ? 4'b0011 : node41239;
																assign node41239 = (inp[8]) ? 4'b0010 : 4'b0011;
													assign node41243 = (inp[12]) ? node41253 : node41244;
														assign node41244 = (inp[4]) ? node41248 : node41245;
															assign node41245 = (inp[8]) ? 4'b0010 : 4'b0011;
															assign node41248 = (inp[8]) ? 4'b0110 : node41249;
																assign node41249 = (inp[7]) ? 4'b0111 : 4'b0110;
														assign node41253 = (inp[4]) ? 4'b0010 : node41254;
															assign node41254 = (inp[7]) ? 4'b0110 : node41255;
																assign node41255 = (inp[8]) ? 4'b0111 : 4'b0110;
										assign node41260 = (inp[5]) ? node41328 : node41261;
											assign node41261 = (inp[4]) ? node41293 : node41262;
												assign node41262 = (inp[9]) ? node41286 : node41263;
													assign node41263 = (inp[12]) ? node41277 : node41264;
														assign node41264 = (inp[7]) ? node41270 : node41265;
															assign node41265 = (inp[14]) ? 4'b0111 : node41266;
																assign node41266 = (inp[8]) ? 4'b0110 : 4'b0111;
															assign node41270 = (inp[8]) ? node41274 : node41271;
																assign node41271 = (inp[14]) ? 4'b0111 : 4'b0110;
																assign node41274 = (inp[14]) ? 4'b0110 : 4'b0111;
														assign node41277 = (inp[14]) ? 4'b0010 : node41278;
															assign node41278 = (inp[7]) ? node41282 : node41279;
																assign node41279 = (inp[8]) ? 4'b0010 : 4'b0011;
																assign node41282 = (inp[8]) ? 4'b0011 : 4'b0010;
													assign node41286 = (inp[12]) ? node41290 : node41287;
														assign node41287 = (inp[7]) ? 4'b0010 : 4'b0011;
														assign node41290 = (inp[14]) ? 4'b0101 : 4'b0100;
												assign node41293 = (inp[12]) ? node41307 : node41294;
													assign node41294 = (inp[9]) ? node41300 : node41295;
														assign node41295 = (inp[8]) ? node41297 : 4'b0011;
															assign node41297 = (inp[7]) ? 4'b0011 : 4'b0010;
														assign node41300 = (inp[14]) ? 4'b0101 : node41301;
															assign node41301 = (inp[8]) ? node41303 : 4'b0100;
																assign node41303 = (inp[7]) ? 4'b0101 : 4'b0100;
													assign node41307 = (inp[9]) ? node41317 : node41308;
														assign node41308 = (inp[14]) ? 4'b0100 : node41309;
															assign node41309 = (inp[8]) ? node41313 : node41310;
																assign node41310 = (inp[7]) ? 4'b0100 : 4'b0101;
																assign node41313 = (inp[7]) ? 4'b0101 : 4'b0100;
														assign node41317 = (inp[14]) ? node41323 : node41318;
															assign node41318 = (inp[7]) ? node41320 : 4'b0000;
																assign node41320 = (inp[8]) ? 4'b0001 : 4'b0000;
															assign node41323 = (inp[7]) ? node41325 : 4'b0001;
																assign node41325 = (inp[8]) ? 4'b0000 : 4'b0001;
											assign node41328 = (inp[7]) ? node41368 : node41329;
												assign node41329 = (inp[9]) ? node41349 : node41330;
													assign node41330 = (inp[4]) ? node41336 : node41331;
														assign node41331 = (inp[12]) ? 4'b0001 : node41332;
															assign node41332 = (inp[14]) ? 4'b0100 : 4'b0101;
														assign node41336 = (inp[12]) ? node41344 : node41337;
															assign node41337 = (inp[8]) ? node41341 : node41338;
																assign node41338 = (inp[14]) ? 4'b0000 : 4'b0001;
																assign node41341 = (inp[14]) ? 4'b0001 : 4'b0000;
															assign node41344 = (inp[8]) ? node41346 : 4'b0100;
																assign node41346 = (inp[14]) ? 4'b0101 : 4'b0100;
													assign node41349 = (inp[8]) ? node41361 : node41350;
														assign node41350 = (inp[14]) ? node41356 : node41351;
															assign node41351 = (inp[12]) ? 4'b0101 : node41352;
																assign node41352 = (inp[4]) ? 4'b0101 : 4'b0001;
															assign node41356 = (inp[4]) ? 4'b0000 : node41357;
																assign node41357 = (inp[12]) ? 4'b0100 : 4'b0000;
														assign node41361 = (inp[4]) ? node41365 : node41362;
															assign node41362 = (inp[12]) ? 4'b0100 : 4'b0000;
															assign node41365 = (inp[12]) ? 4'b0000 : 4'b0100;
												assign node41368 = (inp[9]) ? node41382 : node41369;
													assign node41369 = (inp[4]) ? node41373 : node41370;
														assign node41370 = (inp[12]) ? 4'b0000 : 4'b0100;
														assign node41373 = (inp[12]) ? node41377 : node41374;
															assign node41374 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node41377 = (inp[14]) ? 4'b0100 : node41378;
																assign node41378 = (inp[8]) ? 4'b0101 : 4'b0100;
													assign node41382 = (inp[14]) ? node41396 : node41383;
														assign node41383 = (inp[8]) ? node41391 : node41384;
															assign node41384 = (inp[12]) ? node41388 : node41385;
																assign node41385 = (inp[4]) ? 4'b0100 : 4'b0000;
																assign node41388 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node41391 = (inp[4]) ? node41393 : 4'b0101;
																assign node41393 = (inp[12]) ? 4'b0001 : 4'b0101;
														assign node41396 = (inp[8]) ? 4'b0100 : node41397;
															assign node41397 = (inp[12]) ? node41401 : node41398;
																assign node41398 = (inp[4]) ? 4'b0101 : 4'b0001;
																assign node41401 = (inp[4]) ? 4'b0001 : 4'b0101;
							assign node41405 = (inp[3]) ? node41851 : node41406;
								assign node41406 = (inp[8]) ? node41610 : node41407;
									assign node41407 = (inp[7]) ? node41513 : node41408;
										assign node41408 = (inp[15]) ? node41464 : node41409;
											assign node41409 = (inp[0]) ? node41431 : node41410;
												assign node41410 = (inp[4]) ? node41418 : node41411;
													assign node41411 = (inp[9]) ? node41415 : node41412;
														assign node41412 = (inp[12]) ? 4'b0010 : 4'b0110;
														assign node41415 = (inp[12]) ? 4'b0110 : 4'b0010;
													assign node41418 = (inp[5]) ? node41424 : node41419;
														assign node41419 = (inp[9]) ? node41421 : 4'b0010;
															assign node41421 = (inp[14]) ? 4'b0010 : 4'b0110;
														assign node41424 = (inp[9]) ? node41428 : node41425;
															assign node41425 = (inp[12]) ? 4'b0100 : 4'b0010;
															assign node41428 = (inp[12]) ? 4'b0000 : 4'b0100;
												assign node41431 = (inp[5]) ? node41451 : node41432;
													assign node41432 = (inp[4]) ? node41446 : node41433;
														assign node41433 = (inp[14]) ? node41441 : node41434;
															assign node41434 = (inp[12]) ? node41438 : node41435;
																assign node41435 = (inp[9]) ? 4'b0000 : 4'b0100;
																assign node41438 = (inp[9]) ? 4'b0100 : 4'b0000;
															assign node41441 = (inp[12]) ? 4'b0100 : node41442;
																assign node41442 = (inp[9]) ? 4'b0000 : 4'b0100;
														assign node41446 = (inp[9]) ? node41448 : 4'b0000;
															assign node41448 = (inp[12]) ? 4'b0000 : 4'b0100;
													assign node41451 = (inp[12]) ? node41457 : node41452;
														assign node41452 = (inp[4]) ? 4'b0000 : node41453;
															assign node41453 = (inp[9]) ? 4'b0000 : 4'b0100;
														assign node41457 = (inp[9]) ? node41461 : node41458;
															assign node41458 = (inp[4]) ? 4'b0110 : 4'b0000;
															assign node41461 = (inp[4]) ? 4'b0010 : 4'b0110;
											assign node41464 = (inp[0]) ? node41486 : node41465;
												assign node41465 = (inp[9]) ? node41473 : node41466;
													assign node41466 = (inp[4]) ? node41470 : node41467;
														assign node41467 = (inp[12]) ? 4'b0000 : 4'b0100;
														assign node41470 = (inp[12]) ? 4'b0100 : 4'b0000;
													assign node41473 = (inp[5]) ? node41479 : node41474;
														assign node41474 = (inp[12]) ? 4'b0100 : node41475;
															assign node41475 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node41479 = (inp[4]) ? node41483 : node41480;
															assign node41480 = (inp[12]) ? 4'b0110 : 4'b0000;
															assign node41483 = (inp[12]) ? 4'b0010 : 4'b0110;
												assign node41486 = (inp[5]) ? node41506 : node41487;
													assign node41487 = (inp[4]) ? node41501 : node41488;
														assign node41488 = (inp[14]) ? node41494 : node41489;
															assign node41489 = (inp[9]) ? node41491 : 4'b0010;
																assign node41491 = (inp[12]) ? 4'b0110 : 4'b0010;
															assign node41494 = (inp[9]) ? node41498 : node41495;
																assign node41495 = (inp[12]) ? 4'b0010 : 4'b0110;
																assign node41498 = (inp[12]) ? 4'b0110 : 4'b0010;
														assign node41501 = (inp[9]) ? node41503 : 4'b0110;
															assign node41503 = (inp[12]) ? 4'b0010 : 4'b0110;
													assign node41506 = (inp[4]) ? 4'b0100 : node41507;
														assign node41507 = (inp[12]) ? 4'b0100 : node41508;
															assign node41508 = (inp[9]) ? 4'b0010 : 4'b0110;
										assign node41513 = (inp[0]) ? node41557 : node41514;
											assign node41514 = (inp[15]) ? node41536 : node41515;
												assign node41515 = (inp[4]) ? node41521 : node41516;
													assign node41516 = (inp[14]) ? 4'b0011 : node41517;
														assign node41517 = (inp[12]) ? 4'b0011 : 4'b0111;
													assign node41521 = (inp[5]) ? node41529 : node41522;
														assign node41522 = (inp[12]) ? node41526 : node41523;
															assign node41523 = (inp[9]) ? 4'b0111 : 4'b0011;
															assign node41526 = (inp[9]) ? 4'b0011 : 4'b0111;
														assign node41529 = (inp[9]) ? node41533 : node41530;
															assign node41530 = (inp[12]) ? 4'b0101 : 4'b0011;
															assign node41533 = (inp[12]) ? 4'b0001 : 4'b0101;
												assign node41536 = (inp[12]) ? node41544 : node41537;
													assign node41537 = (inp[14]) ? node41539 : 4'b0001;
														assign node41539 = (inp[9]) ? node41541 : 4'b0001;
															assign node41541 = (inp[4]) ? 4'b0101 : 4'b0001;
													assign node41544 = (inp[5]) ? node41550 : node41545;
														assign node41545 = (inp[4]) ? node41547 : 4'b0101;
															assign node41547 = (inp[9]) ? 4'b0001 : 4'b0101;
														assign node41550 = (inp[4]) ? node41554 : node41551;
															assign node41551 = (inp[9]) ? 4'b0111 : 4'b0001;
															assign node41554 = (inp[9]) ? 4'b0011 : 4'b0111;
											assign node41557 = (inp[15]) ? node41587 : node41558;
												assign node41558 = (inp[5]) ? node41572 : node41559;
													assign node41559 = (inp[4]) ? node41567 : node41560;
														assign node41560 = (inp[12]) ? node41564 : node41561;
															assign node41561 = (inp[9]) ? 4'b0001 : 4'b0101;
															assign node41564 = (inp[9]) ? 4'b0101 : 4'b0001;
														assign node41567 = (inp[14]) ? node41569 : 4'b0101;
															assign node41569 = (inp[12]) ? 4'b0101 : 4'b0001;
													assign node41572 = (inp[4]) ? node41580 : node41573;
														assign node41573 = (inp[9]) ? node41577 : node41574;
															assign node41574 = (inp[12]) ? 4'b0001 : 4'b0101;
															assign node41577 = (inp[12]) ? 4'b0111 : 4'b0001;
														assign node41580 = (inp[12]) ? node41584 : node41581;
															assign node41581 = (inp[9]) ? 4'b0111 : 4'b0001;
															assign node41584 = (inp[9]) ? 4'b0011 : 4'b0111;
												assign node41587 = (inp[9]) ? node41595 : node41588;
													assign node41588 = (inp[12]) ? node41592 : node41589;
														assign node41589 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node41592 = (inp[4]) ? 4'b0111 : 4'b0011;
													assign node41595 = (inp[5]) ? node41605 : node41596;
														assign node41596 = (inp[14]) ? node41598 : 4'b0111;
															assign node41598 = (inp[4]) ? node41602 : node41599;
																assign node41599 = (inp[12]) ? 4'b0111 : 4'b0011;
																assign node41602 = (inp[12]) ? 4'b0011 : 4'b0111;
														assign node41605 = (inp[12]) ? node41607 : 4'b0101;
															assign node41607 = (inp[14]) ? 4'b0001 : 4'b0101;
									assign node41610 = (inp[7]) ? node41738 : node41611;
										assign node41611 = (inp[15]) ? node41675 : node41612;
											assign node41612 = (inp[0]) ? node41650 : node41613;
												assign node41613 = (inp[5]) ? node41633 : node41614;
													assign node41614 = (inp[14]) ? node41620 : node41615;
														assign node41615 = (inp[4]) ? 4'b0011 : node41616;
															assign node41616 = (inp[12]) ? 4'b0111 : 4'b0011;
														assign node41620 = (inp[12]) ? node41626 : node41621;
															assign node41621 = (inp[4]) ? 4'b0111 : node41622;
																assign node41622 = (inp[9]) ? 4'b0011 : 4'b0111;
															assign node41626 = (inp[4]) ? node41630 : node41627;
																assign node41627 = (inp[9]) ? 4'b0111 : 4'b0011;
																assign node41630 = (inp[9]) ? 4'b0011 : 4'b0111;
													assign node41633 = (inp[9]) ? node41641 : node41634;
														assign node41634 = (inp[4]) ? node41638 : node41635;
															assign node41635 = (inp[12]) ? 4'b0011 : 4'b0111;
															assign node41638 = (inp[12]) ? 4'b0101 : 4'b0011;
														assign node41641 = (inp[14]) ? 4'b0101 : node41642;
															assign node41642 = (inp[4]) ? node41646 : node41643;
																assign node41643 = (inp[12]) ? 4'b0101 : 4'b0011;
																assign node41646 = (inp[12]) ? 4'b0001 : 4'b0101;
												assign node41650 = (inp[5]) ? node41662 : node41651;
													assign node41651 = (inp[9]) ? node41657 : node41652;
														assign node41652 = (inp[4]) ? node41654 : 4'b0001;
															assign node41654 = (inp[12]) ? 4'b0101 : 4'b0001;
														assign node41657 = (inp[4]) ? node41659 : 4'b0101;
															assign node41659 = (inp[12]) ? 4'b0001 : 4'b0101;
													assign node41662 = (inp[4]) ? node41668 : node41663;
														assign node41663 = (inp[12]) ? node41665 : 4'b0001;
															assign node41665 = (inp[9]) ? 4'b0111 : 4'b0001;
														assign node41668 = (inp[12]) ? node41672 : node41669;
															assign node41669 = (inp[9]) ? 4'b0111 : 4'b0001;
															assign node41672 = (inp[9]) ? 4'b0011 : 4'b0111;
											assign node41675 = (inp[0]) ? node41707 : node41676;
												assign node41676 = (inp[5]) ? node41692 : node41677;
													assign node41677 = (inp[9]) ? node41685 : node41678;
														assign node41678 = (inp[4]) ? node41682 : node41679;
															assign node41679 = (inp[12]) ? 4'b0001 : 4'b0101;
															assign node41682 = (inp[12]) ? 4'b0101 : 4'b0001;
														assign node41685 = (inp[14]) ? 4'b0001 : node41686;
															assign node41686 = (inp[4]) ? 4'b0001 : node41687;
																assign node41687 = (inp[12]) ? 4'b0101 : 4'b0001;
													assign node41692 = (inp[9]) ? node41700 : node41693;
														assign node41693 = (inp[4]) ? node41697 : node41694;
															assign node41694 = (inp[12]) ? 4'b0001 : 4'b0101;
															assign node41697 = (inp[12]) ? 4'b0111 : 4'b0001;
														assign node41700 = (inp[12]) ? node41704 : node41701;
															assign node41701 = (inp[4]) ? 4'b0111 : 4'b0001;
															assign node41704 = (inp[4]) ? 4'b0011 : 4'b0111;
												assign node41707 = (inp[9]) ? node41729 : node41708;
													assign node41708 = (inp[14]) ? node41718 : node41709;
														assign node41709 = (inp[5]) ? 4'b0111 : node41710;
															assign node41710 = (inp[12]) ? node41714 : node41711;
																assign node41711 = (inp[4]) ? 4'b0011 : 4'b0111;
																assign node41714 = (inp[4]) ? 4'b0111 : 4'b0011;
														assign node41718 = (inp[5]) ? node41724 : node41719;
															assign node41719 = (inp[12]) ? node41721 : 4'b0011;
																assign node41721 = (inp[4]) ? 4'b0111 : 4'b0011;
															assign node41724 = (inp[12]) ? 4'b0011 : node41725;
																assign node41725 = (inp[4]) ? 4'b0011 : 4'b0111;
													assign node41729 = (inp[12]) ? node41733 : node41730;
														assign node41730 = (inp[4]) ? 4'b0111 : 4'b0011;
														assign node41733 = (inp[5]) ? node41735 : 4'b0011;
															assign node41735 = (inp[4]) ? 4'b0001 : 4'b0101;
										assign node41738 = (inp[15]) ? node41804 : node41739;
											assign node41739 = (inp[0]) ? node41769 : node41740;
												assign node41740 = (inp[5]) ? node41752 : node41741;
													assign node41741 = (inp[12]) ? node41747 : node41742;
														assign node41742 = (inp[9]) ? node41744 : 4'b0010;
															assign node41744 = (inp[4]) ? 4'b0110 : 4'b0010;
														assign node41747 = (inp[4]) ? node41749 : 4'b0110;
															assign node41749 = (inp[14]) ? 4'b0010 : 4'b0110;
													assign node41752 = (inp[9]) ? node41762 : node41753;
														assign node41753 = (inp[14]) ? node41759 : node41754;
															assign node41754 = (inp[12]) ? 4'b0010 : node41755;
																assign node41755 = (inp[4]) ? 4'b0010 : 4'b0110;
															assign node41759 = (inp[12]) ? 4'b0100 : 4'b0110;
														assign node41762 = (inp[14]) ? node41764 : 4'b0100;
															assign node41764 = (inp[12]) ? node41766 : 4'b0010;
																assign node41766 = (inp[4]) ? 4'b0000 : 4'b0100;
												assign node41769 = (inp[5]) ? node41795 : node41770;
													assign node41770 = (inp[14]) ? node41786 : node41771;
														assign node41771 = (inp[9]) ? node41779 : node41772;
															assign node41772 = (inp[12]) ? node41776 : node41773;
																assign node41773 = (inp[4]) ? 4'b0000 : 4'b0100;
																assign node41776 = (inp[4]) ? 4'b0100 : 4'b0000;
															assign node41779 = (inp[4]) ? node41783 : node41780;
																assign node41780 = (inp[12]) ? 4'b0100 : 4'b0000;
																assign node41783 = (inp[12]) ? 4'b0000 : 4'b0100;
														assign node41786 = (inp[9]) ? 4'b0100 : node41787;
															assign node41787 = (inp[12]) ? node41791 : node41788;
																assign node41788 = (inp[4]) ? 4'b0000 : 4'b0100;
																assign node41791 = (inp[4]) ? 4'b0100 : 4'b0000;
													assign node41795 = (inp[4]) ? node41797 : 4'b0000;
														assign node41797 = (inp[14]) ? 4'b0010 : node41798;
															assign node41798 = (inp[9]) ? 4'b0110 : node41799;
																assign node41799 = (inp[12]) ? 4'b0110 : 4'b0000;
											assign node41804 = (inp[0]) ? node41826 : node41805;
												assign node41805 = (inp[5]) ? node41813 : node41806;
													assign node41806 = (inp[14]) ? 4'b0000 : node41807;
														assign node41807 = (inp[9]) ? 4'b0100 : node41808;
															assign node41808 = (inp[12]) ? 4'b0000 : 4'b0100;
													assign node41813 = (inp[4]) ? node41821 : node41814;
														assign node41814 = (inp[12]) ? node41818 : node41815;
															assign node41815 = (inp[9]) ? 4'b0000 : 4'b0100;
															assign node41818 = (inp[9]) ? 4'b0110 : 4'b0000;
														assign node41821 = (inp[12]) ? node41823 : 4'b0110;
															assign node41823 = (inp[9]) ? 4'b0010 : 4'b0110;
												assign node41826 = (inp[5]) ? node41840 : node41827;
													assign node41827 = (inp[9]) ? node41835 : node41828;
														assign node41828 = (inp[12]) ? node41832 : node41829;
															assign node41829 = (inp[4]) ? 4'b0010 : 4'b0110;
															assign node41832 = (inp[4]) ? 4'b0110 : 4'b0010;
														assign node41835 = (inp[12]) ? 4'b0010 : node41836;
															assign node41836 = (inp[4]) ? 4'b0110 : 4'b0010;
													assign node41840 = (inp[12]) ? node41846 : node41841;
														assign node41841 = (inp[4]) ? 4'b0010 : node41842;
															assign node41842 = (inp[9]) ? 4'b0010 : 4'b0110;
														assign node41846 = (inp[9]) ? node41848 : 4'b0010;
															assign node41848 = (inp[4]) ? 4'b0000 : 4'b0100;
								assign node41851 = (inp[5]) ? node42153 : node41852;
									assign node41852 = (inp[14]) ? node42000 : node41853;
										assign node41853 = (inp[4]) ? node41913 : node41854;
											assign node41854 = (inp[0]) ? node41886 : node41855;
												assign node41855 = (inp[15]) ? node41867 : node41856;
													assign node41856 = (inp[12]) ? node41864 : node41857;
														assign node41857 = (inp[9]) ? 4'b0011 : node41858;
															assign node41858 = (inp[7]) ? node41860 : 4'b0110;
																assign node41860 = (inp[8]) ? 4'b0110 : 4'b0111;
														assign node41864 = (inp[9]) ? 4'b0101 : 4'b0011;
													assign node41867 = (inp[9]) ? node41879 : node41868;
														assign node41868 = (inp[12]) ? node41874 : node41869;
															assign node41869 = (inp[8]) ? node41871 : 4'b0100;
																assign node41871 = (inp[7]) ? 4'b0100 : 4'b0101;
															assign node41874 = (inp[8]) ? 4'b0001 : node41875;
																assign node41875 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node41879 = (inp[7]) ? node41883 : node41880;
															assign node41880 = (inp[8]) ? 4'b0001 : 4'b0000;
															assign node41883 = (inp[8]) ? 4'b0000 : 4'b0001;
												assign node41886 = (inp[15]) ? node41900 : node41887;
													assign node41887 = (inp[9]) ? node41895 : node41888;
														assign node41888 = (inp[12]) ? node41890 : 4'b0100;
															assign node41890 = (inp[8]) ? 4'b0001 : node41891;
																assign node41891 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node41895 = (inp[12]) ? 4'b0110 : node41896;
															assign node41896 = (inp[7]) ? 4'b0001 : 4'b0000;
													assign node41900 = (inp[12]) ? node41908 : node41901;
														assign node41901 = (inp[9]) ? 4'b0011 : node41902;
															assign node41902 = (inp[8]) ? 4'b0111 : node41903;
																assign node41903 = (inp[7]) ? 4'b0111 : 4'b0110;
														assign node41908 = (inp[9]) ? 4'b0100 : node41909;
															assign node41909 = (inp[8]) ? 4'b0011 : 4'b0010;
											assign node41913 = (inp[12]) ? node41955 : node41914;
												assign node41914 = (inp[9]) ? node41942 : node41915;
													assign node41915 = (inp[8]) ? node41927 : node41916;
														assign node41916 = (inp[7]) ? node41922 : node41917;
															assign node41917 = (inp[0]) ? 4'b0010 : node41918;
																assign node41918 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node41922 = (inp[15]) ? 4'b0011 : node41923;
																assign node41923 = (inp[0]) ? 4'b0001 : 4'b0011;
														assign node41927 = (inp[7]) ? node41935 : node41928;
															assign node41928 = (inp[15]) ? node41932 : node41929;
																assign node41929 = (inp[0]) ? 4'b0001 : 4'b0011;
																assign node41932 = (inp[0]) ? 4'b0011 : 4'b0001;
															assign node41935 = (inp[0]) ? node41939 : node41936;
																assign node41936 = (inp[15]) ? 4'b0000 : 4'b0010;
																assign node41939 = (inp[15]) ? 4'b0010 : 4'b0000;
													assign node41942 = (inp[8]) ? node41950 : node41943;
														assign node41943 = (inp[7]) ? node41945 : 4'b0110;
															assign node41945 = (inp[15]) ? 4'b0111 : node41946;
																assign node41946 = (inp[0]) ? 4'b0111 : 4'b0101;
														assign node41950 = (inp[7]) ? 4'b0110 : node41951;
															assign node41951 = (inp[15]) ? 4'b0101 : 4'b0111;
												assign node41955 = (inp[9]) ? node41977 : node41956;
													assign node41956 = (inp[7]) ? node41964 : node41957;
														assign node41957 = (inp[8]) ? node41959 : 4'b0110;
															assign node41959 = (inp[0]) ? node41961 : 4'b0111;
																assign node41961 = (inp[15]) ? 4'b0101 : 4'b0111;
														assign node41964 = (inp[8]) ? node41972 : node41965;
															assign node41965 = (inp[15]) ? node41969 : node41966;
																assign node41966 = (inp[0]) ? 4'b0111 : 4'b0101;
																assign node41969 = (inp[0]) ? 4'b0101 : 4'b0111;
															assign node41972 = (inp[0]) ? 4'b0110 : node41973;
																assign node41973 = (inp[15]) ? 4'b0110 : 4'b0100;
													assign node41977 = (inp[15]) ? node41991 : node41978;
														assign node41978 = (inp[0]) ? node41986 : node41979;
															assign node41979 = (inp[7]) ? node41983 : node41980;
																assign node41980 = (inp[8]) ? 4'b0001 : 4'b0000;
																assign node41983 = (inp[8]) ? 4'b0000 : 4'b0001;
															assign node41986 = (inp[7]) ? node41988 : 4'b0010;
																assign node41988 = (inp[8]) ? 4'b0010 : 4'b0011;
														assign node41991 = (inp[0]) ? node41997 : node41992;
															assign node41992 = (inp[7]) ? node41994 : 4'b0011;
																assign node41994 = (inp[8]) ? 4'b0010 : 4'b0011;
															assign node41997 = (inp[7]) ? 4'b0001 : 4'b0000;
										assign node42000 = (inp[8]) ? node42070 : node42001;
											assign node42001 = (inp[7]) ? node42027 : node42002;
												assign node42002 = (inp[4]) ? node42012 : node42003;
													assign node42003 = (inp[9]) ? node42007 : node42004;
														assign node42004 = (inp[0]) ? 4'b0000 : 4'b0010;
														assign node42007 = (inp[12]) ? 4'b0100 : node42008;
															assign node42008 = (inp[0]) ? 4'b0010 : 4'b0000;
													assign node42012 = (inp[9]) ? node42020 : node42013;
														assign node42013 = (inp[12]) ? node42015 : 4'b0010;
															assign node42015 = (inp[0]) ? 4'b0110 : node42016;
																assign node42016 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node42020 = (inp[12]) ? 4'b0010 : node42021;
															assign node42021 = (inp[0]) ? node42023 : 4'b0110;
																assign node42023 = (inp[15]) ? 4'b0100 : 4'b0110;
												assign node42027 = (inp[9]) ? node42051 : node42028;
													assign node42028 = (inp[15]) ? node42038 : node42029;
														assign node42029 = (inp[0]) ? 4'b0101 : node42030;
															assign node42030 = (inp[12]) ? node42034 : node42031;
																assign node42031 = (inp[4]) ? 4'b0011 : 4'b0111;
																assign node42034 = (inp[4]) ? 4'b0101 : 4'b0011;
														assign node42038 = (inp[0]) ? node42046 : node42039;
															assign node42039 = (inp[4]) ? node42043 : node42040;
																assign node42040 = (inp[12]) ? 4'b0001 : 4'b0101;
																assign node42043 = (inp[12]) ? 4'b0111 : 4'b0001;
															assign node42046 = (inp[12]) ? node42048 : 4'b0011;
																assign node42048 = (inp[4]) ? 4'b0101 : 4'b0011;
													assign node42051 = (inp[15]) ? node42063 : node42052;
														assign node42052 = (inp[12]) ? node42060 : node42053;
															assign node42053 = (inp[4]) ? node42057 : node42054;
																assign node42054 = (inp[0]) ? 4'b0001 : 4'b0011;
																assign node42057 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node42060 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node42063 = (inp[0]) ? 4'b0101 : node42064;
															assign node42064 = (inp[4]) ? node42066 : 4'b0111;
																assign node42066 = (inp[12]) ? 4'b0011 : 4'b0111;
											assign node42070 = (inp[7]) ? node42106 : node42071;
												assign node42071 = (inp[9]) ? node42089 : node42072;
													assign node42072 = (inp[12]) ? node42080 : node42073;
														assign node42073 = (inp[4]) ? 4'b0011 : node42074;
															assign node42074 = (inp[0]) ? 4'b0111 : node42075;
																assign node42075 = (inp[15]) ? 4'b0101 : 4'b0111;
														assign node42080 = (inp[4]) ? node42082 : 4'b0011;
															assign node42082 = (inp[15]) ? node42086 : node42083;
																assign node42083 = (inp[0]) ? 4'b0111 : 4'b0101;
																assign node42086 = (inp[0]) ? 4'b0101 : 4'b0111;
													assign node42089 = (inp[12]) ? node42099 : node42090;
														assign node42090 = (inp[4]) ? node42092 : 4'b0001;
															assign node42092 = (inp[15]) ? node42096 : node42093;
																assign node42093 = (inp[0]) ? 4'b0111 : 4'b0101;
																assign node42096 = (inp[0]) ? 4'b0101 : 4'b0111;
														assign node42099 = (inp[4]) ? node42101 : 4'b0111;
															assign node42101 = (inp[0]) ? node42103 : 4'b0011;
																assign node42103 = (inp[15]) ? 4'b0001 : 4'b0011;
												assign node42106 = (inp[4]) ? node42124 : node42107;
													assign node42107 = (inp[15]) ? node42115 : node42108;
														assign node42108 = (inp[0]) ? node42112 : node42109;
															assign node42109 = (inp[9]) ? 4'b0010 : 4'b0110;
															assign node42112 = (inp[9]) ? 4'b0110 : 4'b0000;
														assign node42115 = (inp[0]) ? node42119 : node42116;
															assign node42116 = (inp[9]) ? 4'b0110 : 4'b0100;
															assign node42119 = (inp[9]) ? 4'b0100 : node42120;
																assign node42120 = (inp[12]) ? 4'b0010 : 4'b0110;
													assign node42124 = (inp[15]) ? node42140 : node42125;
														assign node42125 = (inp[0]) ? node42133 : node42126;
															assign node42126 = (inp[12]) ? node42130 : node42127;
																assign node42127 = (inp[9]) ? 4'b0100 : 4'b0010;
																assign node42130 = (inp[9]) ? 4'b0000 : 4'b0100;
															assign node42133 = (inp[9]) ? node42137 : node42134;
																assign node42134 = (inp[12]) ? 4'b0110 : 4'b0000;
																assign node42137 = (inp[12]) ? 4'b0010 : 4'b0110;
														assign node42140 = (inp[0]) ? node42146 : node42141;
															assign node42141 = (inp[12]) ? node42143 : 4'b0110;
																assign node42143 = (inp[9]) ? 4'b0010 : 4'b0110;
															assign node42146 = (inp[12]) ? node42150 : node42147;
																assign node42147 = (inp[9]) ? 4'b0100 : 4'b0010;
																assign node42150 = (inp[9]) ? 4'b0000 : 4'b0100;
									assign node42153 = (inp[12]) ? node42287 : node42154;
										assign node42154 = (inp[0]) ? node42216 : node42155;
											assign node42155 = (inp[15]) ? node42173 : node42156;
												assign node42156 = (inp[4]) ? node42164 : node42157;
													assign node42157 = (inp[8]) ? node42161 : node42158;
														assign node42158 = (inp[7]) ? 4'b0101 : 4'b0100;
														assign node42161 = (inp[7]) ? 4'b0100 : 4'b0101;
													assign node42164 = (inp[9]) ? node42166 : 4'b0001;
														assign node42166 = (inp[14]) ? 4'b0101 : node42167;
															assign node42167 = (inp[8]) ? 4'b0100 : node42168;
																assign node42168 = (inp[7]) ? 4'b0101 : 4'b0100;
												assign node42173 = (inp[14]) ? node42193 : node42174;
													assign node42174 = (inp[4]) ? node42186 : node42175;
														assign node42175 = (inp[9]) ? node42183 : node42176;
															assign node42176 = (inp[7]) ? node42180 : node42177;
																assign node42177 = (inp[8]) ? 4'b0111 : 4'b0110;
																assign node42180 = (inp[8]) ? 4'b0110 : 4'b0111;
															assign node42183 = (inp[8]) ? 4'b0010 : 4'b0011;
														assign node42186 = (inp[9]) ? 4'b0110 : node42187;
															assign node42187 = (inp[7]) ? 4'b0010 : node42188;
																assign node42188 = (inp[8]) ? 4'b0011 : 4'b0010;
													assign node42193 = (inp[9]) ? node42203 : node42194;
														assign node42194 = (inp[4]) ? 4'b0011 : node42195;
															assign node42195 = (inp[7]) ? node42199 : node42196;
																assign node42196 = (inp[8]) ? 4'b0111 : 4'b0110;
																assign node42199 = (inp[8]) ? 4'b0110 : 4'b0111;
														assign node42203 = (inp[4]) ? node42209 : node42204;
															assign node42204 = (inp[8]) ? 4'b0011 : node42205;
																assign node42205 = (inp[7]) ? 4'b0011 : 4'b0010;
															assign node42209 = (inp[8]) ? node42213 : node42210;
																assign node42210 = (inp[7]) ? 4'b0111 : 4'b0110;
																assign node42213 = (inp[7]) ? 4'b0110 : 4'b0111;
											assign node42216 = (inp[15]) ? node42254 : node42217;
												assign node42217 = (inp[14]) ? node42241 : node42218;
													assign node42218 = (inp[7]) ? node42228 : node42219;
														assign node42219 = (inp[8]) ? node42223 : node42220;
															assign node42220 = (inp[9]) ? 4'b0110 : 4'b0010;
															assign node42223 = (inp[4]) ? node42225 : 4'b0011;
																assign node42225 = (inp[9]) ? 4'b0111 : 4'b0011;
														assign node42228 = (inp[8]) ? node42236 : node42229;
															assign node42229 = (inp[9]) ? node42233 : node42230;
																assign node42230 = (inp[4]) ? 4'b0011 : 4'b0111;
																assign node42233 = (inp[4]) ? 4'b0111 : 4'b0011;
															assign node42236 = (inp[9]) ? node42238 : 4'b0110;
																assign node42238 = (inp[4]) ? 4'b0110 : 4'b0010;
													assign node42241 = (inp[9]) ? node42249 : node42242;
														assign node42242 = (inp[4]) ? node42244 : 4'b0110;
															assign node42244 = (inp[7]) ? 4'b0010 : node42245;
																assign node42245 = (inp[8]) ? 4'b0011 : 4'b0010;
														assign node42249 = (inp[7]) ? node42251 : 4'b0010;
															assign node42251 = (inp[8]) ? 4'b0110 : 4'b0111;
												assign node42254 = (inp[14]) ? node42270 : node42255;
													assign node42255 = (inp[9]) ? node42265 : node42256;
														assign node42256 = (inp[4]) ? node42262 : node42257;
															assign node42257 = (inp[8]) ? 4'b0101 : node42258;
																assign node42258 = (inp[7]) ? 4'b0101 : 4'b0100;
															assign node42262 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node42265 = (inp[7]) ? node42267 : 4'b0101;
															assign node42267 = (inp[8]) ? 4'b0100 : 4'b0101;
													assign node42270 = (inp[4]) ? node42284 : node42271;
														assign node42271 = (inp[9]) ? node42279 : node42272;
															assign node42272 = (inp[8]) ? node42276 : node42273;
																assign node42273 = (inp[7]) ? 4'b0101 : 4'b0100;
																assign node42276 = (inp[7]) ? 4'b0100 : 4'b0101;
															assign node42279 = (inp[7]) ? 4'b0000 : node42280;
																assign node42280 = (inp[8]) ? 4'b0001 : 4'b0000;
														assign node42284 = (inp[9]) ? 4'b0100 : 4'b0000;
										assign node42287 = (inp[7]) ? node42351 : node42288;
											assign node42288 = (inp[8]) ? node42314 : node42289;
												assign node42289 = (inp[9]) ? node42305 : node42290;
													assign node42290 = (inp[4]) ? node42298 : node42291;
														assign node42291 = (inp[0]) ? node42295 : node42292;
															assign node42292 = (inp[15]) ? 4'b0010 : 4'b0000;
															assign node42295 = (inp[15]) ? 4'b0000 : 4'b0010;
														assign node42298 = (inp[15]) ? node42302 : node42299;
															assign node42299 = (inp[0]) ? 4'b0110 : 4'b0100;
															assign node42302 = (inp[14]) ? 4'b0100 : 4'b0110;
													assign node42305 = (inp[4]) ? node42311 : node42306;
														assign node42306 = (inp[15]) ? node42308 : 4'b0110;
															assign node42308 = (inp[0]) ? 4'b0100 : 4'b0110;
														assign node42311 = (inp[0]) ? 4'b0010 : 4'b0000;
												assign node42314 = (inp[14]) ? node42328 : node42315;
													assign node42315 = (inp[15]) ? node42319 : node42316;
														assign node42316 = (inp[0]) ? 4'b0111 : 4'b0101;
														assign node42319 = (inp[0]) ? node42323 : node42320;
															assign node42320 = (inp[9]) ? 4'b0111 : 4'b0011;
															assign node42323 = (inp[4]) ? 4'b0001 : node42324;
																assign node42324 = (inp[9]) ? 4'b0101 : 4'b0001;
													assign node42328 = (inp[0]) ? node42342 : node42329;
														assign node42329 = (inp[15]) ? node42335 : node42330;
															assign node42330 = (inp[9]) ? 4'b0001 : node42331;
																assign node42331 = (inp[4]) ? 4'b0101 : 4'b0001;
															assign node42335 = (inp[9]) ? node42339 : node42336;
																assign node42336 = (inp[4]) ? 4'b0111 : 4'b0011;
																assign node42339 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node42342 = (inp[15]) ? 4'b0101 : node42343;
															assign node42343 = (inp[9]) ? node42347 : node42344;
																assign node42344 = (inp[4]) ? 4'b0111 : 4'b0011;
																assign node42347 = (inp[4]) ? 4'b0011 : 4'b0111;
											assign node42351 = (inp[8]) ? node42371 : node42352;
												assign node42352 = (inp[4]) ? node42360 : node42353;
													assign node42353 = (inp[9]) ? node42355 : 4'b0001;
														assign node42355 = (inp[0]) ? node42357 : 4'b0101;
															assign node42357 = (inp[15]) ? 4'b0101 : 4'b0111;
													assign node42360 = (inp[9]) ? node42366 : node42361;
														assign node42361 = (inp[15]) ? node42363 : 4'b0101;
															assign node42363 = (inp[0]) ? 4'b0101 : 4'b0111;
														assign node42366 = (inp[0]) ? 4'b0011 : node42367;
															assign node42367 = (inp[15]) ? 4'b0011 : 4'b0001;
												assign node42371 = (inp[15]) ? node42385 : node42372;
													assign node42372 = (inp[0]) ? node42380 : node42373;
														assign node42373 = (inp[9]) ? node42377 : node42374;
															assign node42374 = (inp[4]) ? 4'b0100 : 4'b0000;
															assign node42377 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node42380 = (inp[4]) ? node42382 : 4'b0110;
															assign node42382 = (inp[9]) ? 4'b0010 : 4'b0110;
													assign node42385 = (inp[0]) ? node42397 : node42386;
														assign node42386 = (inp[14]) ? node42392 : node42387;
															assign node42387 = (inp[9]) ? node42389 : 4'b0010;
																assign node42389 = (inp[4]) ? 4'b0010 : 4'b0110;
															assign node42392 = (inp[9]) ? 4'b0110 : node42393;
																assign node42393 = (inp[4]) ? 4'b0110 : 4'b0010;
														assign node42397 = (inp[14]) ? 4'b0000 : node42398;
															assign node42398 = (inp[9]) ? node42402 : node42399;
																assign node42399 = (inp[4]) ? 4'b0100 : 4'b0000;
																assign node42402 = (inp[4]) ? 4'b0000 : 4'b0100;
						assign node42406 = (inp[7]) ? node43276 : node42407;
							assign node42407 = (inp[8]) ? node42935 : node42408;
								assign node42408 = (inp[2]) ? node42670 : node42409;
									assign node42409 = (inp[14]) ? node42543 : node42410;
										assign node42410 = (inp[15]) ? node42488 : node42411;
											assign node42411 = (inp[0]) ? node42455 : node42412;
												assign node42412 = (inp[3]) ? node42432 : node42413;
													assign node42413 = (inp[5]) ? node42417 : node42414;
														assign node42414 = (inp[12]) ? 4'b0011 : 4'b0111;
														assign node42417 = (inp[9]) ? node42425 : node42418;
															assign node42418 = (inp[12]) ? node42422 : node42419;
																assign node42419 = (inp[4]) ? 4'b0011 : 4'b0111;
																assign node42422 = (inp[4]) ? 4'b0101 : 4'b0011;
															assign node42425 = (inp[4]) ? node42429 : node42426;
																assign node42426 = (inp[12]) ? 4'b0101 : 4'b0011;
																assign node42429 = (inp[12]) ? 4'b0001 : 4'b0101;
													assign node42432 = (inp[5]) ? node42442 : node42433;
														assign node42433 = (inp[12]) ? node42435 : 4'b0011;
															assign node42435 = (inp[4]) ? node42439 : node42436;
																assign node42436 = (inp[9]) ? 4'b0101 : 4'b0011;
																assign node42439 = (inp[9]) ? 4'b0001 : 4'b0101;
														assign node42442 = (inp[9]) ? node42450 : node42443;
															assign node42443 = (inp[12]) ? node42447 : node42444;
																assign node42444 = (inp[4]) ? 4'b0001 : 4'b0101;
																assign node42447 = (inp[4]) ? 4'b0101 : 4'b0001;
															assign node42450 = (inp[4]) ? 4'b0101 : node42451;
																assign node42451 = (inp[12]) ? 4'b0101 : 4'b0001;
												assign node42455 = (inp[3]) ? node42475 : node42456;
													assign node42456 = (inp[12]) ? node42462 : node42457;
														assign node42457 = (inp[4]) ? 4'b0001 : node42458;
															assign node42458 = (inp[9]) ? 4'b0001 : 4'b0101;
														assign node42462 = (inp[5]) ? node42468 : node42463;
															assign node42463 = (inp[9]) ? 4'b0101 : node42464;
																assign node42464 = (inp[4]) ? 4'b0101 : 4'b0001;
															assign node42468 = (inp[9]) ? node42472 : node42469;
																assign node42469 = (inp[4]) ? 4'b0111 : 4'b0001;
																assign node42472 = (inp[4]) ? 4'b0011 : 4'b0111;
													assign node42475 = (inp[4]) ? node42483 : node42476;
														assign node42476 = (inp[9]) ? 4'b0111 : node42477;
															assign node42477 = (inp[12]) ? node42479 : 4'b0111;
																assign node42479 = (inp[5]) ? 4'b0011 : 4'b0001;
														assign node42483 = (inp[9]) ? 4'b0011 : node42484;
															assign node42484 = (inp[12]) ? 4'b0111 : 4'b0011;
											assign node42488 = (inp[12]) ? node42516 : node42489;
												assign node42489 = (inp[4]) ? node42507 : node42490;
													assign node42490 = (inp[9]) ? node42500 : node42491;
														assign node42491 = (inp[5]) ? node42493 : 4'b0111;
															assign node42493 = (inp[3]) ? node42497 : node42494;
																assign node42494 = (inp[0]) ? 4'b0111 : 4'b0101;
																assign node42497 = (inp[0]) ? 4'b0101 : 4'b0111;
														assign node42500 = (inp[0]) ? node42502 : 4'b0011;
															assign node42502 = (inp[5]) ? node42504 : 4'b0011;
																assign node42504 = (inp[3]) ? 4'b0001 : 4'b0011;
													assign node42507 = (inp[9]) ? 4'b0101 : node42508;
														assign node42508 = (inp[0]) ? node42510 : 4'b0001;
															assign node42510 = (inp[3]) ? node42512 : 4'b0011;
																assign node42512 = (inp[5]) ? 4'b0001 : 4'b0011;
												assign node42516 = (inp[5]) ? node42538 : node42517;
													assign node42517 = (inp[9]) ? node42529 : node42518;
														assign node42518 = (inp[4]) ? node42522 : node42519;
															assign node42519 = (inp[0]) ? 4'b0011 : 4'b0001;
															assign node42522 = (inp[3]) ? node42526 : node42523;
																assign node42523 = (inp[0]) ? 4'b0111 : 4'b0101;
																assign node42526 = (inp[0]) ? 4'b0101 : 4'b0111;
														assign node42529 = (inp[4]) ? 4'b0011 : node42530;
															assign node42530 = (inp[3]) ? node42534 : node42531;
																assign node42531 = (inp[0]) ? 4'b0111 : 4'b0101;
																assign node42534 = (inp[0]) ? 4'b0101 : 4'b0111;
													assign node42538 = (inp[0]) ? node42540 : 4'b0111;
														assign node42540 = (inp[4]) ? 4'b0001 : 4'b0101;
										assign node42543 = (inp[0]) ? node42597 : node42544;
											assign node42544 = (inp[9]) ? node42564 : node42545;
												assign node42545 = (inp[4]) ? node42557 : node42546;
													assign node42546 = (inp[12]) ? node42550 : node42547;
														assign node42547 = (inp[15]) ? 4'b0100 : 4'b0110;
														assign node42550 = (inp[15]) ? 4'b0000 : node42551;
															assign node42551 = (inp[5]) ? node42553 : 4'b0010;
																assign node42553 = (inp[3]) ? 4'b0000 : 4'b0010;
													assign node42557 = (inp[12]) ? node42559 : 4'b0000;
														assign node42559 = (inp[15]) ? node42561 : 4'b0100;
															assign node42561 = (inp[5]) ? 4'b0110 : 4'b0100;
												assign node42564 = (inp[15]) ? node42578 : node42565;
													assign node42565 = (inp[5]) ? node42573 : node42566;
														assign node42566 = (inp[3]) ? node42568 : 4'b0110;
															assign node42568 = (inp[12]) ? node42570 : 4'b0010;
																assign node42570 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node42573 = (inp[12]) ? node42575 : 4'b0100;
															assign node42575 = (inp[4]) ? 4'b0000 : 4'b0100;
													assign node42578 = (inp[3]) ? node42590 : node42579;
														assign node42579 = (inp[5]) ? node42585 : node42580;
															assign node42580 = (inp[12]) ? node42582 : 4'b0100;
																assign node42582 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node42585 = (inp[4]) ? node42587 : 4'b0000;
																assign node42587 = (inp[12]) ? 4'b0010 : 4'b0110;
														assign node42590 = (inp[4]) ? node42594 : node42591;
															assign node42591 = (inp[12]) ? 4'b0110 : 4'b0010;
															assign node42594 = (inp[12]) ? 4'b0010 : 4'b0110;
											assign node42597 = (inp[15]) ? node42635 : node42598;
												assign node42598 = (inp[5]) ? node42618 : node42599;
													assign node42599 = (inp[3]) ? node42603 : node42600;
														assign node42600 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node42603 = (inp[12]) ? node42611 : node42604;
															assign node42604 = (inp[4]) ? node42608 : node42605;
																assign node42605 = (inp[9]) ? 4'b0000 : 4'b0100;
																assign node42608 = (inp[9]) ? 4'b0110 : 4'b0000;
															assign node42611 = (inp[9]) ? node42615 : node42612;
																assign node42612 = (inp[4]) ? 4'b0110 : 4'b0000;
																assign node42615 = (inp[4]) ? 4'b0010 : 4'b0110;
													assign node42618 = (inp[3]) ? node42624 : node42619;
														assign node42619 = (inp[12]) ? node42621 : 4'b0110;
															assign node42621 = (inp[9]) ? 4'b0010 : 4'b0110;
														assign node42624 = (inp[12]) ? node42630 : node42625;
															assign node42625 = (inp[4]) ? node42627 : 4'b0010;
																assign node42627 = (inp[9]) ? 4'b0110 : 4'b0010;
															assign node42630 = (inp[9]) ? node42632 : 4'b0110;
																assign node42632 = (inp[4]) ? 4'b0010 : 4'b0110;
												assign node42635 = (inp[3]) ? node42653 : node42636;
													assign node42636 = (inp[5]) ? node42644 : node42637;
														assign node42637 = (inp[4]) ? node42639 : 4'b0110;
															assign node42639 = (inp[9]) ? 4'b0010 : node42640;
																assign node42640 = (inp[12]) ? 4'b0110 : 4'b0010;
														assign node42644 = (inp[12]) ? 4'b0100 : node42645;
															assign node42645 = (inp[4]) ? node42649 : node42646;
																assign node42646 = (inp[9]) ? 4'b0010 : 4'b0110;
																assign node42649 = (inp[9]) ? 4'b0100 : 4'b0010;
													assign node42653 = (inp[4]) ? node42665 : node42654;
														assign node42654 = (inp[5]) ? node42660 : node42655;
															assign node42655 = (inp[9]) ? node42657 : 4'b0010;
																assign node42657 = (inp[12]) ? 4'b0100 : 4'b0010;
															assign node42660 = (inp[12]) ? 4'b0100 : node42661;
																assign node42661 = (inp[9]) ? 4'b0000 : 4'b0100;
														assign node42665 = (inp[12]) ? node42667 : 4'b0100;
															assign node42667 = (inp[9]) ? 4'b0000 : 4'b0100;
									assign node42670 = (inp[4]) ? node42796 : node42671;
										assign node42671 = (inp[14]) ? node42735 : node42672;
											assign node42672 = (inp[15]) ? node42704 : node42673;
												assign node42673 = (inp[12]) ? node42689 : node42674;
													assign node42674 = (inp[9]) ? node42680 : node42675;
														assign node42675 = (inp[0]) ? node42677 : 4'b0110;
															assign node42677 = (inp[3]) ? 4'b0110 : 4'b0100;
														assign node42680 = (inp[0]) ? node42686 : node42681;
															assign node42681 = (inp[3]) ? node42683 : 4'b0010;
																assign node42683 = (inp[5]) ? 4'b0000 : 4'b0010;
															assign node42686 = (inp[3]) ? 4'b0010 : 4'b0000;
													assign node42689 = (inp[9]) ? node42693 : node42690;
														assign node42690 = (inp[0]) ? 4'b0000 : 4'b0010;
														assign node42693 = (inp[0]) ? node42699 : node42694;
															assign node42694 = (inp[5]) ? 4'b0100 : node42695;
																assign node42695 = (inp[3]) ? 4'b0100 : 4'b0110;
															assign node42699 = (inp[3]) ? 4'b0110 : node42700;
																assign node42700 = (inp[5]) ? 4'b0110 : 4'b0100;
												assign node42704 = (inp[0]) ? node42722 : node42705;
													assign node42705 = (inp[3]) ? node42717 : node42706;
														assign node42706 = (inp[5]) ? node42714 : node42707;
															assign node42707 = (inp[9]) ? node42711 : node42708;
																assign node42708 = (inp[12]) ? 4'b0000 : 4'b0100;
																assign node42711 = (inp[12]) ? 4'b0100 : 4'b0000;
															assign node42714 = (inp[12]) ? 4'b0110 : 4'b0000;
														assign node42717 = (inp[5]) ? 4'b0110 : node42718;
															assign node42718 = (inp[9]) ? 4'b0110 : 4'b0100;
													assign node42722 = (inp[9]) ? node42730 : node42723;
														assign node42723 = (inp[12]) ? 4'b0010 : node42724;
															assign node42724 = (inp[5]) ? node42726 : 4'b0110;
																assign node42726 = (inp[3]) ? 4'b0100 : 4'b0110;
														assign node42730 = (inp[3]) ? 4'b0100 : node42731;
															assign node42731 = (inp[5]) ? 4'b0100 : 4'b0110;
											assign node42735 = (inp[12]) ? node42771 : node42736;
												assign node42736 = (inp[9]) ? node42752 : node42737;
													assign node42737 = (inp[5]) ? node42745 : node42738;
														assign node42738 = (inp[0]) ? node42742 : node42739;
															assign node42739 = (inp[15]) ? 4'b0100 : 4'b0110;
															assign node42742 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node42745 = (inp[0]) ? 4'b0110 : node42746;
															assign node42746 = (inp[3]) ? 4'b0110 : node42747;
																assign node42747 = (inp[15]) ? 4'b0100 : 4'b0110;
													assign node42752 = (inp[3]) ? node42758 : node42753;
														assign node42753 = (inp[0]) ? 4'b0010 : node42754;
															assign node42754 = (inp[15]) ? 4'b0000 : 4'b0010;
														assign node42758 = (inp[0]) ? node42764 : node42759;
															assign node42759 = (inp[15]) ? node42761 : 4'b0010;
																assign node42761 = (inp[5]) ? 4'b0010 : 4'b0000;
															assign node42764 = (inp[15]) ? node42768 : node42765;
																assign node42765 = (inp[5]) ? 4'b0010 : 4'b0000;
																assign node42768 = (inp[5]) ? 4'b0000 : 4'b0010;
												assign node42771 = (inp[9]) ? node42789 : node42772;
													assign node42772 = (inp[15]) ? node42784 : node42773;
														assign node42773 = (inp[0]) ? node42779 : node42774;
															assign node42774 = (inp[5]) ? node42776 : 4'b0010;
																assign node42776 = (inp[3]) ? 4'b0000 : 4'b0010;
															assign node42779 = (inp[3]) ? node42781 : 4'b0000;
																assign node42781 = (inp[5]) ? 4'b0010 : 4'b0000;
														assign node42784 = (inp[0]) ? 4'b0010 : node42785;
															assign node42785 = (inp[3]) ? 4'b0010 : 4'b0000;
													assign node42789 = (inp[0]) ? 4'b0110 : node42790;
														assign node42790 = (inp[15]) ? 4'b0110 : node42791;
															assign node42791 = (inp[5]) ? 4'b0100 : 4'b0110;
										assign node42796 = (inp[5]) ? node42874 : node42797;
											assign node42797 = (inp[0]) ? node42835 : node42798;
												assign node42798 = (inp[15]) ? node42822 : node42799;
													assign node42799 = (inp[3]) ? node42815 : node42800;
														assign node42800 = (inp[14]) ? node42808 : node42801;
															assign node42801 = (inp[9]) ? node42805 : node42802;
																assign node42802 = (inp[12]) ? 4'b0110 : 4'b0010;
																assign node42805 = (inp[12]) ? 4'b0010 : 4'b0110;
															assign node42808 = (inp[9]) ? node42812 : node42809;
																assign node42809 = (inp[12]) ? 4'b0110 : 4'b0010;
																assign node42812 = (inp[12]) ? 4'b0010 : 4'b0110;
														assign node42815 = (inp[9]) ? node42819 : node42816;
															assign node42816 = (inp[12]) ? 4'b0100 : 4'b0010;
															assign node42819 = (inp[12]) ? 4'b0000 : 4'b0100;
													assign node42822 = (inp[3]) ? node42830 : node42823;
														assign node42823 = (inp[9]) ? node42827 : node42824;
															assign node42824 = (inp[12]) ? 4'b0100 : 4'b0000;
															assign node42827 = (inp[12]) ? 4'b0000 : 4'b0100;
														assign node42830 = (inp[12]) ? node42832 : 4'b0000;
															assign node42832 = (inp[9]) ? 4'b0010 : 4'b0110;
												assign node42835 = (inp[15]) ? node42855 : node42836;
													assign node42836 = (inp[3]) ? node42846 : node42837;
														assign node42837 = (inp[14]) ? node42839 : 4'b0100;
															assign node42839 = (inp[9]) ? node42843 : node42840;
																assign node42840 = (inp[12]) ? 4'b0100 : 4'b0000;
																assign node42843 = (inp[12]) ? 4'b0000 : 4'b0100;
														assign node42846 = (inp[14]) ? node42850 : node42847;
															assign node42847 = (inp[12]) ? 4'b0010 : 4'b0000;
															assign node42850 = (inp[12]) ? node42852 : 4'b0110;
																assign node42852 = (inp[9]) ? 4'b0010 : 4'b0110;
													assign node42855 = (inp[3]) ? node42869 : node42856;
														assign node42856 = (inp[14]) ? node42862 : node42857;
															assign node42857 = (inp[9]) ? 4'b0010 : node42858;
																assign node42858 = (inp[12]) ? 4'b0110 : 4'b0010;
															assign node42862 = (inp[12]) ? node42866 : node42863;
																assign node42863 = (inp[9]) ? 4'b0110 : 4'b0010;
																assign node42866 = (inp[9]) ? 4'b0010 : 4'b0110;
														assign node42869 = (inp[12]) ? 4'b0100 : node42870;
															assign node42870 = (inp[9]) ? 4'b0100 : 4'b0010;
											assign node42874 = (inp[9]) ? node42906 : node42875;
												assign node42875 = (inp[12]) ? node42887 : node42876;
													assign node42876 = (inp[14]) ? node42884 : node42877;
														assign node42877 = (inp[15]) ? node42879 : 4'b0000;
															assign node42879 = (inp[0]) ? 4'b0010 : node42880;
																assign node42880 = (inp[3]) ? 4'b0010 : 4'b0000;
														assign node42884 = (inp[15]) ? 4'b0000 : 4'b0010;
													assign node42887 = (inp[14]) ? node42899 : node42888;
														assign node42888 = (inp[3]) ? node42894 : node42889;
															assign node42889 = (inp[15]) ? node42891 : 4'b0110;
																assign node42891 = (inp[0]) ? 4'b0100 : 4'b0110;
															assign node42894 = (inp[15]) ? node42896 : 4'b0100;
																assign node42896 = (inp[0]) ? 4'b0100 : 4'b0110;
														assign node42899 = (inp[3]) ? node42901 : 4'b0100;
															assign node42901 = (inp[15]) ? node42903 : 4'b0100;
																assign node42903 = (inp[0]) ? 4'b0100 : 4'b0110;
												assign node42906 = (inp[12]) ? node42914 : node42907;
													assign node42907 = (inp[15]) ? node42911 : node42908;
														assign node42908 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node42911 = (inp[0]) ? 4'b0100 : 4'b0110;
													assign node42914 = (inp[3]) ? node42922 : node42915;
														assign node42915 = (inp[15]) ? node42919 : node42916;
															assign node42916 = (inp[0]) ? 4'b0010 : 4'b0000;
															assign node42919 = (inp[0]) ? 4'b0000 : 4'b0010;
														assign node42922 = (inp[14]) ? node42928 : node42923;
															assign node42923 = (inp[15]) ? node42925 : 4'b0010;
																assign node42925 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node42928 = (inp[0]) ? node42932 : node42929;
																assign node42929 = (inp[15]) ? 4'b0010 : 4'b0000;
																assign node42932 = (inp[15]) ? 4'b0000 : 4'b0010;
								assign node42935 = (inp[2]) ? node43165 : node42936;
									assign node42936 = (inp[14]) ? node43076 : node42937;
										assign node42937 = (inp[12]) ? node43005 : node42938;
											assign node42938 = (inp[3]) ? node42964 : node42939;
												assign node42939 = (inp[15]) ? node42949 : node42940;
													assign node42940 = (inp[0]) ? node42946 : node42941;
														assign node42941 = (inp[4]) ? node42943 : 4'b0110;
															assign node42943 = (inp[9]) ? 4'b0110 : 4'b0010;
														assign node42946 = (inp[9]) ? 4'b0000 : 4'b0100;
													assign node42949 = (inp[0]) ? node42959 : node42950;
														assign node42950 = (inp[5]) ? 4'b0000 : node42951;
															assign node42951 = (inp[9]) ? node42955 : node42952;
																assign node42952 = (inp[4]) ? 4'b0000 : 4'b0100;
																assign node42955 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node42959 = (inp[4]) ? node42961 : 4'b0010;
															assign node42961 = (inp[5]) ? 4'b0100 : 4'b0110;
												assign node42964 = (inp[0]) ? node42986 : node42965;
													assign node42965 = (inp[15]) ? node42977 : node42966;
														assign node42966 = (inp[5]) ? node42970 : node42967;
															assign node42967 = (inp[4]) ? 4'b0100 : 4'b0110;
															assign node42970 = (inp[4]) ? node42974 : node42971;
																assign node42971 = (inp[9]) ? 4'b0000 : 4'b0100;
																assign node42974 = (inp[9]) ? 4'b0100 : 4'b0000;
														assign node42977 = (inp[5]) ? 4'b0110 : node42978;
															assign node42978 = (inp[9]) ? node42982 : node42979;
																assign node42979 = (inp[4]) ? 4'b0000 : 4'b0100;
																assign node42982 = (inp[4]) ? 4'b0110 : 4'b0000;
													assign node42986 = (inp[5]) ? node43000 : node42987;
														assign node42987 = (inp[15]) ? node42995 : node42988;
															assign node42988 = (inp[9]) ? node42992 : node42989;
																assign node42989 = (inp[4]) ? 4'b0000 : 4'b0100;
																assign node42992 = (inp[4]) ? 4'b0110 : 4'b0000;
															assign node42995 = (inp[9]) ? 4'b0010 : node42996;
																assign node42996 = (inp[4]) ? 4'b0010 : 4'b0110;
														assign node43000 = (inp[15]) ? 4'b0100 : node43001;
															assign node43001 = (inp[4]) ? 4'b0110 : 4'b0010;
											assign node43005 = (inp[4]) ? node43041 : node43006;
												assign node43006 = (inp[9]) ? node43028 : node43007;
													assign node43007 = (inp[0]) ? node43019 : node43008;
														assign node43008 = (inp[15]) ? node43014 : node43009;
															assign node43009 = (inp[5]) ? node43011 : 4'b0010;
																assign node43011 = (inp[3]) ? 4'b0000 : 4'b0010;
															assign node43014 = (inp[5]) ? node43016 : 4'b0000;
																assign node43016 = (inp[3]) ? 4'b0010 : 4'b0000;
														assign node43019 = (inp[15]) ? node43023 : node43020;
															assign node43020 = (inp[5]) ? 4'b0010 : 4'b0000;
															assign node43023 = (inp[3]) ? node43025 : 4'b0010;
																assign node43025 = (inp[5]) ? 4'b0000 : 4'b0010;
													assign node43028 = (inp[3]) ? node43034 : node43029;
														assign node43029 = (inp[5]) ? node43031 : 4'b0110;
															assign node43031 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node43034 = (inp[0]) ? node43038 : node43035;
															assign node43035 = (inp[15]) ? 4'b0110 : 4'b0100;
															assign node43038 = (inp[15]) ? 4'b0100 : 4'b0110;
												assign node43041 = (inp[9]) ? node43053 : node43042;
													assign node43042 = (inp[0]) ? node43048 : node43043;
														assign node43043 = (inp[15]) ? 4'b0110 : node43044;
															assign node43044 = (inp[5]) ? 4'b0100 : 4'b0110;
														assign node43048 = (inp[15]) ? 4'b0100 : node43049;
															assign node43049 = (inp[3]) ? 4'b0110 : 4'b0100;
													assign node43053 = (inp[3]) ? node43063 : node43054;
														assign node43054 = (inp[15]) ? 4'b0000 : node43055;
															assign node43055 = (inp[5]) ? node43059 : node43056;
																assign node43056 = (inp[0]) ? 4'b0000 : 4'b0010;
																assign node43059 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node43063 = (inp[5]) ? node43069 : node43064;
															assign node43064 = (inp[15]) ? node43066 : 4'b0000;
																assign node43066 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node43069 = (inp[0]) ? node43073 : node43070;
																assign node43070 = (inp[15]) ? 4'b0010 : 4'b0000;
																assign node43073 = (inp[15]) ? 4'b0000 : 4'b0010;
										assign node43076 = (inp[5]) ? node43130 : node43077;
											assign node43077 = (inp[15]) ? node43101 : node43078;
												assign node43078 = (inp[0]) ? node43088 : node43079;
													assign node43079 = (inp[9]) ? node43081 : 4'b1011;
														assign node43081 = (inp[4]) ? node43085 : node43082;
															assign node43082 = (inp[3]) ? 4'b1101 : 4'b1111;
															assign node43085 = (inp[3]) ? 4'b1001 : 4'b1011;
													assign node43088 = (inp[3]) ? node43096 : node43089;
														assign node43089 = (inp[4]) ? node43093 : node43090;
															assign node43090 = (inp[9]) ? 4'b1101 : 4'b1001;
															assign node43093 = (inp[12]) ? 4'b1101 : 4'b1001;
														assign node43096 = (inp[4]) ? node43098 : 4'b1001;
															assign node43098 = (inp[9]) ? 4'b1011 : 4'b1111;
												assign node43101 = (inp[0]) ? node43115 : node43102;
													assign node43102 = (inp[3]) ? node43110 : node43103;
														assign node43103 = (inp[9]) ? node43107 : node43104;
															assign node43104 = (inp[4]) ? 4'b1101 : 4'b1001;
															assign node43107 = (inp[4]) ? 4'b1001 : 4'b1101;
														assign node43110 = (inp[9]) ? node43112 : 4'b1001;
															assign node43112 = (inp[4]) ? 4'b1011 : 4'b1111;
													assign node43115 = (inp[3]) ? node43123 : node43116;
														assign node43116 = (inp[12]) ? 4'b1111 : node43117;
															assign node43117 = (inp[9]) ? 4'b1011 : node43118;
																assign node43118 = (inp[4]) ? 4'b1111 : 4'b1011;
														assign node43123 = (inp[4]) ? node43127 : node43124;
															assign node43124 = (inp[9]) ? 4'b1101 : 4'b1011;
															assign node43127 = (inp[9]) ? 4'b1001 : 4'b1101;
											assign node43130 = (inp[0]) ? node43146 : node43131;
												assign node43131 = (inp[15]) ? node43141 : node43132;
													assign node43132 = (inp[9]) ? node43138 : node43133;
														assign node43133 = (inp[3]) ? node43135 : 4'b1011;
															assign node43135 = (inp[4]) ? 4'b1101 : 4'b1001;
														assign node43138 = (inp[4]) ? 4'b1001 : 4'b1101;
													assign node43141 = (inp[9]) ? node43143 : 4'b1111;
														assign node43143 = (inp[4]) ? 4'b1011 : 4'b1111;
												assign node43146 = (inp[15]) ? node43156 : node43147;
													assign node43147 = (inp[9]) ? node43153 : node43148;
														assign node43148 = (inp[4]) ? 4'b1111 : node43149;
															assign node43149 = (inp[3]) ? 4'b1011 : 4'b1001;
														assign node43153 = (inp[4]) ? 4'b1011 : 4'b1111;
													assign node43156 = (inp[9]) ? node43162 : node43157;
														assign node43157 = (inp[4]) ? 4'b1101 : node43158;
															assign node43158 = (inp[3]) ? 4'b1001 : 4'b1011;
														assign node43162 = (inp[4]) ? 4'b1001 : 4'b1101;
									assign node43165 = (inp[4]) ? node43229 : node43166;
										assign node43166 = (inp[9]) ? node43190 : node43167;
											assign node43167 = (inp[15]) ? node43179 : node43168;
												assign node43168 = (inp[0]) ? node43174 : node43169;
													assign node43169 = (inp[5]) ? node43171 : 4'b1011;
														assign node43171 = (inp[3]) ? 4'b1001 : 4'b1011;
													assign node43174 = (inp[3]) ? node43176 : 4'b1001;
														assign node43176 = (inp[5]) ? 4'b1011 : 4'b1001;
												assign node43179 = (inp[0]) ? node43185 : node43180;
													assign node43180 = (inp[3]) ? node43182 : 4'b1001;
														assign node43182 = (inp[5]) ? 4'b1011 : 4'b1001;
													assign node43185 = (inp[5]) ? node43187 : 4'b1011;
														assign node43187 = (inp[3]) ? 4'b1001 : 4'b1011;
											assign node43190 = (inp[12]) ? node43214 : node43191;
												assign node43191 = (inp[15]) ? node43203 : node43192;
													assign node43192 = (inp[0]) ? node43198 : node43193;
														assign node43193 = (inp[5]) ? 4'b1101 : node43194;
															assign node43194 = (inp[3]) ? 4'b1101 : 4'b1111;
														assign node43198 = (inp[5]) ? 4'b1111 : node43199;
															assign node43199 = (inp[3]) ? 4'b1111 : 4'b1101;
													assign node43203 = (inp[0]) ? node43209 : node43204;
														assign node43204 = (inp[3]) ? 4'b1111 : node43205;
															assign node43205 = (inp[5]) ? 4'b1111 : 4'b1101;
														assign node43209 = (inp[5]) ? 4'b1101 : node43210;
															assign node43210 = (inp[3]) ? 4'b1101 : 4'b1111;
												assign node43214 = (inp[5]) ? node43222 : node43215;
													assign node43215 = (inp[0]) ? node43217 : 4'b1101;
														assign node43217 = (inp[15]) ? node43219 : 4'b1111;
															assign node43219 = (inp[3]) ? 4'b1101 : 4'b1111;
													assign node43222 = (inp[0]) ? node43226 : node43223;
														assign node43223 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node43226 = (inp[15]) ? 4'b1101 : 4'b1111;
										assign node43229 = (inp[9]) ? node43253 : node43230;
											assign node43230 = (inp[0]) ? node43242 : node43231;
												assign node43231 = (inp[15]) ? node43237 : node43232;
													assign node43232 = (inp[3]) ? 4'b1101 : node43233;
														assign node43233 = (inp[5]) ? 4'b1101 : 4'b1111;
													assign node43237 = (inp[3]) ? 4'b1111 : node43238;
														assign node43238 = (inp[5]) ? 4'b1111 : 4'b1101;
												assign node43242 = (inp[15]) ? node43248 : node43243;
													assign node43243 = (inp[5]) ? 4'b1111 : node43244;
														assign node43244 = (inp[3]) ? 4'b1111 : 4'b1101;
													assign node43248 = (inp[12]) ? node43250 : 4'b1101;
														assign node43250 = (inp[3]) ? 4'b1101 : 4'b1111;
											assign node43253 = (inp[15]) ? node43265 : node43254;
												assign node43254 = (inp[0]) ? node43260 : node43255;
													assign node43255 = (inp[5]) ? 4'b1001 : node43256;
														assign node43256 = (inp[3]) ? 4'b1001 : 4'b1011;
													assign node43260 = (inp[3]) ? 4'b1011 : node43261;
														assign node43261 = (inp[5]) ? 4'b1011 : 4'b1001;
												assign node43265 = (inp[0]) ? node43271 : node43266;
													assign node43266 = (inp[5]) ? 4'b1011 : node43267;
														assign node43267 = (inp[3]) ? 4'b1011 : 4'b1001;
													assign node43271 = (inp[3]) ? 4'b1001 : node43272;
														assign node43272 = (inp[5]) ? 4'b1001 : 4'b1011;
							assign node43276 = (inp[8]) ? node43636 : node43277;
								assign node43277 = (inp[2]) ? node43503 : node43278;
									assign node43278 = (inp[14]) ? node43376 : node43279;
										assign node43279 = (inp[12]) ? node43327 : node43280;
											assign node43280 = (inp[4]) ? node43306 : node43281;
												assign node43281 = (inp[9]) ? node43291 : node43282;
													assign node43282 = (inp[0]) ? 4'b0110 : node43283;
														assign node43283 = (inp[15]) ? 4'b0100 : node43284;
															assign node43284 = (inp[5]) ? node43286 : 4'b0110;
																assign node43286 = (inp[3]) ? 4'b0100 : 4'b0110;
													assign node43291 = (inp[0]) ? node43301 : node43292;
														assign node43292 = (inp[3]) ? node43294 : 4'b0010;
															assign node43294 = (inp[15]) ? node43298 : node43295;
																assign node43295 = (inp[5]) ? 4'b0000 : 4'b0010;
																assign node43298 = (inp[5]) ? 4'b0010 : 4'b0000;
														assign node43301 = (inp[15]) ? node43303 : 4'b0000;
															assign node43303 = (inp[5]) ? 4'b0000 : 4'b0010;
												assign node43306 = (inp[9]) ? node43318 : node43307;
													assign node43307 = (inp[3]) ? 4'b0010 : node43308;
														assign node43308 = (inp[5]) ? 4'b0000 : node43309;
															assign node43309 = (inp[15]) ? node43313 : node43310;
																assign node43310 = (inp[0]) ? 4'b0000 : 4'b0010;
																assign node43313 = (inp[0]) ? 4'b0010 : 4'b0000;
													assign node43318 = (inp[15]) ? node43322 : node43319;
														assign node43319 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node43322 = (inp[0]) ? node43324 : 4'b0110;
															assign node43324 = (inp[5]) ? 4'b0100 : 4'b0110;
											assign node43327 = (inp[0]) ? node43345 : node43328;
												assign node43328 = (inp[15]) ? node43336 : node43329;
													assign node43329 = (inp[9]) ? node43333 : node43330;
														assign node43330 = (inp[4]) ? 4'b0100 : 4'b0010;
														assign node43333 = (inp[4]) ? 4'b0000 : 4'b0100;
													assign node43336 = (inp[5]) ? 4'b0110 : node43337;
														assign node43337 = (inp[9]) ? 4'b0110 : node43338;
															assign node43338 = (inp[4]) ? node43340 : 4'b0000;
																assign node43340 = (inp[3]) ? 4'b0110 : 4'b0100;
												assign node43345 = (inp[15]) ? node43363 : node43346;
													assign node43346 = (inp[3]) ? node43352 : node43347;
														assign node43347 = (inp[5]) ? node43349 : 4'b0000;
															assign node43349 = (inp[4]) ? 4'b0110 : 4'b0000;
														assign node43352 = (inp[5]) ? node43358 : node43353;
															assign node43353 = (inp[4]) ? 4'b0110 : node43354;
																assign node43354 = (inp[9]) ? 4'b0110 : 4'b0000;
															assign node43358 = (inp[9]) ? node43360 : 4'b0010;
																assign node43360 = (inp[4]) ? 4'b0010 : 4'b0110;
													assign node43363 = (inp[5]) ? node43369 : node43364;
														assign node43364 = (inp[9]) ? 4'b0100 : node43365;
															assign node43365 = (inp[4]) ? 4'b0110 : 4'b0010;
														assign node43369 = (inp[4]) ? node43373 : node43370;
															assign node43370 = (inp[9]) ? 4'b0100 : 4'b0000;
															assign node43373 = (inp[9]) ? 4'b0000 : 4'b0100;
										assign node43376 = (inp[5]) ? node43456 : node43377;
											assign node43377 = (inp[12]) ? node43413 : node43378;
												assign node43378 = (inp[15]) ? node43396 : node43379;
													assign node43379 = (inp[0]) ? node43389 : node43380;
														assign node43380 = (inp[3]) ? node43384 : node43381;
															assign node43381 = (inp[4]) ? 4'b1011 : 4'b1111;
															assign node43384 = (inp[4]) ? node43386 : 4'b1011;
																assign node43386 = (inp[9]) ? 4'b1001 : 4'b1101;
														assign node43389 = (inp[3]) ? 4'b1111 : node43390;
															assign node43390 = (inp[9]) ? 4'b1001 : node43391;
																assign node43391 = (inp[4]) ? 4'b1101 : 4'b1001;
													assign node43396 = (inp[4]) ? node43406 : node43397;
														assign node43397 = (inp[9]) ? node43401 : node43398;
															assign node43398 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node43401 = (inp[3]) ? 4'b1111 : node43402;
																assign node43402 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node43406 = (inp[3]) ? node43410 : node43407;
															assign node43407 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node43410 = (inp[0]) ? 4'b1101 : 4'b1111;
												assign node43413 = (inp[0]) ? node43433 : node43414;
													assign node43414 = (inp[3]) ? node43422 : node43415;
														assign node43415 = (inp[9]) ? node43419 : node43416;
															assign node43416 = (inp[4]) ? 4'b1111 : 4'b1011;
															assign node43419 = (inp[4]) ? 4'b1011 : 4'b1111;
														assign node43422 = (inp[15]) ? node43428 : node43423;
															assign node43423 = (inp[9]) ? 4'b1101 : node43424;
																assign node43424 = (inp[4]) ? 4'b1101 : 4'b1011;
															assign node43428 = (inp[4]) ? node43430 : 4'b1111;
																assign node43430 = (inp[9]) ? 4'b1011 : 4'b1111;
													assign node43433 = (inp[4]) ? node43443 : node43434;
														assign node43434 = (inp[9]) ? node43436 : 4'b1011;
															assign node43436 = (inp[3]) ? node43440 : node43437;
																assign node43437 = (inp[15]) ? 4'b1111 : 4'b1101;
																assign node43440 = (inp[15]) ? 4'b1101 : 4'b1111;
														assign node43443 = (inp[9]) ? node43449 : node43444;
															assign node43444 = (inp[3]) ? node43446 : 4'b1111;
																assign node43446 = (inp[15]) ? 4'b1101 : 4'b1111;
															assign node43449 = (inp[3]) ? node43453 : node43450;
																assign node43450 = (inp[15]) ? 4'b1011 : 4'b1001;
																assign node43453 = (inp[15]) ? 4'b1001 : 4'b1011;
											assign node43456 = (inp[9]) ? node43480 : node43457;
												assign node43457 = (inp[4]) ? node43467 : node43458;
													assign node43458 = (inp[3]) ? node43460 : 4'b1011;
														assign node43460 = (inp[0]) ? node43464 : node43461;
															assign node43461 = (inp[15]) ? 4'b1011 : 4'b1001;
															assign node43464 = (inp[15]) ? 4'b1001 : 4'b1011;
													assign node43467 = (inp[3]) ? node43473 : node43468;
														assign node43468 = (inp[0]) ? 4'b1111 : node43469;
															assign node43469 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node43473 = (inp[15]) ? node43477 : node43474;
															assign node43474 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node43477 = (inp[0]) ? 4'b1101 : 4'b1111;
												assign node43480 = (inp[4]) ? node43488 : node43481;
													assign node43481 = (inp[15]) ? node43485 : node43482;
														assign node43482 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node43485 = (inp[0]) ? 4'b1101 : 4'b1111;
													assign node43488 = (inp[3]) ? node43494 : node43489;
														assign node43489 = (inp[15]) ? 4'b1001 : node43490;
															assign node43490 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node43494 = (inp[12]) ? 4'b1011 : node43495;
															assign node43495 = (inp[15]) ? node43499 : node43496;
																assign node43496 = (inp[0]) ? 4'b1011 : 4'b1001;
																assign node43499 = (inp[0]) ? 4'b1001 : 4'b1011;
									assign node43503 = (inp[9]) ? node43551 : node43504;
										assign node43504 = (inp[4]) ? node43528 : node43505;
											assign node43505 = (inp[0]) ? node43517 : node43506;
												assign node43506 = (inp[15]) ? node43512 : node43507;
													assign node43507 = (inp[5]) ? node43509 : 4'b1011;
														assign node43509 = (inp[3]) ? 4'b1001 : 4'b1011;
													assign node43512 = (inp[5]) ? node43514 : 4'b1001;
														assign node43514 = (inp[3]) ? 4'b1011 : 4'b1001;
												assign node43517 = (inp[15]) ? node43523 : node43518;
													assign node43518 = (inp[5]) ? node43520 : 4'b1001;
														assign node43520 = (inp[3]) ? 4'b1011 : 4'b1001;
													assign node43523 = (inp[5]) ? node43525 : 4'b1011;
														assign node43525 = (inp[3]) ? 4'b1001 : 4'b1011;
											assign node43528 = (inp[0]) ? node43540 : node43529;
												assign node43529 = (inp[15]) ? node43535 : node43530;
													assign node43530 = (inp[3]) ? 4'b1101 : node43531;
														assign node43531 = (inp[5]) ? 4'b1101 : 4'b1111;
													assign node43535 = (inp[5]) ? 4'b1111 : node43536;
														assign node43536 = (inp[3]) ? 4'b1111 : 4'b1101;
												assign node43540 = (inp[15]) ? node43546 : node43541;
													assign node43541 = (inp[5]) ? 4'b1111 : node43542;
														assign node43542 = (inp[3]) ? 4'b1111 : 4'b1101;
													assign node43546 = (inp[5]) ? 4'b1101 : node43547;
														assign node43547 = (inp[3]) ? 4'b1101 : 4'b1111;
										assign node43551 = (inp[4]) ? node43601 : node43552;
											assign node43552 = (inp[12]) ? node43572 : node43553;
												assign node43553 = (inp[0]) ? node43565 : node43554;
													assign node43554 = (inp[15]) ? node43560 : node43555;
														assign node43555 = (inp[3]) ? 4'b1101 : node43556;
															assign node43556 = (inp[5]) ? 4'b1101 : 4'b1111;
														assign node43560 = (inp[5]) ? 4'b1111 : node43561;
															assign node43561 = (inp[14]) ? 4'b1111 : 4'b1101;
													assign node43565 = (inp[15]) ? 4'b1101 : node43566;
														assign node43566 = (inp[3]) ? 4'b1111 : node43567;
															assign node43567 = (inp[5]) ? 4'b1111 : 4'b1101;
												assign node43572 = (inp[5]) ? node43588 : node43573;
													assign node43573 = (inp[3]) ? node43581 : node43574;
														assign node43574 = (inp[15]) ? node43578 : node43575;
															assign node43575 = (inp[0]) ? 4'b1101 : 4'b1111;
															assign node43578 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node43581 = (inp[15]) ? node43585 : node43582;
															assign node43582 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node43585 = (inp[0]) ? 4'b1101 : 4'b1111;
													assign node43588 = (inp[14]) ? node43596 : node43589;
														assign node43589 = (inp[0]) ? node43593 : node43590;
															assign node43590 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node43593 = (inp[15]) ? 4'b1101 : 4'b1111;
														assign node43596 = (inp[15]) ? node43598 : 4'b1111;
															assign node43598 = (inp[0]) ? 4'b1101 : 4'b1111;
											assign node43601 = (inp[5]) ? node43629 : node43602;
												assign node43602 = (inp[3]) ? node43616 : node43603;
													assign node43603 = (inp[14]) ? node43611 : node43604;
														assign node43604 = (inp[0]) ? node43608 : node43605;
															assign node43605 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node43608 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node43611 = (inp[0]) ? 4'b1001 : node43612;
															assign node43612 = (inp[15]) ? 4'b1001 : 4'b1011;
													assign node43616 = (inp[12]) ? node43624 : node43617;
														assign node43617 = (inp[15]) ? node43621 : node43618;
															assign node43618 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node43621 = (inp[0]) ? 4'b1001 : 4'b1011;
														assign node43624 = (inp[0]) ? node43626 : 4'b1001;
															assign node43626 = (inp[15]) ? 4'b1001 : 4'b1011;
												assign node43629 = (inp[0]) ? node43633 : node43630;
													assign node43630 = (inp[15]) ? 4'b1011 : 4'b1001;
													assign node43633 = (inp[15]) ? 4'b1001 : 4'b1011;
								assign node43636 = (inp[2]) ? node43844 : node43637;
									assign node43637 = (inp[14]) ? node43741 : node43638;
										assign node43638 = (inp[3]) ? node43686 : node43639;
											assign node43639 = (inp[15]) ? node43661 : node43640;
												assign node43640 = (inp[5]) ? node43652 : node43641;
													assign node43641 = (inp[0]) ? node43647 : node43642;
														assign node43642 = (inp[9]) ? node43644 : 4'b1011;
															assign node43644 = (inp[4]) ? 4'b1011 : 4'b1111;
														assign node43647 = (inp[9]) ? node43649 : 4'b1001;
															assign node43649 = (inp[4]) ? 4'b1001 : 4'b1101;
													assign node43652 = (inp[0]) ? node43656 : node43653;
														assign node43653 = (inp[9]) ? 4'b1001 : 4'b1101;
														assign node43656 = (inp[4]) ? 4'b1111 : node43657;
															assign node43657 = (inp[9]) ? 4'b1111 : 4'b1001;
												assign node43661 = (inp[0]) ? node43671 : node43662;
													assign node43662 = (inp[5]) ? node43664 : 4'b1101;
														assign node43664 = (inp[9]) ? node43668 : node43665;
															assign node43665 = (inp[4]) ? 4'b1111 : 4'b1001;
															assign node43668 = (inp[4]) ? 4'b1011 : 4'b1111;
													assign node43671 = (inp[5]) ? node43681 : node43672;
														assign node43672 = (inp[12]) ? 4'b1111 : node43673;
															assign node43673 = (inp[9]) ? node43677 : node43674;
																assign node43674 = (inp[4]) ? 4'b1111 : 4'b1011;
																assign node43677 = (inp[4]) ? 4'b1011 : 4'b1111;
														assign node43681 = (inp[4]) ? node43683 : 4'b1011;
															assign node43683 = (inp[9]) ? 4'b1001 : 4'b1101;
											assign node43686 = (inp[0]) ? node43710 : node43687;
												assign node43687 = (inp[15]) ? node43703 : node43688;
													assign node43688 = (inp[5]) ? node43696 : node43689;
														assign node43689 = (inp[4]) ? node43693 : node43690;
															assign node43690 = (inp[9]) ? 4'b1101 : 4'b1011;
															assign node43693 = (inp[9]) ? 4'b1001 : 4'b1101;
														assign node43696 = (inp[4]) ? node43700 : node43697;
															assign node43697 = (inp[9]) ? 4'b1101 : 4'b1001;
															assign node43700 = (inp[9]) ? 4'b1001 : 4'b1101;
													assign node43703 = (inp[5]) ? 4'b1111 : node43704;
														assign node43704 = (inp[4]) ? node43706 : 4'b1001;
															assign node43706 = (inp[9]) ? 4'b1011 : 4'b1111;
												assign node43710 = (inp[15]) ? node43732 : node43711;
													assign node43711 = (inp[12]) ? node43723 : node43712;
														assign node43712 = (inp[5]) ? node43718 : node43713;
															assign node43713 = (inp[9]) ? node43715 : 4'b1111;
																assign node43715 = (inp[4]) ? 4'b1011 : 4'b1111;
															assign node43718 = (inp[4]) ? node43720 : 4'b1011;
																assign node43720 = (inp[9]) ? 4'b1011 : 4'b1111;
														assign node43723 = (inp[5]) ? node43727 : node43724;
															assign node43724 = (inp[9]) ? 4'b1111 : 4'b1001;
															assign node43727 = (inp[9]) ? node43729 : 4'b1111;
																assign node43729 = (inp[4]) ? 4'b1011 : 4'b1111;
													assign node43732 = (inp[9]) ? node43738 : node43733;
														assign node43733 = (inp[4]) ? 4'b1101 : node43734;
															assign node43734 = (inp[5]) ? 4'b1001 : 4'b1011;
														assign node43738 = (inp[4]) ? 4'b1001 : 4'b1101;
										assign node43741 = (inp[3]) ? node43799 : node43742;
											assign node43742 = (inp[9]) ? node43768 : node43743;
												assign node43743 = (inp[4]) ? node43751 : node43744;
													assign node43744 = (inp[0]) ? node43748 : node43745;
														assign node43745 = (inp[15]) ? 4'b1000 : 4'b1010;
														assign node43748 = (inp[15]) ? 4'b1010 : 4'b1000;
													assign node43751 = (inp[5]) ? node43761 : node43752;
														assign node43752 = (inp[12]) ? node43754 : 4'b1110;
															assign node43754 = (inp[0]) ? node43758 : node43755;
																assign node43755 = (inp[15]) ? 4'b1100 : 4'b1110;
																assign node43758 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node43761 = (inp[12]) ? 4'b1110 : node43762;
															assign node43762 = (inp[0]) ? 4'b1100 : node43763;
																assign node43763 = (inp[15]) ? 4'b1110 : 4'b1100;
												assign node43768 = (inp[4]) ? node43786 : node43769;
													assign node43769 = (inp[0]) ? node43777 : node43770;
														assign node43770 = (inp[5]) ? node43774 : node43771;
															assign node43771 = (inp[15]) ? 4'b1100 : 4'b1110;
															assign node43774 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node43777 = (inp[12]) ? node43779 : 4'b1110;
															assign node43779 = (inp[15]) ? node43783 : node43780;
																assign node43780 = (inp[5]) ? 4'b1110 : 4'b1100;
																assign node43783 = (inp[5]) ? 4'b1100 : 4'b1110;
													assign node43786 = (inp[15]) ? node43792 : node43787;
														assign node43787 = (inp[5]) ? 4'b1010 : node43788;
															assign node43788 = (inp[12]) ? 4'b1000 : 4'b1010;
														assign node43792 = (inp[5]) ? node43796 : node43793;
															assign node43793 = (inp[0]) ? 4'b1010 : 4'b1000;
															assign node43796 = (inp[0]) ? 4'b1000 : 4'b1010;
											assign node43799 = (inp[9]) ? node43829 : node43800;
												assign node43800 = (inp[4]) ? node43816 : node43801;
													assign node43801 = (inp[15]) ? node43809 : node43802;
														assign node43802 = (inp[12]) ? node43804 : 4'b1010;
															assign node43804 = (inp[0]) ? 4'b1000 : node43805;
																assign node43805 = (inp[5]) ? 4'b1000 : 4'b1010;
														assign node43809 = (inp[0]) ? node43813 : node43810;
															assign node43810 = (inp[5]) ? 4'b1010 : 4'b1000;
															assign node43813 = (inp[5]) ? 4'b1000 : 4'b1010;
													assign node43816 = (inp[5]) ? node43824 : node43817;
														assign node43817 = (inp[0]) ? node43821 : node43818;
															assign node43818 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node43821 = (inp[15]) ? 4'b1100 : 4'b1110;
														assign node43824 = (inp[15]) ? 4'b1100 : node43825;
															assign node43825 = (inp[0]) ? 4'b1110 : 4'b1100;
												assign node43829 = (inp[4]) ? node43837 : node43830;
													assign node43830 = (inp[15]) ? node43834 : node43831;
														assign node43831 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node43834 = (inp[0]) ? 4'b1100 : 4'b1110;
													assign node43837 = (inp[0]) ? node43841 : node43838;
														assign node43838 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node43841 = (inp[15]) ? 4'b1000 : 4'b1010;
									assign node43844 = (inp[4]) ? node43928 : node43845;
										assign node43845 = (inp[9]) ? node43889 : node43846;
											assign node43846 = (inp[12]) ? node43868 : node43847;
												assign node43847 = (inp[5]) ? node43855 : node43848;
													assign node43848 = (inp[15]) ? node43852 : node43849;
														assign node43849 = (inp[0]) ? 4'b1000 : 4'b1010;
														assign node43852 = (inp[0]) ? 4'b1010 : 4'b1000;
													assign node43855 = (inp[3]) ? node43863 : node43856;
														assign node43856 = (inp[15]) ? node43860 : node43857;
															assign node43857 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node43860 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node43863 = (inp[15]) ? node43865 : 4'b1000;
															assign node43865 = (inp[0]) ? 4'b1000 : 4'b1010;
												assign node43868 = (inp[5]) ? node43876 : node43869;
													assign node43869 = (inp[15]) ? node43873 : node43870;
														assign node43870 = (inp[0]) ? 4'b1000 : 4'b1010;
														assign node43873 = (inp[0]) ? 4'b1010 : 4'b1000;
													assign node43876 = (inp[3]) ? node43878 : 4'b1010;
														assign node43878 = (inp[14]) ? node43884 : node43879;
															assign node43879 = (inp[0]) ? node43881 : 4'b1010;
																assign node43881 = (inp[15]) ? 4'b1000 : 4'b1010;
															assign node43884 = (inp[15]) ? 4'b1010 : node43885;
																assign node43885 = (inp[0]) ? 4'b1010 : 4'b1000;
											assign node43889 = (inp[5]) ? node43921 : node43890;
												assign node43890 = (inp[12]) ? node43906 : node43891;
													assign node43891 = (inp[15]) ? node43901 : node43892;
														assign node43892 = (inp[14]) ? 4'b1100 : node43893;
															assign node43893 = (inp[3]) ? node43897 : node43894;
																assign node43894 = (inp[0]) ? 4'b1100 : 4'b1110;
																assign node43897 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node43901 = (inp[0]) ? node43903 : 4'b1110;
															assign node43903 = (inp[14]) ? 4'b1110 : 4'b1100;
													assign node43906 = (inp[0]) ? node43914 : node43907;
														assign node43907 = (inp[15]) ? node43911 : node43908;
															assign node43908 = (inp[3]) ? 4'b1100 : 4'b1110;
															assign node43911 = (inp[3]) ? 4'b1110 : 4'b1100;
														assign node43914 = (inp[3]) ? node43918 : node43915;
															assign node43915 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node43918 = (inp[15]) ? 4'b1100 : 4'b1110;
												assign node43921 = (inp[0]) ? node43925 : node43922;
													assign node43922 = (inp[15]) ? 4'b1110 : 4'b1100;
													assign node43925 = (inp[15]) ? 4'b1100 : 4'b1110;
										assign node43928 = (inp[9]) ? node43954 : node43929;
											assign node43929 = (inp[3]) ? node43947 : node43930;
												assign node43930 = (inp[0]) ? node43938 : node43931;
													assign node43931 = (inp[15]) ? node43935 : node43932;
														assign node43932 = (inp[5]) ? 4'b1100 : 4'b1110;
														assign node43935 = (inp[5]) ? 4'b1110 : 4'b1100;
													assign node43938 = (inp[14]) ? 4'b1100 : node43939;
														assign node43939 = (inp[15]) ? node43943 : node43940;
															assign node43940 = (inp[5]) ? 4'b1110 : 4'b1100;
															assign node43943 = (inp[5]) ? 4'b1100 : 4'b1110;
												assign node43947 = (inp[15]) ? node43951 : node43948;
													assign node43948 = (inp[0]) ? 4'b1110 : 4'b1100;
													assign node43951 = (inp[0]) ? 4'b1100 : 4'b1110;
											assign node43954 = (inp[12]) ? node43972 : node43955;
												assign node43955 = (inp[0]) ? node43963 : node43956;
													assign node43956 = (inp[3]) ? 4'b1000 : node43957;
														assign node43957 = (inp[5]) ? 4'b1000 : node43958;
															assign node43958 = (inp[15]) ? 4'b1000 : 4'b1010;
													assign node43963 = (inp[15]) ? node43969 : node43964;
														assign node43964 = (inp[14]) ? 4'b1010 : node43965;
															assign node43965 = (inp[3]) ? 4'b1010 : 4'b1000;
														assign node43969 = (inp[5]) ? 4'b1000 : 4'b1010;
												assign node43972 = (inp[0]) ? node43982 : node43973;
													assign node43973 = (inp[15]) ? node43977 : node43974;
														assign node43974 = (inp[3]) ? 4'b1000 : 4'b1010;
														assign node43977 = (inp[5]) ? 4'b1010 : node43978;
															assign node43978 = (inp[3]) ? 4'b1010 : 4'b1000;
													assign node43982 = (inp[15]) ? node43988 : node43983;
														assign node43983 = (inp[3]) ? 4'b1010 : node43984;
															assign node43984 = (inp[5]) ? 4'b1010 : 4'b1000;
														assign node43988 = (inp[5]) ? 4'b1000 : 4'b1010;
					assign node43991 = (inp[1]) ? node45749 : node43992;
						assign node43992 = (inp[8]) ? node44858 : node43993;
							assign node43993 = (inp[7]) ? node44439 : node43994;
								assign node43994 = (inp[14]) ? node44232 : node43995;
									assign node43995 = (inp[2]) ? node44123 : node43996;
										assign node43996 = (inp[3]) ? node44062 : node43997;
											assign node43997 = (inp[9]) ? node44025 : node43998;
												assign node43998 = (inp[4]) ? node44010 : node43999;
													assign node43999 = (inp[12]) ? node44005 : node44000;
														assign node44000 = (inp[15]) ? node44002 : 4'b0101;
															assign node44002 = (inp[0]) ? 4'b0111 : 4'b0101;
														assign node44005 = (inp[15]) ? node44007 : 4'b0001;
															assign node44007 = (inp[0]) ? 4'b0011 : 4'b0001;
													assign node44010 = (inp[12]) ? node44016 : node44011;
														assign node44011 = (inp[15]) ? node44013 : 4'b0011;
															assign node44013 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node44016 = (inp[15]) ? node44018 : 4'b0111;
															assign node44018 = (inp[5]) ? node44022 : node44019;
																assign node44019 = (inp[0]) ? 4'b0111 : 4'b0101;
																assign node44022 = (inp[0]) ? 4'b0101 : 4'b0111;
												assign node44025 = (inp[15]) ? node44047 : node44026;
													assign node44026 = (inp[12]) ? node44034 : node44027;
														assign node44027 = (inp[4]) ? node44029 : 4'b0011;
															assign node44029 = (inp[0]) ? 4'b0111 : node44030;
																assign node44030 = (inp[5]) ? 4'b0101 : 4'b0111;
														assign node44034 = (inp[4]) ? node44042 : node44035;
															assign node44035 = (inp[0]) ? node44039 : node44036;
																assign node44036 = (inp[5]) ? 4'b0101 : 4'b0111;
																assign node44039 = (inp[5]) ? 4'b0111 : 4'b0101;
															assign node44042 = (inp[0]) ? node44044 : 4'b0011;
																assign node44044 = (inp[5]) ? 4'b0011 : 4'b0001;
													assign node44047 = (inp[0]) ? node44055 : node44048;
														assign node44048 = (inp[12]) ? node44052 : node44049;
															assign node44049 = (inp[4]) ? 4'b0101 : 4'b0001;
															assign node44052 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node44055 = (inp[12]) ? node44059 : node44056;
															assign node44056 = (inp[4]) ? 4'b0111 : 4'b0011;
															assign node44059 = (inp[5]) ? 4'b0001 : 4'b0011;
											assign node44062 = (inp[0]) ? node44096 : node44063;
												assign node44063 = (inp[15]) ? node44081 : node44064;
													assign node44064 = (inp[9]) ? node44072 : node44065;
														assign node44065 = (inp[5]) ? 4'b0001 : node44066;
															assign node44066 = (inp[12]) ? node44068 : 4'b0011;
																assign node44068 = (inp[4]) ? 4'b0101 : 4'b0011;
														assign node44072 = (inp[4]) ? node44078 : node44073;
															assign node44073 = (inp[12]) ? 4'b0101 : node44074;
																assign node44074 = (inp[5]) ? 4'b0001 : 4'b0011;
															assign node44078 = (inp[12]) ? 4'b0001 : 4'b0101;
													assign node44081 = (inp[9]) ? node44087 : node44082;
														assign node44082 = (inp[5]) ? 4'b0111 : node44083;
															assign node44083 = (inp[12]) ? 4'b0111 : 4'b0001;
														assign node44087 = (inp[5]) ? node44089 : 4'b0011;
															assign node44089 = (inp[4]) ? node44093 : node44090;
																assign node44090 = (inp[12]) ? 4'b0111 : 4'b0011;
																assign node44093 = (inp[12]) ? 4'b0011 : 4'b0111;
												assign node44096 = (inp[5]) ? node44110 : node44097;
													assign node44097 = (inp[12]) ? node44105 : node44098;
														assign node44098 = (inp[4]) ? node44102 : node44099;
															assign node44099 = (inp[15]) ? 4'b0111 : 4'b0101;
															assign node44102 = (inp[15]) ? 4'b0011 : 4'b0111;
														assign node44105 = (inp[15]) ? 4'b0101 : node44106;
															assign node44106 = (inp[9]) ? 4'b0111 : 4'b0001;
													assign node44110 = (inp[15]) ? node44112 : 4'b0011;
														assign node44112 = (inp[12]) ? node44118 : node44113;
															assign node44113 = (inp[9]) ? node44115 : 4'b0101;
																assign node44115 = (inp[4]) ? 4'b0101 : 4'b0001;
															assign node44118 = (inp[4]) ? 4'b0001 : node44119;
																assign node44119 = (inp[9]) ? 4'b0101 : 4'b0001;
										assign node44123 = (inp[4]) ? node44177 : node44124;
											assign node44124 = (inp[12]) ? node44146 : node44125;
												assign node44125 = (inp[9]) ? node44139 : node44126;
													assign node44126 = (inp[3]) ? node44132 : node44127;
														assign node44127 = (inp[0]) ? 4'b0100 : node44128;
															assign node44128 = (inp[15]) ? 4'b0100 : 4'b0110;
														assign node44132 = (inp[5]) ? 4'b0110 : node44133;
															assign node44133 = (inp[0]) ? 4'b0110 : node44134;
																assign node44134 = (inp[15]) ? 4'b0100 : 4'b0110;
													assign node44139 = (inp[3]) ? 4'b0010 : node44140;
														assign node44140 = (inp[15]) ? 4'b0000 : node44141;
															assign node44141 = (inp[0]) ? 4'b0000 : 4'b0010;
												assign node44146 = (inp[9]) ? node44166 : node44147;
													assign node44147 = (inp[3]) ? node44153 : node44148;
														assign node44148 = (inp[15]) ? node44150 : 4'b0010;
															assign node44150 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node44153 = (inp[5]) ? node44161 : node44154;
															assign node44154 = (inp[15]) ? node44158 : node44155;
																assign node44155 = (inp[0]) ? 4'b0000 : 4'b0010;
																assign node44158 = (inp[0]) ? 4'b0010 : 4'b0000;
															assign node44161 = (inp[15]) ? node44163 : 4'b0000;
																assign node44163 = (inp[0]) ? 4'b0000 : 4'b0010;
													assign node44166 = (inp[0]) ? node44172 : node44167;
														assign node44167 = (inp[15]) ? 4'b0110 : node44168;
															assign node44168 = (inp[3]) ? 4'b0100 : 4'b0110;
														assign node44172 = (inp[5]) ? 4'b0100 : node44173;
															assign node44173 = (inp[3]) ? 4'b0110 : 4'b0100;
											assign node44177 = (inp[9]) ? node44199 : node44178;
												assign node44178 = (inp[12]) ? node44186 : node44179;
													assign node44179 = (inp[5]) ? node44181 : 4'b0000;
														assign node44181 = (inp[0]) ? node44183 : 4'b0010;
															assign node44183 = (inp[15]) ? 4'b0000 : 4'b0010;
													assign node44186 = (inp[15]) ? node44192 : node44187;
														assign node44187 = (inp[0]) ? 4'b0110 : node44188;
															assign node44188 = (inp[3]) ? 4'b0100 : 4'b0110;
														assign node44192 = (inp[0]) ? 4'b0100 : node44193;
															assign node44193 = (inp[3]) ? 4'b0110 : node44194;
																assign node44194 = (inp[5]) ? 4'b0110 : 4'b0100;
												assign node44199 = (inp[12]) ? node44209 : node44200;
													assign node44200 = (inp[3]) ? 4'b0100 : node44201;
														assign node44201 = (inp[15]) ? 4'b0110 : node44202;
															assign node44202 = (inp[0]) ? 4'b0100 : node44203;
																assign node44203 = (inp[5]) ? 4'b0100 : 4'b0110;
													assign node44209 = (inp[3]) ? node44225 : node44210;
														assign node44210 = (inp[15]) ? node44218 : node44211;
															assign node44211 = (inp[0]) ? node44215 : node44212;
																assign node44212 = (inp[5]) ? 4'b0000 : 4'b0010;
																assign node44215 = (inp[5]) ? 4'b0010 : 4'b0000;
															assign node44218 = (inp[0]) ? node44222 : node44219;
																assign node44219 = (inp[5]) ? 4'b0010 : 4'b0000;
																assign node44222 = (inp[5]) ? 4'b0000 : 4'b0010;
														assign node44225 = (inp[5]) ? 4'b0000 : node44226;
															assign node44226 = (inp[0]) ? 4'b0000 : node44227;
																assign node44227 = (inp[15]) ? 4'b0010 : 4'b0000;
									assign node44232 = (inp[0]) ? node44322 : node44233;
										assign node44233 = (inp[12]) ? node44287 : node44234;
											assign node44234 = (inp[15]) ? node44266 : node44235;
												assign node44235 = (inp[5]) ? node44249 : node44236;
													assign node44236 = (inp[2]) ? node44244 : node44237;
														assign node44237 = (inp[9]) ? node44241 : node44238;
															assign node44238 = (inp[4]) ? 4'b0010 : 4'b0110;
															assign node44241 = (inp[4]) ? 4'b0100 : 4'b0010;
														assign node44244 = (inp[9]) ? node44246 : 4'b0010;
															assign node44246 = (inp[4]) ? 4'b0110 : 4'b0010;
													assign node44249 = (inp[3]) ? node44257 : node44250;
														assign node44250 = (inp[4]) ? node44254 : node44251;
															assign node44251 = (inp[9]) ? 4'b0010 : 4'b0110;
															assign node44254 = (inp[9]) ? 4'b0100 : 4'b0010;
														assign node44257 = (inp[2]) ? 4'b0100 : node44258;
															assign node44258 = (inp[9]) ? node44262 : node44259;
																assign node44259 = (inp[4]) ? 4'b0000 : 4'b0100;
																assign node44262 = (inp[4]) ? 4'b0100 : 4'b0000;
												assign node44266 = (inp[3]) ? node44272 : node44267;
													assign node44267 = (inp[2]) ? node44269 : 4'b0000;
														assign node44269 = (inp[9]) ? 4'b0000 : 4'b0100;
													assign node44272 = (inp[5]) ? node44280 : node44273;
														assign node44273 = (inp[9]) ? node44277 : node44274;
															assign node44274 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node44277 = (inp[4]) ? 4'b0110 : 4'b0000;
														assign node44280 = (inp[4]) ? node44284 : node44281;
															assign node44281 = (inp[9]) ? 4'b0010 : 4'b0110;
															assign node44284 = (inp[9]) ? 4'b0110 : 4'b0010;
											assign node44287 = (inp[4]) ? node44303 : node44288;
												assign node44288 = (inp[9]) ? node44300 : node44289;
													assign node44289 = (inp[15]) ? node44295 : node44290;
														assign node44290 = (inp[5]) ? node44292 : 4'b0010;
															assign node44292 = (inp[3]) ? 4'b0000 : 4'b0010;
														assign node44295 = (inp[5]) ? node44297 : 4'b0000;
															assign node44297 = (inp[3]) ? 4'b0010 : 4'b0000;
													assign node44300 = (inp[5]) ? 4'b0110 : 4'b0100;
												assign node44303 = (inp[9]) ? node44311 : node44304;
													assign node44304 = (inp[15]) ? 4'b0110 : node44305;
														assign node44305 = (inp[5]) ? 4'b0100 : node44306;
															assign node44306 = (inp[3]) ? 4'b0100 : 4'b0110;
													assign node44311 = (inp[15]) ? node44317 : node44312;
														assign node44312 = (inp[5]) ? 4'b0000 : node44313;
															assign node44313 = (inp[3]) ? 4'b0000 : 4'b0010;
														assign node44317 = (inp[3]) ? 4'b0010 : node44318;
															assign node44318 = (inp[5]) ? 4'b0010 : 4'b0000;
										assign node44322 = (inp[5]) ? node44378 : node44323;
											assign node44323 = (inp[15]) ? node44349 : node44324;
												assign node44324 = (inp[3]) ? node44338 : node44325;
													assign node44325 = (inp[9]) ? node44331 : node44326;
														assign node44326 = (inp[4]) ? 4'b0000 : node44327;
															assign node44327 = (inp[12]) ? 4'b0000 : 4'b0100;
														assign node44331 = (inp[12]) ? node44335 : node44332;
															assign node44332 = (inp[4]) ? 4'b0100 : 4'b0000;
															assign node44335 = (inp[4]) ? 4'b0000 : 4'b0100;
													assign node44338 = (inp[4]) ? node44346 : node44339;
														assign node44339 = (inp[2]) ? 4'b0000 : node44340;
															assign node44340 = (inp[9]) ? 4'b0110 : node44341;
																assign node44341 = (inp[12]) ? 4'b0000 : 4'b0100;
														assign node44346 = (inp[12]) ? 4'b0010 : 4'b0110;
												assign node44349 = (inp[3]) ? node44365 : node44350;
													assign node44350 = (inp[9]) ? node44358 : node44351;
														assign node44351 = (inp[2]) ? node44353 : 4'b0110;
															assign node44353 = (inp[4]) ? 4'b0110 : node44354;
																assign node44354 = (inp[12]) ? 4'b0010 : 4'b0110;
														assign node44358 = (inp[12]) ? node44362 : node44359;
															assign node44359 = (inp[4]) ? 4'b0110 : 4'b0010;
															assign node44362 = (inp[4]) ? 4'b0010 : 4'b0110;
													assign node44365 = (inp[12]) ? node44371 : node44366;
														assign node44366 = (inp[4]) ? 4'b0010 : node44367;
															assign node44367 = (inp[9]) ? 4'b0010 : 4'b0110;
														assign node44371 = (inp[4]) ? node44375 : node44372;
															assign node44372 = (inp[2]) ? 4'b0100 : 4'b0010;
															assign node44375 = (inp[9]) ? 4'b0000 : 4'b0100;
											assign node44378 = (inp[15]) ? node44414 : node44379;
												assign node44379 = (inp[3]) ? node44395 : node44380;
													assign node44380 = (inp[12]) ? node44388 : node44381;
														assign node44381 = (inp[9]) ? node44385 : node44382;
															assign node44382 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node44385 = (inp[4]) ? 4'b0110 : 4'b0000;
														assign node44388 = (inp[9]) ? node44392 : node44389;
															assign node44389 = (inp[4]) ? 4'b0110 : 4'b0000;
															assign node44392 = (inp[4]) ? 4'b0010 : 4'b0110;
													assign node44395 = (inp[4]) ? node44405 : node44396;
														assign node44396 = (inp[2]) ? node44398 : 4'b0010;
															assign node44398 = (inp[9]) ? node44402 : node44399;
																assign node44399 = (inp[12]) ? 4'b0010 : 4'b0110;
																assign node44402 = (inp[12]) ? 4'b0110 : 4'b0010;
														assign node44405 = (inp[2]) ? 4'b0110 : node44406;
															assign node44406 = (inp[9]) ? node44410 : node44407;
																assign node44407 = (inp[12]) ? 4'b0110 : 4'b0010;
																assign node44410 = (inp[12]) ? 4'b0010 : 4'b0110;
												assign node44414 = (inp[4]) ? node44426 : node44415;
													assign node44415 = (inp[3]) ? node44419 : node44416;
														assign node44416 = (inp[12]) ? 4'b0010 : 4'b0110;
														assign node44419 = (inp[2]) ? node44421 : 4'b0100;
															assign node44421 = (inp[9]) ? 4'b0100 : node44422;
																assign node44422 = (inp[12]) ? 4'b0000 : 4'b0100;
													assign node44426 = (inp[3]) ? node44432 : node44427;
														assign node44427 = (inp[12]) ? node44429 : 4'b0100;
															assign node44429 = (inp[9]) ? 4'b0000 : 4'b0100;
														assign node44432 = (inp[9]) ? node44436 : node44433;
															assign node44433 = (inp[12]) ? 4'b0100 : 4'b0000;
															assign node44436 = (inp[12]) ? 4'b0000 : 4'b0100;
								assign node44439 = (inp[2]) ? node44669 : node44440;
									assign node44440 = (inp[14]) ? node44572 : node44441;
										assign node44441 = (inp[12]) ? node44505 : node44442;
											assign node44442 = (inp[5]) ? node44478 : node44443;
												assign node44443 = (inp[15]) ? node44463 : node44444;
													assign node44444 = (inp[0]) ? node44452 : node44445;
														assign node44445 = (inp[9]) ? node44449 : node44446;
															assign node44446 = (inp[4]) ? 4'b0010 : 4'b0110;
															assign node44449 = (inp[3]) ? 4'b0100 : 4'b0110;
														assign node44452 = (inp[3]) ? node44458 : node44453;
															assign node44453 = (inp[9]) ? node44455 : 4'b0100;
																assign node44455 = (inp[4]) ? 4'b0100 : 4'b0000;
															assign node44458 = (inp[9]) ? node44460 : 4'b0000;
																assign node44460 = (inp[4]) ? 4'b0110 : 4'b0000;
													assign node44463 = (inp[0]) ? node44471 : node44464;
														assign node44464 = (inp[9]) ? node44466 : 4'b0000;
															assign node44466 = (inp[4]) ? node44468 : 4'b0000;
																assign node44468 = (inp[3]) ? 4'b0110 : 4'b0100;
														assign node44471 = (inp[4]) ? node44475 : node44472;
															assign node44472 = (inp[9]) ? 4'b0010 : 4'b0110;
															assign node44475 = (inp[9]) ? 4'b0110 : 4'b0010;
												assign node44478 = (inp[15]) ? node44492 : node44479;
													assign node44479 = (inp[0]) ? node44481 : 4'b0010;
														assign node44481 = (inp[3]) ? node44485 : node44482;
															assign node44482 = (inp[4]) ? 4'b0110 : 4'b0000;
															assign node44485 = (inp[9]) ? node44489 : node44486;
																assign node44486 = (inp[4]) ? 4'b0010 : 4'b0110;
																assign node44489 = (inp[4]) ? 4'b0110 : 4'b0010;
													assign node44492 = (inp[4]) ? node44502 : node44493;
														assign node44493 = (inp[9]) ? node44499 : node44494;
															assign node44494 = (inp[0]) ? node44496 : 4'b0110;
																assign node44496 = (inp[3]) ? 4'b0100 : 4'b0110;
															assign node44499 = (inp[3]) ? 4'b0010 : 4'b0000;
														assign node44502 = (inp[3]) ? 4'b0000 : 4'b0010;
											assign node44505 = (inp[9]) ? node44543 : node44506;
												assign node44506 = (inp[4]) ? node44528 : node44507;
													assign node44507 = (inp[5]) ? node44515 : node44508;
														assign node44508 = (inp[0]) ? node44512 : node44509;
															assign node44509 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node44512 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node44515 = (inp[3]) ? node44521 : node44516;
															assign node44516 = (inp[0]) ? 4'b0010 : node44517;
																assign node44517 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node44521 = (inp[0]) ? node44525 : node44522;
																assign node44522 = (inp[15]) ? 4'b0010 : 4'b0000;
																assign node44525 = (inp[15]) ? 4'b0000 : 4'b0010;
													assign node44528 = (inp[15]) ? node44534 : node44529;
														assign node44529 = (inp[0]) ? node44531 : 4'b0100;
															assign node44531 = (inp[3]) ? 4'b0110 : 4'b0100;
														assign node44534 = (inp[5]) ? 4'b0110 : node44535;
															assign node44535 = (inp[0]) ? node44539 : node44536;
																assign node44536 = (inp[3]) ? 4'b0110 : 4'b0100;
																assign node44539 = (inp[3]) ? 4'b0100 : 4'b0110;
												assign node44543 = (inp[4]) ? node44555 : node44544;
													assign node44544 = (inp[0]) ? 4'b0100 : node44545;
														assign node44545 = (inp[15]) ? node44551 : node44546;
															assign node44546 = (inp[3]) ? 4'b0100 : node44547;
																assign node44547 = (inp[5]) ? 4'b0100 : 4'b0110;
															assign node44551 = (inp[5]) ? 4'b0110 : 4'b0100;
													assign node44555 = (inp[15]) ? node44563 : node44556;
														assign node44556 = (inp[0]) ? node44560 : node44557;
															assign node44557 = (inp[5]) ? 4'b0000 : 4'b0010;
															assign node44560 = (inp[5]) ? 4'b0010 : 4'b0000;
														assign node44563 = (inp[0]) ? node44567 : node44564;
															assign node44564 = (inp[5]) ? 4'b0010 : 4'b0000;
															assign node44567 = (inp[5]) ? 4'b0000 : node44568;
																assign node44568 = (inp[3]) ? 4'b0000 : 4'b0010;
										assign node44572 = (inp[5]) ? node44632 : node44573;
											assign node44573 = (inp[0]) ? node44605 : node44574;
												assign node44574 = (inp[15]) ? node44590 : node44575;
													assign node44575 = (inp[3]) ? node44583 : node44576;
														assign node44576 = (inp[9]) ? node44580 : node44577;
															assign node44577 = (inp[4]) ? 4'b1111 : 4'b1011;
															assign node44580 = (inp[4]) ? 4'b1011 : 4'b1111;
														assign node44583 = (inp[4]) ? node44587 : node44584;
															assign node44584 = (inp[12]) ? 4'b1011 : 4'b1101;
															assign node44587 = (inp[9]) ? 4'b1001 : 4'b1101;
													assign node44590 = (inp[3]) ? node44598 : node44591;
														assign node44591 = (inp[4]) ? node44595 : node44592;
															assign node44592 = (inp[9]) ? 4'b1101 : 4'b1001;
															assign node44595 = (inp[9]) ? 4'b1001 : 4'b1101;
														assign node44598 = (inp[9]) ? node44602 : node44599;
															assign node44599 = (inp[4]) ? 4'b1111 : 4'b1001;
															assign node44602 = (inp[4]) ? 4'b1011 : 4'b1111;
												assign node44605 = (inp[15]) ? node44615 : node44606;
													assign node44606 = (inp[3]) ? 4'b1111 : node44607;
														assign node44607 = (inp[9]) ? node44611 : node44608;
															assign node44608 = (inp[4]) ? 4'b1101 : 4'b1001;
															assign node44611 = (inp[4]) ? 4'b1001 : 4'b1101;
													assign node44615 = (inp[3]) ? node44625 : node44616;
														assign node44616 = (inp[12]) ? node44620 : node44617;
															assign node44617 = (inp[4]) ? 4'b1111 : 4'b1011;
															assign node44620 = (inp[4]) ? 4'b1011 : node44621;
																assign node44621 = (inp[9]) ? 4'b1111 : 4'b1011;
														assign node44625 = (inp[9]) ? node44629 : node44626;
															assign node44626 = (inp[4]) ? 4'b1101 : 4'b1011;
															assign node44629 = (inp[4]) ? 4'b1001 : 4'b1101;
											assign node44632 = (inp[9]) ? node44654 : node44633;
												assign node44633 = (inp[4]) ? node44647 : node44634;
													assign node44634 = (inp[15]) ? node44642 : node44635;
														assign node44635 = (inp[0]) ? node44639 : node44636;
															assign node44636 = (inp[3]) ? 4'b1001 : 4'b1011;
															assign node44639 = (inp[3]) ? 4'b1011 : 4'b1001;
														assign node44642 = (inp[0]) ? 4'b1001 : node44643;
															assign node44643 = (inp[3]) ? 4'b1011 : 4'b1001;
													assign node44647 = (inp[15]) ? node44651 : node44648;
														assign node44648 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node44651 = (inp[0]) ? 4'b1101 : 4'b1111;
												assign node44654 = (inp[4]) ? node44662 : node44655;
													assign node44655 = (inp[15]) ? node44659 : node44656;
														assign node44656 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node44659 = (inp[0]) ? 4'b1101 : 4'b1111;
													assign node44662 = (inp[15]) ? node44666 : node44663;
														assign node44663 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node44666 = (inp[0]) ? 4'b1001 : 4'b1011;
									assign node44669 = (inp[15]) ? node44769 : node44670;
										assign node44670 = (inp[0]) ? node44716 : node44671;
											assign node44671 = (inp[3]) ? node44695 : node44672;
												assign node44672 = (inp[5]) ? node44688 : node44673;
													assign node44673 = (inp[12]) ? node44681 : node44674;
														assign node44674 = (inp[4]) ? node44678 : node44675;
															assign node44675 = (inp[9]) ? 4'b1111 : 4'b1011;
															assign node44678 = (inp[9]) ? 4'b1011 : 4'b1111;
														assign node44681 = (inp[9]) ? node44685 : node44682;
															assign node44682 = (inp[4]) ? 4'b1111 : 4'b1011;
															assign node44685 = (inp[4]) ? 4'b1011 : 4'b1111;
													assign node44688 = (inp[4]) ? node44692 : node44689;
														assign node44689 = (inp[9]) ? 4'b1101 : 4'b1011;
														assign node44692 = (inp[9]) ? 4'b1001 : 4'b1101;
												assign node44695 = (inp[5]) ? node44703 : node44696;
													assign node44696 = (inp[9]) ? node44700 : node44697;
														assign node44697 = (inp[4]) ? 4'b1101 : 4'b1011;
														assign node44700 = (inp[4]) ? 4'b1001 : 4'b1101;
													assign node44703 = (inp[12]) ? node44709 : node44704;
														assign node44704 = (inp[4]) ? node44706 : 4'b1101;
															assign node44706 = (inp[14]) ? 4'b1001 : 4'b1101;
														assign node44709 = (inp[4]) ? node44713 : node44710;
															assign node44710 = (inp[9]) ? 4'b1101 : 4'b1001;
															assign node44713 = (inp[9]) ? 4'b1001 : 4'b1101;
											assign node44716 = (inp[5]) ? node44730 : node44717;
												assign node44717 = (inp[3]) ? node44723 : node44718;
													assign node44718 = (inp[9]) ? node44720 : 4'b1101;
														assign node44720 = (inp[4]) ? 4'b1001 : 4'b1101;
													assign node44723 = (inp[4]) ? node44727 : node44724;
														assign node44724 = (inp[9]) ? 4'b1111 : 4'b1001;
														assign node44727 = (inp[9]) ? 4'b1011 : 4'b1111;
												assign node44730 = (inp[3]) ? node44738 : node44731;
													assign node44731 = (inp[4]) ? node44735 : node44732;
														assign node44732 = (inp[9]) ? 4'b1111 : 4'b1001;
														assign node44735 = (inp[9]) ? 4'b1011 : 4'b1111;
													assign node44738 = (inp[12]) ? node44754 : node44739;
														assign node44739 = (inp[14]) ? node44747 : node44740;
															assign node44740 = (inp[4]) ? node44744 : node44741;
																assign node44741 = (inp[9]) ? 4'b1111 : 4'b1011;
																assign node44744 = (inp[9]) ? 4'b1011 : 4'b1111;
															assign node44747 = (inp[9]) ? node44751 : node44748;
																assign node44748 = (inp[4]) ? 4'b1111 : 4'b1011;
																assign node44751 = (inp[4]) ? 4'b1011 : 4'b1111;
														assign node44754 = (inp[14]) ? node44762 : node44755;
															assign node44755 = (inp[9]) ? node44759 : node44756;
																assign node44756 = (inp[4]) ? 4'b1111 : 4'b1011;
																assign node44759 = (inp[4]) ? 4'b1011 : 4'b1111;
															assign node44762 = (inp[4]) ? node44766 : node44763;
																assign node44763 = (inp[9]) ? 4'b1111 : 4'b1011;
																assign node44766 = (inp[9]) ? 4'b1011 : 4'b1111;
										assign node44769 = (inp[0]) ? node44807 : node44770;
											assign node44770 = (inp[3]) ? node44792 : node44771;
												assign node44771 = (inp[5]) ? node44785 : node44772;
													assign node44772 = (inp[12]) ? node44780 : node44773;
														assign node44773 = (inp[9]) ? node44777 : node44774;
															assign node44774 = (inp[4]) ? 4'b1101 : 4'b1001;
															assign node44777 = (inp[4]) ? 4'b1001 : 4'b1101;
														assign node44780 = (inp[9]) ? node44782 : 4'b1001;
															assign node44782 = (inp[4]) ? 4'b1001 : 4'b1101;
													assign node44785 = (inp[9]) ? node44789 : node44786;
														assign node44786 = (inp[4]) ? 4'b1111 : 4'b1001;
														assign node44789 = (inp[4]) ? 4'b1011 : 4'b1111;
												assign node44792 = (inp[5]) ? node44800 : node44793;
													assign node44793 = (inp[9]) ? node44797 : node44794;
														assign node44794 = (inp[4]) ? 4'b1111 : 4'b1001;
														assign node44797 = (inp[4]) ? 4'b1011 : 4'b1111;
													assign node44800 = (inp[9]) ? node44804 : node44801;
														assign node44801 = (inp[4]) ? 4'b1111 : 4'b1011;
														assign node44804 = (inp[4]) ? 4'b1011 : 4'b1111;
											assign node44807 = (inp[3]) ? node44827 : node44808;
												assign node44808 = (inp[5]) ? node44820 : node44809;
													assign node44809 = (inp[12]) ? node44815 : node44810;
														assign node44810 = (inp[4]) ? 4'b1111 : node44811;
															assign node44811 = (inp[9]) ? 4'b1111 : 4'b1011;
														assign node44815 = (inp[4]) ? node44817 : 4'b1111;
															assign node44817 = (inp[14]) ? 4'b1111 : 4'b1011;
													assign node44820 = (inp[4]) ? node44824 : node44821;
														assign node44821 = (inp[9]) ? 4'b1101 : 4'b1011;
														assign node44824 = (inp[9]) ? 4'b1001 : 4'b1101;
												assign node44827 = (inp[5]) ? node44835 : node44828;
													assign node44828 = (inp[9]) ? node44832 : node44829;
														assign node44829 = (inp[4]) ? 4'b1101 : 4'b1011;
														assign node44832 = (inp[4]) ? 4'b1001 : 4'b1101;
													assign node44835 = (inp[12]) ? node44851 : node44836;
														assign node44836 = (inp[14]) ? node44844 : node44837;
															assign node44837 = (inp[4]) ? node44841 : node44838;
																assign node44838 = (inp[9]) ? 4'b1101 : 4'b1001;
																assign node44841 = (inp[9]) ? 4'b1001 : 4'b1101;
															assign node44844 = (inp[4]) ? node44848 : node44845;
																assign node44845 = (inp[9]) ? 4'b1101 : 4'b1001;
																assign node44848 = (inp[9]) ? 4'b1001 : 4'b1101;
														assign node44851 = (inp[9]) ? node44855 : node44852;
															assign node44852 = (inp[4]) ? 4'b1101 : 4'b1001;
															assign node44855 = (inp[4]) ? 4'b1001 : 4'b1101;
							assign node44858 = (inp[7]) ? node45324 : node44859;
								assign node44859 = (inp[14]) ? node45117 : node44860;
									assign node44860 = (inp[2]) ? node44986 : node44861;
										assign node44861 = (inp[15]) ? node44921 : node44862;
											assign node44862 = (inp[0]) ? node44898 : node44863;
												assign node44863 = (inp[5]) ? node44881 : node44864;
													assign node44864 = (inp[3]) ? node44868 : node44865;
														assign node44865 = (inp[9]) ? 4'b0010 : 4'b0110;
														assign node44868 = (inp[4]) ? node44874 : node44869;
															assign node44869 = (inp[9]) ? node44871 : 4'b0010;
																assign node44871 = (inp[12]) ? 4'b0100 : 4'b0010;
															assign node44874 = (inp[9]) ? node44878 : node44875;
																assign node44875 = (inp[12]) ? 4'b0100 : 4'b0010;
																assign node44878 = (inp[12]) ? 4'b0000 : 4'b0100;
													assign node44881 = (inp[3]) ? node44893 : node44882;
														assign node44882 = (inp[4]) ? node44888 : node44883;
															assign node44883 = (inp[12]) ? 4'b0100 : node44884;
																assign node44884 = (inp[9]) ? 4'b0010 : 4'b0110;
															assign node44888 = (inp[9]) ? node44890 : 4'b0100;
																assign node44890 = (inp[12]) ? 4'b0000 : 4'b0100;
														assign node44893 = (inp[4]) ? 4'b0000 : node44894;
															assign node44894 = (inp[9]) ? 4'b0000 : 4'b0100;
												assign node44898 = (inp[5]) ? node44908 : node44899;
													assign node44899 = (inp[3]) ? node44901 : 4'b0000;
														assign node44901 = (inp[12]) ? 4'b0010 : node44902;
															assign node44902 = (inp[9]) ? node44904 : 4'b0000;
																assign node44904 = (inp[4]) ? 4'b0110 : 4'b0000;
													assign node44908 = (inp[12]) ? node44916 : node44909;
														assign node44909 = (inp[9]) ? node44913 : node44910;
															assign node44910 = (inp[3]) ? 4'b0010 : 4'b0000;
															assign node44913 = (inp[4]) ? 4'b0110 : 4'b0010;
														assign node44916 = (inp[4]) ? node44918 : 4'b0110;
															assign node44918 = (inp[9]) ? 4'b0010 : 4'b0110;
											assign node44921 = (inp[9]) ? node44959 : node44922;
												assign node44922 = (inp[0]) ? node44944 : node44923;
													assign node44923 = (inp[3]) ? node44933 : node44924;
														assign node44924 = (inp[5]) ? 4'b0000 : node44925;
															assign node44925 = (inp[12]) ? node44929 : node44926;
																assign node44926 = (inp[4]) ? 4'b0000 : 4'b0100;
																assign node44929 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node44933 = (inp[5]) ? node44941 : node44934;
															assign node44934 = (inp[12]) ? node44938 : node44935;
																assign node44935 = (inp[4]) ? 4'b0000 : 4'b0100;
																assign node44938 = (inp[4]) ? 4'b0110 : 4'b0000;
															assign node44941 = (inp[4]) ? 4'b0010 : 4'b0110;
													assign node44944 = (inp[3]) ? node44952 : node44945;
														assign node44945 = (inp[5]) ? node44949 : node44946;
															assign node44946 = (inp[4]) ? 4'b0110 : 4'b0010;
															assign node44949 = (inp[4]) ? 4'b0010 : 4'b0110;
														assign node44952 = (inp[5]) ? 4'b0100 : node44953;
															assign node44953 = (inp[4]) ? node44955 : 4'b0010;
																assign node44955 = (inp[12]) ? 4'b0100 : 4'b0010;
												assign node44959 = (inp[0]) ? node44973 : node44960;
													assign node44960 = (inp[3]) ? node44968 : node44961;
														assign node44961 = (inp[12]) ? node44965 : node44962;
															assign node44962 = (inp[4]) ? 4'b0100 : 4'b0000;
															assign node44965 = (inp[5]) ? 4'b0110 : 4'b0100;
														assign node44968 = (inp[4]) ? node44970 : 4'b0110;
															assign node44970 = (inp[12]) ? 4'b0010 : 4'b0110;
													assign node44973 = (inp[5]) ? node44977 : node44974;
														assign node44974 = (inp[3]) ? 4'b0100 : 4'b0110;
														assign node44977 = (inp[3]) ? node44979 : 4'b0000;
															assign node44979 = (inp[4]) ? node44983 : node44980;
																assign node44980 = (inp[12]) ? 4'b0100 : 4'b0000;
																assign node44983 = (inp[12]) ? 4'b0000 : 4'b0100;
										assign node44986 = (inp[4]) ? node45056 : node44987;
											assign node44987 = (inp[9]) ? node45017 : node44988;
												assign node44988 = (inp[3]) ? node45002 : node44989;
													assign node44989 = (inp[12]) ? node44997 : node44990;
														assign node44990 = (inp[0]) ? node44994 : node44991;
															assign node44991 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node44994 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node44997 = (inp[0]) ? 4'b1001 : node44998;
															assign node44998 = (inp[15]) ? 4'b1001 : 4'b1011;
													assign node45002 = (inp[15]) ? 4'b1011 : node45003;
														assign node45003 = (inp[12]) ? node45011 : node45004;
															assign node45004 = (inp[0]) ? node45008 : node45005;
																assign node45005 = (inp[5]) ? 4'b1001 : 4'b1011;
																assign node45008 = (inp[5]) ? 4'b1011 : 4'b1001;
															assign node45011 = (inp[0]) ? 4'b1011 : node45012;
																assign node45012 = (inp[5]) ? 4'b1001 : 4'b1011;
												assign node45017 = (inp[5]) ? node45035 : node45018;
													assign node45018 = (inp[0]) ? node45024 : node45019;
														assign node45019 = (inp[15]) ? 4'b1111 : node45020;
															assign node45020 = (inp[3]) ? 4'b1101 : 4'b1111;
														assign node45024 = (inp[12]) ? node45030 : node45025;
															assign node45025 = (inp[3]) ? node45027 : 4'b1101;
																assign node45027 = (inp[15]) ? 4'b1101 : 4'b1111;
															assign node45030 = (inp[15]) ? 4'b1111 : node45031;
																assign node45031 = (inp[3]) ? 4'b1111 : 4'b1101;
													assign node45035 = (inp[3]) ? node45043 : node45036;
														assign node45036 = (inp[15]) ? node45040 : node45037;
															assign node45037 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node45040 = (inp[0]) ? 4'b1101 : 4'b1111;
														assign node45043 = (inp[12]) ? node45051 : node45044;
															assign node45044 = (inp[15]) ? node45048 : node45045;
																assign node45045 = (inp[0]) ? 4'b1111 : 4'b1101;
																assign node45048 = (inp[0]) ? 4'b1101 : 4'b1111;
															assign node45051 = (inp[0]) ? node45053 : 4'b1101;
																assign node45053 = (inp[15]) ? 4'b1101 : 4'b1111;
											assign node45056 = (inp[9]) ? node45094 : node45057;
												assign node45057 = (inp[3]) ? node45085 : node45058;
													assign node45058 = (inp[12]) ? node45072 : node45059;
														assign node45059 = (inp[0]) ? node45065 : node45060;
															assign node45060 = (inp[15]) ? node45062 : 4'b1101;
																assign node45062 = (inp[5]) ? 4'b1111 : 4'b1101;
															assign node45065 = (inp[15]) ? node45069 : node45066;
																assign node45066 = (inp[5]) ? 4'b1111 : 4'b1101;
																assign node45069 = (inp[5]) ? 4'b1101 : 4'b1111;
														assign node45072 = (inp[5]) ? node45080 : node45073;
															assign node45073 = (inp[15]) ? node45077 : node45074;
																assign node45074 = (inp[0]) ? 4'b1101 : 4'b1111;
																assign node45077 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node45080 = (inp[15]) ? 4'b1111 : node45081;
																assign node45081 = (inp[0]) ? 4'b1111 : 4'b1101;
													assign node45085 = (inp[5]) ? 4'b1101 : node45086;
														assign node45086 = (inp[0]) ? node45090 : node45087;
															assign node45087 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node45090 = (inp[15]) ? 4'b1101 : 4'b1111;
												assign node45094 = (inp[15]) ? node45106 : node45095;
													assign node45095 = (inp[0]) ? node45101 : node45096;
														assign node45096 = (inp[5]) ? 4'b1001 : node45097;
															assign node45097 = (inp[12]) ? 4'b1011 : 4'b1001;
														assign node45101 = (inp[5]) ? 4'b1011 : node45102;
															assign node45102 = (inp[3]) ? 4'b1011 : 4'b1001;
													assign node45106 = (inp[0]) ? node45110 : node45107;
														assign node45107 = (inp[5]) ? 4'b1011 : 4'b1001;
														assign node45110 = (inp[12]) ? node45112 : 4'b1001;
															assign node45112 = (inp[5]) ? 4'b1001 : node45113;
																assign node45113 = (inp[3]) ? 4'b1001 : 4'b1011;
									assign node45117 = (inp[2]) ? node45213 : node45118;
										assign node45118 = (inp[4]) ? node45160 : node45119;
											assign node45119 = (inp[9]) ? node45141 : node45120;
												assign node45120 = (inp[3]) ? node45128 : node45121;
													assign node45121 = (inp[15]) ? node45125 : node45122;
														assign node45122 = (inp[0]) ? 4'b1001 : 4'b1011;
														assign node45125 = (inp[0]) ? 4'b1011 : 4'b1001;
													assign node45128 = (inp[15]) ? node45134 : node45129;
														assign node45129 = (inp[12]) ? 4'b1001 : node45130;
															assign node45130 = (inp[5]) ? 4'b1011 : 4'b1001;
														assign node45134 = (inp[5]) ? node45138 : node45135;
															assign node45135 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node45138 = (inp[0]) ? 4'b1001 : 4'b1011;
												assign node45141 = (inp[15]) ? node45151 : node45142;
													assign node45142 = (inp[0]) ? node45148 : node45143;
														assign node45143 = (inp[3]) ? 4'b1101 : node45144;
															assign node45144 = (inp[5]) ? 4'b1101 : 4'b1111;
														assign node45148 = (inp[5]) ? 4'b1111 : 4'b1101;
													assign node45151 = (inp[0]) ? node45157 : node45152;
														assign node45152 = (inp[5]) ? 4'b1111 : node45153;
															assign node45153 = (inp[3]) ? 4'b1111 : 4'b1101;
														assign node45157 = (inp[5]) ? 4'b1101 : 4'b1111;
											assign node45160 = (inp[9]) ? node45184 : node45161;
												assign node45161 = (inp[15]) ? node45173 : node45162;
													assign node45162 = (inp[0]) ? node45168 : node45163;
														assign node45163 = (inp[5]) ? 4'b1101 : node45164;
															assign node45164 = (inp[3]) ? 4'b1101 : 4'b1111;
														assign node45168 = (inp[3]) ? 4'b1111 : node45169;
															assign node45169 = (inp[5]) ? 4'b1111 : 4'b1101;
													assign node45173 = (inp[0]) ? node45179 : node45174;
														assign node45174 = (inp[5]) ? 4'b1111 : node45175;
															assign node45175 = (inp[3]) ? 4'b1111 : 4'b1101;
														assign node45179 = (inp[3]) ? 4'b1101 : node45180;
															assign node45180 = (inp[5]) ? 4'b1101 : 4'b1111;
												assign node45184 = (inp[5]) ? node45200 : node45185;
													assign node45185 = (inp[3]) ? node45193 : node45186;
														assign node45186 = (inp[0]) ? node45190 : node45187;
															assign node45187 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node45190 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node45193 = (inp[15]) ? node45197 : node45194;
															assign node45194 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node45197 = (inp[0]) ? 4'b1001 : 4'b1011;
													assign node45200 = (inp[12]) ? node45208 : node45201;
														assign node45201 = (inp[15]) ? node45205 : node45202;
															assign node45202 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node45205 = (inp[0]) ? 4'b1001 : 4'b1011;
														assign node45208 = (inp[15]) ? node45210 : 4'b1001;
															assign node45210 = (inp[0]) ? 4'b1001 : 4'b1011;
										assign node45213 = (inp[5]) ? node45283 : node45214;
											assign node45214 = (inp[0]) ? node45254 : node45215;
												assign node45215 = (inp[15]) ? node45239 : node45216;
													assign node45216 = (inp[3]) ? node45232 : node45217;
														assign node45217 = (inp[12]) ? node45225 : node45218;
															assign node45218 = (inp[4]) ? node45222 : node45219;
																assign node45219 = (inp[9]) ? 4'b1111 : 4'b1011;
																assign node45222 = (inp[9]) ? 4'b1011 : 4'b1111;
															assign node45225 = (inp[4]) ? node45229 : node45226;
																assign node45226 = (inp[9]) ? 4'b1111 : 4'b1011;
																assign node45229 = (inp[9]) ? 4'b1011 : 4'b1111;
														assign node45232 = (inp[4]) ? node45236 : node45233;
															assign node45233 = (inp[9]) ? 4'b1101 : 4'b1011;
															assign node45236 = (inp[9]) ? 4'b1001 : 4'b1101;
													assign node45239 = (inp[3]) ? node45247 : node45240;
														assign node45240 = (inp[4]) ? node45244 : node45241;
															assign node45241 = (inp[9]) ? 4'b1101 : 4'b1001;
															assign node45244 = (inp[9]) ? 4'b1001 : 4'b1101;
														assign node45247 = (inp[4]) ? node45251 : node45248;
															assign node45248 = (inp[9]) ? 4'b1111 : 4'b1001;
															assign node45251 = (inp[9]) ? 4'b1011 : 4'b1111;
												assign node45254 = (inp[12]) ? node45272 : node45255;
													assign node45255 = (inp[9]) ? node45261 : node45256;
														assign node45256 = (inp[4]) ? 4'b1111 : node45257;
															assign node45257 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node45261 = (inp[4]) ? node45269 : node45262;
															assign node45262 = (inp[3]) ? node45266 : node45263;
																assign node45263 = (inp[15]) ? 4'b1111 : 4'b1101;
																assign node45266 = (inp[15]) ? 4'b1101 : 4'b1111;
															assign node45269 = (inp[3]) ? 4'b1011 : 4'b1001;
													assign node45272 = (inp[4]) ? node45276 : node45273;
														assign node45273 = (inp[9]) ? 4'b1101 : 4'b1001;
														assign node45276 = (inp[9]) ? node45278 : 4'b1101;
															assign node45278 = (inp[15]) ? node45280 : 4'b1001;
																assign node45280 = (inp[3]) ? 4'b1001 : 4'b1011;
											assign node45283 = (inp[4]) ? node45303 : node45284;
												assign node45284 = (inp[9]) ? node45298 : node45285;
													assign node45285 = (inp[0]) ? node45291 : node45286;
														assign node45286 = (inp[15]) ? node45288 : 4'b1011;
															assign node45288 = (inp[3]) ? 4'b1011 : 4'b1001;
														assign node45291 = (inp[15]) ? node45295 : node45292;
															assign node45292 = (inp[3]) ? 4'b1011 : 4'b1001;
															assign node45295 = (inp[3]) ? 4'b1001 : 4'b1011;
													assign node45298 = (inp[15]) ? 4'b1111 : node45299;
														assign node45299 = (inp[0]) ? 4'b1111 : 4'b1101;
												assign node45303 = (inp[9]) ? node45309 : node45304;
													assign node45304 = (inp[15]) ? 4'b1101 : node45305;
														assign node45305 = (inp[0]) ? 4'b1111 : 4'b1101;
													assign node45309 = (inp[3]) ? node45317 : node45310;
														assign node45310 = (inp[15]) ? node45314 : node45311;
															assign node45311 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node45314 = (inp[0]) ? 4'b1001 : 4'b1011;
														assign node45317 = (inp[0]) ? node45321 : node45318;
															assign node45318 = (inp[15]) ? 4'b1011 : 4'b1001;
															assign node45321 = (inp[12]) ? 4'b1011 : 4'b1001;
								assign node45324 = (inp[2]) ? node45572 : node45325;
									assign node45325 = (inp[14]) ? node45465 : node45326;
										assign node45326 = (inp[3]) ? node45386 : node45327;
											assign node45327 = (inp[15]) ? node45355 : node45328;
												assign node45328 = (inp[9]) ? node45338 : node45329;
													assign node45329 = (inp[4]) ? node45333 : node45330;
														assign node45330 = (inp[0]) ? 4'b1001 : 4'b1011;
														assign node45333 = (inp[12]) ? node45335 : 4'b1101;
															assign node45335 = (inp[0]) ? 4'b1111 : 4'b1101;
													assign node45338 = (inp[4]) ? node45348 : node45339;
														assign node45339 = (inp[12]) ? 4'b1111 : node45340;
															assign node45340 = (inp[5]) ? node45344 : node45341;
																assign node45341 = (inp[0]) ? 4'b1101 : 4'b1111;
																assign node45344 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node45348 = (inp[5]) ? node45352 : node45349;
															assign node45349 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node45352 = (inp[0]) ? 4'b1011 : 4'b1001;
												assign node45355 = (inp[9]) ? node45373 : node45356;
													assign node45356 = (inp[4]) ? node45360 : node45357;
														assign node45357 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node45360 = (inp[12]) ? node45366 : node45361;
															assign node45361 = (inp[5]) ? node45363 : 4'b1111;
																assign node45363 = (inp[0]) ? 4'b1101 : 4'b1111;
															assign node45366 = (inp[5]) ? node45370 : node45367;
																assign node45367 = (inp[0]) ? 4'b1111 : 4'b1101;
																assign node45370 = (inp[0]) ? 4'b1101 : 4'b1111;
													assign node45373 = (inp[4]) ? node45379 : node45374;
														assign node45374 = (inp[0]) ? 4'b1111 : node45375;
															assign node45375 = (inp[5]) ? 4'b1111 : 4'b1101;
														assign node45379 = (inp[5]) ? node45383 : node45380;
															assign node45380 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node45383 = (inp[0]) ? 4'b1001 : 4'b1011;
											assign node45386 = (inp[12]) ? node45420 : node45387;
												assign node45387 = (inp[9]) ? node45407 : node45388;
													assign node45388 = (inp[4]) ? node45394 : node45389;
														assign node45389 = (inp[15]) ? 4'b1011 : node45390;
															assign node45390 = (inp[0]) ? 4'b1001 : 4'b1011;
														assign node45394 = (inp[5]) ? node45402 : node45395;
															assign node45395 = (inp[0]) ? node45399 : node45396;
																assign node45396 = (inp[15]) ? 4'b1111 : 4'b1101;
																assign node45399 = (inp[15]) ? 4'b1101 : 4'b1111;
															assign node45402 = (inp[15]) ? node45404 : 4'b1111;
																assign node45404 = (inp[0]) ? 4'b1101 : 4'b1111;
													assign node45407 = (inp[4]) ? node45413 : node45408;
														assign node45408 = (inp[0]) ? 4'b1111 : node45409;
															assign node45409 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node45413 = (inp[15]) ? node45417 : node45414;
															assign node45414 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node45417 = (inp[0]) ? 4'b1001 : 4'b1011;
												assign node45420 = (inp[4]) ? node45448 : node45421;
													assign node45421 = (inp[9]) ? node45435 : node45422;
														assign node45422 = (inp[15]) ? node45430 : node45423;
															assign node45423 = (inp[5]) ? node45427 : node45424;
																assign node45424 = (inp[0]) ? 4'b1001 : 4'b1011;
																assign node45427 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node45430 = (inp[5]) ? 4'b1001 : node45431;
																assign node45431 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node45435 = (inp[5]) ? node45441 : node45436;
															assign node45436 = (inp[0]) ? node45438 : 4'b1101;
																assign node45438 = (inp[15]) ? 4'b1101 : 4'b1111;
															assign node45441 = (inp[0]) ? node45445 : node45442;
																assign node45442 = (inp[15]) ? 4'b1111 : 4'b1101;
																assign node45445 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node45448 = (inp[9]) ? node45462 : node45449;
														assign node45449 = (inp[5]) ? node45457 : node45450;
															assign node45450 = (inp[15]) ? node45454 : node45451;
																assign node45451 = (inp[0]) ? 4'b1111 : 4'b1101;
																assign node45454 = (inp[0]) ? 4'b1101 : 4'b1111;
															assign node45457 = (inp[0]) ? 4'b1111 : node45458;
																assign node45458 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node45462 = (inp[15]) ? 4'b1011 : 4'b1001;
										assign node45465 = (inp[0]) ? node45533 : node45466;
											assign node45466 = (inp[15]) ? node45502 : node45467;
												assign node45467 = (inp[3]) ? node45487 : node45468;
													assign node45468 = (inp[5]) ? node45480 : node45469;
														assign node45469 = (inp[12]) ? node45475 : node45470;
															assign node45470 = (inp[9]) ? 4'b1010 : node45471;
																assign node45471 = (inp[4]) ? 4'b1110 : 4'b1010;
															assign node45475 = (inp[4]) ? 4'b1010 : node45476;
																assign node45476 = (inp[9]) ? 4'b1110 : 4'b1010;
														assign node45480 = (inp[9]) ? node45484 : node45481;
															assign node45481 = (inp[4]) ? 4'b1100 : 4'b1010;
															assign node45484 = (inp[4]) ? 4'b1000 : 4'b1100;
													assign node45487 = (inp[12]) ? node45495 : node45488;
														assign node45488 = (inp[5]) ? node45490 : 4'b1100;
															assign node45490 = (inp[9]) ? 4'b1000 : node45491;
																assign node45491 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node45495 = (inp[9]) ? node45499 : node45496;
															assign node45496 = (inp[5]) ? 4'b1000 : 4'b1010;
															assign node45499 = (inp[4]) ? 4'b1000 : 4'b1100;
												assign node45502 = (inp[5]) ? node45518 : node45503;
													assign node45503 = (inp[3]) ? node45513 : node45504;
														assign node45504 = (inp[12]) ? node45506 : 4'b1000;
															assign node45506 = (inp[4]) ? node45510 : node45507;
																assign node45507 = (inp[9]) ? 4'b1100 : 4'b1000;
																assign node45510 = (inp[9]) ? 4'b1000 : 4'b1100;
														assign node45513 = (inp[4]) ? node45515 : 4'b1000;
															assign node45515 = (inp[9]) ? 4'b1010 : 4'b1110;
													assign node45518 = (inp[3]) ? node45526 : node45519;
														assign node45519 = (inp[12]) ? node45521 : 4'b1110;
															assign node45521 = (inp[4]) ? node45523 : 4'b1000;
																assign node45523 = (inp[9]) ? 4'b1010 : 4'b1110;
														assign node45526 = (inp[9]) ? node45530 : node45527;
															assign node45527 = (inp[4]) ? 4'b1110 : 4'b1010;
															assign node45530 = (inp[4]) ? 4'b1010 : 4'b1110;
											assign node45533 = (inp[9]) ? node45551 : node45534;
												assign node45534 = (inp[4]) ? node45540 : node45535;
													assign node45535 = (inp[15]) ? node45537 : 4'b1000;
														assign node45537 = (inp[5]) ? 4'b1000 : 4'b1010;
													assign node45540 = (inp[15]) ? node45546 : node45541;
														assign node45541 = (inp[12]) ? node45543 : 4'b1110;
															assign node45543 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node45546 = (inp[3]) ? 4'b1100 : node45547;
															assign node45547 = (inp[12]) ? 4'b1100 : 4'b1110;
												assign node45551 = (inp[4]) ? node45561 : node45552;
													assign node45552 = (inp[15]) ? node45558 : node45553;
														assign node45553 = (inp[3]) ? 4'b1110 : node45554;
															assign node45554 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node45558 = (inp[3]) ? 4'b1100 : 4'b1110;
													assign node45561 = (inp[15]) ? node45567 : node45562;
														assign node45562 = (inp[5]) ? 4'b1010 : node45563;
															assign node45563 = (inp[3]) ? 4'b1010 : 4'b1000;
														assign node45567 = (inp[3]) ? 4'b1000 : node45568;
															assign node45568 = (inp[5]) ? 4'b1000 : 4'b1010;
									assign node45572 = (inp[9]) ? node45652 : node45573;
										assign node45573 = (inp[4]) ? node45629 : node45574;
											assign node45574 = (inp[3]) ? node45600 : node45575;
												assign node45575 = (inp[12]) ? node45593 : node45576;
													assign node45576 = (inp[5]) ? node45584 : node45577;
														assign node45577 = (inp[0]) ? node45581 : node45578;
															assign node45578 = (inp[15]) ? 4'b1000 : 4'b1010;
															assign node45581 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node45584 = (inp[14]) ? 4'b1010 : node45585;
															assign node45585 = (inp[0]) ? node45589 : node45586;
																assign node45586 = (inp[15]) ? 4'b1000 : 4'b1010;
																assign node45589 = (inp[15]) ? 4'b1010 : 4'b1000;
													assign node45593 = (inp[0]) ? node45597 : node45594;
														assign node45594 = (inp[15]) ? 4'b1000 : 4'b1010;
														assign node45597 = (inp[15]) ? 4'b1010 : 4'b1000;
												assign node45600 = (inp[12]) ? node45616 : node45601;
													assign node45601 = (inp[5]) ? node45609 : node45602;
														assign node45602 = (inp[15]) ? node45606 : node45603;
															assign node45603 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node45606 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node45609 = (inp[0]) ? node45613 : node45610;
															assign node45610 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node45613 = (inp[15]) ? 4'b1000 : 4'b1010;
													assign node45616 = (inp[15]) ? node45624 : node45617;
														assign node45617 = (inp[5]) ? node45621 : node45618;
															assign node45618 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node45621 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node45624 = (inp[14]) ? 4'b1010 : node45625;
															assign node45625 = (inp[5]) ? 4'b1000 : 4'b1010;
											assign node45629 = (inp[0]) ? node45641 : node45630;
												assign node45630 = (inp[15]) ? node45636 : node45631;
													assign node45631 = (inp[5]) ? 4'b1100 : node45632;
														assign node45632 = (inp[3]) ? 4'b1100 : 4'b1110;
													assign node45636 = (inp[5]) ? 4'b1110 : node45637;
														assign node45637 = (inp[3]) ? 4'b1110 : 4'b1100;
												assign node45641 = (inp[15]) ? node45647 : node45642;
													assign node45642 = (inp[3]) ? 4'b1110 : node45643;
														assign node45643 = (inp[5]) ? 4'b1110 : 4'b1100;
													assign node45647 = (inp[3]) ? 4'b1100 : node45648;
														assign node45648 = (inp[5]) ? 4'b1100 : 4'b1110;
										assign node45652 = (inp[4]) ? node45702 : node45653;
											assign node45653 = (inp[5]) ? node45675 : node45654;
												assign node45654 = (inp[3]) ? node45664 : node45655;
													assign node45655 = (inp[12]) ? node45657 : 4'b1110;
														assign node45657 = (inp[15]) ? node45661 : node45658;
															assign node45658 = (inp[0]) ? 4'b1100 : 4'b1110;
															assign node45661 = (inp[0]) ? 4'b1110 : 4'b1100;
													assign node45664 = (inp[14]) ? node45670 : node45665;
														assign node45665 = (inp[0]) ? node45667 : 4'b1110;
															assign node45667 = (inp[15]) ? 4'b1100 : 4'b1110;
														assign node45670 = (inp[0]) ? node45672 : 4'b1100;
															assign node45672 = (inp[15]) ? 4'b1100 : 4'b1110;
												assign node45675 = (inp[12]) ? node45691 : node45676;
													assign node45676 = (inp[14]) ? node45682 : node45677;
														assign node45677 = (inp[15]) ? node45679 : 4'b1100;
															assign node45679 = (inp[0]) ? 4'b1100 : 4'b1110;
														assign node45682 = (inp[3]) ? node45688 : node45683;
															assign node45683 = (inp[0]) ? node45685 : 4'b1100;
																assign node45685 = (inp[15]) ? 4'b1100 : 4'b1110;
															assign node45688 = (inp[15]) ? 4'b1110 : 4'b1100;
													assign node45691 = (inp[3]) ? node45697 : node45692;
														assign node45692 = (inp[0]) ? node45694 : 4'b1110;
															assign node45694 = (inp[15]) ? 4'b1100 : 4'b1110;
														assign node45697 = (inp[15]) ? 4'b1110 : node45698;
															assign node45698 = (inp[0]) ? 4'b1110 : 4'b1100;
											assign node45702 = (inp[12]) ? node45732 : node45703;
												assign node45703 = (inp[14]) ? node45723 : node45704;
													assign node45704 = (inp[0]) ? node45716 : node45705;
														assign node45705 = (inp[15]) ? node45711 : node45706;
															assign node45706 = (inp[5]) ? 4'b1000 : node45707;
																assign node45707 = (inp[3]) ? 4'b1000 : 4'b1010;
															assign node45711 = (inp[5]) ? 4'b1010 : node45712;
																assign node45712 = (inp[3]) ? 4'b1010 : 4'b1000;
														assign node45716 = (inp[15]) ? node45718 : 4'b1010;
															assign node45718 = (inp[3]) ? 4'b1000 : node45719;
																assign node45719 = (inp[5]) ? 4'b1000 : 4'b1010;
													assign node45723 = (inp[3]) ? node45725 : 4'b1010;
														assign node45725 = (inp[0]) ? node45729 : node45726;
															assign node45726 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node45729 = (inp[15]) ? 4'b1000 : 4'b1010;
												assign node45732 = (inp[0]) ? node45738 : node45733;
													assign node45733 = (inp[15]) ? 4'b1010 : node45734;
														assign node45734 = (inp[5]) ? 4'b1000 : 4'b1010;
													assign node45738 = (inp[15]) ? node45744 : node45739;
														assign node45739 = (inp[5]) ? 4'b1010 : node45740;
															assign node45740 = (inp[3]) ? 4'b1010 : 4'b1000;
														assign node45744 = (inp[3]) ? 4'b1000 : node45745;
															assign node45745 = (inp[5]) ? 4'b1000 : 4'b1010;
						assign node45749 = (inp[4]) ? node46613 : node45750;
							assign node45750 = (inp[9]) ? node46170 : node45751;
								assign node45751 = (inp[2]) ? node45983 : node45752;
									assign node45752 = (inp[0]) ? node45858 : node45753;
										assign node45753 = (inp[15]) ? node45815 : node45754;
											assign node45754 = (inp[3]) ? node45778 : node45755;
												assign node45755 = (inp[7]) ? node45763 : node45756;
													assign node45756 = (inp[14]) ? node45760 : node45757;
														assign node45757 = (inp[8]) ? 4'b1010 : 4'b1011;
														assign node45760 = (inp[8]) ? 4'b1011 : 4'b1010;
													assign node45763 = (inp[12]) ? node45771 : node45764;
														assign node45764 = (inp[8]) ? node45768 : node45765;
															assign node45765 = (inp[14]) ? 4'b1011 : 4'b1010;
															assign node45768 = (inp[14]) ? 4'b1010 : 4'b1011;
														assign node45771 = (inp[8]) ? node45775 : node45772;
															assign node45772 = (inp[14]) ? 4'b1011 : 4'b1010;
															assign node45775 = (inp[14]) ? 4'b1010 : 4'b1011;
												assign node45778 = (inp[5]) ? node45796 : node45779;
													assign node45779 = (inp[12]) ? node45785 : node45780;
														assign node45780 = (inp[14]) ? node45782 : 4'b1010;
															assign node45782 = (inp[7]) ? 4'b1010 : 4'b1011;
														assign node45785 = (inp[8]) ? node45791 : node45786;
															assign node45786 = (inp[7]) ? node45788 : 4'b1011;
																assign node45788 = (inp[14]) ? 4'b1011 : 4'b1010;
															assign node45791 = (inp[7]) ? node45793 : 4'b1010;
																assign node45793 = (inp[14]) ? 4'b1010 : 4'b1011;
													assign node45796 = (inp[12]) ? node45806 : node45797;
														assign node45797 = (inp[14]) ? 4'b1000 : node45798;
															assign node45798 = (inp[7]) ? node45802 : node45799;
																assign node45799 = (inp[8]) ? 4'b1000 : 4'b1001;
																assign node45802 = (inp[8]) ? 4'b1001 : 4'b1000;
														assign node45806 = (inp[14]) ? node45808 : 4'b1001;
															assign node45808 = (inp[7]) ? node45812 : node45809;
																assign node45809 = (inp[8]) ? 4'b1001 : 4'b1000;
																assign node45812 = (inp[8]) ? 4'b1000 : 4'b1001;
											assign node45815 = (inp[3]) ? node45833 : node45816;
												assign node45816 = (inp[8]) ? node45824 : node45817;
													assign node45817 = (inp[14]) ? node45821 : node45818;
														assign node45818 = (inp[7]) ? 4'b1000 : 4'b1001;
														assign node45821 = (inp[7]) ? 4'b1001 : 4'b1000;
													assign node45824 = (inp[12]) ? node45826 : 4'b1000;
														assign node45826 = (inp[14]) ? node45830 : node45827;
															assign node45827 = (inp[7]) ? 4'b1001 : 4'b1000;
															assign node45830 = (inp[5]) ? 4'b1001 : 4'b1000;
												assign node45833 = (inp[5]) ? node45849 : node45834;
													assign node45834 = (inp[7]) ? node45844 : node45835;
														assign node45835 = (inp[12]) ? node45841 : node45836;
															assign node45836 = (inp[14]) ? 4'b1001 : node45837;
																assign node45837 = (inp[8]) ? 4'b1000 : 4'b1001;
															assign node45841 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node45844 = (inp[14]) ? 4'b1000 : node45845;
															assign node45845 = (inp[8]) ? 4'b1001 : 4'b1000;
													assign node45849 = (inp[8]) ? 4'b1010 : node45850;
														assign node45850 = (inp[7]) ? node45854 : node45851;
															assign node45851 = (inp[14]) ? 4'b1010 : 4'b1011;
															assign node45854 = (inp[14]) ? 4'b1011 : 4'b1010;
										assign node45858 = (inp[15]) ? node45936 : node45859;
											assign node45859 = (inp[3]) ? node45899 : node45860;
												assign node45860 = (inp[12]) ? node45882 : node45861;
													assign node45861 = (inp[8]) ? node45867 : node45862;
														assign node45862 = (inp[7]) ? node45864 : 4'b1000;
															assign node45864 = (inp[14]) ? 4'b1001 : 4'b1000;
														assign node45867 = (inp[5]) ? node45875 : node45868;
															assign node45868 = (inp[14]) ? node45872 : node45869;
																assign node45869 = (inp[7]) ? 4'b1001 : 4'b1000;
																assign node45872 = (inp[7]) ? 4'b1000 : 4'b1001;
															assign node45875 = (inp[14]) ? node45879 : node45876;
																assign node45876 = (inp[7]) ? 4'b1001 : 4'b1000;
																assign node45879 = (inp[7]) ? 4'b1000 : 4'b1001;
													assign node45882 = (inp[5]) ? node45894 : node45883;
														assign node45883 = (inp[14]) ? node45889 : node45884;
															assign node45884 = (inp[7]) ? node45886 : 4'b1001;
																assign node45886 = (inp[8]) ? 4'b1001 : 4'b1000;
															assign node45889 = (inp[8]) ? 4'b1000 : node45890;
																assign node45890 = (inp[7]) ? 4'b1001 : 4'b1000;
														assign node45894 = (inp[8]) ? node45896 : 4'b1001;
															assign node45896 = (inp[14]) ? 4'b1001 : 4'b1000;
												assign node45899 = (inp[5]) ? node45911 : node45900;
													assign node45900 = (inp[14]) ? node45906 : node45901;
														assign node45901 = (inp[12]) ? node45903 : 4'b1000;
															assign node45903 = (inp[8]) ? 4'b1001 : 4'b1000;
														assign node45906 = (inp[12]) ? node45908 : 4'b1001;
															assign node45908 = (inp[8]) ? 4'b1000 : 4'b1001;
													assign node45911 = (inp[7]) ? node45927 : node45912;
														assign node45912 = (inp[12]) ? node45920 : node45913;
															assign node45913 = (inp[8]) ? node45917 : node45914;
																assign node45914 = (inp[14]) ? 4'b1010 : 4'b1011;
																assign node45917 = (inp[14]) ? 4'b1011 : 4'b1010;
															assign node45920 = (inp[14]) ? node45924 : node45921;
																assign node45921 = (inp[8]) ? 4'b1010 : 4'b1011;
																assign node45924 = (inp[8]) ? 4'b1011 : 4'b1010;
														assign node45927 = (inp[12]) ? node45929 : 4'b1011;
															assign node45929 = (inp[14]) ? node45933 : node45930;
																assign node45930 = (inp[8]) ? 4'b1011 : 4'b1010;
																assign node45933 = (inp[8]) ? 4'b1010 : 4'b1011;
											assign node45936 = (inp[3]) ? node45962 : node45937;
												assign node45937 = (inp[14]) ? node45945 : node45938;
													assign node45938 = (inp[12]) ? node45940 : 4'b1011;
														assign node45940 = (inp[8]) ? node45942 : 4'b1010;
															assign node45942 = (inp[7]) ? 4'b1011 : 4'b1010;
													assign node45945 = (inp[12]) ? node45953 : node45946;
														assign node45946 = (inp[8]) ? node45950 : node45947;
															assign node45947 = (inp[7]) ? 4'b1011 : 4'b1010;
															assign node45950 = (inp[7]) ? 4'b1010 : 4'b1011;
														assign node45953 = (inp[5]) ? node45955 : 4'b1011;
															assign node45955 = (inp[8]) ? node45959 : node45956;
																assign node45956 = (inp[7]) ? 4'b1011 : 4'b1010;
																assign node45959 = (inp[7]) ? 4'b1010 : 4'b1011;
												assign node45962 = (inp[5]) ? node45976 : node45963;
													assign node45963 = (inp[12]) ? 4'b1011 : node45964;
														assign node45964 = (inp[14]) ? node45970 : node45965;
															assign node45965 = (inp[8]) ? node45967 : 4'b1010;
																assign node45967 = (inp[7]) ? 4'b1011 : 4'b1010;
															assign node45970 = (inp[7]) ? node45972 : 4'b1011;
																assign node45972 = (inp[8]) ? 4'b1010 : 4'b1011;
													assign node45976 = (inp[12]) ? node45978 : 4'b1001;
														assign node45978 = (inp[8]) ? 4'b1001 : node45979;
															assign node45979 = (inp[14]) ? 4'b1001 : 4'b1000;
									assign node45983 = (inp[7]) ? node46061 : node45984;
										assign node45984 = (inp[8]) ? node46022 : node45985;
											assign node45985 = (inp[12]) ? node46003 : node45986;
												assign node45986 = (inp[15]) ? node45996 : node45987;
													assign node45987 = (inp[5]) ? node45991 : node45988;
														assign node45988 = (inp[0]) ? 4'b1000 : 4'b1010;
														assign node45991 = (inp[3]) ? node45993 : 4'b1000;
															assign node45993 = (inp[0]) ? 4'b1010 : 4'b1000;
													assign node45996 = (inp[3]) ? node45998 : 4'b1000;
														assign node45998 = (inp[0]) ? 4'b1000 : node45999;
															assign node45999 = (inp[5]) ? 4'b1010 : 4'b1000;
												assign node46003 = (inp[0]) ? node46011 : node46004;
													assign node46004 = (inp[15]) ? 4'b1000 : node46005;
														assign node46005 = (inp[5]) ? node46007 : 4'b1010;
															assign node46007 = (inp[3]) ? 4'b1000 : 4'b1010;
													assign node46011 = (inp[15]) ? node46017 : node46012;
														assign node46012 = (inp[5]) ? node46014 : 4'b1000;
															assign node46014 = (inp[3]) ? 4'b1010 : 4'b1000;
														assign node46017 = (inp[5]) ? node46019 : 4'b1010;
															assign node46019 = (inp[3]) ? 4'b1000 : 4'b1010;
											assign node46022 = (inp[14]) ? node46044 : node46023;
												assign node46023 = (inp[3]) ? node46031 : node46024;
													assign node46024 = (inp[15]) ? node46028 : node46025;
														assign node46025 = (inp[0]) ? 4'b1001 : 4'b1011;
														assign node46028 = (inp[0]) ? 4'b1011 : 4'b1001;
													assign node46031 = (inp[0]) ? node46039 : node46032;
														assign node46032 = (inp[15]) ? node46036 : node46033;
															assign node46033 = (inp[5]) ? 4'b1001 : 4'b1011;
															assign node46036 = (inp[5]) ? 4'b1011 : 4'b1001;
														assign node46039 = (inp[12]) ? node46041 : 4'b1011;
															assign node46041 = (inp[5]) ? 4'b1001 : 4'b1011;
												assign node46044 = (inp[15]) ? node46056 : node46045;
													assign node46045 = (inp[12]) ? node46047 : 4'b1001;
														assign node46047 = (inp[5]) ? node46049 : 4'b1001;
															assign node46049 = (inp[3]) ? node46053 : node46050;
																assign node46050 = (inp[0]) ? 4'b1001 : 4'b1011;
																assign node46053 = (inp[0]) ? 4'b1011 : 4'b1001;
													assign node46056 = (inp[0]) ? 4'b1011 : node46057;
														assign node46057 = (inp[3]) ? 4'b1011 : 4'b1001;
										assign node46061 = (inp[8]) ? node46103 : node46062;
											assign node46062 = (inp[5]) ? node46078 : node46063;
												assign node46063 = (inp[14]) ? node46071 : node46064;
													assign node46064 = (inp[0]) ? node46068 : node46065;
														assign node46065 = (inp[15]) ? 4'b1001 : 4'b1011;
														assign node46068 = (inp[15]) ? 4'b1011 : 4'b1001;
													assign node46071 = (inp[0]) ? node46075 : node46072;
														assign node46072 = (inp[15]) ? 4'b1001 : 4'b1011;
														assign node46075 = (inp[15]) ? 4'b1011 : 4'b1001;
												assign node46078 = (inp[0]) ? node46092 : node46079;
													assign node46079 = (inp[14]) ? node46085 : node46080;
														assign node46080 = (inp[3]) ? node46082 : 4'b1011;
															assign node46082 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node46085 = (inp[15]) ? node46089 : node46086;
															assign node46086 = (inp[3]) ? 4'b1001 : 4'b1011;
															assign node46089 = (inp[3]) ? 4'b1011 : 4'b1001;
													assign node46092 = (inp[14]) ? node46098 : node46093;
														assign node46093 = (inp[15]) ? 4'b1011 : node46094;
															assign node46094 = (inp[3]) ? 4'b1011 : 4'b1001;
														assign node46098 = (inp[15]) ? node46100 : 4'b1011;
															assign node46100 = (inp[3]) ? 4'b1001 : 4'b1011;
											assign node46103 = (inp[12]) ? node46139 : node46104;
												assign node46104 = (inp[3]) ? node46126 : node46105;
													assign node46105 = (inp[5]) ? node46119 : node46106;
														assign node46106 = (inp[14]) ? node46112 : node46107;
															assign node46107 = (inp[0]) ? node46109 : 4'b1010;
																assign node46109 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node46112 = (inp[15]) ? node46116 : node46113;
																assign node46113 = (inp[0]) ? 4'b1000 : 4'b1010;
																assign node46116 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node46119 = (inp[14]) ? 4'b1010 : node46120;
															assign node46120 = (inp[15]) ? node46122 : 4'b1010;
																assign node46122 = (inp[0]) ? 4'b1010 : 4'b1000;
													assign node46126 = (inp[15]) ? node46132 : node46127;
														assign node46127 = (inp[0]) ? node46129 : 4'b1000;
															assign node46129 = (inp[5]) ? 4'b1010 : 4'b1000;
														assign node46132 = (inp[0]) ? node46136 : node46133;
															assign node46133 = (inp[5]) ? 4'b1010 : 4'b1000;
															assign node46136 = (inp[5]) ? 4'b1000 : 4'b1010;
												assign node46139 = (inp[14]) ? node46157 : node46140;
													assign node46140 = (inp[5]) ? node46148 : node46141;
														assign node46141 = (inp[0]) ? node46145 : node46142;
															assign node46142 = (inp[15]) ? 4'b1000 : 4'b1010;
															assign node46145 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node46148 = (inp[0]) ? 4'b1010 : node46149;
															assign node46149 = (inp[3]) ? node46153 : node46150;
																assign node46150 = (inp[15]) ? 4'b1000 : 4'b1010;
																assign node46153 = (inp[15]) ? 4'b1010 : 4'b1000;
													assign node46157 = (inp[15]) ? node46161 : node46158;
														assign node46158 = (inp[0]) ? 4'b1000 : 4'b1010;
														assign node46161 = (inp[0]) ? node46167 : node46162;
															assign node46162 = (inp[5]) ? node46164 : 4'b1000;
																assign node46164 = (inp[3]) ? 4'b1010 : 4'b1000;
															assign node46167 = (inp[3]) ? 4'b1000 : 4'b1010;
								assign node46170 = (inp[5]) ? node46446 : node46171;
									assign node46171 = (inp[2]) ? node46331 : node46172;
										assign node46172 = (inp[0]) ? node46250 : node46173;
											assign node46173 = (inp[14]) ? node46205 : node46174;
												assign node46174 = (inp[15]) ? node46190 : node46175;
													assign node46175 = (inp[3]) ? node46183 : node46176;
														assign node46176 = (inp[8]) ? node46180 : node46177;
															assign node46177 = (inp[12]) ? 4'b1111 : 4'b1110;
															assign node46180 = (inp[7]) ? 4'b1111 : 4'b1110;
														assign node46183 = (inp[8]) ? node46187 : node46184;
															assign node46184 = (inp[7]) ? 4'b1100 : 4'b1101;
															assign node46187 = (inp[7]) ? 4'b1101 : 4'b1100;
													assign node46190 = (inp[3]) ? node46198 : node46191;
														assign node46191 = (inp[8]) ? node46195 : node46192;
															assign node46192 = (inp[7]) ? 4'b1100 : 4'b1101;
															assign node46195 = (inp[7]) ? 4'b1101 : 4'b1100;
														assign node46198 = (inp[8]) ? node46202 : node46199;
															assign node46199 = (inp[7]) ? 4'b1110 : 4'b1111;
															assign node46202 = (inp[7]) ? 4'b1111 : 4'b1110;
												assign node46205 = (inp[12]) ? node46225 : node46206;
													assign node46206 = (inp[15]) ? node46218 : node46207;
														assign node46207 = (inp[3]) ? node46215 : node46208;
															assign node46208 = (inp[7]) ? node46212 : node46209;
																assign node46209 = (inp[8]) ? 4'b1111 : 4'b1110;
																assign node46212 = (inp[8]) ? 4'b1110 : 4'b1111;
															assign node46215 = (inp[7]) ? 4'b1101 : 4'b1100;
														assign node46218 = (inp[3]) ? 4'b1111 : node46219;
															assign node46219 = (inp[7]) ? node46221 : 4'b1101;
																assign node46221 = (inp[8]) ? 4'b1100 : 4'b1101;
													assign node46225 = (inp[8]) ? node46237 : node46226;
														assign node46226 = (inp[7]) ? node46232 : node46227;
															assign node46227 = (inp[3]) ? node46229 : 4'b1110;
																assign node46229 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node46232 = (inp[15]) ? 4'b1111 : node46233;
																assign node46233 = (inp[3]) ? 4'b1101 : 4'b1111;
														assign node46237 = (inp[7]) ? node46245 : node46238;
															assign node46238 = (inp[15]) ? node46242 : node46239;
																assign node46239 = (inp[3]) ? 4'b1101 : 4'b1111;
																assign node46242 = (inp[3]) ? 4'b1111 : 4'b1101;
															assign node46245 = (inp[3]) ? node46247 : 4'b1100;
																assign node46247 = (inp[15]) ? 4'b1110 : 4'b1100;
											assign node46250 = (inp[14]) ? node46286 : node46251;
												assign node46251 = (inp[7]) ? node46267 : node46252;
													assign node46252 = (inp[8]) ? node46260 : node46253;
														assign node46253 = (inp[3]) ? node46257 : node46254;
															assign node46254 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node46257 = (inp[15]) ? 4'b1101 : 4'b1111;
														assign node46260 = (inp[3]) ? node46264 : node46261;
															assign node46261 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node46264 = (inp[15]) ? 4'b1100 : 4'b1110;
													assign node46267 = (inp[8]) ? node46275 : node46268;
														assign node46268 = (inp[3]) ? node46272 : node46269;
															assign node46269 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node46272 = (inp[15]) ? 4'b1100 : 4'b1110;
														assign node46275 = (inp[12]) ? node46281 : node46276;
															assign node46276 = (inp[3]) ? 4'b1101 : node46277;
																assign node46277 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node46281 = (inp[3]) ? node46283 : 4'b1101;
																assign node46283 = (inp[15]) ? 4'b1101 : 4'b1111;
												assign node46286 = (inp[12]) ? node46304 : node46287;
													assign node46287 = (inp[15]) ? node46299 : node46288;
														assign node46288 = (inp[3]) ? node46294 : node46289;
															assign node46289 = (inp[7]) ? 4'b1100 : node46290;
																assign node46290 = (inp[8]) ? 4'b1101 : 4'b1100;
															assign node46294 = (inp[8]) ? node46296 : 4'b1110;
																assign node46296 = (inp[7]) ? 4'b1110 : 4'b1111;
														assign node46299 = (inp[8]) ? 4'b1100 : node46300;
															assign node46300 = (inp[7]) ? 4'b1101 : 4'b1100;
													assign node46304 = (inp[15]) ? node46316 : node46305;
														assign node46305 = (inp[3]) ? node46311 : node46306;
															assign node46306 = (inp[7]) ? 4'b1100 : node46307;
																assign node46307 = (inp[8]) ? 4'b1101 : 4'b1100;
															assign node46311 = (inp[8]) ? 4'b1110 : node46312;
																assign node46312 = (inp[7]) ? 4'b1111 : 4'b1110;
														assign node46316 = (inp[3]) ? node46324 : node46317;
															assign node46317 = (inp[8]) ? node46321 : node46318;
																assign node46318 = (inp[7]) ? 4'b1111 : 4'b1110;
																assign node46321 = (inp[7]) ? 4'b1110 : 4'b1111;
															assign node46324 = (inp[7]) ? node46328 : node46325;
																assign node46325 = (inp[8]) ? 4'b1101 : 4'b1100;
																assign node46328 = (inp[8]) ? 4'b1100 : 4'b1101;
										assign node46331 = (inp[7]) ? node46387 : node46332;
											assign node46332 = (inp[8]) ? node46356 : node46333;
												assign node46333 = (inp[12]) ? node46347 : node46334;
													assign node46334 = (inp[15]) ? node46340 : node46335;
														assign node46335 = (inp[0]) ? 4'b1110 : node46336;
															assign node46336 = (inp[3]) ? 4'b1100 : 4'b1110;
														assign node46340 = (inp[3]) ? node46344 : node46341;
															assign node46341 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node46344 = (inp[0]) ? 4'b1100 : 4'b1110;
													assign node46347 = (inp[0]) ? 4'b1100 : node46348;
														assign node46348 = (inp[3]) ? node46352 : node46349;
															assign node46349 = (inp[15]) ? 4'b1100 : 4'b1110;
															assign node46352 = (inp[15]) ? 4'b1110 : 4'b1100;
												assign node46356 = (inp[14]) ? node46374 : node46357;
													assign node46357 = (inp[15]) ? node46367 : node46358;
														assign node46358 = (inp[12]) ? 4'b1101 : node46359;
															assign node46359 = (inp[0]) ? node46363 : node46360;
																assign node46360 = (inp[3]) ? 4'b1101 : 4'b1111;
																assign node46363 = (inp[3]) ? 4'b1111 : 4'b1101;
														assign node46367 = (inp[12]) ? 4'b1111 : node46368;
															assign node46368 = (inp[3]) ? 4'b1101 : node46369;
																assign node46369 = (inp[0]) ? 4'b1111 : 4'b1101;
													assign node46374 = (inp[3]) ? node46380 : node46375;
														assign node46375 = (inp[15]) ? 4'b1101 : node46376;
															assign node46376 = (inp[0]) ? 4'b1101 : 4'b1111;
														assign node46380 = (inp[0]) ? node46384 : node46381;
															assign node46381 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node46384 = (inp[15]) ? 4'b1101 : 4'b1111;
											assign node46387 = (inp[8]) ? node46425 : node46388;
												assign node46388 = (inp[14]) ? node46404 : node46389;
													assign node46389 = (inp[12]) ? node46397 : node46390;
														assign node46390 = (inp[0]) ? 4'b1101 : node46391;
															assign node46391 = (inp[15]) ? node46393 : 4'b1111;
																assign node46393 = (inp[3]) ? 4'b1111 : 4'b1101;
														assign node46397 = (inp[0]) ? 4'b1111 : node46398;
															assign node46398 = (inp[3]) ? 4'b1101 : node46399;
																assign node46399 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node46404 = (inp[12]) ? node46412 : node46405;
														assign node46405 = (inp[15]) ? node46407 : 4'b1111;
															assign node46407 = (inp[3]) ? node46409 : 4'b1111;
																assign node46409 = (inp[0]) ? 4'b1101 : 4'b1111;
														assign node46412 = (inp[3]) ? node46418 : node46413;
															assign node46413 = (inp[0]) ? node46415 : 4'b1111;
																assign node46415 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node46418 = (inp[0]) ? node46422 : node46419;
																assign node46419 = (inp[15]) ? 4'b1111 : 4'b1101;
																assign node46422 = (inp[15]) ? 4'b1101 : 4'b1111;
												assign node46425 = (inp[0]) ? node46433 : node46426;
													assign node46426 = (inp[3]) ? node46430 : node46427;
														assign node46427 = (inp[15]) ? 4'b1100 : 4'b1110;
														assign node46430 = (inp[15]) ? 4'b1110 : 4'b1100;
													assign node46433 = (inp[14]) ? node46439 : node46434;
														assign node46434 = (inp[3]) ? 4'b1110 : node46435;
															assign node46435 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node46439 = (inp[3]) ? node46443 : node46440;
															assign node46440 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node46443 = (inp[15]) ? 4'b1100 : 4'b1110;
									assign node46446 = (inp[15]) ? node46518 : node46447;
										assign node46447 = (inp[0]) ? node46471 : node46448;
											assign node46448 = (inp[8]) ? node46460 : node46449;
												assign node46449 = (inp[7]) ? node46455 : node46450;
													assign node46450 = (inp[14]) ? 4'b1100 : node46451;
														assign node46451 = (inp[2]) ? 4'b1100 : 4'b1101;
													assign node46455 = (inp[14]) ? 4'b1101 : node46456;
														assign node46456 = (inp[2]) ? 4'b1101 : 4'b1100;
												assign node46460 = (inp[7]) ? node46466 : node46461;
													assign node46461 = (inp[14]) ? 4'b1101 : node46462;
														assign node46462 = (inp[2]) ? 4'b1101 : 4'b1100;
													assign node46466 = (inp[2]) ? 4'b1100 : node46467;
														assign node46467 = (inp[12]) ? 4'b1100 : 4'b1101;
											assign node46471 = (inp[12]) ? node46491 : node46472;
												assign node46472 = (inp[7]) ? node46482 : node46473;
													assign node46473 = (inp[8]) ? node46477 : node46474;
														assign node46474 = (inp[14]) ? 4'b1110 : 4'b1111;
														assign node46477 = (inp[14]) ? 4'b1111 : node46478;
															assign node46478 = (inp[2]) ? 4'b1111 : 4'b1110;
													assign node46482 = (inp[8]) ? node46486 : node46483;
														assign node46483 = (inp[2]) ? 4'b1111 : 4'b1110;
														assign node46486 = (inp[2]) ? 4'b1110 : node46487;
															assign node46487 = (inp[14]) ? 4'b1110 : 4'b1111;
												assign node46491 = (inp[8]) ? node46503 : node46492;
													assign node46492 = (inp[7]) ? node46498 : node46493;
														assign node46493 = (inp[2]) ? 4'b1110 : node46494;
															assign node46494 = (inp[14]) ? 4'b1110 : 4'b1111;
														assign node46498 = (inp[2]) ? 4'b1111 : node46499;
															assign node46499 = (inp[3]) ? 4'b1110 : 4'b1111;
													assign node46503 = (inp[2]) ? 4'b1110 : node46504;
														assign node46504 = (inp[3]) ? node46510 : node46505;
															assign node46505 = (inp[7]) ? 4'b1110 : node46506;
																assign node46506 = (inp[14]) ? 4'b1111 : 4'b1110;
															assign node46510 = (inp[14]) ? node46514 : node46511;
																assign node46511 = (inp[7]) ? 4'b1111 : 4'b1110;
																assign node46514 = (inp[7]) ? 4'b1110 : 4'b1111;
										assign node46518 = (inp[0]) ? node46576 : node46519;
											assign node46519 = (inp[3]) ? node46539 : node46520;
												assign node46520 = (inp[14]) ? node46532 : node46521;
													assign node46521 = (inp[2]) ? node46527 : node46522;
														assign node46522 = (inp[7]) ? 4'b1110 : node46523;
															assign node46523 = (inp[8]) ? 4'b1110 : 4'b1111;
														assign node46527 = (inp[8]) ? 4'b1111 : node46528;
															assign node46528 = (inp[7]) ? 4'b1111 : 4'b1110;
													assign node46532 = (inp[7]) ? node46536 : node46533;
														assign node46533 = (inp[8]) ? 4'b1111 : 4'b1110;
														assign node46536 = (inp[8]) ? 4'b1110 : 4'b1111;
												assign node46539 = (inp[14]) ? node46569 : node46540;
													assign node46540 = (inp[12]) ? node46554 : node46541;
														assign node46541 = (inp[8]) ? node46549 : node46542;
															assign node46542 = (inp[2]) ? node46546 : node46543;
																assign node46543 = (inp[7]) ? 4'b1110 : 4'b1111;
																assign node46546 = (inp[7]) ? 4'b1111 : 4'b1110;
															assign node46549 = (inp[2]) ? 4'b1110 : node46550;
																assign node46550 = (inp[7]) ? 4'b1111 : 4'b1110;
														assign node46554 = (inp[2]) ? node46562 : node46555;
															assign node46555 = (inp[7]) ? node46559 : node46556;
																assign node46556 = (inp[8]) ? 4'b1110 : 4'b1111;
																assign node46559 = (inp[8]) ? 4'b1111 : 4'b1110;
															assign node46562 = (inp[7]) ? node46566 : node46563;
																assign node46563 = (inp[8]) ? 4'b1111 : 4'b1110;
																assign node46566 = (inp[8]) ? 4'b1110 : 4'b1111;
													assign node46569 = (inp[7]) ? node46573 : node46570;
														assign node46570 = (inp[8]) ? 4'b1111 : 4'b1110;
														assign node46573 = (inp[8]) ? 4'b1110 : 4'b1111;
											assign node46576 = (inp[12]) ? node46596 : node46577;
												assign node46577 = (inp[7]) ? node46589 : node46578;
													assign node46578 = (inp[8]) ? node46584 : node46579;
														assign node46579 = (inp[2]) ? 4'b1100 : node46580;
															assign node46580 = (inp[14]) ? 4'b1100 : 4'b1101;
														assign node46584 = (inp[14]) ? 4'b1101 : node46585;
															assign node46585 = (inp[3]) ? 4'b1100 : 4'b1101;
													assign node46589 = (inp[8]) ? 4'b1100 : node46590;
														assign node46590 = (inp[3]) ? 4'b1101 : node46591;
															assign node46591 = (inp[14]) ? 4'b1101 : 4'b1100;
												assign node46596 = (inp[8]) ? node46606 : node46597;
													assign node46597 = (inp[3]) ? node46599 : 4'b1100;
														assign node46599 = (inp[7]) ? node46603 : node46600;
															assign node46600 = (inp[14]) ? 4'b1100 : 4'b1101;
															assign node46603 = (inp[14]) ? 4'b1101 : 4'b1100;
													assign node46606 = (inp[7]) ? node46608 : 4'b1101;
														assign node46608 = (inp[2]) ? 4'b1100 : node46609;
															assign node46609 = (inp[14]) ? 4'b1100 : 4'b1101;
							assign node46613 = (inp[9]) ? node47071 : node46614;
								assign node46614 = (inp[12]) ? node46836 : node46615;
									assign node46615 = (inp[14]) ? node46739 : node46616;
										assign node46616 = (inp[3]) ? node46676 : node46617;
											assign node46617 = (inp[2]) ? node46643 : node46618;
												assign node46618 = (inp[0]) ? node46624 : node46619;
													assign node46619 = (inp[8]) ? 4'b1100 : node46620;
														assign node46620 = (inp[7]) ? 4'b1100 : 4'b1101;
													assign node46624 = (inp[15]) ? node46636 : node46625;
														assign node46625 = (inp[5]) ? node46631 : node46626;
															assign node46626 = (inp[8]) ? 4'b1101 : node46627;
																assign node46627 = (inp[7]) ? 4'b1100 : 4'b1101;
															assign node46631 = (inp[8]) ? node46633 : 4'b1111;
																assign node46633 = (inp[7]) ? 4'b1111 : 4'b1110;
														assign node46636 = (inp[5]) ? 4'b1100 : node46637;
															assign node46637 = (inp[7]) ? 4'b1110 : node46638;
																assign node46638 = (inp[8]) ? 4'b1110 : 4'b1111;
												assign node46643 = (inp[5]) ? node46665 : node46644;
													assign node46644 = (inp[0]) ? node46652 : node46645;
														assign node46645 = (inp[15]) ? 4'b1101 : node46646;
															assign node46646 = (inp[8]) ? 4'b1111 : node46647;
																assign node46647 = (inp[7]) ? 4'b1111 : 4'b1110;
														assign node46652 = (inp[15]) ? node46660 : node46653;
															assign node46653 = (inp[8]) ? node46657 : node46654;
																assign node46654 = (inp[7]) ? 4'b1101 : 4'b1100;
																assign node46657 = (inp[7]) ? 4'b1100 : 4'b1101;
															assign node46660 = (inp[8]) ? 4'b1110 : node46661;
																assign node46661 = (inp[7]) ? 4'b1111 : 4'b1110;
													assign node46665 = (inp[8]) ? node46669 : node46666;
														assign node46666 = (inp[7]) ? 4'b1101 : 4'b1100;
														assign node46669 = (inp[7]) ? 4'b1110 : node46670;
															assign node46670 = (inp[15]) ? 4'b1101 : node46671;
																assign node46671 = (inp[0]) ? 4'b1111 : 4'b1101;
											assign node46676 = (inp[8]) ? node46706 : node46677;
												assign node46677 = (inp[15]) ? node46693 : node46678;
													assign node46678 = (inp[0]) ? node46686 : node46679;
														assign node46679 = (inp[2]) ? node46683 : node46680;
															assign node46680 = (inp[7]) ? 4'b1100 : 4'b1101;
															assign node46683 = (inp[7]) ? 4'b1101 : 4'b1100;
														assign node46686 = (inp[2]) ? node46690 : node46687;
															assign node46687 = (inp[7]) ? 4'b1110 : 4'b1111;
															assign node46690 = (inp[7]) ? 4'b1111 : 4'b1110;
													assign node46693 = (inp[0]) ? node46701 : node46694;
														assign node46694 = (inp[7]) ? node46698 : node46695;
															assign node46695 = (inp[2]) ? 4'b1110 : 4'b1111;
															assign node46698 = (inp[2]) ? 4'b1111 : 4'b1110;
														assign node46701 = (inp[2]) ? node46703 : 4'b1100;
															assign node46703 = (inp[7]) ? 4'b1101 : 4'b1100;
												assign node46706 = (inp[15]) ? node46716 : node46707;
													assign node46707 = (inp[0]) ? node46709 : 4'b1100;
														assign node46709 = (inp[2]) ? node46713 : node46710;
															assign node46710 = (inp[7]) ? 4'b1111 : 4'b1110;
															assign node46713 = (inp[7]) ? 4'b1110 : 4'b1111;
													assign node46716 = (inp[0]) ? node46732 : node46717;
														assign node46717 = (inp[5]) ? node46725 : node46718;
															assign node46718 = (inp[2]) ? node46722 : node46719;
																assign node46719 = (inp[7]) ? 4'b1111 : 4'b1110;
																assign node46722 = (inp[7]) ? 4'b1110 : 4'b1111;
															assign node46725 = (inp[2]) ? node46729 : node46726;
																assign node46726 = (inp[7]) ? 4'b1111 : 4'b1110;
																assign node46729 = (inp[7]) ? 4'b1110 : 4'b1111;
														assign node46732 = (inp[2]) ? node46736 : node46733;
															assign node46733 = (inp[7]) ? 4'b1101 : 4'b1100;
															assign node46736 = (inp[7]) ? 4'b1100 : 4'b1101;
										assign node46739 = (inp[8]) ? node46791 : node46740;
											assign node46740 = (inp[7]) ? node46764 : node46741;
												assign node46741 = (inp[15]) ? node46753 : node46742;
													assign node46742 = (inp[0]) ? node46748 : node46743;
														assign node46743 = (inp[3]) ? 4'b1100 : node46744;
															assign node46744 = (inp[5]) ? 4'b1100 : 4'b1110;
														assign node46748 = (inp[3]) ? 4'b1110 : node46749;
															assign node46749 = (inp[5]) ? 4'b1110 : 4'b1100;
													assign node46753 = (inp[0]) ? node46759 : node46754;
														assign node46754 = (inp[5]) ? 4'b1110 : node46755;
															assign node46755 = (inp[3]) ? 4'b1110 : 4'b1100;
														assign node46759 = (inp[5]) ? 4'b1100 : node46760;
															assign node46760 = (inp[3]) ? 4'b1100 : 4'b1110;
												assign node46764 = (inp[5]) ? node46780 : node46765;
													assign node46765 = (inp[2]) ? node46775 : node46766;
														assign node46766 = (inp[0]) ? node46768 : 4'b1101;
															assign node46768 = (inp[3]) ? node46772 : node46769;
																assign node46769 = (inp[15]) ? 4'b1111 : 4'b1101;
																assign node46772 = (inp[15]) ? 4'b1101 : 4'b1111;
														assign node46775 = (inp[3]) ? node46777 : 4'b1111;
															assign node46777 = (inp[0]) ? 4'b1111 : 4'b1101;
													assign node46780 = (inp[2]) ? node46786 : node46781;
														assign node46781 = (inp[0]) ? node46783 : 4'b1111;
															assign node46783 = (inp[15]) ? 4'b1101 : 4'b1111;
														assign node46786 = (inp[0]) ? 4'b1101 : node46787;
															assign node46787 = (inp[15]) ? 4'b1111 : 4'b1101;
											assign node46791 = (inp[7]) ? node46811 : node46792;
												assign node46792 = (inp[0]) ? node46800 : node46793;
													assign node46793 = (inp[15]) ? node46797 : node46794;
														assign node46794 = (inp[3]) ? 4'b1101 : 4'b1111;
														assign node46797 = (inp[3]) ? 4'b1111 : 4'b1101;
													assign node46800 = (inp[15]) ? node46806 : node46801;
														assign node46801 = (inp[3]) ? 4'b1111 : node46802;
															assign node46802 = (inp[5]) ? 4'b1111 : 4'b1101;
														assign node46806 = (inp[5]) ? 4'b1101 : node46807;
															assign node46807 = (inp[3]) ? 4'b1101 : 4'b1111;
												assign node46811 = (inp[3]) ? node46829 : node46812;
													assign node46812 = (inp[5]) ? node46824 : node46813;
														assign node46813 = (inp[2]) ? node46819 : node46814;
															assign node46814 = (inp[15]) ? 4'b1110 : node46815;
																assign node46815 = (inp[0]) ? 4'b1100 : 4'b1110;
															assign node46819 = (inp[15]) ? node46821 : 4'b1100;
																assign node46821 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node46824 = (inp[0]) ? 4'b1110 : node46825;
															assign node46825 = (inp[15]) ? 4'b1110 : 4'b1100;
													assign node46829 = (inp[15]) ? node46833 : node46830;
														assign node46830 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node46833 = (inp[0]) ? 4'b1100 : 4'b1110;
									assign node46836 = (inp[15]) ? node46970 : node46837;
										assign node46837 = (inp[0]) ? node46903 : node46838;
											assign node46838 = (inp[3]) ? node46864 : node46839;
												assign node46839 = (inp[5]) ? node46851 : node46840;
													assign node46840 = (inp[7]) ? node46848 : node46841;
														assign node46841 = (inp[8]) ? node46845 : node46842;
															assign node46842 = (inp[2]) ? 4'b1110 : 4'b1111;
															assign node46845 = (inp[2]) ? 4'b1111 : 4'b1110;
														assign node46848 = (inp[8]) ? 4'b1110 : 4'b1111;
													assign node46851 = (inp[14]) ? node46857 : node46852;
														assign node46852 = (inp[8]) ? node46854 : 4'b1101;
															assign node46854 = (inp[7]) ? 4'b1101 : 4'b1100;
														assign node46857 = (inp[8]) ? node46861 : node46858;
															assign node46858 = (inp[7]) ? 4'b1101 : 4'b1100;
															assign node46861 = (inp[7]) ? 4'b1100 : 4'b1101;
												assign node46864 = (inp[14]) ? node46890 : node46865;
													assign node46865 = (inp[8]) ? node46881 : node46866;
														assign node46866 = (inp[5]) ? node46874 : node46867;
															assign node46867 = (inp[7]) ? node46871 : node46868;
																assign node46868 = (inp[2]) ? 4'b1100 : 4'b1101;
																assign node46871 = (inp[2]) ? 4'b1101 : 4'b1100;
															assign node46874 = (inp[2]) ? node46878 : node46875;
																assign node46875 = (inp[7]) ? 4'b1100 : 4'b1101;
																assign node46878 = (inp[7]) ? 4'b1101 : 4'b1100;
														assign node46881 = (inp[5]) ? node46883 : 4'b1100;
															assign node46883 = (inp[7]) ? node46887 : node46884;
																assign node46884 = (inp[2]) ? 4'b1101 : 4'b1100;
																assign node46887 = (inp[2]) ? 4'b1100 : 4'b1101;
													assign node46890 = (inp[2]) ? 4'b1101 : node46891;
														assign node46891 = (inp[5]) ? node46897 : node46892;
															assign node46892 = (inp[8]) ? node46894 : 4'b1100;
																assign node46894 = (inp[7]) ? 4'b1100 : 4'b1101;
															assign node46897 = (inp[8]) ? 4'b1101 : node46898;
																assign node46898 = (inp[7]) ? 4'b1101 : 4'b1100;
											assign node46903 = (inp[3]) ? node46947 : node46904;
												assign node46904 = (inp[5]) ? node46930 : node46905;
													assign node46905 = (inp[14]) ? node46919 : node46906;
														assign node46906 = (inp[2]) ? node46914 : node46907;
															assign node46907 = (inp[7]) ? node46911 : node46908;
																assign node46908 = (inp[8]) ? 4'b1100 : 4'b1101;
																assign node46911 = (inp[8]) ? 4'b1101 : 4'b1100;
															assign node46914 = (inp[8]) ? node46916 : 4'b1101;
																assign node46916 = (inp[7]) ? 4'b1100 : 4'b1101;
														assign node46919 = (inp[2]) ? node46925 : node46920;
															assign node46920 = (inp[8]) ? node46922 : 4'b1100;
																assign node46922 = (inp[7]) ? 4'b1100 : 4'b1101;
															assign node46925 = (inp[7]) ? node46927 : 4'b1100;
																assign node46927 = (inp[8]) ? 4'b1100 : 4'b1101;
													assign node46930 = (inp[8]) ? node46938 : node46931;
														assign node46931 = (inp[7]) ? node46933 : 4'b1110;
															assign node46933 = (inp[14]) ? 4'b1111 : node46934;
																assign node46934 = (inp[2]) ? 4'b1111 : 4'b1110;
														assign node46938 = (inp[14]) ? node46944 : node46939;
															assign node46939 = (inp[2]) ? 4'b1111 : node46940;
																assign node46940 = (inp[7]) ? 4'b1111 : 4'b1110;
															assign node46944 = (inp[7]) ? 4'b1110 : 4'b1111;
												assign node46947 = (inp[14]) ? node46963 : node46948;
													assign node46948 = (inp[2]) ? node46954 : node46949;
														assign node46949 = (inp[7]) ? 4'b1111 : node46950;
															assign node46950 = (inp[8]) ? 4'b1110 : 4'b1111;
														assign node46954 = (inp[5]) ? 4'b1110 : node46955;
															assign node46955 = (inp[7]) ? node46959 : node46956;
																assign node46956 = (inp[8]) ? 4'b1111 : 4'b1110;
																assign node46959 = (inp[8]) ? 4'b1110 : 4'b1111;
													assign node46963 = (inp[8]) ? node46967 : node46964;
														assign node46964 = (inp[7]) ? 4'b1111 : 4'b1110;
														assign node46967 = (inp[7]) ? 4'b1110 : 4'b1111;
										assign node46970 = (inp[0]) ? node47014 : node46971;
											assign node46971 = (inp[3]) ? node46997 : node46972;
												assign node46972 = (inp[5]) ? node46982 : node46973;
													assign node46973 = (inp[8]) ? node46977 : node46974;
														assign node46974 = (inp[14]) ? 4'b1100 : 4'b1101;
														assign node46977 = (inp[7]) ? node46979 : 4'b1101;
															assign node46979 = (inp[2]) ? 4'b1100 : 4'b1101;
													assign node46982 = (inp[2]) ? node46990 : node46983;
														assign node46983 = (inp[8]) ? 4'b1110 : node46984;
															assign node46984 = (inp[7]) ? node46986 : 4'b1110;
																assign node46986 = (inp[14]) ? 4'b1111 : 4'b1110;
														assign node46990 = (inp[8]) ? node46994 : node46991;
															assign node46991 = (inp[7]) ? 4'b1111 : 4'b1110;
															assign node46994 = (inp[7]) ? 4'b1110 : 4'b1111;
												assign node46997 = (inp[2]) ? node47007 : node46998;
													assign node46998 = (inp[14]) ? 4'b1111 : node46999;
														assign node46999 = (inp[8]) ? node47003 : node47000;
															assign node47000 = (inp[7]) ? 4'b1110 : 4'b1111;
															assign node47003 = (inp[7]) ? 4'b1111 : 4'b1110;
													assign node47007 = (inp[7]) ? node47011 : node47008;
														assign node47008 = (inp[8]) ? 4'b1111 : 4'b1110;
														assign node47011 = (inp[8]) ? 4'b1110 : 4'b1111;
											assign node47014 = (inp[3]) ? node47046 : node47015;
												assign node47015 = (inp[5]) ? node47037 : node47016;
													assign node47016 = (inp[7]) ? node47026 : node47017;
														assign node47017 = (inp[14]) ? node47023 : node47018;
															assign node47018 = (inp[8]) ? node47020 : 4'b1111;
																assign node47020 = (inp[2]) ? 4'b1111 : 4'b1110;
															assign node47023 = (inp[8]) ? 4'b1111 : 4'b1110;
														assign node47026 = (inp[8]) ? node47032 : node47027;
															assign node47027 = (inp[2]) ? 4'b1111 : node47028;
																assign node47028 = (inp[14]) ? 4'b1111 : 4'b1110;
															assign node47032 = (inp[2]) ? 4'b1110 : node47033;
																assign node47033 = (inp[14]) ? 4'b1110 : 4'b1111;
													assign node47037 = (inp[8]) ? 4'b1100 : node47038;
														assign node47038 = (inp[7]) ? node47042 : node47039;
															assign node47039 = (inp[2]) ? 4'b1100 : 4'b1101;
															assign node47042 = (inp[14]) ? 4'b1101 : 4'b1100;
												assign node47046 = (inp[5]) ? node47060 : node47047;
													assign node47047 = (inp[8]) ? node47053 : node47048;
														assign node47048 = (inp[7]) ? 4'b1101 : node47049;
															assign node47049 = (inp[14]) ? 4'b1100 : 4'b1101;
														assign node47053 = (inp[7]) ? 4'b1100 : node47054;
															assign node47054 = (inp[2]) ? 4'b1101 : node47055;
																assign node47055 = (inp[14]) ? 4'b1101 : 4'b1100;
													assign node47060 = (inp[14]) ? 4'b1100 : node47061;
														assign node47061 = (inp[2]) ? 4'b1100 : node47062;
															assign node47062 = (inp[7]) ? node47066 : node47063;
																assign node47063 = (inp[8]) ? 4'b1100 : 4'b1101;
																assign node47066 = (inp[8]) ? 4'b1101 : 4'b1100;
								assign node47071 = (inp[14]) ? node47261 : node47072;
									assign node47072 = (inp[8]) ? node47172 : node47073;
										assign node47073 = (inp[2]) ? node47121 : node47074;
											assign node47074 = (inp[7]) ? node47100 : node47075;
												assign node47075 = (inp[12]) ? node47089 : node47076;
													assign node47076 = (inp[15]) ? node47084 : node47077;
														assign node47077 = (inp[0]) ? node47081 : node47078;
															assign node47078 = (inp[3]) ? 4'b1001 : 4'b1011;
															assign node47081 = (inp[3]) ? 4'b1011 : 4'b1001;
														assign node47084 = (inp[3]) ? 4'b1011 : node47085;
															assign node47085 = (inp[5]) ? 4'b1001 : 4'b1011;
													assign node47089 = (inp[0]) ? node47093 : node47090;
														assign node47090 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node47093 = (inp[15]) ? 4'b1001 : node47094;
															assign node47094 = (inp[5]) ? 4'b1011 : node47095;
																assign node47095 = (inp[3]) ? 4'b1011 : 4'b1001;
												assign node47100 = (inp[3]) ? node47114 : node47101;
													assign node47101 = (inp[12]) ? node47107 : node47102;
														assign node47102 = (inp[5]) ? 4'b1000 : node47103;
															assign node47103 = (inp[15]) ? 4'b1000 : 4'b1010;
														assign node47107 = (inp[15]) ? node47111 : node47108;
															assign node47108 = (inp[0]) ? 4'b1010 : 4'b1000;
															assign node47111 = (inp[0]) ? 4'b1000 : 4'b1010;
													assign node47114 = (inp[15]) ? node47118 : node47115;
														assign node47115 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node47118 = (inp[0]) ? 4'b1000 : 4'b1010;
											assign node47121 = (inp[7]) ? node47145 : node47122;
												assign node47122 = (inp[15]) ? node47134 : node47123;
													assign node47123 = (inp[0]) ? node47129 : node47124;
														assign node47124 = (inp[5]) ? 4'b1000 : node47125;
															assign node47125 = (inp[3]) ? 4'b1000 : 4'b1010;
														assign node47129 = (inp[5]) ? 4'b1010 : node47130;
															assign node47130 = (inp[3]) ? 4'b1010 : 4'b1000;
													assign node47134 = (inp[0]) ? node47140 : node47135;
														assign node47135 = (inp[5]) ? 4'b1010 : node47136;
															assign node47136 = (inp[3]) ? 4'b1010 : 4'b1000;
														assign node47140 = (inp[3]) ? 4'b1000 : node47141;
															assign node47141 = (inp[5]) ? 4'b1000 : 4'b1010;
												assign node47145 = (inp[3]) ? node47163 : node47146;
													assign node47146 = (inp[0]) ? node47156 : node47147;
														assign node47147 = (inp[12]) ? node47153 : node47148;
															assign node47148 = (inp[5]) ? 4'b1011 : node47149;
																assign node47149 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node47153 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node47156 = (inp[5]) ? node47160 : node47157;
															assign node47157 = (inp[15]) ? 4'b1011 : 4'b1001;
															assign node47160 = (inp[15]) ? 4'b1001 : 4'b1011;
													assign node47163 = (inp[5]) ? 4'b1001 : node47164;
														assign node47164 = (inp[12]) ? 4'b1001 : node47165;
															assign node47165 = (inp[15]) ? node47167 : 4'b1011;
																assign node47167 = (inp[0]) ? 4'b1001 : 4'b1011;
										assign node47172 = (inp[0]) ? node47222 : node47173;
											assign node47173 = (inp[15]) ? node47197 : node47174;
												assign node47174 = (inp[5]) ? node47190 : node47175;
													assign node47175 = (inp[3]) ? node47183 : node47176;
														assign node47176 = (inp[7]) ? node47180 : node47177;
															assign node47177 = (inp[2]) ? 4'b1011 : 4'b1010;
															assign node47180 = (inp[2]) ? 4'b1010 : 4'b1011;
														assign node47183 = (inp[2]) ? node47187 : node47184;
															assign node47184 = (inp[7]) ? 4'b1001 : 4'b1000;
															assign node47187 = (inp[7]) ? 4'b1000 : 4'b1001;
													assign node47190 = (inp[2]) ? node47194 : node47191;
														assign node47191 = (inp[7]) ? 4'b1001 : 4'b1000;
														assign node47194 = (inp[7]) ? 4'b1000 : 4'b1001;
												assign node47197 = (inp[3]) ? node47215 : node47198;
													assign node47198 = (inp[5]) ? node47208 : node47199;
														assign node47199 = (inp[12]) ? node47205 : node47200;
															assign node47200 = (inp[2]) ? 4'b1001 : node47201;
																assign node47201 = (inp[7]) ? 4'b1001 : 4'b1000;
															assign node47205 = (inp[7]) ? 4'b1000 : 4'b1001;
														assign node47208 = (inp[7]) ? node47212 : node47209;
															assign node47209 = (inp[2]) ? 4'b1011 : 4'b1010;
															assign node47212 = (inp[2]) ? 4'b1010 : 4'b1011;
													assign node47215 = (inp[7]) ? node47219 : node47216;
														assign node47216 = (inp[2]) ? 4'b1011 : 4'b1010;
														assign node47219 = (inp[2]) ? 4'b1010 : 4'b1011;
											assign node47222 = (inp[15]) ? node47240 : node47223;
												assign node47223 = (inp[5]) ? node47233 : node47224;
													assign node47224 = (inp[3]) ? node47228 : node47225;
														assign node47225 = (inp[2]) ? 4'b1000 : 4'b1001;
														assign node47228 = (inp[7]) ? node47230 : 4'b1011;
															assign node47230 = (inp[2]) ? 4'b1010 : 4'b1011;
													assign node47233 = (inp[7]) ? node47237 : node47234;
														assign node47234 = (inp[2]) ? 4'b1011 : 4'b1010;
														assign node47237 = (inp[2]) ? 4'b1010 : 4'b1011;
												assign node47240 = (inp[3]) ? node47254 : node47241;
													assign node47241 = (inp[5]) ? node47249 : node47242;
														assign node47242 = (inp[7]) ? node47246 : node47243;
															assign node47243 = (inp[2]) ? 4'b1011 : 4'b1010;
															assign node47246 = (inp[2]) ? 4'b1010 : 4'b1011;
														assign node47249 = (inp[2]) ? node47251 : 4'b1000;
															assign node47251 = (inp[7]) ? 4'b1000 : 4'b1001;
													assign node47254 = (inp[7]) ? node47258 : node47255;
														assign node47255 = (inp[2]) ? 4'b1001 : 4'b1000;
														assign node47258 = (inp[2]) ? 4'b1000 : 4'b1001;
									assign node47261 = (inp[8]) ? node47375 : node47262;
										assign node47262 = (inp[7]) ? node47312 : node47263;
											assign node47263 = (inp[2]) ? node47295 : node47264;
												assign node47264 = (inp[5]) ? node47278 : node47265;
													assign node47265 = (inp[15]) ? node47273 : node47266;
														assign node47266 = (inp[0]) ? node47270 : node47267;
															assign node47267 = (inp[3]) ? 4'b1000 : 4'b1010;
															assign node47270 = (inp[3]) ? 4'b1010 : 4'b1000;
														assign node47273 = (inp[0]) ? 4'b1000 : node47274;
															assign node47274 = (inp[3]) ? 4'b1010 : 4'b1000;
													assign node47278 = (inp[3]) ? 4'b1000 : node47279;
														assign node47279 = (inp[12]) ? node47287 : node47280;
															assign node47280 = (inp[15]) ? node47284 : node47281;
																assign node47281 = (inp[0]) ? 4'b1010 : 4'b1000;
																assign node47284 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node47287 = (inp[15]) ? node47291 : node47288;
																assign node47288 = (inp[0]) ? 4'b1010 : 4'b1000;
																assign node47291 = (inp[0]) ? 4'b1000 : 4'b1010;
												assign node47295 = (inp[15]) ? node47307 : node47296;
													assign node47296 = (inp[0]) ? node47302 : node47297;
														assign node47297 = (inp[5]) ? 4'b1000 : node47298;
															assign node47298 = (inp[3]) ? 4'b1000 : 4'b1010;
														assign node47302 = (inp[5]) ? 4'b1010 : node47303;
															assign node47303 = (inp[3]) ? 4'b1010 : 4'b1000;
													assign node47307 = (inp[0]) ? node47309 : 4'b1010;
														assign node47309 = (inp[3]) ? 4'b1000 : 4'b1010;
											assign node47312 = (inp[3]) ? node47338 : node47313;
												assign node47313 = (inp[0]) ? node47321 : node47314;
													assign node47314 = (inp[12]) ? 4'b1011 : node47315;
														assign node47315 = (inp[15]) ? node47317 : 4'b1011;
															assign node47317 = (inp[5]) ? 4'b1011 : 4'b1001;
													assign node47321 = (inp[12]) ? node47329 : node47322;
														assign node47322 = (inp[15]) ? node47326 : node47323;
															assign node47323 = (inp[5]) ? 4'b1011 : 4'b1001;
															assign node47326 = (inp[5]) ? 4'b1001 : 4'b1011;
														assign node47329 = (inp[2]) ? 4'b1011 : node47330;
															assign node47330 = (inp[15]) ? node47334 : node47331;
																assign node47331 = (inp[5]) ? 4'b1011 : 4'b1001;
																assign node47334 = (inp[5]) ? 4'b1001 : 4'b1011;
												assign node47338 = (inp[2]) ? node47358 : node47339;
													assign node47339 = (inp[12]) ? node47351 : node47340;
														assign node47340 = (inp[5]) ? node47346 : node47341;
															assign node47341 = (inp[15]) ? node47343 : 4'b1011;
																assign node47343 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node47346 = (inp[15]) ? 4'b1011 : node47347;
																assign node47347 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node47351 = (inp[15]) ? node47355 : node47352;
															assign node47352 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node47355 = (inp[0]) ? 4'b1001 : 4'b1011;
													assign node47358 = (inp[12]) ? node47368 : node47359;
														assign node47359 = (inp[5]) ? 4'b1001 : node47360;
															assign node47360 = (inp[0]) ? node47364 : node47361;
																assign node47361 = (inp[15]) ? 4'b1011 : 4'b1001;
																assign node47364 = (inp[15]) ? 4'b1001 : 4'b1011;
														assign node47368 = (inp[5]) ? 4'b1011 : node47369;
															assign node47369 = (inp[0]) ? 4'b1001 : node47370;
																assign node47370 = (inp[15]) ? 4'b1011 : 4'b1001;
										assign node47375 = (inp[7]) ? node47397 : node47376;
											assign node47376 = (inp[15]) ? node47388 : node47377;
												assign node47377 = (inp[0]) ? node47383 : node47378;
													assign node47378 = (inp[5]) ? 4'b1001 : node47379;
														assign node47379 = (inp[3]) ? 4'b1001 : 4'b1011;
													assign node47383 = (inp[5]) ? 4'b1011 : node47384;
														assign node47384 = (inp[3]) ? 4'b1011 : 4'b1001;
												assign node47388 = (inp[3]) ? 4'b1001 : node47389;
													assign node47389 = (inp[0]) ? node47393 : node47390;
														assign node47390 = (inp[5]) ? 4'b1011 : 4'b1001;
														assign node47393 = (inp[5]) ? 4'b1001 : 4'b1011;
											assign node47397 = (inp[15]) ? node47409 : node47398;
												assign node47398 = (inp[0]) ? node47404 : node47399;
													assign node47399 = (inp[5]) ? 4'b1000 : node47400;
														assign node47400 = (inp[3]) ? 4'b1000 : 4'b1010;
													assign node47404 = (inp[5]) ? 4'b1010 : node47405;
														assign node47405 = (inp[3]) ? 4'b1010 : 4'b1000;
												assign node47409 = (inp[0]) ? node47415 : node47410;
													assign node47410 = (inp[3]) ? 4'b1010 : node47411;
														assign node47411 = (inp[5]) ? 4'b1010 : 4'b1000;
													assign node47415 = (inp[5]) ? 4'b1000 : node47416;
														assign node47416 = (inp[3]) ? 4'b1000 : 4'b1010;
			assign node47420 = (inp[6]) ? node54784 : node47421;
				assign node47421 = (inp[13]) ? node51415 : node47422;
					assign node47422 = (inp[1]) ? node49542 : node47423;
						assign node47423 = (inp[8]) ? node48479 : node47424;
							assign node47424 = (inp[7]) ? node47934 : node47425;
								assign node47425 = (inp[2]) ? node47685 : node47426;
									assign node47426 = (inp[14]) ? node47562 : node47427;
										assign node47427 = (inp[9]) ? node47481 : node47428;
											assign node47428 = (inp[4]) ? node47456 : node47429;
												assign node47429 = (inp[12]) ? node47447 : node47430;
													assign node47430 = (inp[3]) ? node47438 : node47431;
														assign node47431 = (inp[15]) ? node47435 : node47432;
															assign node47432 = (inp[0]) ? 4'b0101 : 4'b0111;
															assign node47435 = (inp[0]) ? 4'b0111 : 4'b0101;
														assign node47438 = (inp[5]) ? 4'b0101 : node47439;
															assign node47439 = (inp[0]) ? node47443 : node47440;
																assign node47440 = (inp[15]) ? 4'b0101 : 4'b0111;
																assign node47443 = (inp[15]) ? 4'b0111 : 4'b0101;
													assign node47447 = (inp[5]) ? node47451 : node47448;
														assign node47448 = (inp[3]) ? 4'b0011 : 4'b0001;
														assign node47451 = (inp[15]) ? 4'b0001 : node47452;
															assign node47452 = (inp[3]) ? 4'b0001 : 4'b0011;
												assign node47456 = (inp[12]) ? node47470 : node47457;
													assign node47457 = (inp[5]) ? node47463 : node47458;
														assign node47458 = (inp[15]) ? node47460 : 4'b0001;
															assign node47460 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node47463 = (inp[15]) ? node47465 : 4'b0011;
															assign node47465 = (inp[3]) ? node47467 : 4'b0001;
																assign node47467 = (inp[0]) ? 4'b0001 : 4'b0011;
													assign node47470 = (inp[15]) ? node47478 : node47471;
														assign node47471 = (inp[0]) ? node47473 : 4'b0101;
															assign node47473 = (inp[3]) ? 4'b0111 : node47474;
																assign node47474 = (inp[5]) ? 4'b0111 : 4'b0101;
														assign node47478 = (inp[0]) ? 4'b0101 : 4'b0111;
											assign node47481 = (inp[15]) ? node47519 : node47482;
												assign node47482 = (inp[5]) ? node47504 : node47483;
													assign node47483 = (inp[0]) ? node47491 : node47484;
														assign node47484 = (inp[3]) ? 4'b0001 : node47485;
															assign node47485 = (inp[12]) ? 4'b0011 : node47486;
																assign node47486 = (inp[4]) ? 4'b0111 : 4'b0011;
														assign node47491 = (inp[3]) ? node47497 : node47492;
															assign node47492 = (inp[12]) ? 4'b0001 : node47493;
																assign node47493 = (inp[4]) ? 4'b0101 : 4'b0001;
															assign node47497 = (inp[4]) ? node47501 : node47498;
																assign node47498 = (inp[12]) ? 4'b0111 : 4'b0001;
																assign node47501 = (inp[12]) ? 4'b0011 : 4'b0111;
													assign node47504 = (inp[0]) ? node47514 : node47505;
														assign node47505 = (inp[4]) ? node47511 : node47506;
															assign node47506 = (inp[12]) ? 4'b0101 : node47507;
																assign node47507 = (inp[3]) ? 4'b0001 : 4'b0011;
															assign node47511 = (inp[12]) ? 4'b0001 : 4'b0101;
														assign node47514 = (inp[3]) ? 4'b0011 : node47515;
															assign node47515 = (inp[4]) ? 4'b0111 : 4'b0001;
												assign node47519 = (inp[0]) ? node47543 : node47520;
													assign node47520 = (inp[3]) ? node47532 : node47521;
														assign node47521 = (inp[5]) ? node47527 : node47522;
															assign node47522 = (inp[12]) ? 4'b0001 : node47523;
																assign node47523 = (inp[4]) ? 4'b0101 : 4'b0001;
															assign node47527 = (inp[12]) ? 4'b0111 : node47528;
																assign node47528 = (inp[4]) ? 4'b0111 : 4'b0001;
														assign node47532 = (inp[5]) ? node47538 : node47533;
															assign node47533 = (inp[4]) ? node47535 : 4'b0111;
																assign node47535 = (inp[12]) ? 4'b0011 : 4'b0111;
															assign node47538 = (inp[4]) ? 4'b0011 : node47539;
																assign node47539 = (inp[12]) ? 4'b0111 : 4'b0011;
													assign node47543 = (inp[3]) ? node47553 : node47544;
														assign node47544 = (inp[4]) ? node47548 : node47545;
															assign node47545 = (inp[12]) ? 4'b0111 : 4'b0011;
															assign node47548 = (inp[12]) ? 4'b0001 : node47549;
																assign node47549 = (inp[5]) ? 4'b0101 : 4'b0111;
														assign node47553 = (inp[4]) ? node47559 : node47554;
															assign node47554 = (inp[12]) ? 4'b0101 : node47555;
																assign node47555 = (inp[5]) ? 4'b0001 : 4'b0011;
															assign node47559 = (inp[12]) ? 4'b0001 : 4'b0101;
										assign node47562 = (inp[9]) ? node47626 : node47563;
											assign node47563 = (inp[3]) ? node47599 : node47564;
												assign node47564 = (inp[0]) ? node47580 : node47565;
													assign node47565 = (inp[15]) ? node47573 : node47566;
														assign node47566 = (inp[4]) ? node47570 : node47567;
															assign node47567 = (inp[12]) ? 4'b0010 : 4'b0110;
															assign node47570 = (inp[12]) ? 4'b0100 : 4'b0010;
														assign node47573 = (inp[4]) ? node47577 : node47574;
															assign node47574 = (inp[12]) ? 4'b0000 : 4'b0100;
															assign node47577 = (inp[12]) ? 4'b0110 : 4'b0000;
													assign node47580 = (inp[15]) ? node47594 : node47581;
														assign node47581 = (inp[5]) ? node47587 : node47582;
															assign node47582 = (inp[4]) ? node47584 : 4'b0000;
																assign node47584 = (inp[12]) ? 4'b0100 : 4'b0000;
															assign node47587 = (inp[12]) ? node47591 : node47588;
																assign node47588 = (inp[4]) ? 4'b0000 : 4'b0100;
																assign node47591 = (inp[4]) ? 4'b0110 : 4'b0000;
														assign node47594 = (inp[5]) ? 4'b0110 : node47595;
															assign node47595 = (inp[12]) ? 4'b0110 : 4'b0010;
												assign node47599 = (inp[12]) ? node47611 : node47600;
													assign node47600 = (inp[4]) ? node47604 : node47601;
														assign node47601 = (inp[5]) ? 4'b0110 : 4'b0100;
														assign node47604 = (inp[0]) ? node47606 : 4'b0010;
															assign node47606 = (inp[5]) ? node47608 : 4'b0010;
																assign node47608 = (inp[15]) ? 4'b0000 : 4'b0010;
													assign node47611 = (inp[4]) ? node47621 : node47612;
														assign node47612 = (inp[15]) ? 4'b0010 : node47613;
															assign node47613 = (inp[5]) ? node47617 : node47614;
																assign node47614 = (inp[0]) ? 4'b0000 : 4'b0010;
																assign node47617 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node47621 = (inp[5]) ? 4'b0100 : node47622;
															assign node47622 = (inp[15]) ? 4'b0110 : 4'b0100;
											assign node47626 = (inp[15]) ? node47652 : node47627;
												assign node47627 = (inp[0]) ? node47639 : node47628;
													assign node47628 = (inp[3]) ? node47632 : node47629;
														assign node47629 = (inp[5]) ? 4'b0100 : 4'b0110;
														assign node47632 = (inp[4]) ? node47636 : node47633;
															assign node47633 = (inp[12]) ? 4'b0100 : 4'b0000;
															assign node47636 = (inp[12]) ? 4'b0000 : 4'b0100;
													assign node47639 = (inp[3]) ? node47647 : node47640;
														assign node47640 = (inp[4]) ? 4'b0000 : node47641;
															assign node47641 = (inp[12]) ? node47643 : 4'b0000;
																assign node47643 = (inp[5]) ? 4'b0110 : 4'b0100;
														assign node47647 = (inp[4]) ? 4'b0110 : node47648;
															assign node47648 = (inp[12]) ? 4'b0110 : 4'b0000;
												assign node47652 = (inp[5]) ? node47670 : node47653;
													assign node47653 = (inp[12]) ? node47663 : node47654;
														assign node47654 = (inp[4]) ? node47658 : node47655;
															assign node47655 = (inp[0]) ? 4'b0010 : 4'b0000;
															assign node47658 = (inp[0]) ? 4'b0100 : node47659;
																assign node47659 = (inp[3]) ? 4'b0110 : 4'b0100;
														assign node47663 = (inp[4]) ? node47665 : 4'b0110;
															assign node47665 = (inp[3]) ? 4'b0010 : node47666;
																assign node47666 = (inp[0]) ? 4'b0010 : 4'b0000;
													assign node47670 = (inp[0]) ? node47676 : node47671;
														assign node47671 = (inp[4]) ? node47673 : 4'b0000;
															assign node47673 = (inp[12]) ? 4'b0010 : 4'b0110;
														assign node47676 = (inp[12]) ? node47682 : node47677;
															assign node47677 = (inp[4]) ? 4'b0100 : node47678;
																assign node47678 = (inp[3]) ? 4'b0000 : 4'b0010;
															assign node47682 = (inp[4]) ? 4'b0000 : 4'b0100;
									assign node47685 = (inp[15]) ? node47811 : node47686;
										assign node47686 = (inp[3]) ? node47752 : node47687;
											assign node47687 = (inp[0]) ? node47713 : node47688;
												assign node47688 = (inp[5]) ? node47704 : node47689;
													assign node47689 = (inp[14]) ? node47695 : node47690;
														assign node47690 = (inp[9]) ? 4'b0110 : node47691;
															assign node47691 = (inp[4]) ? 4'b0110 : 4'b0010;
														assign node47695 = (inp[9]) ? 4'b0010 : node47696;
															assign node47696 = (inp[4]) ? node47700 : node47697;
																assign node47697 = (inp[12]) ? 4'b0010 : 4'b0110;
																assign node47700 = (inp[12]) ? 4'b0110 : 4'b0010;
													assign node47704 = (inp[9]) ? node47706 : 4'b0100;
														assign node47706 = (inp[12]) ? node47710 : node47707;
															assign node47707 = (inp[4]) ? 4'b0100 : 4'b0010;
															assign node47710 = (inp[4]) ? 4'b0000 : 4'b0100;
												assign node47713 = (inp[5]) ? node47741 : node47714;
													assign node47714 = (inp[14]) ? node47728 : node47715;
														assign node47715 = (inp[9]) ? node47721 : node47716;
															assign node47716 = (inp[4]) ? node47718 : 4'b0100;
																assign node47718 = (inp[12]) ? 4'b0100 : 4'b0000;
															assign node47721 = (inp[12]) ? node47725 : node47722;
																assign node47722 = (inp[4]) ? 4'b0100 : 4'b0000;
																assign node47725 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node47728 = (inp[9]) ? node47736 : node47729;
															assign node47729 = (inp[12]) ? node47733 : node47730;
																assign node47730 = (inp[4]) ? 4'b0000 : 4'b0100;
																assign node47733 = (inp[4]) ? 4'b0100 : 4'b0000;
															assign node47736 = (inp[12]) ? node47738 : 4'b0000;
																assign node47738 = (inp[4]) ? 4'b0000 : 4'b0100;
													assign node47741 = (inp[12]) ? node47747 : node47742;
														assign node47742 = (inp[4]) ? 4'b0000 : node47743;
															assign node47743 = (inp[9]) ? 4'b0000 : 4'b0100;
														assign node47747 = (inp[4]) ? node47749 : 4'b0110;
															assign node47749 = (inp[9]) ? 4'b0010 : 4'b0110;
											assign node47752 = (inp[0]) ? node47784 : node47753;
												assign node47753 = (inp[5]) ? node47767 : node47754;
													assign node47754 = (inp[12]) ? node47760 : node47755;
														assign node47755 = (inp[14]) ? 4'b0010 : node47756;
															assign node47756 = (inp[9]) ? 4'b0100 : 4'b0010;
														assign node47760 = (inp[9]) ? node47764 : node47761;
															assign node47761 = (inp[4]) ? 4'b0100 : 4'b0010;
															assign node47764 = (inp[4]) ? 4'b0000 : 4'b0100;
													assign node47767 = (inp[12]) ? node47773 : node47768;
														assign node47768 = (inp[9]) ? 4'b0100 : node47769;
															assign node47769 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node47773 = (inp[14]) ? node47779 : node47774;
															assign node47774 = (inp[4]) ? node47776 : 4'b0000;
																assign node47776 = (inp[9]) ? 4'b0000 : 4'b0100;
															assign node47779 = (inp[4]) ? 4'b0000 : node47780;
																assign node47780 = (inp[9]) ? 4'b0100 : 4'b0000;
												assign node47784 = (inp[5]) ? node47798 : node47785;
													assign node47785 = (inp[4]) ? node47791 : node47786;
														assign node47786 = (inp[14]) ? node47788 : 4'b0000;
															assign node47788 = (inp[12]) ? 4'b0000 : 4'b0100;
														assign node47791 = (inp[12]) ? node47795 : node47792;
															assign node47792 = (inp[9]) ? 4'b0110 : 4'b0000;
															assign node47795 = (inp[9]) ? 4'b0010 : 4'b0110;
													assign node47798 = (inp[4]) ? node47806 : node47799;
														assign node47799 = (inp[12]) ? node47803 : node47800;
															assign node47800 = (inp[9]) ? 4'b0010 : 4'b0110;
															assign node47803 = (inp[9]) ? 4'b0110 : 4'b0010;
														assign node47806 = (inp[12]) ? 4'b0110 : node47807;
															assign node47807 = (inp[9]) ? 4'b0110 : 4'b0010;
										assign node47811 = (inp[5]) ? node47869 : node47812;
											assign node47812 = (inp[0]) ? node47842 : node47813;
												assign node47813 = (inp[3]) ? node47829 : node47814;
													assign node47814 = (inp[4]) ? node47824 : node47815;
														assign node47815 = (inp[14]) ? node47821 : node47816;
															assign node47816 = (inp[12]) ? node47818 : 4'b0000;
																assign node47818 = (inp[9]) ? 4'b0100 : 4'b0000;
															assign node47821 = (inp[9]) ? 4'b0000 : 4'b0100;
														assign node47824 = (inp[12]) ? 4'b0100 : node47825;
															assign node47825 = (inp[9]) ? 4'b0100 : 4'b0000;
													assign node47829 = (inp[9]) ? node47837 : node47830;
														assign node47830 = (inp[4]) ? node47834 : node47831;
															assign node47831 = (inp[12]) ? 4'b0000 : 4'b0100;
															assign node47834 = (inp[12]) ? 4'b0110 : 4'b0000;
														assign node47837 = (inp[14]) ? node47839 : 4'b0110;
															assign node47839 = (inp[4]) ? 4'b0010 : 4'b0110;
												assign node47842 = (inp[3]) ? node47858 : node47843;
													assign node47843 = (inp[4]) ? node47849 : node47844;
														assign node47844 = (inp[12]) ? node47846 : 4'b0010;
															assign node47846 = (inp[9]) ? 4'b0110 : 4'b0010;
														assign node47849 = (inp[14]) ? node47853 : node47850;
															assign node47850 = (inp[12]) ? 4'b0110 : 4'b0010;
															assign node47853 = (inp[9]) ? node47855 : 4'b0110;
																assign node47855 = (inp[12]) ? 4'b0010 : 4'b0110;
													assign node47858 = (inp[12]) ? node47866 : node47859;
														assign node47859 = (inp[4]) ? node47863 : node47860;
															assign node47860 = (inp[9]) ? 4'b0010 : 4'b0110;
															assign node47863 = (inp[9]) ? 4'b0100 : 4'b0010;
														assign node47866 = (inp[14]) ? 4'b0000 : 4'b0100;
											assign node47869 = (inp[0]) ? node47895 : node47870;
												assign node47870 = (inp[3]) ? node47880 : node47871;
													assign node47871 = (inp[9]) ? 4'b0110 : node47872;
														assign node47872 = (inp[4]) ? node47876 : node47873;
															assign node47873 = (inp[12]) ? 4'b0000 : 4'b0100;
															assign node47876 = (inp[12]) ? 4'b0110 : 4'b0000;
													assign node47880 = (inp[9]) ? node47886 : node47881;
														assign node47881 = (inp[4]) ? node47883 : 4'b0110;
															assign node47883 = (inp[12]) ? 4'b0110 : 4'b0010;
														assign node47886 = (inp[14]) ? node47892 : node47887;
															assign node47887 = (inp[12]) ? node47889 : 4'b0110;
																assign node47889 = (inp[4]) ? 4'b0010 : 4'b0110;
															assign node47892 = (inp[4]) ? 4'b0110 : 4'b0010;
												assign node47895 = (inp[3]) ? node47907 : node47896;
													assign node47896 = (inp[14]) ? 4'b0100 : node47897;
														assign node47897 = (inp[4]) ? node47903 : node47898;
															assign node47898 = (inp[12]) ? 4'b0010 : node47899;
																assign node47899 = (inp[9]) ? 4'b0010 : 4'b0110;
															assign node47903 = (inp[12]) ? 4'b0000 : 4'b0100;
													assign node47907 = (inp[14]) ? node47921 : node47908;
														assign node47908 = (inp[4]) ? node47916 : node47909;
															assign node47909 = (inp[12]) ? node47913 : node47910;
																assign node47910 = (inp[9]) ? 4'b0000 : 4'b0100;
																assign node47913 = (inp[9]) ? 4'b0100 : 4'b0000;
															assign node47916 = (inp[9]) ? node47918 : 4'b0000;
																assign node47918 = (inp[12]) ? 4'b0000 : 4'b0100;
														assign node47921 = (inp[4]) ? node47927 : node47922;
															assign node47922 = (inp[12]) ? 4'b0100 : node47923;
																assign node47923 = (inp[9]) ? 4'b0000 : 4'b0100;
															assign node47927 = (inp[12]) ? node47931 : node47928;
																assign node47928 = (inp[9]) ? 4'b0100 : 4'b0000;
																assign node47931 = (inp[9]) ? 4'b0000 : 4'b0100;
								assign node47934 = (inp[14]) ? node48214 : node47935;
									assign node47935 = (inp[2]) ? node48089 : node47936;
										assign node47936 = (inp[5]) ? node48012 : node47937;
											assign node47937 = (inp[15]) ? node47967 : node47938;
												assign node47938 = (inp[0]) ? node47954 : node47939;
													assign node47939 = (inp[3]) ? node47947 : node47940;
														assign node47940 = (inp[12]) ? node47942 : 4'b0110;
															assign node47942 = (inp[4]) ? node47944 : 4'b0110;
																assign node47944 = (inp[9]) ? 4'b0010 : 4'b0110;
														assign node47947 = (inp[4]) ? node47949 : 4'b0010;
															assign node47949 = (inp[12]) ? 4'b0100 : node47950;
																assign node47950 = (inp[9]) ? 4'b0100 : 4'b0010;
													assign node47954 = (inp[9]) ? node47960 : node47955;
														assign node47955 = (inp[4]) ? 4'b0100 : node47956;
															assign node47956 = (inp[3]) ? 4'b0100 : 4'b0000;
														assign node47960 = (inp[3]) ? node47962 : 4'b0100;
															assign node47962 = (inp[4]) ? node47964 : 4'b0110;
																assign node47964 = (inp[12]) ? 4'b0010 : 4'b0110;
												assign node47967 = (inp[0]) ? node47991 : node47968;
													assign node47968 = (inp[3]) ? node47982 : node47969;
														assign node47969 = (inp[12]) ? node47975 : node47970;
															assign node47970 = (inp[9]) ? 4'b0000 : node47971;
																assign node47971 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node47975 = (inp[9]) ? node47979 : node47976;
																assign node47976 = (inp[4]) ? 4'b0100 : 4'b0000;
																assign node47979 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node47982 = (inp[4]) ? node47986 : node47983;
															assign node47983 = (inp[9]) ? 4'b0000 : 4'b0100;
															assign node47986 = (inp[12]) ? node47988 : 4'b0110;
																assign node47988 = (inp[9]) ? 4'b0010 : 4'b0110;
													assign node47991 = (inp[3]) ? node47999 : node47992;
														assign node47992 = (inp[9]) ? node47994 : 4'b0110;
															assign node47994 = (inp[4]) ? node47996 : 4'b0010;
																assign node47996 = (inp[12]) ? 4'b0010 : 4'b0110;
														assign node47999 = (inp[4]) ? node48007 : node48000;
															assign node48000 = (inp[12]) ? node48004 : node48001;
																assign node48001 = (inp[9]) ? 4'b0010 : 4'b0110;
																assign node48004 = (inp[9]) ? 4'b0100 : 4'b0010;
															assign node48007 = (inp[9]) ? 4'b0100 : node48008;
																assign node48008 = (inp[12]) ? 4'b0100 : 4'b0010;
											assign node48012 = (inp[15]) ? node48056 : node48013;
												assign node48013 = (inp[0]) ? node48035 : node48014;
													assign node48014 = (inp[3]) ? node48026 : node48015;
														assign node48015 = (inp[4]) ? node48023 : node48016;
															assign node48016 = (inp[9]) ? node48020 : node48017;
																assign node48017 = (inp[12]) ? 4'b0010 : 4'b0110;
																assign node48020 = (inp[12]) ? 4'b0100 : 4'b0010;
															assign node48023 = (inp[12]) ? 4'b0000 : 4'b0100;
														assign node48026 = (inp[12]) ? node48028 : 4'b0100;
															assign node48028 = (inp[4]) ? node48032 : node48029;
																assign node48029 = (inp[9]) ? 4'b0100 : 4'b0000;
																assign node48032 = (inp[9]) ? 4'b0000 : 4'b0100;
													assign node48035 = (inp[3]) ? node48049 : node48036;
														assign node48036 = (inp[12]) ? node48042 : node48037;
															assign node48037 = (inp[9]) ? 4'b0000 : node48038;
																assign node48038 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node48042 = (inp[9]) ? node48046 : node48043;
																assign node48043 = (inp[4]) ? 4'b0110 : 4'b0000;
																assign node48046 = (inp[4]) ? 4'b0010 : 4'b0110;
														assign node48049 = (inp[12]) ? 4'b0110 : node48050;
															assign node48050 = (inp[4]) ? 4'b0010 : node48051;
																assign node48051 = (inp[9]) ? 4'b0010 : 4'b0110;
												assign node48056 = (inp[0]) ? node48074 : node48057;
													assign node48057 = (inp[3]) ? node48069 : node48058;
														assign node48058 = (inp[4]) ? node48064 : node48059;
															assign node48059 = (inp[12]) ? 4'b0110 : node48060;
																assign node48060 = (inp[9]) ? 4'b0000 : 4'b0100;
															assign node48064 = (inp[12]) ? node48066 : 4'b0110;
																assign node48066 = (inp[9]) ? 4'b0010 : 4'b0110;
														assign node48069 = (inp[9]) ? node48071 : 4'b0010;
															assign node48071 = (inp[12]) ? 4'b0110 : 4'b0010;
													assign node48074 = (inp[3]) ? node48080 : node48075;
														assign node48075 = (inp[9]) ? node48077 : 4'b0010;
															assign node48077 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node48080 = (inp[12]) ? node48082 : 4'b0000;
															assign node48082 = (inp[9]) ? node48086 : node48083;
																assign node48083 = (inp[4]) ? 4'b0100 : 4'b0000;
																assign node48086 = (inp[4]) ? 4'b0000 : 4'b0100;
										assign node48089 = (inp[0]) ? node48151 : node48090;
											assign node48090 = (inp[4]) ? node48122 : node48091;
												assign node48091 = (inp[15]) ? node48103 : node48092;
													assign node48092 = (inp[3]) ? node48098 : node48093;
														assign node48093 = (inp[12]) ? 4'b0011 : node48094;
															assign node48094 = (inp[9]) ? 4'b0011 : 4'b0111;
														assign node48098 = (inp[5]) ? 4'b0101 : node48099;
															assign node48099 = (inp[12]) ? 4'b0101 : 4'b0011;
													assign node48103 = (inp[3]) ? node48111 : node48104;
														assign node48104 = (inp[5]) ? node48106 : 4'b0101;
															assign node48106 = (inp[9]) ? 4'b0001 : node48107;
																assign node48107 = (inp[12]) ? 4'b0001 : 4'b0101;
														assign node48111 = (inp[5]) ? node48117 : node48112;
															assign node48112 = (inp[12]) ? 4'b0001 : node48113;
																assign node48113 = (inp[9]) ? 4'b0001 : 4'b0101;
															assign node48117 = (inp[9]) ? 4'b0011 : node48118;
																assign node48118 = (inp[12]) ? 4'b0011 : 4'b0111;
												assign node48122 = (inp[15]) ? node48140 : node48123;
													assign node48123 = (inp[5]) ? node48131 : node48124;
														assign node48124 = (inp[9]) ? node48126 : 4'b0011;
															assign node48126 = (inp[3]) ? 4'b0101 : node48127;
																assign node48127 = (inp[12]) ? 4'b0011 : 4'b0111;
														assign node48131 = (inp[3]) ? 4'b0001 : node48132;
															assign node48132 = (inp[9]) ? node48136 : node48133;
																assign node48133 = (inp[12]) ? 4'b0101 : 4'b0011;
																assign node48136 = (inp[12]) ? 4'b0001 : 4'b0101;
													assign node48140 = (inp[9]) ? 4'b0011 : node48141;
														assign node48141 = (inp[12]) ? node48145 : node48142;
															assign node48142 = (inp[3]) ? 4'b0011 : 4'b0001;
															assign node48145 = (inp[5]) ? 4'b0111 : node48146;
																assign node48146 = (inp[3]) ? 4'b0111 : 4'b0101;
											assign node48151 = (inp[15]) ? node48187 : node48152;
												assign node48152 = (inp[3]) ? node48170 : node48153;
													assign node48153 = (inp[9]) ? node48161 : node48154;
														assign node48154 = (inp[4]) ? node48158 : node48155;
															assign node48155 = (inp[12]) ? 4'b0001 : 4'b0101;
															assign node48158 = (inp[12]) ? 4'b0101 : 4'b0001;
														assign node48161 = (inp[4]) ? node48165 : node48162;
															assign node48162 = (inp[12]) ? 4'b0101 : 4'b0001;
															assign node48165 = (inp[5]) ? node48167 : 4'b0001;
																assign node48167 = (inp[12]) ? 4'b0011 : 4'b0111;
													assign node48170 = (inp[12]) ? node48180 : node48171;
														assign node48171 = (inp[5]) ? 4'b0011 : node48172;
															assign node48172 = (inp[9]) ? node48176 : node48173;
																assign node48173 = (inp[4]) ? 4'b0001 : 4'b0101;
																assign node48176 = (inp[4]) ? 4'b0111 : 4'b0001;
														assign node48180 = (inp[9]) ? node48184 : node48181;
															assign node48181 = (inp[4]) ? 4'b0111 : 4'b0011;
															assign node48184 = (inp[5]) ? 4'b0111 : 4'b0011;
												assign node48187 = (inp[5]) ? node48197 : node48188;
													assign node48188 = (inp[4]) ? node48194 : node48189;
														assign node48189 = (inp[3]) ? node48191 : 4'b0111;
															assign node48191 = (inp[12]) ? 4'b0011 : 4'b0111;
														assign node48194 = (inp[3]) ? 4'b0101 : 4'b0111;
													assign node48197 = (inp[4]) ? node48209 : node48198;
														assign node48198 = (inp[3]) ? node48202 : node48199;
															assign node48199 = (inp[12]) ? 4'b0011 : 4'b0111;
															assign node48202 = (inp[9]) ? node48206 : node48203;
																assign node48203 = (inp[12]) ? 4'b0001 : 4'b0101;
																assign node48206 = (inp[12]) ? 4'b0101 : 4'b0001;
														assign node48209 = (inp[9]) ? node48211 : 4'b0101;
															assign node48211 = (inp[12]) ? 4'b0001 : 4'b0101;
									assign node48214 = (inp[0]) ? node48332 : node48215;
										assign node48215 = (inp[12]) ? node48259 : node48216;
											assign node48216 = (inp[15]) ? node48238 : node48217;
												assign node48217 = (inp[3]) ? node48225 : node48218;
													assign node48218 = (inp[4]) ? node48222 : node48219;
														assign node48219 = (inp[9]) ? 4'b0011 : 4'b0111;
														assign node48222 = (inp[9]) ? 4'b0111 : 4'b0011;
													assign node48225 = (inp[5]) ? node48233 : node48226;
														assign node48226 = (inp[2]) ? node48228 : 4'b0011;
															assign node48228 = (inp[4]) ? 4'b0101 : node48229;
																assign node48229 = (inp[9]) ? 4'b0011 : 4'b0111;
														assign node48233 = (inp[9]) ? node48235 : 4'b0001;
															assign node48235 = (inp[4]) ? 4'b0101 : 4'b0001;
												assign node48238 = (inp[3]) ? node48246 : node48239;
													assign node48239 = (inp[2]) ? node48241 : 4'b0001;
														assign node48241 = (inp[4]) ? 4'b0001 : node48242;
															assign node48242 = (inp[9]) ? 4'b0001 : 4'b0101;
													assign node48246 = (inp[5]) ? node48254 : node48247;
														assign node48247 = (inp[9]) ? node48251 : node48248;
															assign node48248 = (inp[4]) ? 4'b0001 : 4'b0101;
															assign node48251 = (inp[4]) ? 4'b0111 : 4'b0001;
														assign node48254 = (inp[4]) ? 4'b0111 : node48255;
															assign node48255 = (inp[9]) ? 4'b0011 : 4'b0111;
											assign node48259 = (inp[15]) ? node48289 : node48260;
												assign node48260 = (inp[3]) ? node48274 : node48261;
													assign node48261 = (inp[5]) ? node48267 : node48262;
														assign node48262 = (inp[4]) ? node48264 : 4'b0011;
															assign node48264 = (inp[9]) ? 4'b0011 : 4'b0111;
														assign node48267 = (inp[4]) ? node48271 : node48268;
															assign node48268 = (inp[9]) ? 4'b0101 : 4'b0011;
															assign node48271 = (inp[9]) ? 4'b0001 : 4'b0101;
													assign node48274 = (inp[5]) ? node48280 : node48275;
														assign node48275 = (inp[9]) ? node48277 : 4'b0101;
															assign node48277 = (inp[4]) ? 4'b0001 : 4'b0101;
														assign node48280 = (inp[2]) ? node48286 : node48281;
															assign node48281 = (inp[9]) ? 4'b0001 : node48282;
																assign node48282 = (inp[4]) ? 4'b0101 : 4'b0001;
															assign node48286 = (inp[9]) ? 4'b0101 : 4'b0001;
												assign node48289 = (inp[5]) ? node48313 : node48290;
													assign node48290 = (inp[3]) ? node48306 : node48291;
														assign node48291 = (inp[2]) ? node48299 : node48292;
															assign node48292 = (inp[9]) ? node48296 : node48293;
																assign node48293 = (inp[4]) ? 4'b0101 : 4'b0001;
																assign node48296 = (inp[4]) ? 4'b0001 : 4'b0101;
															assign node48299 = (inp[4]) ? node48303 : node48300;
																assign node48300 = (inp[9]) ? 4'b0101 : 4'b0001;
																assign node48303 = (inp[9]) ? 4'b0001 : 4'b0101;
														assign node48306 = (inp[4]) ? node48310 : node48307;
															assign node48307 = (inp[9]) ? 4'b0111 : 4'b0001;
															assign node48310 = (inp[9]) ? 4'b0011 : 4'b0111;
													assign node48313 = (inp[3]) ? node48321 : node48314;
														assign node48314 = (inp[9]) ? node48318 : node48315;
															assign node48315 = (inp[4]) ? 4'b0111 : 4'b0001;
															assign node48318 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node48321 = (inp[2]) ? node48327 : node48322;
															assign node48322 = (inp[9]) ? 4'b0011 : node48323;
																assign node48323 = (inp[4]) ? 4'b0111 : 4'b0011;
															assign node48327 = (inp[9]) ? node48329 : 4'b0011;
																assign node48329 = (inp[4]) ? 4'b0011 : 4'b0111;
										assign node48332 = (inp[2]) ? node48414 : node48333;
											assign node48333 = (inp[9]) ? node48373 : node48334;
												assign node48334 = (inp[15]) ? node48350 : node48335;
													assign node48335 = (inp[3]) ? node48341 : node48336;
														assign node48336 = (inp[12]) ? 4'b0001 : node48337;
															assign node48337 = (inp[4]) ? 4'b0001 : 4'b0101;
														assign node48341 = (inp[4]) ? node48347 : node48342;
															assign node48342 = (inp[5]) ? 4'b0111 : node48343;
																assign node48343 = (inp[12]) ? 4'b0001 : 4'b0101;
															assign node48347 = (inp[12]) ? 4'b0111 : 4'b0011;
													assign node48350 = (inp[5]) ? node48360 : node48351;
														assign node48351 = (inp[4]) ? node48355 : node48352;
															assign node48352 = (inp[12]) ? 4'b0011 : 4'b0111;
															assign node48355 = (inp[12]) ? node48357 : 4'b0011;
																assign node48357 = (inp[3]) ? 4'b0101 : 4'b0111;
														assign node48360 = (inp[3]) ? node48368 : node48361;
															assign node48361 = (inp[12]) ? node48365 : node48362;
																assign node48362 = (inp[4]) ? 4'b0011 : 4'b0111;
																assign node48365 = (inp[4]) ? 4'b0101 : 4'b0011;
															assign node48368 = (inp[4]) ? 4'b0001 : node48369;
																assign node48369 = (inp[12]) ? 4'b0001 : 4'b0101;
												assign node48373 = (inp[15]) ? node48395 : node48374;
													assign node48374 = (inp[5]) ? node48388 : node48375;
														assign node48375 = (inp[3]) ? node48383 : node48376;
															assign node48376 = (inp[4]) ? node48380 : node48377;
																assign node48377 = (inp[12]) ? 4'b0101 : 4'b0001;
																assign node48380 = (inp[12]) ? 4'b0001 : 4'b0101;
															assign node48383 = (inp[12]) ? node48385 : 4'b0001;
																assign node48385 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node48388 = (inp[4]) ? node48392 : node48389;
															assign node48389 = (inp[12]) ? 4'b0111 : 4'b0011;
															assign node48392 = (inp[12]) ? 4'b0011 : 4'b0111;
													assign node48395 = (inp[5]) ? node48407 : node48396;
														assign node48396 = (inp[3]) ? node48402 : node48397;
															assign node48397 = (inp[12]) ? 4'b0111 : node48398;
																assign node48398 = (inp[4]) ? 4'b0111 : 4'b0011;
															assign node48402 = (inp[4]) ? node48404 : 4'b0101;
																assign node48404 = (inp[12]) ? 4'b0001 : 4'b0101;
														assign node48407 = (inp[12]) ? node48411 : node48408;
															assign node48408 = (inp[4]) ? 4'b0101 : 4'b0001;
															assign node48411 = (inp[4]) ? 4'b0001 : 4'b0101;
											assign node48414 = (inp[9]) ? node48450 : node48415;
												assign node48415 = (inp[15]) ? node48435 : node48416;
													assign node48416 = (inp[5]) ? node48426 : node48417;
														assign node48417 = (inp[4]) ? node48421 : node48418;
															assign node48418 = (inp[12]) ? 4'b0001 : 4'b0101;
															assign node48421 = (inp[12]) ? node48423 : 4'b0001;
																assign node48423 = (inp[3]) ? 4'b0111 : 4'b0101;
														assign node48426 = (inp[3]) ? node48430 : node48427;
															assign node48427 = (inp[4]) ? 4'b0111 : 4'b0001;
															assign node48430 = (inp[12]) ? 4'b0111 : node48431;
																assign node48431 = (inp[4]) ? 4'b0011 : 4'b0111;
													assign node48435 = (inp[5]) ? node48443 : node48436;
														assign node48436 = (inp[3]) ? node48438 : 4'b0111;
															assign node48438 = (inp[12]) ? 4'b0011 : node48439;
																assign node48439 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node48443 = (inp[4]) ? 4'b0101 : node48444;
															assign node48444 = (inp[12]) ? 4'b0011 : node48445;
																assign node48445 = (inp[3]) ? 4'b0101 : 4'b0111;
												assign node48450 = (inp[15]) ? node48464 : node48451;
													assign node48451 = (inp[3]) ? node48457 : node48452;
														assign node48452 = (inp[12]) ? node48454 : 4'b0001;
															assign node48454 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node48457 = (inp[5]) ? node48461 : node48458;
															assign node48458 = (inp[4]) ? 4'b0011 : 4'b0111;
															assign node48461 = (inp[4]) ? 4'b0111 : 4'b0011;
													assign node48464 = (inp[3]) ? node48470 : node48465;
														assign node48465 = (inp[12]) ? 4'b0001 : node48466;
															assign node48466 = (inp[4]) ? 4'b0111 : 4'b0011;
														assign node48470 = (inp[4]) ? node48476 : node48471;
															assign node48471 = (inp[12]) ? 4'b0101 : node48472;
																assign node48472 = (inp[5]) ? 4'b0001 : 4'b0011;
															assign node48476 = (inp[12]) ? 4'b0001 : 4'b0101;
							assign node48479 = (inp[7]) ? node49021 : node48480;
								assign node48480 = (inp[2]) ? node48786 : node48481;
									assign node48481 = (inp[14]) ? node48639 : node48482;
										assign node48482 = (inp[15]) ? node48574 : node48483;
											assign node48483 = (inp[0]) ? node48519 : node48484;
												assign node48484 = (inp[5]) ? node48500 : node48485;
													assign node48485 = (inp[12]) ? node48493 : node48486;
														assign node48486 = (inp[4]) ? node48490 : node48487;
															assign node48487 = (inp[9]) ? 4'b0010 : 4'b0110;
															assign node48490 = (inp[9]) ? 4'b0110 : 4'b0010;
														assign node48493 = (inp[4]) ? node48495 : 4'b0010;
															assign node48495 = (inp[9]) ? node48497 : 4'b0100;
																assign node48497 = (inp[3]) ? 4'b0000 : 4'b0010;
													assign node48500 = (inp[3]) ? node48512 : node48501;
														assign node48501 = (inp[9]) ? node48507 : node48502;
															assign node48502 = (inp[4]) ? 4'b0010 : node48503;
																assign node48503 = (inp[12]) ? 4'b0010 : 4'b0110;
															assign node48507 = (inp[4]) ? node48509 : 4'b0010;
																assign node48509 = (inp[12]) ? 4'b0000 : 4'b0100;
														assign node48512 = (inp[12]) ? 4'b0000 : node48513;
															assign node48513 = (inp[9]) ? 4'b0000 : node48514;
																assign node48514 = (inp[4]) ? 4'b0000 : 4'b0100;
												assign node48519 = (inp[3]) ? node48549 : node48520;
													assign node48520 = (inp[5]) ? node48534 : node48521;
														assign node48521 = (inp[12]) ? node48529 : node48522;
															assign node48522 = (inp[9]) ? node48526 : node48523;
																assign node48523 = (inp[4]) ? 4'b0000 : 4'b0100;
																assign node48526 = (inp[4]) ? 4'b0100 : 4'b0000;
															assign node48529 = (inp[4]) ? node48531 : 4'b0100;
																assign node48531 = (inp[9]) ? 4'b0000 : 4'b0100;
														assign node48534 = (inp[9]) ? node48542 : node48535;
															assign node48535 = (inp[4]) ? node48539 : node48536;
																assign node48536 = (inp[12]) ? 4'b0000 : 4'b0100;
																assign node48539 = (inp[12]) ? 4'b0110 : 4'b0000;
															assign node48542 = (inp[12]) ? node48546 : node48543;
																assign node48543 = (inp[4]) ? 4'b0110 : 4'b0000;
																assign node48546 = (inp[4]) ? 4'b0010 : 4'b0110;
													assign node48549 = (inp[5]) ? node48559 : node48550;
														assign node48550 = (inp[12]) ? node48552 : 4'b0100;
															assign node48552 = (inp[9]) ? node48556 : node48553;
																assign node48553 = (inp[4]) ? 4'b0110 : 4'b0000;
																assign node48556 = (inp[4]) ? 4'b0010 : 4'b0110;
														assign node48559 = (inp[4]) ? node48567 : node48560;
															assign node48560 = (inp[9]) ? node48564 : node48561;
																assign node48561 = (inp[12]) ? 4'b0010 : 4'b0110;
																assign node48564 = (inp[12]) ? 4'b0110 : 4'b0010;
															assign node48567 = (inp[12]) ? node48571 : node48568;
																assign node48568 = (inp[9]) ? 4'b0110 : 4'b0010;
																assign node48571 = (inp[9]) ? 4'b0010 : 4'b0110;
											assign node48574 = (inp[5]) ? node48608 : node48575;
												assign node48575 = (inp[0]) ? node48597 : node48576;
													assign node48576 = (inp[3]) ? node48586 : node48577;
														assign node48577 = (inp[9]) ? 4'b0100 : node48578;
															assign node48578 = (inp[12]) ? node48582 : node48579;
																assign node48579 = (inp[4]) ? 4'b0000 : 4'b0100;
																assign node48582 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node48586 = (inp[4]) ? node48592 : node48587;
															assign node48587 = (inp[9]) ? 4'b0000 : node48588;
																assign node48588 = (inp[12]) ? 4'b0000 : 4'b0100;
															assign node48592 = (inp[9]) ? node48594 : 4'b0000;
																assign node48594 = (inp[12]) ? 4'b0010 : 4'b0110;
													assign node48597 = (inp[3]) ? node48599 : 4'b0010;
														assign node48599 = (inp[9]) ? node48603 : node48600;
															assign node48600 = (inp[12]) ? 4'b0010 : 4'b0110;
															assign node48603 = (inp[4]) ? node48605 : 4'b0100;
																assign node48605 = (inp[12]) ? 4'b0000 : 4'b0100;
												assign node48608 = (inp[0]) ? node48622 : node48609;
													assign node48609 = (inp[12]) ? node48615 : node48610;
														assign node48610 = (inp[3]) ? 4'b0010 : node48611;
															assign node48611 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node48615 = (inp[3]) ? 4'b0110 : node48616;
															assign node48616 = (inp[4]) ? 4'b0110 : node48617;
																assign node48617 = (inp[9]) ? 4'b0110 : 4'b0000;
													assign node48622 = (inp[3]) ? node48632 : node48623;
														assign node48623 = (inp[12]) ? 4'b0100 : node48624;
															assign node48624 = (inp[9]) ? node48628 : node48625;
																assign node48625 = (inp[4]) ? 4'b0010 : 4'b0110;
																assign node48628 = (inp[4]) ? 4'b0100 : 4'b0010;
														assign node48632 = (inp[9]) ? node48634 : 4'b0100;
															assign node48634 = (inp[12]) ? node48636 : 4'b0100;
																assign node48636 = (inp[4]) ? 4'b0000 : 4'b0100;
										assign node48639 = (inp[12]) ? node48719 : node48640;
											assign node48640 = (inp[3]) ? node48670 : node48641;
												assign node48641 = (inp[4]) ? node48653 : node48642;
													assign node48642 = (inp[9]) ? node48650 : node48643;
														assign node48643 = (inp[15]) ? node48647 : node48644;
															assign node48644 = (inp[0]) ? 4'b0101 : 4'b0111;
															assign node48647 = (inp[0]) ? 4'b0111 : 4'b0101;
														assign node48650 = (inp[5]) ? 4'b0001 : 4'b0011;
													assign node48653 = (inp[9]) ? node48661 : node48654;
														assign node48654 = (inp[5]) ? 4'b0011 : node48655;
															assign node48655 = (inp[0]) ? node48657 : 4'b0001;
																assign node48657 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node48661 = (inp[0]) ? node48663 : 4'b0111;
															assign node48663 = (inp[15]) ? node48667 : node48664;
																assign node48664 = (inp[5]) ? 4'b0111 : 4'b0101;
																assign node48667 = (inp[5]) ? 4'b0101 : 4'b0111;
												assign node48670 = (inp[5]) ? node48698 : node48671;
													assign node48671 = (inp[15]) ? node48685 : node48672;
														assign node48672 = (inp[0]) ? node48680 : node48673;
															assign node48673 = (inp[4]) ? node48677 : node48674;
																assign node48674 = (inp[9]) ? 4'b0011 : 4'b0111;
																assign node48677 = (inp[9]) ? 4'b0101 : 4'b0011;
															assign node48680 = (inp[9]) ? 4'b0111 : node48681;
																assign node48681 = (inp[4]) ? 4'b0001 : 4'b0101;
														assign node48685 = (inp[0]) ? node48691 : node48686;
															assign node48686 = (inp[4]) ? 4'b0111 : node48687;
																assign node48687 = (inp[9]) ? 4'b0001 : 4'b0101;
															assign node48691 = (inp[4]) ? node48695 : node48692;
																assign node48692 = (inp[9]) ? 4'b0011 : 4'b0111;
																assign node48695 = (inp[9]) ? 4'b0101 : 4'b0011;
													assign node48698 = (inp[4]) ? node48706 : node48699;
														assign node48699 = (inp[9]) ? node48701 : 4'b0111;
															assign node48701 = (inp[15]) ? node48703 : 4'b0001;
																assign node48703 = (inp[0]) ? 4'b0001 : 4'b0011;
														assign node48706 = (inp[9]) ? node48712 : node48707;
															assign node48707 = (inp[0]) ? node48709 : 4'b0001;
																assign node48709 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node48712 = (inp[0]) ? node48716 : node48713;
																assign node48713 = (inp[15]) ? 4'b0111 : 4'b0101;
																assign node48716 = (inp[15]) ? 4'b0101 : 4'b0111;
											assign node48719 = (inp[5]) ? node48759 : node48720;
												assign node48720 = (inp[4]) ? node48738 : node48721;
													assign node48721 = (inp[9]) ? node48729 : node48722;
														assign node48722 = (inp[15]) ? node48726 : node48723;
															assign node48723 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node48726 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node48729 = (inp[15]) ? node48731 : 4'b0101;
															assign node48731 = (inp[0]) ? node48735 : node48732;
																assign node48732 = (inp[3]) ? 4'b0111 : 4'b0101;
																assign node48735 = (inp[3]) ? 4'b0101 : 4'b0111;
													assign node48738 = (inp[9]) ? node48746 : node48739;
														assign node48739 = (inp[0]) ? node48741 : 4'b0101;
															assign node48741 = (inp[15]) ? 4'b0111 : node48742;
																assign node48742 = (inp[3]) ? 4'b0111 : 4'b0101;
														assign node48746 = (inp[3]) ? node48754 : node48747;
															assign node48747 = (inp[15]) ? node48751 : node48748;
																assign node48748 = (inp[0]) ? 4'b0001 : 4'b0011;
																assign node48751 = (inp[0]) ? 4'b0011 : 4'b0001;
															assign node48754 = (inp[15]) ? node48756 : 4'b0011;
																assign node48756 = (inp[0]) ? 4'b0001 : 4'b0011;
												assign node48759 = (inp[15]) ? node48775 : node48760;
													assign node48760 = (inp[0]) ? node48768 : node48761;
														assign node48761 = (inp[3]) ? node48765 : node48762;
															assign node48762 = (inp[9]) ? 4'b0001 : 4'b0011;
															assign node48765 = (inp[4]) ? 4'b0101 : 4'b0001;
														assign node48768 = (inp[9]) ? node48772 : node48769;
															assign node48769 = (inp[4]) ? 4'b0111 : 4'b0011;
															assign node48772 = (inp[4]) ? 4'b0011 : 4'b0111;
													assign node48775 = (inp[0]) ? node48781 : node48776;
														assign node48776 = (inp[9]) ? node48778 : 4'b0111;
															assign node48778 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node48781 = (inp[4]) ? node48783 : 4'b0101;
															assign node48783 = (inp[9]) ? 4'b0001 : 4'b0101;
									assign node48786 = (inp[9]) ? node48894 : node48787;
										assign node48787 = (inp[0]) ? node48843 : node48788;
											assign node48788 = (inp[15]) ? node48816 : node48789;
												assign node48789 = (inp[5]) ? node48799 : node48790;
													assign node48790 = (inp[4]) ? node48794 : node48791;
														assign node48791 = (inp[12]) ? 4'b0011 : 4'b0111;
														assign node48794 = (inp[12]) ? node48796 : 4'b0011;
															assign node48796 = (inp[3]) ? 4'b0101 : 4'b0111;
													assign node48799 = (inp[3]) ? node48809 : node48800;
														assign node48800 = (inp[14]) ? 4'b0011 : node48801;
															assign node48801 = (inp[4]) ? node48805 : node48802;
																assign node48802 = (inp[12]) ? 4'b0011 : 4'b0111;
																assign node48805 = (inp[12]) ? 4'b0101 : 4'b0011;
														assign node48809 = (inp[12]) ? node48813 : node48810;
															assign node48810 = (inp[4]) ? 4'b0001 : 4'b0101;
															assign node48813 = (inp[4]) ? 4'b0101 : 4'b0001;
												assign node48816 = (inp[5]) ? node48832 : node48817;
													assign node48817 = (inp[3]) ? node48825 : node48818;
														assign node48818 = (inp[4]) ? node48822 : node48819;
															assign node48819 = (inp[12]) ? 4'b0001 : 4'b0101;
															assign node48822 = (inp[12]) ? 4'b0101 : 4'b0001;
														assign node48825 = (inp[4]) ? node48829 : node48826;
															assign node48826 = (inp[12]) ? 4'b0001 : 4'b0101;
															assign node48829 = (inp[12]) ? 4'b0111 : 4'b0001;
													assign node48832 = (inp[3]) ? node48836 : node48833;
														assign node48833 = (inp[14]) ? 4'b0111 : 4'b0001;
														assign node48836 = (inp[12]) ? node48840 : node48837;
															assign node48837 = (inp[4]) ? 4'b0011 : 4'b0111;
															assign node48840 = (inp[4]) ? 4'b0111 : 4'b0011;
											assign node48843 = (inp[15]) ? node48863 : node48844;
												assign node48844 = (inp[4]) ? node48852 : node48845;
													assign node48845 = (inp[12]) ? 4'b0001 : node48846;
														assign node48846 = (inp[5]) ? node48848 : 4'b0101;
															assign node48848 = (inp[3]) ? 4'b0111 : 4'b0101;
													assign node48852 = (inp[12]) ? node48858 : node48853;
														assign node48853 = (inp[3]) ? node48855 : 4'b0001;
															assign node48855 = (inp[5]) ? 4'b0011 : 4'b0001;
														assign node48858 = (inp[14]) ? node48860 : 4'b0111;
															assign node48860 = (inp[3]) ? 4'b0111 : 4'b0101;
												assign node48863 = (inp[3]) ? node48873 : node48864;
													assign node48864 = (inp[4]) ? node48868 : node48865;
														assign node48865 = (inp[12]) ? 4'b0011 : 4'b0111;
														assign node48868 = (inp[12]) ? node48870 : 4'b0011;
															assign node48870 = (inp[5]) ? 4'b0101 : 4'b0111;
													assign node48873 = (inp[5]) ? node48881 : node48874;
														assign node48874 = (inp[12]) ? node48878 : node48875;
															assign node48875 = (inp[4]) ? 4'b0011 : 4'b0111;
															assign node48878 = (inp[4]) ? 4'b0101 : 4'b0011;
														assign node48881 = (inp[14]) ? node48889 : node48882;
															assign node48882 = (inp[12]) ? node48886 : node48883;
																assign node48883 = (inp[4]) ? 4'b0001 : 4'b0101;
																assign node48886 = (inp[4]) ? 4'b0101 : 4'b0001;
															assign node48889 = (inp[12]) ? node48891 : 4'b0001;
																assign node48891 = (inp[4]) ? 4'b0101 : 4'b0001;
										assign node48894 = (inp[3]) ? node48964 : node48895;
											assign node48895 = (inp[5]) ? node48919 : node48896;
												assign node48896 = (inp[15]) ? node48910 : node48897;
													assign node48897 = (inp[0]) ? node48905 : node48898;
														assign node48898 = (inp[12]) ? node48902 : node48899;
															assign node48899 = (inp[4]) ? 4'b0111 : 4'b0011;
															assign node48902 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node48905 = (inp[4]) ? node48907 : 4'b0101;
															assign node48907 = (inp[14]) ? 4'b0101 : 4'b0001;
													assign node48910 = (inp[0]) ? node48912 : 4'b0001;
														assign node48912 = (inp[4]) ? node48916 : node48913;
															assign node48913 = (inp[12]) ? 4'b0111 : 4'b0011;
															assign node48916 = (inp[12]) ? 4'b0011 : 4'b0111;
												assign node48919 = (inp[12]) ? node48943 : node48920;
													assign node48920 = (inp[4]) ? node48930 : node48921;
														assign node48921 = (inp[14]) ? node48923 : 4'b0001;
															assign node48923 = (inp[0]) ? node48927 : node48924;
																assign node48924 = (inp[15]) ? 4'b0001 : 4'b0011;
																assign node48927 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node48930 = (inp[14]) ? node48936 : node48931;
															assign node48931 = (inp[0]) ? node48933 : 4'b0101;
																assign node48933 = (inp[15]) ? 4'b0101 : 4'b0111;
															assign node48936 = (inp[0]) ? node48940 : node48937;
																assign node48937 = (inp[15]) ? 4'b0111 : 4'b0101;
																assign node48940 = (inp[15]) ? 4'b0101 : 4'b0111;
													assign node48943 = (inp[4]) ? node48951 : node48944;
														assign node48944 = (inp[0]) ? node48948 : node48945;
															assign node48945 = (inp[15]) ? 4'b0111 : 4'b0101;
															assign node48948 = (inp[15]) ? 4'b0101 : 4'b0111;
														assign node48951 = (inp[14]) ? node48959 : node48952;
															assign node48952 = (inp[15]) ? node48956 : node48953;
																assign node48953 = (inp[0]) ? 4'b0011 : 4'b0001;
																assign node48956 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node48959 = (inp[0]) ? 4'b0011 : node48960;
																assign node48960 = (inp[15]) ? 4'b0011 : 4'b0001;
											assign node48964 = (inp[5]) ? node48992 : node48965;
												assign node48965 = (inp[0]) ? node48975 : node48966;
													assign node48966 = (inp[15]) ? node48968 : 4'b0101;
														assign node48968 = (inp[12]) ? node48972 : node48969;
															assign node48969 = (inp[4]) ? 4'b0111 : 4'b0001;
															assign node48972 = (inp[4]) ? 4'b0011 : 4'b0111;
													assign node48975 = (inp[15]) ? node48985 : node48976;
														assign node48976 = (inp[14]) ? node48978 : 4'b0111;
															assign node48978 = (inp[4]) ? node48982 : node48979;
																assign node48979 = (inp[12]) ? 4'b0111 : 4'b0001;
																assign node48982 = (inp[12]) ? 4'b0011 : 4'b0111;
														assign node48985 = (inp[4]) ? node48989 : node48986;
															assign node48986 = (inp[12]) ? 4'b0101 : 4'b0011;
															assign node48989 = (inp[12]) ? 4'b0001 : 4'b0101;
												assign node48992 = (inp[12]) ? node49008 : node48993;
													assign node48993 = (inp[4]) ? node49001 : node48994;
														assign node48994 = (inp[15]) ? node48998 : node48995;
															assign node48995 = (inp[0]) ? 4'b0011 : 4'b0001;
															assign node48998 = (inp[0]) ? 4'b0001 : 4'b0011;
														assign node49001 = (inp[15]) ? node49005 : node49002;
															assign node49002 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node49005 = (inp[0]) ? 4'b0101 : 4'b0111;
													assign node49008 = (inp[4]) ? node49016 : node49009;
														assign node49009 = (inp[0]) ? node49013 : node49010;
															assign node49010 = (inp[15]) ? 4'b0111 : 4'b0101;
															assign node49013 = (inp[15]) ? 4'b0101 : 4'b0111;
														assign node49016 = (inp[14]) ? node49018 : 4'b0011;
															assign node49018 = (inp[0]) ? 4'b0011 : 4'b0001;
								assign node49021 = (inp[14]) ? node49301 : node49022;
									assign node49022 = (inp[2]) ? node49172 : node49023;
										assign node49023 = (inp[15]) ? node49097 : node49024;
											assign node49024 = (inp[12]) ? node49054 : node49025;
												assign node49025 = (inp[5]) ? node49039 : node49026;
													assign node49026 = (inp[9]) ? node49030 : node49027;
														assign node49027 = (inp[4]) ? 4'b0001 : 4'b0101;
														assign node49030 = (inp[4]) ? node49034 : node49031;
															assign node49031 = (inp[3]) ? 4'b0001 : 4'b0011;
															assign node49034 = (inp[3]) ? node49036 : 4'b0101;
																assign node49036 = (inp[0]) ? 4'b0111 : 4'b0101;
													assign node49039 = (inp[0]) ? node49047 : node49040;
														assign node49040 = (inp[3]) ? 4'b0101 : node49041;
															assign node49041 = (inp[9]) ? 4'b0101 : node49042;
																assign node49042 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node49047 = (inp[9]) ? node49049 : 4'b0001;
															assign node49049 = (inp[4]) ? 4'b0111 : node49050;
																assign node49050 = (inp[3]) ? 4'b0011 : 4'b0001;
												assign node49054 = (inp[5]) ? node49086 : node49055;
													assign node49055 = (inp[0]) ? node49071 : node49056;
														assign node49056 = (inp[3]) ? node49064 : node49057;
															assign node49057 = (inp[4]) ? node49061 : node49058;
																assign node49058 = (inp[9]) ? 4'b0111 : 4'b0011;
																assign node49061 = (inp[9]) ? 4'b0011 : 4'b0111;
															assign node49064 = (inp[9]) ? node49068 : node49065;
																assign node49065 = (inp[4]) ? 4'b0101 : 4'b0011;
																assign node49068 = (inp[4]) ? 4'b0001 : 4'b0101;
														assign node49071 = (inp[3]) ? node49079 : node49072;
															assign node49072 = (inp[4]) ? node49076 : node49073;
																assign node49073 = (inp[9]) ? 4'b0101 : 4'b0001;
																assign node49076 = (inp[9]) ? 4'b0001 : 4'b0101;
															assign node49079 = (inp[4]) ? node49083 : node49080;
																assign node49080 = (inp[9]) ? 4'b0111 : 4'b0001;
																assign node49083 = (inp[9]) ? 4'b0011 : 4'b0111;
													assign node49086 = (inp[0]) ? node49092 : node49087;
														assign node49087 = (inp[9]) ? 4'b0001 : node49088;
															assign node49088 = (inp[3]) ? 4'b0001 : 4'b0011;
														assign node49092 = (inp[9]) ? node49094 : 4'b0001;
															assign node49094 = (inp[4]) ? 4'b0011 : 4'b0111;
											assign node49097 = (inp[4]) ? node49127 : node49098;
												assign node49098 = (inp[5]) ? node49118 : node49099;
													assign node49099 = (inp[0]) ? node49109 : node49100;
														assign node49100 = (inp[12]) ? node49104 : node49101;
															assign node49101 = (inp[9]) ? 4'b0001 : 4'b0101;
															assign node49104 = (inp[9]) ? node49106 : 4'b0001;
																assign node49106 = (inp[3]) ? 4'b0111 : 4'b0101;
														assign node49109 = (inp[9]) ? node49113 : node49110;
															assign node49110 = (inp[12]) ? 4'b0011 : 4'b0111;
															assign node49113 = (inp[12]) ? node49115 : 4'b0011;
																assign node49115 = (inp[3]) ? 4'b0101 : 4'b0111;
													assign node49118 = (inp[9]) ? node49122 : node49119;
														assign node49119 = (inp[12]) ? 4'b0011 : 4'b0111;
														assign node49122 = (inp[12]) ? node49124 : 4'b0011;
															assign node49124 = (inp[0]) ? 4'b0101 : 4'b0111;
												assign node49127 = (inp[3]) ? node49155 : node49128;
													assign node49128 = (inp[0]) ? node49142 : node49129;
														assign node49129 = (inp[5]) ? node49135 : node49130;
															assign node49130 = (inp[12]) ? 4'b0101 : node49131;
																assign node49131 = (inp[9]) ? 4'b0101 : 4'b0001;
															assign node49135 = (inp[12]) ? node49139 : node49136;
																assign node49136 = (inp[9]) ? 4'b0111 : 4'b0001;
																assign node49139 = (inp[9]) ? 4'b0011 : 4'b0111;
														assign node49142 = (inp[5]) ? node49150 : node49143;
															assign node49143 = (inp[9]) ? node49147 : node49144;
																assign node49144 = (inp[12]) ? 4'b0111 : 4'b0011;
																assign node49147 = (inp[12]) ? 4'b0011 : 4'b0111;
															assign node49150 = (inp[12]) ? node49152 : 4'b0011;
																assign node49152 = (inp[9]) ? 4'b0001 : 4'b0101;
													assign node49155 = (inp[0]) ? node49163 : node49156;
														assign node49156 = (inp[5]) ? 4'b0111 : node49157;
															assign node49157 = (inp[12]) ? node49159 : 4'b0001;
																assign node49159 = (inp[9]) ? 4'b0011 : 4'b0111;
														assign node49163 = (inp[5]) ? node49165 : 4'b0101;
															assign node49165 = (inp[12]) ? node49169 : node49166;
																assign node49166 = (inp[9]) ? 4'b0101 : 4'b0001;
																assign node49169 = (inp[9]) ? 4'b0001 : 4'b0101;
										assign node49172 = (inp[12]) ? node49254 : node49173;
											assign node49173 = (inp[5]) ? node49217 : node49174;
												assign node49174 = (inp[3]) ? node49188 : node49175;
													assign node49175 = (inp[4]) ? node49181 : node49176;
														assign node49176 = (inp[9]) ? node49178 : 4'b0100;
															assign node49178 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node49181 = (inp[0]) ? node49185 : node49182;
															assign node49182 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node49185 = (inp[15]) ? 4'b0010 : 4'b0000;
													assign node49188 = (inp[9]) ? node49202 : node49189;
														assign node49189 = (inp[4]) ? node49195 : node49190;
															assign node49190 = (inp[15]) ? node49192 : 4'b0110;
																assign node49192 = (inp[0]) ? 4'b0110 : 4'b0100;
															assign node49195 = (inp[15]) ? node49199 : node49196;
																assign node49196 = (inp[0]) ? 4'b0000 : 4'b0010;
																assign node49199 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node49202 = (inp[4]) ? node49210 : node49203;
															assign node49203 = (inp[15]) ? node49207 : node49204;
																assign node49204 = (inp[0]) ? 4'b0000 : 4'b0010;
																assign node49207 = (inp[0]) ? 4'b0010 : 4'b0000;
															assign node49210 = (inp[15]) ? node49214 : node49211;
																assign node49211 = (inp[0]) ? 4'b0110 : 4'b0100;
																assign node49214 = (inp[0]) ? 4'b0100 : 4'b0110;
												assign node49217 = (inp[9]) ? node49237 : node49218;
													assign node49218 = (inp[4]) ? node49232 : node49219;
														assign node49219 = (inp[0]) ? node49227 : node49220;
															assign node49220 = (inp[3]) ? node49224 : node49221;
																assign node49221 = (inp[15]) ? 4'b0100 : 4'b0110;
																assign node49224 = (inp[15]) ? 4'b0110 : 4'b0100;
															assign node49227 = (inp[15]) ? node49229 : 4'b0110;
																assign node49229 = (inp[3]) ? 4'b0100 : 4'b0110;
														assign node49232 = (inp[0]) ? 4'b0000 : node49233;
															assign node49233 = (inp[15]) ? 4'b0010 : 4'b0000;
													assign node49237 = (inp[4]) ? node49247 : node49238;
														assign node49238 = (inp[0]) ? node49240 : 4'b0000;
															assign node49240 = (inp[3]) ? node49244 : node49241;
																assign node49241 = (inp[15]) ? 4'b0010 : 4'b0000;
																assign node49244 = (inp[15]) ? 4'b0000 : 4'b0010;
														assign node49247 = (inp[0]) ? node49251 : node49248;
															assign node49248 = (inp[15]) ? 4'b0110 : 4'b0100;
															assign node49251 = (inp[15]) ? 4'b0100 : 4'b0110;
											assign node49254 = (inp[4]) ? node49272 : node49255;
												assign node49255 = (inp[9]) ? node49263 : node49256;
													assign node49256 = (inp[0]) ? 4'b0010 : node49257;
														assign node49257 = (inp[15]) ? 4'b0000 : node49258;
															assign node49258 = (inp[5]) ? 4'b0000 : 4'b0010;
													assign node49263 = (inp[3]) ? node49265 : 4'b0110;
														assign node49265 = (inp[0]) ? node49269 : node49266;
															assign node49266 = (inp[15]) ? 4'b0110 : 4'b0100;
															assign node49269 = (inp[15]) ? 4'b0100 : 4'b0110;
												assign node49272 = (inp[9]) ? node49290 : node49273;
													assign node49273 = (inp[5]) ? node49285 : node49274;
														assign node49274 = (inp[15]) ? node49280 : node49275;
															assign node49275 = (inp[0]) ? 4'b0100 : node49276;
																assign node49276 = (inp[3]) ? 4'b0100 : 4'b0110;
															assign node49280 = (inp[3]) ? node49282 : 4'b0110;
																assign node49282 = (inp[0]) ? 4'b0100 : 4'b0110;
														assign node49285 = (inp[0]) ? 4'b0110 : node49286;
															assign node49286 = (inp[15]) ? 4'b0110 : 4'b0100;
													assign node49290 = (inp[15]) ? node49296 : node49291;
														assign node49291 = (inp[0]) ? 4'b0010 : node49292;
															assign node49292 = (inp[5]) ? 4'b0000 : 4'b0010;
														assign node49296 = (inp[0]) ? 4'b0000 : node49297;
															assign node49297 = (inp[5]) ? 4'b0010 : 4'b0000;
									assign node49301 = (inp[9]) ? node49443 : node49302;
										assign node49302 = (inp[3]) ? node49386 : node49303;
											assign node49303 = (inp[2]) ? node49353 : node49304;
												assign node49304 = (inp[5]) ? node49328 : node49305;
													assign node49305 = (inp[0]) ? node49317 : node49306;
														assign node49306 = (inp[15]) ? node49312 : node49307;
															assign node49307 = (inp[12]) ? node49309 : 4'b0010;
																assign node49309 = (inp[4]) ? 4'b0110 : 4'b0010;
															assign node49312 = (inp[4]) ? 4'b0100 : node49313;
																assign node49313 = (inp[12]) ? 4'b0000 : 4'b0100;
														assign node49317 = (inp[15]) ? node49323 : node49318;
															assign node49318 = (inp[12]) ? 4'b0100 : node49319;
																assign node49319 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node49323 = (inp[12]) ? 4'b0010 : node49324;
																assign node49324 = (inp[4]) ? 4'b0010 : 4'b0110;
													assign node49328 = (inp[0]) ? node49342 : node49329;
														assign node49329 = (inp[15]) ? node49335 : node49330;
															assign node49330 = (inp[4]) ? 4'b0100 : node49331;
																assign node49331 = (inp[12]) ? 4'b0010 : 4'b0110;
															assign node49335 = (inp[4]) ? node49339 : node49336;
																assign node49336 = (inp[12]) ? 4'b0000 : 4'b0100;
																assign node49339 = (inp[12]) ? 4'b0110 : 4'b0000;
														assign node49342 = (inp[15]) ? node49348 : node49343;
															assign node49343 = (inp[4]) ? 4'b0110 : node49344;
																assign node49344 = (inp[12]) ? 4'b0000 : 4'b0100;
															assign node49348 = (inp[12]) ? 4'b0100 : node49349;
																assign node49349 = (inp[4]) ? 4'b0010 : 4'b0110;
												assign node49353 = (inp[15]) ? node49371 : node49354;
													assign node49354 = (inp[0]) ? node49364 : node49355;
														assign node49355 = (inp[4]) ? node49359 : node49356;
															assign node49356 = (inp[12]) ? 4'b0010 : 4'b0110;
															assign node49359 = (inp[12]) ? node49361 : 4'b0010;
																assign node49361 = (inp[5]) ? 4'b0100 : 4'b0110;
														assign node49364 = (inp[4]) ? node49366 : 4'b0000;
															assign node49366 = (inp[12]) ? node49368 : 4'b0000;
																assign node49368 = (inp[5]) ? 4'b0110 : 4'b0100;
													assign node49371 = (inp[0]) ? node49377 : node49372;
														assign node49372 = (inp[12]) ? 4'b0110 : node49373;
															assign node49373 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node49377 = (inp[5]) ? node49383 : node49378;
															assign node49378 = (inp[12]) ? node49380 : 4'b0110;
																assign node49380 = (inp[4]) ? 4'b0110 : 4'b0010;
															assign node49383 = (inp[4]) ? 4'b0010 : 4'b0110;
											assign node49386 = (inp[15]) ? node49416 : node49387;
												assign node49387 = (inp[12]) ? node49407 : node49388;
													assign node49388 = (inp[4]) ? node49400 : node49389;
														assign node49389 = (inp[2]) ? node49395 : node49390;
															assign node49390 = (inp[5]) ? node49392 : 4'b0100;
																assign node49392 = (inp[0]) ? 4'b0110 : 4'b0100;
															assign node49395 = (inp[5]) ? 4'b0100 : node49396;
																assign node49396 = (inp[0]) ? 4'b0100 : 4'b0110;
														assign node49400 = (inp[0]) ? node49404 : node49401;
															assign node49401 = (inp[5]) ? 4'b0000 : 4'b0010;
															assign node49404 = (inp[5]) ? 4'b0010 : 4'b0000;
													assign node49407 = (inp[4]) ? node49413 : node49408;
														assign node49408 = (inp[5]) ? 4'b0010 : node49409;
															assign node49409 = (inp[0]) ? 4'b0000 : 4'b0010;
														assign node49413 = (inp[0]) ? 4'b0110 : 4'b0100;
												assign node49416 = (inp[5]) ? node49434 : node49417;
													assign node49417 = (inp[0]) ? node49427 : node49418;
														assign node49418 = (inp[2]) ? node49422 : node49419;
															assign node49419 = (inp[4]) ? 4'b0110 : 4'b0000;
															assign node49422 = (inp[4]) ? 4'b0000 : node49423;
																assign node49423 = (inp[12]) ? 4'b0000 : 4'b0100;
														assign node49427 = (inp[12]) ? node49431 : node49428;
															assign node49428 = (inp[4]) ? 4'b0010 : 4'b0110;
															assign node49431 = (inp[4]) ? 4'b0100 : 4'b0010;
													assign node49434 = (inp[0]) ? 4'b0000 : node49435;
														assign node49435 = (inp[4]) ? node49439 : node49436;
															assign node49436 = (inp[12]) ? 4'b0010 : 4'b0110;
															assign node49439 = (inp[12]) ? 4'b0110 : 4'b0010;
										assign node49443 = (inp[12]) ? node49487 : node49444;
											assign node49444 = (inp[4]) ? node49468 : node49445;
												assign node49445 = (inp[15]) ? node49457 : node49446;
													assign node49446 = (inp[0]) ? node49452 : node49447;
														assign node49447 = (inp[3]) ? node49449 : 4'b0010;
															assign node49449 = (inp[5]) ? 4'b0000 : 4'b0010;
														assign node49452 = (inp[5]) ? node49454 : 4'b0000;
															assign node49454 = (inp[3]) ? 4'b0010 : 4'b0000;
													assign node49457 = (inp[0]) ? node49463 : node49458;
														assign node49458 = (inp[5]) ? node49460 : 4'b0000;
															assign node49460 = (inp[3]) ? 4'b0010 : 4'b0000;
														assign node49463 = (inp[5]) ? node49465 : 4'b0010;
															assign node49465 = (inp[3]) ? 4'b0000 : 4'b0010;
												assign node49468 = (inp[2]) ? node49484 : node49469;
													assign node49469 = (inp[5]) ? node49479 : node49470;
														assign node49470 = (inp[3]) ? 4'b0100 : node49471;
															assign node49471 = (inp[0]) ? node49475 : node49472;
																assign node49472 = (inp[15]) ? 4'b0100 : 4'b0110;
																assign node49475 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node49479 = (inp[0]) ? 4'b0110 : node49480;
															assign node49480 = (inp[15]) ? 4'b0110 : 4'b0100;
													assign node49484 = (inp[3]) ? 4'b0110 : 4'b0100;
											assign node49487 = (inp[4]) ? node49519 : node49488;
												assign node49488 = (inp[5]) ? node49512 : node49489;
													assign node49489 = (inp[2]) ? node49499 : node49490;
														assign node49490 = (inp[15]) ? node49492 : 4'b0100;
															assign node49492 = (inp[0]) ? node49496 : node49493;
																assign node49493 = (inp[3]) ? 4'b0110 : 4'b0100;
																assign node49496 = (inp[3]) ? 4'b0100 : 4'b0110;
														assign node49499 = (inp[3]) ? node49505 : node49500;
															assign node49500 = (inp[15]) ? node49502 : 4'b0110;
																assign node49502 = (inp[0]) ? 4'b0110 : 4'b0100;
															assign node49505 = (inp[0]) ? node49509 : node49506;
																assign node49506 = (inp[15]) ? 4'b0110 : 4'b0100;
																assign node49509 = (inp[15]) ? 4'b0100 : 4'b0110;
													assign node49512 = (inp[15]) ? node49516 : node49513;
														assign node49513 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node49516 = (inp[0]) ? 4'b0100 : 4'b0110;
												assign node49519 = (inp[15]) ? node49531 : node49520;
													assign node49520 = (inp[0]) ? node49526 : node49521;
														assign node49521 = (inp[3]) ? 4'b0000 : node49522;
															assign node49522 = (inp[5]) ? 4'b0000 : 4'b0010;
														assign node49526 = (inp[5]) ? 4'b0010 : node49527;
															assign node49527 = (inp[3]) ? 4'b0010 : 4'b0000;
													assign node49531 = (inp[0]) ? node49537 : node49532;
														assign node49532 = (inp[2]) ? node49534 : 4'b0010;
															assign node49534 = (inp[3]) ? 4'b0010 : 4'b0000;
														assign node49537 = (inp[5]) ? 4'b0000 : node49538;
															assign node49538 = (inp[3]) ? 4'b0000 : 4'b0010;
						assign node49542 = (inp[7]) ? node50588 : node49543;
							assign node49543 = (inp[8]) ? node50083 : node49544;
								assign node49544 = (inp[14]) ? node49854 : node49545;
									assign node49545 = (inp[2]) ? node49707 : node49546;
										assign node49546 = (inp[9]) ? node49622 : node49547;
											assign node49547 = (inp[12]) ? node49587 : node49548;
												assign node49548 = (inp[4]) ? node49564 : node49549;
													assign node49549 = (inp[5]) ? node49559 : node49550;
														assign node49550 = (inp[3]) ? 4'b0111 : node49551;
															assign node49551 = (inp[0]) ? node49555 : node49552;
																assign node49552 = (inp[15]) ? 4'b0101 : 4'b0111;
																assign node49555 = (inp[15]) ? 4'b0111 : 4'b0101;
														assign node49559 = (inp[3]) ? node49561 : 4'b0101;
															assign node49561 = (inp[15]) ? 4'b0101 : 4'b0111;
													assign node49564 = (inp[3]) ? node49574 : node49565;
														assign node49565 = (inp[5]) ? 4'b0011 : node49566;
															assign node49566 = (inp[0]) ? node49570 : node49567;
																assign node49567 = (inp[15]) ? 4'b0001 : 4'b0011;
																assign node49570 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node49574 = (inp[15]) ? node49580 : node49575;
															assign node49575 = (inp[0]) ? 4'b0001 : node49576;
																assign node49576 = (inp[5]) ? 4'b0001 : 4'b0011;
															assign node49580 = (inp[0]) ? node49584 : node49581;
																assign node49581 = (inp[5]) ? 4'b0011 : 4'b0001;
																assign node49584 = (inp[5]) ? 4'b0001 : 4'b0011;
												assign node49587 = (inp[4]) ? node49605 : node49588;
													assign node49588 = (inp[15]) ? node49600 : node49589;
														assign node49589 = (inp[0]) ? node49595 : node49590;
															assign node49590 = (inp[3]) ? node49592 : 4'b0011;
																assign node49592 = (inp[5]) ? 4'b0001 : 4'b0011;
															assign node49595 = (inp[5]) ? node49597 : 4'b0001;
																assign node49597 = (inp[3]) ? 4'b0011 : 4'b0001;
														assign node49600 = (inp[0]) ? node49602 : 4'b0001;
															assign node49602 = (inp[5]) ? 4'b0001 : 4'b0011;
													assign node49605 = (inp[5]) ? node49615 : node49606;
														assign node49606 = (inp[3]) ? node49608 : 4'b0101;
															assign node49608 = (inp[0]) ? node49612 : node49609;
																assign node49609 = (inp[15]) ? 4'b0111 : 4'b0101;
																assign node49612 = (inp[15]) ? 4'b0101 : 4'b0111;
														assign node49615 = (inp[15]) ? node49619 : node49616;
															assign node49616 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node49619 = (inp[0]) ? 4'b0101 : 4'b0111;
											assign node49622 = (inp[3]) ? node49666 : node49623;
												assign node49623 = (inp[4]) ? node49647 : node49624;
													assign node49624 = (inp[12]) ? node49632 : node49625;
														assign node49625 = (inp[15]) ? node49629 : node49626;
															assign node49626 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node49629 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node49632 = (inp[0]) ? node49640 : node49633;
															assign node49633 = (inp[5]) ? node49637 : node49634;
																assign node49634 = (inp[15]) ? 4'b0101 : 4'b0111;
																assign node49637 = (inp[15]) ? 4'b0111 : 4'b0101;
															assign node49640 = (inp[5]) ? node49644 : node49641;
																assign node49641 = (inp[15]) ? 4'b0111 : 4'b0101;
																assign node49644 = (inp[15]) ? 4'b0101 : 4'b0111;
													assign node49647 = (inp[12]) ? node49651 : node49648;
														assign node49648 = (inp[0]) ? 4'b0101 : 4'b0111;
														assign node49651 = (inp[15]) ? node49659 : node49652;
															assign node49652 = (inp[5]) ? node49656 : node49653;
																assign node49653 = (inp[0]) ? 4'b0001 : 4'b0011;
																assign node49656 = (inp[0]) ? 4'b0011 : 4'b0001;
															assign node49659 = (inp[5]) ? node49663 : node49660;
																assign node49660 = (inp[0]) ? 4'b0011 : 4'b0001;
																assign node49663 = (inp[0]) ? 4'b0001 : 4'b0011;
												assign node49666 = (inp[0]) ? node49684 : node49667;
													assign node49667 = (inp[15]) ? node49673 : node49668;
														assign node49668 = (inp[5]) ? node49670 : 4'b0101;
															assign node49670 = (inp[12]) ? 4'b0001 : 4'b0101;
														assign node49673 = (inp[5]) ? node49679 : node49674;
															assign node49674 = (inp[12]) ? node49676 : 4'b0111;
																assign node49676 = (inp[4]) ? 4'b0011 : 4'b0111;
															assign node49679 = (inp[12]) ? 4'b0111 : node49680;
																assign node49680 = (inp[4]) ? 4'b0111 : 4'b0011;
													assign node49684 = (inp[15]) ? node49700 : node49685;
														assign node49685 = (inp[5]) ? node49693 : node49686;
															assign node49686 = (inp[12]) ? node49690 : node49687;
																assign node49687 = (inp[4]) ? 4'b0111 : 4'b0001;
																assign node49690 = (inp[4]) ? 4'b0011 : 4'b0111;
															assign node49693 = (inp[12]) ? node49697 : node49694;
																assign node49694 = (inp[4]) ? 4'b0111 : 4'b0011;
																assign node49697 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node49700 = (inp[12]) ? 4'b0101 : node49701;
															assign node49701 = (inp[4]) ? 4'b0101 : node49702;
																assign node49702 = (inp[5]) ? 4'b0001 : 4'b0011;
										assign node49707 = (inp[5]) ? node49783 : node49708;
											assign node49708 = (inp[12]) ? node49738 : node49709;
												assign node49709 = (inp[15]) ? node49723 : node49710;
													assign node49710 = (inp[0]) ? node49718 : node49711;
														assign node49711 = (inp[3]) ? node49713 : 4'b0010;
															assign node49713 = (inp[9]) ? 4'b0100 : node49714;
																assign node49714 = (inp[4]) ? 4'b0010 : 4'b0110;
														assign node49718 = (inp[4]) ? 4'b0000 : node49719;
															assign node49719 = (inp[9]) ? 4'b0000 : 4'b0100;
													assign node49723 = (inp[0]) ? node49733 : node49724;
														assign node49724 = (inp[3]) ? 4'b0000 : node49725;
															assign node49725 = (inp[9]) ? node49729 : node49726;
																assign node49726 = (inp[4]) ? 4'b0000 : 4'b0100;
																assign node49729 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node49733 = (inp[4]) ? node49735 : 4'b0010;
															assign node49735 = (inp[9]) ? 4'b0100 : 4'b0010;
												assign node49738 = (inp[3]) ? node49768 : node49739;
													assign node49739 = (inp[0]) ? node49755 : node49740;
														assign node49740 = (inp[15]) ? node49748 : node49741;
															assign node49741 = (inp[9]) ? node49745 : node49742;
																assign node49742 = (inp[4]) ? 4'b0110 : 4'b0010;
																assign node49745 = (inp[4]) ? 4'b0010 : 4'b0110;
															assign node49748 = (inp[4]) ? node49752 : node49749;
																assign node49749 = (inp[9]) ? 4'b0100 : 4'b0000;
																assign node49752 = (inp[9]) ? 4'b0000 : 4'b0100;
														assign node49755 = (inp[15]) ? node49763 : node49756;
															assign node49756 = (inp[4]) ? node49760 : node49757;
																assign node49757 = (inp[9]) ? 4'b0100 : 4'b0000;
																assign node49760 = (inp[9]) ? 4'b0000 : 4'b0100;
															assign node49763 = (inp[4]) ? node49765 : 4'b0010;
																assign node49765 = (inp[9]) ? 4'b0010 : 4'b0110;
													assign node49768 = (inp[0]) ? node49774 : node49769;
														assign node49769 = (inp[15]) ? node49771 : 4'b0100;
															assign node49771 = (inp[4]) ? 4'b0010 : 4'b0110;
														assign node49774 = (inp[15]) ? node49778 : node49775;
															assign node49775 = (inp[4]) ? 4'b0110 : 4'b0000;
															assign node49778 = (inp[4]) ? node49780 : 4'b0100;
																assign node49780 = (inp[9]) ? 4'b0000 : 4'b0100;
											assign node49783 = (inp[4]) ? node49817 : node49784;
												assign node49784 = (inp[12]) ? node49802 : node49785;
													assign node49785 = (inp[9]) ? node49793 : node49786;
														assign node49786 = (inp[3]) ? node49788 : 4'b0100;
															assign node49788 = (inp[0]) ? node49790 : 4'b0110;
																assign node49790 = (inp[15]) ? 4'b0100 : 4'b0110;
														assign node49793 = (inp[0]) ? node49795 : 4'b0000;
															assign node49795 = (inp[3]) ? node49799 : node49796;
																assign node49796 = (inp[15]) ? 4'b0010 : 4'b0000;
																assign node49799 = (inp[15]) ? 4'b0000 : 4'b0010;
													assign node49802 = (inp[9]) ? node49810 : node49803;
														assign node49803 = (inp[3]) ? node49805 : 4'b0010;
															assign node49805 = (inp[15]) ? node49807 : 4'b0000;
																assign node49807 = (inp[0]) ? 4'b0000 : 4'b0010;
														assign node49810 = (inp[0]) ? node49814 : node49811;
															assign node49811 = (inp[15]) ? 4'b0110 : 4'b0100;
															assign node49814 = (inp[15]) ? 4'b0100 : 4'b0110;
												assign node49817 = (inp[15]) ? node49841 : node49818;
													assign node49818 = (inp[0]) ? node49828 : node49819;
														assign node49819 = (inp[9]) ? node49825 : node49820;
															assign node49820 = (inp[12]) ? 4'b0100 : node49821;
																assign node49821 = (inp[3]) ? 4'b0000 : 4'b0010;
															assign node49825 = (inp[12]) ? 4'b0000 : 4'b0100;
														assign node49828 = (inp[3]) ? node49834 : node49829;
															assign node49829 = (inp[12]) ? 4'b0110 : node49830;
																assign node49830 = (inp[9]) ? 4'b0110 : 4'b0000;
															assign node49834 = (inp[9]) ? node49838 : node49835;
																assign node49835 = (inp[12]) ? 4'b0110 : 4'b0010;
																assign node49838 = (inp[12]) ? 4'b0010 : 4'b0110;
													assign node49841 = (inp[0]) ? node49849 : node49842;
														assign node49842 = (inp[9]) ? node49846 : node49843;
															assign node49843 = (inp[12]) ? 4'b0110 : 4'b0010;
															assign node49846 = (inp[12]) ? 4'b0010 : 4'b0110;
														assign node49849 = (inp[12]) ? node49851 : 4'b0010;
															assign node49851 = (inp[9]) ? 4'b0000 : 4'b0100;
									assign node49854 = (inp[9]) ? node49976 : node49855;
										assign node49855 = (inp[15]) ? node49921 : node49856;
											assign node49856 = (inp[0]) ? node49884 : node49857;
												assign node49857 = (inp[5]) ? node49871 : node49858;
													assign node49858 = (inp[2]) ? node49864 : node49859;
														assign node49859 = (inp[4]) ? node49861 : 4'b0010;
															assign node49861 = (inp[3]) ? 4'b0100 : 4'b0110;
														assign node49864 = (inp[4]) ? node49868 : node49865;
															assign node49865 = (inp[12]) ? 4'b0010 : 4'b0110;
															assign node49868 = (inp[12]) ? 4'b0110 : 4'b0010;
													assign node49871 = (inp[3]) ? node49877 : node49872;
														assign node49872 = (inp[2]) ? node49874 : 4'b0010;
															assign node49874 = (inp[4]) ? 4'b0100 : 4'b0010;
														assign node49877 = (inp[4]) ? node49881 : node49878;
															assign node49878 = (inp[12]) ? 4'b0000 : 4'b0100;
															assign node49881 = (inp[12]) ? 4'b0100 : 4'b0000;
												assign node49884 = (inp[3]) ? node49902 : node49885;
													assign node49885 = (inp[2]) ? node49893 : node49886;
														assign node49886 = (inp[5]) ? 4'b0000 : node49887;
															assign node49887 = (inp[12]) ? 4'b0000 : node49888;
																assign node49888 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node49893 = (inp[4]) ? node49897 : node49894;
															assign node49894 = (inp[12]) ? 4'b0000 : 4'b0100;
															assign node49897 = (inp[12]) ? node49899 : 4'b0000;
																assign node49899 = (inp[5]) ? 4'b0110 : 4'b0100;
													assign node49902 = (inp[5]) ? node49910 : node49903;
														assign node49903 = (inp[4]) ? node49907 : node49904;
															assign node49904 = (inp[12]) ? 4'b0000 : 4'b0100;
															assign node49907 = (inp[12]) ? 4'b0110 : 4'b0000;
														assign node49910 = (inp[2]) ? node49916 : node49911;
															assign node49911 = (inp[4]) ? 4'b0010 : node49912;
																assign node49912 = (inp[12]) ? 4'b0010 : 4'b0110;
															assign node49916 = (inp[4]) ? node49918 : 4'b0110;
																assign node49918 = (inp[12]) ? 4'b0110 : 4'b0010;
											assign node49921 = (inp[0]) ? node49949 : node49922;
												assign node49922 = (inp[5]) ? node49932 : node49923;
													assign node49923 = (inp[12]) ? node49927 : node49924;
														assign node49924 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node49927 = (inp[4]) ? node49929 : 4'b0000;
															assign node49929 = (inp[3]) ? 4'b0110 : 4'b0100;
													assign node49932 = (inp[3]) ? node49942 : node49933;
														assign node49933 = (inp[2]) ? node49939 : node49934;
															assign node49934 = (inp[12]) ? node49936 : 4'b0000;
																assign node49936 = (inp[4]) ? 4'b0110 : 4'b0000;
															assign node49939 = (inp[12]) ? 4'b0110 : 4'b0100;
														assign node49942 = (inp[4]) ? node49946 : node49943;
															assign node49943 = (inp[12]) ? 4'b0010 : 4'b0110;
															assign node49946 = (inp[12]) ? 4'b0110 : 4'b0010;
												assign node49949 = (inp[3]) ? node49957 : node49950;
													assign node49950 = (inp[2]) ? 4'b0110 : node49951;
														assign node49951 = (inp[12]) ? 4'b0010 : node49952;
															assign node49952 = (inp[4]) ? 4'b0010 : 4'b0110;
													assign node49957 = (inp[5]) ? node49965 : node49958;
														assign node49958 = (inp[12]) ? node49962 : node49959;
															assign node49959 = (inp[4]) ? 4'b0010 : 4'b0110;
															assign node49962 = (inp[4]) ? 4'b0100 : 4'b0010;
														assign node49965 = (inp[2]) ? node49971 : node49966;
															assign node49966 = (inp[12]) ? node49968 : 4'b0100;
																assign node49968 = (inp[4]) ? 4'b0100 : 4'b0000;
															assign node49971 = (inp[12]) ? 4'b0000 : node49972;
																assign node49972 = (inp[4]) ? 4'b0000 : 4'b0100;
										assign node49976 = (inp[0]) ? node50030 : node49977;
											assign node49977 = (inp[15]) ? node50001 : node49978;
												assign node49978 = (inp[5]) ? node49994 : node49979;
													assign node49979 = (inp[3]) ? node49987 : node49980;
														assign node49980 = (inp[4]) ? node49984 : node49981;
															assign node49981 = (inp[12]) ? 4'b0110 : 4'b0010;
															assign node49984 = (inp[12]) ? 4'b0010 : 4'b0110;
														assign node49987 = (inp[4]) ? node49991 : node49988;
															assign node49988 = (inp[12]) ? 4'b0100 : 4'b0010;
															assign node49991 = (inp[12]) ? 4'b0000 : 4'b0100;
													assign node49994 = (inp[12]) ? node49998 : node49995;
														assign node49995 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node49998 = (inp[4]) ? 4'b0000 : 4'b0100;
												assign node50001 = (inp[3]) ? node50021 : node50002;
													assign node50002 = (inp[5]) ? node50016 : node50003;
														assign node50003 = (inp[2]) ? node50011 : node50004;
															assign node50004 = (inp[4]) ? node50008 : node50005;
																assign node50005 = (inp[12]) ? 4'b0100 : 4'b0000;
																assign node50008 = (inp[12]) ? 4'b0000 : 4'b0100;
															assign node50011 = (inp[12]) ? 4'b0100 : node50012;
																assign node50012 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node50016 = (inp[12]) ? node50018 : 4'b0000;
															assign node50018 = (inp[4]) ? 4'b0010 : 4'b0110;
													assign node50021 = (inp[12]) ? node50027 : node50022;
														assign node50022 = (inp[4]) ? 4'b0110 : node50023;
															assign node50023 = (inp[5]) ? 4'b0010 : 4'b0000;
														assign node50027 = (inp[4]) ? 4'b0010 : 4'b0110;
											assign node50030 = (inp[15]) ? node50056 : node50031;
												assign node50031 = (inp[5]) ? node50049 : node50032;
													assign node50032 = (inp[3]) ? node50040 : node50033;
														assign node50033 = (inp[4]) ? node50037 : node50034;
															assign node50034 = (inp[12]) ? 4'b0100 : 4'b0000;
															assign node50037 = (inp[12]) ? 4'b0000 : 4'b0100;
														assign node50040 = (inp[2]) ? node50046 : node50041;
															assign node50041 = (inp[4]) ? node50043 : 4'b0110;
																assign node50043 = (inp[12]) ? 4'b0010 : 4'b0110;
															assign node50046 = (inp[4]) ? 4'b0010 : 4'b0000;
													assign node50049 = (inp[12]) ? node50053 : node50050;
														assign node50050 = (inp[4]) ? 4'b0110 : 4'b0010;
														assign node50053 = (inp[4]) ? 4'b0010 : 4'b0110;
												assign node50056 = (inp[5]) ? node50074 : node50057;
													assign node50057 = (inp[3]) ? node50067 : node50058;
														assign node50058 = (inp[2]) ? 4'b0010 : node50059;
															assign node50059 = (inp[4]) ? node50063 : node50060;
																assign node50060 = (inp[12]) ? 4'b0110 : 4'b0010;
																assign node50063 = (inp[12]) ? 4'b0010 : 4'b0110;
														assign node50067 = (inp[4]) ? node50071 : node50068;
															assign node50068 = (inp[12]) ? 4'b0100 : 4'b0010;
															assign node50071 = (inp[12]) ? 4'b0000 : 4'b0100;
													assign node50074 = (inp[12]) ? node50080 : node50075;
														assign node50075 = (inp[2]) ? 4'b0100 : node50076;
															assign node50076 = (inp[3]) ? 4'b0000 : 4'b0010;
														assign node50080 = (inp[4]) ? 4'b0000 : 4'b0100;
								assign node50083 = (inp[2]) ? node50373 : node50084;
									assign node50084 = (inp[14]) ? node50242 : node50085;
										assign node50085 = (inp[5]) ? node50171 : node50086;
											assign node50086 = (inp[3]) ? node50136 : node50087;
												assign node50087 = (inp[9]) ? node50111 : node50088;
													assign node50088 = (inp[0]) ? node50098 : node50089;
														assign node50089 = (inp[15]) ? node50091 : 4'b0010;
															assign node50091 = (inp[12]) ? node50095 : node50092;
																assign node50092 = (inp[4]) ? 4'b0000 : 4'b0100;
																assign node50095 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node50098 = (inp[15]) ? node50106 : node50099;
															assign node50099 = (inp[4]) ? node50103 : node50100;
																assign node50100 = (inp[12]) ? 4'b0000 : 4'b0100;
																assign node50103 = (inp[12]) ? 4'b0100 : 4'b0000;
															assign node50106 = (inp[4]) ? 4'b0010 : node50107;
																assign node50107 = (inp[12]) ? 4'b0010 : 4'b0110;
													assign node50111 = (inp[12]) ? node50123 : node50112;
														assign node50112 = (inp[4]) ? node50118 : node50113;
															assign node50113 = (inp[15]) ? 4'b0000 : node50114;
																assign node50114 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node50118 = (inp[0]) ? 4'b0100 : node50119;
																assign node50119 = (inp[15]) ? 4'b0100 : 4'b0110;
														assign node50123 = (inp[4]) ? node50131 : node50124;
															assign node50124 = (inp[0]) ? node50128 : node50125;
																assign node50125 = (inp[15]) ? 4'b0100 : 4'b0110;
																assign node50128 = (inp[15]) ? 4'b0110 : 4'b0100;
															assign node50131 = (inp[15]) ? node50133 : 4'b0000;
																assign node50133 = (inp[0]) ? 4'b0010 : 4'b0000;
												assign node50136 = (inp[12]) ? node50154 : node50137;
													assign node50137 = (inp[15]) ? node50151 : node50138;
														assign node50138 = (inp[0]) ? node50146 : node50139;
															assign node50139 = (inp[9]) ? node50143 : node50140;
																assign node50140 = (inp[4]) ? 4'b0010 : 4'b0110;
																assign node50143 = (inp[4]) ? 4'b0100 : 4'b0010;
															assign node50146 = (inp[9]) ? 4'b0000 : node50147;
																assign node50147 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node50151 = (inp[0]) ? 4'b0010 : 4'b0000;
													assign node50154 = (inp[4]) ? node50160 : node50155;
														assign node50155 = (inp[9]) ? node50157 : 4'b0000;
															assign node50157 = (inp[0]) ? 4'b0100 : 4'b0110;
														assign node50160 = (inp[9]) ? node50166 : node50161;
															assign node50161 = (inp[15]) ? 4'b0110 : node50162;
																assign node50162 = (inp[0]) ? 4'b0110 : 4'b0100;
															assign node50166 = (inp[15]) ? 4'b0010 : node50167;
																assign node50167 = (inp[0]) ? 4'b0010 : 4'b0000;
											assign node50171 = (inp[15]) ? node50207 : node50172;
												assign node50172 = (inp[0]) ? node50190 : node50173;
													assign node50173 = (inp[3]) ? node50183 : node50174;
														assign node50174 = (inp[12]) ? 4'b0100 : node50175;
															assign node50175 = (inp[4]) ? node50179 : node50176;
																assign node50176 = (inp[9]) ? 4'b0010 : 4'b0110;
																assign node50179 = (inp[9]) ? 4'b0100 : 4'b0010;
														assign node50183 = (inp[4]) ? node50185 : 4'b0100;
															assign node50185 = (inp[12]) ? 4'b0000 : node50186;
																assign node50186 = (inp[9]) ? 4'b0100 : 4'b0000;
													assign node50190 = (inp[3]) ? node50198 : node50191;
														assign node50191 = (inp[4]) ? node50193 : 4'b0100;
															assign node50193 = (inp[12]) ? node50195 : 4'b0110;
																assign node50195 = (inp[9]) ? 4'b0010 : 4'b0110;
														assign node50198 = (inp[12]) ? 4'b0110 : node50199;
															assign node50199 = (inp[4]) ? node50203 : node50200;
																assign node50200 = (inp[9]) ? 4'b0010 : 4'b0110;
																assign node50203 = (inp[9]) ? 4'b0110 : 4'b0010;
												assign node50207 = (inp[0]) ? node50227 : node50208;
													assign node50208 = (inp[3]) ? node50218 : node50209;
														assign node50209 = (inp[9]) ? node50215 : node50210;
															assign node50210 = (inp[12]) ? 4'b0000 : node50211;
																assign node50211 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node50215 = (inp[4]) ? 4'b0010 : 4'b0110;
														assign node50218 = (inp[4]) ? node50220 : 4'b0110;
															assign node50220 = (inp[12]) ? node50224 : node50221;
																assign node50221 = (inp[9]) ? 4'b0110 : 4'b0010;
																assign node50224 = (inp[9]) ? 4'b0010 : 4'b0110;
													assign node50227 = (inp[3]) ? node50235 : node50228;
														assign node50228 = (inp[4]) ? node50230 : 4'b0010;
															assign node50230 = (inp[9]) ? node50232 : 4'b0010;
																assign node50232 = (inp[12]) ? 4'b0000 : 4'b0100;
														assign node50235 = (inp[9]) ? 4'b0000 : node50236;
															assign node50236 = (inp[12]) ? node50238 : 4'b0100;
																assign node50238 = (inp[4]) ? 4'b0100 : 4'b0000;
										assign node50242 = (inp[5]) ? node50306 : node50243;
											assign node50243 = (inp[9]) ? node50269 : node50244;
												assign node50244 = (inp[4]) ? node50254 : node50245;
													assign node50245 = (inp[12]) ? node50247 : 4'b1011;
														assign node50247 = (inp[0]) ? node50251 : node50248;
															assign node50248 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node50251 = (inp[15]) ? 4'b1011 : 4'b1001;
													assign node50254 = (inp[3]) ? node50262 : node50255;
														assign node50255 = (inp[0]) ? node50259 : node50256;
															assign node50256 = (inp[15]) ? 4'b1101 : 4'b1111;
															assign node50259 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node50262 = (inp[12]) ? 4'b1111 : node50263;
															assign node50263 = (inp[15]) ? node50265 : 4'b1111;
																assign node50265 = (inp[0]) ? 4'b1101 : 4'b1111;
												assign node50269 = (inp[4]) ? node50285 : node50270;
													assign node50270 = (inp[15]) ? node50278 : node50271;
														assign node50271 = (inp[0]) ? node50275 : node50272;
															assign node50272 = (inp[3]) ? 4'b1101 : 4'b1111;
															assign node50275 = (inp[3]) ? 4'b1111 : 4'b1101;
														assign node50278 = (inp[0]) ? node50282 : node50279;
															assign node50279 = (inp[3]) ? 4'b1111 : 4'b1101;
															assign node50282 = (inp[3]) ? 4'b1101 : 4'b1111;
													assign node50285 = (inp[15]) ? node50301 : node50286;
														assign node50286 = (inp[12]) ? node50294 : node50287;
															assign node50287 = (inp[3]) ? node50291 : node50288;
																assign node50288 = (inp[0]) ? 4'b1001 : 4'b1011;
																assign node50291 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node50294 = (inp[0]) ? node50298 : node50295;
																assign node50295 = (inp[3]) ? 4'b1001 : 4'b1011;
																assign node50298 = (inp[3]) ? 4'b1011 : 4'b1001;
														assign node50301 = (inp[3]) ? 4'b1001 : node50302;
															assign node50302 = (inp[0]) ? 4'b1011 : 4'b1001;
											assign node50306 = (inp[3]) ? node50344 : node50307;
												assign node50307 = (inp[12]) ? node50329 : node50308;
													assign node50308 = (inp[15]) ? node50320 : node50309;
														assign node50309 = (inp[0]) ? node50317 : node50310;
															assign node50310 = (inp[9]) ? node50314 : node50311;
																assign node50311 = (inp[4]) ? 4'b1101 : 4'b1011;
																assign node50314 = (inp[4]) ? 4'b1001 : 4'b1101;
															assign node50317 = (inp[9]) ? 4'b1011 : 4'b1001;
														assign node50320 = (inp[0]) ? node50324 : node50321;
															assign node50321 = (inp[9]) ? 4'b1011 : 4'b1001;
															assign node50324 = (inp[4]) ? node50326 : 4'b1011;
																assign node50326 = (inp[9]) ? 4'b1001 : 4'b1101;
													assign node50329 = (inp[15]) ? node50333 : node50330;
														assign node50330 = (inp[9]) ? 4'b1111 : 4'b1011;
														assign node50333 = (inp[9]) ? node50341 : node50334;
															assign node50334 = (inp[4]) ? node50338 : node50335;
																assign node50335 = (inp[0]) ? 4'b1011 : 4'b1001;
																assign node50338 = (inp[0]) ? 4'b1101 : 4'b1111;
															assign node50341 = (inp[0]) ? 4'b1001 : 4'b1011;
												assign node50344 = (inp[9]) ? node50358 : node50345;
													assign node50345 = (inp[4]) ? node50349 : node50346;
														assign node50346 = (inp[15]) ? 4'b1001 : 4'b1011;
														assign node50349 = (inp[12]) ? node50351 : 4'b1101;
															assign node50351 = (inp[15]) ? node50355 : node50352;
																assign node50352 = (inp[0]) ? 4'b1111 : 4'b1101;
																assign node50355 = (inp[0]) ? 4'b1101 : 4'b1111;
													assign node50358 = (inp[4]) ? node50364 : node50359;
														assign node50359 = (inp[12]) ? 4'b1101 : node50360;
															assign node50360 = (inp[0]) ? 4'b1101 : 4'b1111;
														assign node50364 = (inp[12]) ? node50366 : 4'b1011;
															assign node50366 = (inp[15]) ? node50370 : node50367;
																assign node50367 = (inp[0]) ? 4'b1011 : 4'b1001;
																assign node50370 = (inp[0]) ? 4'b1001 : 4'b1011;
									assign node50373 = (inp[14]) ? node50487 : node50374;
										assign node50374 = (inp[15]) ? node50438 : node50375;
											assign node50375 = (inp[0]) ? node50407 : node50376;
												assign node50376 = (inp[3]) ? node50394 : node50377;
													assign node50377 = (inp[5]) ? node50389 : node50378;
														assign node50378 = (inp[12]) ? node50384 : node50379;
															assign node50379 = (inp[4]) ? 4'b1111 : node50380;
																assign node50380 = (inp[9]) ? 4'b1111 : 4'b1011;
															assign node50384 = (inp[4]) ? 4'b1011 : node50385;
																assign node50385 = (inp[9]) ? 4'b1111 : 4'b1011;
														assign node50389 = (inp[4]) ? node50391 : 4'b1011;
															assign node50391 = (inp[9]) ? 4'b1001 : 4'b1101;
													assign node50394 = (inp[5]) ? node50400 : node50395;
														assign node50395 = (inp[4]) ? node50397 : 4'b1101;
															assign node50397 = (inp[9]) ? 4'b1001 : 4'b1101;
														assign node50400 = (inp[9]) ? node50404 : node50401;
															assign node50401 = (inp[4]) ? 4'b1101 : 4'b1001;
															assign node50404 = (inp[4]) ? 4'b1001 : 4'b1101;
												assign node50407 = (inp[3]) ? node50423 : node50408;
													assign node50408 = (inp[5]) ? node50416 : node50409;
														assign node50409 = (inp[4]) ? node50413 : node50410;
															assign node50410 = (inp[9]) ? 4'b1101 : 4'b1001;
															assign node50413 = (inp[9]) ? 4'b1001 : 4'b1101;
														assign node50416 = (inp[12]) ? 4'b1111 : node50417;
															assign node50417 = (inp[9]) ? 4'b1111 : node50418;
																assign node50418 = (inp[4]) ? 4'b1111 : 4'b1001;
													assign node50423 = (inp[5]) ? node50429 : node50424;
														assign node50424 = (inp[4]) ? node50426 : 4'b1111;
															assign node50426 = (inp[9]) ? 4'b1011 : 4'b1111;
														assign node50429 = (inp[12]) ? node50431 : 4'b1111;
															assign node50431 = (inp[4]) ? node50435 : node50432;
																assign node50432 = (inp[9]) ? 4'b1111 : 4'b1011;
																assign node50435 = (inp[9]) ? 4'b1011 : 4'b1111;
											assign node50438 = (inp[0]) ? node50460 : node50439;
												assign node50439 = (inp[5]) ? node50451 : node50440;
													assign node50440 = (inp[4]) ? node50444 : node50441;
														assign node50441 = (inp[9]) ? 4'b1101 : 4'b1001;
														assign node50444 = (inp[3]) ? node50448 : node50445;
															assign node50445 = (inp[9]) ? 4'b1001 : 4'b1101;
															assign node50448 = (inp[9]) ? 4'b1011 : 4'b1111;
													assign node50451 = (inp[9]) ? node50457 : node50452;
														assign node50452 = (inp[4]) ? 4'b1111 : node50453;
															assign node50453 = (inp[3]) ? 4'b1011 : 4'b1001;
														assign node50457 = (inp[4]) ? 4'b1011 : 4'b1111;
												assign node50460 = (inp[3]) ? node50478 : node50461;
													assign node50461 = (inp[5]) ? node50471 : node50462;
														assign node50462 = (inp[12]) ? node50468 : node50463;
															assign node50463 = (inp[4]) ? node50465 : 4'b1111;
																assign node50465 = (inp[9]) ? 4'b1011 : 4'b1111;
															assign node50468 = (inp[4]) ? 4'b1111 : 4'b1011;
														assign node50471 = (inp[4]) ? node50475 : node50472;
															assign node50472 = (inp[9]) ? 4'b1101 : 4'b1011;
															assign node50475 = (inp[9]) ? 4'b1001 : 4'b1101;
													assign node50478 = (inp[9]) ? node50484 : node50479;
														assign node50479 = (inp[4]) ? 4'b1101 : node50480;
															assign node50480 = (inp[5]) ? 4'b1001 : 4'b1011;
														assign node50484 = (inp[4]) ? 4'b1001 : 4'b1101;
										assign node50487 = (inp[9]) ? node50545 : node50488;
											assign node50488 = (inp[4]) ? node50520 : node50489;
												assign node50489 = (inp[12]) ? node50505 : node50490;
													assign node50490 = (inp[0]) ? node50496 : node50491;
														assign node50491 = (inp[5]) ? 4'b1001 : node50492;
															assign node50492 = (inp[15]) ? 4'b1001 : 4'b1011;
														assign node50496 = (inp[15]) ? node50502 : node50497;
															assign node50497 = (inp[5]) ? node50499 : 4'b1001;
																assign node50499 = (inp[3]) ? 4'b1011 : 4'b1001;
															assign node50502 = (inp[3]) ? 4'b1001 : 4'b1011;
													assign node50505 = (inp[5]) ? node50513 : node50506;
														assign node50506 = (inp[0]) ? node50510 : node50507;
															assign node50507 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node50510 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node50513 = (inp[3]) ? node50515 : 4'b1011;
															assign node50515 = (inp[0]) ? 4'b1011 : node50516;
																assign node50516 = (inp[15]) ? 4'b1011 : 4'b1001;
												assign node50520 = (inp[5]) ? node50542 : node50521;
													assign node50521 = (inp[3]) ? node50537 : node50522;
														assign node50522 = (inp[12]) ? node50530 : node50523;
															assign node50523 = (inp[15]) ? node50527 : node50524;
																assign node50524 = (inp[0]) ? 4'b1101 : 4'b1111;
																assign node50527 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node50530 = (inp[0]) ? node50534 : node50531;
																assign node50531 = (inp[15]) ? 4'b1101 : 4'b1111;
																assign node50534 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node50537 = (inp[0]) ? 4'b1111 : node50538;
															assign node50538 = (inp[15]) ? 4'b1111 : 4'b1101;
													assign node50542 = (inp[0]) ? 4'b1101 : 4'b1111;
											assign node50545 = (inp[4]) ? node50561 : node50546;
												assign node50546 = (inp[15]) ? node50554 : node50547;
													assign node50547 = (inp[0]) ? 4'b1111 : node50548;
														assign node50548 = (inp[5]) ? 4'b1101 : node50549;
															assign node50549 = (inp[12]) ? 4'b1111 : 4'b1101;
													assign node50554 = (inp[0]) ? node50556 : 4'b1111;
														assign node50556 = (inp[3]) ? 4'b1101 : node50557;
															assign node50557 = (inp[5]) ? 4'b1101 : 4'b1111;
												assign node50561 = (inp[5]) ? node50581 : node50562;
													assign node50562 = (inp[15]) ? node50570 : node50563;
														assign node50563 = (inp[12]) ? 4'b1011 : node50564;
															assign node50564 = (inp[3]) ? 4'b1001 : node50565;
																assign node50565 = (inp[0]) ? 4'b1001 : 4'b1011;
														assign node50570 = (inp[12]) ? node50576 : node50571;
															assign node50571 = (inp[3]) ? node50573 : 4'b1001;
																assign node50573 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node50576 = (inp[0]) ? node50578 : 4'b1001;
																assign node50578 = (inp[3]) ? 4'b1001 : 4'b1011;
													assign node50581 = (inp[3]) ? 4'b1011 : node50582;
														assign node50582 = (inp[0]) ? node50584 : 4'b1011;
															assign node50584 = (inp[15]) ? 4'b1001 : 4'b1011;
							assign node50588 = (inp[8]) ? node51018 : node50589;
								assign node50589 = (inp[2]) ? node50831 : node50590;
									assign node50590 = (inp[14]) ? node50732 : node50591;
										assign node50591 = (inp[0]) ? node50677 : node50592;
											assign node50592 = (inp[3]) ? node50642 : node50593;
												assign node50593 = (inp[15]) ? node50619 : node50594;
													assign node50594 = (inp[5]) ? node50610 : node50595;
														assign node50595 = (inp[4]) ? node50603 : node50596;
															assign node50596 = (inp[12]) ? node50600 : node50597;
																assign node50597 = (inp[9]) ? 4'b0010 : 4'b0110;
																assign node50600 = (inp[9]) ? 4'b0110 : 4'b0010;
															assign node50603 = (inp[12]) ? node50607 : node50604;
																assign node50604 = (inp[9]) ? 4'b0110 : 4'b0010;
																assign node50607 = (inp[9]) ? 4'b0010 : 4'b0110;
														assign node50610 = (inp[4]) ? 4'b0100 : node50611;
															assign node50611 = (inp[12]) ? node50615 : node50612;
																assign node50612 = (inp[9]) ? 4'b0010 : 4'b0110;
																assign node50615 = (inp[9]) ? 4'b0100 : 4'b0010;
													assign node50619 = (inp[5]) ? node50631 : node50620;
														assign node50620 = (inp[4]) ? node50626 : node50621;
															assign node50621 = (inp[12]) ? node50623 : 4'b0100;
																assign node50623 = (inp[9]) ? 4'b0100 : 4'b0000;
															assign node50626 = (inp[9]) ? 4'b0000 : node50627;
																assign node50627 = (inp[12]) ? 4'b0100 : 4'b0000;
														assign node50631 = (inp[9]) ? node50637 : node50632;
															assign node50632 = (inp[12]) ? 4'b0110 : node50633;
																assign node50633 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node50637 = (inp[4]) ? node50639 : 4'b0110;
																assign node50639 = (inp[12]) ? 4'b0010 : 4'b0110;
												assign node50642 = (inp[15]) ? node50652 : node50643;
													assign node50643 = (inp[4]) ? node50645 : 4'b0000;
														assign node50645 = (inp[9]) ? node50649 : node50646;
															assign node50646 = (inp[12]) ? 4'b0100 : 4'b0010;
															assign node50649 = (inp[12]) ? 4'b0000 : 4'b0100;
													assign node50652 = (inp[5]) ? node50662 : node50653;
														assign node50653 = (inp[4]) ? node50659 : node50654;
															assign node50654 = (inp[9]) ? 4'b0000 : node50655;
																assign node50655 = (inp[12]) ? 4'b0000 : 4'b0100;
															assign node50659 = (inp[9]) ? 4'b0010 : 4'b0110;
														assign node50662 = (inp[12]) ? node50670 : node50663;
															assign node50663 = (inp[9]) ? node50667 : node50664;
																assign node50664 = (inp[4]) ? 4'b0010 : 4'b0110;
																assign node50667 = (inp[4]) ? 4'b0110 : 4'b0010;
															assign node50670 = (inp[4]) ? node50674 : node50671;
																assign node50671 = (inp[9]) ? 4'b0110 : 4'b0010;
																assign node50674 = (inp[9]) ? 4'b0010 : 4'b0110;
											assign node50677 = (inp[12]) ? node50717 : node50678;
												assign node50678 = (inp[15]) ? node50698 : node50679;
													assign node50679 = (inp[3]) ? node50683 : node50680;
														assign node50680 = (inp[9]) ? 4'b0000 : 4'b0100;
														assign node50683 = (inp[5]) ? node50691 : node50684;
															assign node50684 = (inp[9]) ? node50688 : node50685;
																assign node50685 = (inp[4]) ? 4'b0000 : 4'b0100;
																assign node50688 = (inp[4]) ? 4'b0110 : 4'b0000;
															assign node50691 = (inp[9]) ? node50695 : node50692;
																assign node50692 = (inp[4]) ? 4'b0010 : 4'b0110;
																assign node50695 = (inp[4]) ? 4'b0110 : 4'b0010;
													assign node50698 = (inp[3]) ? node50706 : node50699;
														assign node50699 = (inp[5]) ? 4'b0010 : node50700;
															assign node50700 = (inp[9]) ? 4'b0110 : node50701;
																assign node50701 = (inp[4]) ? 4'b0010 : 4'b0110;
														assign node50706 = (inp[5]) ? node50712 : node50707;
															assign node50707 = (inp[9]) ? node50709 : 4'b0010;
																assign node50709 = (inp[4]) ? 4'b0100 : 4'b0010;
															assign node50712 = (inp[4]) ? node50714 : 4'b0000;
																assign node50714 = (inp[9]) ? 4'b0100 : 4'b0000;
												assign node50717 = (inp[4]) ? node50725 : node50718;
													assign node50718 = (inp[9]) ? node50722 : node50719;
														assign node50719 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node50722 = (inp[5]) ? 4'b0100 : 4'b0110;
													assign node50725 = (inp[9]) ? 4'b0000 : node50726;
														assign node50726 = (inp[15]) ? 4'b0100 : node50727;
															assign node50727 = (inp[3]) ? 4'b0110 : 4'b0100;
										assign node50732 = (inp[9]) ? node50796 : node50733;
											assign node50733 = (inp[4]) ? node50767 : node50734;
												assign node50734 = (inp[3]) ? node50754 : node50735;
													assign node50735 = (inp[5]) ? node50743 : node50736;
														assign node50736 = (inp[0]) ? node50740 : node50737;
															assign node50737 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node50740 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node50743 = (inp[12]) ? node50749 : node50744;
															assign node50744 = (inp[15]) ? node50746 : 4'b1001;
																assign node50746 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node50749 = (inp[15]) ? 4'b1001 : node50750;
																assign node50750 = (inp[0]) ? 4'b1001 : 4'b1011;
													assign node50754 = (inp[0]) ? node50762 : node50755;
														assign node50755 = (inp[12]) ? node50757 : 4'b1011;
															assign node50757 = (inp[5]) ? node50759 : 4'b1011;
																assign node50759 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node50762 = (inp[15]) ? 4'b1001 : node50763;
															assign node50763 = (inp[5]) ? 4'b1011 : 4'b1001;
												assign node50767 = (inp[3]) ? node50789 : node50768;
													assign node50768 = (inp[5]) ? node50782 : node50769;
														assign node50769 = (inp[12]) ? node50777 : node50770;
															assign node50770 = (inp[15]) ? node50774 : node50771;
																assign node50771 = (inp[0]) ? 4'b1101 : 4'b1111;
																assign node50774 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node50777 = (inp[0]) ? 4'b1111 : node50778;
																assign node50778 = (inp[15]) ? 4'b1101 : 4'b1111;
														assign node50782 = (inp[15]) ? node50786 : node50783;
															assign node50783 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node50786 = (inp[0]) ? 4'b1101 : 4'b1111;
													assign node50789 = (inp[0]) ? node50793 : node50790;
														assign node50790 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node50793 = (inp[15]) ? 4'b1101 : 4'b1111;
											assign node50796 = (inp[4]) ? node50816 : node50797;
												assign node50797 = (inp[5]) ? node50811 : node50798;
													assign node50798 = (inp[12]) ? node50806 : node50799;
														assign node50799 = (inp[3]) ? node50801 : 4'b1101;
															assign node50801 = (inp[0]) ? 4'b1111 : node50802;
																assign node50802 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node50806 = (inp[3]) ? node50808 : 4'b1111;
															assign node50808 = (inp[0]) ? 4'b1101 : 4'b1111;
													assign node50811 = (inp[15]) ? 4'b1111 : node50812;
														assign node50812 = (inp[0]) ? 4'b1111 : 4'b1101;
												assign node50816 = (inp[0]) ? node50822 : node50817;
													assign node50817 = (inp[15]) ? node50819 : 4'b1001;
														assign node50819 = (inp[3]) ? 4'b1011 : 4'b1001;
													assign node50822 = (inp[5]) ? 4'b1011 : node50823;
														assign node50823 = (inp[12]) ? node50825 : 4'b1011;
															assign node50825 = (inp[3]) ? 4'b1011 : node50826;
																assign node50826 = (inp[15]) ? 4'b1011 : 4'b1001;
									assign node50831 = (inp[5]) ? node50931 : node50832;
										assign node50832 = (inp[9]) ? node50864 : node50833;
											assign node50833 = (inp[4]) ? node50841 : node50834;
												assign node50834 = (inp[15]) ? node50838 : node50835;
													assign node50835 = (inp[0]) ? 4'b1001 : 4'b1011;
													assign node50838 = (inp[0]) ? 4'b1011 : 4'b1001;
												assign node50841 = (inp[3]) ? node50857 : node50842;
													assign node50842 = (inp[12]) ? node50850 : node50843;
														assign node50843 = (inp[14]) ? 4'b1111 : node50844;
															assign node50844 = (inp[0]) ? node50846 : 4'b1111;
																assign node50846 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node50850 = (inp[14]) ? node50852 : 4'b1111;
															assign node50852 = (inp[15]) ? node50854 : 4'b1101;
																assign node50854 = (inp[0]) ? 4'b1111 : 4'b1101;
													assign node50857 = (inp[15]) ? node50861 : node50858;
														assign node50858 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node50861 = (inp[0]) ? 4'b1101 : 4'b1111;
											assign node50864 = (inp[4]) ? node50898 : node50865;
												assign node50865 = (inp[14]) ? node50883 : node50866;
													assign node50866 = (inp[0]) ? node50876 : node50867;
														assign node50867 = (inp[12]) ? 4'b1111 : node50868;
															assign node50868 = (inp[15]) ? node50872 : node50869;
																assign node50869 = (inp[3]) ? 4'b1101 : 4'b1111;
																assign node50872 = (inp[3]) ? 4'b1111 : 4'b1101;
														assign node50876 = (inp[3]) ? node50880 : node50877;
															assign node50877 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node50880 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node50883 = (inp[0]) ? node50891 : node50884;
														assign node50884 = (inp[3]) ? node50888 : node50885;
															assign node50885 = (inp[15]) ? 4'b1101 : 4'b1111;
															assign node50888 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node50891 = (inp[3]) ? node50895 : node50892;
															assign node50892 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node50895 = (inp[15]) ? 4'b1101 : 4'b1111;
												assign node50898 = (inp[12]) ? node50912 : node50899;
													assign node50899 = (inp[14]) ? node50905 : node50900;
														assign node50900 = (inp[3]) ? node50902 : 4'b1011;
															assign node50902 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node50905 = (inp[3]) ? node50907 : 4'b1001;
															assign node50907 = (inp[15]) ? node50909 : 4'b1001;
																assign node50909 = (inp[0]) ? 4'b1001 : 4'b1011;
													assign node50912 = (inp[14]) ? node50924 : node50913;
														assign node50913 = (inp[15]) ? node50919 : node50914;
															assign node50914 = (inp[3]) ? node50916 : 4'b1011;
																assign node50916 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node50919 = (inp[3]) ? 4'b1001 : node50920;
																assign node50920 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node50924 = (inp[3]) ? 4'b1011 : node50925;
															assign node50925 = (inp[15]) ? node50927 : 4'b1011;
																assign node50927 = (inp[0]) ? 4'b1011 : 4'b1001;
										assign node50931 = (inp[4]) ? node50979 : node50932;
											assign node50932 = (inp[9]) ? node50972 : node50933;
												assign node50933 = (inp[14]) ? node50961 : node50934;
													assign node50934 = (inp[12]) ? node50948 : node50935;
														assign node50935 = (inp[0]) ? node50941 : node50936;
															assign node50936 = (inp[15]) ? 4'b1001 : node50937;
																assign node50937 = (inp[3]) ? 4'b1001 : 4'b1011;
															assign node50941 = (inp[15]) ? node50945 : node50942;
																assign node50942 = (inp[3]) ? 4'b1011 : 4'b1001;
																assign node50945 = (inp[3]) ? 4'b1001 : 4'b1011;
														assign node50948 = (inp[3]) ? node50954 : node50949;
															assign node50949 = (inp[15]) ? 4'b1011 : node50950;
																assign node50950 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node50954 = (inp[15]) ? node50958 : node50955;
																assign node50955 = (inp[0]) ? 4'b1011 : 4'b1001;
																assign node50958 = (inp[0]) ? 4'b1001 : 4'b1011;
													assign node50961 = (inp[0]) ? node50963 : 4'b1011;
														assign node50963 = (inp[12]) ? node50965 : 4'b1011;
															assign node50965 = (inp[3]) ? node50969 : node50966;
																assign node50966 = (inp[15]) ? 4'b1011 : 4'b1001;
																assign node50969 = (inp[15]) ? 4'b1001 : 4'b1011;
												assign node50972 = (inp[0]) ? node50976 : node50973;
													assign node50973 = (inp[15]) ? 4'b1111 : 4'b1101;
													assign node50976 = (inp[15]) ? 4'b1101 : 4'b1111;
											assign node50979 = (inp[9]) ? node50997 : node50980;
												assign node50980 = (inp[3]) ? node50990 : node50981;
													assign node50981 = (inp[12]) ? node50983 : 4'b1111;
														assign node50983 = (inp[15]) ? node50987 : node50984;
															assign node50984 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node50987 = (inp[0]) ? 4'b1101 : 4'b1111;
													assign node50990 = (inp[14]) ? 4'b1101 : node50991;
														assign node50991 = (inp[0]) ? node50993 : 4'b1101;
															assign node50993 = (inp[12]) ? 4'b1101 : 4'b1111;
												assign node50997 = (inp[12]) ? node51009 : node50998;
													assign node50998 = (inp[14]) ? node51006 : node50999;
														assign node50999 = (inp[0]) ? node51003 : node51000;
															assign node51000 = (inp[15]) ? 4'b1011 : 4'b1001;
															assign node51003 = (inp[15]) ? 4'b1001 : 4'b1011;
														assign node51006 = (inp[3]) ? 4'b1001 : 4'b1011;
													assign node51009 = (inp[3]) ? node51011 : 4'b1001;
														assign node51011 = (inp[15]) ? node51015 : node51012;
															assign node51012 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node51015 = (inp[0]) ? 4'b1001 : 4'b1011;
								assign node51018 = (inp[14]) ? node51270 : node51019;
									assign node51019 = (inp[2]) ? node51169 : node51020;
										assign node51020 = (inp[12]) ? node51094 : node51021;
											assign node51021 = (inp[5]) ? node51055 : node51022;
												assign node51022 = (inp[9]) ? node51042 : node51023;
													assign node51023 = (inp[4]) ? node51031 : node51024;
														assign node51024 = (inp[0]) ? node51028 : node51025;
															assign node51025 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node51028 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node51031 = (inp[15]) ? node51037 : node51032;
															assign node51032 = (inp[3]) ? node51034 : 4'b1111;
																assign node51034 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node51037 = (inp[0]) ? 4'b1101 : node51038;
																assign node51038 = (inp[3]) ? 4'b1111 : 4'b1101;
													assign node51042 = (inp[4]) ? 4'b1001 : node51043;
														assign node51043 = (inp[3]) ? node51049 : node51044;
															assign node51044 = (inp[0]) ? node51046 : 4'b1111;
																assign node51046 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node51049 = (inp[0]) ? 4'b1101 : node51050;
																assign node51050 = (inp[15]) ? 4'b1111 : 4'b1101;
												assign node51055 = (inp[15]) ? node51077 : node51056;
													assign node51056 = (inp[0]) ? node51062 : node51057;
														assign node51057 = (inp[9]) ? node51059 : 4'b1011;
															assign node51059 = (inp[4]) ? 4'b1001 : 4'b1101;
														assign node51062 = (inp[3]) ? node51070 : node51063;
															assign node51063 = (inp[9]) ? node51067 : node51064;
																assign node51064 = (inp[4]) ? 4'b1111 : 4'b1001;
																assign node51067 = (inp[4]) ? 4'b1011 : 4'b1111;
															assign node51070 = (inp[4]) ? node51074 : node51071;
																assign node51071 = (inp[9]) ? 4'b1111 : 4'b1011;
																assign node51074 = (inp[9]) ? 4'b1011 : 4'b1111;
													assign node51077 = (inp[0]) ? node51087 : node51078;
														assign node51078 = (inp[9]) ? node51084 : node51079;
															assign node51079 = (inp[4]) ? 4'b1111 : node51080;
																assign node51080 = (inp[3]) ? 4'b1011 : 4'b1001;
															assign node51084 = (inp[4]) ? 4'b1011 : 4'b1111;
														assign node51087 = (inp[4]) ? node51091 : node51088;
															assign node51088 = (inp[3]) ? 4'b1001 : 4'b1011;
															assign node51091 = (inp[9]) ? 4'b1001 : 4'b1101;
											assign node51094 = (inp[3]) ? node51126 : node51095;
												assign node51095 = (inp[9]) ? node51105 : node51096;
													assign node51096 = (inp[4]) ? 4'b1101 : node51097;
														assign node51097 = (inp[0]) ? node51101 : node51098;
															assign node51098 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node51101 = (inp[15]) ? 4'b1011 : 4'b1001;
													assign node51105 = (inp[4]) ? node51113 : node51106;
														assign node51106 = (inp[0]) ? 4'b1111 : node51107;
															assign node51107 = (inp[5]) ? 4'b1101 : node51108;
																assign node51108 = (inp[15]) ? 4'b1101 : 4'b1111;
														assign node51113 = (inp[15]) ? node51119 : node51114;
															assign node51114 = (inp[5]) ? 4'b1011 : node51115;
																assign node51115 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node51119 = (inp[5]) ? node51123 : node51120;
																assign node51120 = (inp[0]) ? 4'b1011 : 4'b1001;
																assign node51123 = (inp[0]) ? 4'b1001 : 4'b1011;
												assign node51126 = (inp[5]) ? node51150 : node51127;
													assign node51127 = (inp[15]) ? node51135 : node51128;
														assign node51128 = (inp[0]) ? node51132 : node51129;
															assign node51129 = (inp[4]) ? 4'b1001 : 4'b1101;
															assign node51132 = (inp[4]) ? 4'b1111 : 4'b1001;
														assign node51135 = (inp[0]) ? node51143 : node51136;
															assign node51136 = (inp[9]) ? node51140 : node51137;
																assign node51137 = (inp[4]) ? 4'b1111 : 4'b1001;
																assign node51140 = (inp[4]) ? 4'b1011 : 4'b1111;
															assign node51143 = (inp[9]) ? node51147 : node51144;
																assign node51144 = (inp[4]) ? 4'b1101 : 4'b1011;
																assign node51147 = (inp[4]) ? 4'b1001 : 4'b1101;
													assign node51150 = (inp[0]) ? node51158 : node51151;
														assign node51151 = (inp[15]) ? 4'b1011 : node51152;
															assign node51152 = (inp[9]) ? 4'b1001 : node51153;
																assign node51153 = (inp[4]) ? 4'b1101 : 4'b1001;
														assign node51158 = (inp[15]) ? node51164 : node51159;
															assign node51159 = (inp[9]) ? node51161 : 4'b1011;
																assign node51161 = (inp[4]) ? 4'b1011 : 4'b1111;
															assign node51164 = (inp[9]) ? node51166 : 4'b1101;
																assign node51166 = (inp[4]) ? 4'b1001 : 4'b1101;
										assign node51169 = (inp[4]) ? node51217 : node51170;
											assign node51170 = (inp[9]) ? node51184 : node51171;
												assign node51171 = (inp[15]) ? node51177 : node51172;
													assign node51172 = (inp[0]) ? 4'b1000 : node51173;
														assign node51173 = (inp[3]) ? 4'b1000 : 4'b1010;
													assign node51177 = (inp[0]) ? node51179 : 4'b1000;
														assign node51179 = (inp[5]) ? node51181 : 4'b1010;
															assign node51181 = (inp[3]) ? 4'b1000 : 4'b1010;
												assign node51184 = (inp[12]) ? node51204 : node51185;
													assign node51185 = (inp[0]) ? node51193 : node51186;
														assign node51186 = (inp[15]) ? node51188 : 4'b1100;
															assign node51188 = (inp[5]) ? 4'b1110 : node51189;
																assign node51189 = (inp[3]) ? 4'b1110 : 4'b1100;
														assign node51193 = (inp[15]) ? node51199 : node51194;
															assign node51194 = (inp[3]) ? 4'b1110 : node51195;
																assign node51195 = (inp[5]) ? 4'b1110 : 4'b1100;
															assign node51199 = (inp[3]) ? 4'b1100 : node51200;
																assign node51200 = (inp[5]) ? 4'b1100 : 4'b1110;
													assign node51204 = (inp[15]) ? 4'b1100 : node51205;
														assign node51205 = (inp[0]) ? node51211 : node51206;
															assign node51206 = (inp[3]) ? 4'b1100 : node51207;
																assign node51207 = (inp[5]) ? 4'b1100 : 4'b1110;
															assign node51211 = (inp[3]) ? 4'b1110 : node51212;
																assign node51212 = (inp[5]) ? 4'b1110 : 4'b1100;
											assign node51217 = (inp[9]) ? node51239 : node51218;
												assign node51218 = (inp[3]) ? node51226 : node51219;
													assign node51219 = (inp[5]) ? 4'b1110 : node51220;
														assign node51220 = (inp[0]) ? 4'b1100 : node51221;
															assign node51221 = (inp[15]) ? 4'b1100 : 4'b1110;
													assign node51226 = (inp[5]) ? node51234 : node51227;
														assign node51227 = (inp[0]) ? node51231 : node51228;
															assign node51228 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node51231 = (inp[15]) ? 4'b1100 : 4'b1110;
														assign node51234 = (inp[15]) ? node51236 : 4'b1100;
															assign node51236 = (inp[0]) ? 4'b1100 : 4'b1110;
												assign node51239 = (inp[5]) ? node51253 : node51240;
													assign node51240 = (inp[3]) ? node51246 : node51241;
														assign node51241 = (inp[0]) ? node51243 : 4'b1010;
															assign node51243 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node51246 = (inp[15]) ? node51250 : node51247;
															assign node51247 = (inp[0]) ? 4'b1010 : 4'b1000;
															assign node51250 = (inp[0]) ? 4'b1000 : 4'b1010;
													assign node51253 = (inp[12]) ? node51263 : node51254;
														assign node51254 = (inp[3]) ? node51260 : node51255;
															assign node51255 = (inp[15]) ? 4'b1000 : node51256;
																assign node51256 = (inp[0]) ? 4'b1010 : 4'b1000;
															assign node51260 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node51263 = (inp[15]) ? node51267 : node51264;
															assign node51264 = (inp[3]) ? 4'b1000 : 4'b1010;
															assign node51267 = (inp[0]) ? 4'b1000 : 4'b1010;
									assign node51270 = (inp[4]) ? node51330 : node51271;
										assign node51271 = (inp[9]) ? node51295 : node51272;
											assign node51272 = (inp[15]) ? node51284 : node51273;
												assign node51273 = (inp[0]) ? node51279 : node51274;
													assign node51274 = (inp[3]) ? node51276 : 4'b1010;
														assign node51276 = (inp[5]) ? 4'b1000 : 4'b1010;
													assign node51279 = (inp[5]) ? node51281 : 4'b1000;
														assign node51281 = (inp[3]) ? 4'b1010 : 4'b1000;
												assign node51284 = (inp[0]) ? node51290 : node51285;
													assign node51285 = (inp[5]) ? node51287 : 4'b1000;
														assign node51287 = (inp[3]) ? 4'b1010 : 4'b1000;
													assign node51290 = (inp[3]) ? node51292 : 4'b1010;
														assign node51292 = (inp[5]) ? 4'b1000 : 4'b1010;
											assign node51295 = (inp[2]) ? node51315 : node51296;
												assign node51296 = (inp[15]) ? node51308 : node51297;
													assign node51297 = (inp[0]) ? node51303 : node51298;
														assign node51298 = (inp[3]) ? 4'b1100 : node51299;
															assign node51299 = (inp[5]) ? 4'b1100 : 4'b1110;
														assign node51303 = (inp[3]) ? 4'b1110 : node51304;
															assign node51304 = (inp[5]) ? 4'b1110 : 4'b1100;
													assign node51308 = (inp[0]) ? 4'b1100 : node51309;
														assign node51309 = (inp[5]) ? 4'b1110 : node51310;
															assign node51310 = (inp[12]) ? 4'b1110 : 4'b1100;
												assign node51315 = (inp[0]) ? node51319 : node51316;
													assign node51316 = (inp[15]) ? 4'b1110 : 4'b1100;
													assign node51319 = (inp[15]) ? node51325 : node51320;
														assign node51320 = (inp[5]) ? 4'b1110 : node51321;
															assign node51321 = (inp[3]) ? 4'b1110 : 4'b1100;
														assign node51325 = (inp[3]) ? 4'b1100 : node51326;
															assign node51326 = (inp[5]) ? 4'b1100 : 4'b1110;
										assign node51330 = (inp[9]) ? node51396 : node51331;
											assign node51331 = (inp[2]) ? node51369 : node51332;
												assign node51332 = (inp[12]) ? node51354 : node51333;
													assign node51333 = (inp[3]) ? node51345 : node51334;
														assign node51334 = (inp[5]) ? node51340 : node51335;
															assign node51335 = (inp[0]) ? node51337 : 4'b1100;
																assign node51337 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node51340 = (inp[15]) ? node51342 : 4'b1110;
																assign node51342 = (inp[0]) ? 4'b1100 : 4'b1110;
														assign node51345 = (inp[5]) ? node51347 : 4'b1110;
															assign node51347 = (inp[15]) ? node51351 : node51348;
																assign node51348 = (inp[0]) ? 4'b1110 : 4'b1100;
																assign node51351 = (inp[0]) ? 4'b1100 : 4'b1110;
													assign node51354 = (inp[5]) ? node51362 : node51355;
														assign node51355 = (inp[3]) ? node51357 : 4'b1100;
															assign node51357 = (inp[0]) ? 4'b1100 : node51358;
																assign node51358 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node51362 = (inp[15]) ? node51366 : node51363;
															assign node51363 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node51366 = (inp[0]) ? 4'b1100 : 4'b1110;
												assign node51369 = (inp[5]) ? node51391 : node51370;
													assign node51370 = (inp[12]) ? node51380 : node51371;
														assign node51371 = (inp[0]) ? node51373 : 4'b1100;
															assign node51373 = (inp[3]) ? node51377 : node51374;
																assign node51374 = (inp[15]) ? 4'b1110 : 4'b1100;
																assign node51377 = (inp[15]) ? 4'b1100 : 4'b1110;
														assign node51380 = (inp[0]) ? node51386 : node51381;
															assign node51381 = (inp[3]) ? 4'b1110 : node51382;
																assign node51382 = (inp[15]) ? 4'b1100 : 4'b1110;
															assign node51386 = (inp[3]) ? 4'b1100 : node51387;
																assign node51387 = (inp[15]) ? 4'b1110 : 4'b1100;
													assign node51391 = (inp[15]) ? node51393 : 4'b1100;
														assign node51393 = (inp[0]) ? 4'b1100 : 4'b1110;
											assign node51396 = (inp[15]) ? node51408 : node51397;
												assign node51397 = (inp[0]) ? node51403 : node51398;
													assign node51398 = (inp[5]) ? 4'b1000 : node51399;
														assign node51399 = (inp[3]) ? 4'b1000 : 4'b1010;
													assign node51403 = (inp[5]) ? 4'b1010 : node51404;
														assign node51404 = (inp[3]) ? 4'b1010 : 4'b1000;
												assign node51408 = (inp[0]) ? node51410 : 4'b1010;
													assign node51410 = (inp[3]) ? 4'b1000 : node51411;
														assign node51411 = (inp[5]) ? 4'b1000 : 4'b1010;
					assign node51415 = (inp[1]) ? node53179 : node51416;
						assign node51416 = (inp[7]) ? node52328 : node51417;
							assign node51417 = (inp[8]) ? node51935 : node51418;
								assign node51418 = (inp[14]) ? node51716 : node51419;
									assign node51419 = (inp[2]) ? node51563 : node51420;
										assign node51420 = (inp[15]) ? node51480 : node51421;
											assign node51421 = (inp[3]) ? node51459 : node51422;
												assign node51422 = (inp[0]) ? node51442 : node51423;
													assign node51423 = (inp[5]) ? node51431 : node51424;
														assign node51424 = (inp[9]) ? 4'b0011 : node51425;
															assign node51425 = (inp[12]) ? node51427 : 4'b0111;
																assign node51427 = (inp[4]) ? 4'b0111 : 4'b0011;
														assign node51431 = (inp[4]) ? node51437 : node51432;
															assign node51432 = (inp[9]) ? 4'b0101 : node51433;
																assign node51433 = (inp[12]) ? 4'b0011 : 4'b0111;
															assign node51437 = (inp[12]) ? node51439 : 4'b0101;
																assign node51439 = (inp[9]) ? 4'b0001 : 4'b0101;
													assign node51442 = (inp[5]) ? node51454 : node51443;
														assign node51443 = (inp[9]) ? node51449 : node51444;
															assign node51444 = (inp[12]) ? 4'b0101 : node51445;
																assign node51445 = (inp[4]) ? 4'b0001 : 4'b0101;
															assign node51449 = (inp[4]) ? node51451 : 4'b0001;
																assign node51451 = (inp[12]) ? 4'b0001 : 4'b0101;
														assign node51454 = (inp[9]) ? 4'b0111 : node51455;
															assign node51455 = (inp[4]) ? 4'b0111 : 4'b0001;
												assign node51459 = (inp[0]) ? node51471 : node51460;
													assign node51460 = (inp[12]) ? 4'b0101 : node51461;
														assign node51461 = (inp[9]) ? node51465 : node51462;
															assign node51462 = (inp[5]) ? 4'b0101 : 4'b0111;
															assign node51465 = (inp[4]) ? 4'b0101 : node51466;
																assign node51466 = (inp[5]) ? 4'b0001 : 4'b0011;
													assign node51471 = (inp[4]) ? node51475 : node51472;
														assign node51472 = (inp[12]) ? 4'b0111 : 4'b0101;
														assign node51475 = (inp[9]) ? node51477 : 4'b0011;
															assign node51477 = (inp[12]) ? 4'b0011 : 4'b0111;
											assign node51480 = (inp[5]) ? node51518 : node51481;
												assign node51481 = (inp[0]) ? node51499 : node51482;
													assign node51482 = (inp[9]) ? node51490 : node51483;
														assign node51483 = (inp[12]) ? node51487 : node51484;
															assign node51484 = (inp[4]) ? 4'b0001 : 4'b0101;
															assign node51487 = (inp[4]) ? 4'b0101 : 4'b0001;
														assign node51490 = (inp[3]) ? node51492 : 4'b0001;
															assign node51492 = (inp[4]) ? node51496 : node51493;
																assign node51493 = (inp[12]) ? 4'b0111 : 4'b0001;
																assign node51496 = (inp[12]) ? 4'b0011 : 4'b0111;
													assign node51499 = (inp[3]) ? node51507 : node51500;
														assign node51500 = (inp[4]) ? node51502 : 4'b0111;
															assign node51502 = (inp[12]) ? 4'b0011 : node51503;
																assign node51503 = (inp[9]) ? 4'b0111 : 4'b0011;
														assign node51507 = (inp[9]) ? node51513 : node51508;
															assign node51508 = (inp[12]) ? node51510 : 4'b0011;
																assign node51510 = (inp[4]) ? 4'b0101 : 4'b0011;
															assign node51513 = (inp[12]) ? node51515 : 4'b0101;
																assign node51515 = (inp[4]) ? 4'b0001 : 4'b0101;
												assign node51518 = (inp[0]) ? node51546 : node51519;
													assign node51519 = (inp[3]) ? node51533 : node51520;
														assign node51520 = (inp[4]) ? node51528 : node51521;
															assign node51521 = (inp[9]) ? node51525 : node51522;
																assign node51522 = (inp[12]) ? 4'b0001 : 4'b0101;
																assign node51525 = (inp[12]) ? 4'b0111 : 4'b0001;
															assign node51528 = (inp[12]) ? node51530 : 4'b0111;
																assign node51530 = (inp[9]) ? 4'b0011 : 4'b0111;
														assign node51533 = (inp[4]) ? node51541 : node51534;
															assign node51534 = (inp[12]) ? node51538 : node51535;
																assign node51535 = (inp[9]) ? 4'b0011 : 4'b0111;
																assign node51538 = (inp[9]) ? 4'b0111 : 4'b0011;
															assign node51541 = (inp[12]) ? node51543 : 4'b0011;
																assign node51543 = (inp[9]) ? 4'b0011 : 4'b0111;
													assign node51546 = (inp[12]) ? node51558 : node51547;
														assign node51547 = (inp[3]) ? node51553 : node51548;
															assign node51548 = (inp[9]) ? 4'b0011 : node51549;
																assign node51549 = (inp[4]) ? 4'b0011 : 4'b0111;
															assign node51553 = (inp[4]) ? node51555 : 4'b0001;
																assign node51555 = (inp[9]) ? 4'b0101 : 4'b0001;
														assign node51558 = (inp[9]) ? node51560 : 4'b0101;
															assign node51560 = (inp[4]) ? 4'b0001 : 4'b0101;
										assign node51563 = (inp[3]) ? node51643 : node51564;
											assign node51564 = (inp[5]) ? node51608 : node51565;
												assign node51565 = (inp[0]) ? node51589 : node51566;
													assign node51566 = (inp[15]) ? node51580 : node51567;
														assign node51567 = (inp[4]) ? node51573 : node51568;
															assign node51568 = (inp[12]) ? node51570 : 4'b0110;
																assign node51570 = (inp[9]) ? 4'b0110 : 4'b0010;
															assign node51573 = (inp[12]) ? node51577 : node51574;
																assign node51574 = (inp[9]) ? 4'b0110 : 4'b0010;
																assign node51577 = (inp[9]) ? 4'b0010 : 4'b0110;
														assign node51580 = (inp[9]) ? 4'b0000 : node51581;
															assign node51581 = (inp[4]) ? node51585 : node51582;
																assign node51582 = (inp[12]) ? 4'b0000 : 4'b0100;
																assign node51585 = (inp[12]) ? 4'b0100 : 4'b0000;
													assign node51589 = (inp[15]) ? node51599 : node51590;
														assign node51590 = (inp[9]) ? node51592 : 4'b0100;
															assign node51592 = (inp[12]) ? node51596 : node51593;
																assign node51593 = (inp[4]) ? 4'b0100 : 4'b0000;
																assign node51596 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node51599 = (inp[4]) ? 4'b0110 : node51600;
															assign node51600 = (inp[9]) ? node51604 : node51601;
																assign node51601 = (inp[12]) ? 4'b0010 : 4'b0110;
																assign node51604 = (inp[12]) ? 4'b0110 : 4'b0010;
												assign node51608 = (inp[15]) ? node51628 : node51609;
													assign node51609 = (inp[9]) ? node51619 : node51610;
														assign node51610 = (inp[0]) ? node51614 : node51611;
															assign node51611 = (inp[12]) ? 4'b0010 : 4'b0110;
															assign node51614 = (inp[4]) ? 4'b0110 : node51615;
																assign node51615 = (inp[12]) ? 4'b0000 : 4'b0100;
														assign node51619 = (inp[0]) ? node51625 : node51620;
															assign node51620 = (inp[12]) ? node51622 : 4'b0100;
																assign node51622 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node51625 = (inp[12]) ? 4'b0110 : 4'b0000;
													assign node51628 = (inp[0]) ? node51638 : node51629;
														assign node51629 = (inp[12]) ? 4'b0110 : node51630;
															assign node51630 = (inp[4]) ? node51634 : node51631;
																assign node51631 = (inp[9]) ? 4'b0000 : 4'b0100;
																assign node51634 = (inp[9]) ? 4'b0110 : 4'b0000;
														assign node51638 = (inp[4]) ? 4'b0100 : node51639;
															assign node51639 = (inp[9]) ? 4'b0100 : 4'b0110;
											assign node51643 = (inp[12]) ? node51685 : node51644;
												assign node51644 = (inp[15]) ? node51668 : node51645;
													assign node51645 = (inp[0]) ? node51653 : node51646;
														assign node51646 = (inp[9]) ? node51650 : node51647;
															assign node51647 = (inp[5]) ? 4'b0100 : 4'b0010;
															assign node51650 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node51653 = (inp[5]) ? node51661 : node51654;
															assign node51654 = (inp[9]) ? node51658 : node51655;
																assign node51655 = (inp[4]) ? 4'b0000 : 4'b0100;
																assign node51658 = (inp[4]) ? 4'b0110 : 4'b0000;
															assign node51661 = (inp[4]) ? node51665 : node51662;
																assign node51662 = (inp[9]) ? 4'b0010 : 4'b0110;
																assign node51665 = (inp[9]) ? 4'b0110 : 4'b0010;
													assign node51668 = (inp[0]) ? node51676 : node51669;
														assign node51669 = (inp[5]) ? 4'b0010 : node51670;
															assign node51670 = (inp[4]) ? node51672 : 4'b0000;
																assign node51672 = (inp[9]) ? 4'b0110 : 4'b0000;
														assign node51676 = (inp[5]) ? node51678 : 4'b0100;
															assign node51678 = (inp[9]) ? node51682 : node51679;
																assign node51679 = (inp[4]) ? 4'b0000 : 4'b0100;
																assign node51682 = (inp[4]) ? 4'b0100 : 4'b0000;
												assign node51685 = (inp[0]) ? node51701 : node51686;
													assign node51686 = (inp[15]) ? node51692 : node51687;
														assign node51687 = (inp[5]) ? 4'b0000 : node51688;
															assign node51688 = (inp[9]) ? 4'b0100 : 4'b0010;
														assign node51692 = (inp[4]) ? node51698 : node51693;
															assign node51693 = (inp[5]) ? node51695 : 4'b0000;
																assign node51695 = (inp[9]) ? 4'b0110 : 4'b0010;
															assign node51698 = (inp[9]) ? 4'b0010 : 4'b0110;
													assign node51701 = (inp[15]) ? node51709 : node51702;
														assign node51702 = (inp[9]) ? node51706 : node51703;
															assign node51703 = (inp[4]) ? 4'b0110 : 4'b0000;
															assign node51706 = (inp[4]) ? 4'b0010 : 4'b0110;
														assign node51709 = (inp[9]) ? node51713 : node51710;
															assign node51710 = (inp[4]) ? 4'b0100 : 4'b0010;
															assign node51713 = (inp[4]) ? 4'b0000 : 4'b0100;
									assign node51716 = (inp[3]) ? node51838 : node51717;
										assign node51717 = (inp[0]) ? node51775 : node51718;
											assign node51718 = (inp[15]) ? node51742 : node51719;
												assign node51719 = (inp[9]) ? node51731 : node51720;
													assign node51720 = (inp[2]) ? node51726 : node51721;
														assign node51721 = (inp[12]) ? node51723 : 4'b0010;
															assign node51723 = (inp[4]) ? 4'b0110 : 4'b0010;
														assign node51726 = (inp[12]) ? 4'b0010 : node51727;
															assign node51727 = (inp[4]) ? 4'b0010 : 4'b0110;
													assign node51731 = (inp[5]) ? node51735 : node51732;
														assign node51732 = (inp[4]) ? 4'b0110 : 4'b0010;
														assign node51735 = (inp[12]) ? node51739 : node51736;
															assign node51736 = (inp[4]) ? 4'b0100 : 4'b0010;
															assign node51739 = (inp[4]) ? 4'b0000 : 4'b0100;
												assign node51742 = (inp[5]) ? node51760 : node51743;
													assign node51743 = (inp[4]) ? node51745 : 4'b0000;
														assign node51745 = (inp[2]) ? node51753 : node51746;
															assign node51746 = (inp[9]) ? node51750 : node51747;
																assign node51747 = (inp[12]) ? 4'b0100 : 4'b0000;
																assign node51750 = (inp[12]) ? 4'b0000 : 4'b0100;
															assign node51753 = (inp[9]) ? node51757 : node51754;
																assign node51754 = (inp[12]) ? 4'b0100 : 4'b0000;
																assign node51757 = (inp[12]) ? 4'b0000 : 4'b0100;
													assign node51760 = (inp[9]) ? node51768 : node51761;
														assign node51761 = (inp[4]) ? node51765 : node51762;
															assign node51762 = (inp[12]) ? 4'b0000 : 4'b0100;
															assign node51765 = (inp[12]) ? 4'b0110 : 4'b0000;
														assign node51768 = (inp[4]) ? node51772 : node51769;
															assign node51769 = (inp[12]) ? 4'b0110 : 4'b0000;
															assign node51772 = (inp[12]) ? 4'b0010 : 4'b0110;
											assign node51775 = (inp[15]) ? node51811 : node51776;
												assign node51776 = (inp[5]) ? node51796 : node51777;
													assign node51777 = (inp[4]) ? node51791 : node51778;
														assign node51778 = (inp[2]) ? node51786 : node51779;
															assign node51779 = (inp[9]) ? node51783 : node51780;
																assign node51780 = (inp[12]) ? 4'b0000 : 4'b0100;
																assign node51783 = (inp[12]) ? 4'b0100 : 4'b0000;
															assign node51786 = (inp[12]) ? 4'b0000 : node51787;
																assign node51787 = (inp[9]) ? 4'b0000 : 4'b0100;
														assign node51791 = (inp[9]) ? node51793 : 4'b0100;
															assign node51793 = (inp[12]) ? 4'b0000 : 4'b0100;
													assign node51796 = (inp[4]) ? node51802 : node51797;
														assign node51797 = (inp[9]) ? 4'b0000 : node51798;
															assign node51798 = (inp[12]) ? 4'b0000 : 4'b0100;
														assign node51802 = (inp[2]) ? node51804 : 4'b0000;
															assign node51804 = (inp[12]) ? node51808 : node51805;
																assign node51805 = (inp[9]) ? 4'b0110 : 4'b0000;
																assign node51808 = (inp[9]) ? 4'b0010 : 4'b0110;
												assign node51811 = (inp[5]) ? node51829 : node51812;
													assign node51812 = (inp[4]) ? node51822 : node51813;
														assign node51813 = (inp[2]) ? 4'b0110 : node51814;
															assign node51814 = (inp[12]) ? node51818 : node51815;
																assign node51815 = (inp[9]) ? 4'b0010 : 4'b0110;
																assign node51818 = (inp[9]) ? 4'b0110 : 4'b0010;
														assign node51822 = (inp[2]) ? 4'b0010 : node51823;
															assign node51823 = (inp[12]) ? 4'b0110 : node51824;
																assign node51824 = (inp[9]) ? 4'b0110 : 4'b0010;
													assign node51829 = (inp[9]) ? 4'b0100 : node51830;
														assign node51830 = (inp[4]) ? node51834 : node51831;
															assign node51831 = (inp[12]) ? 4'b0010 : 4'b0110;
															assign node51834 = (inp[12]) ? 4'b0100 : 4'b0010;
										assign node51838 = (inp[12]) ? node51896 : node51839;
											assign node51839 = (inp[5]) ? node51873 : node51840;
												assign node51840 = (inp[9]) ? node51854 : node51841;
													assign node51841 = (inp[4]) ? node51849 : node51842;
														assign node51842 = (inp[15]) ? node51846 : node51843;
															assign node51843 = (inp[0]) ? 4'b0100 : 4'b0110;
															assign node51846 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node51849 = (inp[15]) ? node51851 : 4'b0000;
															assign node51851 = (inp[0]) ? 4'b0010 : 4'b0000;
													assign node51854 = (inp[4]) ? node51868 : node51855;
														assign node51855 = (inp[2]) ? node51863 : node51856;
															assign node51856 = (inp[0]) ? node51860 : node51857;
																assign node51857 = (inp[15]) ? 4'b0000 : 4'b0010;
																assign node51860 = (inp[15]) ? 4'b0010 : 4'b0000;
															assign node51863 = (inp[15]) ? 4'b0010 : node51864;
																assign node51864 = (inp[0]) ? 4'b0000 : 4'b0010;
														assign node51868 = (inp[0]) ? node51870 : 4'b0100;
															assign node51870 = (inp[15]) ? 4'b0100 : 4'b0110;
												assign node51873 = (inp[15]) ? node51883 : node51874;
													assign node51874 = (inp[0]) ? node51876 : 4'b0000;
														assign node51876 = (inp[9]) ? node51880 : node51877;
															assign node51877 = (inp[4]) ? 4'b0010 : 4'b0110;
															assign node51880 = (inp[4]) ? 4'b0110 : 4'b0010;
													assign node51883 = (inp[0]) ? node51891 : node51884;
														assign node51884 = (inp[9]) ? node51888 : node51885;
															assign node51885 = (inp[2]) ? 4'b0010 : 4'b0110;
															assign node51888 = (inp[4]) ? 4'b0110 : 4'b0010;
														assign node51891 = (inp[9]) ? 4'b0000 : node51892;
															assign node51892 = (inp[4]) ? 4'b0000 : 4'b0100;
											assign node51896 = (inp[0]) ? node51916 : node51897;
												assign node51897 = (inp[15]) ? node51907 : node51898;
													assign node51898 = (inp[9]) ? node51904 : node51899;
														assign node51899 = (inp[4]) ? 4'b0100 : node51900;
															assign node51900 = (inp[5]) ? 4'b0000 : 4'b0010;
														assign node51904 = (inp[4]) ? 4'b0000 : 4'b0100;
													assign node51907 = (inp[9]) ? node51913 : node51908;
														assign node51908 = (inp[4]) ? 4'b0110 : node51909;
															assign node51909 = (inp[5]) ? 4'b0010 : 4'b0000;
														assign node51913 = (inp[4]) ? 4'b0010 : 4'b0110;
												assign node51916 = (inp[15]) ? node51926 : node51917;
													assign node51917 = (inp[5]) ? node51919 : 4'b0110;
														assign node51919 = (inp[9]) ? node51923 : node51920;
															assign node51920 = (inp[4]) ? 4'b0110 : 4'b0010;
															assign node51923 = (inp[4]) ? 4'b0010 : 4'b0110;
													assign node51926 = (inp[9]) ? node51932 : node51927;
														assign node51927 = (inp[4]) ? 4'b0100 : node51928;
															assign node51928 = (inp[5]) ? 4'b0000 : 4'b0010;
														assign node51932 = (inp[4]) ? 4'b0000 : 4'b0100;
								assign node51935 = (inp[14]) ? node52169 : node51936;
									assign node51936 = (inp[2]) ? node52084 : node51937;
										assign node51937 = (inp[9]) ? node52011 : node51938;
											assign node51938 = (inp[5]) ? node51974 : node51939;
												assign node51939 = (inp[3]) ? node51957 : node51940;
													assign node51940 = (inp[15]) ? node51948 : node51941;
														assign node51941 = (inp[0]) ? 4'b0000 : node51942;
															assign node51942 = (inp[12]) ? 4'b0010 : node51943;
																assign node51943 = (inp[4]) ? 4'b0010 : 4'b0110;
														assign node51948 = (inp[0]) ? node51950 : 4'b0100;
															assign node51950 = (inp[12]) ? node51954 : node51951;
																assign node51951 = (inp[4]) ? 4'b0010 : 4'b0110;
																assign node51954 = (inp[4]) ? 4'b0110 : 4'b0010;
													assign node51957 = (inp[15]) ? node51959 : 4'b0100;
														assign node51959 = (inp[0]) ? node51967 : node51960;
															assign node51960 = (inp[12]) ? node51964 : node51961;
																assign node51961 = (inp[4]) ? 4'b0000 : 4'b0100;
																assign node51964 = (inp[4]) ? 4'b0110 : 4'b0000;
															assign node51967 = (inp[4]) ? node51971 : node51968;
																assign node51968 = (inp[12]) ? 4'b0010 : 4'b0110;
																assign node51971 = (inp[12]) ? 4'b0100 : 4'b0010;
												assign node51974 = (inp[0]) ? node51996 : node51975;
													assign node51975 = (inp[15]) ? node51985 : node51976;
														assign node51976 = (inp[4]) ? 4'b0100 : node51977;
															assign node51977 = (inp[3]) ? node51981 : node51978;
																assign node51978 = (inp[12]) ? 4'b0010 : 4'b0110;
																assign node51981 = (inp[12]) ? 4'b0000 : 4'b0100;
														assign node51985 = (inp[3]) ? node51993 : node51986;
															assign node51986 = (inp[4]) ? node51990 : node51987;
																assign node51987 = (inp[12]) ? 4'b0000 : 4'b0100;
																assign node51990 = (inp[12]) ? 4'b0110 : 4'b0000;
															assign node51993 = (inp[4]) ? 4'b0010 : 4'b0110;
													assign node51996 = (inp[15]) ? node52006 : node51997;
														assign node51997 = (inp[3]) ? 4'b0110 : node51998;
															assign node51998 = (inp[4]) ? node52002 : node51999;
																assign node51999 = (inp[12]) ? 4'b0000 : 4'b0100;
																assign node52002 = (inp[12]) ? 4'b0110 : 4'b0000;
														assign node52006 = (inp[3]) ? node52008 : 4'b0100;
															assign node52008 = (inp[4]) ? 4'b0000 : 4'b0100;
											assign node52011 = (inp[15]) ? node52043 : node52012;
												assign node52012 = (inp[0]) ? node52030 : node52013;
													assign node52013 = (inp[5]) ? node52027 : node52014;
														assign node52014 = (inp[3]) ? node52022 : node52015;
															assign node52015 = (inp[12]) ? node52019 : node52016;
																assign node52016 = (inp[4]) ? 4'b0110 : 4'b0010;
																assign node52019 = (inp[4]) ? 4'b0010 : 4'b0110;
															assign node52022 = (inp[12]) ? node52024 : 4'b0010;
																assign node52024 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node52027 = (inp[12]) ? 4'b0000 : 4'b0100;
													assign node52030 = (inp[4]) ? node52040 : node52031;
														assign node52031 = (inp[12]) ? node52035 : node52032;
															assign node52032 = (inp[5]) ? 4'b0010 : 4'b0000;
															assign node52035 = (inp[3]) ? 4'b0110 : node52036;
																assign node52036 = (inp[5]) ? 4'b0110 : 4'b0100;
														assign node52040 = (inp[12]) ? 4'b0010 : 4'b0110;
												assign node52043 = (inp[0]) ? node52067 : node52044;
													assign node52044 = (inp[5]) ? node52056 : node52045;
														assign node52045 = (inp[3]) ? node52051 : node52046;
															assign node52046 = (inp[12]) ? node52048 : 4'b0100;
																assign node52048 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node52051 = (inp[4]) ? node52053 : 4'b0000;
																assign node52053 = (inp[12]) ? 4'b0010 : 4'b0110;
														assign node52056 = (inp[3]) ? node52062 : node52057;
															assign node52057 = (inp[12]) ? node52059 : 4'b0000;
																assign node52059 = (inp[4]) ? 4'b0010 : 4'b0110;
															assign node52062 = (inp[4]) ? node52064 : 4'b0110;
																assign node52064 = (inp[12]) ? 4'b0010 : 4'b0110;
													assign node52067 = (inp[5]) ? node52075 : node52068;
														assign node52068 = (inp[3]) ? node52070 : 4'b0010;
															assign node52070 = (inp[4]) ? node52072 : 4'b0010;
																assign node52072 = (inp[12]) ? 4'b0000 : 4'b0100;
														assign node52075 = (inp[3]) ? 4'b0000 : node52076;
															assign node52076 = (inp[12]) ? node52080 : node52077;
																assign node52077 = (inp[4]) ? 4'b0100 : 4'b0010;
																assign node52080 = (inp[4]) ? 4'b0000 : 4'b0100;
										assign node52084 = (inp[0]) ? node52118 : node52085;
											assign node52085 = (inp[4]) ? node52103 : node52086;
												assign node52086 = (inp[9]) ? node52098 : node52087;
													assign node52087 = (inp[15]) ? node52093 : node52088;
														assign node52088 = (inp[3]) ? node52090 : 4'b1011;
															assign node52090 = (inp[5]) ? 4'b1001 : 4'b1011;
														assign node52093 = (inp[3]) ? node52095 : 4'b1001;
															assign node52095 = (inp[5]) ? 4'b1011 : 4'b1001;
													assign node52098 = (inp[15]) ? node52100 : 4'b1101;
														assign node52100 = (inp[5]) ? 4'b1111 : 4'b1101;
												assign node52103 = (inp[9]) ? node52113 : node52104;
													assign node52104 = (inp[15]) ? node52110 : node52105;
														assign node52105 = (inp[5]) ? 4'b1101 : node52106;
															assign node52106 = (inp[3]) ? 4'b1101 : 4'b1111;
														assign node52110 = (inp[12]) ? 4'b1101 : 4'b1111;
													assign node52113 = (inp[5]) ? node52115 : 4'b1011;
														assign node52115 = (inp[15]) ? 4'b1011 : 4'b1001;
											assign node52118 = (inp[15]) ? node52146 : node52119;
												assign node52119 = (inp[3]) ? node52137 : node52120;
													assign node52120 = (inp[5]) ? node52126 : node52121;
														assign node52121 = (inp[4]) ? 4'b1001 : node52122;
															assign node52122 = (inp[9]) ? 4'b1101 : 4'b1001;
														assign node52126 = (inp[12]) ? node52132 : node52127;
															assign node52127 = (inp[9]) ? node52129 : 4'b1111;
																assign node52129 = (inp[4]) ? 4'b1011 : 4'b1111;
															assign node52132 = (inp[9]) ? node52134 : 4'b1001;
																assign node52134 = (inp[4]) ? 4'b1011 : 4'b1111;
													assign node52137 = (inp[4]) ? node52143 : node52138;
														assign node52138 = (inp[9]) ? 4'b1111 : node52139;
															assign node52139 = (inp[5]) ? 4'b1011 : 4'b1001;
														assign node52143 = (inp[9]) ? 4'b1011 : 4'b1111;
												assign node52146 = (inp[3]) ? node52154 : node52147;
													assign node52147 = (inp[9]) ? node52151 : node52148;
														assign node52148 = (inp[4]) ? 4'b1111 : 4'b1011;
														assign node52151 = (inp[5]) ? 4'b1101 : 4'b1111;
													assign node52154 = (inp[12]) ? node52160 : node52155;
														assign node52155 = (inp[9]) ? node52157 : 4'b1101;
															assign node52157 = (inp[4]) ? 4'b1001 : 4'b1101;
														assign node52160 = (inp[5]) ? node52164 : node52161;
															assign node52161 = (inp[9]) ? 4'b1101 : 4'b1011;
															assign node52164 = (inp[4]) ? node52166 : 4'b1001;
																assign node52166 = (inp[9]) ? 4'b1001 : 4'b1101;
									assign node52169 = (inp[3]) ? node52249 : node52170;
										assign node52170 = (inp[0]) ? node52214 : node52171;
											assign node52171 = (inp[15]) ? node52193 : node52172;
												assign node52172 = (inp[5]) ? node52186 : node52173;
													assign node52173 = (inp[2]) ? node52181 : node52174;
														assign node52174 = (inp[9]) ? node52178 : node52175;
															assign node52175 = (inp[4]) ? 4'b1111 : 4'b1011;
															assign node52178 = (inp[4]) ? 4'b1011 : 4'b1111;
														assign node52181 = (inp[12]) ? node52183 : 4'b1111;
															assign node52183 = (inp[9]) ? 4'b1011 : 4'b1111;
													assign node52186 = (inp[9]) ? node52190 : node52187;
														assign node52187 = (inp[4]) ? 4'b1101 : 4'b1011;
														assign node52190 = (inp[4]) ? 4'b1001 : 4'b1101;
												assign node52193 = (inp[5]) ? node52201 : node52194;
													assign node52194 = (inp[4]) ? node52198 : node52195;
														assign node52195 = (inp[9]) ? 4'b1101 : 4'b1001;
														assign node52198 = (inp[9]) ? 4'b1001 : 4'b1101;
													assign node52201 = (inp[12]) ? node52207 : node52202;
														assign node52202 = (inp[2]) ? node52204 : 4'b1111;
															assign node52204 = (inp[4]) ? 4'b1011 : 4'b1111;
														assign node52207 = (inp[4]) ? node52211 : node52208;
															assign node52208 = (inp[9]) ? 4'b1111 : 4'b1001;
															assign node52211 = (inp[9]) ? 4'b1011 : 4'b1111;
											assign node52214 = (inp[15]) ? node52234 : node52215;
												assign node52215 = (inp[5]) ? node52227 : node52216;
													assign node52216 = (inp[2]) ? node52222 : node52217;
														assign node52217 = (inp[12]) ? node52219 : 4'b1101;
															assign node52219 = (inp[4]) ? 4'b1101 : 4'b1001;
														assign node52222 = (inp[4]) ? 4'b1001 : node52223;
															assign node52223 = (inp[9]) ? 4'b1101 : 4'b1001;
													assign node52227 = (inp[9]) ? node52231 : node52228;
														assign node52228 = (inp[4]) ? 4'b1111 : 4'b1001;
														assign node52231 = (inp[4]) ? 4'b1011 : 4'b1111;
												assign node52234 = (inp[5]) ? node52242 : node52235;
													assign node52235 = (inp[4]) ? node52239 : node52236;
														assign node52236 = (inp[9]) ? 4'b1111 : 4'b1011;
														assign node52239 = (inp[9]) ? 4'b1011 : 4'b1111;
													assign node52242 = (inp[4]) ? node52246 : node52243;
														assign node52243 = (inp[9]) ? 4'b1101 : 4'b1011;
														assign node52246 = (inp[9]) ? 4'b1001 : 4'b1101;
										assign node52249 = (inp[2]) ? node52289 : node52250;
											assign node52250 = (inp[9]) ? node52274 : node52251;
												assign node52251 = (inp[4]) ? node52267 : node52252;
													assign node52252 = (inp[15]) ? node52260 : node52253;
														assign node52253 = (inp[0]) ? node52257 : node52254;
															assign node52254 = (inp[5]) ? 4'b1001 : 4'b1011;
															assign node52257 = (inp[5]) ? 4'b1011 : 4'b1001;
														assign node52260 = (inp[0]) ? node52264 : node52261;
															assign node52261 = (inp[5]) ? 4'b1011 : 4'b1001;
															assign node52264 = (inp[5]) ? 4'b1001 : 4'b1011;
													assign node52267 = (inp[0]) ? node52271 : node52268;
														assign node52268 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node52271 = (inp[15]) ? 4'b1101 : 4'b1111;
												assign node52274 = (inp[4]) ? node52282 : node52275;
													assign node52275 = (inp[15]) ? node52279 : node52276;
														assign node52276 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node52279 = (inp[0]) ? 4'b1101 : 4'b1111;
													assign node52282 = (inp[15]) ? node52286 : node52283;
														assign node52283 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node52286 = (inp[0]) ? 4'b1001 : 4'b1011;
											assign node52289 = (inp[15]) ? node52309 : node52290;
												assign node52290 = (inp[0]) ? node52300 : node52291;
													assign node52291 = (inp[4]) ? node52297 : node52292;
														assign node52292 = (inp[9]) ? 4'b1101 : node52293;
															assign node52293 = (inp[5]) ? 4'b1001 : 4'b1011;
														assign node52297 = (inp[9]) ? 4'b1001 : 4'b1101;
													assign node52300 = (inp[4]) ? node52306 : node52301;
														assign node52301 = (inp[9]) ? 4'b1111 : node52302;
															assign node52302 = (inp[5]) ? 4'b1011 : 4'b1001;
														assign node52306 = (inp[9]) ? 4'b1011 : 4'b1111;
												assign node52309 = (inp[0]) ? node52319 : node52310;
													assign node52310 = (inp[4]) ? node52316 : node52311;
														assign node52311 = (inp[9]) ? 4'b1111 : node52312;
															assign node52312 = (inp[5]) ? 4'b1011 : 4'b1001;
														assign node52316 = (inp[9]) ? 4'b1011 : 4'b1111;
													assign node52319 = (inp[9]) ? node52325 : node52320;
														assign node52320 = (inp[4]) ? 4'b1101 : node52321;
															assign node52321 = (inp[5]) ? 4'b1001 : 4'b1011;
														assign node52325 = (inp[4]) ? 4'b1001 : 4'b1101;
							assign node52328 = (inp[8]) ? node52724 : node52329;
								assign node52329 = (inp[2]) ? node52553 : node52330;
									assign node52330 = (inp[14]) ? node52448 : node52331;
										assign node52331 = (inp[4]) ? node52395 : node52332;
											assign node52332 = (inp[0]) ? node52354 : node52333;
												assign node52333 = (inp[15]) ? node52347 : node52334;
													assign node52334 = (inp[9]) ? node52342 : node52335;
														assign node52335 = (inp[12]) ? node52337 : 4'b0110;
															assign node52337 = (inp[3]) ? node52339 : 4'b0010;
																assign node52339 = (inp[5]) ? 4'b0000 : 4'b0010;
														assign node52342 = (inp[12]) ? 4'b0100 : node52343;
															assign node52343 = (inp[3]) ? 4'b0000 : 4'b0010;
													assign node52347 = (inp[9]) ? node52351 : node52348;
														assign node52348 = (inp[12]) ? 4'b0000 : 4'b0100;
														assign node52351 = (inp[12]) ? 4'b0110 : 4'b0000;
												assign node52354 = (inp[15]) ? node52376 : node52355;
													assign node52355 = (inp[3]) ? node52367 : node52356;
														assign node52356 = (inp[5]) ? node52362 : node52357;
															assign node52357 = (inp[12]) ? 4'b0100 : node52358;
																assign node52358 = (inp[9]) ? 4'b0000 : 4'b0100;
															assign node52362 = (inp[12]) ? 4'b0000 : node52363;
																assign node52363 = (inp[9]) ? 4'b0000 : 4'b0100;
														assign node52367 = (inp[5]) ? node52369 : 4'b0000;
															assign node52369 = (inp[9]) ? node52373 : node52370;
																assign node52370 = (inp[12]) ? 4'b0010 : 4'b0110;
																assign node52373 = (inp[12]) ? 4'b0110 : 4'b0010;
													assign node52376 = (inp[5]) ? node52382 : node52377;
														assign node52377 = (inp[3]) ? node52379 : 4'b0010;
															assign node52379 = (inp[12]) ? 4'b0010 : 4'b0110;
														assign node52382 = (inp[3]) ? node52390 : node52383;
															assign node52383 = (inp[9]) ? node52387 : node52384;
																assign node52384 = (inp[12]) ? 4'b0010 : 4'b0110;
																assign node52387 = (inp[12]) ? 4'b0100 : 4'b0010;
															assign node52390 = (inp[12]) ? node52392 : 4'b0000;
																assign node52392 = (inp[9]) ? 4'b0100 : 4'b0000;
											assign node52395 = (inp[9]) ? node52425 : node52396;
												assign node52396 = (inp[12]) ? node52408 : node52397;
													assign node52397 = (inp[0]) ? node52403 : node52398;
														assign node52398 = (inp[5]) ? 4'b0010 : node52399;
															assign node52399 = (inp[15]) ? 4'b0000 : 4'b0010;
														assign node52403 = (inp[15]) ? node52405 : 4'b0000;
															assign node52405 = (inp[5]) ? 4'b0000 : 4'b0010;
													assign node52408 = (inp[5]) ? node52418 : node52409;
														assign node52409 = (inp[15]) ? node52411 : 4'b0100;
															assign node52411 = (inp[0]) ? node52415 : node52412;
																assign node52412 = (inp[3]) ? 4'b0110 : 4'b0100;
																assign node52415 = (inp[3]) ? 4'b0100 : 4'b0110;
														assign node52418 = (inp[0]) ? node52422 : node52419;
															assign node52419 = (inp[3]) ? 4'b0110 : 4'b0100;
															assign node52422 = (inp[15]) ? 4'b0100 : 4'b0110;
												assign node52425 = (inp[12]) ? node52435 : node52426;
													assign node52426 = (inp[0]) ? node52428 : 4'b0110;
														assign node52428 = (inp[5]) ? 4'b0100 : node52429;
															assign node52429 = (inp[15]) ? node52431 : 4'b0110;
																assign node52431 = (inp[3]) ? 4'b0100 : 4'b0110;
													assign node52435 = (inp[3]) ? node52439 : node52436;
														assign node52436 = (inp[5]) ? 4'b0000 : 4'b0010;
														assign node52439 = (inp[5]) ? 4'b0010 : node52440;
															assign node52440 = (inp[15]) ? node52444 : node52441;
																assign node52441 = (inp[0]) ? 4'b0010 : 4'b0000;
																assign node52444 = (inp[0]) ? 4'b0000 : 4'b0010;
										assign node52448 = (inp[5]) ? node52500 : node52449;
											assign node52449 = (inp[3]) ? node52471 : node52450;
												assign node52450 = (inp[9]) ? node52462 : node52451;
													assign node52451 = (inp[4]) ? node52455 : node52452;
														assign node52452 = (inp[12]) ? 4'b1001 : 4'b1011;
														assign node52455 = (inp[15]) ? node52459 : node52456;
															assign node52456 = (inp[0]) ? 4'b1101 : 4'b1111;
															assign node52459 = (inp[0]) ? 4'b1111 : 4'b1101;
													assign node52462 = (inp[4]) ? node52468 : node52463;
														assign node52463 = (inp[15]) ? 4'b1101 : node52464;
															assign node52464 = (inp[0]) ? 4'b1101 : 4'b1111;
														assign node52468 = (inp[12]) ? 4'b1011 : 4'b1001;
												assign node52471 = (inp[0]) ? node52485 : node52472;
													assign node52472 = (inp[15]) ? node52480 : node52473;
														assign node52473 = (inp[12]) ? node52475 : 4'b1011;
															assign node52475 = (inp[4]) ? 4'b1101 : node52476;
																assign node52476 = (inp[9]) ? 4'b1101 : 4'b1011;
														assign node52480 = (inp[9]) ? node52482 : 4'b1111;
															assign node52482 = (inp[4]) ? 4'b1011 : 4'b1111;
													assign node52485 = (inp[15]) ? node52493 : node52486;
														assign node52486 = (inp[4]) ? node52490 : node52487;
															assign node52487 = (inp[9]) ? 4'b1111 : 4'b1001;
															assign node52490 = (inp[9]) ? 4'b1011 : 4'b1111;
														assign node52493 = (inp[9]) ? node52497 : node52494;
															assign node52494 = (inp[4]) ? 4'b1101 : 4'b1011;
															assign node52497 = (inp[4]) ? 4'b1001 : 4'b1101;
											assign node52500 = (inp[0]) ? node52526 : node52501;
												assign node52501 = (inp[15]) ? node52517 : node52502;
													assign node52502 = (inp[12]) ? node52512 : node52503;
														assign node52503 = (inp[4]) ? node52509 : node52504;
															assign node52504 = (inp[9]) ? 4'b1101 : node52505;
																assign node52505 = (inp[3]) ? 4'b1001 : 4'b1011;
															assign node52509 = (inp[9]) ? 4'b1001 : 4'b1101;
														assign node52512 = (inp[3]) ? 4'b1001 : node52513;
															assign node52513 = (inp[9]) ? 4'b1001 : 4'b1101;
													assign node52517 = (inp[9]) ? node52523 : node52518;
														assign node52518 = (inp[4]) ? 4'b1111 : node52519;
															assign node52519 = (inp[3]) ? 4'b1011 : 4'b1001;
														assign node52523 = (inp[4]) ? 4'b1011 : 4'b1111;
												assign node52526 = (inp[15]) ? node52544 : node52527;
													assign node52527 = (inp[12]) ? node52535 : node52528;
														assign node52528 = (inp[4]) ? node52532 : node52529;
															assign node52529 = (inp[3]) ? 4'b1011 : 4'b1001;
															assign node52532 = (inp[9]) ? 4'b1011 : 4'b1111;
														assign node52535 = (inp[3]) ? node52539 : node52536;
															assign node52536 = (inp[9]) ? 4'b1011 : 4'b1111;
															assign node52539 = (inp[4]) ? 4'b1011 : node52540;
																assign node52540 = (inp[9]) ? 4'b1111 : 4'b1011;
													assign node52544 = (inp[3]) ? node52548 : node52545;
														assign node52545 = (inp[4]) ? 4'b1001 : 4'b1011;
														assign node52548 = (inp[4]) ? node52550 : 4'b1001;
															assign node52550 = (inp[9]) ? 4'b1001 : 4'b1101;
									assign node52553 = (inp[4]) ? node52633 : node52554;
										assign node52554 = (inp[9]) ? node52578 : node52555;
											assign node52555 = (inp[3]) ? node52563 : node52556;
												assign node52556 = (inp[0]) ? node52560 : node52557;
													assign node52557 = (inp[15]) ? 4'b1001 : 4'b1011;
													assign node52560 = (inp[15]) ? 4'b1011 : 4'b1001;
												assign node52563 = (inp[15]) ? node52571 : node52564;
													assign node52564 = (inp[14]) ? node52566 : 4'b1011;
														assign node52566 = (inp[0]) ? 4'b1011 : node52567;
															assign node52567 = (inp[5]) ? 4'b1001 : 4'b1011;
													assign node52571 = (inp[0]) ? node52575 : node52572;
														assign node52572 = (inp[5]) ? 4'b1011 : 4'b1001;
														assign node52575 = (inp[5]) ? 4'b1001 : 4'b1011;
											assign node52578 = (inp[12]) ? node52600 : node52579;
												assign node52579 = (inp[14]) ? node52587 : node52580;
													assign node52580 = (inp[5]) ? node52582 : 4'b1111;
														assign node52582 = (inp[0]) ? node52584 : 4'b1111;
															assign node52584 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node52587 = (inp[3]) ? node52595 : node52588;
														assign node52588 = (inp[5]) ? 4'b1111 : node52589;
															assign node52589 = (inp[0]) ? 4'b1101 : node52590;
																assign node52590 = (inp[15]) ? 4'b1101 : 4'b1111;
														assign node52595 = (inp[0]) ? 4'b1101 : node52596;
															assign node52596 = (inp[15]) ? 4'b1111 : 4'b1101;
												assign node52600 = (inp[5]) ? node52620 : node52601;
													assign node52601 = (inp[3]) ? node52615 : node52602;
														assign node52602 = (inp[14]) ? node52610 : node52603;
															assign node52603 = (inp[0]) ? node52607 : node52604;
																assign node52604 = (inp[15]) ? 4'b1101 : 4'b1111;
																assign node52607 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node52610 = (inp[15]) ? node52612 : 4'b1101;
																assign node52612 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node52615 = (inp[15]) ? 4'b1111 : node52616;
															assign node52616 = (inp[0]) ? 4'b1111 : 4'b1101;
													assign node52620 = (inp[14]) ? node52626 : node52621;
														assign node52621 = (inp[15]) ? 4'b1101 : node52622;
															assign node52622 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node52626 = (inp[0]) ? node52630 : node52627;
															assign node52627 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node52630 = (inp[15]) ? 4'b1101 : 4'b1111;
										assign node52633 = (inp[9]) ? node52657 : node52634;
											assign node52634 = (inp[0]) ? node52646 : node52635;
												assign node52635 = (inp[15]) ? node52641 : node52636;
													assign node52636 = (inp[5]) ? 4'b1101 : node52637;
														assign node52637 = (inp[3]) ? 4'b1101 : 4'b1111;
													assign node52641 = (inp[5]) ? 4'b1111 : node52642;
														assign node52642 = (inp[3]) ? 4'b1111 : 4'b1101;
												assign node52646 = (inp[15]) ? node52652 : node52647;
													assign node52647 = (inp[5]) ? 4'b1111 : node52648;
														assign node52648 = (inp[3]) ? 4'b1111 : 4'b1101;
													assign node52652 = (inp[3]) ? 4'b1101 : node52653;
														assign node52653 = (inp[5]) ? 4'b1101 : 4'b1111;
											assign node52657 = (inp[14]) ? node52687 : node52658;
												assign node52658 = (inp[12]) ? node52672 : node52659;
													assign node52659 = (inp[15]) ? node52665 : node52660;
														assign node52660 = (inp[0]) ? 4'b1011 : node52661;
															assign node52661 = (inp[3]) ? 4'b1001 : 4'b1011;
														assign node52665 = (inp[3]) ? node52669 : node52666;
															assign node52666 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node52669 = (inp[0]) ? 4'b1001 : 4'b1011;
													assign node52672 = (inp[0]) ? node52678 : node52673;
														assign node52673 = (inp[3]) ? node52675 : 4'b1011;
															assign node52675 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node52678 = (inp[3]) ? 4'b1001 : node52679;
															assign node52679 = (inp[5]) ? node52683 : node52680;
																assign node52680 = (inp[15]) ? 4'b1011 : 4'b1001;
																assign node52683 = (inp[15]) ? 4'b1001 : 4'b1011;
												assign node52687 = (inp[5]) ? node52707 : node52688;
													assign node52688 = (inp[12]) ? node52698 : node52689;
														assign node52689 = (inp[3]) ? 4'b1001 : node52690;
															assign node52690 = (inp[15]) ? node52694 : node52691;
																assign node52691 = (inp[0]) ? 4'b1001 : 4'b1011;
																assign node52694 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node52698 = (inp[3]) ? node52700 : 4'b1001;
															assign node52700 = (inp[0]) ? node52704 : node52701;
																assign node52701 = (inp[15]) ? 4'b1011 : 4'b1001;
																assign node52704 = (inp[15]) ? 4'b1001 : 4'b1011;
													assign node52707 = (inp[3]) ? node52717 : node52708;
														assign node52708 = (inp[12]) ? node52712 : node52709;
															assign node52709 = (inp[15]) ? 4'b1011 : 4'b1001;
															assign node52712 = (inp[0]) ? node52714 : 4'b1001;
																assign node52714 = (inp[15]) ? 4'b1001 : 4'b1011;
														assign node52717 = (inp[0]) ? node52721 : node52718;
															assign node52718 = (inp[15]) ? 4'b1011 : 4'b1001;
															assign node52721 = (inp[15]) ? 4'b1001 : 4'b1011;
								assign node52724 = (inp[2]) ? node52974 : node52725;
									assign node52725 = (inp[14]) ? node52845 : node52726;
										assign node52726 = (inp[12]) ? node52780 : node52727;
											assign node52727 = (inp[9]) ? node52749 : node52728;
												assign node52728 = (inp[4]) ? node52740 : node52729;
													assign node52729 = (inp[0]) ? node52735 : node52730;
														assign node52730 = (inp[15]) ? node52732 : 4'b1011;
															assign node52732 = (inp[5]) ? 4'b1011 : 4'b1001;
														assign node52735 = (inp[15]) ? node52737 : 4'b1001;
															assign node52737 = (inp[5]) ? 4'b1001 : 4'b1011;
													assign node52740 = (inp[3]) ? 4'b1101 : node52741;
														assign node52741 = (inp[5]) ? node52743 : 4'b1111;
															assign node52743 = (inp[15]) ? node52745 : 4'b1111;
																assign node52745 = (inp[0]) ? 4'b1101 : 4'b1111;
												assign node52749 = (inp[4]) ? node52761 : node52750;
													assign node52750 = (inp[0]) ? node52756 : node52751;
														assign node52751 = (inp[3]) ? node52753 : 4'b1101;
															assign node52753 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node52756 = (inp[15]) ? node52758 : 4'b1111;
															assign node52758 = (inp[3]) ? 4'b1101 : 4'b1111;
													assign node52761 = (inp[3]) ? node52769 : node52762;
														assign node52762 = (inp[5]) ? 4'b1001 : node52763;
															assign node52763 = (inp[15]) ? node52765 : 4'b1001;
																assign node52765 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node52769 = (inp[5]) ? node52775 : node52770;
															assign node52770 = (inp[0]) ? node52772 : 4'b1011;
																assign node52772 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node52775 = (inp[0]) ? 4'b1001 : node52776;
																assign node52776 = (inp[15]) ? 4'b1011 : 4'b1001;
											assign node52780 = (inp[9]) ? node52816 : node52781;
												assign node52781 = (inp[4]) ? node52795 : node52782;
													assign node52782 = (inp[15]) ? node52792 : node52783;
														assign node52783 = (inp[3]) ? node52785 : 4'b1001;
															assign node52785 = (inp[5]) ? node52789 : node52786;
																assign node52786 = (inp[0]) ? 4'b1001 : 4'b1011;
																assign node52789 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node52792 = (inp[0]) ? 4'b1011 : 4'b1001;
													assign node52795 = (inp[5]) ? node52807 : node52796;
														assign node52796 = (inp[3]) ? node52802 : node52797;
															assign node52797 = (inp[15]) ? 4'b1101 : node52798;
																assign node52798 = (inp[0]) ? 4'b1101 : 4'b1111;
															assign node52802 = (inp[15]) ? 4'b1111 : node52803;
																assign node52803 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node52807 = (inp[3]) ? 4'b1101 : node52808;
															assign node52808 = (inp[0]) ? node52812 : node52809;
																assign node52809 = (inp[15]) ? 4'b1111 : 4'b1101;
																assign node52812 = (inp[15]) ? 4'b1101 : 4'b1111;
												assign node52816 = (inp[4]) ? node52834 : node52817;
													assign node52817 = (inp[0]) ? node52825 : node52818;
														assign node52818 = (inp[15]) ? 4'b1111 : node52819;
															assign node52819 = (inp[3]) ? 4'b1101 : node52820;
																assign node52820 = (inp[5]) ? 4'b1101 : 4'b1111;
														assign node52825 = (inp[5]) ? 4'b1101 : node52826;
															assign node52826 = (inp[15]) ? node52830 : node52827;
																assign node52827 = (inp[3]) ? 4'b1111 : 4'b1101;
																assign node52830 = (inp[3]) ? 4'b1101 : 4'b1111;
													assign node52834 = (inp[0]) ? node52842 : node52835;
														assign node52835 = (inp[15]) ? node52839 : node52836;
															assign node52836 = (inp[3]) ? 4'b1001 : 4'b1011;
															assign node52839 = (inp[5]) ? 4'b1011 : 4'b1001;
														assign node52842 = (inp[15]) ? 4'b1001 : 4'b1011;
										assign node52845 = (inp[12]) ? node52909 : node52846;
											assign node52846 = (inp[4]) ? node52876 : node52847;
												assign node52847 = (inp[9]) ? node52861 : node52848;
													assign node52848 = (inp[5]) ? node52854 : node52849;
														assign node52849 = (inp[15]) ? 4'b1000 : node52850;
															assign node52850 = (inp[0]) ? 4'b1000 : 4'b1010;
														assign node52854 = (inp[15]) ? node52858 : node52855;
															assign node52855 = (inp[3]) ? 4'b1010 : 4'b1000;
															assign node52858 = (inp[3]) ? 4'b1000 : 4'b1010;
													assign node52861 = (inp[15]) ? node52867 : node52862;
														assign node52862 = (inp[0]) ? 4'b1110 : node52863;
															assign node52863 = (inp[3]) ? 4'b1100 : 4'b1110;
														assign node52867 = (inp[0]) ? node52871 : node52868;
															assign node52868 = (inp[5]) ? 4'b1110 : 4'b1100;
															assign node52871 = (inp[5]) ? 4'b1100 : node52872;
																assign node52872 = (inp[3]) ? 4'b1100 : 4'b1110;
												assign node52876 = (inp[9]) ? node52896 : node52877;
													assign node52877 = (inp[0]) ? node52887 : node52878;
														assign node52878 = (inp[3]) ? 4'b1110 : node52879;
															assign node52879 = (inp[15]) ? node52883 : node52880;
																assign node52880 = (inp[5]) ? 4'b1100 : 4'b1110;
																assign node52883 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node52887 = (inp[15]) ? node52893 : node52888;
															assign node52888 = (inp[3]) ? 4'b1110 : node52889;
																assign node52889 = (inp[5]) ? 4'b1110 : 4'b1100;
															assign node52893 = (inp[3]) ? 4'b1100 : 4'b1110;
													assign node52896 = (inp[5]) ? node52904 : node52897;
														assign node52897 = (inp[3]) ? 4'b1010 : node52898;
															assign node52898 = (inp[0]) ? node52900 : 4'b1010;
																assign node52900 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node52904 = (inp[0]) ? 4'b1000 : node52905;
															assign node52905 = (inp[15]) ? 4'b1010 : 4'b1000;
											assign node52909 = (inp[0]) ? node52937 : node52910;
												assign node52910 = (inp[4]) ? node52924 : node52911;
													assign node52911 = (inp[9]) ? node52917 : node52912;
														assign node52912 = (inp[15]) ? 4'b1000 : node52913;
															assign node52913 = (inp[3]) ? 4'b1000 : 4'b1010;
														assign node52917 = (inp[3]) ? 4'b1100 : node52918;
															assign node52918 = (inp[15]) ? 4'b1100 : node52919;
																assign node52919 = (inp[5]) ? 4'b1100 : 4'b1110;
													assign node52924 = (inp[9]) ? node52928 : node52925;
														assign node52925 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node52928 = (inp[15]) ? node52934 : node52929;
															assign node52929 = (inp[3]) ? 4'b1000 : node52930;
																assign node52930 = (inp[5]) ? 4'b1000 : 4'b1010;
															assign node52934 = (inp[3]) ? 4'b1010 : 4'b1000;
												assign node52937 = (inp[15]) ? node52953 : node52938;
													assign node52938 = (inp[5]) ? node52946 : node52939;
														assign node52939 = (inp[4]) ? node52943 : node52940;
															assign node52940 = (inp[9]) ? 4'b1110 : 4'b1000;
															assign node52943 = (inp[9]) ? 4'b1000 : 4'b1100;
														assign node52946 = (inp[9]) ? node52950 : node52947;
															assign node52947 = (inp[4]) ? 4'b1110 : 4'b1010;
															assign node52950 = (inp[4]) ? 4'b1010 : 4'b1110;
													assign node52953 = (inp[5]) ? node52965 : node52954;
														assign node52954 = (inp[3]) ? node52960 : node52955;
															assign node52955 = (inp[4]) ? node52957 : 4'b1110;
																assign node52957 = (inp[9]) ? 4'b1010 : 4'b1110;
															assign node52960 = (inp[4]) ? node52962 : 4'b1010;
																assign node52962 = (inp[9]) ? 4'b1000 : 4'b1100;
														assign node52965 = (inp[4]) ? node52971 : node52966;
															assign node52966 = (inp[9]) ? 4'b1100 : node52967;
																assign node52967 = (inp[3]) ? 4'b1000 : 4'b1010;
															assign node52971 = (inp[9]) ? 4'b1000 : 4'b1100;
									assign node52974 = (inp[4]) ? node53080 : node52975;
										assign node52975 = (inp[9]) ? node53013 : node52976;
											assign node52976 = (inp[14]) ? node52996 : node52977;
												assign node52977 = (inp[0]) ? node52987 : node52978;
													assign node52978 = (inp[15]) ? node52982 : node52979;
														assign node52979 = (inp[3]) ? 4'b1000 : 4'b1010;
														assign node52982 = (inp[3]) ? node52984 : 4'b1000;
															assign node52984 = (inp[5]) ? 4'b1010 : 4'b1000;
													assign node52987 = (inp[15]) ? node52991 : node52988;
														assign node52988 = (inp[5]) ? 4'b1010 : 4'b1000;
														assign node52991 = (inp[5]) ? node52993 : 4'b1010;
															assign node52993 = (inp[3]) ? 4'b1000 : 4'b1010;
												assign node52996 = (inp[15]) ? node53004 : node52997;
													assign node52997 = (inp[0]) ? node52999 : 4'b1010;
														assign node52999 = (inp[5]) ? node53001 : 4'b1000;
															assign node53001 = (inp[3]) ? 4'b1010 : 4'b1000;
													assign node53004 = (inp[0]) ? node53010 : node53005;
														assign node53005 = (inp[3]) ? node53007 : 4'b1000;
															assign node53007 = (inp[5]) ? 4'b1010 : 4'b1000;
														assign node53010 = (inp[5]) ? 4'b1000 : 4'b1010;
											assign node53013 = (inp[5]) ? node53051 : node53014;
												assign node53014 = (inp[12]) ? node53034 : node53015;
													assign node53015 = (inp[3]) ? node53021 : node53016;
														assign node53016 = (inp[15]) ? 4'b1110 : node53017;
															assign node53017 = (inp[0]) ? 4'b1100 : 4'b1110;
														assign node53021 = (inp[14]) ? node53029 : node53022;
															assign node53022 = (inp[0]) ? node53026 : node53023;
																assign node53023 = (inp[15]) ? 4'b1110 : 4'b1100;
																assign node53026 = (inp[15]) ? 4'b1100 : 4'b1110;
															assign node53029 = (inp[0]) ? node53031 : 4'b1100;
																assign node53031 = (inp[15]) ? 4'b1100 : 4'b1110;
													assign node53034 = (inp[15]) ? node53044 : node53035;
														assign node53035 = (inp[14]) ? node53037 : 4'b1100;
															assign node53037 = (inp[0]) ? node53041 : node53038;
																assign node53038 = (inp[3]) ? 4'b1100 : 4'b1110;
																assign node53041 = (inp[3]) ? 4'b1110 : 4'b1100;
														assign node53044 = (inp[14]) ? 4'b1100 : node53045;
															assign node53045 = (inp[3]) ? node53047 : 4'b1100;
																assign node53047 = (inp[0]) ? 4'b1100 : 4'b1110;
												assign node53051 = (inp[3]) ? node53065 : node53052;
													assign node53052 = (inp[12]) ? node53060 : node53053;
														assign node53053 = (inp[14]) ? 4'b1100 : node53054;
															assign node53054 = (inp[15]) ? 4'b1100 : node53055;
																assign node53055 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node53060 = (inp[0]) ? 4'b1110 : node53061;
															assign node53061 = (inp[15]) ? 4'b1110 : 4'b1100;
													assign node53065 = (inp[14]) ? node53073 : node53066;
														assign node53066 = (inp[0]) ? node53070 : node53067;
															assign node53067 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node53070 = (inp[15]) ? 4'b1100 : 4'b1110;
														assign node53073 = (inp[15]) ? node53077 : node53074;
															assign node53074 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node53077 = (inp[0]) ? 4'b1100 : 4'b1110;
										assign node53080 = (inp[9]) ? node53120 : node53081;
											assign node53081 = (inp[5]) ? node53109 : node53082;
												assign node53082 = (inp[15]) ? node53094 : node53083;
													assign node53083 = (inp[14]) ? node53089 : node53084;
														assign node53084 = (inp[0]) ? node53086 : 4'b1100;
															assign node53086 = (inp[3]) ? 4'b1110 : 4'b1100;
														assign node53089 = (inp[0]) ? 4'b1100 : node53090;
															assign node53090 = (inp[3]) ? 4'b1100 : 4'b1110;
													assign node53094 = (inp[14]) ? node53102 : node53095;
														assign node53095 = (inp[3]) ? node53099 : node53096;
															assign node53096 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node53099 = (inp[0]) ? 4'b1100 : 4'b1110;
														assign node53102 = (inp[0]) ? node53106 : node53103;
															assign node53103 = (inp[3]) ? 4'b1110 : 4'b1100;
															assign node53106 = (inp[3]) ? 4'b1100 : 4'b1110;
												assign node53109 = (inp[12]) ? node53115 : node53110;
													assign node53110 = (inp[0]) ? 4'b1110 : node53111;
														assign node53111 = (inp[15]) ? 4'b1110 : 4'b1100;
													assign node53115 = (inp[15]) ? node53117 : 4'b1110;
														assign node53117 = (inp[0]) ? 4'b1100 : 4'b1110;
											assign node53120 = (inp[12]) ? node53152 : node53121;
												assign node53121 = (inp[5]) ? node53145 : node53122;
													assign node53122 = (inp[0]) ? node53130 : node53123;
														assign node53123 = (inp[15]) ? node53127 : node53124;
															assign node53124 = (inp[3]) ? 4'b1000 : 4'b1010;
															assign node53127 = (inp[3]) ? 4'b1010 : 4'b1000;
														assign node53130 = (inp[14]) ? node53138 : node53131;
															assign node53131 = (inp[15]) ? node53135 : node53132;
																assign node53132 = (inp[3]) ? 4'b1010 : 4'b1000;
																assign node53135 = (inp[3]) ? 4'b1000 : 4'b1010;
															assign node53138 = (inp[15]) ? node53142 : node53139;
																assign node53139 = (inp[3]) ? 4'b1010 : 4'b1000;
																assign node53142 = (inp[3]) ? 4'b1000 : 4'b1010;
													assign node53145 = (inp[15]) ? node53149 : node53146;
														assign node53146 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node53149 = (inp[0]) ? 4'b1000 : 4'b1010;
												assign node53152 = (inp[3]) ? node53172 : node53153;
													assign node53153 = (inp[14]) ? node53163 : node53154;
														assign node53154 = (inp[15]) ? node53156 : 4'b1010;
															assign node53156 = (inp[5]) ? node53160 : node53157;
																assign node53157 = (inp[0]) ? 4'b1010 : 4'b1000;
																assign node53160 = (inp[0]) ? 4'b1000 : 4'b1010;
														assign node53163 = (inp[15]) ? 4'b1010 : node53164;
															assign node53164 = (inp[5]) ? node53168 : node53165;
																assign node53165 = (inp[0]) ? 4'b1000 : 4'b1010;
																assign node53168 = (inp[0]) ? 4'b1010 : 4'b1000;
													assign node53172 = (inp[15]) ? node53176 : node53173;
														assign node53173 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node53176 = (inp[0]) ? 4'b1000 : 4'b1010;
						assign node53179 = (inp[9]) ? node53977 : node53180;
							assign node53180 = (inp[4]) ? node53640 : node53181;
								assign node53181 = (inp[5]) ? node53409 : node53182;
									assign node53182 = (inp[12]) ? node53276 : node53183;
										assign node53183 = (inp[15]) ? node53217 : node53184;
											assign node53184 = (inp[0]) ? node53200 : node53185;
												assign node53185 = (inp[7]) ? node53195 : node53186;
													assign node53186 = (inp[8]) ? node53190 : node53187;
														assign node53187 = (inp[14]) ? 4'b1010 : 4'b1011;
														assign node53190 = (inp[14]) ? 4'b1011 : node53191;
															assign node53191 = (inp[2]) ? 4'b1011 : 4'b1010;
													assign node53195 = (inp[3]) ? 4'b1010 : node53196;
														assign node53196 = (inp[14]) ? 4'b1010 : 4'b1011;
												assign node53200 = (inp[2]) ? node53210 : node53201;
													assign node53201 = (inp[14]) ? node53203 : 4'b1001;
														assign node53203 = (inp[7]) ? node53207 : node53204;
															assign node53204 = (inp[8]) ? 4'b1001 : 4'b1000;
															assign node53207 = (inp[8]) ? 4'b1000 : 4'b1001;
													assign node53210 = (inp[8]) ? node53214 : node53211;
														assign node53211 = (inp[7]) ? 4'b1001 : 4'b1000;
														assign node53214 = (inp[7]) ? 4'b1000 : 4'b1001;
											assign node53217 = (inp[0]) ? node53239 : node53218;
												assign node53218 = (inp[8]) ? node53230 : node53219;
													assign node53219 = (inp[2]) ? 4'b1000 : node53220;
														assign node53220 = (inp[3]) ? node53226 : node53221;
															assign node53221 = (inp[14]) ? 4'b1000 : node53222;
																assign node53222 = (inp[7]) ? 4'b1000 : 4'b1001;
															assign node53226 = (inp[14]) ? 4'b1001 : 4'b1000;
													assign node53230 = (inp[7]) ? node53236 : node53231;
														assign node53231 = (inp[2]) ? 4'b1001 : node53232;
															assign node53232 = (inp[14]) ? 4'b1001 : 4'b1000;
														assign node53236 = (inp[14]) ? 4'b1000 : 4'b1001;
												assign node53239 = (inp[2]) ? node53261 : node53240;
													assign node53240 = (inp[3]) ? node53246 : node53241;
														assign node53241 = (inp[8]) ? 4'b1010 : node53242;
															assign node53242 = (inp[14]) ? 4'b1011 : 4'b1010;
														assign node53246 = (inp[8]) ? node53254 : node53247;
															assign node53247 = (inp[14]) ? node53251 : node53248;
																assign node53248 = (inp[7]) ? 4'b1010 : 4'b1011;
																assign node53251 = (inp[7]) ? 4'b1011 : 4'b1010;
															assign node53254 = (inp[7]) ? node53258 : node53255;
																assign node53255 = (inp[14]) ? 4'b1011 : 4'b1010;
																assign node53258 = (inp[14]) ? 4'b1010 : 4'b1011;
													assign node53261 = (inp[14]) ? node53269 : node53262;
														assign node53262 = (inp[8]) ? node53266 : node53263;
															assign node53263 = (inp[7]) ? 4'b1011 : 4'b1010;
															assign node53266 = (inp[7]) ? 4'b1010 : 4'b1011;
														assign node53269 = (inp[7]) ? node53273 : node53270;
															assign node53270 = (inp[8]) ? 4'b1011 : 4'b1010;
															assign node53273 = (inp[8]) ? 4'b1010 : 4'b1011;
										assign node53276 = (inp[14]) ? node53344 : node53277;
											assign node53277 = (inp[8]) ? node53317 : node53278;
												assign node53278 = (inp[2]) ? node53304 : node53279;
													assign node53279 = (inp[7]) ? node53295 : node53280;
														assign node53280 = (inp[3]) ? node53288 : node53281;
															assign node53281 = (inp[15]) ? node53285 : node53282;
																assign node53282 = (inp[0]) ? 4'b1001 : 4'b1011;
																assign node53285 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node53288 = (inp[15]) ? node53292 : node53289;
																assign node53289 = (inp[0]) ? 4'b1001 : 4'b1011;
																assign node53292 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node53295 = (inp[3]) ? node53301 : node53296;
															assign node53296 = (inp[15]) ? node53298 : 4'b1010;
																assign node53298 = (inp[0]) ? 4'b1010 : 4'b1000;
															assign node53301 = (inp[0]) ? 4'b1000 : 4'b1010;
													assign node53304 = (inp[7]) ? node53312 : node53305;
														assign node53305 = (inp[15]) ? node53309 : node53306;
															assign node53306 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node53309 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node53312 = (inp[15]) ? 4'b1001 : node53313;
															assign node53313 = (inp[3]) ? 4'b1001 : 4'b1011;
												assign node53317 = (inp[2]) ? node53329 : node53318;
													assign node53318 = (inp[7]) ? node53326 : node53319;
														assign node53319 = (inp[15]) ? node53323 : node53320;
															assign node53320 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node53323 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node53326 = (inp[3]) ? 4'b1001 : 4'b1011;
													assign node53329 = (inp[7]) ? node53339 : node53330;
														assign node53330 = (inp[3]) ? node53332 : 4'b1001;
															assign node53332 = (inp[15]) ? node53336 : node53333;
																assign node53333 = (inp[0]) ? 4'b1001 : 4'b1011;
																assign node53336 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node53339 = (inp[15]) ? node53341 : 4'b1000;
															assign node53341 = (inp[0]) ? 4'b1010 : 4'b1000;
											assign node53344 = (inp[3]) ? node53378 : node53345;
												assign node53345 = (inp[15]) ? node53367 : node53346;
													assign node53346 = (inp[0]) ? node53354 : node53347;
														assign node53347 = (inp[2]) ? 4'b1010 : node53348;
															assign node53348 = (inp[7]) ? node53350 : 4'b1011;
																assign node53350 = (inp[8]) ? 4'b1010 : 4'b1011;
														assign node53354 = (inp[2]) ? node53360 : node53355;
															assign node53355 = (inp[8]) ? 4'b1001 : node53356;
																assign node53356 = (inp[7]) ? 4'b1001 : 4'b1000;
															assign node53360 = (inp[8]) ? node53364 : node53361;
																assign node53361 = (inp[7]) ? 4'b1001 : 4'b1000;
																assign node53364 = (inp[7]) ? 4'b1000 : 4'b1001;
													assign node53367 = (inp[0]) ? node53373 : node53368;
														assign node53368 = (inp[7]) ? 4'b1001 : node53369;
															assign node53369 = (inp[8]) ? 4'b1001 : 4'b1000;
														assign node53373 = (inp[8]) ? node53375 : 4'b1011;
															assign node53375 = (inp[7]) ? 4'b1010 : 4'b1011;
												assign node53378 = (inp[8]) ? node53398 : node53379;
													assign node53379 = (inp[7]) ? node53391 : node53380;
														assign node53380 = (inp[2]) ? node53386 : node53381;
															assign node53381 = (inp[15]) ? 4'b1010 : node53382;
																assign node53382 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node53386 = (inp[0]) ? node53388 : 4'b1000;
																assign node53388 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node53391 = (inp[0]) ? node53395 : node53392;
															assign node53392 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node53395 = (inp[15]) ? 4'b1011 : 4'b1001;
													assign node53398 = (inp[7]) ? node53406 : node53399;
														assign node53399 = (inp[15]) ? node53403 : node53400;
															assign node53400 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node53403 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node53406 = (inp[15]) ? 4'b1000 : 4'b1010;
									assign node53409 = (inp[2]) ? node53531 : node53410;
										assign node53410 = (inp[7]) ? node53478 : node53411;
											assign node53411 = (inp[8]) ? node53443 : node53412;
												assign node53412 = (inp[14]) ? node53432 : node53413;
													assign node53413 = (inp[3]) ? node53427 : node53414;
														assign node53414 = (inp[12]) ? node53420 : node53415;
															assign node53415 = (inp[0]) ? 4'b1011 : node53416;
																assign node53416 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node53420 = (inp[15]) ? node53424 : node53421;
																assign node53421 = (inp[0]) ? 4'b1001 : 4'b1011;
																assign node53424 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node53427 = (inp[15]) ? 4'b1011 : node53428;
															assign node53428 = (inp[0]) ? 4'b1011 : 4'b1001;
													assign node53432 = (inp[0]) ? node53438 : node53433;
														assign node53433 = (inp[3]) ? node53435 : 4'b1010;
															assign node53435 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node53438 = (inp[3]) ? node53440 : 4'b1000;
															assign node53440 = (inp[15]) ? 4'b1000 : 4'b1010;
												assign node53443 = (inp[14]) ? node53467 : node53444;
													assign node53444 = (inp[12]) ? node53458 : node53445;
														assign node53445 = (inp[0]) ? node53453 : node53446;
															assign node53446 = (inp[15]) ? node53450 : node53447;
																assign node53447 = (inp[3]) ? 4'b1000 : 4'b1010;
																assign node53450 = (inp[3]) ? 4'b1010 : 4'b1000;
															assign node53453 = (inp[3]) ? 4'b1000 : node53454;
																assign node53454 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node53458 = (inp[15]) ? node53460 : 4'b1010;
															assign node53460 = (inp[0]) ? node53464 : node53461;
																assign node53461 = (inp[3]) ? 4'b1010 : 4'b1000;
																assign node53464 = (inp[3]) ? 4'b1000 : 4'b1010;
													assign node53467 = (inp[12]) ? node53473 : node53468;
														assign node53468 = (inp[3]) ? node53470 : 4'b1001;
															assign node53470 = (inp[15]) ? 4'b1001 : 4'b1011;
														assign node53473 = (inp[3]) ? 4'b1011 : node53474;
															assign node53474 = (inp[15]) ? 4'b1001 : 4'b1011;
											assign node53478 = (inp[3]) ? node53512 : node53479;
												assign node53479 = (inp[14]) ? node53493 : node53480;
													assign node53480 = (inp[8]) ? node53486 : node53481;
														assign node53481 = (inp[0]) ? node53483 : 4'b1010;
															assign node53483 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node53486 = (inp[12]) ? 4'b1001 : node53487;
															assign node53487 = (inp[15]) ? 4'b1001 : node53488;
																assign node53488 = (inp[0]) ? 4'b1001 : 4'b1011;
													assign node53493 = (inp[8]) ? node53507 : node53494;
														assign node53494 = (inp[12]) ? node53502 : node53495;
															assign node53495 = (inp[0]) ? node53499 : node53496;
																assign node53496 = (inp[15]) ? 4'b1001 : 4'b1011;
																assign node53499 = (inp[15]) ? 4'b1011 : 4'b1001;
															assign node53502 = (inp[0]) ? node53504 : 4'b1011;
																assign node53504 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node53507 = (inp[15]) ? node53509 : 4'b1010;
															assign node53509 = (inp[0]) ? 4'b1010 : 4'b1000;
												assign node53512 = (inp[14]) ? node53524 : node53513;
													assign node53513 = (inp[8]) ? node53517 : node53514;
														assign node53514 = (inp[15]) ? 4'b1000 : 4'b1010;
														assign node53517 = (inp[0]) ? node53521 : node53518;
															assign node53518 = (inp[15]) ? 4'b1011 : 4'b1001;
															assign node53521 = (inp[12]) ? 4'b1001 : 4'b1011;
													assign node53524 = (inp[8]) ? node53526 : 4'b1001;
														assign node53526 = (inp[15]) ? node53528 : 4'b1000;
															assign node53528 = (inp[0]) ? 4'b1000 : 4'b1010;
										assign node53531 = (inp[12]) ? node53585 : node53532;
											assign node53532 = (inp[8]) ? node53558 : node53533;
												assign node53533 = (inp[7]) ? node53543 : node53534;
													assign node53534 = (inp[0]) ? node53536 : 4'b1010;
														assign node53536 = (inp[3]) ? node53540 : node53537;
															assign node53537 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node53540 = (inp[15]) ? 4'b1000 : 4'b1010;
													assign node53543 = (inp[15]) ? node53549 : node53544;
														assign node53544 = (inp[0]) ? 4'b1011 : node53545;
															assign node53545 = (inp[3]) ? 4'b1001 : 4'b1011;
														assign node53549 = (inp[14]) ? node53553 : node53550;
															assign node53550 = (inp[3]) ? 4'b1011 : 4'b1001;
															assign node53553 = (inp[3]) ? node53555 : 4'b1011;
																assign node53555 = (inp[0]) ? 4'b1001 : 4'b1011;
												assign node53558 = (inp[7]) ? node53580 : node53559;
													assign node53559 = (inp[3]) ? node53567 : node53560;
														assign node53560 = (inp[0]) ? node53564 : node53561;
															assign node53561 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node53564 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node53567 = (inp[14]) ? node53575 : node53568;
															assign node53568 = (inp[0]) ? node53572 : node53569;
																assign node53569 = (inp[15]) ? 4'b1011 : 4'b1001;
																assign node53572 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node53575 = (inp[15]) ? 4'b1011 : node53576;
																assign node53576 = (inp[0]) ? 4'b1011 : 4'b1001;
													assign node53580 = (inp[0]) ? node53582 : 4'b1010;
														assign node53582 = (inp[3]) ? 4'b1010 : 4'b1000;
											assign node53585 = (inp[7]) ? node53617 : node53586;
												assign node53586 = (inp[8]) ? node53602 : node53587;
													assign node53587 = (inp[15]) ? node53595 : node53588;
														assign node53588 = (inp[14]) ? node53590 : 4'b1000;
															assign node53590 = (inp[3]) ? node53592 : 4'b1000;
																assign node53592 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node53595 = (inp[3]) ? node53599 : node53596;
															assign node53596 = (inp[14]) ? 4'b1000 : 4'b1010;
															assign node53599 = (inp[14]) ? 4'b1010 : 4'b1000;
													assign node53602 = (inp[3]) ? node53610 : node53603;
														assign node53603 = (inp[15]) ? node53607 : node53604;
															assign node53604 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node53607 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node53610 = (inp[14]) ? 4'b1011 : node53611;
															assign node53611 = (inp[0]) ? node53613 : 4'b1011;
																assign node53613 = (inp[15]) ? 4'b1001 : 4'b1011;
												assign node53617 = (inp[8]) ? node53629 : node53618;
													assign node53618 = (inp[14]) ? node53620 : 4'b1011;
														assign node53620 = (inp[0]) ? 4'b1011 : node53621;
															assign node53621 = (inp[15]) ? node53625 : node53622;
																assign node53622 = (inp[3]) ? 4'b1001 : 4'b1011;
																assign node53625 = (inp[3]) ? 4'b1011 : 4'b1001;
													assign node53629 = (inp[0]) ? node53633 : node53630;
														assign node53630 = (inp[14]) ? 4'b1010 : 4'b1000;
														assign node53633 = (inp[3]) ? node53637 : node53634;
															assign node53634 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node53637 = (inp[15]) ? 4'b1000 : 4'b1010;
								assign node53640 = (inp[8]) ? node53784 : node53641;
									assign node53641 = (inp[7]) ? node53715 : node53642;
										assign node53642 = (inp[2]) ? node53688 : node53643;
											assign node53643 = (inp[14]) ? node53667 : node53644;
												assign node53644 = (inp[0]) ? node53656 : node53645;
													assign node53645 = (inp[15]) ? node53651 : node53646;
														assign node53646 = (inp[12]) ? 4'b1101 : node53647;
															assign node53647 = (inp[5]) ? 4'b1101 : 4'b1111;
														assign node53651 = (inp[5]) ? 4'b1111 : node53652;
															assign node53652 = (inp[3]) ? 4'b1111 : 4'b1101;
													assign node53656 = (inp[15]) ? node53662 : node53657;
														assign node53657 = (inp[3]) ? 4'b1111 : node53658;
															assign node53658 = (inp[5]) ? 4'b1111 : 4'b1101;
														assign node53662 = (inp[3]) ? 4'b1101 : node53663;
															assign node53663 = (inp[5]) ? 4'b1101 : 4'b1111;
												assign node53667 = (inp[5]) ? node53681 : node53668;
													assign node53668 = (inp[15]) ? node53676 : node53669;
														assign node53669 = (inp[12]) ? 4'b1100 : node53670;
															assign node53670 = (inp[3]) ? 4'b1110 : node53671;
																assign node53671 = (inp[0]) ? 4'b1100 : 4'b1110;
														assign node53676 = (inp[0]) ? node53678 : 4'b1100;
															assign node53678 = (inp[3]) ? 4'b1100 : 4'b1110;
													assign node53681 = (inp[0]) ? node53685 : node53682;
														assign node53682 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node53685 = (inp[15]) ? 4'b1100 : 4'b1110;
											assign node53688 = (inp[3]) ? node53708 : node53689;
												assign node53689 = (inp[15]) ? node53701 : node53690;
													assign node53690 = (inp[14]) ? node53696 : node53691;
														assign node53691 = (inp[5]) ? node53693 : 4'b1110;
															assign node53693 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node53696 = (inp[12]) ? node53698 : 4'b1110;
															assign node53698 = (inp[0]) ? 4'b1100 : 4'b1110;
													assign node53701 = (inp[0]) ? node53705 : node53702;
														assign node53702 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node53705 = (inp[5]) ? 4'b1100 : 4'b1110;
												assign node53708 = (inp[0]) ? node53712 : node53709;
													assign node53709 = (inp[15]) ? 4'b1110 : 4'b1100;
													assign node53712 = (inp[15]) ? 4'b1100 : 4'b1110;
										assign node53715 = (inp[14]) ? node53761 : node53716;
											assign node53716 = (inp[2]) ? node53738 : node53717;
												assign node53717 = (inp[0]) ? node53727 : node53718;
													assign node53718 = (inp[15]) ? node53722 : node53719;
														assign node53719 = (inp[5]) ? 4'b1100 : 4'b1110;
														assign node53722 = (inp[5]) ? 4'b1110 : node53723;
															assign node53723 = (inp[3]) ? 4'b1110 : 4'b1100;
													assign node53727 = (inp[15]) ? node53733 : node53728;
														assign node53728 = (inp[5]) ? 4'b1110 : node53729;
															assign node53729 = (inp[3]) ? 4'b1110 : 4'b1100;
														assign node53733 = (inp[3]) ? 4'b1100 : node53734;
															assign node53734 = (inp[5]) ? 4'b1100 : 4'b1110;
												assign node53738 = (inp[3]) ? node53754 : node53739;
													assign node53739 = (inp[5]) ? node53749 : node53740;
														assign node53740 = (inp[12]) ? 4'b1111 : node53741;
															assign node53741 = (inp[0]) ? node53745 : node53742;
																assign node53742 = (inp[15]) ? 4'b1101 : 4'b1111;
																assign node53745 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node53749 = (inp[15]) ? 4'b1111 : node53750;
															assign node53750 = (inp[0]) ? 4'b1111 : 4'b1101;
													assign node53754 = (inp[0]) ? node53758 : node53755;
														assign node53755 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node53758 = (inp[15]) ? 4'b1101 : 4'b1111;
											assign node53761 = (inp[0]) ? node53773 : node53762;
												assign node53762 = (inp[15]) ? node53768 : node53763;
													assign node53763 = (inp[5]) ? 4'b1101 : node53764;
														assign node53764 = (inp[3]) ? 4'b1101 : 4'b1111;
													assign node53768 = (inp[5]) ? 4'b1111 : node53769;
														assign node53769 = (inp[3]) ? 4'b1111 : 4'b1101;
												assign node53773 = (inp[15]) ? node53779 : node53774;
													assign node53774 = (inp[3]) ? 4'b1111 : node53775;
														assign node53775 = (inp[5]) ? 4'b1111 : 4'b1101;
													assign node53779 = (inp[3]) ? 4'b1101 : node53780;
														assign node53780 = (inp[5]) ? 4'b1101 : 4'b1111;
									assign node53784 = (inp[7]) ? node53886 : node53785;
										assign node53785 = (inp[14]) ? node53859 : node53786;
											assign node53786 = (inp[2]) ? node53824 : node53787;
												assign node53787 = (inp[12]) ? node53805 : node53788;
													assign node53788 = (inp[0]) ? node53794 : node53789;
														assign node53789 = (inp[15]) ? node53791 : 4'b1100;
															assign node53791 = (inp[3]) ? 4'b1110 : 4'b1100;
														assign node53794 = (inp[15]) ? node53800 : node53795;
															assign node53795 = (inp[3]) ? 4'b1110 : node53796;
																assign node53796 = (inp[5]) ? 4'b1110 : 4'b1100;
															assign node53800 = (inp[5]) ? 4'b1100 : node53801;
																assign node53801 = (inp[3]) ? 4'b1100 : 4'b1110;
													assign node53805 = (inp[3]) ? node53819 : node53806;
														assign node53806 = (inp[15]) ? node53814 : node53807;
															assign node53807 = (inp[0]) ? node53811 : node53808;
																assign node53808 = (inp[5]) ? 4'b1100 : 4'b1110;
																assign node53811 = (inp[5]) ? 4'b1110 : 4'b1100;
															assign node53814 = (inp[0]) ? node53816 : 4'b1110;
																assign node53816 = (inp[5]) ? 4'b1100 : 4'b1110;
														assign node53819 = (inp[0]) ? node53821 : 4'b1110;
															assign node53821 = (inp[15]) ? 4'b1100 : 4'b1110;
												assign node53824 = (inp[5]) ? node53838 : node53825;
													assign node53825 = (inp[12]) ? node53831 : node53826;
														assign node53826 = (inp[15]) ? 4'b1111 : node53827;
															assign node53827 = (inp[0]) ? 4'b1101 : 4'b1111;
														assign node53831 = (inp[0]) ? 4'b1101 : node53832;
															assign node53832 = (inp[3]) ? 4'b1101 : node53833;
																assign node53833 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node53838 = (inp[12]) ? node53854 : node53839;
														assign node53839 = (inp[3]) ? node53847 : node53840;
															assign node53840 = (inp[15]) ? node53844 : node53841;
																assign node53841 = (inp[0]) ? 4'b1111 : 4'b1101;
																assign node53844 = (inp[0]) ? 4'b1101 : 4'b1111;
															assign node53847 = (inp[0]) ? node53851 : node53848;
																assign node53848 = (inp[15]) ? 4'b1111 : 4'b1101;
																assign node53851 = (inp[15]) ? 4'b1101 : 4'b1111;
														assign node53854 = (inp[15]) ? 4'b1111 : node53855;
															assign node53855 = (inp[0]) ? 4'b1111 : 4'b1101;
											assign node53859 = (inp[5]) ? node53879 : node53860;
												assign node53860 = (inp[15]) ? node53868 : node53861;
													assign node53861 = (inp[0]) ? node53865 : node53862;
														assign node53862 = (inp[3]) ? 4'b1101 : 4'b1111;
														assign node53865 = (inp[3]) ? 4'b1111 : 4'b1101;
													assign node53868 = (inp[12]) ? node53874 : node53869;
														assign node53869 = (inp[3]) ? 4'b1101 : node53870;
															assign node53870 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node53874 = (inp[0]) ? 4'b1101 : node53875;
															assign node53875 = (inp[3]) ? 4'b1111 : 4'b1101;
												assign node53879 = (inp[0]) ? node53883 : node53880;
													assign node53880 = (inp[15]) ? 4'b1111 : 4'b1101;
													assign node53883 = (inp[15]) ? 4'b1101 : 4'b1111;
										assign node53886 = (inp[14]) ? node53940 : node53887;
											assign node53887 = (inp[2]) ? node53919 : node53888;
												assign node53888 = (inp[5]) ? node53906 : node53889;
													assign node53889 = (inp[12]) ? node53893 : node53890;
														assign node53890 = (inp[3]) ? 4'b1111 : 4'b1101;
														assign node53893 = (inp[0]) ? node53901 : node53894;
															assign node53894 = (inp[3]) ? node53898 : node53895;
																assign node53895 = (inp[15]) ? 4'b1101 : 4'b1111;
																assign node53898 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node53901 = (inp[3]) ? 4'b1101 : node53902;
																assign node53902 = (inp[15]) ? 4'b1111 : 4'b1101;
													assign node53906 = (inp[12]) ? node53912 : node53907;
														assign node53907 = (inp[3]) ? 4'b1101 : node53908;
															assign node53908 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node53912 = (inp[0]) ? node53916 : node53913;
															assign node53913 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node53916 = (inp[15]) ? 4'b1101 : 4'b1111;
												assign node53919 = (inp[5]) ? node53933 : node53920;
													assign node53920 = (inp[15]) ? node53926 : node53921;
														assign node53921 = (inp[12]) ? 4'b1100 : node53922;
															assign node53922 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node53926 = (inp[0]) ? node53930 : node53927;
															assign node53927 = (inp[3]) ? 4'b1110 : 4'b1100;
															assign node53930 = (inp[3]) ? 4'b1100 : 4'b1110;
													assign node53933 = (inp[0]) ? node53937 : node53934;
														assign node53934 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node53937 = (inp[15]) ? 4'b1100 : 4'b1110;
											assign node53940 = (inp[5]) ? node53970 : node53941;
												assign node53941 = (inp[12]) ? node53957 : node53942;
													assign node53942 = (inp[15]) ? 4'b1100 : node53943;
														assign node53943 = (inp[2]) ? node53949 : node53944;
															assign node53944 = (inp[0]) ? 4'b1100 : node53945;
																assign node53945 = (inp[3]) ? 4'b1100 : 4'b1110;
															assign node53949 = (inp[0]) ? node53953 : node53950;
																assign node53950 = (inp[3]) ? 4'b1100 : 4'b1110;
																assign node53953 = (inp[3]) ? 4'b1110 : 4'b1100;
													assign node53957 = (inp[15]) ? node53963 : node53958;
														assign node53958 = (inp[0]) ? node53960 : 4'b1100;
															assign node53960 = (inp[3]) ? 4'b1110 : 4'b1100;
														assign node53963 = (inp[3]) ? node53967 : node53964;
															assign node53964 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node53967 = (inp[0]) ? 4'b1100 : 4'b1110;
												assign node53970 = (inp[0]) ? node53974 : node53971;
													assign node53971 = (inp[15]) ? 4'b1110 : 4'b1100;
													assign node53974 = (inp[15]) ? 4'b1100 : 4'b1110;
							assign node53977 = (inp[4]) ? node54415 : node53978;
								assign node53978 = (inp[12]) ? node54210 : node53979;
									assign node53979 = (inp[15]) ? node54091 : node53980;
										assign node53980 = (inp[0]) ? node54036 : node53981;
											assign node53981 = (inp[5]) ? node54015 : node53982;
												assign node53982 = (inp[3]) ? node54008 : node53983;
													assign node53983 = (inp[14]) ? node53997 : node53984;
														assign node53984 = (inp[7]) ? node53990 : node53985;
															assign node53985 = (inp[2]) ? 4'b1110 : node53986;
																assign node53986 = (inp[8]) ? 4'b1110 : 4'b1111;
															assign node53990 = (inp[2]) ? node53994 : node53991;
																assign node53991 = (inp[8]) ? 4'b1111 : 4'b1110;
																assign node53994 = (inp[8]) ? 4'b1110 : 4'b1111;
														assign node53997 = (inp[2]) ? node54003 : node53998;
															assign node53998 = (inp[7]) ? node54000 : 4'b1111;
																assign node54000 = (inp[8]) ? 4'b1110 : 4'b1111;
															assign node54003 = (inp[8]) ? 4'b1111 : node54004;
																assign node54004 = (inp[7]) ? 4'b1111 : 4'b1110;
													assign node54008 = (inp[14]) ? node54010 : 4'b1100;
														assign node54010 = (inp[7]) ? 4'b1101 : node54011;
															assign node54011 = (inp[8]) ? 4'b1101 : 4'b1100;
												assign node54015 = (inp[3]) ? node54027 : node54016;
													assign node54016 = (inp[7]) ? node54018 : 4'b1101;
														assign node54018 = (inp[14]) ? node54024 : node54019;
															assign node54019 = (inp[2]) ? 4'b1101 : node54020;
																assign node54020 = (inp[8]) ? 4'b1101 : 4'b1100;
															assign node54024 = (inp[8]) ? 4'b1100 : 4'b1101;
													assign node54027 = (inp[8]) ? node54029 : 4'b1100;
														assign node54029 = (inp[2]) ? 4'b1101 : node54030;
															assign node54030 = (inp[7]) ? 4'b1100 : node54031;
																assign node54031 = (inp[14]) ? 4'b1101 : 4'b1100;
											assign node54036 = (inp[5]) ? node54076 : node54037;
												assign node54037 = (inp[3]) ? node54053 : node54038;
													assign node54038 = (inp[2]) ? node54048 : node54039;
														assign node54039 = (inp[8]) ? node54041 : 4'b1101;
															assign node54041 = (inp[14]) ? node54045 : node54042;
																assign node54042 = (inp[7]) ? 4'b1101 : 4'b1100;
																assign node54045 = (inp[7]) ? 4'b1100 : 4'b1101;
														assign node54048 = (inp[7]) ? node54050 : 4'b1100;
															assign node54050 = (inp[8]) ? 4'b1100 : 4'b1101;
													assign node54053 = (inp[2]) ? node54069 : node54054;
														assign node54054 = (inp[7]) ? node54062 : node54055;
															assign node54055 = (inp[14]) ? node54059 : node54056;
																assign node54056 = (inp[8]) ? 4'b1110 : 4'b1111;
																assign node54059 = (inp[8]) ? 4'b1111 : 4'b1110;
															assign node54062 = (inp[8]) ? node54066 : node54063;
																assign node54063 = (inp[14]) ? 4'b1111 : 4'b1110;
																assign node54066 = (inp[14]) ? 4'b1110 : 4'b1111;
														assign node54069 = (inp[7]) ? node54073 : node54070;
															assign node54070 = (inp[8]) ? 4'b1111 : 4'b1110;
															assign node54073 = (inp[8]) ? 4'b1110 : 4'b1111;
												assign node54076 = (inp[7]) ? node54084 : node54077;
													assign node54077 = (inp[8]) ? 4'b1111 : node54078;
														assign node54078 = (inp[14]) ? 4'b1110 : node54079;
															assign node54079 = (inp[2]) ? 4'b1110 : 4'b1111;
													assign node54084 = (inp[8]) ? 4'b1110 : node54085;
														assign node54085 = (inp[14]) ? 4'b1111 : node54086;
															assign node54086 = (inp[2]) ? 4'b1111 : 4'b1110;
										assign node54091 = (inp[0]) ? node54167 : node54092;
											assign node54092 = (inp[5]) ? node54126 : node54093;
												assign node54093 = (inp[3]) ? node54107 : node54094;
													assign node54094 = (inp[8]) ? node54100 : node54095;
														assign node54095 = (inp[7]) ? 4'b1101 : node54096;
															assign node54096 = (inp[2]) ? 4'b1100 : 4'b1101;
														assign node54100 = (inp[7]) ? 4'b1100 : node54101;
															assign node54101 = (inp[2]) ? 4'b1101 : node54102;
																assign node54102 = (inp[14]) ? 4'b1101 : 4'b1100;
													assign node54107 = (inp[14]) ? node54121 : node54108;
														assign node54108 = (inp[2]) ? node54116 : node54109;
															assign node54109 = (inp[7]) ? node54113 : node54110;
																assign node54110 = (inp[8]) ? 4'b1110 : 4'b1111;
																assign node54113 = (inp[8]) ? 4'b1111 : 4'b1110;
															assign node54116 = (inp[7]) ? 4'b1110 : node54117;
																assign node54117 = (inp[8]) ? 4'b1111 : 4'b1110;
														assign node54121 = (inp[2]) ? node54123 : 4'b1110;
															assign node54123 = (inp[7]) ? 4'b1111 : 4'b1110;
												assign node54126 = (inp[3]) ? node54146 : node54127;
													assign node54127 = (inp[2]) ? node54141 : node54128;
														assign node54128 = (inp[14]) ? node54136 : node54129;
															assign node54129 = (inp[7]) ? node54133 : node54130;
																assign node54130 = (inp[8]) ? 4'b1110 : 4'b1111;
																assign node54133 = (inp[8]) ? 4'b1111 : 4'b1110;
															assign node54136 = (inp[8]) ? node54138 : 4'b1111;
																assign node54138 = (inp[7]) ? 4'b1110 : 4'b1111;
														assign node54141 = (inp[7]) ? 4'b1111 : node54142;
															assign node54142 = (inp[8]) ? 4'b1111 : 4'b1110;
													assign node54146 = (inp[14]) ? node54160 : node54147;
														assign node54147 = (inp[2]) ? node54153 : node54148;
															assign node54148 = (inp[8]) ? node54150 : 4'b1111;
																assign node54150 = (inp[7]) ? 4'b1111 : 4'b1110;
															assign node54153 = (inp[7]) ? node54157 : node54154;
																assign node54154 = (inp[8]) ? 4'b1111 : 4'b1110;
																assign node54157 = (inp[8]) ? 4'b1110 : 4'b1111;
														assign node54160 = (inp[7]) ? node54164 : node54161;
															assign node54161 = (inp[2]) ? 4'b1111 : 4'b1110;
															assign node54164 = (inp[8]) ? 4'b1110 : 4'b1111;
											assign node54167 = (inp[5]) ? node54189 : node54168;
												assign node54168 = (inp[3]) ? node54178 : node54169;
													assign node54169 = (inp[7]) ? 4'b1110 : node54170;
														assign node54170 = (inp[2]) ? 4'b1110 : node54171;
															assign node54171 = (inp[14]) ? 4'b1111 : node54172;
																assign node54172 = (inp[8]) ? 4'b1110 : 4'b1111;
													assign node54178 = (inp[14]) ? node54180 : 4'b1101;
														assign node54180 = (inp[2]) ? node54182 : 4'b1100;
															assign node54182 = (inp[7]) ? node54186 : node54183;
																assign node54183 = (inp[8]) ? 4'b1101 : 4'b1100;
																assign node54186 = (inp[8]) ? 4'b1100 : 4'b1101;
												assign node54189 = (inp[2]) ? node54203 : node54190;
													assign node54190 = (inp[7]) ? node54198 : node54191;
														assign node54191 = (inp[14]) ? node54195 : node54192;
															assign node54192 = (inp[8]) ? 4'b1100 : 4'b1101;
															assign node54195 = (inp[8]) ? 4'b1101 : 4'b1100;
														assign node54198 = (inp[8]) ? 4'b1101 : node54199;
															assign node54199 = (inp[3]) ? 4'b1100 : 4'b1101;
													assign node54203 = (inp[7]) ? node54207 : node54204;
														assign node54204 = (inp[8]) ? 4'b1101 : 4'b1100;
														assign node54207 = (inp[8]) ? 4'b1100 : 4'b1101;
									assign node54210 = (inp[2]) ? node54316 : node54211;
										assign node54211 = (inp[0]) ? node54269 : node54212;
											assign node54212 = (inp[15]) ? node54242 : node54213;
												assign node54213 = (inp[3]) ? node54225 : node54214;
													assign node54214 = (inp[5]) ? 4'b1101 : node54215;
														assign node54215 = (inp[7]) ? 4'b1110 : node54216;
															assign node54216 = (inp[8]) ? node54220 : node54217;
																assign node54217 = (inp[14]) ? 4'b1110 : 4'b1111;
																assign node54220 = (inp[14]) ? 4'b1111 : 4'b1110;
													assign node54225 = (inp[5]) ? node54233 : node54226;
														assign node54226 = (inp[7]) ? 4'b1101 : node54227;
															assign node54227 = (inp[14]) ? 4'b1101 : node54228;
																assign node54228 = (inp[8]) ? 4'b1100 : 4'b1101;
														assign node54233 = (inp[8]) ? 4'b1101 : node54234;
															assign node54234 = (inp[7]) ? node54238 : node54235;
																assign node54235 = (inp[14]) ? 4'b1100 : 4'b1101;
																assign node54238 = (inp[14]) ? 4'b1101 : 4'b1100;
												assign node54242 = (inp[3]) ? node54248 : node54243;
													assign node54243 = (inp[5]) ? node54245 : 4'b1101;
														assign node54245 = (inp[14]) ? 4'b1110 : 4'b1111;
													assign node54248 = (inp[5]) ? node54260 : node54249;
														assign node54249 = (inp[7]) ? node54255 : node54250;
															assign node54250 = (inp[8]) ? node54252 : 4'b1110;
																assign node54252 = (inp[14]) ? 4'b1111 : 4'b1110;
															assign node54255 = (inp[14]) ? node54257 : 4'b1111;
																assign node54257 = (inp[8]) ? 4'b1110 : 4'b1111;
														assign node54260 = (inp[7]) ? node54262 : 4'b1111;
															assign node54262 = (inp[8]) ? node54266 : node54263;
																assign node54263 = (inp[14]) ? 4'b1111 : 4'b1110;
																assign node54266 = (inp[14]) ? 4'b1110 : 4'b1111;
											assign node54269 = (inp[15]) ? node54295 : node54270;
												assign node54270 = (inp[3]) ? node54282 : node54271;
													assign node54271 = (inp[5]) ? node54275 : node54272;
														assign node54272 = (inp[7]) ? 4'b1100 : 4'b1101;
														assign node54275 = (inp[8]) ? node54279 : node54276;
															assign node54276 = (inp[7]) ? 4'b1110 : 4'b1111;
															assign node54279 = (inp[7]) ? 4'b1111 : 4'b1110;
													assign node54282 = (inp[5]) ? node54284 : 4'b1111;
														assign node54284 = (inp[14]) ? node54290 : node54285;
															assign node54285 = (inp[8]) ? 4'b1110 : node54286;
																assign node54286 = (inp[7]) ? 4'b1110 : 4'b1111;
															assign node54290 = (inp[7]) ? 4'b1111 : node54291;
																assign node54291 = (inp[8]) ? 4'b1111 : 4'b1110;
												assign node54295 = (inp[3]) ? node54303 : node54296;
													assign node54296 = (inp[5]) ? node54300 : node54297;
														assign node54297 = (inp[14]) ? 4'b1110 : 4'b1111;
														assign node54300 = (inp[14]) ? 4'b1101 : 4'b1100;
													assign node54303 = (inp[8]) ? node54309 : node54304;
														assign node54304 = (inp[7]) ? node54306 : 4'b1100;
															assign node54306 = (inp[14]) ? 4'b1101 : 4'b1100;
														assign node54309 = (inp[7]) ? node54313 : node54310;
															assign node54310 = (inp[14]) ? 4'b1101 : 4'b1100;
															assign node54313 = (inp[14]) ? 4'b1100 : 4'b1101;
										assign node54316 = (inp[7]) ? node54370 : node54317;
											assign node54317 = (inp[8]) ? node54335 : node54318;
												assign node54318 = (inp[0]) ? node54330 : node54319;
													assign node54319 = (inp[15]) ? node54325 : node54320;
														assign node54320 = (inp[5]) ? 4'b1100 : node54321;
															assign node54321 = (inp[3]) ? 4'b1100 : 4'b1110;
														assign node54325 = (inp[3]) ? 4'b1110 : node54326;
															assign node54326 = (inp[5]) ? 4'b1110 : 4'b1100;
													assign node54330 = (inp[15]) ? 4'b1100 : node54331;
														assign node54331 = (inp[5]) ? 4'b1110 : 4'b1100;
												assign node54335 = (inp[14]) ? node54349 : node54336;
													assign node54336 = (inp[0]) ? node54346 : node54337;
														assign node54337 = (inp[3]) ? node54343 : node54338;
															assign node54338 = (inp[5]) ? 4'b1111 : node54339;
																assign node54339 = (inp[15]) ? 4'b1101 : 4'b1111;
															assign node54343 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node54346 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node54349 = (inp[5]) ? node54357 : node54350;
														assign node54350 = (inp[3]) ? 4'b1101 : node54351;
															assign node54351 = (inp[0]) ? node54353 : 4'b1101;
																assign node54353 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node54357 = (inp[3]) ? node54363 : node54358;
															assign node54358 = (inp[0]) ? node54360 : 4'b1101;
																assign node54360 = (inp[15]) ? 4'b1101 : 4'b1111;
															assign node54363 = (inp[15]) ? node54367 : node54364;
																assign node54364 = (inp[0]) ? 4'b1111 : 4'b1101;
																assign node54367 = (inp[0]) ? 4'b1101 : 4'b1111;
											assign node54370 = (inp[8]) ? node54390 : node54371;
												assign node54371 = (inp[15]) ? node54379 : node54372;
													assign node54372 = (inp[0]) ? 4'b1111 : node54373;
														assign node54373 = (inp[5]) ? 4'b1101 : node54374;
															assign node54374 = (inp[3]) ? 4'b1101 : 4'b1111;
													assign node54379 = (inp[0]) ? node54385 : node54380;
														assign node54380 = (inp[3]) ? 4'b1111 : node54381;
															assign node54381 = (inp[5]) ? 4'b1111 : 4'b1101;
														assign node54385 = (inp[5]) ? 4'b1101 : node54386;
															assign node54386 = (inp[3]) ? 4'b1101 : 4'b1111;
												assign node54390 = (inp[3]) ? node54408 : node54391;
													assign node54391 = (inp[14]) ? node54403 : node54392;
														assign node54392 = (inp[5]) ? node54398 : node54393;
															assign node54393 = (inp[15]) ? node54395 : 4'b1100;
																assign node54395 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node54398 = (inp[0]) ? node54400 : 4'b1110;
																assign node54400 = (inp[15]) ? 4'b1100 : 4'b1110;
														assign node54403 = (inp[0]) ? 4'b1100 : node54404;
															assign node54404 = (inp[15]) ? 4'b1100 : 4'b1110;
													assign node54408 = (inp[15]) ? node54412 : node54409;
														assign node54409 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node54412 = (inp[0]) ? 4'b1100 : 4'b1110;
								assign node54415 = (inp[8]) ? node54589 : node54416;
									assign node54416 = (inp[7]) ? node54508 : node54417;
										assign node54417 = (inp[2]) ? node54475 : node54418;
											assign node54418 = (inp[14]) ? node54442 : node54419;
												assign node54419 = (inp[0]) ? node54431 : node54420;
													assign node54420 = (inp[15]) ? node54426 : node54421;
														assign node54421 = (inp[3]) ? 4'b1001 : node54422;
															assign node54422 = (inp[5]) ? 4'b1001 : 4'b1011;
														assign node54426 = (inp[3]) ? 4'b1011 : node54427;
															assign node54427 = (inp[5]) ? 4'b1011 : 4'b1001;
													assign node54431 = (inp[15]) ? node54437 : node54432;
														assign node54432 = (inp[5]) ? 4'b1011 : node54433;
															assign node54433 = (inp[12]) ? 4'b1011 : 4'b1001;
														assign node54437 = (inp[5]) ? 4'b1001 : node54438;
															assign node54438 = (inp[3]) ? 4'b1001 : 4'b1011;
												assign node54442 = (inp[12]) ? node54456 : node54443;
													assign node54443 = (inp[15]) ? node54453 : node54444;
														assign node54444 = (inp[0]) ? node54448 : node54445;
															assign node54445 = (inp[5]) ? 4'b1000 : 4'b1010;
															assign node54448 = (inp[3]) ? 4'b1010 : node54449;
																assign node54449 = (inp[5]) ? 4'b1010 : 4'b1000;
														assign node54453 = (inp[0]) ? 4'b1000 : 4'b1010;
													assign node54456 = (inp[15]) ? node54464 : node54457;
														assign node54457 = (inp[0]) ? 4'b1010 : node54458;
															assign node54458 = (inp[3]) ? 4'b1000 : node54459;
																assign node54459 = (inp[5]) ? 4'b1000 : 4'b1010;
														assign node54464 = (inp[0]) ? node54470 : node54465;
															assign node54465 = (inp[3]) ? 4'b1010 : node54466;
																assign node54466 = (inp[5]) ? 4'b1010 : 4'b1000;
															assign node54470 = (inp[3]) ? 4'b1000 : node54471;
																assign node54471 = (inp[5]) ? 4'b1000 : 4'b1010;
											assign node54475 = (inp[3]) ? node54493 : node54476;
												assign node54476 = (inp[15]) ? node54486 : node54477;
													assign node54477 = (inp[14]) ? 4'b1010 : node54478;
														assign node54478 = (inp[5]) ? node54482 : node54479;
															assign node54479 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node54482 = (inp[0]) ? 4'b1010 : 4'b1000;
													assign node54486 = (inp[0]) ? node54490 : node54487;
														assign node54487 = (inp[5]) ? 4'b1010 : 4'b1000;
														assign node54490 = (inp[5]) ? 4'b1000 : 4'b1010;
												assign node54493 = (inp[14]) ? node54501 : node54494;
													assign node54494 = (inp[0]) ? node54498 : node54495;
														assign node54495 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node54498 = (inp[15]) ? 4'b1000 : 4'b1010;
													assign node54501 = (inp[0]) ? node54505 : node54502;
														assign node54502 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node54505 = (inp[15]) ? 4'b1000 : 4'b1010;
										assign node54508 = (inp[14]) ? node54566 : node54509;
											assign node54509 = (inp[2]) ? node54549 : node54510;
												assign node54510 = (inp[5]) ? node54532 : node54511;
													assign node54511 = (inp[12]) ? node54525 : node54512;
														assign node54512 = (inp[3]) ? node54520 : node54513;
															assign node54513 = (inp[15]) ? node54517 : node54514;
																assign node54514 = (inp[0]) ? 4'b1000 : 4'b1010;
																assign node54517 = (inp[0]) ? 4'b1010 : 4'b1000;
															assign node54520 = (inp[0]) ? node54522 : 4'b1000;
																assign node54522 = (inp[15]) ? 4'b1000 : 4'b1010;
														assign node54525 = (inp[0]) ? node54527 : 4'b1000;
															assign node54527 = (inp[15]) ? node54529 : 4'b1000;
																assign node54529 = (inp[3]) ? 4'b1000 : 4'b1010;
													assign node54532 = (inp[3]) ? node54540 : node54533;
														assign node54533 = (inp[15]) ? node54537 : node54534;
															assign node54534 = (inp[0]) ? 4'b1010 : 4'b1000;
															assign node54537 = (inp[0]) ? 4'b1000 : 4'b1010;
														assign node54540 = (inp[12]) ? node54542 : 4'b1010;
															assign node54542 = (inp[0]) ? node54546 : node54543;
																assign node54543 = (inp[15]) ? 4'b1010 : 4'b1000;
																assign node54546 = (inp[15]) ? 4'b1000 : 4'b1010;
												assign node54549 = (inp[3]) ? node54559 : node54550;
													assign node54550 = (inp[0]) ? 4'b1001 : node54551;
														assign node54551 = (inp[12]) ? node54553 : 4'b1011;
															assign node54553 = (inp[15]) ? 4'b1001 : node54554;
																assign node54554 = (inp[5]) ? 4'b1001 : 4'b1011;
													assign node54559 = (inp[0]) ? node54563 : node54560;
														assign node54560 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node54563 = (inp[15]) ? 4'b1001 : 4'b1011;
											assign node54566 = (inp[15]) ? node54578 : node54567;
												assign node54567 = (inp[0]) ? node54573 : node54568;
													assign node54568 = (inp[5]) ? 4'b1001 : node54569;
														assign node54569 = (inp[3]) ? 4'b1001 : 4'b1011;
													assign node54573 = (inp[3]) ? 4'b1011 : node54574;
														assign node54574 = (inp[5]) ? 4'b1011 : 4'b1001;
												assign node54578 = (inp[0]) ? node54584 : node54579;
													assign node54579 = (inp[3]) ? 4'b1011 : node54580;
														assign node54580 = (inp[5]) ? 4'b1011 : 4'b1001;
													assign node54584 = (inp[5]) ? 4'b1001 : node54585;
														assign node54585 = (inp[3]) ? 4'b1001 : 4'b1011;
									assign node54589 = (inp[7]) ? node54695 : node54590;
										assign node54590 = (inp[14]) ? node54656 : node54591;
											assign node54591 = (inp[2]) ? node54627 : node54592;
												assign node54592 = (inp[12]) ? node54612 : node54593;
													assign node54593 = (inp[3]) ? node54607 : node54594;
														assign node54594 = (inp[5]) ? node54600 : node54595;
															assign node54595 = (inp[0]) ? node54597 : 4'b1000;
																assign node54597 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node54600 = (inp[0]) ? node54604 : node54601;
																assign node54601 = (inp[15]) ? 4'b1010 : 4'b1000;
																assign node54604 = (inp[15]) ? 4'b1000 : 4'b1010;
														assign node54607 = (inp[0]) ? node54609 : 4'b1010;
															assign node54609 = (inp[15]) ? 4'b1000 : 4'b1010;
													assign node54612 = (inp[5]) ? node54620 : node54613;
														assign node54613 = (inp[0]) ? 4'b1010 : node54614;
															assign node54614 = (inp[15]) ? 4'b1010 : node54615;
																assign node54615 = (inp[3]) ? 4'b1000 : 4'b1010;
														assign node54620 = (inp[0]) ? node54624 : node54621;
															assign node54621 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node54624 = (inp[15]) ? 4'b1000 : 4'b1010;
												assign node54627 = (inp[3]) ? node54645 : node54628;
													assign node54628 = (inp[15]) ? node54638 : node54629;
														assign node54629 = (inp[12]) ? node54635 : node54630;
															assign node54630 = (inp[0]) ? node54632 : 4'b1001;
																assign node54632 = (inp[5]) ? 4'b1011 : 4'b1001;
															assign node54635 = (inp[5]) ? 4'b1001 : 4'b1011;
														assign node54638 = (inp[5]) ? node54642 : node54639;
															assign node54639 = (inp[12]) ? 4'b1001 : 4'b1011;
															assign node54642 = (inp[0]) ? 4'b1001 : 4'b1011;
													assign node54645 = (inp[5]) ? 4'b1011 : node54646;
														assign node54646 = (inp[12]) ? node54650 : node54647;
															assign node54647 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node54650 = (inp[15]) ? 4'b1011 : node54651;
																assign node54651 = (inp[0]) ? 4'b1011 : 4'b1001;
											assign node54656 = (inp[3]) ? node54688 : node54657;
												assign node54657 = (inp[0]) ? node54673 : node54658;
													assign node54658 = (inp[12]) ? node54660 : 4'b1011;
														assign node54660 = (inp[2]) ? node54668 : node54661;
															assign node54661 = (inp[15]) ? node54665 : node54662;
																assign node54662 = (inp[5]) ? 4'b1001 : 4'b1011;
																assign node54665 = (inp[5]) ? 4'b1011 : 4'b1001;
															assign node54668 = (inp[5]) ? node54670 : 4'b1011;
																assign node54670 = (inp[15]) ? 4'b1011 : 4'b1001;
													assign node54673 = (inp[12]) ? node54681 : node54674;
														assign node54674 = (inp[15]) ? node54678 : node54675;
															assign node54675 = (inp[5]) ? 4'b1011 : 4'b1001;
															assign node54678 = (inp[5]) ? 4'b1001 : 4'b1011;
														assign node54681 = (inp[15]) ? node54685 : node54682;
															assign node54682 = (inp[5]) ? 4'b1011 : 4'b1001;
															assign node54685 = (inp[5]) ? 4'b1001 : 4'b1011;
												assign node54688 = (inp[0]) ? node54692 : node54689;
													assign node54689 = (inp[15]) ? 4'b1011 : 4'b1001;
													assign node54692 = (inp[15]) ? 4'b1001 : 4'b1011;
										assign node54695 = (inp[2]) ? node54761 : node54696;
											assign node54696 = (inp[14]) ? node54734 : node54697;
												assign node54697 = (inp[5]) ? node54713 : node54698;
													assign node54698 = (inp[15]) ? node54708 : node54699;
														assign node54699 = (inp[12]) ? node54701 : 4'b1011;
															assign node54701 = (inp[3]) ? node54705 : node54702;
																assign node54702 = (inp[0]) ? 4'b1001 : 4'b1011;
																assign node54705 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node54708 = (inp[0]) ? 4'b1011 : node54709;
															assign node54709 = (inp[3]) ? 4'b1011 : 4'b1001;
													assign node54713 = (inp[12]) ? node54727 : node54714;
														assign node54714 = (inp[3]) ? node54722 : node54715;
															assign node54715 = (inp[15]) ? node54719 : node54716;
																assign node54716 = (inp[0]) ? 4'b1011 : 4'b1001;
																assign node54719 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node54722 = (inp[15]) ? node54724 : 4'b1001;
																assign node54724 = (inp[0]) ? 4'b1001 : 4'b1011;
														assign node54727 = (inp[15]) ? node54731 : node54728;
															assign node54728 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node54731 = (inp[0]) ? 4'b1001 : 4'b1011;
												assign node54734 = (inp[12]) ? node54750 : node54735;
													assign node54735 = (inp[5]) ? node54743 : node54736;
														assign node54736 = (inp[3]) ? node54738 : 4'b1010;
															assign node54738 = (inp[0]) ? 4'b1000 : node54739;
																assign node54739 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node54743 = (inp[15]) ? node54747 : node54744;
															assign node54744 = (inp[0]) ? 4'b1010 : 4'b1000;
															assign node54747 = (inp[0]) ? 4'b1000 : 4'b1010;
													assign node54750 = (inp[3]) ? 4'b1010 : node54751;
														assign node54751 = (inp[0]) ? 4'b1010 : node54752;
															assign node54752 = (inp[15]) ? node54756 : node54753;
																assign node54753 = (inp[5]) ? 4'b1000 : 4'b1010;
																assign node54756 = (inp[5]) ? 4'b1010 : 4'b1000;
											assign node54761 = (inp[0]) ? node54773 : node54762;
												assign node54762 = (inp[15]) ? node54768 : node54763;
													assign node54763 = (inp[3]) ? 4'b1000 : node54764;
														assign node54764 = (inp[5]) ? 4'b1000 : 4'b1010;
													assign node54768 = (inp[3]) ? 4'b1010 : node54769;
														assign node54769 = (inp[5]) ? 4'b1010 : 4'b1000;
												assign node54773 = (inp[15]) ? node54779 : node54774;
													assign node54774 = (inp[5]) ? 4'b1010 : node54775;
														assign node54775 = (inp[3]) ? 4'b1010 : 4'b1000;
													assign node54779 = (inp[3]) ? 4'b1000 : node54780;
														assign node54780 = (inp[5]) ? 4'b1000 : 4'b1010;
				assign node54784 = (inp[13]) ? node58044 : node54785;
					assign node54785 = (inp[1]) ? node56447 : node54786;
						assign node54786 = (inp[9]) ? node55514 : node54787;
							assign node54787 = (inp[4]) ? node55121 : node54788;
								assign node54788 = (inp[15]) ? node54954 : node54789;
									assign node54789 = (inp[0]) ? node54869 : node54790;
										assign node54790 = (inp[5]) ? node54814 : node54791;
											assign node54791 = (inp[7]) ? node54803 : node54792;
												assign node54792 = (inp[8]) ? node54798 : node54793;
													assign node54793 = (inp[2]) ? 4'b1010 : node54794;
														assign node54794 = (inp[14]) ? 4'b1010 : 4'b1011;
													assign node54798 = (inp[14]) ? 4'b1011 : node54799;
														assign node54799 = (inp[2]) ? 4'b1011 : 4'b1010;
												assign node54803 = (inp[8]) ? node54809 : node54804;
													assign node54804 = (inp[2]) ? 4'b1011 : node54805;
														assign node54805 = (inp[14]) ? 4'b1011 : 4'b1010;
													assign node54809 = (inp[14]) ? 4'b1010 : node54810;
														assign node54810 = (inp[2]) ? 4'b1010 : 4'b1011;
											assign node54814 = (inp[3]) ? node54838 : node54815;
												assign node54815 = (inp[2]) ? node54831 : node54816;
													assign node54816 = (inp[7]) ? node54824 : node54817;
														assign node54817 = (inp[14]) ? node54821 : node54818;
															assign node54818 = (inp[8]) ? 4'b1010 : 4'b1011;
															assign node54821 = (inp[8]) ? 4'b1011 : 4'b1010;
														assign node54824 = (inp[12]) ? 4'b1010 : node54825;
															assign node54825 = (inp[8]) ? node54827 : 4'b1010;
																assign node54827 = (inp[14]) ? 4'b1010 : 4'b1011;
													assign node54831 = (inp[7]) ? node54835 : node54832;
														assign node54832 = (inp[8]) ? 4'b1011 : 4'b1010;
														assign node54835 = (inp[8]) ? 4'b1010 : 4'b1011;
												assign node54838 = (inp[12]) ? node54854 : node54839;
													assign node54839 = (inp[2]) ? node54847 : node54840;
														assign node54840 = (inp[14]) ? 4'b1000 : node54841;
															assign node54841 = (inp[7]) ? 4'b1001 : node54842;
																assign node54842 = (inp[8]) ? 4'b1000 : 4'b1001;
														assign node54847 = (inp[14]) ? 4'b1001 : node54848;
															assign node54848 = (inp[7]) ? node54850 : 4'b1001;
																assign node54850 = (inp[8]) ? 4'b1000 : 4'b1001;
													assign node54854 = (inp[14]) ? 4'b1000 : node54855;
														assign node54855 = (inp[8]) ? node54863 : node54856;
															assign node54856 = (inp[2]) ? node54860 : node54857;
																assign node54857 = (inp[7]) ? 4'b1000 : 4'b1001;
																assign node54860 = (inp[7]) ? 4'b1001 : 4'b1000;
															assign node54863 = (inp[2]) ? node54865 : 4'b1001;
																assign node54865 = (inp[7]) ? 4'b1000 : 4'b1001;
										assign node54869 = (inp[3]) ? node54893 : node54870;
											assign node54870 = (inp[7]) ? node54882 : node54871;
												assign node54871 = (inp[8]) ? node54877 : node54872;
													assign node54872 = (inp[14]) ? 4'b1000 : node54873;
														assign node54873 = (inp[2]) ? 4'b1000 : 4'b1001;
													assign node54877 = (inp[2]) ? 4'b1001 : node54878;
														assign node54878 = (inp[14]) ? 4'b1001 : 4'b1000;
												assign node54882 = (inp[8]) ? node54888 : node54883;
													assign node54883 = (inp[2]) ? 4'b1001 : node54884;
														assign node54884 = (inp[14]) ? 4'b1001 : 4'b1000;
													assign node54888 = (inp[14]) ? 4'b1000 : node54889;
														assign node54889 = (inp[2]) ? 4'b1000 : 4'b1001;
											assign node54893 = (inp[5]) ? node54923 : node54894;
												assign node54894 = (inp[2]) ? node54908 : node54895;
													assign node54895 = (inp[8]) ? node54901 : node54896;
														assign node54896 = (inp[7]) ? 4'b1000 : node54897;
															assign node54897 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node54901 = (inp[7]) ? node54905 : node54902;
															assign node54902 = (inp[14]) ? 4'b1001 : 4'b1000;
															assign node54905 = (inp[14]) ? 4'b1000 : 4'b1001;
													assign node54908 = (inp[12]) ? node54916 : node54909;
														assign node54909 = (inp[7]) ? node54913 : node54910;
															assign node54910 = (inp[8]) ? 4'b1001 : 4'b1000;
															assign node54913 = (inp[8]) ? 4'b1000 : 4'b1001;
														assign node54916 = (inp[7]) ? node54920 : node54917;
															assign node54917 = (inp[8]) ? 4'b1001 : 4'b1000;
															assign node54920 = (inp[8]) ? 4'b1000 : 4'b1001;
												assign node54923 = (inp[2]) ? node54935 : node54924;
													assign node54924 = (inp[7]) ? node54926 : 4'b1011;
														assign node54926 = (inp[12]) ? 4'b1011 : node54927;
															assign node54927 = (inp[14]) ? node54931 : node54928;
																assign node54928 = (inp[8]) ? 4'b1011 : 4'b1010;
																assign node54931 = (inp[8]) ? 4'b1010 : 4'b1011;
													assign node54935 = (inp[14]) ? node54949 : node54936;
														assign node54936 = (inp[12]) ? node54944 : node54937;
															assign node54937 = (inp[8]) ? node54941 : node54938;
																assign node54938 = (inp[7]) ? 4'b1011 : 4'b1010;
																assign node54941 = (inp[7]) ? 4'b1010 : 4'b1011;
															assign node54944 = (inp[7]) ? 4'b1011 : node54945;
																assign node54945 = (inp[8]) ? 4'b1011 : 4'b1010;
														assign node54949 = (inp[7]) ? 4'b1010 : node54950;
															assign node54950 = (inp[8]) ? 4'b1011 : 4'b1010;
									assign node54954 = (inp[0]) ? node55050 : node54955;
										assign node54955 = (inp[3]) ? node54987 : node54956;
											assign node54956 = (inp[2]) ? node54980 : node54957;
												assign node54957 = (inp[7]) ? node54975 : node54958;
													assign node54958 = (inp[5]) ? node54966 : node54959;
														assign node54959 = (inp[14]) ? node54963 : node54960;
															assign node54960 = (inp[8]) ? 4'b1000 : 4'b1001;
															assign node54963 = (inp[8]) ? 4'b1001 : 4'b1000;
														assign node54966 = (inp[12]) ? node54968 : 4'b1000;
															assign node54968 = (inp[14]) ? node54972 : node54969;
																assign node54969 = (inp[8]) ? 4'b1000 : 4'b1001;
																assign node54972 = (inp[8]) ? 4'b1001 : 4'b1000;
													assign node54975 = (inp[14]) ? node54977 : 4'b1000;
														assign node54977 = (inp[8]) ? 4'b1000 : 4'b1001;
												assign node54980 = (inp[8]) ? node54984 : node54981;
													assign node54981 = (inp[7]) ? 4'b1001 : 4'b1000;
													assign node54984 = (inp[7]) ? 4'b1000 : 4'b1001;
											assign node54987 = (inp[5]) ? node55015 : node54988;
												assign node54988 = (inp[2]) ? node54998 : node54989;
													assign node54989 = (inp[8]) ? 4'b1000 : node54990;
														assign node54990 = (inp[14]) ? node54994 : node54991;
															assign node54991 = (inp[7]) ? 4'b1000 : 4'b1001;
															assign node54994 = (inp[7]) ? 4'b1001 : 4'b1000;
													assign node54998 = (inp[12]) ? node55008 : node54999;
														assign node54999 = (inp[14]) ? node55001 : 4'b1000;
															assign node55001 = (inp[7]) ? node55005 : node55002;
																assign node55002 = (inp[8]) ? 4'b1001 : 4'b1000;
																assign node55005 = (inp[8]) ? 4'b1000 : 4'b1001;
														assign node55008 = (inp[8]) ? node55012 : node55009;
															assign node55009 = (inp[7]) ? 4'b1001 : 4'b1000;
															assign node55012 = (inp[7]) ? 4'b1000 : 4'b1001;
												assign node55015 = (inp[12]) ? node55035 : node55016;
													assign node55016 = (inp[2]) ? node55022 : node55017;
														assign node55017 = (inp[14]) ? 4'b1011 : node55018;
															assign node55018 = (inp[7]) ? 4'b1011 : 4'b1010;
														assign node55022 = (inp[14]) ? node55030 : node55023;
															assign node55023 = (inp[8]) ? node55027 : node55024;
																assign node55024 = (inp[7]) ? 4'b1011 : 4'b1010;
																assign node55027 = (inp[7]) ? 4'b1010 : 4'b1011;
															assign node55030 = (inp[7]) ? node55032 : 4'b1010;
																assign node55032 = (inp[8]) ? 4'b1010 : 4'b1011;
													assign node55035 = (inp[14]) ? node55043 : node55036;
														assign node55036 = (inp[8]) ? 4'b1010 : node55037;
															assign node55037 = (inp[7]) ? 4'b1010 : node55038;
																assign node55038 = (inp[2]) ? 4'b1010 : 4'b1011;
														assign node55043 = (inp[7]) ? node55047 : node55044;
															assign node55044 = (inp[8]) ? 4'b1011 : 4'b1010;
															assign node55047 = (inp[8]) ? 4'b1010 : 4'b1011;
										assign node55050 = (inp[5]) ? node55074 : node55051;
											assign node55051 = (inp[8]) ? node55063 : node55052;
												assign node55052 = (inp[7]) ? node55058 : node55053;
													assign node55053 = (inp[2]) ? 4'b1010 : node55054;
														assign node55054 = (inp[14]) ? 4'b1010 : 4'b1011;
													assign node55058 = (inp[2]) ? 4'b1011 : node55059;
														assign node55059 = (inp[14]) ? 4'b1011 : 4'b1010;
												assign node55063 = (inp[7]) ? node55069 : node55064;
													assign node55064 = (inp[14]) ? 4'b1011 : node55065;
														assign node55065 = (inp[2]) ? 4'b1011 : 4'b1010;
													assign node55069 = (inp[14]) ? 4'b1010 : node55070;
														assign node55070 = (inp[2]) ? 4'b1010 : 4'b1011;
											assign node55074 = (inp[3]) ? node55096 : node55075;
												assign node55075 = (inp[7]) ? node55087 : node55076;
													assign node55076 = (inp[8]) ? node55082 : node55077;
														assign node55077 = (inp[2]) ? 4'b1010 : node55078;
															assign node55078 = (inp[12]) ? 4'b1011 : 4'b1010;
														assign node55082 = (inp[2]) ? 4'b1011 : node55083;
															assign node55083 = (inp[14]) ? 4'b1011 : 4'b1010;
													assign node55087 = (inp[8]) ? node55093 : node55088;
														assign node55088 = (inp[2]) ? 4'b1011 : node55089;
															assign node55089 = (inp[14]) ? 4'b1011 : 4'b1010;
														assign node55093 = (inp[2]) ? 4'b1010 : 4'b1011;
												assign node55096 = (inp[14]) ? node55106 : node55097;
													assign node55097 = (inp[8]) ? node55099 : 4'b1000;
														assign node55099 = (inp[2]) ? node55103 : node55100;
															assign node55100 = (inp[7]) ? 4'b1001 : 4'b1000;
															assign node55103 = (inp[7]) ? 4'b1000 : 4'b1001;
													assign node55106 = (inp[12]) ? node55116 : node55107;
														assign node55107 = (inp[2]) ? 4'b1000 : node55108;
															assign node55108 = (inp[8]) ? node55112 : node55109;
																assign node55109 = (inp[7]) ? 4'b1001 : 4'b1000;
																assign node55112 = (inp[7]) ? 4'b1000 : 4'b1001;
														assign node55116 = (inp[8]) ? node55118 : 4'b1001;
															assign node55118 = (inp[7]) ? 4'b1000 : 4'b1001;
								assign node55121 = (inp[0]) ? node55303 : node55122;
									assign node55122 = (inp[15]) ? node55222 : node55123;
										assign node55123 = (inp[5]) ? node55167 : node55124;
											assign node55124 = (inp[3]) ? node55144 : node55125;
												assign node55125 = (inp[7]) ? node55137 : node55126;
													assign node55126 = (inp[8]) ? node55132 : node55127;
														assign node55127 = (inp[2]) ? 4'b1110 : node55128;
															assign node55128 = (inp[14]) ? 4'b1110 : 4'b1111;
														assign node55132 = (inp[2]) ? 4'b1111 : node55133;
															assign node55133 = (inp[12]) ? 4'b1111 : 4'b1110;
													assign node55137 = (inp[8]) ? 4'b1110 : node55138;
														assign node55138 = (inp[14]) ? 4'b1111 : node55139;
															assign node55139 = (inp[2]) ? 4'b1111 : 4'b1110;
												assign node55144 = (inp[14]) ? node55160 : node55145;
													assign node55145 = (inp[7]) ? node55151 : node55146;
														assign node55146 = (inp[8]) ? 4'b1100 : node55147;
															assign node55147 = (inp[2]) ? 4'b1100 : 4'b1101;
														assign node55151 = (inp[12]) ? node55157 : node55152;
															assign node55152 = (inp[2]) ? 4'b1100 : node55153;
																assign node55153 = (inp[8]) ? 4'b1101 : 4'b1100;
															assign node55157 = (inp[2]) ? 4'b1101 : 4'b1100;
													assign node55160 = (inp[7]) ? node55164 : node55161;
														assign node55161 = (inp[8]) ? 4'b1101 : 4'b1100;
														assign node55164 = (inp[8]) ? 4'b1100 : 4'b1101;
											assign node55167 = (inp[2]) ? node55195 : node55168;
												assign node55168 = (inp[7]) ? node55180 : node55169;
													assign node55169 = (inp[12]) ? node55175 : node55170;
														assign node55170 = (inp[8]) ? node55172 : 4'b1100;
															assign node55172 = (inp[14]) ? 4'b1101 : 4'b1100;
														assign node55175 = (inp[14]) ? 4'b1100 : node55176;
															assign node55176 = (inp[8]) ? 4'b1100 : 4'b1101;
													assign node55180 = (inp[3]) ? node55188 : node55181;
														assign node55181 = (inp[8]) ? node55185 : node55182;
															assign node55182 = (inp[14]) ? 4'b1101 : 4'b1100;
															assign node55185 = (inp[14]) ? 4'b1100 : 4'b1101;
														assign node55188 = (inp[8]) ? node55192 : node55189;
															assign node55189 = (inp[14]) ? 4'b1101 : 4'b1100;
															assign node55192 = (inp[14]) ? 4'b1100 : 4'b1101;
												assign node55195 = (inp[14]) ? node55215 : node55196;
													assign node55196 = (inp[12]) ? node55208 : node55197;
														assign node55197 = (inp[3]) ? node55203 : node55198;
															assign node55198 = (inp[7]) ? 4'b1100 : node55199;
																assign node55199 = (inp[8]) ? 4'b1101 : 4'b1100;
															assign node55203 = (inp[7]) ? node55205 : 4'b1100;
																assign node55205 = (inp[8]) ? 4'b1100 : 4'b1101;
														assign node55208 = (inp[8]) ? node55212 : node55209;
															assign node55209 = (inp[7]) ? 4'b1101 : 4'b1100;
															assign node55212 = (inp[7]) ? 4'b1100 : 4'b1101;
													assign node55215 = (inp[8]) ? node55219 : node55216;
														assign node55216 = (inp[7]) ? 4'b1101 : 4'b1100;
														assign node55219 = (inp[7]) ? 4'b1100 : 4'b1101;
										assign node55222 = (inp[3]) ? node55280 : node55223;
											assign node55223 = (inp[5]) ? node55249 : node55224;
												assign node55224 = (inp[14]) ? node55238 : node55225;
													assign node55225 = (inp[2]) ? node55233 : node55226;
														assign node55226 = (inp[8]) ? node55230 : node55227;
															assign node55227 = (inp[7]) ? 4'b1100 : 4'b1101;
															assign node55230 = (inp[7]) ? 4'b1101 : 4'b1100;
														assign node55233 = (inp[12]) ? node55235 : 4'b1100;
															assign node55235 = (inp[7]) ? 4'b1101 : 4'b1100;
													assign node55238 = (inp[12]) ? node55244 : node55239;
														assign node55239 = (inp[8]) ? 4'b1101 : node55240;
															assign node55240 = (inp[7]) ? 4'b1101 : 4'b1100;
														assign node55244 = (inp[7]) ? node55246 : 4'b1101;
															assign node55246 = (inp[8]) ? 4'b1100 : 4'b1101;
												assign node55249 = (inp[2]) ? node55265 : node55250;
													assign node55250 = (inp[14]) ? node55256 : node55251;
														assign node55251 = (inp[7]) ? 4'b1110 : node55252;
															assign node55252 = (inp[8]) ? 4'b1110 : 4'b1111;
														assign node55256 = (inp[12]) ? node55262 : node55257;
															assign node55257 = (inp[8]) ? node55259 : 4'b1111;
																assign node55259 = (inp[7]) ? 4'b1110 : 4'b1111;
															assign node55262 = (inp[7]) ? 4'b1111 : 4'b1110;
													assign node55265 = (inp[14]) ? node55275 : node55266;
														assign node55266 = (inp[12]) ? node55270 : node55267;
															assign node55267 = (inp[7]) ? 4'b1110 : 4'b1111;
															assign node55270 = (inp[7]) ? 4'b1111 : node55271;
																assign node55271 = (inp[8]) ? 4'b1111 : 4'b1110;
														assign node55275 = (inp[8]) ? node55277 : 4'b1111;
															assign node55277 = (inp[7]) ? 4'b1110 : 4'b1111;
											assign node55280 = (inp[7]) ? node55292 : node55281;
												assign node55281 = (inp[8]) ? node55287 : node55282;
													assign node55282 = (inp[2]) ? 4'b1110 : node55283;
														assign node55283 = (inp[14]) ? 4'b1110 : 4'b1111;
													assign node55287 = (inp[14]) ? 4'b1111 : node55288;
														assign node55288 = (inp[2]) ? 4'b1111 : 4'b1110;
												assign node55292 = (inp[8]) ? node55298 : node55293;
													assign node55293 = (inp[2]) ? 4'b1111 : node55294;
														assign node55294 = (inp[14]) ? 4'b1111 : 4'b1110;
													assign node55298 = (inp[2]) ? 4'b1110 : node55299;
														assign node55299 = (inp[14]) ? 4'b1110 : 4'b1111;
									assign node55303 = (inp[15]) ? node55387 : node55304;
										assign node55304 = (inp[5]) ? node55364 : node55305;
											assign node55305 = (inp[3]) ? node55333 : node55306;
												assign node55306 = (inp[2]) ? node55326 : node55307;
													assign node55307 = (inp[8]) ? node55317 : node55308;
														assign node55308 = (inp[12]) ? 4'b1101 : node55309;
															assign node55309 = (inp[7]) ? node55313 : node55310;
																assign node55310 = (inp[14]) ? 4'b1100 : 4'b1101;
																assign node55313 = (inp[14]) ? 4'b1101 : 4'b1100;
														assign node55317 = (inp[12]) ? node55319 : 4'b1101;
															assign node55319 = (inp[7]) ? node55323 : node55320;
																assign node55320 = (inp[14]) ? 4'b1101 : 4'b1100;
																assign node55323 = (inp[14]) ? 4'b1100 : 4'b1101;
													assign node55326 = (inp[8]) ? node55330 : node55327;
														assign node55327 = (inp[7]) ? 4'b1101 : 4'b1100;
														assign node55330 = (inp[7]) ? 4'b1100 : 4'b1101;
												assign node55333 = (inp[14]) ? node55357 : node55334;
													assign node55334 = (inp[8]) ? node55344 : node55335;
														assign node55335 = (inp[12]) ? 4'b1111 : node55336;
															assign node55336 = (inp[2]) ? node55340 : node55337;
																assign node55337 = (inp[7]) ? 4'b1110 : 4'b1111;
																assign node55340 = (inp[7]) ? 4'b1111 : 4'b1110;
														assign node55344 = (inp[12]) ? node55352 : node55345;
															assign node55345 = (inp[2]) ? node55349 : node55346;
																assign node55346 = (inp[7]) ? 4'b1111 : 4'b1110;
																assign node55349 = (inp[7]) ? 4'b1110 : 4'b1111;
															assign node55352 = (inp[2]) ? 4'b1110 : node55353;
																assign node55353 = (inp[7]) ? 4'b1111 : 4'b1110;
													assign node55357 = (inp[8]) ? node55361 : node55358;
														assign node55358 = (inp[7]) ? 4'b1111 : 4'b1110;
														assign node55361 = (inp[7]) ? 4'b1110 : 4'b1111;
											assign node55364 = (inp[7]) ? node55376 : node55365;
												assign node55365 = (inp[8]) ? node55371 : node55366;
													assign node55366 = (inp[14]) ? 4'b1110 : node55367;
														assign node55367 = (inp[2]) ? 4'b1110 : 4'b1111;
													assign node55371 = (inp[2]) ? 4'b1111 : node55372;
														assign node55372 = (inp[14]) ? 4'b1111 : 4'b1110;
												assign node55376 = (inp[8]) ? node55382 : node55377;
													assign node55377 = (inp[14]) ? 4'b1111 : node55378;
														assign node55378 = (inp[2]) ? 4'b1111 : 4'b1110;
													assign node55382 = (inp[2]) ? 4'b1110 : node55383;
														assign node55383 = (inp[14]) ? 4'b1110 : 4'b1111;
										assign node55387 = (inp[3]) ? node55453 : node55388;
											assign node55388 = (inp[5]) ? node55426 : node55389;
												assign node55389 = (inp[12]) ? node55407 : node55390;
													assign node55390 = (inp[2]) ? node55402 : node55391;
														assign node55391 = (inp[7]) ? node55397 : node55392;
															assign node55392 = (inp[8]) ? 4'b1110 : node55393;
																assign node55393 = (inp[14]) ? 4'b1110 : 4'b1111;
															assign node55397 = (inp[8]) ? node55399 : 4'b1111;
																assign node55399 = (inp[14]) ? 4'b1110 : 4'b1111;
														assign node55402 = (inp[8]) ? 4'b1111 : node55403;
															assign node55403 = (inp[7]) ? 4'b1111 : 4'b1110;
													assign node55407 = (inp[8]) ? node55417 : node55408;
														assign node55408 = (inp[14]) ? 4'b1110 : node55409;
															assign node55409 = (inp[7]) ? node55413 : node55410;
																assign node55410 = (inp[2]) ? 4'b1110 : 4'b1111;
																assign node55413 = (inp[2]) ? 4'b1111 : 4'b1110;
														assign node55417 = (inp[7]) ? node55423 : node55418;
															assign node55418 = (inp[2]) ? 4'b1111 : node55419;
																assign node55419 = (inp[14]) ? 4'b1111 : 4'b1110;
															assign node55423 = (inp[2]) ? 4'b1110 : 4'b1111;
												assign node55426 = (inp[2]) ? node55442 : node55427;
													assign node55427 = (inp[7]) ? node55435 : node55428;
														assign node55428 = (inp[14]) ? node55432 : node55429;
															assign node55429 = (inp[8]) ? 4'b1100 : 4'b1101;
															assign node55432 = (inp[8]) ? 4'b1101 : 4'b1100;
														assign node55435 = (inp[8]) ? node55439 : node55436;
															assign node55436 = (inp[14]) ? 4'b1101 : 4'b1100;
															assign node55439 = (inp[14]) ? 4'b1100 : 4'b1101;
													assign node55442 = (inp[14]) ? node55444 : 4'b1101;
														assign node55444 = (inp[12]) ? 4'b1101 : node55445;
															assign node55445 = (inp[8]) ? node55449 : node55446;
																assign node55446 = (inp[7]) ? 4'b1101 : 4'b1100;
																assign node55449 = (inp[7]) ? 4'b1100 : 4'b1101;
											assign node55453 = (inp[2]) ? node55483 : node55454;
												assign node55454 = (inp[12]) ? node55464 : node55455;
													assign node55455 = (inp[14]) ? 4'b1101 : node55456;
														assign node55456 = (inp[8]) ? node55460 : node55457;
															assign node55457 = (inp[7]) ? 4'b1100 : 4'b1101;
															assign node55460 = (inp[7]) ? 4'b1101 : 4'b1100;
													assign node55464 = (inp[7]) ? node55476 : node55465;
														assign node55465 = (inp[5]) ? node55471 : node55466;
															assign node55466 = (inp[8]) ? node55468 : 4'b1101;
																assign node55468 = (inp[14]) ? 4'b1101 : 4'b1100;
															assign node55471 = (inp[14]) ? node55473 : 4'b1101;
																assign node55473 = (inp[8]) ? 4'b1101 : 4'b1100;
														assign node55476 = (inp[8]) ? node55480 : node55477;
															assign node55477 = (inp[14]) ? 4'b1101 : 4'b1100;
															assign node55480 = (inp[14]) ? 4'b1100 : 4'b1101;
												assign node55483 = (inp[14]) ? node55495 : node55484;
													assign node55484 = (inp[5]) ? node55490 : node55485;
														assign node55485 = (inp[7]) ? 4'b1100 : node55486;
															assign node55486 = (inp[8]) ? 4'b1101 : 4'b1100;
														assign node55490 = (inp[7]) ? 4'b1101 : node55491;
															assign node55491 = (inp[8]) ? 4'b1101 : 4'b1100;
													assign node55495 = (inp[5]) ? node55503 : node55496;
														assign node55496 = (inp[7]) ? node55500 : node55497;
															assign node55497 = (inp[8]) ? 4'b1101 : 4'b1100;
															assign node55500 = (inp[8]) ? 4'b1100 : 4'b1101;
														assign node55503 = (inp[12]) ? node55509 : node55504;
															assign node55504 = (inp[7]) ? node55506 : 4'b1100;
																assign node55506 = (inp[8]) ? 4'b1100 : 4'b1101;
															assign node55509 = (inp[7]) ? 4'b1100 : node55510;
																assign node55510 = (inp[8]) ? 4'b1101 : 4'b1100;
							assign node55514 = (inp[4]) ? node55998 : node55515;
								assign node55515 = (inp[3]) ? node55801 : node55516;
									assign node55516 = (inp[15]) ? node55650 : node55517;
										assign node55517 = (inp[2]) ? node55587 : node55518;
											assign node55518 = (inp[12]) ? node55552 : node55519;
												assign node55519 = (inp[7]) ? node55535 : node55520;
													assign node55520 = (inp[14]) ? node55528 : node55521;
														assign node55521 = (inp[8]) ? 4'b1110 : node55522;
															assign node55522 = (inp[5]) ? node55524 : 4'b1111;
																assign node55524 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node55528 = (inp[8]) ? node55530 : 4'b1110;
															assign node55530 = (inp[0]) ? 4'b1101 : node55531;
																assign node55531 = (inp[5]) ? 4'b1101 : 4'b1111;
													assign node55535 = (inp[14]) ? node55543 : node55536;
														assign node55536 = (inp[8]) ? node55538 : 4'b1100;
															assign node55538 = (inp[0]) ? node55540 : 4'b1101;
																assign node55540 = (inp[5]) ? 4'b1111 : 4'b1101;
														assign node55543 = (inp[8]) ? node55549 : node55544;
															assign node55544 = (inp[5]) ? node55546 : 4'b1111;
																assign node55546 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node55549 = (inp[0]) ? 4'b1100 : 4'b1110;
												assign node55552 = (inp[14]) ? node55568 : node55553;
													assign node55553 = (inp[0]) ? node55561 : node55554;
														assign node55554 = (inp[5]) ? 4'b1100 : node55555;
															assign node55555 = (inp[8]) ? node55557 : 4'b1110;
																assign node55557 = (inp[7]) ? 4'b1111 : 4'b1110;
														assign node55561 = (inp[5]) ? node55563 : 4'b1100;
															assign node55563 = (inp[7]) ? node55565 : 4'b1111;
																assign node55565 = (inp[8]) ? 4'b1111 : 4'b1110;
													assign node55568 = (inp[0]) ? node55574 : node55569;
														assign node55569 = (inp[8]) ? 4'b1100 : node55570;
															assign node55570 = (inp[7]) ? 4'b1101 : 4'b1100;
														assign node55574 = (inp[5]) ? node55580 : node55575;
															assign node55575 = (inp[8]) ? 4'b1100 : node55576;
																assign node55576 = (inp[7]) ? 4'b1101 : 4'b1100;
															assign node55580 = (inp[7]) ? node55584 : node55581;
																assign node55581 = (inp[8]) ? 4'b1111 : 4'b1110;
																assign node55584 = (inp[8]) ? 4'b1110 : 4'b1111;
											assign node55587 = (inp[14]) ? node55619 : node55588;
												assign node55588 = (inp[5]) ? node55608 : node55589;
													assign node55589 = (inp[0]) ? node55595 : node55590;
														assign node55590 = (inp[8]) ? node55592 : 4'b1111;
															assign node55592 = (inp[7]) ? 4'b1110 : 4'b1111;
														assign node55595 = (inp[12]) ? node55603 : node55596;
															assign node55596 = (inp[7]) ? node55600 : node55597;
																assign node55597 = (inp[8]) ? 4'b1101 : 4'b1100;
																assign node55600 = (inp[8]) ? 4'b1100 : 4'b1101;
															assign node55603 = (inp[8]) ? 4'b1101 : node55604;
																assign node55604 = (inp[7]) ? 4'b1101 : 4'b1100;
													assign node55608 = (inp[0]) ? node55616 : node55609;
														assign node55609 = (inp[8]) ? node55613 : node55610;
															assign node55610 = (inp[7]) ? 4'b1101 : 4'b1100;
															assign node55613 = (inp[7]) ? 4'b1100 : 4'b1101;
														assign node55616 = (inp[7]) ? 4'b1111 : 4'b1110;
												assign node55619 = (inp[7]) ? node55633 : node55620;
													assign node55620 = (inp[8]) ? node55622 : 4'b1110;
														assign node55622 = (inp[12]) ? node55628 : node55623;
															assign node55623 = (inp[0]) ? 4'b1111 : node55624;
																assign node55624 = (inp[5]) ? 4'b1101 : 4'b1111;
															assign node55628 = (inp[5]) ? 4'b1111 : node55629;
																assign node55629 = (inp[0]) ? 4'b1101 : 4'b1111;
													assign node55633 = (inp[8]) ? node55641 : node55634;
														assign node55634 = (inp[0]) ? node55638 : node55635;
															assign node55635 = (inp[5]) ? 4'b1101 : 4'b1111;
															assign node55638 = (inp[5]) ? 4'b1111 : 4'b1101;
														assign node55641 = (inp[12]) ? node55643 : 4'b1100;
															assign node55643 = (inp[0]) ? node55647 : node55644;
																assign node55644 = (inp[5]) ? 4'b1100 : 4'b1110;
																assign node55647 = (inp[5]) ? 4'b1110 : 4'b1100;
										assign node55650 = (inp[12]) ? node55724 : node55651;
											assign node55651 = (inp[2]) ? node55697 : node55652;
												assign node55652 = (inp[8]) ? node55672 : node55653;
													assign node55653 = (inp[5]) ? node55663 : node55654;
														assign node55654 = (inp[0]) ? node55658 : node55655;
															assign node55655 = (inp[14]) ? 4'b1101 : 4'b1100;
															assign node55658 = (inp[14]) ? node55660 : 4'b1110;
																assign node55660 = (inp[7]) ? 4'b1111 : 4'b1110;
														assign node55663 = (inp[0]) ? 4'b1101 : node55664;
															assign node55664 = (inp[7]) ? node55668 : node55665;
																assign node55665 = (inp[14]) ? 4'b1110 : 4'b1111;
																assign node55668 = (inp[14]) ? 4'b1111 : 4'b1110;
													assign node55672 = (inp[0]) ? node55682 : node55673;
														assign node55673 = (inp[5]) ? node55675 : 4'b1101;
															assign node55675 = (inp[14]) ? node55679 : node55676;
																assign node55676 = (inp[7]) ? 4'b1111 : 4'b1110;
																assign node55679 = (inp[7]) ? 4'b1110 : 4'b1111;
														assign node55682 = (inp[5]) ? node55690 : node55683;
															assign node55683 = (inp[14]) ? node55687 : node55684;
																assign node55684 = (inp[7]) ? 4'b1111 : 4'b1110;
																assign node55687 = (inp[7]) ? 4'b1110 : 4'b1111;
															assign node55690 = (inp[14]) ? node55694 : node55691;
																assign node55691 = (inp[7]) ? 4'b1101 : 4'b1100;
																assign node55694 = (inp[7]) ? 4'b1100 : 4'b1101;
												assign node55697 = (inp[0]) ? node55711 : node55698;
													assign node55698 = (inp[5]) ? node55704 : node55699;
														assign node55699 = (inp[7]) ? node55701 : 4'b1100;
															assign node55701 = (inp[8]) ? 4'b1100 : 4'b1101;
														assign node55704 = (inp[8]) ? node55708 : node55705;
															assign node55705 = (inp[7]) ? 4'b1111 : 4'b1110;
															assign node55708 = (inp[7]) ? 4'b1110 : 4'b1111;
													assign node55711 = (inp[5]) ? node55719 : node55712;
														assign node55712 = (inp[7]) ? node55716 : node55713;
															assign node55713 = (inp[8]) ? 4'b1111 : 4'b1110;
															assign node55716 = (inp[8]) ? 4'b1110 : 4'b1111;
														assign node55719 = (inp[7]) ? 4'b1100 : node55720;
															assign node55720 = (inp[8]) ? 4'b1101 : 4'b1100;
											assign node55724 = (inp[7]) ? node55772 : node55725;
												assign node55725 = (inp[8]) ? node55743 : node55726;
													assign node55726 = (inp[2]) ? node55736 : node55727;
														assign node55727 = (inp[14]) ? node55733 : node55728;
															assign node55728 = (inp[5]) ? 4'b1111 : node55729;
																assign node55729 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node55733 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node55736 = (inp[5]) ? node55740 : node55737;
															assign node55737 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node55740 = (inp[0]) ? 4'b1100 : 4'b1110;
													assign node55743 = (inp[14]) ? node55757 : node55744;
														assign node55744 = (inp[2]) ? node55752 : node55745;
															assign node55745 = (inp[5]) ? node55749 : node55746;
																assign node55746 = (inp[0]) ? 4'b1110 : 4'b1100;
																assign node55749 = (inp[0]) ? 4'b1100 : 4'b1110;
															assign node55752 = (inp[0]) ? 4'b1101 : node55753;
																assign node55753 = (inp[5]) ? 4'b1111 : 4'b1101;
														assign node55757 = (inp[2]) ? node55765 : node55758;
															assign node55758 = (inp[0]) ? node55762 : node55759;
																assign node55759 = (inp[5]) ? 4'b1111 : 4'b1101;
																assign node55762 = (inp[5]) ? 4'b1101 : 4'b1111;
															assign node55765 = (inp[0]) ? node55769 : node55766;
																assign node55766 = (inp[5]) ? 4'b1111 : 4'b1101;
																assign node55769 = (inp[5]) ? 4'b1101 : 4'b1111;
												assign node55772 = (inp[8]) ? node55780 : node55773;
													assign node55773 = (inp[14]) ? 4'b1101 : node55774;
														assign node55774 = (inp[2]) ? 4'b1111 : node55775;
															assign node55775 = (inp[0]) ? 4'b1110 : 4'b1100;
													assign node55780 = (inp[14]) ? node55790 : node55781;
														assign node55781 = (inp[2]) ? node55787 : node55782;
															assign node55782 = (inp[0]) ? node55784 : 4'b1101;
																assign node55784 = (inp[5]) ? 4'b1101 : 4'b1111;
															assign node55787 = (inp[0]) ? 4'b1100 : 4'b1110;
														assign node55790 = (inp[2]) ? node55796 : node55791;
															assign node55791 = (inp[5]) ? 4'b1110 : node55792;
																assign node55792 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node55796 = (inp[0]) ? node55798 : 4'b1100;
																assign node55798 = (inp[5]) ? 4'b1100 : 4'b1110;
									assign node55801 = (inp[2]) ? node55921 : node55802;
										assign node55802 = (inp[12]) ? node55864 : node55803;
											assign node55803 = (inp[8]) ? node55835 : node55804;
												assign node55804 = (inp[7]) ? node55822 : node55805;
													assign node55805 = (inp[14]) ? node55815 : node55806;
														assign node55806 = (inp[5]) ? node55810 : node55807;
															assign node55807 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node55810 = (inp[15]) ? 4'b1101 : node55811;
																assign node55811 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node55815 = (inp[15]) ? node55819 : node55816;
															assign node55816 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node55819 = (inp[0]) ? 4'b1100 : 4'b1110;
													assign node55822 = (inp[14]) ? node55828 : node55823;
														assign node55823 = (inp[5]) ? node55825 : 4'b1100;
															assign node55825 = (inp[15]) ? 4'b1100 : 4'b1110;
														assign node55828 = (inp[0]) ? node55832 : node55829;
															assign node55829 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node55832 = (inp[15]) ? 4'b1101 : 4'b1111;
												assign node55835 = (inp[14]) ? node55849 : node55836;
													assign node55836 = (inp[7]) ? node55842 : node55837;
														assign node55837 = (inp[0]) ? 4'b1110 : node55838;
															assign node55838 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node55842 = (inp[15]) ? node55846 : node55843;
															assign node55843 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node55846 = (inp[0]) ? 4'b1101 : 4'b1111;
													assign node55849 = (inp[7]) ? node55857 : node55850;
														assign node55850 = (inp[15]) ? node55854 : node55851;
															assign node55851 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node55854 = (inp[0]) ? 4'b1101 : 4'b1111;
														assign node55857 = (inp[5]) ? 4'b1100 : node55858;
															assign node55858 = (inp[0]) ? node55860 : 4'b1100;
																assign node55860 = (inp[15]) ? 4'b1100 : 4'b1110;
											assign node55864 = (inp[7]) ? node55888 : node55865;
												assign node55865 = (inp[15]) ? node55875 : node55866;
													assign node55866 = (inp[0]) ? node55870 : node55867;
														assign node55867 = (inp[14]) ? 4'b1101 : 4'b1100;
														assign node55870 = (inp[14]) ? 4'b1110 : node55871;
															assign node55871 = (inp[8]) ? 4'b1110 : 4'b1111;
													assign node55875 = (inp[0]) ? node55881 : node55876;
														assign node55876 = (inp[8]) ? node55878 : 4'b1110;
															assign node55878 = (inp[14]) ? 4'b1111 : 4'b1110;
														assign node55881 = (inp[8]) ? node55885 : node55882;
															assign node55882 = (inp[14]) ? 4'b1100 : 4'b1101;
															assign node55885 = (inp[14]) ? 4'b1101 : 4'b1100;
												assign node55888 = (inp[15]) ? node55908 : node55889;
													assign node55889 = (inp[0]) ? node55895 : node55890;
														assign node55890 = (inp[14]) ? node55892 : 4'b1101;
															assign node55892 = (inp[8]) ? 4'b1100 : 4'b1101;
														assign node55895 = (inp[5]) ? node55901 : node55896;
															assign node55896 = (inp[8]) ? node55898 : 4'b1111;
																assign node55898 = (inp[14]) ? 4'b1110 : 4'b1111;
															assign node55901 = (inp[14]) ? node55905 : node55902;
																assign node55902 = (inp[8]) ? 4'b1111 : 4'b1110;
																assign node55905 = (inp[8]) ? 4'b1110 : 4'b1111;
													assign node55908 = (inp[0]) ? node55916 : node55909;
														assign node55909 = (inp[8]) ? node55913 : node55910;
															assign node55910 = (inp[14]) ? 4'b1111 : 4'b1110;
															assign node55913 = (inp[14]) ? 4'b1110 : 4'b1111;
														assign node55916 = (inp[5]) ? node55918 : 4'b1100;
															assign node55918 = (inp[8]) ? 4'b1100 : 4'b1101;
										assign node55921 = (inp[7]) ? node55951 : node55922;
											assign node55922 = (inp[8]) ? node55938 : node55923;
												assign node55923 = (inp[14]) ? node55931 : node55924;
													assign node55924 = (inp[15]) ? node55928 : node55925;
														assign node55925 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node55928 = (inp[0]) ? 4'b1100 : 4'b1110;
													assign node55931 = (inp[0]) ? node55935 : node55932;
														assign node55932 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node55935 = (inp[15]) ? 4'b1100 : 4'b1110;
												assign node55938 = (inp[14]) ? node55946 : node55939;
													assign node55939 = (inp[0]) ? node55943 : node55940;
														assign node55940 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node55943 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node55946 = (inp[15]) ? 4'b1111 : node55947;
														assign node55947 = (inp[0]) ? 4'b1111 : 4'b1101;
											assign node55951 = (inp[8]) ? node55967 : node55952;
												assign node55952 = (inp[14]) ? node55960 : node55953;
													assign node55953 = (inp[15]) ? node55957 : node55954;
														assign node55954 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node55957 = (inp[0]) ? 4'b1101 : 4'b1111;
													assign node55960 = (inp[15]) ? node55964 : node55961;
														assign node55961 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node55964 = (inp[0]) ? 4'b1101 : 4'b1111;
												assign node55967 = (inp[12]) ? node55991 : node55968;
													assign node55968 = (inp[14]) ? node55984 : node55969;
														assign node55969 = (inp[5]) ? node55977 : node55970;
															assign node55970 = (inp[15]) ? node55974 : node55971;
																assign node55971 = (inp[0]) ? 4'b1110 : 4'b1100;
																assign node55974 = (inp[0]) ? 4'b1100 : 4'b1110;
															assign node55977 = (inp[15]) ? node55981 : node55978;
																assign node55978 = (inp[0]) ? 4'b1110 : 4'b1100;
																assign node55981 = (inp[0]) ? 4'b1100 : 4'b1110;
														assign node55984 = (inp[0]) ? node55988 : node55985;
															assign node55985 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node55988 = (inp[15]) ? 4'b1100 : 4'b1110;
													assign node55991 = (inp[15]) ? node55995 : node55992;
														assign node55992 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node55995 = (inp[0]) ? 4'b1100 : 4'b1110;
								assign node55998 = (inp[3]) ? node56298 : node55999;
									assign node55999 = (inp[12]) ? node56133 : node56000;
										assign node56000 = (inp[2]) ? node56080 : node56001;
											assign node56001 = (inp[14]) ? node56045 : node56002;
												assign node56002 = (inp[15]) ? node56018 : node56003;
													assign node56003 = (inp[8]) ? node56015 : node56004;
														assign node56004 = (inp[7]) ? node56010 : node56005;
															assign node56005 = (inp[0]) ? node56007 : 4'b1011;
																assign node56007 = (inp[5]) ? 4'b1011 : 4'b1001;
															assign node56010 = (inp[0]) ? 4'b1000 : node56011;
																assign node56011 = (inp[5]) ? 4'b1000 : 4'b1010;
														assign node56015 = (inp[7]) ? 4'b1011 : 4'b1010;
													assign node56018 = (inp[7]) ? node56030 : node56019;
														assign node56019 = (inp[8]) ? node56025 : node56020;
															assign node56020 = (inp[5]) ? 4'b1001 : node56021;
																assign node56021 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node56025 = (inp[0]) ? 4'b1000 : node56026;
																assign node56026 = (inp[5]) ? 4'b1010 : 4'b1000;
														assign node56030 = (inp[8]) ? node56038 : node56031;
															assign node56031 = (inp[5]) ? node56035 : node56032;
																assign node56032 = (inp[0]) ? 4'b1010 : 4'b1000;
																assign node56035 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node56038 = (inp[0]) ? node56042 : node56039;
																assign node56039 = (inp[5]) ? 4'b1011 : 4'b1001;
																assign node56042 = (inp[5]) ? 4'b1001 : 4'b1011;
												assign node56045 = (inp[5]) ? node56063 : node56046;
													assign node56046 = (inp[15]) ? node56054 : node56047;
														assign node56047 = (inp[0]) ? node56049 : 4'b1010;
															assign node56049 = (inp[7]) ? 4'b1000 : node56050;
																assign node56050 = (inp[8]) ? 4'b1001 : 4'b1000;
														assign node56054 = (inp[0]) ? node56058 : node56055;
															assign node56055 = (inp[7]) ? 4'b1001 : 4'b1000;
															assign node56058 = (inp[7]) ? 4'b1010 : node56059;
																assign node56059 = (inp[8]) ? 4'b1011 : 4'b1010;
													assign node56063 = (inp[7]) ? node56069 : node56064;
														assign node56064 = (inp[8]) ? 4'b1001 : node56065;
															assign node56065 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node56069 = (inp[8]) ? node56075 : node56070;
															assign node56070 = (inp[15]) ? 4'b1001 : node56071;
																assign node56071 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node56075 = (inp[0]) ? node56077 : 4'b1010;
																assign node56077 = (inp[15]) ? 4'b1000 : 4'b1010;
											assign node56080 = (inp[8]) ? node56108 : node56081;
												assign node56081 = (inp[7]) ? node56093 : node56082;
													assign node56082 = (inp[5]) ? node56088 : node56083;
														assign node56083 = (inp[15]) ? node56085 : 4'b1000;
															assign node56085 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node56088 = (inp[14]) ? 4'b1010 : node56089;
															assign node56089 = (inp[15]) ? 4'b1010 : 4'b1000;
													assign node56093 = (inp[15]) ? node56101 : node56094;
														assign node56094 = (inp[5]) ? node56098 : node56095;
															assign node56095 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node56098 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node56101 = (inp[5]) ? node56105 : node56102;
															assign node56102 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node56105 = (inp[0]) ? 4'b1001 : 4'b1011;
												assign node56108 = (inp[7]) ? node56120 : node56109;
													assign node56109 = (inp[15]) ? node56117 : node56110;
														assign node56110 = (inp[5]) ? node56114 : node56111;
															assign node56111 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node56114 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node56117 = (inp[5]) ? 4'b1011 : 4'b1001;
													assign node56120 = (inp[5]) ? node56130 : node56121;
														assign node56121 = (inp[14]) ? node56123 : 4'b1000;
															assign node56123 = (inp[0]) ? node56127 : node56124;
																assign node56124 = (inp[15]) ? 4'b1000 : 4'b1010;
																assign node56127 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node56130 = (inp[14]) ? 4'b1000 : 4'b1010;
										assign node56133 = (inp[0]) ? node56225 : node56134;
											assign node56134 = (inp[2]) ? node56180 : node56135;
												assign node56135 = (inp[14]) ? node56157 : node56136;
													assign node56136 = (inp[7]) ? node56146 : node56137;
														assign node56137 = (inp[8]) ? node56139 : 4'b1001;
															assign node56139 = (inp[5]) ? node56143 : node56140;
																assign node56140 = (inp[15]) ? 4'b1000 : 4'b1010;
																assign node56143 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node56146 = (inp[8]) ? node56152 : node56147;
															assign node56147 = (inp[15]) ? 4'b1010 : node56148;
																assign node56148 = (inp[5]) ? 4'b1000 : 4'b1010;
															assign node56152 = (inp[5]) ? node56154 : 4'b1001;
																assign node56154 = (inp[15]) ? 4'b1011 : 4'b1001;
													assign node56157 = (inp[15]) ? node56167 : node56158;
														assign node56158 = (inp[5]) ? 4'b1001 : node56159;
															assign node56159 = (inp[7]) ? node56163 : node56160;
																assign node56160 = (inp[8]) ? 4'b1011 : 4'b1010;
																assign node56163 = (inp[8]) ? 4'b1010 : 4'b1011;
														assign node56167 = (inp[5]) ? node56175 : node56168;
															assign node56168 = (inp[7]) ? node56172 : node56169;
																assign node56169 = (inp[8]) ? 4'b1001 : 4'b1000;
																assign node56172 = (inp[8]) ? 4'b1000 : 4'b1001;
															assign node56175 = (inp[7]) ? 4'b1010 : node56176;
																assign node56176 = (inp[8]) ? 4'b1011 : 4'b1010;
												assign node56180 = (inp[14]) ? node56198 : node56181;
													assign node56181 = (inp[8]) ? node56189 : node56182;
														assign node56182 = (inp[7]) ? 4'b1011 : node56183;
															assign node56183 = (inp[5]) ? node56185 : 4'b1010;
																assign node56185 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node56189 = (inp[7]) ? node56195 : node56190;
															assign node56190 = (inp[15]) ? 4'b1011 : node56191;
																assign node56191 = (inp[5]) ? 4'b1001 : 4'b1011;
															assign node56195 = (inp[15]) ? 4'b1000 : 4'b1010;
													assign node56198 = (inp[7]) ? node56210 : node56199;
														assign node56199 = (inp[8]) ? node56205 : node56200;
															assign node56200 = (inp[5]) ? node56202 : 4'b1010;
																assign node56202 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node56205 = (inp[15]) ? node56207 : 4'b1011;
																assign node56207 = (inp[5]) ? 4'b1011 : 4'b1001;
														assign node56210 = (inp[8]) ? node56218 : node56211;
															assign node56211 = (inp[5]) ? node56215 : node56212;
																assign node56212 = (inp[15]) ? 4'b1001 : 4'b1011;
																assign node56215 = (inp[15]) ? 4'b1011 : 4'b1001;
															assign node56218 = (inp[15]) ? node56222 : node56219;
																assign node56219 = (inp[5]) ? 4'b1000 : 4'b1010;
																assign node56222 = (inp[5]) ? 4'b1010 : 4'b1000;
											assign node56225 = (inp[2]) ? node56259 : node56226;
												assign node56226 = (inp[15]) ? node56244 : node56227;
													assign node56227 = (inp[5]) ? node56231 : node56228;
														assign node56228 = (inp[7]) ? 4'b1001 : 4'b1000;
														assign node56231 = (inp[8]) ? node56237 : node56232;
															assign node56232 = (inp[14]) ? node56234 : 4'b1010;
																assign node56234 = (inp[7]) ? 4'b1011 : 4'b1010;
															assign node56237 = (inp[7]) ? node56241 : node56238;
																assign node56238 = (inp[14]) ? 4'b1011 : 4'b1010;
																assign node56241 = (inp[14]) ? 4'b1010 : 4'b1011;
													assign node56244 = (inp[5]) ? 4'b1001 : node56245;
														assign node56245 = (inp[7]) ? node56253 : node56246;
															assign node56246 = (inp[8]) ? node56250 : node56247;
																assign node56247 = (inp[14]) ? 4'b1010 : 4'b1011;
																assign node56250 = (inp[14]) ? 4'b1011 : 4'b1010;
															assign node56253 = (inp[14]) ? node56255 : 4'b1011;
																assign node56255 = (inp[8]) ? 4'b1010 : 4'b1011;
												assign node56259 = (inp[8]) ? node56281 : node56260;
													assign node56260 = (inp[7]) ? node56268 : node56261;
														assign node56261 = (inp[5]) ? node56265 : node56262;
															assign node56262 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node56265 = (inp[15]) ? 4'b1000 : 4'b1010;
														assign node56268 = (inp[14]) ? node56276 : node56269;
															assign node56269 = (inp[15]) ? node56273 : node56270;
																assign node56270 = (inp[5]) ? 4'b1011 : 4'b1001;
																assign node56273 = (inp[5]) ? 4'b1001 : 4'b1011;
															assign node56276 = (inp[15]) ? 4'b1001 : node56277;
																assign node56277 = (inp[5]) ? 4'b1011 : 4'b1001;
													assign node56281 = (inp[7]) ? node56291 : node56282;
														assign node56282 = (inp[14]) ? node56284 : 4'b1011;
															assign node56284 = (inp[15]) ? node56288 : node56285;
																assign node56285 = (inp[5]) ? 4'b1011 : 4'b1001;
																assign node56288 = (inp[5]) ? 4'b1001 : 4'b1011;
														assign node56291 = (inp[15]) ? node56295 : node56292;
															assign node56292 = (inp[5]) ? 4'b1010 : 4'b1000;
															assign node56295 = (inp[5]) ? 4'b1000 : 4'b1010;
									assign node56298 = (inp[0]) ? node56384 : node56299;
										assign node56299 = (inp[15]) ? node56323 : node56300;
											assign node56300 = (inp[8]) ? node56312 : node56301;
												assign node56301 = (inp[7]) ? node56307 : node56302;
													assign node56302 = (inp[14]) ? 4'b1000 : node56303;
														assign node56303 = (inp[2]) ? 4'b1000 : 4'b1001;
													assign node56307 = (inp[2]) ? 4'b1001 : node56308;
														assign node56308 = (inp[14]) ? 4'b1001 : 4'b1000;
												assign node56312 = (inp[7]) ? node56318 : node56313;
													assign node56313 = (inp[2]) ? 4'b1001 : node56314;
														assign node56314 = (inp[14]) ? 4'b1001 : 4'b1000;
													assign node56318 = (inp[2]) ? 4'b1000 : node56319;
														assign node56319 = (inp[14]) ? 4'b1000 : 4'b1001;
											assign node56323 = (inp[2]) ? node56361 : node56324;
												assign node56324 = (inp[5]) ? node56338 : node56325;
													assign node56325 = (inp[8]) ? node56333 : node56326;
														assign node56326 = (inp[7]) ? node56330 : node56327;
															assign node56327 = (inp[14]) ? 4'b1010 : 4'b1011;
															assign node56330 = (inp[14]) ? 4'b1011 : 4'b1010;
														assign node56333 = (inp[7]) ? node56335 : 4'b1011;
															assign node56335 = (inp[14]) ? 4'b1010 : 4'b1011;
													assign node56338 = (inp[8]) ? node56346 : node56339;
														assign node56339 = (inp[7]) ? node56343 : node56340;
															assign node56340 = (inp[14]) ? 4'b1010 : 4'b1011;
															assign node56343 = (inp[14]) ? 4'b1011 : 4'b1010;
														assign node56346 = (inp[12]) ? node56354 : node56347;
															assign node56347 = (inp[7]) ? node56351 : node56348;
																assign node56348 = (inp[14]) ? 4'b1011 : 4'b1010;
																assign node56351 = (inp[14]) ? 4'b1010 : 4'b1011;
															assign node56354 = (inp[14]) ? node56358 : node56355;
																assign node56355 = (inp[7]) ? 4'b1011 : 4'b1010;
																assign node56358 = (inp[7]) ? 4'b1010 : 4'b1011;
												assign node56361 = (inp[14]) ? node56377 : node56362;
													assign node56362 = (inp[5]) ? node56370 : node56363;
														assign node56363 = (inp[7]) ? node56367 : node56364;
															assign node56364 = (inp[8]) ? 4'b1011 : 4'b1010;
															assign node56367 = (inp[8]) ? 4'b1010 : 4'b1011;
														assign node56370 = (inp[7]) ? node56374 : node56371;
															assign node56371 = (inp[8]) ? 4'b1011 : 4'b1010;
															assign node56374 = (inp[8]) ? 4'b1010 : 4'b1011;
													assign node56377 = (inp[7]) ? node56381 : node56378;
														assign node56378 = (inp[8]) ? 4'b1011 : 4'b1010;
														assign node56381 = (inp[8]) ? 4'b1010 : 4'b1011;
										assign node56384 = (inp[15]) ? node56424 : node56385;
											assign node56385 = (inp[5]) ? node56409 : node56386;
												assign node56386 = (inp[8]) ? node56398 : node56387;
													assign node56387 = (inp[7]) ? node56393 : node56388;
														assign node56388 = (inp[2]) ? 4'b1010 : node56389;
															assign node56389 = (inp[14]) ? 4'b1010 : 4'b1011;
														assign node56393 = (inp[14]) ? 4'b1011 : node56394;
															assign node56394 = (inp[2]) ? 4'b1011 : 4'b1010;
													assign node56398 = (inp[12]) ? node56406 : node56399;
														assign node56399 = (inp[14]) ? 4'b1011 : node56400;
															assign node56400 = (inp[2]) ? 4'b1011 : node56401;
																assign node56401 = (inp[7]) ? 4'b1011 : 4'b1010;
														assign node56406 = (inp[2]) ? 4'b1010 : 4'b1011;
												assign node56409 = (inp[8]) ? node56419 : node56410;
													assign node56410 = (inp[2]) ? node56416 : node56411;
														assign node56411 = (inp[7]) ? node56413 : 4'b1011;
															assign node56413 = (inp[14]) ? 4'b1011 : 4'b1010;
														assign node56416 = (inp[7]) ? 4'b1011 : 4'b1010;
													assign node56419 = (inp[7]) ? 4'b1010 : node56420;
														assign node56420 = (inp[2]) ? 4'b1011 : 4'b1010;
											assign node56424 = (inp[7]) ? node56436 : node56425;
												assign node56425 = (inp[8]) ? node56431 : node56426;
													assign node56426 = (inp[14]) ? 4'b1000 : node56427;
														assign node56427 = (inp[2]) ? 4'b1000 : 4'b1001;
													assign node56431 = (inp[14]) ? 4'b1001 : node56432;
														assign node56432 = (inp[2]) ? 4'b1001 : 4'b1000;
												assign node56436 = (inp[8]) ? node56442 : node56437;
													assign node56437 = (inp[2]) ? 4'b1001 : node56438;
														assign node56438 = (inp[14]) ? 4'b1001 : 4'b1000;
													assign node56442 = (inp[2]) ? 4'b1000 : node56443;
														assign node56443 = (inp[14]) ? 4'b1000 : 4'b1001;
						assign node56447 = (inp[8]) ? node57249 : node56448;
							assign node56448 = (inp[7]) ? node56828 : node56449;
								assign node56449 = (inp[2]) ? node56635 : node56450;
									assign node56450 = (inp[14]) ? node56538 : node56451;
										assign node56451 = (inp[9]) ? node56501 : node56452;
											assign node56452 = (inp[4]) ? node56474 : node56453;
												assign node56453 = (inp[15]) ? node56465 : node56454;
													assign node56454 = (inp[0]) ? node56460 : node56455;
														assign node56455 = (inp[3]) ? node56457 : 4'b1011;
															assign node56457 = (inp[5]) ? 4'b1001 : 4'b1011;
														assign node56460 = (inp[3]) ? node56462 : 4'b1001;
															assign node56462 = (inp[5]) ? 4'b1011 : 4'b1001;
													assign node56465 = (inp[0]) ? node56471 : node56466;
														assign node56466 = (inp[3]) ? node56468 : 4'b1001;
															assign node56468 = (inp[5]) ? 4'b1011 : 4'b1001;
														assign node56471 = (inp[3]) ? 4'b1001 : 4'b1011;
												assign node56474 = (inp[5]) ? node56494 : node56475;
													assign node56475 = (inp[3]) ? node56485 : node56476;
														assign node56476 = (inp[12]) ? node56482 : node56477;
															assign node56477 = (inp[15]) ? 4'b1111 : node56478;
																assign node56478 = (inp[0]) ? 4'b1101 : 4'b1111;
															assign node56482 = (inp[15]) ? 4'b1101 : 4'b1111;
														assign node56485 = (inp[12]) ? node56489 : node56486;
															assign node56486 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node56489 = (inp[0]) ? node56491 : 4'b1101;
																assign node56491 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node56494 = (inp[3]) ? node56498 : node56495;
														assign node56495 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node56498 = (inp[0]) ? 4'b1101 : 4'b1111;
											assign node56501 = (inp[4]) ? node56519 : node56502;
												assign node56502 = (inp[3]) ? node56510 : node56503;
													assign node56503 = (inp[5]) ? node56505 : 4'b1111;
														assign node56505 = (inp[0]) ? node56507 : 4'b1111;
															assign node56507 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node56510 = (inp[12]) ? node56512 : 4'b1111;
														assign node56512 = (inp[15]) ? node56516 : node56513;
															assign node56513 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node56516 = (inp[0]) ? 4'b1101 : 4'b1111;
												assign node56519 = (inp[15]) ? node56529 : node56520;
													assign node56520 = (inp[0]) ? node56526 : node56521;
														assign node56521 = (inp[3]) ? 4'b1001 : node56522;
															assign node56522 = (inp[5]) ? 4'b1001 : 4'b1011;
														assign node56526 = (inp[5]) ? 4'b1011 : 4'b1001;
													assign node56529 = (inp[0]) ? node56531 : 4'b1011;
														assign node56531 = (inp[12]) ? 4'b1011 : node56532;
															assign node56532 = (inp[3]) ? 4'b1001 : node56533;
																assign node56533 = (inp[5]) ? 4'b1001 : 4'b1011;
										assign node56538 = (inp[0]) ? node56586 : node56539;
											assign node56539 = (inp[15]) ? node56561 : node56540;
												assign node56540 = (inp[3]) ? node56554 : node56541;
													assign node56541 = (inp[5]) ? node56549 : node56542;
														assign node56542 = (inp[9]) ? node56546 : node56543;
															assign node56543 = (inp[4]) ? 4'b1110 : 4'b1010;
															assign node56546 = (inp[4]) ? 4'b1010 : 4'b1110;
														assign node56549 = (inp[4]) ? 4'b1100 : node56550;
															assign node56550 = (inp[12]) ? 4'b1100 : 4'b1010;
													assign node56554 = (inp[9]) ? node56558 : node56555;
														assign node56555 = (inp[4]) ? 4'b1100 : 4'b1010;
														assign node56558 = (inp[4]) ? 4'b1000 : 4'b1100;
												assign node56561 = (inp[3]) ? node56575 : node56562;
													assign node56562 = (inp[5]) ? node56568 : node56563;
														assign node56563 = (inp[9]) ? node56565 : 4'b1100;
															assign node56565 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node56568 = (inp[12]) ? node56570 : 4'b1110;
															assign node56570 = (inp[4]) ? node56572 : 4'b1000;
																assign node56572 = (inp[9]) ? 4'b1010 : 4'b1110;
													assign node56575 = (inp[5]) ? node56581 : node56576;
														assign node56576 = (inp[4]) ? node56578 : 4'b1110;
															assign node56578 = (inp[9]) ? 4'b1010 : 4'b1110;
														assign node56581 = (inp[9]) ? 4'b1110 : node56582;
															assign node56582 = (inp[4]) ? 4'b1110 : 4'b1010;
											assign node56586 = (inp[15]) ? node56614 : node56587;
												assign node56587 = (inp[5]) ? node56603 : node56588;
													assign node56588 = (inp[3]) ? node56596 : node56589;
														assign node56589 = (inp[12]) ? node56591 : 4'b1000;
															assign node56591 = (inp[9]) ? 4'b1100 : node56592;
																assign node56592 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node56596 = (inp[9]) ? node56600 : node56597;
															assign node56597 = (inp[4]) ? 4'b1110 : 4'b1000;
															assign node56600 = (inp[4]) ? 4'b1010 : 4'b1110;
													assign node56603 = (inp[12]) ? node56605 : 4'b1110;
														assign node56605 = (inp[3]) ? 4'b1010 : node56606;
															assign node56606 = (inp[9]) ? node56610 : node56607;
																assign node56607 = (inp[4]) ? 4'b1110 : 4'b1000;
																assign node56610 = (inp[4]) ? 4'b1010 : 4'b1110;
												assign node56614 = (inp[5]) ? node56628 : node56615;
													assign node56615 = (inp[3]) ? node56621 : node56616;
														assign node56616 = (inp[9]) ? 4'b1110 : node56617;
															assign node56617 = (inp[4]) ? 4'b1110 : 4'b1010;
														assign node56621 = (inp[4]) ? node56625 : node56622;
															assign node56622 = (inp[9]) ? 4'b1100 : 4'b1010;
															assign node56625 = (inp[9]) ? 4'b1000 : 4'b1100;
													assign node56628 = (inp[4]) ? node56632 : node56629;
														assign node56629 = (inp[9]) ? 4'b1100 : 4'b1000;
														assign node56632 = (inp[9]) ? 4'b1000 : 4'b1100;
									assign node56635 = (inp[12]) ? node56739 : node56636;
										assign node56636 = (inp[0]) ? node56692 : node56637;
											assign node56637 = (inp[15]) ? node56663 : node56638;
												assign node56638 = (inp[3]) ? node56654 : node56639;
													assign node56639 = (inp[5]) ? node56647 : node56640;
														assign node56640 = (inp[9]) ? node56644 : node56641;
															assign node56641 = (inp[4]) ? 4'b1110 : 4'b1010;
															assign node56644 = (inp[4]) ? 4'b1010 : 4'b1110;
														assign node56647 = (inp[4]) ? node56651 : node56648;
															assign node56648 = (inp[9]) ? 4'b1100 : 4'b1010;
															assign node56651 = (inp[9]) ? 4'b1000 : 4'b1100;
													assign node56654 = (inp[9]) ? node56660 : node56655;
														assign node56655 = (inp[4]) ? 4'b1100 : node56656;
															assign node56656 = (inp[5]) ? 4'b1000 : 4'b1010;
														assign node56660 = (inp[4]) ? 4'b1000 : 4'b1100;
												assign node56663 = (inp[5]) ? node56677 : node56664;
													assign node56664 = (inp[3]) ? node56672 : node56665;
														assign node56665 = (inp[4]) ? node56669 : node56666;
															assign node56666 = (inp[9]) ? 4'b1100 : 4'b1000;
															assign node56669 = (inp[9]) ? 4'b1000 : 4'b1100;
														assign node56672 = (inp[9]) ? node56674 : 4'b1000;
															assign node56674 = (inp[4]) ? 4'b1010 : 4'b1110;
													assign node56677 = (inp[3]) ? node56685 : node56678;
														assign node56678 = (inp[9]) ? node56682 : node56679;
															assign node56679 = (inp[4]) ? 4'b1110 : 4'b1000;
															assign node56682 = (inp[4]) ? 4'b1010 : 4'b1110;
														assign node56685 = (inp[9]) ? node56689 : node56686;
															assign node56686 = (inp[4]) ? 4'b1110 : 4'b1010;
															assign node56689 = (inp[4]) ? 4'b1010 : 4'b1110;
											assign node56692 = (inp[3]) ? node56716 : node56693;
												assign node56693 = (inp[4]) ? node56703 : node56694;
													assign node56694 = (inp[9]) ? node56698 : node56695;
														assign node56695 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node56698 = (inp[5]) ? 4'b1100 : node56699;
															assign node56699 = (inp[15]) ? 4'b1110 : 4'b1100;
													assign node56703 = (inp[9]) ? node56709 : node56704;
														assign node56704 = (inp[14]) ? node56706 : 4'b1100;
															assign node56706 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node56709 = (inp[15]) ? node56713 : node56710;
															assign node56710 = (inp[5]) ? 4'b1010 : 4'b1000;
															assign node56713 = (inp[5]) ? 4'b1000 : 4'b1010;
												assign node56716 = (inp[15]) ? node56726 : node56717;
													assign node56717 = (inp[9]) ? node56723 : node56718;
														assign node56718 = (inp[4]) ? 4'b1110 : node56719;
															assign node56719 = (inp[5]) ? 4'b1010 : 4'b1000;
														assign node56723 = (inp[4]) ? 4'b1010 : 4'b1110;
													assign node56726 = (inp[5]) ? node56734 : node56727;
														assign node56727 = (inp[4]) ? node56731 : node56728;
															assign node56728 = (inp[9]) ? 4'b1100 : 4'b1010;
															assign node56731 = (inp[9]) ? 4'b1000 : 4'b1100;
														assign node56734 = (inp[4]) ? 4'b1100 : node56735;
															assign node56735 = (inp[14]) ? 4'b1100 : 4'b1000;
										assign node56739 = (inp[3]) ? node56791 : node56740;
											assign node56740 = (inp[9]) ? node56760 : node56741;
												assign node56741 = (inp[4]) ? node56747 : node56742;
													assign node56742 = (inp[15]) ? node56744 : 4'b1010;
														assign node56744 = (inp[0]) ? 4'b1010 : 4'b1000;
													assign node56747 = (inp[5]) ? node56755 : node56748;
														assign node56748 = (inp[15]) ? node56752 : node56749;
															assign node56749 = (inp[0]) ? 4'b1100 : 4'b1110;
															assign node56752 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node56755 = (inp[0]) ? 4'b1100 : node56756;
															assign node56756 = (inp[15]) ? 4'b1110 : 4'b1100;
												assign node56760 = (inp[4]) ? node56772 : node56761;
													assign node56761 = (inp[15]) ? 4'b1110 : node56762;
														assign node56762 = (inp[14]) ? 4'b1100 : node56763;
															assign node56763 = (inp[5]) ? node56767 : node56764;
																assign node56764 = (inp[0]) ? 4'b1100 : 4'b1110;
																assign node56767 = (inp[0]) ? 4'b1110 : 4'b1100;
													assign node56772 = (inp[14]) ? node56782 : node56773;
														assign node56773 = (inp[5]) ? 4'b1000 : node56774;
															assign node56774 = (inp[15]) ? node56778 : node56775;
																assign node56775 = (inp[0]) ? 4'b1000 : 4'b1010;
																assign node56778 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node56782 = (inp[5]) ? node56784 : 4'b1010;
															assign node56784 = (inp[15]) ? node56788 : node56785;
																assign node56785 = (inp[0]) ? 4'b1010 : 4'b1000;
																assign node56788 = (inp[0]) ? 4'b1000 : 4'b1010;
											assign node56791 = (inp[15]) ? node56815 : node56792;
												assign node56792 = (inp[0]) ? node56800 : node56793;
													assign node56793 = (inp[4]) ? node56797 : node56794;
														assign node56794 = (inp[9]) ? 4'b1100 : 4'b1010;
														assign node56797 = (inp[9]) ? 4'b1000 : 4'b1100;
													assign node56800 = (inp[5]) ? node56808 : node56801;
														assign node56801 = (inp[14]) ? node56803 : 4'b1110;
															assign node56803 = (inp[4]) ? 4'b1110 : node56804;
																assign node56804 = (inp[9]) ? 4'b1110 : 4'b1000;
														assign node56808 = (inp[14]) ? node56810 : 4'b1010;
															assign node56810 = (inp[4]) ? 4'b1010 : node56811;
																assign node56811 = (inp[9]) ? 4'b1110 : 4'b1010;
												assign node56815 = (inp[0]) ? node56823 : node56816;
													assign node56816 = (inp[4]) ? node56820 : node56817;
														assign node56817 = (inp[9]) ? 4'b1110 : 4'b1000;
														assign node56820 = (inp[9]) ? 4'b1010 : 4'b1110;
													assign node56823 = (inp[9]) ? 4'b1100 : node56824;
														assign node56824 = (inp[4]) ? 4'b1100 : 4'b1010;
								assign node56828 = (inp[14]) ? node57056 : node56829;
									assign node56829 = (inp[2]) ? node56943 : node56830;
										assign node56830 = (inp[0]) ? node56892 : node56831;
											assign node56831 = (inp[15]) ? node56863 : node56832;
												assign node56832 = (inp[5]) ? node56856 : node56833;
													assign node56833 = (inp[3]) ? node56849 : node56834;
														assign node56834 = (inp[12]) ? node56842 : node56835;
															assign node56835 = (inp[9]) ? node56839 : node56836;
																assign node56836 = (inp[4]) ? 4'b1110 : 4'b1010;
																assign node56839 = (inp[4]) ? 4'b1010 : 4'b1110;
															assign node56842 = (inp[9]) ? node56846 : node56843;
																assign node56843 = (inp[4]) ? 4'b1110 : 4'b1010;
																assign node56846 = (inp[4]) ? 4'b1010 : 4'b1110;
														assign node56849 = (inp[9]) ? node56853 : node56850;
															assign node56850 = (inp[4]) ? 4'b1100 : 4'b1010;
															assign node56853 = (inp[4]) ? 4'b1000 : 4'b1100;
													assign node56856 = (inp[3]) ? node56858 : 4'b1100;
														assign node56858 = (inp[4]) ? node56860 : 4'b1000;
															assign node56860 = (inp[9]) ? 4'b1000 : 4'b1100;
												assign node56863 = (inp[3]) ? node56879 : node56864;
													assign node56864 = (inp[5]) ? node56872 : node56865;
														assign node56865 = (inp[4]) ? node56869 : node56866;
															assign node56866 = (inp[9]) ? 4'b1100 : 4'b1000;
															assign node56869 = (inp[9]) ? 4'b1000 : 4'b1100;
														assign node56872 = (inp[9]) ? node56876 : node56873;
															assign node56873 = (inp[4]) ? 4'b1110 : 4'b1000;
															assign node56876 = (inp[4]) ? 4'b1010 : 4'b1110;
													assign node56879 = (inp[5]) ? node56887 : node56880;
														assign node56880 = (inp[4]) ? node56884 : node56881;
															assign node56881 = (inp[9]) ? 4'b1110 : 4'b1000;
															assign node56884 = (inp[9]) ? 4'b1010 : 4'b1110;
														assign node56887 = (inp[4]) ? 4'b1010 : node56888;
															assign node56888 = (inp[9]) ? 4'b1110 : 4'b1010;
											assign node56892 = (inp[15]) ? node56914 : node56893;
												assign node56893 = (inp[9]) ? node56905 : node56894;
													assign node56894 = (inp[4]) ? node56900 : node56895;
														assign node56895 = (inp[5]) ? node56897 : 4'b1000;
															assign node56897 = (inp[3]) ? 4'b1010 : 4'b1000;
														assign node56900 = (inp[3]) ? 4'b1110 : node56901;
															assign node56901 = (inp[5]) ? 4'b1110 : 4'b1100;
													assign node56905 = (inp[4]) ? node56907 : 4'b1110;
														assign node56907 = (inp[12]) ? 4'b1010 : node56908;
															assign node56908 = (inp[5]) ? 4'b1010 : node56909;
																assign node56909 = (inp[3]) ? 4'b1010 : 4'b1000;
												assign node56914 = (inp[3]) ? node56930 : node56915;
													assign node56915 = (inp[5]) ? node56923 : node56916;
														assign node56916 = (inp[9]) ? node56920 : node56917;
															assign node56917 = (inp[4]) ? 4'b1110 : 4'b1010;
															assign node56920 = (inp[4]) ? 4'b1010 : 4'b1110;
														assign node56923 = (inp[12]) ? node56925 : 4'b1100;
															assign node56925 = (inp[4]) ? node56927 : 4'b1010;
																assign node56927 = (inp[9]) ? 4'b1000 : 4'b1100;
													assign node56930 = (inp[5]) ? node56938 : node56931;
														assign node56931 = (inp[4]) ? node56935 : node56932;
															assign node56932 = (inp[9]) ? 4'b1100 : 4'b1010;
															assign node56935 = (inp[9]) ? 4'b1000 : 4'b1100;
														assign node56938 = (inp[4]) ? 4'b1100 : node56939;
															assign node56939 = (inp[9]) ? 4'b1100 : 4'b1000;
										assign node56943 = (inp[5]) ? node57001 : node56944;
											assign node56944 = (inp[9]) ? node56970 : node56945;
												assign node56945 = (inp[4]) ? node56953 : node56946;
													assign node56946 = (inp[15]) ? node56950 : node56947;
														assign node56947 = (inp[0]) ? 4'b0001 : 4'b0011;
														assign node56950 = (inp[0]) ? 4'b0011 : 4'b0001;
													assign node56953 = (inp[0]) ? node56963 : node56954;
														assign node56954 = (inp[12]) ? node56956 : 4'b0101;
															assign node56956 = (inp[15]) ? node56960 : node56957;
																assign node56957 = (inp[3]) ? 4'b0101 : 4'b0111;
																assign node56960 = (inp[3]) ? 4'b0111 : 4'b0101;
														assign node56963 = (inp[15]) ? node56967 : node56964;
															assign node56964 = (inp[3]) ? 4'b0111 : 4'b0101;
															assign node56967 = (inp[3]) ? 4'b0101 : 4'b0111;
												assign node56970 = (inp[4]) ? node56980 : node56971;
													assign node56971 = (inp[12]) ? 4'b0111 : node56972;
														assign node56972 = (inp[3]) ? 4'b0111 : node56973;
															assign node56973 = (inp[15]) ? node56975 : 4'b0101;
																assign node56975 = (inp[0]) ? 4'b0111 : 4'b0101;
													assign node56980 = (inp[12]) ? node56988 : node56981;
														assign node56981 = (inp[15]) ? node56983 : 4'b0011;
															assign node56983 = (inp[3]) ? 4'b0011 : node56984;
																assign node56984 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node56988 = (inp[0]) ? node56996 : node56989;
															assign node56989 = (inp[3]) ? node56993 : node56990;
																assign node56990 = (inp[15]) ? 4'b0001 : 4'b0011;
																assign node56993 = (inp[15]) ? 4'b0011 : 4'b0001;
															assign node56996 = (inp[15]) ? node56998 : 4'b0011;
																assign node56998 = (inp[3]) ? 4'b0001 : 4'b0011;
											assign node57001 = (inp[0]) ? node57023 : node57002;
												assign node57002 = (inp[15]) ? node57016 : node57003;
													assign node57003 = (inp[3]) ? node57011 : node57004;
														assign node57004 = (inp[4]) ? node57008 : node57005;
															assign node57005 = (inp[9]) ? 4'b0101 : 4'b0011;
															assign node57008 = (inp[9]) ? 4'b0001 : 4'b0101;
														assign node57011 = (inp[4]) ? node57013 : 4'b0001;
															assign node57013 = (inp[9]) ? 4'b0001 : 4'b0101;
													assign node57016 = (inp[9]) ? node57020 : node57017;
														assign node57017 = (inp[4]) ? 4'b0111 : 4'b0001;
														assign node57020 = (inp[4]) ? 4'b0011 : 4'b0111;
												assign node57023 = (inp[15]) ? node57033 : node57024;
													assign node57024 = (inp[3]) ? node57030 : node57025;
														assign node57025 = (inp[4]) ? node57027 : 4'b0001;
															assign node57027 = (inp[9]) ? 4'b0011 : 4'b0111;
														assign node57030 = (inp[9]) ? 4'b0111 : 4'b0011;
													assign node57033 = (inp[3]) ? node57041 : node57034;
														assign node57034 = (inp[4]) ? node57038 : node57035;
															assign node57035 = (inp[9]) ? 4'b0101 : 4'b0011;
															assign node57038 = (inp[9]) ? 4'b0001 : 4'b0101;
														assign node57041 = (inp[12]) ? node57049 : node57042;
															assign node57042 = (inp[4]) ? node57046 : node57043;
																assign node57043 = (inp[9]) ? 4'b0101 : 4'b0001;
																assign node57046 = (inp[9]) ? 4'b0001 : 4'b0101;
															assign node57049 = (inp[9]) ? node57053 : node57050;
																assign node57050 = (inp[4]) ? 4'b0101 : 4'b0001;
																assign node57053 = (inp[4]) ? 4'b0001 : 4'b0101;
									assign node57056 = (inp[12]) ? node57164 : node57057;
										assign node57057 = (inp[2]) ? node57115 : node57058;
											assign node57058 = (inp[3]) ? node57086 : node57059;
												assign node57059 = (inp[0]) ? node57073 : node57060;
													assign node57060 = (inp[4]) ? node57066 : node57061;
														assign node57061 = (inp[9]) ? 4'b0101 : node57062;
															assign node57062 = (inp[15]) ? 4'b0001 : 4'b0011;
														assign node57066 = (inp[9]) ? 4'b0011 : node57067;
															assign node57067 = (inp[5]) ? node57069 : 4'b0111;
																assign node57069 = (inp[15]) ? 4'b0111 : 4'b0101;
													assign node57073 = (inp[5]) ? node57077 : node57074;
														assign node57074 = (inp[15]) ? 4'b0111 : 4'b0101;
														assign node57077 = (inp[15]) ? node57079 : 4'b0111;
															assign node57079 = (inp[9]) ? node57083 : node57080;
																assign node57080 = (inp[4]) ? 4'b0101 : 4'b0011;
																assign node57083 = (inp[4]) ? 4'b0001 : 4'b0101;
												assign node57086 = (inp[9]) ? node57104 : node57087;
													assign node57087 = (inp[4]) ? node57097 : node57088;
														assign node57088 = (inp[0]) ? 4'b0001 : node57089;
															assign node57089 = (inp[5]) ? node57093 : node57090;
																assign node57090 = (inp[15]) ? 4'b0001 : 4'b0011;
																assign node57093 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node57097 = (inp[0]) ? node57101 : node57098;
															assign node57098 = (inp[15]) ? 4'b0111 : 4'b0101;
															assign node57101 = (inp[15]) ? 4'b0101 : 4'b0111;
													assign node57104 = (inp[4]) ? node57112 : node57105;
														assign node57105 = (inp[15]) ? node57109 : node57106;
															assign node57106 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node57109 = (inp[0]) ? 4'b0101 : 4'b0111;
														assign node57112 = (inp[15]) ? 4'b0001 : 4'b0011;
											assign node57115 = (inp[9]) ? node57151 : node57116;
												assign node57116 = (inp[4]) ? node57138 : node57117;
													assign node57117 = (inp[5]) ? node57125 : node57118;
														assign node57118 = (inp[15]) ? node57122 : node57119;
															assign node57119 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node57122 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node57125 = (inp[0]) ? node57133 : node57126;
															assign node57126 = (inp[3]) ? node57130 : node57127;
																assign node57127 = (inp[15]) ? 4'b0001 : 4'b0011;
																assign node57130 = (inp[15]) ? 4'b0011 : 4'b0001;
															assign node57133 = (inp[15]) ? 4'b0011 : node57134;
																assign node57134 = (inp[3]) ? 4'b0011 : 4'b0001;
													assign node57138 = (inp[15]) ? 4'b0111 : node57139;
														assign node57139 = (inp[0]) ? node57145 : node57140;
															assign node57140 = (inp[3]) ? 4'b0101 : node57141;
																assign node57141 = (inp[5]) ? 4'b0101 : 4'b0111;
															assign node57145 = (inp[3]) ? 4'b0111 : node57146;
																assign node57146 = (inp[5]) ? 4'b0111 : 4'b0101;
												assign node57151 = (inp[4]) ? node57157 : node57152;
													assign node57152 = (inp[0]) ? 4'b0111 : node57153;
														assign node57153 = (inp[5]) ? 4'b0111 : 4'b0101;
													assign node57157 = (inp[15]) ? 4'b0011 : node57158;
														assign node57158 = (inp[5]) ? 4'b0011 : node57159;
															assign node57159 = (inp[3]) ? 4'b0011 : 4'b0001;
										assign node57164 = (inp[15]) ? node57210 : node57165;
											assign node57165 = (inp[0]) ? node57183 : node57166;
												assign node57166 = (inp[5]) ? node57174 : node57167;
													assign node57167 = (inp[3]) ? 4'b0101 : node57168;
														assign node57168 = (inp[9]) ? node57170 : 4'b0111;
															assign node57170 = (inp[4]) ? 4'b0011 : 4'b0111;
													assign node57174 = (inp[4]) ? node57180 : node57175;
														assign node57175 = (inp[9]) ? 4'b0101 : node57176;
															assign node57176 = (inp[3]) ? 4'b0001 : 4'b0011;
														assign node57180 = (inp[9]) ? 4'b0001 : 4'b0101;
												assign node57183 = (inp[5]) ? node57201 : node57184;
													assign node57184 = (inp[3]) ? node57194 : node57185;
														assign node57185 = (inp[2]) ? 4'b0101 : node57186;
															assign node57186 = (inp[4]) ? node57190 : node57187;
																assign node57187 = (inp[9]) ? 4'b0101 : 4'b0001;
																assign node57190 = (inp[9]) ? 4'b0001 : 4'b0101;
														assign node57194 = (inp[9]) ? node57198 : node57195;
															assign node57195 = (inp[4]) ? 4'b0111 : 4'b0001;
															assign node57198 = (inp[4]) ? 4'b0011 : 4'b0111;
													assign node57201 = (inp[4]) ? node57207 : node57202;
														assign node57202 = (inp[9]) ? 4'b0111 : node57203;
															assign node57203 = (inp[2]) ? 4'b0001 : 4'b0011;
														assign node57207 = (inp[9]) ? 4'b0011 : 4'b0111;
											assign node57210 = (inp[0]) ? node57236 : node57211;
												assign node57211 = (inp[3]) ? node57227 : node57212;
													assign node57212 = (inp[5]) ? node57220 : node57213;
														assign node57213 = (inp[2]) ? node57215 : 4'b0101;
															assign node57215 = (inp[9]) ? node57217 : 4'b0101;
																assign node57217 = (inp[4]) ? 4'b0001 : 4'b0101;
														assign node57220 = (inp[4]) ? node57224 : node57221;
															assign node57221 = (inp[9]) ? 4'b0111 : 4'b0001;
															assign node57224 = (inp[2]) ? 4'b0111 : 4'b0011;
													assign node57227 = (inp[9]) ? node57233 : node57228;
														assign node57228 = (inp[4]) ? 4'b0111 : node57229;
															assign node57229 = (inp[5]) ? 4'b0011 : 4'b0001;
														assign node57233 = (inp[4]) ? 4'b0011 : 4'b0111;
												assign node57236 = (inp[4]) ? node57246 : node57237;
													assign node57237 = (inp[9]) ? node57243 : node57238;
														assign node57238 = (inp[5]) ? node57240 : 4'b0011;
															assign node57240 = (inp[3]) ? 4'b0001 : 4'b0011;
														assign node57243 = (inp[3]) ? 4'b0101 : 4'b0111;
													assign node57246 = (inp[9]) ? 4'b0001 : 4'b0101;
							assign node57249 = (inp[7]) ? node57627 : node57250;
								assign node57250 = (inp[2]) ? node57468 : node57251;
									assign node57251 = (inp[14]) ? node57365 : node57252;
										assign node57252 = (inp[3]) ? node57312 : node57253;
											assign node57253 = (inp[4]) ? node57279 : node57254;
												assign node57254 = (inp[9]) ? node57264 : node57255;
													assign node57255 = (inp[5]) ? node57257 : 4'b1000;
														assign node57257 = (inp[0]) ? node57261 : node57258;
															assign node57258 = (inp[15]) ? 4'b1000 : 4'b1010;
															assign node57261 = (inp[15]) ? 4'b1010 : 4'b1000;
													assign node57264 = (inp[15]) ? node57272 : node57265;
														assign node57265 = (inp[12]) ? 4'b1110 : node57266;
															assign node57266 = (inp[5]) ? node57268 : 4'b1100;
																assign node57268 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node57272 = (inp[5]) ? node57276 : node57273;
															assign node57273 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node57276 = (inp[0]) ? 4'b1100 : 4'b1110;
												assign node57279 = (inp[9]) ? node57301 : node57280;
													assign node57280 = (inp[0]) ? node57288 : node57281;
														assign node57281 = (inp[5]) ? node57285 : node57282;
															assign node57282 = (inp[15]) ? 4'b1100 : 4'b1110;
															assign node57285 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node57288 = (inp[12]) ? node57294 : node57289;
															assign node57289 = (inp[5]) ? node57291 : 4'b1100;
																assign node57291 = (inp[15]) ? 4'b1100 : 4'b1110;
															assign node57294 = (inp[5]) ? node57298 : node57295;
																assign node57295 = (inp[15]) ? 4'b1110 : 4'b1100;
																assign node57298 = (inp[15]) ? 4'b1100 : 4'b1110;
													assign node57301 = (inp[5]) ? node57307 : node57302;
														assign node57302 = (inp[15]) ? 4'b1000 : node57303;
															assign node57303 = (inp[0]) ? 4'b1000 : 4'b1010;
														assign node57307 = (inp[12]) ? 4'b1010 : node57308;
															assign node57308 = (inp[15]) ? 4'b1010 : 4'b1000;
											assign node57312 = (inp[0]) ? node57334 : node57313;
												assign node57313 = (inp[15]) ? node57327 : node57314;
													assign node57314 = (inp[5]) ? node57320 : node57315;
														assign node57315 = (inp[4]) ? node57317 : 4'b1010;
															assign node57317 = (inp[9]) ? 4'b1000 : 4'b1100;
														assign node57320 = (inp[9]) ? node57324 : node57321;
															assign node57321 = (inp[4]) ? 4'b1100 : 4'b1000;
															assign node57324 = (inp[4]) ? 4'b1000 : 4'b1100;
													assign node57327 = (inp[4]) ? node57331 : node57328;
														assign node57328 = (inp[9]) ? 4'b1110 : 4'b1000;
														assign node57331 = (inp[9]) ? 4'b1010 : 4'b1110;
												assign node57334 = (inp[15]) ? node57352 : node57335;
													assign node57335 = (inp[5]) ? node57343 : node57336;
														assign node57336 = (inp[9]) ? node57340 : node57337;
															assign node57337 = (inp[4]) ? 4'b1110 : 4'b1000;
															assign node57340 = (inp[4]) ? 4'b1010 : 4'b1110;
														assign node57343 = (inp[12]) ? node57345 : 4'b1010;
															assign node57345 = (inp[4]) ? node57349 : node57346;
																assign node57346 = (inp[9]) ? 4'b1110 : 4'b1010;
																assign node57349 = (inp[9]) ? 4'b1010 : 4'b1110;
													assign node57352 = (inp[5]) ? 4'b1000 : node57353;
														assign node57353 = (inp[12]) ? node57359 : node57354;
															assign node57354 = (inp[4]) ? node57356 : 4'b1010;
																assign node57356 = (inp[9]) ? 4'b1000 : 4'b1100;
															assign node57359 = (inp[4]) ? node57361 : 4'b1100;
																assign node57361 = (inp[9]) ? 4'b1000 : 4'b1100;
										assign node57365 = (inp[3]) ? node57419 : node57366;
											assign node57366 = (inp[15]) ? node57392 : node57367;
												assign node57367 = (inp[0]) ? node57379 : node57368;
													assign node57368 = (inp[5]) ? node57374 : node57369;
														assign node57369 = (inp[9]) ? node57371 : 4'b0111;
															assign node57371 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node57374 = (inp[9]) ? 4'b0101 : node57375;
															assign node57375 = (inp[4]) ? 4'b0101 : 4'b0011;
													assign node57379 = (inp[5]) ? node57387 : node57380;
														assign node57380 = (inp[4]) ? node57384 : node57381;
															assign node57381 = (inp[9]) ? 4'b0101 : 4'b0001;
															assign node57384 = (inp[9]) ? 4'b0001 : 4'b0101;
														assign node57387 = (inp[4]) ? node57389 : 4'b0111;
															assign node57389 = (inp[9]) ? 4'b0011 : 4'b0111;
												assign node57392 = (inp[5]) ? node57404 : node57393;
													assign node57393 = (inp[0]) ? node57399 : node57394;
														assign node57394 = (inp[4]) ? node57396 : 4'b0101;
															assign node57396 = (inp[12]) ? 4'b0001 : 4'b0101;
														assign node57399 = (inp[4]) ? 4'b0111 : node57400;
															assign node57400 = (inp[9]) ? 4'b0111 : 4'b0011;
													assign node57404 = (inp[0]) ? node57412 : node57405;
														assign node57405 = (inp[9]) ? node57409 : node57406;
															assign node57406 = (inp[4]) ? 4'b0111 : 4'b0001;
															assign node57409 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node57412 = (inp[9]) ? node57416 : node57413;
															assign node57413 = (inp[4]) ? 4'b0101 : 4'b0011;
															assign node57416 = (inp[4]) ? 4'b0001 : 4'b0101;
											assign node57419 = (inp[0]) ? node57441 : node57420;
												assign node57420 = (inp[15]) ? node57432 : node57421;
													assign node57421 = (inp[12]) ? node57423 : 4'b0101;
														assign node57423 = (inp[5]) ? node57427 : node57424;
															assign node57424 = (inp[4]) ? 4'b0001 : 4'b0011;
															assign node57427 = (inp[4]) ? node57429 : 4'b0101;
																assign node57429 = (inp[9]) ? 4'b0001 : 4'b0101;
													assign node57432 = (inp[4]) ? node57438 : node57433;
														assign node57433 = (inp[9]) ? 4'b0111 : node57434;
															assign node57434 = (inp[5]) ? 4'b0011 : 4'b0001;
														assign node57438 = (inp[9]) ? 4'b0011 : 4'b0111;
												assign node57441 = (inp[15]) ? node57461 : node57442;
													assign node57442 = (inp[5]) ? node57450 : node57443;
														assign node57443 = (inp[9]) ? node57447 : node57444;
															assign node57444 = (inp[4]) ? 4'b0111 : 4'b0001;
															assign node57447 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node57450 = (inp[12]) ? node57456 : node57451;
															assign node57451 = (inp[4]) ? node57453 : 4'b0011;
																assign node57453 = (inp[9]) ? 4'b0011 : 4'b0111;
															assign node57456 = (inp[9]) ? node57458 : 4'b0011;
																assign node57458 = (inp[4]) ? 4'b0011 : 4'b0111;
													assign node57461 = (inp[9]) ? node57465 : node57462;
														assign node57462 = (inp[4]) ? 4'b0101 : 4'b0001;
														assign node57465 = (inp[4]) ? 4'b0001 : 4'b0101;
									assign node57468 = (inp[0]) ? node57554 : node57469;
										assign node57469 = (inp[15]) ? node57529 : node57470;
											assign node57470 = (inp[3]) ? node57500 : node57471;
												assign node57471 = (inp[5]) ? node57493 : node57472;
													assign node57472 = (inp[14]) ? node57488 : node57473;
														assign node57473 = (inp[12]) ? node57481 : node57474;
															assign node57474 = (inp[4]) ? node57478 : node57475;
																assign node57475 = (inp[9]) ? 4'b0111 : 4'b0011;
																assign node57478 = (inp[9]) ? 4'b0011 : 4'b0111;
															assign node57481 = (inp[9]) ? node57485 : node57482;
																assign node57482 = (inp[4]) ? 4'b0111 : 4'b0011;
																assign node57485 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node57488 = (inp[4]) ? 4'b0111 : node57489;
															assign node57489 = (inp[9]) ? 4'b0111 : 4'b0011;
													assign node57493 = (inp[4]) ? node57497 : node57494;
														assign node57494 = (inp[9]) ? 4'b0101 : 4'b0011;
														assign node57497 = (inp[9]) ? 4'b0001 : 4'b0101;
												assign node57500 = (inp[5]) ? node57510 : node57501;
													assign node57501 = (inp[12]) ? node57503 : 4'b0101;
														assign node57503 = (inp[4]) ? node57507 : node57504;
															assign node57504 = (inp[9]) ? 4'b0101 : 4'b0011;
															assign node57507 = (inp[9]) ? 4'b0001 : 4'b0101;
													assign node57510 = (inp[12]) ? node57516 : node57511;
														assign node57511 = (inp[4]) ? 4'b0001 : node57512;
															assign node57512 = (inp[9]) ? 4'b0101 : 4'b0001;
														assign node57516 = (inp[14]) ? node57522 : node57517;
															assign node57517 = (inp[4]) ? 4'b0101 : node57518;
																assign node57518 = (inp[9]) ? 4'b0101 : 4'b0001;
															assign node57522 = (inp[4]) ? node57526 : node57523;
																assign node57523 = (inp[9]) ? 4'b0101 : 4'b0001;
																assign node57526 = (inp[9]) ? 4'b0001 : 4'b0101;
											assign node57529 = (inp[3]) ? node57545 : node57530;
												assign node57530 = (inp[5]) ? node57538 : node57531;
													assign node57531 = (inp[4]) ? node57535 : node57532;
														assign node57532 = (inp[9]) ? 4'b0101 : 4'b0001;
														assign node57535 = (inp[9]) ? 4'b0001 : 4'b0101;
													assign node57538 = (inp[9]) ? node57542 : node57539;
														assign node57539 = (inp[4]) ? 4'b0111 : 4'b0001;
														assign node57542 = (inp[4]) ? 4'b0011 : 4'b0111;
												assign node57545 = (inp[9]) ? node57551 : node57546;
													assign node57546 = (inp[4]) ? 4'b0111 : node57547;
														assign node57547 = (inp[5]) ? 4'b0011 : 4'b0001;
													assign node57551 = (inp[4]) ? 4'b0011 : 4'b0111;
										assign node57554 = (inp[15]) ? node57594 : node57555;
											assign node57555 = (inp[3]) ? node57571 : node57556;
												assign node57556 = (inp[5]) ? node57564 : node57557;
													assign node57557 = (inp[4]) ? node57561 : node57558;
														assign node57558 = (inp[9]) ? 4'b0101 : 4'b0001;
														assign node57561 = (inp[9]) ? 4'b0001 : 4'b0101;
													assign node57564 = (inp[4]) ? node57568 : node57565;
														assign node57565 = (inp[9]) ? 4'b0111 : 4'b0001;
														assign node57568 = (inp[9]) ? 4'b0011 : 4'b0111;
												assign node57571 = (inp[12]) ? node57579 : node57572;
													assign node57572 = (inp[9]) ? node57576 : node57573;
														assign node57573 = (inp[5]) ? 4'b0011 : 4'b0111;
														assign node57576 = (inp[5]) ? 4'b0111 : 4'b0011;
													assign node57579 = (inp[5]) ? node57587 : node57580;
														assign node57580 = (inp[4]) ? node57584 : node57581;
															assign node57581 = (inp[9]) ? 4'b0111 : 4'b0001;
															assign node57584 = (inp[9]) ? 4'b0011 : 4'b0111;
														assign node57587 = (inp[9]) ? node57591 : node57588;
															assign node57588 = (inp[4]) ? 4'b0111 : 4'b0011;
															assign node57591 = (inp[4]) ? 4'b0011 : 4'b0111;
											assign node57594 = (inp[5]) ? node57612 : node57595;
												assign node57595 = (inp[3]) ? node57605 : node57596;
													assign node57596 = (inp[14]) ? 4'b0011 : node57597;
														assign node57597 = (inp[4]) ? node57601 : node57598;
															assign node57598 = (inp[9]) ? 4'b0111 : 4'b0011;
															assign node57601 = (inp[9]) ? 4'b0011 : 4'b0111;
													assign node57605 = (inp[9]) ? node57609 : node57606;
														assign node57606 = (inp[4]) ? 4'b0101 : 4'b0011;
														assign node57609 = (inp[4]) ? 4'b0001 : 4'b0101;
												assign node57612 = (inp[3]) ? node57620 : node57613;
													assign node57613 = (inp[9]) ? node57617 : node57614;
														assign node57614 = (inp[4]) ? 4'b0101 : 4'b0011;
														assign node57617 = (inp[4]) ? 4'b0001 : 4'b0101;
													assign node57620 = (inp[4]) ? node57624 : node57621;
														assign node57621 = (inp[9]) ? 4'b0101 : 4'b0001;
														assign node57624 = (inp[9]) ? 4'b0001 : 4'b0101;
								assign node57627 = (inp[2]) ? node57843 : node57628;
									assign node57628 = (inp[14]) ? node57720 : node57629;
										assign node57629 = (inp[15]) ? node57685 : node57630;
											assign node57630 = (inp[0]) ? node57654 : node57631;
												assign node57631 = (inp[5]) ? node57645 : node57632;
													assign node57632 = (inp[3]) ? node57640 : node57633;
														assign node57633 = (inp[12]) ? node57635 : 4'b0011;
															assign node57635 = (inp[9]) ? node57637 : 4'b0111;
																assign node57637 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node57640 = (inp[4]) ? node57642 : 4'b0011;
															assign node57642 = (inp[9]) ? 4'b0001 : 4'b0101;
													assign node57645 = (inp[4]) ? node57651 : node57646;
														assign node57646 = (inp[9]) ? 4'b0101 : node57647;
															assign node57647 = (inp[3]) ? 4'b0001 : 4'b0011;
														assign node57651 = (inp[9]) ? 4'b0001 : 4'b0101;
												assign node57654 = (inp[5]) ? node57676 : node57655;
													assign node57655 = (inp[3]) ? node57669 : node57656;
														assign node57656 = (inp[12]) ? node57664 : node57657;
															assign node57657 = (inp[9]) ? node57661 : node57658;
																assign node57658 = (inp[4]) ? 4'b0101 : 4'b0001;
																assign node57661 = (inp[4]) ? 4'b0001 : 4'b0101;
															assign node57664 = (inp[4]) ? node57666 : 4'b0101;
																assign node57666 = (inp[9]) ? 4'b0001 : 4'b0101;
														assign node57669 = (inp[9]) ? node57673 : node57670;
															assign node57670 = (inp[4]) ? 4'b0111 : 4'b0001;
															assign node57673 = (inp[4]) ? 4'b0011 : 4'b0111;
													assign node57676 = (inp[4]) ? node57682 : node57677;
														assign node57677 = (inp[9]) ? 4'b0111 : node57678;
															assign node57678 = (inp[3]) ? 4'b0011 : 4'b0001;
														assign node57682 = (inp[9]) ? 4'b0011 : 4'b0111;
											assign node57685 = (inp[0]) ? node57703 : node57686;
												assign node57686 = (inp[3]) ? node57698 : node57687;
													assign node57687 = (inp[5]) ? node57693 : node57688;
														assign node57688 = (inp[4]) ? node57690 : 4'b0001;
															assign node57690 = (inp[9]) ? 4'b0001 : 4'b0101;
														assign node57693 = (inp[4]) ? 4'b0111 : node57694;
															assign node57694 = (inp[9]) ? 4'b0111 : 4'b0001;
													assign node57698 = (inp[4]) ? node57700 : 4'b0111;
														assign node57700 = (inp[9]) ? 4'b0011 : 4'b0111;
												assign node57703 = (inp[5]) ? node57713 : node57704;
													assign node57704 = (inp[3]) ? node57708 : node57705;
														assign node57705 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node57708 = (inp[4]) ? node57710 : 4'b0101;
															assign node57710 = (inp[9]) ? 4'b0001 : 4'b0101;
													assign node57713 = (inp[9]) ? node57717 : node57714;
														assign node57714 = (inp[4]) ? 4'b0101 : 4'b0001;
														assign node57717 = (inp[4]) ? 4'b0001 : 4'b0101;
										assign node57720 = (inp[5]) ? node57794 : node57721;
											assign node57721 = (inp[12]) ? node57761 : node57722;
												assign node57722 = (inp[0]) ? node57742 : node57723;
													assign node57723 = (inp[4]) ? node57729 : node57724;
														assign node57724 = (inp[15]) ? 4'b0000 : node57725;
															assign node57725 = (inp[9]) ? 4'b0110 : 4'b0010;
														assign node57729 = (inp[9]) ? node57735 : node57730;
															assign node57730 = (inp[15]) ? node57732 : 4'b0100;
																assign node57732 = (inp[3]) ? 4'b0110 : 4'b0100;
															assign node57735 = (inp[15]) ? node57739 : node57736;
																assign node57736 = (inp[3]) ? 4'b0000 : 4'b0010;
																assign node57739 = (inp[3]) ? 4'b0010 : 4'b0000;
													assign node57742 = (inp[15]) ? node57754 : node57743;
														assign node57743 = (inp[3]) ? node57751 : node57744;
															assign node57744 = (inp[9]) ? node57748 : node57745;
																assign node57745 = (inp[4]) ? 4'b0100 : 4'b0000;
																assign node57748 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node57751 = (inp[9]) ? 4'b0110 : 4'b0000;
														assign node57754 = (inp[9]) ? node57758 : node57755;
															assign node57755 = (inp[4]) ? 4'b0110 : 4'b0010;
															assign node57758 = (inp[4]) ? 4'b0010 : 4'b0100;
												assign node57761 = (inp[9]) ? node57777 : node57762;
													assign node57762 = (inp[4]) ? node57772 : node57763;
														assign node57763 = (inp[3]) ? 4'b0000 : node57764;
															assign node57764 = (inp[0]) ? node57768 : node57765;
																assign node57765 = (inp[15]) ? 4'b0000 : 4'b0010;
																assign node57768 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node57772 = (inp[15]) ? node57774 : 4'b0110;
															assign node57774 = (inp[0]) ? 4'b0110 : 4'b0100;
													assign node57777 = (inp[4]) ? node57787 : node57778;
														assign node57778 = (inp[15]) ? 4'b0100 : node57779;
															assign node57779 = (inp[3]) ? node57783 : node57780;
																assign node57780 = (inp[0]) ? 4'b0100 : 4'b0110;
																assign node57783 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node57787 = (inp[0]) ? 4'b0000 : node57788;
															assign node57788 = (inp[15]) ? 4'b0000 : node57789;
																assign node57789 = (inp[3]) ? 4'b0000 : 4'b0010;
											assign node57794 = (inp[0]) ? node57818 : node57795;
												assign node57795 = (inp[15]) ? node57809 : node57796;
													assign node57796 = (inp[3]) ? node57802 : node57797;
														assign node57797 = (inp[9]) ? node57799 : 4'b0010;
															assign node57799 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node57802 = (inp[4]) ? node57806 : node57803;
															assign node57803 = (inp[9]) ? 4'b0100 : 4'b0000;
															assign node57806 = (inp[9]) ? 4'b0000 : 4'b0100;
													assign node57809 = (inp[4]) ? node57815 : node57810;
														assign node57810 = (inp[9]) ? 4'b0110 : node57811;
															assign node57811 = (inp[3]) ? 4'b0010 : 4'b0000;
														assign node57815 = (inp[9]) ? 4'b0010 : 4'b0110;
												assign node57818 = (inp[15]) ? node57834 : node57819;
													assign node57819 = (inp[12]) ? node57821 : 4'b0110;
														assign node57821 = (inp[3]) ? node57827 : node57822;
															assign node57822 = (inp[4]) ? 4'b0110 : node57823;
																assign node57823 = (inp[9]) ? 4'b0110 : 4'b0000;
															assign node57827 = (inp[9]) ? node57831 : node57828;
																assign node57828 = (inp[4]) ? 4'b0110 : 4'b0010;
																assign node57831 = (inp[4]) ? 4'b0010 : 4'b0110;
													assign node57834 = (inp[4]) ? node57840 : node57835;
														assign node57835 = (inp[9]) ? 4'b0100 : node57836;
															assign node57836 = (inp[3]) ? 4'b0000 : 4'b0010;
														assign node57840 = (inp[9]) ? 4'b0000 : 4'b0100;
									assign node57843 = (inp[4]) ? node57959 : node57844;
										assign node57844 = (inp[9]) ? node57908 : node57845;
											assign node57845 = (inp[14]) ? node57865 : node57846;
												assign node57846 = (inp[0]) ? node57856 : node57847;
													assign node57847 = (inp[15]) ? node57853 : node57848;
														assign node57848 = (inp[5]) ? node57850 : 4'b0010;
															assign node57850 = (inp[3]) ? 4'b0000 : 4'b0010;
														assign node57853 = (inp[5]) ? 4'b0010 : 4'b0000;
													assign node57856 = (inp[15]) ? node57860 : node57857;
														assign node57857 = (inp[3]) ? 4'b0010 : 4'b0000;
														assign node57860 = (inp[3]) ? node57862 : 4'b0010;
															assign node57862 = (inp[5]) ? 4'b0000 : 4'b0010;
												assign node57865 = (inp[12]) ? node57889 : node57866;
													assign node57866 = (inp[0]) ? node57878 : node57867;
														assign node57867 = (inp[15]) ? node57873 : node57868;
															assign node57868 = (inp[5]) ? node57870 : 4'b0010;
																assign node57870 = (inp[3]) ? 4'b0000 : 4'b0010;
															assign node57873 = (inp[5]) ? node57875 : 4'b0000;
																assign node57875 = (inp[3]) ? 4'b0010 : 4'b0000;
														assign node57878 = (inp[15]) ? node57884 : node57879;
															assign node57879 = (inp[3]) ? node57881 : 4'b0000;
																assign node57881 = (inp[5]) ? 4'b0010 : 4'b0000;
															assign node57884 = (inp[5]) ? node57886 : 4'b0010;
																assign node57886 = (inp[3]) ? 4'b0000 : 4'b0010;
													assign node57889 = (inp[5]) ? node57895 : node57890;
														assign node57890 = (inp[0]) ? node57892 : 4'b0010;
															assign node57892 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node57895 = (inp[0]) ? node57903 : node57896;
															assign node57896 = (inp[15]) ? node57900 : node57897;
																assign node57897 = (inp[3]) ? 4'b0000 : 4'b0010;
																assign node57900 = (inp[3]) ? 4'b0010 : 4'b0000;
															assign node57903 = (inp[15]) ? node57905 : 4'b0000;
																assign node57905 = (inp[3]) ? 4'b0000 : 4'b0010;
											assign node57908 = (inp[3]) ? node57944 : node57909;
												assign node57909 = (inp[5]) ? node57929 : node57910;
													assign node57910 = (inp[12]) ? node57918 : node57911;
														assign node57911 = (inp[14]) ? node57913 : 4'b0100;
															assign node57913 = (inp[0]) ? 4'b0100 : node57914;
																assign node57914 = (inp[15]) ? 4'b0100 : 4'b0110;
														assign node57918 = (inp[14]) ? node57924 : node57919;
															assign node57919 = (inp[15]) ? node57921 : 4'b0110;
																assign node57921 = (inp[0]) ? 4'b0110 : 4'b0100;
															assign node57924 = (inp[15]) ? node57926 : 4'b0100;
																assign node57926 = (inp[0]) ? 4'b0110 : 4'b0100;
													assign node57929 = (inp[12]) ? node57937 : node57930;
														assign node57930 = (inp[15]) ? node57934 : node57931;
															assign node57931 = (inp[0]) ? 4'b0110 : 4'b0100;
															assign node57934 = (inp[0]) ? 4'b0100 : 4'b0110;
														assign node57937 = (inp[15]) ? node57941 : node57938;
															assign node57938 = (inp[0]) ? 4'b0110 : 4'b0100;
															assign node57941 = (inp[0]) ? 4'b0100 : 4'b0110;
												assign node57944 = (inp[12]) ? node57952 : node57945;
													assign node57945 = (inp[15]) ? node57949 : node57946;
														assign node57946 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node57949 = (inp[0]) ? 4'b0100 : 4'b0110;
													assign node57952 = (inp[0]) ? node57956 : node57953;
														assign node57953 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node57956 = (inp[15]) ? 4'b0100 : 4'b0110;
										assign node57959 = (inp[9]) ? node58023 : node57960;
											assign node57960 = (inp[12]) ? node58000 : node57961;
												assign node57961 = (inp[5]) ? node57977 : node57962;
													assign node57962 = (inp[15]) ? node57970 : node57963;
														assign node57963 = (inp[14]) ? node57965 : 4'b0110;
															assign node57965 = (inp[3]) ? node57967 : 4'b0110;
																assign node57967 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node57970 = (inp[3]) ? node57974 : node57971;
															assign node57971 = (inp[0]) ? 4'b0110 : 4'b0100;
															assign node57974 = (inp[0]) ? 4'b0100 : 4'b0110;
													assign node57977 = (inp[3]) ? node57987 : node57978;
														assign node57978 = (inp[14]) ? node57984 : node57979;
															assign node57979 = (inp[0]) ? node57981 : 4'b0110;
																assign node57981 = (inp[15]) ? 4'b0100 : 4'b0110;
															assign node57984 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node57987 = (inp[14]) ? node57995 : node57988;
															assign node57988 = (inp[0]) ? node57992 : node57989;
																assign node57989 = (inp[15]) ? 4'b0110 : 4'b0100;
																assign node57992 = (inp[15]) ? 4'b0100 : 4'b0110;
															assign node57995 = (inp[0]) ? node57997 : 4'b0100;
																assign node57997 = (inp[15]) ? 4'b0100 : 4'b0110;
												assign node58000 = (inp[0]) ? node58012 : node58001;
													assign node58001 = (inp[15]) ? node58007 : node58002;
														assign node58002 = (inp[3]) ? 4'b0100 : node58003;
															assign node58003 = (inp[5]) ? 4'b0100 : 4'b0110;
														assign node58007 = (inp[5]) ? 4'b0110 : node58008;
															assign node58008 = (inp[14]) ? 4'b0100 : 4'b0110;
													assign node58012 = (inp[15]) ? node58018 : node58013;
														assign node58013 = (inp[3]) ? 4'b0110 : node58014;
															assign node58014 = (inp[5]) ? 4'b0110 : 4'b0100;
														assign node58018 = (inp[3]) ? 4'b0100 : node58019;
															assign node58019 = (inp[5]) ? 4'b0100 : 4'b0110;
											assign node58023 = (inp[15]) ? node58033 : node58024;
												assign node58024 = (inp[0]) ? node58028 : node58025;
													assign node58025 = (inp[5]) ? 4'b0000 : 4'b0010;
													assign node58028 = (inp[5]) ? 4'b0010 : node58029;
														assign node58029 = (inp[3]) ? 4'b0010 : 4'b0000;
												assign node58033 = (inp[0]) ? node58039 : node58034;
													assign node58034 = (inp[5]) ? 4'b0010 : node58035;
														assign node58035 = (inp[3]) ? 4'b0010 : 4'b0000;
													assign node58039 = (inp[3]) ? 4'b0000 : node58040;
														assign node58040 = (inp[5]) ? 4'b0000 : 4'b0010;
					assign node58044 = (inp[1]) ? node59688 : node58045;
						assign node58045 = (inp[8]) ? node58827 : node58046;
							assign node58046 = (inp[7]) ? node58466 : node58047;
								assign node58047 = (inp[14]) ? node58225 : node58048;
									assign node58048 = (inp[2]) ? node58136 : node58049;
										assign node58049 = (inp[5]) ? node58097 : node58050;
											assign node58050 = (inp[4]) ? node58072 : node58051;
												assign node58051 = (inp[9]) ? node58059 : node58052;
													assign node58052 = (inp[0]) ? node58056 : node58053;
														assign node58053 = (inp[15]) ? 4'b1001 : 4'b1011;
														assign node58056 = (inp[15]) ? 4'b1011 : 4'b1001;
													assign node58059 = (inp[15]) ? node58067 : node58060;
														assign node58060 = (inp[3]) ? node58064 : node58061;
															assign node58061 = (inp[0]) ? 4'b1101 : 4'b1111;
															assign node58064 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node58067 = (inp[3]) ? node58069 : 4'b1111;
															assign node58069 = (inp[0]) ? 4'b1101 : 4'b1111;
												assign node58072 = (inp[9]) ? node58086 : node58073;
													assign node58073 = (inp[0]) ? node58079 : node58074;
														assign node58074 = (inp[15]) ? node58076 : 4'b1111;
															assign node58076 = (inp[3]) ? 4'b1111 : 4'b1101;
														assign node58079 = (inp[3]) ? node58083 : node58080;
															assign node58080 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node58083 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node58086 = (inp[3]) ? node58092 : node58087;
														assign node58087 = (inp[0]) ? node58089 : 4'b1011;
															assign node58089 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node58092 = (inp[15]) ? 4'b1001 : node58093;
															assign node58093 = (inp[0]) ? 4'b1011 : 4'b1001;
											assign node58097 = (inp[4]) ? node58121 : node58098;
												assign node58098 = (inp[9]) ? node58108 : node58099;
													assign node58099 = (inp[0]) ? 4'b1001 : node58100;
														assign node58100 = (inp[3]) ? node58104 : node58101;
															assign node58101 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node58104 = (inp[15]) ? 4'b1011 : 4'b1001;
													assign node58108 = (inp[12]) ? node58114 : node58109;
														assign node58109 = (inp[0]) ? node58111 : 4'b1111;
															assign node58111 = (inp[15]) ? 4'b1101 : 4'b1111;
														assign node58114 = (inp[0]) ? node58118 : node58115;
															assign node58115 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node58118 = (inp[15]) ? 4'b1101 : 4'b1111;
												assign node58121 = (inp[9]) ? node58129 : node58122;
													assign node58122 = (inp[0]) ? node58126 : node58123;
														assign node58123 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node58126 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node58129 = (inp[15]) ? node58133 : node58130;
														assign node58130 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node58133 = (inp[0]) ? 4'b1001 : 4'b1011;
										assign node58136 = (inp[0]) ? node58180 : node58137;
											assign node58137 = (inp[5]) ? node58163 : node58138;
												assign node58138 = (inp[15]) ? node58152 : node58139;
													assign node58139 = (inp[3]) ? node58145 : node58140;
														assign node58140 = (inp[4]) ? 4'b1010 : node58141;
															assign node58141 = (inp[9]) ? 4'b1110 : 4'b1010;
														assign node58145 = (inp[9]) ? node58149 : node58146;
															assign node58146 = (inp[4]) ? 4'b1100 : 4'b1010;
															assign node58149 = (inp[4]) ? 4'b1000 : 4'b1100;
													assign node58152 = (inp[3]) ? node58158 : node58153;
														assign node58153 = (inp[9]) ? 4'b1000 : node58154;
															assign node58154 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node58158 = (inp[4]) ? node58160 : 4'b1000;
															assign node58160 = (inp[9]) ? 4'b1010 : 4'b1110;
												assign node58163 = (inp[15]) ? node58171 : node58164;
													assign node58164 = (inp[4]) ? node58168 : node58165;
														assign node58165 = (inp[9]) ? 4'b1100 : 4'b1010;
														assign node58168 = (inp[9]) ? 4'b1000 : 4'b1100;
													assign node58171 = (inp[4]) ? node58177 : node58172;
														assign node58172 = (inp[9]) ? 4'b1110 : node58173;
															assign node58173 = (inp[3]) ? 4'b1010 : 4'b1000;
														assign node58177 = (inp[9]) ? 4'b1010 : 4'b1110;
											assign node58180 = (inp[15]) ? node58198 : node58181;
												assign node58181 = (inp[9]) ? node58191 : node58182;
													assign node58182 = (inp[4]) ? node58186 : node58183;
														assign node58183 = (inp[12]) ? 4'b1000 : 4'b1010;
														assign node58186 = (inp[3]) ? 4'b1110 : node58187;
															assign node58187 = (inp[5]) ? 4'b1110 : 4'b1100;
													assign node58191 = (inp[4]) ? node58193 : 4'b1110;
														assign node58193 = (inp[3]) ? 4'b1010 : node58194;
															assign node58194 = (inp[5]) ? 4'b1010 : 4'b1000;
												assign node58198 = (inp[5]) ? node58210 : node58199;
													assign node58199 = (inp[9]) ? node58203 : node58200;
														assign node58200 = (inp[4]) ? 4'b1110 : 4'b1010;
														assign node58203 = (inp[4]) ? node58207 : node58204;
															assign node58204 = (inp[3]) ? 4'b1100 : 4'b1110;
															assign node58207 = (inp[3]) ? 4'b1000 : 4'b1010;
													assign node58210 = (inp[12]) ? node58218 : node58211;
														assign node58211 = (inp[9]) ? node58215 : node58212;
															assign node58212 = (inp[4]) ? 4'b1100 : 4'b1000;
															assign node58215 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node58218 = (inp[9]) ? node58222 : node58219;
															assign node58219 = (inp[3]) ? 4'b1000 : 4'b1010;
															assign node58222 = (inp[4]) ? 4'b1000 : 4'b1100;
									assign node58225 = (inp[3]) ? node58339 : node58226;
										assign node58226 = (inp[12]) ? node58290 : node58227;
											assign node58227 = (inp[2]) ? node58261 : node58228;
												assign node58228 = (inp[9]) ? node58242 : node58229;
													assign node58229 = (inp[4]) ? node58231 : 4'b1000;
														assign node58231 = (inp[5]) ? node58237 : node58232;
															assign node58232 = (inp[15]) ? 4'b1100 : node58233;
																assign node58233 = (inp[0]) ? 4'b1100 : 4'b1110;
															assign node58237 = (inp[0]) ? 4'b1110 : node58238;
																assign node58238 = (inp[15]) ? 4'b1110 : 4'b1100;
													assign node58242 = (inp[4]) ? node58252 : node58243;
														assign node58243 = (inp[0]) ? 4'b1110 : node58244;
															assign node58244 = (inp[5]) ? node58248 : node58245;
																assign node58245 = (inp[15]) ? 4'b1100 : 4'b1110;
																assign node58248 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node58252 = (inp[15]) ? 4'b1010 : node58253;
															assign node58253 = (inp[0]) ? node58257 : node58254;
																assign node58254 = (inp[5]) ? 4'b1000 : 4'b1010;
																assign node58257 = (inp[5]) ? 4'b1010 : 4'b1000;
												assign node58261 = (inp[9]) ? node58277 : node58262;
													assign node58262 = (inp[4]) ? node58268 : node58263;
														assign node58263 = (inp[15]) ? node58265 : 4'b1010;
															assign node58265 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node58268 = (inp[0]) ? node58270 : 4'b1110;
															assign node58270 = (inp[5]) ? node58274 : node58271;
																assign node58271 = (inp[15]) ? 4'b1110 : 4'b1100;
																assign node58274 = (inp[15]) ? 4'b1100 : 4'b1110;
													assign node58277 = (inp[4]) ? node58287 : node58278;
														assign node58278 = (inp[5]) ? 4'b1110 : node58279;
															assign node58279 = (inp[0]) ? node58283 : node58280;
																assign node58280 = (inp[15]) ? 4'b1100 : 4'b1110;
																assign node58283 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node58287 = (inp[15]) ? 4'b1010 : 4'b1000;
											assign node58290 = (inp[0]) ? node58314 : node58291;
												assign node58291 = (inp[15]) ? node58303 : node58292;
													assign node58292 = (inp[5]) ? node58298 : node58293;
														assign node58293 = (inp[4]) ? 4'b1010 : node58294;
															assign node58294 = (inp[9]) ? 4'b1110 : 4'b1010;
														assign node58298 = (inp[9]) ? 4'b1100 : node58299;
															assign node58299 = (inp[4]) ? 4'b1100 : 4'b1010;
													assign node58303 = (inp[5]) ? node58309 : node58304;
														assign node58304 = (inp[9]) ? node58306 : 4'b1100;
															assign node58306 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node58309 = (inp[4]) ? node58311 : 4'b1000;
															assign node58311 = (inp[9]) ? 4'b1010 : 4'b1110;
												assign node58314 = (inp[15]) ? node58328 : node58315;
													assign node58315 = (inp[5]) ? node58323 : node58316;
														assign node58316 = (inp[9]) ? node58320 : node58317;
															assign node58317 = (inp[4]) ? 4'b1100 : 4'b1000;
															assign node58320 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node58323 = (inp[4]) ? 4'b1110 : node58324;
															assign node58324 = (inp[9]) ? 4'b1110 : 4'b1000;
													assign node58328 = (inp[5]) ? node58334 : node58329;
														assign node58329 = (inp[9]) ? node58331 : 4'b1110;
															assign node58331 = (inp[4]) ? 4'b1010 : 4'b1110;
														assign node58334 = (inp[9]) ? node58336 : 4'b1100;
															assign node58336 = (inp[4]) ? 4'b1000 : 4'b1100;
										assign node58339 = (inp[2]) ? node58411 : node58340;
											assign node58340 = (inp[12]) ? node58374 : node58341;
												assign node58341 = (inp[9]) ? node58361 : node58342;
													assign node58342 = (inp[4]) ? node58354 : node58343;
														assign node58343 = (inp[0]) ? node58349 : node58344;
															assign node58344 = (inp[15]) ? 4'b1010 : node58345;
																assign node58345 = (inp[5]) ? 4'b1000 : 4'b1010;
															assign node58349 = (inp[5]) ? node58351 : 4'b1000;
																assign node58351 = (inp[15]) ? 4'b1000 : 4'b1010;
														assign node58354 = (inp[0]) ? node58358 : node58355;
															assign node58355 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node58358 = (inp[15]) ? 4'b1100 : 4'b1110;
													assign node58361 = (inp[4]) ? node58367 : node58362;
														assign node58362 = (inp[0]) ? 4'b1110 : node58363;
															assign node58363 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node58367 = (inp[0]) ? node58371 : node58368;
															assign node58368 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node58371 = (inp[15]) ? 4'b1000 : 4'b1010;
												assign node58374 = (inp[15]) ? node58392 : node58375;
													assign node58375 = (inp[0]) ? node58383 : node58376;
														assign node58376 = (inp[4]) ? node58380 : node58377;
															assign node58377 = (inp[5]) ? 4'b1000 : 4'b1010;
															assign node58380 = (inp[9]) ? 4'b1000 : 4'b1100;
														assign node58383 = (inp[9]) ? node58389 : node58384;
															assign node58384 = (inp[4]) ? 4'b1110 : node58385;
																assign node58385 = (inp[5]) ? 4'b1010 : 4'b1000;
															assign node58389 = (inp[4]) ? 4'b1010 : 4'b1110;
													assign node58392 = (inp[0]) ? node58408 : node58393;
														assign node58393 = (inp[5]) ? node58401 : node58394;
															assign node58394 = (inp[9]) ? node58398 : node58395;
																assign node58395 = (inp[4]) ? 4'b1110 : 4'b1000;
																assign node58398 = (inp[4]) ? 4'b1010 : 4'b1110;
															assign node58401 = (inp[9]) ? node58405 : node58402;
																assign node58402 = (inp[4]) ? 4'b1110 : 4'b1010;
																assign node58405 = (inp[4]) ? 4'b1010 : 4'b1110;
														assign node58408 = (inp[9]) ? 4'b1000 : 4'b1010;
											assign node58411 = (inp[5]) ? node58439 : node58412;
												assign node58412 = (inp[0]) ? node58424 : node58413;
													assign node58413 = (inp[15]) ? node58419 : node58414;
														assign node58414 = (inp[9]) ? node58416 : 4'b1100;
															assign node58416 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node58419 = (inp[9]) ? node58421 : 4'b1000;
															assign node58421 = (inp[4]) ? 4'b1010 : 4'b1110;
													assign node58424 = (inp[15]) ? node58432 : node58425;
														assign node58425 = (inp[9]) ? node58429 : node58426;
															assign node58426 = (inp[4]) ? 4'b1110 : 4'b1000;
															assign node58429 = (inp[4]) ? 4'b1010 : 4'b1110;
														assign node58432 = (inp[9]) ? node58436 : node58433;
															assign node58433 = (inp[4]) ? 4'b1100 : 4'b1010;
															assign node58436 = (inp[4]) ? 4'b1000 : 4'b1100;
												assign node58439 = (inp[0]) ? node58453 : node58440;
													assign node58440 = (inp[15]) ? node58446 : node58441;
														assign node58441 = (inp[4]) ? 4'b1100 : node58442;
															assign node58442 = (inp[9]) ? 4'b1100 : 4'b1000;
														assign node58446 = (inp[9]) ? node58450 : node58447;
															assign node58447 = (inp[4]) ? 4'b1110 : 4'b1010;
															assign node58450 = (inp[4]) ? 4'b1010 : 4'b1110;
													assign node58453 = (inp[15]) ? node58459 : node58454;
														assign node58454 = (inp[4]) ? node58456 : 4'b1110;
															assign node58456 = (inp[9]) ? 4'b1010 : 4'b1110;
														assign node58459 = (inp[12]) ? node58461 : 4'b1000;
															assign node58461 = (inp[4]) ? node58463 : 4'b1000;
																assign node58463 = (inp[9]) ? 4'b1000 : 4'b1100;
								assign node58466 = (inp[14]) ? node58702 : node58467;
									assign node58467 = (inp[2]) ? node58567 : node58468;
										assign node58468 = (inp[15]) ? node58524 : node58469;
											assign node58469 = (inp[0]) ? node58499 : node58470;
												assign node58470 = (inp[5]) ? node58488 : node58471;
													assign node58471 = (inp[3]) ? node58483 : node58472;
														assign node58472 = (inp[12]) ? node58478 : node58473;
															assign node58473 = (inp[9]) ? node58475 : 4'b1110;
																assign node58475 = (inp[4]) ? 4'b1010 : 4'b1110;
															assign node58478 = (inp[9]) ? 4'b1010 : node58479;
																assign node58479 = (inp[4]) ? 4'b1110 : 4'b1010;
														assign node58483 = (inp[4]) ? node58485 : 4'b1010;
															assign node58485 = (inp[9]) ? 4'b1000 : 4'b1100;
													assign node58488 = (inp[12]) ? 4'b1100 : node58489;
														assign node58489 = (inp[3]) ? 4'b1000 : node58490;
															assign node58490 = (inp[4]) ? node58494 : node58491;
																assign node58491 = (inp[9]) ? 4'b1100 : 4'b1010;
																assign node58494 = (inp[9]) ? 4'b1000 : 4'b1100;
												assign node58499 = (inp[3]) ? node58515 : node58500;
													assign node58500 = (inp[5]) ? node58508 : node58501;
														assign node58501 = (inp[9]) ? node58505 : node58502;
															assign node58502 = (inp[4]) ? 4'b1100 : 4'b1000;
															assign node58505 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node58508 = (inp[4]) ? node58512 : node58509;
															assign node58509 = (inp[9]) ? 4'b1110 : 4'b1000;
															assign node58512 = (inp[9]) ? 4'b1010 : 4'b1110;
													assign node58515 = (inp[9]) ? node58521 : node58516;
														assign node58516 = (inp[4]) ? 4'b1110 : node58517;
															assign node58517 = (inp[5]) ? 4'b1010 : 4'b1000;
														assign node58521 = (inp[4]) ? 4'b1010 : 4'b1110;
											assign node58524 = (inp[0]) ? node58550 : node58525;
												assign node58525 = (inp[5]) ? node58541 : node58526;
													assign node58526 = (inp[3]) ? node58534 : node58527;
														assign node58527 = (inp[9]) ? node58531 : node58528;
															assign node58528 = (inp[4]) ? 4'b1100 : 4'b1000;
															assign node58531 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node58534 = (inp[9]) ? node58538 : node58535;
															assign node58535 = (inp[4]) ? 4'b1110 : 4'b1000;
															assign node58538 = (inp[4]) ? 4'b1010 : 4'b1110;
													assign node58541 = (inp[4]) ? node58547 : node58542;
														assign node58542 = (inp[9]) ? 4'b1110 : node58543;
															assign node58543 = (inp[12]) ? 4'b1000 : 4'b1010;
														assign node58547 = (inp[9]) ? 4'b1010 : 4'b1110;
												assign node58550 = (inp[3]) ? node58562 : node58551;
													assign node58551 = (inp[5]) ? node58557 : node58552;
														assign node58552 = (inp[12]) ? node58554 : 4'b1010;
															assign node58554 = (inp[9]) ? 4'b1010 : 4'b1110;
														assign node58557 = (inp[4]) ? node58559 : 4'b1010;
															assign node58559 = (inp[9]) ? 4'b1000 : 4'b1100;
													assign node58562 = (inp[4]) ? node58564 : 4'b1100;
														assign node58564 = (inp[9]) ? 4'b1000 : 4'b1100;
										assign node58567 = (inp[12]) ? node58637 : node58568;
											assign node58568 = (inp[5]) ? node58606 : node58569;
												assign node58569 = (inp[0]) ? node58589 : node58570;
													assign node58570 = (inp[15]) ? node58578 : node58571;
														assign node58571 = (inp[3]) ? node58573 : 4'b0111;
															assign node58573 = (inp[4]) ? node58575 : 4'b0101;
																assign node58575 = (inp[9]) ? 4'b0001 : 4'b0101;
														assign node58578 = (inp[3]) ? node58586 : node58579;
															assign node58579 = (inp[9]) ? node58583 : node58580;
																assign node58580 = (inp[4]) ? 4'b0101 : 4'b0001;
																assign node58583 = (inp[4]) ? 4'b0001 : 4'b0101;
															assign node58586 = (inp[4]) ? 4'b0111 : 4'b0001;
													assign node58589 = (inp[9]) ? node58597 : node58590;
														assign node58590 = (inp[4]) ? node58592 : 4'b0011;
															assign node58592 = (inp[3]) ? 4'b0101 : node58593;
																assign node58593 = (inp[15]) ? 4'b0111 : 4'b0101;
														assign node58597 = (inp[4]) ? 4'b0011 : node58598;
															assign node58598 = (inp[15]) ? node58602 : node58599;
																assign node58599 = (inp[3]) ? 4'b0111 : 4'b0101;
																assign node58602 = (inp[3]) ? 4'b0101 : 4'b0111;
												assign node58606 = (inp[4]) ? node58616 : node58607;
													assign node58607 = (inp[9]) ? 4'b0101 : node58608;
														assign node58608 = (inp[0]) ? 4'b0001 : node58609;
															assign node58609 = (inp[15]) ? node58611 : 4'b0011;
																assign node58611 = (inp[3]) ? 4'b0011 : 4'b0001;
													assign node58616 = (inp[9]) ? node58624 : node58617;
														assign node58617 = (inp[3]) ? 4'b0111 : node58618;
															assign node58618 = (inp[0]) ? 4'b0101 : node58619;
																assign node58619 = (inp[15]) ? 4'b0111 : 4'b0101;
														assign node58624 = (inp[3]) ? node58632 : node58625;
															assign node58625 = (inp[0]) ? node58629 : node58626;
																assign node58626 = (inp[15]) ? 4'b0011 : 4'b0001;
																assign node58629 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node58632 = (inp[15]) ? node58634 : 4'b0011;
																assign node58634 = (inp[0]) ? 4'b0001 : 4'b0011;
											assign node58637 = (inp[15]) ? node58671 : node58638;
												assign node58638 = (inp[0]) ? node58650 : node58639;
													assign node58639 = (inp[3]) ? node58643 : node58640;
														assign node58640 = (inp[9]) ? 4'b0111 : 4'b0011;
														assign node58643 = (inp[4]) ? node58647 : node58644;
															assign node58644 = (inp[9]) ? 4'b0101 : 4'b0001;
															assign node58647 = (inp[9]) ? 4'b0001 : 4'b0101;
													assign node58650 = (inp[3]) ? node58658 : node58651;
														assign node58651 = (inp[9]) ? 4'b0111 : node58652;
															assign node58652 = (inp[4]) ? node58654 : 4'b0001;
																assign node58654 = (inp[5]) ? 4'b0111 : 4'b0101;
														assign node58658 = (inp[5]) ? node58664 : node58659;
															assign node58659 = (inp[9]) ? node58661 : 4'b0111;
																assign node58661 = (inp[4]) ? 4'b0011 : 4'b0111;
															assign node58664 = (inp[4]) ? node58668 : node58665;
																assign node58665 = (inp[9]) ? 4'b0111 : 4'b0011;
																assign node58668 = (inp[9]) ? 4'b0011 : 4'b0111;
												assign node58671 = (inp[0]) ? node58687 : node58672;
													assign node58672 = (inp[5]) ? node58678 : node58673;
														assign node58673 = (inp[3]) ? node58675 : 4'b0101;
															assign node58675 = (inp[4]) ? 4'b0011 : 4'b0001;
														assign node58678 = (inp[3]) ? node58680 : 4'b0111;
															assign node58680 = (inp[4]) ? node58684 : node58681;
																assign node58681 = (inp[9]) ? 4'b0111 : 4'b0011;
																assign node58684 = (inp[9]) ? 4'b0011 : 4'b0111;
													assign node58687 = (inp[5]) ? node58695 : node58688;
														assign node58688 = (inp[9]) ? node58692 : node58689;
															assign node58689 = (inp[3]) ? 4'b0011 : 4'b0111;
															assign node58692 = (inp[3]) ? 4'b0001 : 4'b0011;
														assign node58695 = (inp[9]) ? node58699 : node58696;
															assign node58696 = (inp[3]) ? 4'b0001 : 4'b0011;
															assign node58699 = (inp[4]) ? 4'b0001 : 4'b0101;
									assign node58702 = (inp[15]) ? node58768 : node58703;
										assign node58703 = (inp[0]) ? node58737 : node58704;
											assign node58704 = (inp[5]) ? node58728 : node58705;
												assign node58705 = (inp[3]) ? node58721 : node58706;
													assign node58706 = (inp[2]) ? node58714 : node58707;
														assign node58707 = (inp[4]) ? node58711 : node58708;
															assign node58708 = (inp[9]) ? 4'b0111 : 4'b0011;
															assign node58711 = (inp[9]) ? 4'b0011 : 4'b0111;
														assign node58714 = (inp[9]) ? node58718 : node58715;
															assign node58715 = (inp[4]) ? 4'b0111 : 4'b0011;
															assign node58718 = (inp[4]) ? 4'b0011 : 4'b0111;
													assign node58721 = (inp[4]) ? node58725 : node58722;
														assign node58722 = (inp[2]) ? 4'b0101 : 4'b0011;
														assign node58725 = (inp[9]) ? 4'b0001 : 4'b0101;
												assign node58728 = (inp[9]) ? node58734 : node58729;
													assign node58729 = (inp[4]) ? 4'b0101 : node58730;
														assign node58730 = (inp[3]) ? 4'b0001 : 4'b0011;
													assign node58734 = (inp[4]) ? 4'b0001 : 4'b0101;
											assign node58737 = (inp[5]) ? node58759 : node58738;
												assign node58738 = (inp[3]) ? node58752 : node58739;
													assign node58739 = (inp[2]) ? node58745 : node58740;
														assign node58740 = (inp[12]) ? node58742 : 4'b0001;
															assign node58742 = (inp[9]) ? 4'b0101 : 4'b0001;
														assign node58745 = (inp[12]) ? node58747 : 4'b0101;
															assign node58747 = (inp[9]) ? node58749 : 4'b0001;
																assign node58749 = (inp[4]) ? 4'b0001 : 4'b0101;
													assign node58752 = (inp[4]) ? node58756 : node58753;
														assign node58753 = (inp[9]) ? 4'b0111 : 4'b0001;
														assign node58756 = (inp[9]) ? 4'b0011 : 4'b0111;
												assign node58759 = (inp[4]) ? node58765 : node58760;
													assign node58760 = (inp[9]) ? 4'b0111 : node58761;
														assign node58761 = (inp[3]) ? 4'b0011 : 4'b0001;
													assign node58765 = (inp[9]) ? 4'b0011 : 4'b0111;
										assign node58768 = (inp[0]) ? node58794 : node58769;
											assign node58769 = (inp[5]) ? node58785 : node58770;
												assign node58770 = (inp[3]) ? node58778 : node58771;
													assign node58771 = (inp[4]) ? node58775 : node58772;
														assign node58772 = (inp[9]) ? 4'b0101 : 4'b0001;
														assign node58775 = (inp[9]) ? 4'b0001 : 4'b0101;
													assign node58778 = (inp[4]) ? node58782 : node58779;
														assign node58779 = (inp[9]) ? 4'b0111 : 4'b0001;
														assign node58782 = (inp[9]) ? 4'b0011 : 4'b0111;
												assign node58785 = (inp[4]) ? node58791 : node58786;
													assign node58786 = (inp[9]) ? 4'b0111 : node58787;
														assign node58787 = (inp[3]) ? 4'b0011 : 4'b0001;
													assign node58791 = (inp[9]) ? 4'b0011 : 4'b0111;
											assign node58794 = (inp[5]) ? node58804 : node58795;
												assign node58795 = (inp[9]) ? node58801 : node58796;
													assign node58796 = (inp[4]) ? node58798 : 4'b0011;
														assign node58798 = (inp[3]) ? 4'b0101 : 4'b0111;
													assign node58801 = (inp[3]) ? 4'b0101 : 4'b0111;
												assign node58804 = (inp[3]) ? node58812 : node58805;
													assign node58805 = (inp[4]) ? node58809 : node58806;
														assign node58806 = (inp[9]) ? 4'b0101 : 4'b0011;
														assign node58809 = (inp[9]) ? 4'b0001 : 4'b0101;
													assign node58812 = (inp[12]) ? node58820 : node58813;
														assign node58813 = (inp[9]) ? node58817 : node58814;
															assign node58814 = (inp[4]) ? 4'b0101 : 4'b0001;
															assign node58817 = (inp[4]) ? 4'b0001 : 4'b0101;
														assign node58820 = (inp[4]) ? node58824 : node58821;
															assign node58821 = (inp[9]) ? 4'b0101 : 4'b0001;
															assign node58824 = (inp[9]) ? 4'b0001 : 4'b0101;
							assign node58827 = (inp[7]) ? node59211 : node58828;
								assign node58828 = (inp[14]) ? node59068 : node58829;
									assign node58829 = (inp[2]) ? node58925 : node58830;
										assign node58830 = (inp[5]) ? node58894 : node58831;
											assign node58831 = (inp[15]) ? node58869 : node58832;
												assign node58832 = (inp[0]) ? node58852 : node58833;
													assign node58833 = (inp[3]) ? node58845 : node58834;
														assign node58834 = (inp[12]) ? node58840 : node58835;
															assign node58835 = (inp[4]) ? 4'b1010 : node58836;
																assign node58836 = (inp[9]) ? 4'b1110 : 4'b1010;
															assign node58840 = (inp[9]) ? node58842 : 4'b1110;
																assign node58842 = (inp[4]) ? 4'b1010 : 4'b1110;
														assign node58845 = (inp[4]) ? node58849 : node58846;
															assign node58846 = (inp[9]) ? 4'b1100 : 4'b1010;
															assign node58849 = (inp[9]) ? 4'b1000 : 4'b1100;
													assign node58852 = (inp[3]) ? node58860 : node58853;
														assign node58853 = (inp[9]) ? node58857 : node58854;
															assign node58854 = (inp[4]) ? 4'b1100 : 4'b1000;
															assign node58857 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node58860 = (inp[12]) ? node58864 : node58861;
															assign node58861 = (inp[9]) ? 4'b1110 : 4'b1000;
															assign node58864 = (inp[9]) ? node58866 : 4'b1110;
																assign node58866 = (inp[4]) ? 4'b1010 : 4'b1110;
												assign node58869 = (inp[0]) ? node58883 : node58870;
													assign node58870 = (inp[3]) ? node58878 : node58871;
														assign node58871 = (inp[4]) ? node58875 : node58872;
															assign node58872 = (inp[9]) ? 4'b1100 : 4'b1000;
															assign node58875 = (inp[9]) ? 4'b1000 : 4'b1100;
														assign node58878 = (inp[9]) ? 4'b1110 : node58879;
															assign node58879 = (inp[4]) ? 4'b1110 : 4'b1000;
													assign node58883 = (inp[3]) ? node58889 : node58884;
														assign node58884 = (inp[12]) ? node58886 : 4'b1110;
															assign node58886 = (inp[4]) ? 4'b1010 : 4'b1110;
														assign node58889 = (inp[4]) ? node58891 : 4'b1010;
															assign node58891 = (inp[9]) ? 4'b1000 : 4'b1100;
											assign node58894 = (inp[9]) ? node58910 : node58895;
												assign node58895 = (inp[4]) ? node58903 : node58896;
													assign node58896 = (inp[3]) ? 4'b1010 : node58897;
														assign node58897 = (inp[15]) ? 4'b1010 : node58898;
															assign node58898 = (inp[0]) ? 4'b1000 : 4'b1010;
													assign node58903 = (inp[0]) ? node58907 : node58904;
														assign node58904 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node58907 = (inp[15]) ? 4'b1100 : 4'b1110;
												assign node58910 = (inp[4]) ? node58918 : node58911;
													assign node58911 = (inp[0]) ? node58915 : node58912;
														assign node58912 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node58915 = (inp[15]) ? 4'b1100 : 4'b1110;
													assign node58918 = (inp[15]) ? node58922 : node58919;
														assign node58919 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node58922 = (inp[0]) ? 4'b1000 : 4'b1010;
										assign node58925 = (inp[12]) ? node58987 : node58926;
											assign node58926 = (inp[9]) ? node58954 : node58927;
												assign node58927 = (inp[4]) ? node58937 : node58928;
													assign node58928 = (inp[15]) ? node58932 : node58929;
														assign node58929 = (inp[0]) ? 4'b0001 : 4'b0011;
														assign node58932 = (inp[0]) ? node58934 : 4'b0001;
															assign node58934 = (inp[5]) ? 4'b0001 : 4'b0011;
													assign node58937 = (inp[3]) ? 4'b0111 : node58938;
														assign node58938 = (inp[5]) ? node58946 : node58939;
															assign node58939 = (inp[0]) ? node58943 : node58940;
																assign node58940 = (inp[15]) ? 4'b0101 : 4'b0111;
																assign node58943 = (inp[15]) ? 4'b0111 : 4'b0101;
															assign node58946 = (inp[15]) ? node58950 : node58947;
																assign node58947 = (inp[0]) ? 4'b0111 : 4'b0101;
																assign node58950 = (inp[0]) ? 4'b0101 : 4'b0111;
												assign node58954 = (inp[4]) ? node58966 : node58955;
													assign node58955 = (inp[3]) ? node58961 : node58956;
														assign node58956 = (inp[15]) ? 4'b0111 : node58957;
															assign node58957 = (inp[5]) ? 4'b0101 : 4'b0111;
														assign node58961 = (inp[0]) ? node58963 : 4'b0101;
															assign node58963 = (inp[15]) ? 4'b0101 : 4'b0111;
													assign node58966 = (inp[5]) ? node58980 : node58967;
														assign node58967 = (inp[3]) ? node58973 : node58968;
															assign node58968 = (inp[15]) ? node58970 : 4'b0001;
																assign node58970 = (inp[0]) ? 4'b0011 : 4'b0001;
															assign node58973 = (inp[15]) ? node58977 : node58974;
																assign node58974 = (inp[0]) ? 4'b0011 : 4'b0001;
																assign node58977 = (inp[0]) ? 4'b0001 : 4'b0011;
														assign node58980 = (inp[15]) ? node58984 : node58981;
															assign node58981 = (inp[0]) ? 4'b0011 : 4'b0001;
															assign node58984 = (inp[0]) ? 4'b0001 : 4'b0011;
											assign node58987 = (inp[3]) ? node59025 : node58988;
												assign node58988 = (inp[9]) ? node59004 : node58989;
													assign node58989 = (inp[4]) ? node58997 : node58990;
														assign node58990 = (inp[15]) ? node58994 : node58991;
															assign node58991 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node58994 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node58997 = (inp[0]) ? node58999 : 4'b0101;
															assign node58999 = (inp[5]) ? 4'b0111 : node59000;
																assign node59000 = (inp[15]) ? 4'b0111 : 4'b0101;
													assign node59004 = (inp[4]) ? node59020 : node59005;
														assign node59005 = (inp[5]) ? node59013 : node59006;
															assign node59006 = (inp[15]) ? node59010 : node59007;
																assign node59007 = (inp[0]) ? 4'b0101 : 4'b0111;
																assign node59010 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node59013 = (inp[0]) ? node59017 : node59014;
																assign node59014 = (inp[15]) ? 4'b0111 : 4'b0101;
																assign node59017 = (inp[15]) ? 4'b0101 : 4'b0111;
														assign node59020 = (inp[15]) ? 4'b0001 : node59021;
															assign node59021 = (inp[5]) ? 4'b0011 : 4'b0001;
												assign node59025 = (inp[5]) ? node59045 : node59026;
													assign node59026 = (inp[9]) ? node59038 : node59027;
														assign node59027 = (inp[4]) ? node59033 : node59028;
															assign node59028 = (inp[0]) ? node59030 : 4'b0011;
																assign node59030 = (inp[15]) ? 4'b0011 : 4'b0001;
															assign node59033 = (inp[0]) ? 4'b0101 : node59034;
																assign node59034 = (inp[15]) ? 4'b0111 : 4'b0101;
														assign node59038 = (inp[4]) ? node59040 : 4'b0101;
															assign node59040 = (inp[15]) ? node59042 : 4'b0001;
																assign node59042 = (inp[0]) ? 4'b0001 : 4'b0011;
													assign node59045 = (inp[15]) ? node59059 : node59046;
														assign node59046 = (inp[0]) ? node59054 : node59047;
															assign node59047 = (inp[9]) ? node59051 : node59048;
																assign node59048 = (inp[4]) ? 4'b0101 : 4'b0001;
																assign node59051 = (inp[4]) ? 4'b0001 : 4'b0101;
															assign node59054 = (inp[4]) ? node59056 : 4'b0111;
																assign node59056 = (inp[9]) ? 4'b0011 : 4'b0111;
														assign node59059 = (inp[0]) ? node59061 : 4'b0111;
															assign node59061 = (inp[4]) ? node59065 : node59062;
																assign node59062 = (inp[9]) ? 4'b0101 : 4'b0001;
																assign node59065 = (inp[9]) ? 4'b0001 : 4'b0101;
									assign node59068 = (inp[0]) ? node59126 : node59069;
										assign node59069 = (inp[15]) ? node59101 : node59070;
											assign node59070 = (inp[5]) ? node59086 : node59071;
												assign node59071 = (inp[3]) ? node59079 : node59072;
													assign node59072 = (inp[4]) ? node59076 : node59073;
														assign node59073 = (inp[9]) ? 4'b0111 : 4'b0011;
														assign node59076 = (inp[9]) ? 4'b0011 : 4'b0111;
													assign node59079 = (inp[9]) ? node59083 : node59080;
														assign node59080 = (inp[4]) ? 4'b0101 : 4'b0011;
														assign node59083 = (inp[4]) ? 4'b0001 : 4'b0101;
												assign node59086 = (inp[3]) ? node59094 : node59087;
													assign node59087 = (inp[4]) ? node59091 : node59088;
														assign node59088 = (inp[9]) ? 4'b0101 : 4'b0011;
														assign node59091 = (inp[9]) ? 4'b0001 : 4'b0101;
													assign node59094 = (inp[4]) ? node59098 : node59095;
														assign node59095 = (inp[9]) ? 4'b0101 : 4'b0001;
														assign node59098 = (inp[9]) ? 4'b0001 : 4'b0101;
											assign node59101 = (inp[3]) ? node59117 : node59102;
												assign node59102 = (inp[5]) ? node59110 : node59103;
													assign node59103 = (inp[9]) ? node59107 : node59104;
														assign node59104 = (inp[4]) ? 4'b0101 : 4'b0001;
														assign node59107 = (inp[4]) ? 4'b0001 : 4'b0101;
													assign node59110 = (inp[9]) ? node59114 : node59111;
														assign node59111 = (inp[4]) ? 4'b0111 : 4'b0001;
														assign node59114 = (inp[4]) ? 4'b0011 : 4'b0111;
												assign node59117 = (inp[4]) ? node59123 : node59118;
													assign node59118 = (inp[9]) ? 4'b0111 : node59119;
														assign node59119 = (inp[5]) ? 4'b0011 : 4'b0001;
													assign node59123 = (inp[9]) ? 4'b0011 : 4'b0111;
										assign node59126 = (inp[15]) ? node59170 : node59127;
											assign node59127 = (inp[5]) ? node59153 : node59128;
												assign node59128 = (inp[3]) ? node59146 : node59129;
													assign node59129 = (inp[12]) ? node59137 : node59130;
														assign node59130 = (inp[9]) ? node59134 : node59131;
															assign node59131 = (inp[4]) ? 4'b0101 : 4'b0001;
															assign node59134 = (inp[4]) ? 4'b0001 : 4'b0101;
														assign node59137 = (inp[2]) ? node59143 : node59138;
															assign node59138 = (inp[9]) ? 4'b0101 : node59139;
																assign node59139 = (inp[4]) ? 4'b0101 : 4'b0001;
															assign node59143 = (inp[4]) ? 4'b0001 : 4'b0101;
													assign node59146 = (inp[9]) ? node59150 : node59147;
														assign node59147 = (inp[4]) ? 4'b0111 : 4'b0001;
														assign node59150 = (inp[4]) ? 4'b0011 : 4'b0111;
												assign node59153 = (inp[2]) ? node59161 : node59154;
													assign node59154 = (inp[4]) ? node59158 : node59155;
														assign node59155 = (inp[9]) ? 4'b0111 : 4'b0011;
														assign node59158 = (inp[9]) ? 4'b0011 : 4'b0111;
													assign node59161 = (inp[4]) ? node59167 : node59162;
														assign node59162 = (inp[9]) ? 4'b0111 : node59163;
															assign node59163 = (inp[3]) ? 4'b0011 : 4'b0001;
														assign node59167 = (inp[9]) ? 4'b0011 : 4'b0111;
											assign node59170 = (inp[5]) ? node59202 : node59171;
												assign node59171 = (inp[3]) ? node59195 : node59172;
													assign node59172 = (inp[12]) ? node59188 : node59173;
														assign node59173 = (inp[2]) ? node59181 : node59174;
															assign node59174 = (inp[9]) ? node59178 : node59175;
																assign node59175 = (inp[4]) ? 4'b0111 : 4'b0011;
																assign node59178 = (inp[4]) ? 4'b0011 : 4'b0111;
															assign node59181 = (inp[9]) ? node59185 : node59182;
																assign node59182 = (inp[4]) ? 4'b0111 : 4'b0011;
																assign node59185 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node59188 = (inp[2]) ? node59190 : 4'b0011;
															assign node59190 = (inp[9]) ? 4'b0011 : node59191;
																assign node59191 = (inp[4]) ? 4'b0111 : 4'b0011;
													assign node59195 = (inp[4]) ? node59199 : node59196;
														assign node59196 = (inp[9]) ? 4'b0101 : 4'b0011;
														assign node59199 = (inp[9]) ? 4'b0001 : 4'b0101;
												assign node59202 = (inp[9]) ? node59208 : node59203;
													assign node59203 = (inp[4]) ? 4'b0101 : node59204;
														assign node59204 = (inp[3]) ? 4'b0001 : 4'b0011;
													assign node59208 = (inp[4]) ? 4'b0001 : 4'b0101;
								assign node59211 = (inp[14]) ? node59467 : node59212;
									assign node59212 = (inp[2]) ? node59334 : node59213;
										assign node59213 = (inp[3]) ? node59267 : node59214;
											assign node59214 = (inp[4]) ? node59232 : node59215;
												assign node59215 = (inp[9]) ? node59223 : node59216;
													assign node59216 = (inp[0]) ? node59220 : node59217;
														assign node59217 = (inp[15]) ? 4'b0001 : 4'b0011;
														assign node59220 = (inp[15]) ? 4'b0011 : 4'b0001;
													assign node59223 = (inp[15]) ? 4'b0101 : node59224;
														assign node59224 = (inp[5]) ? node59228 : node59225;
															assign node59225 = (inp[0]) ? 4'b0101 : 4'b0111;
															assign node59228 = (inp[0]) ? 4'b0111 : 4'b0101;
												assign node59232 = (inp[9]) ? node59246 : node59233;
													assign node59233 = (inp[15]) ? node59239 : node59234;
														assign node59234 = (inp[0]) ? node59236 : 4'b0101;
															assign node59236 = (inp[5]) ? 4'b0111 : 4'b0101;
														assign node59239 = (inp[5]) ? node59243 : node59240;
															assign node59240 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node59243 = (inp[0]) ? 4'b0101 : 4'b0111;
													assign node59246 = (inp[5]) ? node59252 : node59247;
														assign node59247 = (inp[0]) ? 4'b0011 : node59248;
															assign node59248 = (inp[15]) ? 4'b0001 : 4'b0011;
														assign node59252 = (inp[12]) ? node59260 : node59253;
															assign node59253 = (inp[0]) ? node59257 : node59254;
																assign node59254 = (inp[15]) ? 4'b0011 : 4'b0001;
																assign node59257 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node59260 = (inp[15]) ? node59264 : node59261;
																assign node59261 = (inp[0]) ? 4'b0011 : 4'b0001;
																assign node59264 = (inp[0]) ? 4'b0001 : 4'b0011;
											assign node59267 = (inp[4]) ? node59305 : node59268;
												assign node59268 = (inp[9]) ? node59290 : node59269;
													assign node59269 = (inp[5]) ? node59277 : node59270;
														assign node59270 = (inp[0]) ? node59274 : node59271;
															assign node59271 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node59274 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node59277 = (inp[12]) ? node59285 : node59278;
															assign node59278 = (inp[0]) ? node59282 : node59279;
																assign node59279 = (inp[15]) ? 4'b0011 : 4'b0001;
																assign node59282 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node59285 = (inp[15]) ? node59287 : 4'b0001;
																assign node59287 = (inp[0]) ? 4'b0001 : 4'b0011;
													assign node59290 = (inp[5]) ? node59298 : node59291;
														assign node59291 = (inp[0]) ? node59295 : node59292;
															assign node59292 = (inp[15]) ? 4'b0111 : 4'b0101;
															assign node59295 = (inp[15]) ? 4'b0101 : 4'b0111;
														assign node59298 = (inp[15]) ? node59302 : node59299;
															assign node59299 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node59302 = (inp[0]) ? 4'b0101 : 4'b0111;
												assign node59305 = (inp[9]) ? node59327 : node59306;
													assign node59306 = (inp[12]) ? node59322 : node59307;
														assign node59307 = (inp[5]) ? node59315 : node59308;
															assign node59308 = (inp[15]) ? node59312 : node59309;
																assign node59309 = (inp[0]) ? 4'b0111 : 4'b0101;
																assign node59312 = (inp[0]) ? 4'b0101 : 4'b0111;
															assign node59315 = (inp[0]) ? node59319 : node59316;
																assign node59316 = (inp[15]) ? 4'b0111 : 4'b0101;
																assign node59319 = (inp[15]) ? 4'b0101 : 4'b0111;
														assign node59322 = (inp[0]) ? 4'b0111 : node59323;
															assign node59323 = (inp[5]) ? 4'b0111 : 4'b0101;
													assign node59327 = (inp[15]) ? node59331 : node59328;
														assign node59328 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node59331 = (inp[0]) ? 4'b0001 : 4'b0011;
										assign node59334 = (inp[3]) ? node59406 : node59335;
											assign node59335 = (inp[15]) ? node59361 : node59336;
												assign node59336 = (inp[9]) ? node59350 : node59337;
													assign node59337 = (inp[4]) ? node59341 : node59338;
														assign node59338 = (inp[0]) ? 4'b0000 : 4'b0010;
														assign node59341 = (inp[12]) ? node59343 : 4'b0110;
															assign node59343 = (inp[5]) ? node59347 : node59344;
																assign node59344 = (inp[0]) ? 4'b0100 : 4'b0110;
																assign node59347 = (inp[0]) ? 4'b0110 : 4'b0100;
													assign node59350 = (inp[4]) ? 4'b0000 : node59351;
														assign node59351 = (inp[12]) ? 4'b0100 : node59352;
															assign node59352 = (inp[0]) ? node59356 : node59353;
																assign node59353 = (inp[5]) ? 4'b0100 : 4'b0110;
																assign node59356 = (inp[5]) ? 4'b0110 : 4'b0100;
												assign node59361 = (inp[12]) ? node59385 : node59362;
													assign node59362 = (inp[0]) ? node59370 : node59363;
														assign node59363 = (inp[5]) ? node59365 : 4'b0100;
															assign node59365 = (inp[9]) ? node59367 : 4'b0110;
																assign node59367 = (inp[4]) ? 4'b0010 : 4'b0110;
														assign node59370 = (inp[5]) ? node59378 : node59371;
															assign node59371 = (inp[9]) ? node59375 : node59372;
																assign node59372 = (inp[4]) ? 4'b0110 : 4'b0010;
																assign node59375 = (inp[4]) ? 4'b0010 : 4'b0110;
															assign node59378 = (inp[9]) ? node59382 : node59379;
																assign node59379 = (inp[4]) ? 4'b0100 : 4'b0010;
																assign node59382 = (inp[4]) ? 4'b0000 : 4'b0100;
													assign node59385 = (inp[0]) ? node59395 : node59386;
														assign node59386 = (inp[4]) ? node59390 : node59387;
															assign node59387 = (inp[9]) ? 4'b0100 : 4'b0000;
															assign node59390 = (inp[5]) ? node59392 : 4'b0000;
																assign node59392 = (inp[9]) ? 4'b0010 : 4'b0110;
														assign node59395 = (inp[5]) ? node59403 : node59396;
															assign node59396 = (inp[9]) ? node59400 : node59397;
																assign node59397 = (inp[4]) ? 4'b0110 : 4'b0010;
																assign node59400 = (inp[4]) ? 4'b0010 : 4'b0110;
															assign node59403 = (inp[9]) ? 4'b0000 : 4'b0010;
											assign node59406 = (inp[12]) ? node59442 : node59407;
												assign node59407 = (inp[4]) ? node59423 : node59408;
													assign node59408 = (inp[9]) ? node59418 : node59409;
														assign node59409 = (inp[5]) ? node59411 : 4'b0010;
															assign node59411 = (inp[15]) ? node59415 : node59412;
																assign node59412 = (inp[0]) ? 4'b0010 : 4'b0000;
																assign node59415 = (inp[0]) ? 4'b0000 : 4'b0010;
														assign node59418 = (inp[15]) ? 4'b0100 : node59419;
															assign node59419 = (inp[0]) ? 4'b0110 : 4'b0100;
													assign node59423 = (inp[9]) ? node59429 : node59424;
														assign node59424 = (inp[15]) ? node59426 : 4'b0100;
															assign node59426 = (inp[0]) ? 4'b0100 : 4'b0110;
														assign node59429 = (inp[5]) ? node59437 : node59430;
															assign node59430 = (inp[0]) ? node59434 : node59431;
																assign node59431 = (inp[15]) ? 4'b0010 : 4'b0000;
																assign node59434 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node59437 = (inp[15]) ? 4'b0000 : node59438;
																assign node59438 = (inp[0]) ? 4'b0010 : 4'b0000;
												assign node59442 = (inp[5]) ? node59456 : node59443;
													assign node59443 = (inp[9]) ? node59451 : node59444;
														assign node59444 = (inp[4]) ? 4'b0100 : node59445;
															assign node59445 = (inp[15]) ? node59447 : 4'b0000;
																assign node59447 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node59451 = (inp[15]) ? node59453 : 4'b0010;
															assign node59453 = (inp[0]) ? 4'b0100 : 4'b0110;
													assign node59456 = (inp[4]) ? node59464 : node59457;
														assign node59457 = (inp[9]) ? 4'b0110 : node59458;
															assign node59458 = (inp[0]) ? 4'b0010 : node59459;
																assign node59459 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node59464 = (inp[9]) ? 4'b0010 : 4'b0110;
									assign node59467 = (inp[12]) ? node59545 : node59468;
										assign node59468 = (inp[9]) ? node59510 : node59469;
											assign node59469 = (inp[4]) ? node59485 : node59470;
												assign node59470 = (inp[0]) ? node59480 : node59471;
													assign node59471 = (inp[15]) ? node59477 : node59472;
														assign node59472 = (inp[5]) ? node59474 : 4'b0010;
															assign node59474 = (inp[3]) ? 4'b0000 : 4'b0010;
														assign node59477 = (inp[3]) ? 4'b0010 : 4'b0000;
													assign node59480 = (inp[15]) ? 4'b0010 : node59481;
														assign node59481 = (inp[5]) ? 4'b0010 : 4'b0000;
												assign node59485 = (inp[3]) ? node59505 : node59486;
													assign node59486 = (inp[2]) ? node59496 : node59487;
														assign node59487 = (inp[15]) ? 4'b0110 : node59488;
															assign node59488 = (inp[5]) ? node59492 : node59489;
																assign node59489 = (inp[0]) ? 4'b0100 : 4'b0110;
																assign node59492 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node59496 = (inp[15]) ? node59498 : 4'b0110;
															assign node59498 = (inp[0]) ? node59502 : node59499;
																assign node59499 = (inp[5]) ? 4'b0110 : 4'b0100;
																assign node59502 = (inp[5]) ? 4'b0100 : 4'b0110;
													assign node59505 = (inp[0]) ? 4'b0100 : node59506;
														assign node59506 = (inp[15]) ? 4'b0110 : 4'b0100;
											assign node59510 = (inp[4]) ? node59528 : node59511;
												assign node59511 = (inp[15]) ? node59521 : node59512;
													assign node59512 = (inp[0]) ? node59516 : node59513;
														assign node59513 = (inp[5]) ? 4'b0100 : 4'b0110;
														assign node59516 = (inp[3]) ? 4'b0110 : node59517;
															assign node59517 = (inp[5]) ? 4'b0110 : 4'b0100;
													assign node59521 = (inp[0]) ? 4'b0100 : node59522;
														assign node59522 = (inp[3]) ? 4'b0110 : node59523;
															assign node59523 = (inp[5]) ? 4'b0110 : 4'b0100;
												assign node59528 = (inp[0]) ? node59536 : node59529;
													assign node59529 = (inp[3]) ? 4'b0010 : node59530;
														assign node59530 = (inp[5]) ? 4'b0010 : node59531;
															assign node59531 = (inp[15]) ? 4'b0000 : 4'b0010;
													assign node59536 = (inp[5]) ? node59542 : node59537;
														assign node59537 = (inp[3]) ? 4'b0010 : node59538;
															assign node59538 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node59542 = (inp[15]) ? 4'b0000 : 4'b0010;
										assign node59545 = (inp[2]) ? node59615 : node59546;
											assign node59546 = (inp[9]) ? node59584 : node59547;
												assign node59547 = (inp[4]) ? node59567 : node59548;
													assign node59548 = (inp[0]) ? node59560 : node59549;
														assign node59549 = (inp[15]) ? node59555 : node59550;
															assign node59550 = (inp[3]) ? node59552 : 4'b0010;
																assign node59552 = (inp[5]) ? 4'b0000 : 4'b0010;
															assign node59555 = (inp[5]) ? node59557 : 4'b0000;
																assign node59557 = (inp[3]) ? 4'b0010 : 4'b0000;
														assign node59560 = (inp[15]) ? node59562 : 4'b0000;
															assign node59562 = (inp[5]) ? node59564 : 4'b0010;
																assign node59564 = (inp[3]) ? 4'b0000 : 4'b0010;
													assign node59567 = (inp[3]) ? node59577 : node59568;
														assign node59568 = (inp[15]) ? 4'b0110 : node59569;
															assign node59569 = (inp[5]) ? node59573 : node59570;
																assign node59570 = (inp[0]) ? 4'b0100 : 4'b0110;
																assign node59573 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node59577 = (inp[15]) ? node59581 : node59578;
															assign node59578 = (inp[0]) ? 4'b0110 : 4'b0100;
															assign node59581 = (inp[0]) ? 4'b0100 : 4'b0110;
												assign node59584 = (inp[4]) ? node59596 : node59585;
													assign node59585 = (inp[15]) ? node59591 : node59586;
														assign node59586 = (inp[3]) ? node59588 : 4'b0100;
															assign node59588 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node59591 = (inp[0]) ? 4'b0100 : node59592;
															assign node59592 = (inp[5]) ? 4'b0110 : 4'b0100;
													assign node59596 = (inp[0]) ? node59606 : node59597;
														assign node59597 = (inp[3]) ? 4'b0000 : node59598;
															assign node59598 = (inp[5]) ? node59602 : node59599;
																assign node59599 = (inp[15]) ? 4'b0000 : 4'b0010;
																assign node59602 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node59606 = (inp[15]) ? node59610 : node59607;
															assign node59607 = (inp[3]) ? 4'b0010 : 4'b0000;
															assign node59610 = (inp[5]) ? 4'b0000 : node59611;
																assign node59611 = (inp[3]) ? 4'b0000 : 4'b0010;
											assign node59615 = (inp[3]) ? node59655 : node59616;
												assign node59616 = (inp[4]) ? node59636 : node59617;
													assign node59617 = (inp[9]) ? node59625 : node59618;
														assign node59618 = (inp[0]) ? node59622 : node59619;
															assign node59619 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node59622 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node59625 = (inp[0]) ? node59631 : node59626;
															assign node59626 = (inp[15]) ? node59628 : 4'b0100;
																assign node59628 = (inp[5]) ? 4'b0110 : 4'b0100;
															assign node59631 = (inp[15]) ? node59633 : 4'b0110;
																assign node59633 = (inp[5]) ? 4'b0100 : 4'b0110;
													assign node59636 = (inp[9]) ? node59646 : node59637;
														assign node59637 = (inp[0]) ? 4'b0100 : node59638;
															assign node59638 = (inp[5]) ? node59642 : node59639;
																assign node59639 = (inp[15]) ? 4'b0100 : 4'b0110;
																assign node59642 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node59646 = (inp[5]) ? 4'b0000 : node59647;
															assign node59647 = (inp[15]) ? node59651 : node59648;
																assign node59648 = (inp[0]) ? 4'b0000 : 4'b0010;
																assign node59651 = (inp[0]) ? 4'b0010 : 4'b0000;
												assign node59655 = (inp[15]) ? node59673 : node59656;
													assign node59656 = (inp[0]) ? node59666 : node59657;
														assign node59657 = (inp[4]) ? node59663 : node59658;
															assign node59658 = (inp[9]) ? 4'b0100 : node59659;
																assign node59659 = (inp[5]) ? 4'b0000 : 4'b0010;
															assign node59663 = (inp[9]) ? 4'b0000 : 4'b0100;
														assign node59666 = (inp[4]) ? node59670 : node59667;
															assign node59667 = (inp[9]) ? 4'b0110 : 4'b0010;
															assign node59670 = (inp[9]) ? 4'b0010 : 4'b0110;
													assign node59673 = (inp[0]) ? node59683 : node59674;
														assign node59674 = (inp[5]) ? node59676 : 4'b0110;
															assign node59676 = (inp[9]) ? node59680 : node59677;
																assign node59677 = (inp[4]) ? 4'b0110 : 4'b0010;
																assign node59680 = (inp[4]) ? 4'b0010 : 4'b0110;
														assign node59683 = (inp[4]) ? 4'b0100 : node59684;
															assign node59684 = (inp[9]) ? 4'b0100 : 4'b0000;
						assign node59688 = (inp[9]) ? node60554 : node59689;
							assign node59689 = (inp[4]) ? node60053 : node59690;
								assign node59690 = (inp[7]) ? node59906 : node59691;
									assign node59691 = (inp[8]) ? node59797 : node59692;
										assign node59692 = (inp[14]) ? node59736 : node59693;
											assign node59693 = (inp[2]) ? node59719 : node59694;
												assign node59694 = (inp[12]) ? node59704 : node59695;
													assign node59695 = (inp[15]) ? node59697 : 4'b0001;
														assign node59697 = (inp[0]) ? node59699 : 4'b0001;
															assign node59699 = (inp[3]) ? node59701 : 4'b0011;
																assign node59701 = (inp[5]) ? 4'b0001 : 4'b0011;
													assign node59704 = (inp[0]) ? node59712 : node59705;
														assign node59705 = (inp[15]) ? 4'b0001 : node59706;
															assign node59706 = (inp[3]) ? node59708 : 4'b0011;
																assign node59708 = (inp[5]) ? 4'b0001 : 4'b0011;
														assign node59712 = (inp[15]) ? 4'b0011 : node59713;
															assign node59713 = (inp[3]) ? node59715 : 4'b0001;
																assign node59715 = (inp[5]) ? 4'b0011 : 4'b0001;
												assign node59719 = (inp[5]) ? node59727 : node59720;
													assign node59720 = (inp[15]) ? node59724 : node59721;
														assign node59721 = (inp[0]) ? 4'b0000 : 4'b0010;
														assign node59724 = (inp[0]) ? 4'b0010 : 4'b0000;
													assign node59727 = (inp[0]) ? node59729 : 4'b0000;
														assign node59729 = (inp[12]) ? 4'b0000 : node59730;
															assign node59730 = (inp[3]) ? node59732 : 4'b0010;
																assign node59732 = (inp[15]) ? 4'b0000 : 4'b0010;
											assign node59736 = (inp[2]) ? node59770 : node59737;
												assign node59737 = (inp[12]) ? node59753 : node59738;
													assign node59738 = (inp[15]) ? node59746 : node59739;
														assign node59739 = (inp[0]) ? node59741 : 4'b0010;
															assign node59741 = (inp[5]) ? node59743 : 4'b0000;
																assign node59743 = (inp[3]) ? 4'b0010 : 4'b0000;
														assign node59746 = (inp[0]) ? node59750 : node59747;
															assign node59747 = (inp[3]) ? 4'b0010 : 4'b0000;
															assign node59750 = (inp[3]) ? 4'b0000 : 4'b0010;
													assign node59753 = (inp[5]) ? node59763 : node59754;
														assign node59754 = (inp[3]) ? 4'b0010 : node59755;
															assign node59755 = (inp[15]) ? node59759 : node59756;
																assign node59756 = (inp[0]) ? 4'b0000 : 4'b0010;
																assign node59759 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node59763 = (inp[0]) ? node59765 : 4'b0010;
															assign node59765 = (inp[3]) ? node59767 : 4'b0010;
																assign node59767 = (inp[15]) ? 4'b0000 : 4'b0010;
												assign node59770 = (inp[12]) ? node59788 : node59771;
													assign node59771 = (inp[0]) ? node59781 : node59772;
														assign node59772 = (inp[15]) ? node59778 : node59773;
															assign node59773 = (inp[5]) ? node59775 : 4'b0010;
																assign node59775 = (inp[3]) ? 4'b0000 : 4'b0010;
															assign node59778 = (inp[5]) ? 4'b0010 : 4'b0000;
														assign node59781 = (inp[15]) ? node59785 : node59782;
															assign node59782 = (inp[3]) ? 4'b0010 : 4'b0000;
															assign node59785 = (inp[3]) ? 4'b0000 : 4'b0010;
													assign node59788 = (inp[5]) ? node59790 : 4'b0000;
														assign node59790 = (inp[3]) ? node59792 : 4'b0010;
															assign node59792 = (inp[0]) ? 4'b0000 : node59793;
																assign node59793 = (inp[15]) ? 4'b0010 : 4'b0000;
										assign node59797 = (inp[2]) ? node59853 : node59798;
											assign node59798 = (inp[14]) ? node59830 : node59799;
												assign node59799 = (inp[12]) ? node59809 : node59800;
													assign node59800 = (inp[15]) ? node59804 : node59801;
														assign node59801 = (inp[0]) ? 4'b0000 : 4'b0010;
														assign node59804 = (inp[0]) ? 4'b0010 : node59805;
															assign node59805 = (inp[3]) ? 4'b0010 : 4'b0000;
													assign node59809 = (inp[15]) ? node59821 : node59810;
														assign node59810 = (inp[0]) ? node59816 : node59811;
															assign node59811 = (inp[3]) ? node59813 : 4'b0010;
																assign node59813 = (inp[5]) ? 4'b0000 : 4'b0010;
															assign node59816 = (inp[3]) ? node59818 : 4'b0000;
																assign node59818 = (inp[5]) ? 4'b0010 : 4'b0000;
														assign node59821 = (inp[0]) ? node59827 : node59822;
															assign node59822 = (inp[3]) ? node59824 : 4'b0000;
																assign node59824 = (inp[5]) ? 4'b0010 : 4'b0000;
															assign node59827 = (inp[5]) ? 4'b0000 : 4'b0010;
												assign node59830 = (inp[15]) ? node59842 : node59831;
													assign node59831 = (inp[0]) ? node59837 : node59832;
														assign node59832 = (inp[3]) ? node59834 : 4'b0011;
															assign node59834 = (inp[5]) ? 4'b0001 : 4'b0011;
														assign node59837 = (inp[3]) ? node59839 : 4'b0001;
															assign node59839 = (inp[5]) ? 4'b0011 : 4'b0001;
													assign node59842 = (inp[0]) ? node59848 : node59843;
														assign node59843 = (inp[3]) ? node59845 : 4'b0001;
															assign node59845 = (inp[5]) ? 4'b0011 : 4'b0001;
														assign node59848 = (inp[5]) ? node59850 : 4'b0011;
															assign node59850 = (inp[3]) ? 4'b0001 : 4'b0011;
											assign node59853 = (inp[14]) ? node59875 : node59854;
												assign node59854 = (inp[0]) ? node59864 : node59855;
													assign node59855 = (inp[15]) ? node59859 : node59856;
														assign node59856 = (inp[5]) ? 4'b0001 : 4'b0011;
														assign node59859 = (inp[5]) ? node59861 : 4'b0001;
															assign node59861 = (inp[3]) ? 4'b0011 : 4'b0001;
													assign node59864 = (inp[15]) ? node59870 : node59865;
														assign node59865 = (inp[3]) ? node59867 : 4'b0001;
															assign node59867 = (inp[5]) ? 4'b0011 : 4'b0001;
														assign node59870 = (inp[3]) ? node59872 : 4'b0011;
															assign node59872 = (inp[5]) ? 4'b0001 : 4'b0011;
												assign node59875 = (inp[3]) ? node59893 : node59876;
													assign node59876 = (inp[5]) ? node59884 : node59877;
														assign node59877 = (inp[0]) ? node59881 : node59878;
															assign node59878 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node59881 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node59884 = (inp[12]) ? 4'b0001 : node59885;
															assign node59885 = (inp[0]) ? node59889 : node59886;
																assign node59886 = (inp[15]) ? 4'b0001 : 4'b0011;
																assign node59889 = (inp[15]) ? 4'b0011 : 4'b0001;
													assign node59893 = (inp[15]) ? node59901 : node59894;
														assign node59894 = (inp[5]) ? node59898 : node59895;
															assign node59895 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node59898 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node59901 = (inp[5]) ? node59903 : 4'b0011;
															assign node59903 = (inp[0]) ? 4'b0001 : 4'b0011;
									assign node59906 = (inp[8]) ? node59972 : node59907;
										assign node59907 = (inp[14]) ? node59949 : node59908;
											assign node59908 = (inp[2]) ? node59934 : node59909;
												assign node59909 = (inp[3]) ? node59917 : node59910;
													assign node59910 = (inp[15]) ? node59914 : node59911;
														assign node59911 = (inp[0]) ? 4'b0000 : 4'b0010;
														assign node59914 = (inp[0]) ? 4'b0010 : 4'b0000;
													assign node59917 = (inp[0]) ? node59927 : node59918;
														assign node59918 = (inp[12]) ? node59924 : node59919;
															assign node59919 = (inp[15]) ? node59921 : 4'b0000;
																assign node59921 = (inp[5]) ? 4'b0010 : 4'b0000;
															assign node59924 = (inp[5]) ? 4'b0000 : 4'b0010;
														assign node59927 = (inp[15]) ? node59931 : node59928;
															assign node59928 = (inp[5]) ? 4'b0010 : 4'b0000;
															assign node59931 = (inp[5]) ? 4'b0000 : 4'b0010;
												assign node59934 = (inp[0]) ? node59944 : node59935;
													assign node59935 = (inp[15]) ? node59941 : node59936;
														assign node59936 = (inp[3]) ? node59938 : 4'b0011;
															assign node59938 = (inp[5]) ? 4'b0001 : 4'b0011;
														assign node59941 = (inp[5]) ? 4'b0011 : 4'b0001;
													assign node59944 = (inp[15]) ? 4'b0011 : node59945;
														assign node59945 = (inp[5]) ? 4'b0011 : 4'b0001;
											assign node59949 = (inp[0]) ? node59961 : node59950;
												assign node59950 = (inp[15]) ? node59956 : node59951;
													assign node59951 = (inp[5]) ? node59953 : 4'b0011;
														assign node59953 = (inp[3]) ? 4'b0001 : 4'b0011;
													assign node59956 = (inp[5]) ? node59958 : 4'b0001;
														assign node59958 = (inp[3]) ? 4'b0011 : 4'b0001;
												assign node59961 = (inp[15]) ? node59967 : node59962;
													assign node59962 = (inp[3]) ? node59964 : 4'b0001;
														assign node59964 = (inp[5]) ? 4'b0011 : 4'b0001;
													assign node59967 = (inp[5]) ? node59969 : 4'b0011;
														assign node59969 = (inp[3]) ? 4'b0001 : 4'b0011;
										assign node59972 = (inp[14]) ? node60030 : node59973;
											assign node59973 = (inp[2]) ? node59999 : node59974;
												assign node59974 = (inp[3]) ? node59982 : node59975;
													assign node59975 = (inp[0]) ? node59979 : node59976;
														assign node59976 = (inp[15]) ? 4'b0001 : 4'b0011;
														assign node59979 = (inp[15]) ? 4'b0011 : 4'b0001;
													assign node59982 = (inp[0]) ? node59990 : node59983;
														assign node59983 = (inp[5]) ? node59987 : node59984;
															assign node59984 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node59987 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node59990 = (inp[12]) ? 4'b0001 : node59991;
															assign node59991 = (inp[5]) ? node59995 : node59992;
																assign node59992 = (inp[15]) ? 4'b0011 : 4'b0001;
																assign node59995 = (inp[15]) ? 4'b0001 : 4'b0011;
												assign node59999 = (inp[3]) ? node60015 : node60000;
													assign node60000 = (inp[5]) ? node60010 : node60001;
														assign node60001 = (inp[12]) ? node60003 : 4'b0010;
															assign node60003 = (inp[0]) ? node60007 : node60004;
																assign node60004 = (inp[15]) ? 4'b0000 : 4'b0010;
																assign node60007 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node60010 = (inp[15]) ? node60012 : 4'b0000;
															assign node60012 = (inp[0]) ? 4'b0010 : 4'b0000;
													assign node60015 = (inp[5]) ? node60023 : node60016;
														assign node60016 = (inp[15]) ? node60020 : node60017;
															assign node60017 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node60020 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node60023 = (inp[12]) ? 4'b0010 : node60024;
															assign node60024 = (inp[0]) ? node60026 : 4'b0010;
																assign node60026 = (inp[15]) ? 4'b0000 : 4'b0010;
											assign node60030 = (inp[15]) ? node60042 : node60031;
												assign node60031 = (inp[0]) ? node60037 : node60032;
													assign node60032 = (inp[3]) ? node60034 : 4'b0010;
														assign node60034 = (inp[5]) ? 4'b0000 : 4'b0010;
													assign node60037 = (inp[3]) ? node60039 : 4'b0000;
														assign node60039 = (inp[5]) ? 4'b0010 : 4'b0000;
												assign node60042 = (inp[0]) ? node60048 : node60043;
													assign node60043 = (inp[3]) ? node60045 : 4'b0000;
														assign node60045 = (inp[5]) ? 4'b0010 : 4'b0000;
													assign node60048 = (inp[5]) ? node60050 : 4'b0010;
														assign node60050 = (inp[3]) ? 4'b0000 : 4'b0010;
								assign node60053 = (inp[5]) ? node60331 : node60054;
									assign node60054 = (inp[12]) ? node60200 : node60055;
										assign node60055 = (inp[15]) ? node60131 : node60056;
											assign node60056 = (inp[8]) ? node60094 : node60057;
												assign node60057 = (inp[7]) ? node60075 : node60058;
													assign node60058 = (inp[2]) ? node60068 : node60059;
														assign node60059 = (inp[14]) ? node60065 : node60060;
															assign node60060 = (inp[0]) ? 4'b0111 : node60061;
																assign node60061 = (inp[3]) ? 4'b0101 : 4'b0111;
															assign node60065 = (inp[0]) ? 4'b0100 : 4'b0110;
														assign node60068 = (inp[3]) ? node60072 : node60069;
															assign node60069 = (inp[0]) ? 4'b0100 : 4'b0110;
															assign node60072 = (inp[0]) ? 4'b0110 : 4'b0100;
													assign node60075 = (inp[14]) ? node60087 : node60076;
														assign node60076 = (inp[2]) ? node60082 : node60077;
															assign node60077 = (inp[3]) ? 4'b0110 : node60078;
																assign node60078 = (inp[0]) ? 4'b0100 : 4'b0110;
															assign node60082 = (inp[3]) ? node60084 : 4'b0111;
																assign node60084 = (inp[0]) ? 4'b0111 : 4'b0101;
														assign node60087 = (inp[0]) ? node60091 : node60088;
															assign node60088 = (inp[3]) ? 4'b0101 : 4'b0111;
															assign node60091 = (inp[3]) ? 4'b0111 : 4'b0101;
												assign node60094 = (inp[7]) ? node60110 : node60095;
													assign node60095 = (inp[14]) ? node60105 : node60096;
														assign node60096 = (inp[2]) ? node60102 : node60097;
															assign node60097 = (inp[0]) ? 4'b0100 : node60098;
																assign node60098 = (inp[3]) ? 4'b0100 : 4'b0110;
															assign node60102 = (inp[3]) ? 4'b0111 : 4'b0101;
														assign node60105 = (inp[0]) ? node60107 : 4'b0111;
															assign node60107 = (inp[3]) ? 4'b0111 : 4'b0101;
													assign node60110 = (inp[14]) ? node60124 : node60111;
														assign node60111 = (inp[2]) ? node60117 : node60112;
															assign node60112 = (inp[3]) ? 4'b0101 : node60113;
																assign node60113 = (inp[0]) ? 4'b0101 : 4'b0111;
															assign node60117 = (inp[3]) ? node60121 : node60118;
																assign node60118 = (inp[0]) ? 4'b0100 : 4'b0110;
																assign node60121 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node60124 = (inp[3]) ? node60128 : node60125;
															assign node60125 = (inp[0]) ? 4'b0100 : 4'b0110;
															assign node60128 = (inp[0]) ? 4'b0110 : 4'b0100;
											assign node60131 = (inp[14]) ? node60171 : node60132;
												assign node60132 = (inp[7]) ? node60150 : node60133;
													assign node60133 = (inp[3]) ? node60143 : node60134;
														assign node60134 = (inp[0]) ? node60140 : node60135;
															assign node60135 = (inp[2]) ? node60137 : 4'b0100;
																assign node60137 = (inp[8]) ? 4'b0101 : 4'b0100;
															assign node60140 = (inp[2]) ? 4'b0110 : 4'b0111;
														assign node60143 = (inp[0]) ? 4'b0101 : node60144;
															assign node60144 = (inp[2]) ? 4'b0111 : node60145;
																assign node60145 = (inp[8]) ? 4'b0110 : 4'b0111;
													assign node60150 = (inp[3]) ? node60164 : node60151;
														assign node60151 = (inp[0]) ? node60159 : node60152;
															assign node60152 = (inp[8]) ? node60156 : node60153;
																assign node60153 = (inp[2]) ? 4'b0101 : 4'b0100;
																assign node60156 = (inp[2]) ? 4'b0100 : 4'b0101;
															assign node60159 = (inp[8]) ? node60161 : 4'b0111;
																assign node60161 = (inp[2]) ? 4'b0110 : 4'b0111;
														assign node60164 = (inp[0]) ? node60166 : 4'b0110;
															assign node60166 = (inp[2]) ? node60168 : 4'b0100;
																assign node60168 = (inp[8]) ? 4'b0100 : 4'b0101;
												assign node60171 = (inp[7]) ? node60185 : node60172;
													assign node60172 = (inp[8]) ? node60178 : node60173;
														assign node60173 = (inp[3]) ? 4'b0100 : node60174;
															assign node60174 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node60178 = (inp[0]) ? node60182 : node60179;
															assign node60179 = (inp[3]) ? 4'b0111 : 4'b0101;
															assign node60182 = (inp[3]) ? 4'b0101 : 4'b0111;
													assign node60185 = (inp[8]) ? node60195 : node60186;
														assign node60186 = (inp[2]) ? 4'b0111 : node60187;
															assign node60187 = (inp[3]) ? node60191 : node60188;
																assign node60188 = (inp[0]) ? 4'b0111 : 4'b0101;
																assign node60191 = (inp[0]) ? 4'b0101 : 4'b0111;
														assign node60195 = (inp[3]) ? node60197 : 4'b0110;
															assign node60197 = (inp[0]) ? 4'b0100 : 4'b0110;
										assign node60200 = (inp[15]) ? node60258 : node60201;
											assign node60201 = (inp[0]) ? node60233 : node60202;
												assign node60202 = (inp[3]) ? node60214 : node60203;
													assign node60203 = (inp[2]) ? 4'b0111 : node60204;
														assign node60204 = (inp[7]) ? node60206 : 4'b0111;
															assign node60206 = (inp[14]) ? node60210 : node60207;
																assign node60207 = (inp[8]) ? 4'b0111 : 4'b0110;
																assign node60210 = (inp[8]) ? 4'b0110 : 4'b0111;
													assign node60214 = (inp[2]) ? node60228 : node60215;
														assign node60215 = (inp[7]) ? node60223 : node60216;
															assign node60216 = (inp[8]) ? node60220 : node60217;
																assign node60217 = (inp[14]) ? 4'b0100 : 4'b0101;
																assign node60220 = (inp[14]) ? 4'b0101 : 4'b0100;
															assign node60223 = (inp[14]) ? node60225 : 4'b0101;
																assign node60225 = (inp[8]) ? 4'b0100 : 4'b0101;
														assign node60228 = (inp[8]) ? 4'b0100 : node60229;
															assign node60229 = (inp[7]) ? 4'b0101 : 4'b0100;
												assign node60233 = (inp[3]) ? node60253 : node60234;
													assign node60234 = (inp[7]) ? node60242 : node60235;
														assign node60235 = (inp[8]) ? 4'b0101 : node60236;
															assign node60236 = (inp[14]) ? 4'b0100 : node60237;
																assign node60237 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node60242 = (inp[8]) ? node60248 : node60243;
															assign node60243 = (inp[14]) ? 4'b0101 : node60244;
																assign node60244 = (inp[2]) ? 4'b0101 : 4'b0100;
															assign node60248 = (inp[2]) ? 4'b0100 : node60249;
																assign node60249 = (inp[14]) ? 4'b0100 : 4'b0101;
													assign node60253 = (inp[8]) ? 4'b0111 : node60254;
														assign node60254 = (inp[7]) ? 4'b0111 : 4'b0110;
											assign node60258 = (inp[2]) ? node60286 : node60259;
												assign node60259 = (inp[0]) ? node60275 : node60260;
													assign node60260 = (inp[3]) ? node60272 : node60261;
														assign node60261 = (inp[7]) ? node60267 : node60262;
															assign node60262 = (inp[14]) ? node60264 : 4'b0100;
																assign node60264 = (inp[8]) ? 4'b0101 : 4'b0100;
															assign node60267 = (inp[8]) ? node60269 : 4'b0101;
																assign node60269 = (inp[14]) ? 4'b0100 : 4'b0101;
														assign node60272 = (inp[14]) ? 4'b0110 : 4'b0111;
													assign node60275 = (inp[3]) ? node60279 : node60276;
														assign node60276 = (inp[8]) ? 4'b0110 : 4'b0111;
														assign node60279 = (inp[8]) ? 4'b0101 : node60280;
															assign node60280 = (inp[14]) ? 4'b0101 : node60281;
																assign node60281 = (inp[7]) ? 4'b0100 : 4'b0101;
												assign node60286 = (inp[14]) ? node60308 : node60287;
													assign node60287 = (inp[8]) ? node60297 : node60288;
														assign node60288 = (inp[7]) ? 4'b0101 : node60289;
															assign node60289 = (inp[3]) ? node60293 : node60290;
																assign node60290 = (inp[0]) ? 4'b0110 : 4'b0100;
																assign node60293 = (inp[0]) ? 4'b0100 : 4'b0110;
														assign node60297 = (inp[7]) ? node60301 : node60298;
															assign node60298 = (inp[3]) ? 4'b0111 : 4'b0101;
															assign node60301 = (inp[0]) ? node60305 : node60302;
																assign node60302 = (inp[3]) ? 4'b0110 : 4'b0100;
																assign node60305 = (inp[3]) ? 4'b0100 : 4'b0110;
													assign node60308 = (inp[3]) ? node60322 : node60309;
														assign node60309 = (inp[0]) ? node60315 : node60310;
															assign node60310 = (inp[7]) ? node60312 : 4'b0101;
																assign node60312 = (inp[8]) ? 4'b0100 : 4'b0101;
															assign node60315 = (inp[8]) ? node60319 : node60316;
																assign node60316 = (inp[7]) ? 4'b0111 : 4'b0110;
																assign node60319 = (inp[7]) ? 4'b0110 : 4'b0111;
														assign node60322 = (inp[0]) ? 4'b0100 : node60323;
															assign node60323 = (inp[8]) ? node60327 : node60324;
																assign node60324 = (inp[7]) ? 4'b0111 : 4'b0110;
																assign node60327 = (inp[7]) ? 4'b0110 : 4'b0111;
									assign node60331 = (inp[14]) ? node60479 : node60332;
										assign node60332 = (inp[3]) ? node60404 : node60333;
											assign node60333 = (inp[0]) ? node60373 : node60334;
												assign node60334 = (inp[15]) ? node60352 : node60335;
													assign node60335 = (inp[2]) ? node60343 : node60336;
														assign node60336 = (inp[8]) ? node60340 : node60337;
															assign node60337 = (inp[7]) ? 4'b0100 : 4'b0101;
															assign node60340 = (inp[7]) ? 4'b0101 : 4'b0100;
														assign node60343 = (inp[12]) ? 4'b0101 : node60344;
															assign node60344 = (inp[8]) ? node60348 : node60345;
																assign node60345 = (inp[7]) ? 4'b0101 : 4'b0100;
																assign node60348 = (inp[7]) ? 4'b0100 : 4'b0101;
													assign node60352 = (inp[12]) ? node60360 : node60353;
														assign node60353 = (inp[7]) ? node60355 : 4'b0111;
															assign node60355 = (inp[2]) ? node60357 : 4'b0111;
																assign node60357 = (inp[8]) ? 4'b0110 : 4'b0111;
														assign node60360 = (inp[2]) ? node60366 : node60361;
															assign node60361 = (inp[8]) ? node60363 : 4'b0110;
																assign node60363 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node60366 = (inp[8]) ? node60370 : node60367;
																assign node60367 = (inp[7]) ? 4'b0111 : 4'b0110;
																assign node60370 = (inp[7]) ? 4'b0110 : 4'b0111;
												assign node60373 = (inp[15]) ? node60395 : node60374;
													assign node60374 = (inp[7]) ? node60388 : node60375;
														assign node60375 = (inp[12]) ? node60381 : node60376;
															assign node60376 = (inp[2]) ? node60378 : 4'b0111;
																assign node60378 = (inp[8]) ? 4'b0111 : 4'b0110;
															assign node60381 = (inp[8]) ? node60385 : node60382;
																assign node60382 = (inp[2]) ? 4'b0110 : 4'b0111;
																assign node60385 = (inp[2]) ? 4'b0111 : 4'b0110;
														assign node60388 = (inp[12]) ? 4'b0111 : node60389;
															assign node60389 = (inp[2]) ? node60391 : 4'b0111;
																assign node60391 = (inp[8]) ? 4'b0110 : 4'b0111;
													assign node60395 = (inp[7]) ? 4'b0101 : node60396;
														assign node60396 = (inp[12]) ? node60398 : 4'b0101;
															assign node60398 = (inp[2]) ? 4'b0100 : node60399;
																assign node60399 = (inp[8]) ? 4'b0100 : 4'b0101;
											assign node60404 = (inp[12]) ? node60440 : node60405;
												assign node60405 = (inp[8]) ? node60421 : node60406;
													assign node60406 = (inp[0]) ? node60418 : node60407;
														assign node60407 = (inp[15]) ? node60413 : node60408;
															assign node60408 = (inp[2]) ? 4'b0101 : node60409;
																assign node60409 = (inp[7]) ? 4'b0100 : 4'b0101;
															assign node60413 = (inp[7]) ? 4'b0110 : node60414;
																assign node60414 = (inp[2]) ? 4'b0110 : 4'b0111;
														assign node60418 = (inp[15]) ? 4'b0100 : 4'b0110;
													assign node60421 = (inp[15]) ? node60429 : node60422;
														assign node60422 = (inp[7]) ? node60426 : node60423;
															assign node60423 = (inp[2]) ? 4'b0111 : 4'b0110;
															assign node60426 = (inp[2]) ? 4'b0110 : 4'b0111;
														assign node60429 = (inp[0]) ? node60437 : node60430;
															assign node60430 = (inp[7]) ? node60434 : node60431;
																assign node60431 = (inp[2]) ? 4'b0111 : 4'b0110;
																assign node60434 = (inp[2]) ? 4'b0110 : 4'b0111;
															assign node60437 = (inp[2]) ? 4'b0100 : 4'b0101;
												assign node60440 = (inp[7]) ? node60458 : node60441;
													assign node60441 = (inp[15]) ? node60449 : node60442;
														assign node60442 = (inp[0]) ? node60444 : 4'b0101;
															assign node60444 = (inp[2]) ? node60446 : 4'b0111;
																assign node60446 = (inp[8]) ? 4'b0111 : 4'b0110;
														assign node60449 = (inp[0]) ? node60453 : node60450;
															assign node60450 = (inp[2]) ? 4'b0111 : 4'b0110;
															assign node60453 = (inp[8]) ? node60455 : 4'b0101;
																assign node60455 = (inp[2]) ? 4'b0101 : 4'b0100;
													assign node60458 = (inp[0]) ? node60470 : node60459;
														assign node60459 = (inp[15]) ? node60465 : node60460;
															assign node60460 = (inp[8]) ? node60462 : 4'b0101;
																assign node60462 = (inp[2]) ? 4'b0100 : 4'b0101;
															assign node60465 = (inp[2]) ? node60467 : 4'b0111;
																assign node60467 = (inp[8]) ? 4'b0110 : 4'b0111;
														assign node60470 = (inp[15]) ? node60472 : 4'b0110;
															assign node60472 = (inp[2]) ? node60476 : node60473;
																assign node60473 = (inp[8]) ? 4'b0101 : 4'b0100;
																assign node60476 = (inp[8]) ? 4'b0100 : 4'b0101;
										assign node60479 = (inp[0]) ? node60521 : node60480;
											assign node60480 = (inp[15]) ? node60488 : node60481;
												assign node60481 = (inp[7]) ? node60485 : node60482;
													assign node60482 = (inp[8]) ? 4'b0101 : 4'b0100;
													assign node60485 = (inp[8]) ? 4'b0100 : 4'b0101;
												assign node60488 = (inp[12]) ? node60514 : node60489;
													assign node60489 = (inp[3]) ? node60501 : node60490;
														assign node60490 = (inp[2]) ? node60496 : node60491;
															assign node60491 = (inp[8]) ? 4'b0110 : node60492;
																assign node60492 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node60496 = (inp[8]) ? node60498 : 4'b0110;
																assign node60498 = (inp[7]) ? 4'b0110 : 4'b0111;
														assign node60501 = (inp[2]) ? node60509 : node60502;
															assign node60502 = (inp[8]) ? node60506 : node60503;
																assign node60503 = (inp[7]) ? 4'b0111 : 4'b0110;
																assign node60506 = (inp[7]) ? 4'b0110 : 4'b0111;
															assign node60509 = (inp[8]) ? node60511 : 4'b0110;
																assign node60511 = (inp[7]) ? 4'b0110 : 4'b0111;
													assign node60514 = (inp[7]) ? node60518 : node60515;
														assign node60515 = (inp[8]) ? 4'b0111 : 4'b0110;
														assign node60518 = (inp[8]) ? 4'b0110 : 4'b0111;
											assign node60521 = (inp[15]) ? node60547 : node60522;
												assign node60522 = (inp[12]) ? node60530 : node60523;
													assign node60523 = (inp[8]) ? node60527 : node60524;
														assign node60524 = (inp[7]) ? 4'b0111 : 4'b0110;
														assign node60527 = (inp[7]) ? 4'b0110 : 4'b0111;
													assign node60530 = (inp[3]) ? node60540 : node60531;
														assign node60531 = (inp[2]) ? node60533 : 4'b0110;
															assign node60533 = (inp[7]) ? node60537 : node60534;
																assign node60534 = (inp[8]) ? 4'b0111 : 4'b0110;
																assign node60537 = (inp[8]) ? 4'b0110 : 4'b0111;
														assign node60540 = (inp[2]) ? node60542 : 4'b0111;
															assign node60542 = (inp[8]) ? node60544 : 4'b0110;
																assign node60544 = (inp[7]) ? 4'b0110 : 4'b0111;
												assign node60547 = (inp[8]) ? node60551 : node60548;
													assign node60548 = (inp[7]) ? 4'b0101 : 4'b0100;
													assign node60551 = (inp[7]) ? 4'b0100 : 4'b0101;
							assign node60554 = (inp[4]) ? node60952 : node60555;
								assign node60555 = (inp[7]) ? node60761 : node60556;
									assign node60556 = (inp[8]) ? node60668 : node60557;
										assign node60557 = (inp[2]) ? node60609 : node60558;
											assign node60558 = (inp[14]) ? node60584 : node60559;
												assign node60559 = (inp[15]) ? node60571 : node60560;
													assign node60560 = (inp[0]) ? node60566 : node60561;
														assign node60561 = (inp[3]) ? 4'b0101 : node60562;
															assign node60562 = (inp[5]) ? 4'b0101 : 4'b0111;
														assign node60566 = (inp[5]) ? 4'b0111 : node60567;
															assign node60567 = (inp[3]) ? 4'b0111 : 4'b0101;
													assign node60571 = (inp[3]) ? 4'b0101 : node60572;
														assign node60572 = (inp[12]) ? node60578 : node60573;
															assign node60573 = (inp[5]) ? 4'b0111 : node60574;
																assign node60574 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node60578 = (inp[0]) ? node60580 : 4'b0101;
																assign node60580 = (inp[5]) ? 4'b0101 : 4'b0111;
												assign node60584 = (inp[0]) ? node60594 : node60585;
													assign node60585 = (inp[15]) ? node60589 : node60586;
														assign node60586 = (inp[5]) ? 4'b0100 : 4'b0110;
														assign node60589 = (inp[5]) ? 4'b0110 : node60590;
															assign node60590 = (inp[3]) ? 4'b0110 : 4'b0100;
													assign node60594 = (inp[3]) ? 4'b0100 : node60595;
														assign node60595 = (inp[12]) ? node60601 : node60596;
															assign node60596 = (inp[5]) ? 4'b0100 : node60597;
																assign node60597 = (inp[15]) ? 4'b0110 : 4'b0100;
															assign node60601 = (inp[15]) ? node60605 : node60602;
																assign node60602 = (inp[5]) ? 4'b0110 : 4'b0100;
																assign node60605 = (inp[5]) ? 4'b0100 : 4'b0110;
											assign node60609 = (inp[3]) ? node60651 : node60610;
												assign node60610 = (inp[12]) ? node60630 : node60611;
													assign node60611 = (inp[14]) ? node60625 : node60612;
														assign node60612 = (inp[15]) ? node60620 : node60613;
															assign node60613 = (inp[0]) ? node60617 : node60614;
																assign node60614 = (inp[5]) ? 4'b0100 : 4'b0110;
																assign node60617 = (inp[5]) ? 4'b0110 : 4'b0100;
															assign node60620 = (inp[0]) ? node60622 : 4'b0100;
																assign node60622 = (inp[5]) ? 4'b0100 : 4'b0110;
														assign node60625 = (inp[0]) ? 4'b0110 : node60626;
															assign node60626 = (inp[5]) ? 4'b0110 : 4'b0100;
													assign node60630 = (inp[5]) ? node60644 : node60631;
														assign node60631 = (inp[14]) ? node60637 : node60632;
															assign node60632 = (inp[15]) ? 4'b0100 : node60633;
																assign node60633 = (inp[0]) ? 4'b0100 : 4'b0110;
															assign node60637 = (inp[15]) ? node60641 : node60638;
																assign node60638 = (inp[0]) ? 4'b0100 : 4'b0110;
																assign node60641 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node60644 = (inp[14]) ? 4'b0100 : node60645;
															assign node60645 = (inp[15]) ? node60647 : 4'b0100;
																assign node60647 = (inp[0]) ? 4'b0100 : 4'b0110;
												assign node60651 = (inp[5]) ? node60659 : node60652;
													assign node60652 = (inp[0]) ? node60656 : node60653;
														assign node60653 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node60656 = (inp[15]) ? 4'b0100 : 4'b0110;
													assign node60659 = (inp[14]) ? node60661 : 4'b0110;
														assign node60661 = (inp[15]) ? node60665 : node60662;
															assign node60662 = (inp[0]) ? 4'b0110 : 4'b0100;
															assign node60665 = (inp[0]) ? 4'b0100 : 4'b0110;
										assign node60668 = (inp[14]) ? node60706 : node60669;
											assign node60669 = (inp[2]) ? node60687 : node60670;
												assign node60670 = (inp[15]) ? node60678 : node60671;
													assign node60671 = (inp[0]) ? node60673 : 4'b0100;
														assign node60673 = (inp[3]) ? 4'b0110 : node60674;
															assign node60674 = (inp[5]) ? 4'b0110 : 4'b0100;
													assign node60678 = (inp[0]) ? node60680 : 4'b0110;
														assign node60680 = (inp[12]) ? 4'b0100 : node60681;
															assign node60681 = (inp[3]) ? 4'b0100 : node60682;
																assign node60682 = (inp[5]) ? 4'b0100 : 4'b0110;
												assign node60687 = (inp[0]) ? node60699 : node60688;
													assign node60688 = (inp[15]) ? node60694 : node60689;
														assign node60689 = (inp[3]) ? 4'b0101 : node60690;
															assign node60690 = (inp[5]) ? 4'b0101 : 4'b0111;
														assign node60694 = (inp[5]) ? 4'b0111 : node60695;
															assign node60695 = (inp[3]) ? 4'b0111 : 4'b0101;
													assign node60699 = (inp[15]) ? 4'b0101 : node60700;
														assign node60700 = (inp[3]) ? 4'b0111 : node60701;
															assign node60701 = (inp[5]) ? 4'b0111 : 4'b0101;
											assign node60706 = (inp[3]) ? node60740 : node60707;
												assign node60707 = (inp[15]) ? node60733 : node60708;
													assign node60708 = (inp[12]) ? node60720 : node60709;
														assign node60709 = (inp[2]) ? node60715 : node60710;
															assign node60710 = (inp[5]) ? node60712 : 4'b0101;
																assign node60712 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node60715 = (inp[5]) ? 4'b0101 : node60716;
																assign node60716 = (inp[0]) ? 4'b0101 : 4'b0111;
														assign node60720 = (inp[2]) ? node60728 : node60721;
															assign node60721 = (inp[0]) ? node60725 : node60722;
																assign node60722 = (inp[5]) ? 4'b0101 : 4'b0111;
																assign node60725 = (inp[5]) ? 4'b0111 : 4'b0101;
															assign node60728 = (inp[5]) ? node60730 : 4'b0111;
																assign node60730 = (inp[0]) ? 4'b0111 : 4'b0101;
													assign node60733 = (inp[0]) ? node60737 : node60734;
														assign node60734 = (inp[5]) ? 4'b0111 : 4'b0101;
														assign node60737 = (inp[5]) ? 4'b0101 : 4'b0111;
												assign node60740 = (inp[5]) ? node60748 : node60741;
													assign node60741 = (inp[15]) ? node60745 : node60742;
														assign node60742 = (inp[0]) ? 4'b0111 : 4'b0101;
														assign node60745 = (inp[0]) ? 4'b0101 : 4'b0111;
													assign node60748 = (inp[2]) ? node60754 : node60749;
														assign node60749 = (inp[0]) ? 4'b0101 : node60750;
															assign node60750 = (inp[15]) ? 4'b0111 : 4'b0101;
														assign node60754 = (inp[0]) ? node60758 : node60755;
															assign node60755 = (inp[15]) ? 4'b0111 : 4'b0101;
															assign node60758 = (inp[15]) ? 4'b0101 : 4'b0111;
									assign node60761 = (inp[8]) ? node60837 : node60762;
										assign node60762 = (inp[2]) ? node60814 : node60763;
											assign node60763 = (inp[14]) ? node60793 : node60764;
												assign node60764 = (inp[12]) ? node60780 : node60765;
													assign node60765 = (inp[3]) ? 4'b0110 : node60766;
														assign node60766 = (inp[15]) ? node60774 : node60767;
															assign node60767 = (inp[5]) ? node60771 : node60768;
																assign node60768 = (inp[0]) ? 4'b0100 : 4'b0110;
																assign node60771 = (inp[0]) ? 4'b0110 : 4'b0100;
															assign node60774 = (inp[0]) ? node60776 : 4'b0110;
																assign node60776 = (inp[5]) ? 4'b0100 : 4'b0110;
													assign node60780 = (inp[0]) ? node60782 : 4'b0100;
														assign node60782 = (inp[15]) ? node60788 : node60783;
															assign node60783 = (inp[3]) ? 4'b0110 : node60784;
																assign node60784 = (inp[5]) ? 4'b0110 : 4'b0100;
															assign node60788 = (inp[3]) ? 4'b0100 : node60789;
																assign node60789 = (inp[5]) ? 4'b0100 : 4'b0110;
												assign node60793 = (inp[5]) ? node60807 : node60794;
													assign node60794 = (inp[3]) ? node60802 : node60795;
														assign node60795 = (inp[15]) ? node60799 : node60796;
															assign node60796 = (inp[0]) ? 4'b0101 : 4'b0111;
															assign node60799 = (inp[0]) ? 4'b0111 : 4'b0101;
														assign node60802 = (inp[0]) ? 4'b0101 : node60803;
															assign node60803 = (inp[15]) ? 4'b0111 : 4'b0101;
													assign node60807 = (inp[15]) ? node60811 : node60808;
														assign node60808 = (inp[0]) ? 4'b0111 : 4'b0101;
														assign node60811 = (inp[0]) ? 4'b0101 : 4'b0111;
											assign node60814 = (inp[15]) ? node60826 : node60815;
												assign node60815 = (inp[0]) ? node60821 : node60816;
													assign node60816 = (inp[5]) ? 4'b0101 : node60817;
														assign node60817 = (inp[14]) ? 4'b0111 : 4'b0101;
													assign node60821 = (inp[5]) ? 4'b0111 : node60822;
														assign node60822 = (inp[3]) ? 4'b0111 : 4'b0101;
												assign node60826 = (inp[0]) ? node60832 : node60827;
													assign node60827 = (inp[5]) ? 4'b0111 : node60828;
														assign node60828 = (inp[3]) ? 4'b0111 : 4'b0101;
													assign node60832 = (inp[5]) ? 4'b0101 : node60833;
														assign node60833 = (inp[3]) ? 4'b0101 : 4'b0111;
										assign node60837 = (inp[14]) ? node60897 : node60838;
											assign node60838 = (inp[2]) ? node60858 : node60839;
												assign node60839 = (inp[0]) ? node60851 : node60840;
													assign node60840 = (inp[15]) ? node60846 : node60841;
														assign node60841 = (inp[3]) ? 4'b0101 : node60842;
															assign node60842 = (inp[12]) ? 4'b0101 : 4'b0111;
														assign node60846 = (inp[5]) ? 4'b0111 : node60847;
															assign node60847 = (inp[3]) ? 4'b0111 : 4'b0101;
													assign node60851 = (inp[15]) ? node60853 : 4'b0111;
														assign node60853 = (inp[5]) ? 4'b0101 : node60854;
															assign node60854 = (inp[3]) ? 4'b0101 : 4'b0111;
												assign node60858 = (inp[12]) ? node60880 : node60859;
													assign node60859 = (inp[5]) ? node60869 : node60860;
														assign node60860 = (inp[3]) ? node60862 : 4'b0110;
															assign node60862 = (inp[0]) ? node60866 : node60863;
																assign node60863 = (inp[15]) ? 4'b0110 : 4'b0100;
																assign node60866 = (inp[15]) ? 4'b0100 : 4'b0110;
														assign node60869 = (inp[3]) ? node60875 : node60870;
															assign node60870 = (inp[15]) ? 4'b0100 : node60871;
																assign node60871 = (inp[0]) ? 4'b0110 : 4'b0100;
															assign node60875 = (inp[15]) ? 4'b0110 : node60876;
																assign node60876 = (inp[0]) ? 4'b0110 : 4'b0100;
													assign node60880 = (inp[3]) ? node60890 : node60881;
														assign node60881 = (inp[5]) ? 4'b0110 : node60882;
															assign node60882 = (inp[0]) ? node60886 : node60883;
																assign node60883 = (inp[15]) ? 4'b0100 : 4'b0110;
																assign node60886 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node60890 = (inp[5]) ? 4'b0100 : node60891;
															assign node60891 = (inp[0]) ? 4'b0100 : node60892;
																assign node60892 = (inp[15]) ? 4'b0110 : 4'b0100;
											assign node60897 = (inp[12]) ? node60919 : node60898;
												assign node60898 = (inp[15]) ? node60910 : node60899;
													assign node60899 = (inp[0]) ? node60905 : node60900;
														assign node60900 = (inp[5]) ? 4'b0100 : node60901;
															assign node60901 = (inp[3]) ? 4'b0100 : 4'b0110;
														assign node60905 = (inp[3]) ? 4'b0110 : node60906;
															assign node60906 = (inp[5]) ? 4'b0110 : 4'b0100;
													assign node60910 = (inp[0]) ? node60914 : node60911;
														assign node60911 = (inp[3]) ? 4'b0110 : 4'b0100;
														assign node60914 = (inp[5]) ? 4'b0100 : node60915;
															assign node60915 = (inp[3]) ? 4'b0100 : 4'b0110;
												assign node60919 = (inp[2]) ? node60935 : node60920;
													assign node60920 = (inp[15]) ? node60928 : node60921;
														assign node60921 = (inp[0]) ? node60923 : 4'b0100;
															assign node60923 = (inp[5]) ? 4'b0110 : node60924;
																assign node60924 = (inp[3]) ? 4'b0110 : 4'b0100;
														assign node60928 = (inp[0]) ? node60930 : 4'b0110;
															assign node60930 = (inp[5]) ? 4'b0100 : node60931;
																assign node60931 = (inp[3]) ? 4'b0100 : 4'b0110;
													assign node60935 = (inp[0]) ? node60947 : node60936;
														assign node60936 = (inp[15]) ? node60942 : node60937;
															assign node60937 = (inp[5]) ? 4'b0100 : node60938;
																assign node60938 = (inp[3]) ? 4'b0100 : 4'b0110;
															assign node60942 = (inp[3]) ? 4'b0110 : node60943;
																assign node60943 = (inp[5]) ? 4'b0110 : 4'b0100;
														assign node60947 = (inp[15]) ? node60949 : 4'b0110;
															assign node60949 = (inp[5]) ? 4'b0100 : 4'b0110;
								assign node60952 = (inp[5]) ? node61202 : node60953;
									assign node60953 = (inp[8]) ? node61077 : node60954;
										assign node60954 = (inp[7]) ? node61022 : node60955;
											assign node60955 = (inp[2]) ? node60993 : node60956;
												assign node60956 = (inp[14]) ? node60976 : node60957;
													assign node60957 = (inp[12]) ? node60969 : node60958;
														assign node60958 = (inp[15]) ? node60964 : node60959;
															assign node60959 = (inp[3]) ? node60961 : 4'b0001;
																assign node60961 = (inp[0]) ? 4'b0011 : 4'b0001;
															assign node60964 = (inp[3]) ? node60966 : 4'b0011;
																assign node60966 = (inp[0]) ? 4'b0001 : 4'b0011;
														assign node60969 = (inp[3]) ? node60971 : 4'b0001;
															assign node60971 = (inp[15]) ? node60973 : 4'b0001;
																assign node60973 = (inp[0]) ? 4'b0001 : 4'b0011;
													assign node60976 = (inp[15]) ? node60986 : node60977;
														assign node60977 = (inp[12]) ? node60979 : 4'b0010;
															assign node60979 = (inp[0]) ? node60983 : node60980;
																assign node60980 = (inp[3]) ? 4'b0000 : 4'b0010;
																assign node60983 = (inp[3]) ? 4'b0010 : 4'b0000;
														assign node60986 = (inp[3]) ? node60990 : node60987;
															assign node60987 = (inp[0]) ? 4'b0010 : 4'b0000;
															assign node60990 = (inp[0]) ? 4'b0000 : 4'b0010;
												assign node60993 = (inp[12]) ? node61009 : node60994;
													assign node60994 = (inp[3]) ? node61004 : node60995;
														assign node60995 = (inp[14]) ? node60999 : node60996;
															assign node60996 = (inp[15]) ? 4'b0010 : 4'b0000;
															assign node60999 = (inp[15]) ? 4'b0000 : node61000;
																assign node61000 = (inp[0]) ? 4'b0000 : 4'b0010;
														assign node61004 = (inp[0]) ? node61006 : 4'b0000;
															assign node61006 = (inp[15]) ? 4'b0000 : 4'b0010;
													assign node61009 = (inp[0]) ? node61017 : node61010;
														assign node61010 = (inp[15]) ? node61014 : node61011;
															assign node61011 = (inp[3]) ? 4'b0000 : 4'b0010;
															assign node61014 = (inp[3]) ? 4'b0010 : 4'b0000;
														assign node61017 = (inp[3]) ? node61019 : 4'b0010;
															assign node61019 = (inp[15]) ? 4'b0000 : 4'b0010;
											assign node61022 = (inp[14]) ? node61052 : node61023;
												assign node61023 = (inp[2]) ? node61037 : node61024;
													assign node61024 = (inp[12]) ? node61030 : node61025;
														assign node61025 = (inp[0]) ? 4'b0010 : node61026;
															assign node61026 = (inp[3]) ? 4'b0000 : 4'b0010;
														assign node61030 = (inp[3]) ? 4'b0000 : node61031;
															assign node61031 = (inp[0]) ? 4'b0000 : node61032;
																assign node61032 = (inp[15]) ? 4'b0000 : 4'b0010;
													assign node61037 = (inp[12]) ? node61043 : node61038;
														assign node61038 = (inp[15]) ? 4'b0001 : node61039;
															assign node61039 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node61043 = (inp[0]) ? 4'b0011 : node61044;
															assign node61044 = (inp[15]) ? node61048 : node61045;
																assign node61045 = (inp[3]) ? 4'b0001 : 4'b0011;
																assign node61048 = (inp[3]) ? 4'b0011 : 4'b0001;
												assign node61052 = (inp[2]) ? node61068 : node61053;
													assign node61053 = (inp[3]) ? node61059 : node61054;
														assign node61054 = (inp[15]) ? node61056 : 4'b0001;
															assign node61056 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node61059 = (inp[12]) ? node61063 : node61060;
															assign node61060 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node61063 = (inp[0]) ? node61065 : 4'b0001;
																assign node61065 = (inp[15]) ? 4'b0001 : 4'b0011;
													assign node61068 = (inp[12]) ? 4'b0001 : node61069;
														assign node61069 = (inp[15]) ? node61071 : 4'b0001;
															assign node61071 = (inp[3]) ? 4'b0001 : node61072;
																assign node61072 = (inp[0]) ? 4'b0011 : 4'b0001;
										assign node61077 = (inp[7]) ? node61149 : node61078;
											assign node61078 = (inp[14]) ? node61114 : node61079;
												assign node61079 = (inp[2]) ? node61095 : node61080;
													assign node61080 = (inp[0]) ? node61088 : node61081;
														assign node61081 = (inp[3]) ? node61085 : node61082;
															assign node61082 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node61085 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node61088 = (inp[3]) ? node61092 : node61089;
															assign node61089 = (inp[15]) ? 4'b0010 : 4'b0000;
															assign node61092 = (inp[15]) ? 4'b0000 : 4'b0010;
													assign node61095 = (inp[15]) ? node61109 : node61096;
														assign node61096 = (inp[12]) ? node61104 : node61097;
															assign node61097 = (inp[0]) ? node61101 : node61098;
																assign node61098 = (inp[3]) ? 4'b0001 : 4'b0011;
																assign node61101 = (inp[3]) ? 4'b0011 : 4'b0001;
															assign node61104 = (inp[0]) ? 4'b0011 : node61105;
																assign node61105 = (inp[3]) ? 4'b0001 : 4'b0011;
														assign node61109 = (inp[0]) ? 4'b0001 : node61110;
															assign node61110 = (inp[3]) ? 4'b0011 : 4'b0001;
												assign node61114 = (inp[2]) ? node61136 : node61115;
													assign node61115 = (inp[12]) ? node61125 : node61116;
														assign node61116 = (inp[3]) ? 4'b0001 : node61117;
															assign node61117 = (inp[0]) ? node61121 : node61118;
																assign node61118 = (inp[15]) ? 4'b0001 : 4'b0011;
																assign node61121 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node61125 = (inp[15]) ? node61131 : node61126;
															assign node61126 = (inp[0]) ? node61128 : 4'b0001;
																assign node61128 = (inp[3]) ? 4'b0011 : 4'b0001;
															assign node61131 = (inp[0]) ? node61133 : 4'b0011;
																assign node61133 = (inp[3]) ? 4'b0001 : 4'b0011;
													assign node61136 = (inp[12]) ? node61142 : node61137;
														assign node61137 = (inp[15]) ? 4'b0011 : node61138;
															assign node61138 = (inp[3]) ? 4'b0001 : 4'b0011;
														assign node61142 = (inp[3]) ? node61146 : node61143;
															assign node61143 = (inp[15]) ? 4'b0011 : 4'b0001;
															assign node61146 = (inp[15]) ? 4'b0001 : 4'b0011;
											assign node61149 = (inp[2]) ? node61175 : node61150;
												assign node61150 = (inp[14]) ? node61164 : node61151;
													assign node61151 = (inp[3]) ? node61159 : node61152;
														assign node61152 = (inp[0]) ? node61156 : node61153;
															assign node61153 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node61156 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node61159 = (inp[12]) ? 4'b0001 : node61160;
															assign node61160 = (inp[15]) ? 4'b0011 : 4'b0001;
													assign node61164 = (inp[0]) ? node61166 : 4'b0010;
														assign node61166 = (inp[12]) ? node61168 : 4'b0000;
															assign node61168 = (inp[3]) ? node61172 : node61169;
																assign node61169 = (inp[15]) ? 4'b0010 : 4'b0000;
																assign node61172 = (inp[15]) ? 4'b0000 : 4'b0010;
												assign node61175 = (inp[3]) ? node61183 : node61176;
													assign node61176 = (inp[0]) ? node61180 : node61177;
														assign node61177 = (inp[15]) ? 4'b0000 : 4'b0010;
														assign node61180 = (inp[15]) ? 4'b0010 : 4'b0000;
													assign node61183 = (inp[14]) ? node61193 : node61184;
														assign node61184 = (inp[12]) ? node61186 : 4'b0010;
															assign node61186 = (inp[0]) ? node61190 : node61187;
																assign node61187 = (inp[15]) ? 4'b0010 : 4'b0000;
																assign node61190 = (inp[15]) ? 4'b0000 : 4'b0010;
														assign node61193 = (inp[12]) ? 4'b0010 : node61194;
															assign node61194 = (inp[0]) ? node61198 : node61195;
																assign node61195 = (inp[15]) ? 4'b0010 : 4'b0000;
																assign node61198 = (inp[15]) ? 4'b0000 : 4'b0010;
									assign node61202 = (inp[12]) ? node61350 : node61203;
										assign node61203 = (inp[3]) ? node61281 : node61204;
											assign node61204 = (inp[7]) ? node61244 : node61205;
												assign node61205 = (inp[8]) ? node61225 : node61206;
													assign node61206 = (inp[14]) ? node61218 : node61207;
														assign node61207 = (inp[2]) ? node61215 : node61208;
															assign node61208 = (inp[15]) ? node61212 : node61209;
																assign node61209 = (inp[0]) ? 4'b0011 : 4'b0001;
																assign node61212 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node61215 = (inp[0]) ? 4'b0000 : 4'b0010;
														assign node61218 = (inp[2]) ? 4'b0010 : node61219;
															assign node61219 = (inp[0]) ? node61221 : 4'b0000;
																assign node61221 = (inp[15]) ? 4'b0000 : 4'b0010;
													assign node61225 = (inp[2]) ? node61237 : node61226;
														assign node61226 = (inp[14]) ? node61232 : node61227;
															assign node61227 = (inp[15]) ? node61229 : 4'b0000;
																assign node61229 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node61232 = (inp[0]) ? node61234 : 4'b0011;
																assign node61234 = (inp[15]) ? 4'b0001 : 4'b0011;
														assign node61237 = (inp[0]) ? node61241 : node61238;
															assign node61238 = (inp[15]) ? 4'b0011 : 4'b0001;
															assign node61241 = (inp[15]) ? 4'b0001 : 4'b0011;
												assign node61244 = (inp[8]) ? node61264 : node61245;
													assign node61245 = (inp[14]) ? node61259 : node61246;
														assign node61246 = (inp[2]) ? node61254 : node61247;
															assign node61247 = (inp[15]) ? node61251 : node61248;
																assign node61248 = (inp[0]) ? 4'b0010 : 4'b0000;
																assign node61251 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node61254 = (inp[0]) ? 4'b0001 : node61255;
																assign node61255 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node61259 = (inp[15]) ? 4'b0001 : node61260;
															assign node61260 = (inp[0]) ? 4'b0011 : 4'b0001;
													assign node61264 = (inp[2]) ? node61274 : node61265;
														assign node61265 = (inp[14]) ? node61267 : 4'b0001;
															assign node61267 = (inp[0]) ? node61271 : node61268;
																assign node61268 = (inp[15]) ? 4'b0010 : 4'b0000;
																assign node61271 = (inp[15]) ? 4'b0000 : 4'b0010;
														assign node61274 = (inp[15]) ? node61278 : node61275;
															assign node61275 = (inp[0]) ? 4'b0010 : 4'b0000;
															assign node61278 = (inp[0]) ? 4'b0000 : 4'b0010;
											assign node61281 = (inp[0]) ? node61321 : node61282;
												assign node61282 = (inp[15]) ? node61302 : node61283;
													assign node61283 = (inp[7]) ? node61295 : node61284;
														assign node61284 = (inp[8]) ? node61290 : node61285;
															assign node61285 = (inp[14]) ? 4'b0000 : node61286;
																assign node61286 = (inp[2]) ? 4'b0000 : 4'b0001;
															assign node61290 = (inp[14]) ? 4'b0001 : node61291;
																assign node61291 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node61295 = (inp[2]) ? 4'b0000 : node61296;
															assign node61296 = (inp[14]) ? 4'b0000 : node61297;
																assign node61297 = (inp[8]) ? 4'b0001 : 4'b0000;
													assign node61302 = (inp[14]) ? node61314 : node61303;
														assign node61303 = (inp[8]) ? node61309 : node61304;
															assign node61304 = (inp[7]) ? node61306 : 4'b0011;
																assign node61306 = (inp[2]) ? 4'b0011 : 4'b0010;
															assign node61309 = (inp[2]) ? 4'b0010 : node61310;
																assign node61310 = (inp[7]) ? 4'b0011 : 4'b0010;
														assign node61314 = (inp[7]) ? node61318 : node61315;
															assign node61315 = (inp[8]) ? 4'b0011 : 4'b0010;
															assign node61318 = (inp[8]) ? 4'b0010 : 4'b0011;
												assign node61321 = (inp[15]) ? node61335 : node61322;
													assign node61322 = (inp[8]) ? node61328 : node61323;
														assign node61323 = (inp[14]) ? node61325 : 4'b0010;
															assign node61325 = (inp[2]) ? 4'b0010 : 4'b0011;
														assign node61328 = (inp[7]) ? node61332 : node61329;
															assign node61329 = (inp[2]) ? 4'b0011 : 4'b0010;
															assign node61332 = (inp[2]) ? 4'b0010 : 4'b0011;
													assign node61335 = (inp[7]) ? node61345 : node61336;
														assign node61336 = (inp[8]) ? node61342 : node61337;
															assign node61337 = (inp[2]) ? 4'b0000 : node61338;
																assign node61338 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node61342 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node61345 = (inp[8]) ? node61347 : 4'b0001;
															assign node61347 = (inp[2]) ? 4'b0000 : 4'b0001;
										assign node61350 = (inp[8]) ? node61390 : node61351;
											assign node61351 = (inp[7]) ? node61373 : node61352;
												assign node61352 = (inp[14]) ? node61368 : node61353;
													assign node61353 = (inp[2]) ? node61361 : node61354;
														assign node61354 = (inp[0]) ? node61358 : node61355;
															assign node61355 = (inp[15]) ? 4'b0011 : 4'b0001;
															assign node61358 = (inp[15]) ? 4'b0001 : 4'b0011;
														assign node61361 = (inp[3]) ? node61363 : 4'b0010;
															assign node61363 = (inp[0]) ? 4'b0000 : node61364;
																assign node61364 = (inp[15]) ? 4'b0010 : 4'b0000;
													assign node61368 = (inp[0]) ? 4'b0010 : node61369;
														assign node61369 = (inp[15]) ? 4'b0010 : 4'b0000;
												assign node61373 = (inp[14]) ? node61383 : node61374;
													assign node61374 = (inp[2]) ? node61380 : node61375;
														assign node61375 = (inp[3]) ? node61377 : 4'b0010;
															assign node61377 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node61380 = (inp[0]) ? 4'b0011 : 4'b0001;
													assign node61383 = (inp[15]) ? node61387 : node61384;
														assign node61384 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node61387 = (inp[0]) ? 4'b0001 : 4'b0011;
											assign node61390 = (inp[7]) ? node61424 : node61391;
												assign node61391 = (inp[14]) ? node61403 : node61392;
													assign node61392 = (inp[2]) ? node61398 : node61393;
														assign node61393 = (inp[0]) ? node61395 : 4'b0010;
															assign node61395 = (inp[15]) ? 4'b0000 : 4'b0010;
														assign node61398 = (inp[0]) ? node61400 : 4'b0001;
															assign node61400 = (inp[15]) ? 4'b0001 : 4'b0011;
													assign node61403 = (inp[3]) ? node61411 : node61404;
														assign node61404 = (inp[0]) ? node61408 : node61405;
															assign node61405 = (inp[15]) ? 4'b0011 : 4'b0001;
															assign node61408 = (inp[15]) ? 4'b0001 : 4'b0011;
														assign node61411 = (inp[2]) ? node61417 : node61412;
															assign node61412 = (inp[0]) ? 4'b0011 : node61413;
																assign node61413 = (inp[15]) ? 4'b0011 : 4'b0001;
															assign node61417 = (inp[15]) ? node61421 : node61418;
																assign node61418 = (inp[0]) ? 4'b0011 : 4'b0001;
																assign node61421 = (inp[0]) ? 4'b0001 : 4'b0011;
												assign node61424 = (inp[14]) ? node61436 : node61425;
													assign node61425 = (inp[2]) ? 4'b0000 : node61426;
														assign node61426 = (inp[3]) ? 4'b0011 : node61427;
															assign node61427 = (inp[0]) ? node61431 : node61428;
																assign node61428 = (inp[15]) ? 4'b0011 : 4'b0001;
																assign node61431 = (inp[15]) ? 4'b0001 : 4'b0011;
													assign node61436 = (inp[0]) ? node61440 : node61437;
														assign node61437 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node61440 = (inp[15]) ? 4'b0000 : 4'b0010;

endmodule