module dtc_split75_bm14 (
	input  wire [13-1:0] inp,
	output wire [1-1:0] outp
);

	wire [1-1:0] node1;
	wire [1-1:0] node2;
	wire [1-1:0] node3;
	wire [1-1:0] node4;
	wire [1-1:0] node5;
	wire [1-1:0] node7;
	wire [1-1:0] node10;
	wire [1-1:0] node11;
	wire [1-1:0] node14;
	wire [1-1:0] node17;
	wire [1-1:0] node18;
	wire [1-1:0] node19;
	wire [1-1:0] node22;
	wire [1-1:0] node25;
	wire [1-1:0] node26;
	wire [1-1:0] node29;
	wire [1-1:0] node32;
	wire [1-1:0] node33;
	wire [1-1:0] node34;
	wire [1-1:0] node35;
	wire [1-1:0] node38;
	wire [1-1:0] node41;
	wire [1-1:0] node42;
	wire [1-1:0] node45;
	wire [1-1:0] node48;
	wire [1-1:0] node49;
	wire [1-1:0] node50;
	wire [1-1:0] node53;
	wire [1-1:0] node56;
	wire [1-1:0] node57;
	wire [1-1:0] node60;
	wire [1-1:0] node63;
	wire [1-1:0] node64;
	wire [1-1:0] node65;
	wire [1-1:0] node66;
	wire [1-1:0] node67;
	wire [1-1:0] node70;
	wire [1-1:0] node73;
	wire [1-1:0] node74;
	wire [1-1:0] node77;
	wire [1-1:0] node80;
	wire [1-1:0] node81;
	wire [1-1:0] node82;
	wire [1-1:0] node85;
	wire [1-1:0] node88;
	wire [1-1:0] node89;
	wire [1-1:0] node92;
	wire [1-1:0] node95;
	wire [1-1:0] node96;
	wire [1-1:0] node97;
	wire [1-1:0] node98;
	wire [1-1:0] node101;
	wire [1-1:0] node104;
	wire [1-1:0] node105;
	wire [1-1:0] node108;
	wire [1-1:0] node111;
	wire [1-1:0] node112;
	wire [1-1:0] node113;
	wire [1-1:0] node116;
	wire [1-1:0] node119;
	wire [1-1:0] node120;
	wire [1-1:0] node123;
	wire [1-1:0] node126;
	wire [1-1:0] node127;
	wire [1-1:0] node128;
	wire [1-1:0] node129;
	wire [1-1:0] node130;
	wire [1-1:0] node131;
	wire [1-1:0] node134;
	wire [1-1:0] node137;
	wire [1-1:0] node138;
	wire [1-1:0] node141;
	wire [1-1:0] node144;
	wire [1-1:0] node145;
	wire [1-1:0] node146;
	wire [1-1:0] node149;
	wire [1-1:0] node152;
	wire [1-1:0] node153;
	wire [1-1:0] node156;
	wire [1-1:0] node159;
	wire [1-1:0] node160;
	wire [1-1:0] node161;
	wire [1-1:0] node162;
	wire [1-1:0] node165;
	wire [1-1:0] node168;
	wire [1-1:0] node169;
	wire [1-1:0] node172;
	wire [1-1:0] node175;
	wire [1-1:0] node176;
	wire [1-1:0] node177;
	wire [1-1:0] node180;
	wire [1-1:0] node183;
	wire [1-1:0] node184;
	wire [1-1:0] node187;
	wire [1-1:0] node190;
	wire [1-1:0] node191;
	wire [1-1:0] node192;
	wire [1-1:0] node193;
	wire [1-1:0] node194;
	wire [1-1:0] node197;
	wire [1-1:0] node200;
	wire [1-1:0] node201;
	wire [1-1:0] node204;
	wire [1-1:0] node207;
	wire [1-1:0] node208;
	wire [1-1:0] node209;
	wire [1-1:0] node212;
	wire [1-1:0] node215;
	wire [1-1:0] node216;
	wire [1-1:0] node219;
	wire [1-1:0] node222;
	wire [1-1:0] node223;
	wire [1-1:0] node224;
	wire [1-1:0] node225;
	wire [1-1:0] node228;
	wire [1-1:0] node231;
	wire [1-1:0] node232;
	wire [1-1:0] node235;
	wire [1-1:0] node238;
	wire [1-1:0] node239;
	wire [1-1:0] node240;
	wire [1-1:0] node243;
	wire [1-1:0] node246;
	wire [1-1:0] node247;

	assign outp = (inp[1]) ? node126 : node1;
		assign node1 = (inp[7]) ? node63 : node2;
			assign node2 = (inp[9]) ? node32 : node3;
				assign node3 = (inp[10]) ? node17 : node4;
					assign node4 = (inp[6]) ? node10 : node5;
						assign node5 = (inp[2]) ? node7 : 1'b1;
							assign node7 = (inp[0]) ? 1'b1 : 1'b1;
						assign node10 = (inp[8]) ? node14 : node11;
							assign node11 = (inp[11]) ? 1'b1 : 1'b1;
							assign node14 = (inp[2]) ? 1'b1 : 1'b1;
					assign node17 = (inp[2]) ? node25 : node18;
						assign node18 = (inp[6]) ? node22 : node19;
							assign node19 = (inp[3]) ? 1'b1 : 1'b1;
							assign node22 = (inp[0]) ? 1'b1 : 1'b1;
						assign node25 = (inp[11]) ? node29 : node26;
							assign node26 = (inp[0]) ? 1'b1 : 1'b1;
							assign node29 = (inp[8]) ? 1'b0 : 1'b1;
				assign node32 = (inp[6]) ? node48 : node33;
					assign node33 = (inp[8]) ? node41 : node34;
						assign node34 = (inp[10]) ? node38 : node35;
							assign node35 = (inp[5]) ? 1'b1 : 1'b1;
							assign node38 = (inp[12]) ? 1'b1 : 1'b1;
						assign node41 = (inp[5]) ? node45 : node42;
							assign node42 = (inp[10]) ? 1'b1 : 1'b1;
							assign node45 = (inp[11]) ? 1'b0 : 1'b1;
					assign node48 = (inp[4]) ? node56 : node49;
						assign node49 = (inp[5]) ? node53 : node50;
							assign node50 = (inp[12]) ? 1'b1 : 1'b1;
							assign node53 = (inp[3]) ? 1'b0 : 1'b1;
						assign node56 = (inp[3]) ? node60 : node57;
							assign node57 = (inp[8]) ? 1'b0 : 1'b1;
							assign node60 = (inp[11]) ? 1'b0 : 1'b0;
			assign node63 = (inp[6]) ? node95 : node64;
				assign node64 = (inp[11]) ? node80 : node65;
					assign node65 = (inp[5]) ? node73 : node66;
						assign node66 = (inp[12]) ? node70 : node67;
							assign node67 = (inp[3]) ? 1'b1 : 1'b1;
							assign node70 = (inp[4]) ? 1'b1 : 1'b1;
						assign node73 = (inp[10]) ? node77 : node74;
							assign node74 = (inp[9]) ? 1'b1 : 1'b1;
							assign node77 = (inp[0]) ? 1'b0 : 1'b1;
					assign node80 = (inp[9]) ? node88 : node81;
						assign node81 = (inp[4]) ? node85 : node82;
							assign node82 = (inp[8]) ? 1'b1 : 1'b1;
							assign node85 = (inp[3]) ? 1'b0 : 1'b1;
						assign node88 = (inp[2]) ? node92 : node89;
							assign node89 = (inp[5]) ? 1'b0 : 1'b1;
							assign node92 = (inp[8]) ? 1'b0 : 1'b0;
				assign node95 = (inp[2]) ? node111 : node96;
					assign node96 = (inp[12]) ? node104 : node97;
						assign node97 = (inp[9]) ? node101 : node98;
							assign node98 = (inp[4]) ? 1'b1 : 1'b1;
							assign node101 = (inp[10]) ? 1'b0 : 1'b1;
						assign node104 = (inp[11]) ? node108 : node105;
							assign node105 = (inp[5]) ? 1'b0 : 1'b1;
							assign node108 = (inp[3]) ? 1'b0 : 1'b0;
					assign node111 = (inp[11]) ? node119 : node112;
						assign node112 = (inp[12]) ? node116 : node113;
							assign node113 = (inp[9]) ? 1'b0 : 1'b1;
							assign node116 = (inp[3]) ? 1'b0 : 1'b0;
						assign node119 = (inp[8]) ? node123 : node120;
							assign node120 = (inp[10]) ? 1'b0 : 1'b0;
							assign node123 = (inp[3]) ? 1'b0 : 1'b0;
		assign node126 = (inp[12]) ? node190 : node127;
			assign node127 = (inp[11]) ? node159 : node128;
				assign node128 = (inp[2]) ? node144 : node129;
					assign node129 = (inp[5]) ? node137 : node130;
						assign node130 = (inp[10]) ? node134 : node131;
							assign node131 = (inp[4]) ? 1'b1 : 1'b1;
							assign node134 = (inp[4]) ? 1'b1 : 1'b1;
						assign node137 = (inp[6]) ? node141 : node138;
							assign node138 = (inp[0]) ? 1'b1 : 1'b1;
							assign node141 = (inp[3]) ? 1'b0 : 1'b1;
					assign node144 = (inp[0]) ? node152 : node145;
						assign node145 = (inp[5]) ? node149 : node146;
							assign node146 = (inp[9]) ? 1'b1 : 1'b1;
							assign node149 = (inp[4]) ? 1'b0 : 1'b1;
						assign node152 = (inp[6]) ? node156 : node153;
							assign node153 = (inp[10]) ? 1'b0 : 1'b1;
							assign node156 = (inp[7]) ? 1'b0 : 1'b0;
				assign node159 = (inp[0]) ? node175 : node160;
					assign node160 = (inp[9]) ? node168 : node161;
						assign node161 = (inp[6]) ? node165 : node162;
							assign node162 = (inp[7]) ? 1'b1 : 1'b1;
							assign node165 = (inp[8]) ? 1'b0 : 1'b1;
						assign node168 = (inp[5]) ? node172 : node169;
							assign node169 = (inp[7]) ? 1'b0 : 1'b1;
							assign node172 = (inp[4]) ? 1'b0 : 1'b0;
					assign node175 = (inp[5]) ? node183 : node176;
						assign node176 = (inp[3]) ? node180 : node177;
							assign node177 = (inp[4]) ? 1'b0 : 1'b1;
							assign node180 = (inp[2]) ? 1'b0 : 1'b0;
						assign node183 = (inp[8]) ? node187 : node184;
							assign node184 = (inp[9]) ? 1'b0 : 1'b0;
							assign node187 = (inp[9]) ? 1'b0 : 1'b0;
			assign node190 = (inp[8]) ? node222 : node191;
				assign node191 = (inp[9]) ? node207 : node192;
					assign node192 = (inp[0]) ? node200 : node193;
						assign node193 = (inp[10]) ? node197 : node194;
							assign node194 = (inp[4]) ? 1'b1 : 1'b1;
							assign node197 = (inp[11]) ? 1'b0 : 1'b1;
						assign node200 = (inp[10]) ? node204 : node201;
							assign node201 = (inp[2]) ? 1'b0 : 1'b1;
							assign node204 = (inp[6]) ? 1'b0 : 1'b0;
					assign node207 = (inp[7]) ? node215 : node208;
						assign node208 = (inp[2]) ? node212 : node209;
							assign node209 = (inp[4]) ? 1'b0 : 1'b1;
							assign node212 = (inp[11]) ? 1'b0 : 1'b0;
						assign node215 = (inp[6]) ? node219 : node216;
							assign node216 = (inp[5]) ? 1'b0 : 1'b0;
							assign node219 = (inp[3]) ? 1'b0 : 1'b0;
				assign node222 = (inp[4]) ? node238 : node223;
					assign node223 = (inp[5]) ? node231 : node224;
						assign node224 = (inp[10]) ? node228 : node225;
							assign node225 = (inp[6]) ? 1'b0 : 1'b1;
							assign node228 = (inp[9]) ? 1'b0 : 1'b0;
						assign node231 = (inp[3]) ? node235 : node232;
							assign node232 = (inp[9]) ? 1'b0 : 1'b0;
							assign node235 = (inp[6]) ? 1'b0 : 1'b0;
					assign node238 = (inp[3]) ? node246 : node239;
						assign node239 = (inp[9]) ? node243 : node240;
							assign node240 = (inp[5]) ? 1'b0 : 1'b0;
							assign node243 = (inp[6]) ? 1'b0 : 1'b0;
						assign node246 = (inp[7]) ? 1'b0 : node247;
							assign node247 = (inp[0]) ? 1'b0 : 1'b0;

endmodule