module dtc_split66_bm93 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node7;
	wire [3-1:0] node11;
	wire [3-1:0] node12;
	wire [3-1:0] node13;
	wire [3-1:0] node17;
	wire [3-1:0] node19;
	wire [3-1:0] node24;
	wire [3-1:0] node25;
	wire [3-1:0] node26;
	wire [3-1:0] node27;
	wire [3-1:0] node28;
	wire [3-1:0] node29;
	wire [3-1:0] node34;
	wire [3-1:0] node35;
	wire [3-1:0] node36;
	wire [3-1:0] node37;
	wire [3-1:0] node38;
	wire [3-1:0] node42;
	wire [3-1:0] node44;
	wire [3-1:0] node45;
	wire [3-1:0] node49;
	wire [3-1:0] node51;
	wire [3-1:0] node55;
	wire [3-1:0] node56;
	wire [3-1:0] node57;
	wire [3-1:0] node59;
	wire [3-1:0] node63;
	wire [3-1:0] node64;
	wire [3-1:0] node65;
	wire [3-1:0] node66;
	wire [3-1:0] node67;
	wire [3-1:0] node69;
	wire [3-1:0] node70;
	wire [3-1:0] node78;
	wire [3-1:0] node80;
	wire [3-1:0] node81;
	wire [3-1:0] node83;
	wire [3-1:0] node85;
	wire [3-1:0] node86;
	wire [3-1:0] node87;
	wire [3-1:0] node88;
	wire [3-1:0] node90;
	wire [3-1:0] node94;
	wire [3-1:0] node97;
	wire [3-1:0] node99;
	wire [3-1:0] node100;
	wire [3-1:0] node102;
	wire [3-1:0] node106;
	wire [3-1:0] node107;
	wire [3-1:0] node108;
	wire [3-1:0] node109;
	wire [3-1:0] node111;
	wire [3-1:0] node114;
	wire [3-1:0] node116;
	wire [3-1:0] node119;
	wire [3-1:0] node120;
	wire [3-1:0] node122;
	wire [3-1:0] node126;
	wire [3-1:0] node127;
	wire [3-1:0] node129;
	wire [3-1:0] node131;
	wire [3-1:0] node133;
	wire [3-1:0] node135;

	assign outp = (inp[0]) ? node24 : node1;
		assign node1 = (inp[3]) ? node3 : 3'b000;
			assign node3 = (inp[7]) ? 3'b000 : node4;
				assign node4 = (inp[6]) ? 3'b000 : node5;
					assign node5 = (inp[5]) ? node11 : node6;
						assign node6 = (inp[8]) ? 3'b000 : node7;
							assign node7 = (inp[4]) ? 3'b100 : 3'b000;
						assign node11 = (inp[8]) ? node17 : node12;
							assign node12 = (inp[10]) ? 3'b010 : node13;
								assign node13 = (inp[4]) ? 3'b100 : 3'b010;
							assign node17 = (inp[4]) ? node19 : 3'b100;
								assign node19 = (inp[10]) ? 3'b100 : 3'b000;
		assign node24 = (inp[7]) ? node78 : node25;
			assign node25 = (inp[3]) ? node55 : node26;
				assign node26 = (inp[5]) ? node34 : node27;
					assign node27 = (inp[8]) ? 3'b000 : node28;
						assign node28 = (inp[6]) ? 3'b000 : node29;
							assign node29 = (inp[4]) ? 3'b110 : 3'b000;
					assign node34 = (inp[6]) ? 3'b100 : node35;
						assign node35 = (inp[8]) ? node49 : node36;
							assign node36 = (inp[4]) ? node42 : node37;
								assign node37 = (inp[1]) ? 3'b100 : node38;
									assign node38 = (inp[2]) ? 3'b100 : 3'b000;
								assign node42 = (inp[10]) ? node44 : 3'b110;
									assign node44 = (inp[2]) ? 3'b100 : node45;
										assign node45 = (inp[1]) ? 3'b100 : 3'b000;
							assign node49 = (inp[4]) ? node51 : 3'b110;
								assign node51 = (inp[10]) ? 3'b110 : 3'b100;
				assign node55 = (inp[5]) ? node63 : node56;
					assign node56 = (inp[6]) ? 3'b011 : node57;
						assign node57 = (inp[4]) ? node59 : 3'b011;
							assign node59 = (inp[8]) ? 3'b011 : 3'b111;
					assign node63 = (inp[6]) ? 3'b110 : node64;
						assign node64 = (inp[8]) ? 3'b111 : node65;
							assign node65 = (inp[1]) ? 3'b111 : node66;
								assign node66 = (inp[2]) ? 3'b111 : node67;
									assign node67 = (inp[4]) ? node69 : 3'b011;
										assign node69 = (inp[10]) ? 3'b011 : node70;
											assign node70 = (inp[11]) ? 3'b011 : 3'b101;
			assign node78 = (inp[5]) ? node80 : 3'b000;
				assign node80 = (inp[3]) ? node106 : node81;
					assign node81 = (inp[2]) ? node83 : 3'b000;
						assign node83 = (inp[1]) ? node85 : 3'b000;
							assign node85 = (inp[6]) ? node97 : node86;
								assign node86 = (inp[11]) ? node94 : node87;
									assign node87 = (inp[8]) ? 3'b100 : node88;
										assign node88 = (inp[4]) ? node90 : 3'b100;
											assign node90 = (inp[10]) ? 3'b100 : 3'b000;
									assign node94 = (inp[8]) ? 3'b000 : 3'b100;
								assign node97 = (inp[4]) ? node99 : 3'b000;
									assign node99 = (inp[10]) ? 3'b000 : node100;
										assign node100 = (inp[9]) ? node102 : 3'b000;
											assign node102 = (inp[8]) ? 3'b100 : 3'b000;
					assign node106 = (inp[6]) ? node126 : node107;
						assign node107 = (inp[11]) ? node119 : node108;
							assign node108 = (inp[8]) ? node114 : node109;
								assign node109 = (inp[2]) ? node111 : 3'b011;
									assign node111 = (inp[1]) ? 3'b111 : 3'b011;
								assign node114 = (inp[1]) ? node116 : 3'b001;
									assign node116 = (inp[2]) ? 3'b101 : 3'b001;
							assign node119 = (inp[8]) ? 3'b011 : node120;
								assign node120 = (inp[1]) ? node122 : 3'b011;
									assign node122 = (inp[2]) ? 3'b111 : 3'b011;
						assign node126 = (inp[10]) ? 3'b000 : node127;
							assign node127 = (inp[1]) ? node129 : 3'b000;
								assign node129 = (inp[9]) ? node131 : 3'b000;
									assign node131 = (inp[2]) ? node133 : 3'b000;
										assign node133 = (inp[8]) ? node135 : 3'b000;
											assign node135 = (inp[4]) ? 3'b100 : 3'b000;

endmodule