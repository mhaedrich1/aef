module dtc_split33_bm6 (
	input  wire [12-1:0] inp,
	output wire [1-1:0] outp
);

	wire [1-1:0] node1;
	wire [1-1:0] node2;
	wire [1-1:0] node3;
	wire [1-1:0] node4;
	wire [1-1:0] node5;
	wire [1-1:0] node6;
	wire [1-1:0] node7;
	wire [1-1:0] node10;
	wire [1-1:0] node13;
	wire [1-1:0] node14;
	wire [1-1:0] node17;
	wire [1-1:0] node20;
	wire [1-1:0] node21;
	wire [1-1:0] node23;
	wire [1-1:0] node26;
	wire [1-1:0] node27;
	wire [1-1:0] node30;
	wire [1-1:0] node33;
	wire [1-1:0] node34;
	wire [1-1:0] node35;
	wire [1-1:0] node36;
	wire [1-1:0] node39;
	wire [1-1:0] node42;
	wire [1-1:0] node43;
	wire [1-1:0] node46;
	wire [1-1:0] node49;
	wire [1-1:0] node50;
	wire [1-1:0] node51;
	wire [1-1:0] node55;
	wire [1-1:0] node56;
	wire [1-1:0] node59;
	wire [1-1:0] node62;
	wire [1-1:0] node63;
	wire [1-1:0] node64;
	wire [1-1:0] node65;
	wire [1-1:0] node66;
	wire [1-1:0] node69;
	wire [1-1:0] node72;
	wire [1-1:0] node73;
	wire [1-1:0] node76;
	wire [1-1:0] node79;
	wire [1-1:0] node80;
	wire [1-1:0] node81;
	wire [1-1:0] node84;
	wire [1-1:0] node87;
	wire [1-1:0] node88;
	wire [1-1:0] node91;
	wire [1-1:0] node94;
	wire [1-1:0] node95;
	wire [1-1:0] node96;
	wire [1-1:0] node97;
	wire [1-1:0] node100;
	wire [1-1:0] node103;
	wire [1-1:0] node104;
	wire [1-1:0] node107;
	wire [1-1:0] node110;
	wire [1-1:0] node111;
	wire [1-1:0] node112;
	wire [1-1:0] node115;
	wire [1-1:0] node118;
	wire [1-1:0] node119;
	wire [1-1:0] node122;
	wire [1-1:0] node125;
	wire [1-1:0] node126;
	wire [1-1:0] node127;
	wire [1-1:0] node128;
	wire [1-1:0] node129;
	wire [1-1:0] node130;
	wire [1-1:0] node133;
	wire [1-1:0] node136;
	wire [1-1:0] node137;
	wire [1-1:0] node140;
	wire [1-1:0] node143;
	wire [1-1:0] node144;
	wire [1-1:0] node145;
	wire [1-1:0] node148;
	wire [1-1:0] node151;
	wire [1-1:0] node152;
	wire [1-1:0] node155;
	wire [1-1:0] node158;
	wire [1-1:0] node159;
	wire [1-1:0] node160;
	wire [1-1:0] node161;
	wire [1-1:0] node164;
	wire [1-1:0] node167;
	wire [1-1:0] node168;
	wire [1-1:0] node171;
	wire [1-1:0] node174;
	wire [1-1:0] node175;
	wire [1-1:0] node176;
	wire [1-1:0] node179;
	wire [1-1:0] node182;
	wire [1-1:0] node183;
	wire [1-1:0] node187;
	wire [1-1:0] node188;
	wire [1-1:0] node189;
	wire [1-1:0] node190;
	wire [1-1:0] node192;
	wire [1-1:0] node195;
	wire [1-1:0] node196;
	wire [1-1:0] node199;
	wire [1-1:0] node202;
	wire [1-1:0] node203;
	wire [1-1:0] node204;
	wire [1-1:0] node207;
	wire [1-1:0] node210;
	wire [1-1:0] node211;
	wire [1-1:0] node214;
	wire [1-1:0] node217;
	wire [1-1:0] node218;
	wire [1-1:0] node219;
	wire [1-1:0] node220;
	wire [1-1:0] node223;
	wire [1-1:0] node226;
	wire [1-1:0] node227;
	wire [1-1:0] node230;
	wire [1-1:0] node233;
	wire [1-1:0] node234;
	wire [1-1:0] node235;
	wire [1-1:0] node238;
	wire [1-1:0] node241;
	wire [1-1:0] node242;
	wire [1-1:0] node245;
	wire [1-1:0] node248;
	wire [1-1:0] node249;
	wire [1-1:0] node250;
	wire [1-1:0] node251;
	wire [1-1:0] node252;
	wire [1-1:0] node253;
	wire [1-1:0] node254;
	wire [1-1:0] node257;
	wire [1-1:0] node260;
	wire [1-1:0] node261;
	wire [1-1:0] node264;
	wire [1-1:0] node267;
	wire [1-1:0] node268;
	wire [1-1:0] node270;
	wire [1-1:0] node273;
	wire [1-1:0] node274;
	wire [1-1:0] node277;
	wire [1-1:0] node280;
	wire [1-1:0] node281;
	wire [1-1:0] node282;
	wire [1-1:0] node283;
	wire [1-1:0] node286;
	wire [1-1:0] node289;
	wire [1-1:0] node290;
	wire [1-1:0] node293;
	wire [1-1:0] node296;
	wire [1-1:0] node297;
	wire [1-1:0] node298;
	wire [1-1:0] node301;
	wire [1-1:0] node304;
	wire [1-1:0] node305;
	wire [1-1:0] node308;
	wire [1-1:0] node311;
	wire [1-1:0] node312;
	wire [1-1:0] node313;
	wire [1-1:0] node314;
	wire [1-1:0] node315;
	wire [1-1:0] node318;
	wire [1-1:0] node321;
	wire [1-1:0] node322;
	wire [1-1:0] node325;
	wire [1-1:0] node328;
	wire [1-1:0] node329;
	wire [1-1:0] node330;
	wire [1-1:0] node333;
	wire [1-1:0] node336;
	wire [1-1:0] node337;
	wire [1-1:0] node340;
	wire [1-1:0] node343;
	wire [1-1:0] node344;
	wire [1-1:0] node345;
	wire [1-1:0] node346;
	wire [1-1:0] node349;
	wire [1-1:0] node352;
	wire [1-1:0] node353;
	wire [1-1:0] node356;
	wire [1-1:0] node359;
	wire [1-1:0] node360;
	wire [1-1:0] node361;
	wire [1-1:0] node364;
	wire [1-1:0] node367;
	wire [1-1:0] node368;
	wire [1-1:0] node371;
	wire [1-1:0] node374;
	wire [1-1:0] node375;
	wire [1-1:0] node376;
	wire [1-1:0] node377;
	wire [1-1:0] node378;
	wire [1-1:0] node379;
	wire [1-1:0] node382;
	wire [1-1:0] node385;
	wire [1-1:0] node386;
	wire [1-1:0] node389;
	wire [1-1:0] node392;
	wire [1-1:0] node393;
	wire [1-1:0] node394;
	wire [1-1:0] node397;
	wire [1-1:0] node400;
	wire [1-1:0] node401;
	wire [1-1:0] node404;
	wire [1-1:0] node407;
	wire [1-1:0] node408;
	wire [1-1:0] node409;
	wire [1-1:0] node410;
	wire [1-1:0] node413;
	wire [1-1:0] node416;
	wire [1-1:0] node417;
	wire [1-1:0] node420;
	wire [1-1:0] node423;
	wire [1-1:0] node424;
	wire [1-1:0] node425;
	wire [1-1:0] node428;
	wire [1-1:0] node431;
	wire [1-1:0] node432;
	wire [1-1:0] node435;
	wire [1-1:0] node438;
	wire [1-1:0] node439;
	wire [1-1:0] node440;
	wire [1-1:0] node441;
	wire [1-1:0] node442;
	wire [1-1:0] node445;
	wire [1-1:0] node448;
	wire [1-1:0] node449;
	wire [1-1:0] node452;
	wire [1-1:0] node455;
	wire [1-1:0] node456;
	wire [1-1:0] node457;
	wire [1-1:0] node460;
	wire [1-1:0] node463;
	wire [1-1:0] node464;
	wire [1-1:0] node467;
	wire [1-1:0] node470;
	wire [1-1:0] node471;
	wire [1-1:0] node472;
	wire [1-1:0] node473;
	wire [1-1:0] node476;
	wire [1-1:0] node479;
	wire [1-1:0] node480;
	wire [1-1:0] node483;
	wire [1-1:0] node486;
	wire [1-1:0] node487;
	wire [1-1:0] node488;
	wire [1-1:0] node491;
	wire [1-1:0] node494;
	wire [1-1:0] node495;
	wire [1-1:0] node498;

	assign outp = (inp[10]) ? node248 : node1;
		assign node1 = (inp[9]) ? node125 : node2;
			assign node2 = (inp[8]) ? node62 : node3;
				assign node3 = (inp[2]) ? node33 : node4;
					assign node4 = (inp[4]) ? node20 : node5;
						assign node5 = (inp[7]) ? node13 : node6;
							assign node6 = (inp[0]) ? node10 : node7;
								assign node7 = (inp[1]) ? 1'b0 : 1'b1;
								assign node10 = (inp[6]) ? 1'b0 : 1'b0;
							assign node13 = (inp[11]) ? node17 : node14;
								assign node14 = (inp[6]) ? 1'b1 : 1'b1;
								assign node17 = (inp[5]) ? 1'b1 : 1'b0;
						assign node20 = (inp[7]) ? node26 : node21;
							assign node21 = (inp[1]) ? node23 : 1'b1;
								assign node23 = (inp[11]) ? 1'b1 : 1'b0;
							assign node26 = (inp[5]) ? node30 : node27;
								assign node27 = (inp[1]) ? 1'b0 : 1'b0;
								assign node30 = (inp[0]) ? 1'b0 : 1'b1;
					assign node33 = (inp[5]) ? node49 : node34;
						assign node34 = (inp[11]) ? node42 : node35;
							assign node35 = (inp[1]) ? node39 : node36;
								assign node36 = (inp[0]) ? 1'b0 : 1'b0;
								assign node39 = (inp[7]) ? 1'b1 : 1'b0;
							assign node42 = (inp[1]) ? node46 : node43;
								assign node43 = (inp[3]) ? 1'b1 : 1'b1;
								assign node46 = (inp[0]) ? 1'b0 : 1'b1;
						assign node49 = (inp[0]) ? node55 : node50;
							assign node50 = (inp[11]) ? 1'b0 : node51;
								assign node51 = (inp[4]) ? 1'b0 : 1'b0;
							assign node55 = (inp[11]) ? node59 : node56;
								assign node56 = (inp[3]) ? 1'b0 : 1'b1;
								assign node59 = (inp[3]) ? 1'b1 : 1'b0;
				assign node62 = (inp[3]) ? node94 : node63;
					assign node63 = (inp[0]) ? node79 : node64;
						assign node64 = (inp[7]) ? node72 : node65;
							assign node65 = (inp[11]) ? node69 : node66;
								assign node66 = (inp[2]) ? 1'b0 : 1'b1;
								assign node69 = (inp[1]) ? 1'b1 : 1'b0;
							assign node72 = (inp[1]) ? node76 : node73;
								assign node73 = (inp[6]) ? 1'b1 : 1'b0;
								assign node76 = (inp[2]) ? 1'b0 : 1'b0;
						assign node79 = (inp[1]) ? node87 : node80;
							assign node80 = (inp[2]) ? node84 : node81;
								assign node81 = (inp[6]) ? 1'b0 : 1'b1;
								assign node84 = (inp[4]) ? 1'b0 : 1'b0;
							assign node87 = (inp[6]) ? node91 : node88;
								assign node88 = (inp[2]) ? 1'b1 : 1'b0;
								assign node91 = (inp[7]) ? 1'b1 : 1'b1;
					assign node94 = (inp[2]) ? node110 : node95;
						assign node95 = (inp[7]) ? node103 : node96;
							assign node96 = (inp[5]) ? node100 : node97;
								assign node97 = (inp[11]) ? 1'b0 : 1'b0;
								assign node100 = (inp[6]) ? 1'b0 : 1'b1;
							assign node103 = (inp[11]) ? node107 : node104;
								assign node104 = (inp[1]) ? 1'b0 : 1'b1;
								assign node107 = (inp[5]) ? 1'b1 : 1'b1;
						assign node110 = (inp[7]) ? node118 : node111;
							assign node111 = (inp[4]) ? node115 : node112;
								assign node112 = (inp[11]) ? 1'b1 : 1'b0;
								assign node115 = (inp[6]) ? 1'b1 : 1'b1;
							assign node118 = (inp[4]) ? node122 : node119;
								assign node119 = (inp[5]) ? 1'b0 : 1'b1;
								assign node122 = (inp[5]) ? 1'b0 : 1'b0;
			assign node125 = (inp[2]) ? node187 : node126;
				assign node126 = (inp[8]) ? node158 : node127;
					assign node127 = (inp[0]) ? node143 : node128;
						assign node128 = (inp[11]) ? node136 : node129;
							assign node129 = (inp[6]) ? node133 : node130;
								assign node130 = (inp[1]) ? 1'b1 : 1'b0;
								assign node133 = (inp[3]) ? 1'b0 : 1'b1;
							assign node136 = (inp[4]) ? node140 : node137;
								assign node137 = (inp[6]) ? 1'b1 : 1'b1;
								assign node140 = (inp[5]) ? 1'b0 : 1'b1;
						assign node143 = (inp[3]) ? node151 : node144;
							assign node144 = (inp[11]) ? node148 : node145;
								assign node145 = (inp[7]) ? 1'b0 : 1'b0;
								assign node148 = (inp[1]) ? 1'b1 : 1'b0;
							assign node151 = (inp[6]) ? node155 : node152;
								assign node152 = (inp[7]) ? 1'b1 : 1'b0;
								assign node155 = (inp[5]) ? 1'b0 : 1'b0;
					assign node158 = (inp[3]) ? node174 : node159;
						assign node159 = (inp[7]) ? node167 : node160;
							assign node160 = (inp[6]) ? node164 : node161;
								assign node161 = (inp[1]) ? 1'b0 : 1'b0;
								assign node164 = (inp[0]) ? 1'b1 : 1'b0;
							assign node167 = (inp[5]) ? node171 : node168;
								assign node168 = (inp[4]) ? 1'b0 : 1'b0;
								assign node171 = (inp[4]) ? 1'b1 : 1'b0;
						assign node174 = (inp[0]) ? node182 : node175;
							assign node175 = (inp[11]) ? node179 : node176;
								assign node176 = (inp[4]) ? 1'b0 : 1'b0;
								assign node179 = (inp[4]) ? 1'b1 : 1'b0;
							assign node182 = (inp[11]) ? 1'b0 : node183;
								assign node183 = (inp[4]) ? 1'b0 : 1'b1;
				assign node187 = (inp[11]) ? node217 : node188;
					assign node188 = (inp[5]) ? node202 : node189;
						assign node189 = (inp[7]) ? node195 : node190;
							assign node190 = (inp[0]) ? node192 : 1'b1;
								assign node192 = (inp[1]) ? 1'b0 : 1'b1;
							assign node195 = (inp[0]) ? node199 : node196;
								assign node196 = (inp[6]) ? 1'b0 : 1'b0;
								assign node199 = (inp[6]) ? 1'b1 : 1'b1;
						assign node202 = (inp[1]) ? node210 : node203;
							assign node203 = (inp[4]) ? node207 : node204;
								assign node204 = (inp[0]) ? 1'b0 : 1'b1;
								assign node207 = (inp[0]) ? 1'b1 : 1'b0;
							assign node210 = (inp[8]) ? node214 : node211;
								assign node211 = (inp[6]) ? 1'b0 : 1'b1;
								assign node214 = (inp[6]) ? 1'b1 : 1'b0;
					assign node217 = (inp[8]) ? node233 : node218;
						assign node218 = (inp[1]) ? node226 : node219;
							assign node219 = (inp[4]) ? node223 : node220;
								assign node220 = (inp[5]) ? 1'b1 : 1'b1;
								assign node223 = (inp[3]) ? 1'b0 : 1'b0;
							assign node226 = (inp[0]) ? node230 : node227;
								assign node227 = (inp[7]) ? 1'b0 : 1'b0;
								assign node230 = (inp[7]) ? 1'b0 : 1'b0;
						assign node233 = (inp[1]) ? node241 : node234;
							assign node234 = (inp[4]) ? node238 : node235;
								assign node235 = (inp[0]) ? 1'b0 : 1'b0;
								assign node238 = (inp[0]) ? 1'b0 : 1'b1;
							assign node241 = (inp[3]) ? node245 : node242;
								assign node242 = (inp[0]) ? 1'b1 : 1'b1;
								assign node245 = (inp[7]) ? 1'b0 : 1'b1;
		assign node248 = (inp[7]) ? node374 : node249;
			assign node249 = (inp[9]) ? node311 : node250;
				assign node250 = (inp[0]) ? node280 : node251;
					assign node251 = (inp[4]) ? node267 : node252;
						assign node252 = (inp[8]) ? node260 : node253;
							assign node253 = (inp[11]) ? node257 : node254;
								assign node254 = (inp[5]) ? 1'b0 : 1'b1;
								assign node257 = (inp[5]) ? 1'b0 : 1'b0;
							assign node260 = (inp[1]) ? node264 : node261;
								assign node261 = (inp[2]) ? 1'b0 : 1'b0;
								assign node264 = (inp[2]) ? 1'b1 : 1'b0;
						assign node267 = (inp[3]) ? node273 : node268;
							assign node268 = (inp[5]) ? node270 : 1'b0;
								assign node270 = (inp[1]) ? 1'b0 : 1'b0;
							assign node273 = (inp[1]) ? node277 : node274;
								assign node274 = (inp[8]) ? 1'b0 : 1'b0;
								assign node277 = (inp[8]) ? 1'b1 : 1'b0;
					assign node280 = (inp[4]) ? node296 : node281;
						assign node281 = (inp[3]) ? node289 : node282;
							assign node282 = (inp[6]) ? node286 : node283;
								assign node283 = (inp[8]) ? 1'b0 : 1'b0;
								assign node286 = (inp[11]) ? 1'b0 : 1'b1;
							assign node289 = (inp[1]) ? node293 : node290;
								assign node290 = (inp[11]) ? 1'b1 : 1'b0;
								assign node293 = (inp[2]) ? 1'b1 : 1'b1;
						assign node296 = (inp[1]) ? node304 : node297;
							assign node297 = (inp[5]) ? node301 : node298;
								assign node298 = (inp[2]) ? 1'b1 : 1'b1;
								assign node301 = (inp[3]) ? 1'b0 : 1'b1;
							assign node304 = (inp[5]) ? node308 : node305;
								assign node305 = (inp[6]) ? 1'b0 : 1'b0;
								assign node308 = (inp[6]) ? 1'b0 : 1'b1;
				assign node311 = (inp[5]) ? node343 : node312;
					assign node312 = (inp[6]) ? node328 : node313;
						assign node313 = (inp[1]) ? node321 : node314;
							assign node314 = (inp[4]) ? node318 : node315;
								assign node315 = (inp[11]) ? 1'b0 : 1'b0;
								assign node318 = (inp[2]) ? 1'b0 : 1'b0;
							assign node321 = (inp[2]) ? node325 : node322;
								assign node322 = (inp[11]) ? 1'b1 : 1'b0;
								assign node325 = (inp[11]) ? 1'b0 : 1'b0;
						assign node328 = (inp[4]) ? node336 : node329;
							assign node329 = (inp[11]) ? node333 : node330;
								assign node330 = (inp[1]) ? 1'b0 : 1'b0;
								assign node333 = (inp[2]) ? 1'b1 : 1'b0;
							assign node336 = (inp[0]) ? node340 : node337;
								assign node337 = (inp[2]) ? 1'b1 : 1'b1;
								assign node340 = (inp[3]) ? 1'b1 : 1'b0;
					assign node343 = (inp[11]) ? node359 : node344;
						assign node344 = (inp[2]) ? node352 : node345;
							assign node345 = (inp[6]) ? node349 : node346;
								assign node346 = (inp[0]) ? 1'b1 : 1'b1;
								assign node349 = (inp[1]) ? 1'b0 : 1'b0;
							assign node352 = (inp[0]) ? node356 : node353;
								assign node353 = (inp[3]) ? 1'b0 : 1'b1;
								assign node356 = (inp[1]) ? 1'b1 : 1'b1;
						assign node359 = (inp[0]) ? node367 : node360;
							assign node360 = (inp[4]) ? node364 : node361;
								assign node361 = (inp[8]) ? 1'b1 : 1'b0;
								assign node364 = (inp[3]) ? 1'b0 : 1'b1;
							assign node367 = (inp[8]) ? node371 : node368;
								assign node368 = (inp[6]) ? 1'b0 : 1'b1;
								assign node371 = (inp[2]) ? 1'b0 : 1'b0;
			assign node374 = (inp[1]) ? node438 : node375;
				assign node375 = (inp[2]) ? node407 : node376;
					assign node376 = (inp[4]) ? node392 : node377;
						assign node377 = (inp[8]) ? node385 : node378;
							assign node378 = (inp[6]) ? node382 : node379;
								assign node379 = (inp[0]) ? 1'b0 : 1'b1;
								assign node382 = (inp[5]) ? 1'b0 : 1'b1;
							assign node385 = (inp[3]) ? node389 : node386;
								assign node386 = (inp[11]) ? 1'b1 : 1'b1;
								assign node389 = (inp[0]) ? 1'b1 : 1'b0;
						assign node392 = (inp[8]) ? node400 : node393;
							assign node393 = (inp[9]) ? node397 : node394;
								assign node394 = (inp[0]) ? 1'b1 : 1'b1;
								assign node397 = (inp[11]) ? 1'b1 : 1'b1;
							assign node400 = (inp[3]) ? node404 : node401;
								assign node401 = (inp[9]) ? 1'b0 : 1'b0;
								assign node404 = (inp[0]) ? 1'b1 : 1'b0;
					assign node407 = (inp[9]) ? node423 : node408;
						assign node408 = (inp[0]) ? node416 : node409;
							assign node409 = (inp[3]) ? node413 : node410;
								assign node410 = (inp[8]) ? 1'b1 : 1'b0;
								assign node413 = (inp[11]) ? 1'b1 : 1'b0;
							assign node416 = (inp[5]) ? node420 : node417;
								assign node417 = (inp[6]) ? 1'b1 : 1'b0;
								assign node420 = (inp[8]) ? 1'b1 : 1'b1;
						assign node423 = (inp[4]) ? node431 : node424;
							assign node424 = (inp[5]) ? node428 : node425;
								assign node425 = (inp[11]) ? 1'b0 : 1'b1;
								assign node428 = (inp[0]) ? 1'b1 : 1'b1;
							assign node431 = (inp[5]) ? node435 : node432;
								assign node432 = (inp[3]) ? 1'b1 : 1'b0;
								assign node435 = (inp[3]) ? 1'b0 : 1'b0;
				assign node438 = (inp[9]) ? node470 : node439;
					assign node439 = (inp[6]) ? node455 : node440;
						assign node440 = (inp[11]) ? node448 : node441;
							assign node441 = (inp[8]) ? node445 : node442;
								assign node442 = (inp[5]) ? 1'b1 : 1'b1;
								assign node445 = (inp[2]) ? 1'b0 : 1'b1;
							assign node448 = (inp[3]) ? node452 : node449;
								assign node449 = (inp[8]) ? 1'b1 : 1'b0;
								assign node452 = (inp[5]) ? 1'b1 : 1'b0;
						assign node455 = (inp[4]) ? node463 : node456;
							assign node456 = (inp[5]) ? node460 : node457;
								assign node457 = (inp[0]) ? 1'b1 : 1'b0;
								assign node460 = (inp[3]) ? 1'b0 : 1'b0;
							assign node463 = (inp[5]) ? node467 : node464;
								assign node464 = (inp[2]) ? 1'b1 : 1'b1;
								assign node467 = (inp[2]) ? 1'b0 : 1'b1;
					assign node470 = (inp[5]) ? node486 : node471;
						assign node471 = (inp[2]) ? node479 : node472;
							assign node472 = (inp[4]) ? node476 : node473;
								assign node473 = (inp[11]) ? 1'b1 : 1'b0;
								assign node476 = (inp[6]) ? 1'b0 : 1'b0;
							assign node479 = (inp[8]) ? node483 : node480;
								assign node480 = (inp[3]) ? 1'b0 : 1'b0;
								assign node483 = (inp[11]) ? 1'b0 : 1'b0;
						assign node486 = (inp[2]) ? node494 : node487;
							assign node487 = (inp[11]) ? node491 : node488;
								assign node488 = (inp[3]) ? 1'b0 : 1'b1;
								assign node491 = (inp[0]) ? 1'b0 : 1'b0;
							assign node494 = (inp[0]) ? node498 : node495;
								assign node495 = (inp[11]) ? 1'b1 : 1'b0;
								assign node498 = (inp[8]) ? 1'b1 : 1'b1;

endmodule