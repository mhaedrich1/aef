module dtc_split33_bm66 (
	input  wire [16-1:0] inp,
	output wire [4-1:0] outp
);

	wire [4-1:0] node1;
	wire [4-1:0] node2;
	wire [4-1:0] node3;
	wire [4-1:0] node4;
	wire [4-1:0] node6;
	wire [4-1:0] node7;
	wire [4-1:0] node9;
	wire [4-1:0] node11;
	wire [4-1:0] node13;
	wire [4-1:0] node14;
	wire [4-1:0] node16;
	wire [4-1:0] node18;
	wire [4-1:0] node20;
	wire [4-1:0] node23;
	wire [4-1:0] node24;
	wire [4-1:0] node26;
	wire [4-1:0] node28;
	wire [4-1:0] node32;
	wire [4-1:0] node33;
	wire [4-1:0] node34;
	wire [4-1:0] node36;
	wire [4-1:0] node39;
	wire [4-1:0] node40;
	wire [4-1:0] node41;
	wire [4-1:0] node42;
	wire [4-1:0] node44;
	wire [4-1:0] node46;
	wire [4-1:0] node53;
	wire [4-1:0] node54;
	wire [4-1:0] node56;
	wire [4-1:0] node58;
	wire [4-1:0] node60;
	wire [4-1:0] node62;
	wire [4-1:0] node65;
	wire [4-1:0] node66;
	wire [4-1:0] node68;
	wire [4-1:0] node70;
	wire [4-1:0] node72;
	wire [4-1:0] node73;
	wire [4-1:0] node75;
	wire [4-1:0] node79;
	wire [4-1:0] node80;
	wire [4-1:0] node81;
	wire [4-1:0] node82;
	wire [4-1:0] node84;
	wire [4-1:0] node86;
	wire [4-1:0] node92;
	wire [4-1:0] node93;
	wire [4-1:0] node94;
	wire [4-1:0] node95;
	wire [4-1:0] node97;
	wire [4-1:0] node99;
	wire [4-1:0] node101;
	wire [4-1:0] node102;
	wire [4-1:0] node103;
	wire [4-1:0] node105;
	wire [4-1:0] node110;
	wire [4-1:0] node111;
	wire [4-1:0] node113;
	wire [4-1:0] node114;
	wire [4-1:0] node116;
	wire [4-1:0] node117;
	wire [4-1:0] node118;
	wire [4-1:0] node120;
	wire [4-1:0] node127;
	wire [4-1:0] node128;
	wire [4-1:0] node130;
	wire [4-1:0] node132;
	wire [4-1:0] node133;
	wire [4-1:0] node135;
	wire [4-1:0] node137;
	wire [4-1:0] node141;
	wire [4-1:0] node142;
	wire [4-1:0] node143;
	wire [4-1:0] node145;
	wire [4-1:0] node147;
	wire [4-1:0] node149;
	wire [4-1:0] node154;
	wire [4-1:0] node155;
	wire [4-1:0] node156;
	wire [4-1:0] node158;
	wire [4-1:0] node160;
	wire [4-1:0] node161;
	wire [4-1:0] node162;
	wire [4-1:0] node164;
	wire [4-1:0] node166;
	wire [4-1:0] node171;
	wire [4-1:0] node172;
	wire [4-1:0] node173;
	wire [4-1:0] node174;
	wire [4-1:0] node176;
	wire [4-1:0] node178;
	wire [4-1:0] node180;
	wire [4-1:0] node182;
	wire [4-1:0] node188;
	wire [4-1:0] node189;
	wire [4-1:0] node191;
	wire [4-1:0] node194;
	wire [4-1:0] node196;
	wire [4-1:0] node198;
	wire [4-1:0] node199;
	wire [4-1:0] node201;
	wire [4-1:0] node203;
	wire [4-1:0] node205;
	wire [4-1:0] node207;
	wire [4-1:0] node211;
	wire [4-1:0] node212;
	wire [4-1:0] node213;
	wire [4-1:0] node214;
	wire [4-1:0] node215;
	wire [4-1:0] node216;
	wire [4-1:0] node217;
	wire [4-1:0] node219;
	wire [4-1:0] node220;
	wire [4-1:0] node222;
	wire [4-1:0] node224;
	wire [4-1:0] node226;
	wire [4-1:0] node231;
	wire [4-1:0] node232;
	wire [4-1:0] node234;
	wire [4-1:0] node236;
	wire [4-1:0] node238;
	wire [4-1:0] node239;
	wire [4-1:0] node243;
	wire [4-1:0] node246;
	wire [4-1:0] node247;
	wire [4-1:0] node249;
	wire [4-1:0] node251;
	wire [4-1:0] node254;
	wire [4-1:0] node255;
	wire [4-1:0] node256;
	wire [4-1:0] node258;
	wire [4-1:0] node259;
	wire [4-1:0] node261;
	wire [4-1:0] node267;
	wire [4-1:0] node269;
	wire [4-1:0] node270;
	wire [4-1:0] node272;
	wire [4-1:0] node274;
	wire [4-1:0] node276;
	wire [4-1:0] node278;
	wire [4-1:0] node281;
	wire [4-1:0] node284;
	wire [4-1:0] node285;
	wire [4-1:0] node286;
	wire [4-1:0] node287;
	wire [4-1:0] node289;
	wire [4-1:0] node291;
	wire [4-1:0] node292;
	wire [4-1:0] node294;
	wire [4-1:0] node296;
	wire [4-1:0] node301;
	wire [4-1:0] node302;
	wire [4-1:0] node303;
	wire [4-1:0] node305;
	wire [4-1:0] node306;
	wire [4-1:0] node308;
	wire [4-1:0] node310;
	wire [4-1:0] node312;
	wire [4-1:0] node316;
	wire [4-1:0] node320;
	wire [4-1:0] node321;
	wire [4-1:0] node322;
	wire [4-1:0] node323;
	wire [4-1:0] node324;
	wire [4-1:0] node326;
	wire [4-1:0] node328;
	wire [4-1:0] node333;
	wire [4-1:0] node335;
	wire [4-1:0] node336;
	wire [4-1:0] node337;
	wire [4-1:0] node338;
	wire [4-1:0] node340;
	wire [4-1:0] node342;
	wire [4-1:0] node348;
	wire [4-1:0] node350;
	wire [4-1:0] node351;
	wire [4-1:0] node352;
	wire [4-1:0] node354;
	wire [4-1:0] node355;
	wire [4-1:0] node357;
	wire [4-1:0] node363;
	wire [4-1:0] node364;
	wire [4-1:0] node365;
	wire [4-1:0] node366;
	wire [4-1:0] node367;
	wire [4-1:0] node368;
	wire [4-1:0] node371;
	wire [4-1:0] node373;
	wire [4-1:0] node375;
	wire [4-1:0] node376;
	wire [4-1:0] node378;
	wire [4-1:0] node382;
	wire [4-1:0] node383;
	wire [4-1:0] node384;
	wire [4-1:0] node386;
	wire [4-1:0] node388;
	wire [4-1:0] node392;
	wire [4-1:0] node395;
	wire [4-1:0] node396;
	wire [4-1:0] node398;
	wire [4-1:0] node399;
	wire [4-1:0] node403;
	wire [4-1:0] node405;
	wire [4-1:0] node406;
	wire [4-1:0] node408;
	wire [4-1:0] node410;
	wire [4-1:0] node414;
	wire [4-1:0] node415;
	wire [4-1:0] node416;
	wire [4-1:0] node418;
	wire [4-1:0] node420;
	wire [4-1:0] node423;
	wire [4-1:0] node425;
	wire [4-1:0] node427;
	wire [4-1:0] node428;
	wire [4-1:0] node429;
	wire [4-1:0] node431;
	wire [4-1:0] node436;
	wire [4-1:0] node438;
	wire [4-1:0] node440;
	wire [4-1:0] node442;
	wire [4-1:0] node445;
	wire [4-1:0] node446;
	wire [4-1:0] node447;
	wire [4-1:0] node448;
	wire [4-1:0] node449;
	wire [4-1:0] node450;
	wire [4-1:0] node451;
	wire [4-1:0] node452;
	wire [4-1:0] node453;
	wire [4-1:0] node455;
	wire [4-1:0] node462;
	wire [4-1:0] node463;
	wire [4-1:0] node465;
	wire [4-1:0] node467;
	wire [4-1:0] node469;
	wire [4-1:0] node471;
	wire [4-1:0] node474;
	wire [4-1:0] node478;
	wire [4-1:0] node480;
	wire [4-1:0] node481;
	wire [4-1:0] node483;
	wire [4-1:0] node485;
	wire [4-1:0] node489;
	wire [4-1:0] node490;
	wire [4-1:0] node491;
	wire [4-1:0] node492;
	wire [4-1:0] node493;
	wire [4-1:0] node495;
	wire [4-1:0] node497;
	wire [4-1:0] node502;
	wire [4-1:0] node505;
	wire [4-1:0] node507;
	wire [4-1:0] node508;
	wire [4-1:0] node510;
	wire [4-1:0] node512;
	wire [4-1:0] node514;
	wire [4-1:0] node518;
	wire [4-1:0] node519;
	wire [4-1:0] node520;
	wire [4-1:0] node521;
	wire [4-1:0] node522;
	wire [4-1:0] node523;
	wire [4-1:0] node524;
	wire [4-1:0] node526;
	wire [4-1:0] node528;
	wire [4-1:0] node529;
	wire [4-1:0] node533;
	wire [4-1:0] node535;
	wire [4-1:0] node536;
	wire [4-1:0] node538;
	wire [4-1:0] node540;
	wire [4-1:0] node544;
	wire [4-1:0] node546;
	wire [4-1:0] node548;
	wire [4-1:0] node550;
	wire [4-1:0] node553;
	wire [4-1:0] node554;
	wire [4-1:0] node556;
	wire [4-1:0] node557;
	wire [4-1:0] node558;
	wire [4-1:0] node560;
	wire [4-1:0] node561;
	wire [4-1:0] node563;
	wire [4-1:0] node569;
	wire [4-1:0] node571;
	wire [4-1:0] node572;
	wire [4-1:0] node574;
	wire [4-1:0] node576;
	wire [4-1:0] node577;
	wire [4-1:0] node579;
	wire [4-1:0] node584;
	wire [4-1:0] node585;
	wire [4-1:0] node586;
	wire [4-1:0] node587;
	wire [4-1:0] node589;
	wire [4-1:0] node591;
	wire [4-1:0] node594;
	wire [4-1:0] node596;
	wire [4-1:0] node598;
	wire [4-1:0] node600;
	wire [4-1:0] node602;
	wire [4-1:0] node606;
	wire [4-1:0] node607;
	wire [4-1:0] node608;
	wire [4-1:0] node610;
	wire [4-1:0] node612;
	wire [4-1:0] node614;
	wire [4-1:0] node616;
	wire [4-1:0] node618;
	wire [4-1:0] node620;
	wire [4-1:0] node623;
	wire [4-1:0] node624;
	wire [4-1:0] node625;
	wire [4-1:0] node626;
	wire [4-1:0] node633;
	wire [4-1:0] node634;
	wire [4-1:0] node635;
	wire [4-1:0] node636;
	wire [4-1:0] node637;
	wire [4-1:0] node638;
	wire [4-1:0] node639;
	wire [4-1:0] node641;
	wire [4-1:0] node643;
	wire [4-1:0] node648;
	wire [4-1:0] node650;
	wire [4-1:0] node652;
	wire [4-1:0] node653;
	wire [4-1:0] node655;
	wire [4-1:0] node657;
	wire [4-1:0] node661;
	wire [4-1:0] node663;
	wire [4-1:0] node666;
	wire [4-1:0] node667;
	wire [4-1:0] node668;
	wire [4-1:0] node669;
	wire [4-1:0] node672;
	wire [4-1:0] node673;
	wire [4-1:0] node674;
	wire [4-1:0] node679;
	wire [4-1:0] node680;
	wire [4-1:0] node683;
	wire [4-1:0] node684;
	wire [4-1:0] node685;
	wire [4-1:0] node687;
	wire [4-1:0] node692;
	wire [4-1:0] node693;
	wire [4-1:0] node695;
	wire [4-1:0] node697;
	wire [4-1:0] node698;
	wire [4-1:0] node700;
	wire [4-1:0] node702;
	wire [4-1:0] node706;
	wire [4-1:0] node707;
	wire [4-1:0] node708;
	wire [4-1:0] node709;
	wire [4-1:0] node710;
	wire [4-1:0] node712;
	wire [4-1:0] node714;
	wire [4-1:0] node721;
	wire [4-1:0] node722;
	wire [4-1:0] node723;
	wire [4-1:0] node725;
	wire [4-1:0] node726;
	wire [4-1:0] node728;
	wire [4-1:0] node730;
	wire [4-1:0] node732;
	wire [4-1:0] node734;
	wire [4-1:0] node738;
	wire [4-1:0] node739;
	wire [4-1:0] node741;
	wire [4-1:0] node743;
	wire [4-1:0] node745;
	wire [4-1:0] node747;
	wire [4-1:0] node751;
	wire [4-1:0] node752;
	wire [4-1:0] node753;
	wire [4-1:0] node754;
	wire [4-1:0] node756;
	wire [4-1:0] node758;
	wire [4-1:0] node759;
	wire [4-1:0] node761;
	wire [4-1:0] node766;
	wire [4-1:0] node768;
	wire [4-1:0] node770;
	wire [4-1:0] node773;
	wire [4-1:0] node775;
	wire [4-1:0] node776;
	wire [4-1:0] node778;
	wire [4-1:0] node779;
	wire [4-1:0] node780;
	wire [4-1:0] node782;
	wire [4-1:0] node788;
	wire [4-1:0] node789;
	wire [4-1:0] node790;
	wire [4-1:0] node791;
	wire [4-1:0] node792;
	wire [4-1:0] node794;
	wire [4-1:0] node796;
	wire [4-1:0] node798;
	wire [4-1:0] node800;
	wire [4-1:0] node801;
	wire [4-1:0] node803;
	wire [4-1:0] node805;
	wire [4-1:0] node809;
	wire [4-1:0] node810;
	wire [4-1:0] node811;
	wire [4-1:0] node813;
	wire [4-1:0] node816;
	wire [4-1:0] node817;
	wire [4-1:0] node818;
	wire [4-1:0] node819;
	wire [4-1:0] node821;
	wire [4-1:0] node823;
	wire [4-1:0] node829;
	wire [4-1:0] node831;
	wire [4-1:0] node833;
	wire [4-1:0] node836;
	wire [4-1:0] node837;
	wire [4-1:0] node839;
	wire [4-1:0] node841;
	wire [4-1:0] node843;
	wire [4-1:0] node844;
	wire [4-1:0] node846;
	wire [4-1:0] node850;
	wire [4-1:0] node851;
	wire [4-1:0] node852;
	wire [4-1:0] node853;
	wire [4-1:0] node855;
	wire [4-1:0] node857;
	wire [4-1:0] node862;
	wire [4-1:0] node864;
	wire [4-1:0] node865;
	wire [4-1:0] node867;
	wire [4-1:0] node868;
	wire [4-1:0] node870;
	wire [4-1:0] node872;
	wire [4-1:0] node877;
	wire [4-1:0] node878;
	wire [4-1:0] node879;
	wire [4-1:0] node880;
	wire [4-1:0] node882;
	wire [4-1:0] node884;
	wire [4-1:0] node885;
	wire [4-1:0] node886;
	wire [4-1:0] node888;
	wire [4-1:0] node893;
	wire [4-1:0] node894;
	wire [4-1:0] node896;
	wire [4-1:0] node898;
	wire [4-1:0] node900;
	wire [4-1:0] node904;
	wire [4-1:0] node905;
	wire [4-1:0] node906;
	wire [4-1:0] node908;
	wire [4-1:0] node909;
	wire [4-1:0] node911;
	wire [4-1:0] node915;
	wire [4-1:0] node916;
	wire [4-1:0] node920;
	wire [4-1:0] node921;
	wire [4-1:0] node922;
	wire [4-1:0] node923;
	wire [4-1:0] node924;
	wire [4-1:0] node925;
	wire [4-1:0] node929;
	wire [4-1:0] node930;
	wire [4-1:0] node933;
	wire [4-1:0] node934;
	wire [4-1:0] node938;
	wire [4-1:0] node940;
	wire [4-1:0] node941;
	wire [4-1:0] node942;
	wire [4-1:0] node945;
	wire [4-1:0] node948;
	wire [4-1:0] node950;
	wire [4-1:0] node953;
	wire [4-1:0] node954;
	wire [4-1:0] node956;
	wire [4-1:0] node959;
	wire [4-1:0] node961;
	wire [4-1:0] node964;
	wire [4-1:0] node965;
	wire [4-1:0] node967;
	wire [4-1:0] node968;
	wire [4-1:0] node970;
	wire [4-1:0] node972;
	wire [4-1:0] node976;
	wire [4-1:0] node977;
	wire [4-1:0] node981;
	wire [4-1:0] node982;
	wire [4-1:0] node983;
	wire [4-1:0] node985;
	wire [4-1:0] node986;
	wire [4-1:0] node990;
	wire [4-1:0] node993;
	wire [4-1:0] node994;
	wire [4-1:0] node996;
	wire [4-1:0] node997;
	wire [4-1:0] node999;
	wire [4-1:0] node1001;
	wire [4-1:0] node1003;
	wire [4-1:0] node1007;
	wire [4-1:0] node1008;
	wire [4-1:0] node1010;
	wire [4-1:0] node1012;
	wire [4-1:0] node1014;
	wire [4-1:0] node1018;
	wire [4-1:0] node1019;
	wire [4-1:0] node1020;
	wire [4-1:0] node1021;
	wire [4-1:0] node1022;
	wire [4-1:0] node1023;
	wire [4-1:0] node1024;
	wire [4-1:0] node1028;
	wire [4-1:0] node1029;
	wire [4-1:0] node1030;
	wire [4-1:0] node1031;
	wire [4-1:0] node1033;
	wire [4-1:0] node1038;
	wire [4-1:0] node1041;
	wire [4-1:0] node1042;
	wire [4-1:0] node1043;
	wire [4-1:0] node1044;
	wire [4-1:0] node1046;
	wire [4-1:0] node1048;
	wire [4-1:0] node1053;
	wire [4-1:0] node1054;
	wire [4-1:0] node1056;
	wire [4-1:0] node1058;
	wire [4-1:0] node1062;
	wire [4-1:0] node1063;
	wire [4-1:0] node1065;
	wire [4-1:0] node1066;
	wire [4-1:0] node1067;
	wire [4-1:0] node1072;
	wire [4-1:0] node1073;
	wire [4-1:0] node1075;
	wire [4-1:0] node1076;
	wire [4-1:0] node1077;
	wire [4-1:0] node1079;
	wire [4-1:0] node1084;
	wire [4-1:0] node1086;
	wire [4-1:0] node1089;
	wire [4-1:0] node1090;
	wire [4-1:0] node1091;
	wire [4-1:0] node1092;
	wire [4-1:0] node1093;
	wire [4-1:0] node1095;
	wire [4-1:0] node1097;
	wire [4-1:0] node1102;
	wire [4-1:0] node1104;
	wire [4-1:0] node1106;
	wire [4-1:0] node1107;
	wire [4-1:0] node1108;
	wire [4-1:0] node1110;
	wire [4-1:0] node1112;
	wire [4-1:0] node1116;
	wire [4-1:0] node1118;
	wire [4-1:0] node1120;
	wire [4-1:0] node1122;
	wire [4-1:0] node1125;
	wire [4-1:0] node1126;
	wire [4-1:0] node1127;
	wire [4-1:0] node1129;
	wire [4-1:0] node1133;
	wire [4-1:0] node1135;
	wire [4-1:0] node1137;
	wire [4-1:0] node1138;
	wire [4-1:0] node1140;
	wire [4-1:0] node1144;
	wire [4-1:0] node1145;
	wire [4-1:0] node1146;
	wire [4-1:0] node1147;
	wire [4-1:0] node1149;
	wire [4-1:0] node1151;
	wire [4-1:0] node1152;
	wire [4-1:0] node1154;
	wire [4-1:0] node1156;
	wire [4-1:0] node1159;
	wire [4-1:0] node1160;
	wire [4-1:0] node1162;
	wire [4-1:0] node1166;
	wire [4-1:0] node1168;
	wire [4-1:0] node1170;
	wire [4-1:0] node1171;
	wire [4-1:0] node1173;
	wire [4-1:0] node1177;
	wire [4-1:0] node1178;
	wire [4-1:0] node1179;
	wire [4-1:0] node1180;
	wire [4-1:0] node1182;
	wire [4-1:0] node1183;
	wire [4-1:0] node1185;
	wire [4-1:0] node1187;
	wire [4-1:0] node1191;
	wire [4-1:0] node1193;
	wire [4-1:0] node1194;
	wire [4-1:0] node1198;
	wire [4-1:0] node1199;
	wire [4-1:0] node1202;
	wire [4-1:0] node1205;
	wire [4-1:0] node1206;
	wire [4-1:0] node1208;
	wire [4-1:0] node1209;
	wire [4-1:0] node1211;
	wire [4-1:0] node1213;
	wire [4-1:0] node1216;
	wire [4-1:0] node1218;
	wire [4-1:0] node1220;
	wire [4-1:0] node1223;
	wire [4-1:0] node1225;
	wire [4-1:0] node1227;
	wire [4-1:0] node1228;
	wire [4-1:0] node1232;
	wire [4-1:0] node1233;
	wire [4-1:0] node1234;
	wire [4-1:0] node1235;
	wire [4-1:0] node1237;
	wire [4-1:0] node1238;
	wire [4-1:0] node1240;
	wire [4-1:0] node1242;
	wire [4-1:0] node1246;
	wire [4-1:0] node1247;
	wire [4-1:0] node1248;
	wire [4-1:0] node1249;
	wire [4-1:0] node1251;
	wire [4-1:0] node1257;
	wire [4-1:0] node1258;
	wire [4-1:0] node1259;
	wire [4-1:0] node1261;
	wire [4-1:0] node1263;
	wire [4-1:0] node1267;
	wire [4-1:0] node1269;
	wire [4-1:0] node1270;
	wire [4-1:0] node1272;
	wire [4-1:0] node1274;
	wire [4-1:0] node1276;
	wire [4-1:0] node1280;
	wire [4-1:0] node1281;
	wire [4-1:0] node1282;
	wire [4-1:0] node1284;
	wire [4-1:0] node1285;
	wire [4-1:0] node1287;
	wire [4-1:0] node1289;
	wire [4-1:0] node1292;
	wire [4-1:0] node1295;
	wire [4-1:0] node1297;
	wire [4-1:0] node1298;
	wire [4-1:0] node1300;
	wire [4-1:0] node1304;
	wire [4-1:0] node1305;
	wire [4-1:0] node1306;
	wire [4-1:0] node1307;
	wire [4-1:0] node1309;
	wire [4-1:0] node1311;
	wire [4-1:0] node1314;
	wire [4-1:0] node1316;
	wire [4-1:0] node1318;
	wire [4-1:0] node1321;
	wire [4-1:0] node1323;
	wire [4-1:0] node1324;
	wire [4-1:0] node1328;
	wire [4-1:0] node1329;
	wire [4-1:0] node1330;
	wire [4-1:0] node1331;
	wire [4-1:0] node1333;
	wire [4-1:0] node1335;
	wire [4-1:0] node1339;
	wire [4-1:0] node1341;
	wire [4-1:0] node1344;
	wire [4-1:0] node1345;
	wire [4-1:0] node1346;
	wire [4-1:0] node1348;
	wire [4-1:0] node1352;
	wire [4-1:0] node1354;
	wire [4-1:0] node1356;
	wire [4-1:0] node1358;

	assign outp = (inp[10]) ? node518 : node1;
		assign node1 = (inp[5]) ? node211 : node2;
			assign node2 = (inp[4]) ? node92 : node3;
				assign node3 = (inp[14]) ? node53 : node4;
					assign node4 = (inp[13]) ? node6 : 4'b1111;
						assign node6 = (inp[12]) ? node32 : node7;
							assign node7 = (inp[9]) ? node9 : 4'b1111;
								assign node9 = (inp[2]) ? node11 : 4'b1111;
									assign node11 = (inp[8]) ? node13 : 4'b1111;
										assign node13 = (inp[6]) ? node23 : node14;
											assign node14 = (inp[15]) ? node16 : 4'b1111;
												assign node16 = (inp[7]) ? node18 : 4'b1111;
													assign node18 = (inp[1]) ? node20 : 4'b1111;
														assign node20 = (inp[11]) ? 4'b1101 : 4'b1111;
											assign node23 = (inp[7]) ? 4'b1101 : node24;
												assign node24 = (inp[11]) ? node26 : 4'b1111;
													assign node26 = (inp[0]) ? node28 : 4'b1111;
														assign node28 = (inp[15]) ? 4'b1101 : 4'b1111;
							assign node32 = (inp[2]) ? 4'b1101 : node33;
								assign node33 = (inp[6]) ? node39 : node34;
									assign node34 = (inp[8]) ? node36 : 4'b1111;
										assign node36 = (inp[9]) ? 4'b1101 : 4'b1111;
									assign node39 = (inp[9]) ? 4'b1101 : node40;
										assign node40 = (inp[8]) ? 4'b1101 : node41;
											assign node41 = (inp[7]) ? 4'b1101 : node42;
												assign node42 = (inp[1]) ? node44 : 4'b1111;
													assign node44 = (inp[11]) ? node46 : 4'b1111;
														assign node46 = (inp[0]) ? 4'b1101 : 4'b1111;
					assign node53 = (inp[13]) ? node65 : node54;
						assign node54 = (inp[9]) ? node56 : 4'b1101;
							assign node56 = (inp[6]) ? node58 : 4'b1101;
								assign node58 = (inp[8]) ? node60 : 4'b1101;
									assign node60 = (inp[12]) ? node62 : 4'b1101;
										assign node62 = (inp[2]) ? 4'b1011 : 4'b1101;
						assign node65 = (inp[12]) ? node79 : node66;
							assign node66 = (inp[8]) ? node68 : 4'b1101;
								assign node68 = (inp[2]) ? node70 : 4'b1101;
									assign node70 = (inp[9]) ? node72 : 4'b1101;
										assign node72 = (inp[6]) ? 4'b1011 : node73;
											assign node73 = (inp[7]) ? node75 : 4'b1101;
												assign node75 = (inp[15]) ? 4'b1111 : 4'b1101;
							assign node79 = (inp[6]) ? 4'b1011 : node80;
								assign node80 = (inp[9]) ? 4'b1111 : node81;
									assign node81 = (inp[2]) ? 4'b1111 : node82;
										assign node82 = (inp[8]) ? node84 : 4'b1101;
											assign node84 = (inp[15]) ? node86 : 4'b1101;
												assign node86 = (inp[7]) ? 4'b1111 : 4'b1101;
				assign node92 = (inp[6]) ? node154 : node93;
					assign node93 = (inp[14]) ? node127 : node94;
						assign node94 = (inp[12]) ? node110 : node95;
							assign node95 = (inp[2]) ? node97 : 4'b1011;
								assign node97 = (inp[13]) ? node99 : 4'b1011;
									assign node99 = (inp[9]) ? node101 : 4'b1011;
										assign node101 = (inp[8]) ? 4'b1001 : node102;
											assign node102 = (inp[7]) ? 4'b1001 : node103;
												assign node103 = (inp[11]) ? node105 : 4'b1011;
													assign node105 = (inp[15]) ? 4'b1001 : 4'b1011;
							assign node110 = (inp[13]) ? 4'b1001 : node111;
								assign node111 = (inp[2]) ? node113 : 4'b1011;
									assign node113 = (inp[9]) ? 4'b1001 : node114;
										assign node114 = (inp[8]) ? node116 : 4'b1011;
											assign node116 = (inp[7]) ? 4'b1001 : node117;
												assign node117 = (inp[0]) ? 4'b1011 : node118;
													assign node118 = (inp[15]) ? node120 : 4'b1011;
														assign node120 = (inp[1]) ? 4'b1001 : 4'b1011;
						assign node127 = (inp[12]) ? node141 : node128;
							assign node128 = (inp[13]) ? node130 : 4'b1001;
								assign node130 = (inp[2]) ? node132 : 4'b1001;
									assign node132 = (inp[9]) ? 4'b1011 : node133;
										assign node133 = (inp[8]) ? node135 : 4'b1001;
											assign node135 = (inp[7]) ? node137 : 4'b1001;
												assign node137 = (inp[15]) ? 4'b1011 : 4'b1001;
							assign node141 = (inp[13]) ? 4'b1011 : node142;
								assign node142 = (inp[2]) ? 4'b1011 : node143;
									assign node143 = (inp[15]) ? node145 : 4'b1001;
										assign node145 = (inp[8]) ? node147 : 4'b1001;
											assign node147 = (inp[9]) ? node149 : 4'b1001;
												assign node149 = (inp[7]) ? 4'b1011 : 4'b1001;
					assign node154 = (inp[14]) ? node188 : node155;
						assign node155 = (inp[12]) ? node171 : node156;
							assign node156 = (inp[2]) ? node158 : 4'b1011;
								assign node158 = (inp[13]) ? node160 : 4'b1011;
									assign node160 = (inp[9]) ? 4'b1001 : node161;
										assign node161 = (inp[8]) ? 4'b1001 : node162;
											assign node162 = (inp[11]) ? node164 : 4'b1011;
												assign node164 = (inp[15]) ? node166 : 4'b1011;
													assign node166 = (inp[1]) ? 4'b1001 : 4'b1011;
							assign node171 = (inp[9]) ? 4'b1001 : node172;
								assign node172 = (inp[13]) ? 4'b1001 : node173;
									assign node173 = (inp[2]) ? 4'b1001 : node174;
										assign node174 = (inp[11]) ? node176 : 4'b1011;
											assign node176 = (inp[7]) ? node178 : 4'b1011;
												assign node178 = (inp[15]) ? node180 : 4'b1011;
													assign node180 = (inp[8]) ? node182 : 4'b1011;
														assign node182 = (inp[1]) ? 4'b1001 : 4'b1011;
						assign node188 = (inp[12]) ? node194 : node189;
							assign node189 = (inp[2]) ? node191 : 4'b1001;
								assign node191 = (inp[13]) ? 4'b1111 : 4'b1001;
							assign node194 = (inp[13]) ? node196 : 4'b1110;
								assign node196 = (inp[2]) ? node198 : 4'b1110;
									assign node198 = (inp[9]) ? 4'b1100 : node199;
										assign node199 = (inp[15]) ? node201 : 4'b1110;
											assign node201 = (inp[1]) ? node203 : 4'b1110;
												assign node203 = (inp[7]) ? node205 : 4'b1110;
													assign node205 = (inp[3]) ? node207 : 4'b1110;
														assign node207 = (inp[8]) ? 4'b1100 : 4'b1110;
			assign node211 = (inp[12]) ? node363 : node212;
				assign node212 = (inp[6]) ? node284 : node213;
					assign node213 = (inp[13]) ? node267 : node214;
						assign node214 = (inp[4]) ? node246 : node215;
							assign node215 = (inp[2]) ? node231 : node216;
								assign node216 = (inp[9]) ? 4'b1001 : node217;
									assign node217 = (inp[14]) ? node219 : 4'b1001;
										assign node219 = (inp[8]) ? 4'b1001 : node220;
											assign node220 = (inp[1]) ? node222 : 4'b1011;
												assign node222 = (inp[7]) ? node224 : 4'b1011;
													assign node224 = (inp[11]) ? node226 : 4'b1011;
														assign node226 = (inp[15]) ? 4'b1001 : 4'b1011;
								assign node231 = (inp[9]) ? node243 : node232;
									assign node232 = (inp[3]) ? node234 : 4'b1001;
										assign node234 = (inp[15]) ? node236 : 4'b1001;
											assign node236 = (inp[8]) ? node238 : 4'b1001;
												assign node238 = (inp[14]) ? 4'b1001 : node239;
													assign node239 = (inp[7]) ? 4'b1011 : 4'b1001;
									assign node243 = (inp[14]) ? 4'b1001 : 4'b1011;
							assign node246 = (inp[14]) ? node254 : node247;
								assign node247 = (inp[2]) ? node249 : 4'b1101;
									assign node249 = (inp[9]) ? node251 : 4'b1101;
										assign node251 = (inp[8]) ? 4'b1011 : 4'b1101;
								assign node254 = (inp[9]) ? 4'b1001 : node255;
									assign node255 = (inp[2]) ? 4'b1001 : node256;
										assign node256 = (inp[8]) ? node258 : 4'b1011;
											assign node258 = (inp[7]) ? 4'b1001 : node259;
												assign node259 = (inp[11]) ? node261 : 4'b1011;
													assign node261 = (inp[1]) ? 4'b1001 : 4'b1011;
						assign node267 = (inp[14]) ? node269 : 4'b1011;
							assign node269 = (inp[2]) ? node281 : node270;
								assign node270 = (inp[15]) ? node272 : 4'b1001;
									assign node272 = (inp[9]) ? node274 : 4'b1001;
										assign node274 = (inp[4]) ? node276 : 4'b1001;
											assign node276 = (inp[8]) ? node278 : 4'b1001;
												assign node278 = (inp[7]) ? 4'b1011 : 4'b1001;
								assign node281 = (inp[4]) ? 4'b1011 : 4'b1111;
					assign node284 = (inp[14]) ? node320 : node285;
						assign node285 = (inp[4]) ? node301 : node286;
							assign node286 = (inp[13]) ? 4'b1101 : node287;
								assign node287 = (inp[2]) ? node289 : 4'b1111;
									assign node289 = (inp[9]) ? node291 : 4'b1111;
										assign node291 = (inp[8]) ? 4'b1101 : node292;
											assign node292 = (inp[1]) ? node294 : 4'b1111;
												assign node294 = (inp[7]) ? node296 : 4'b1111;
													assign node296 = (inp[15]) ? 4'b1101 : 4'b1111;
							assign node301 = (inp[13]) ? 4'b1001 : node302;
								assign node302 = (inp[9]) ? node316 : node303;
									assign node303 = (inp[15]) ? node305 : 4'b1011;
										assign node305 = (inp[3]) ? 4'b1011 : node306;
											assign node306 = (inp[7]) ? node308 : 4'b1011;
												assign node308 = (inp[8]) ? node310 : 4'b1011;
													assign node310 = (inp[2]) ? node312 : 4'b1011;
														assign node312 = (inp[11]) ? 4'b1001 : 4'b1011;
									assign node316 = (inp[2]) ? 4'b1001 : 4'b1011;
						assign node320 = (inp[4]) ? node348 : node321;
							assign node321 = (inp[13]) ? node333 : node322;
								assign node322 = (inp[9]) ? 4'b1111 : node323;
									assign node323 = (inp[2]) ? 4'b1111 : node324;
										assign node324 = (inp[15]) ? node326 : 4'b1101;
											assign node326 = (inp[7]) ? node328 : 4'b1101;
												assign node328 = (inp[8]) ? 4'b1111 : 4'b1101;
								assign node333 = (inp[2]) ? node335 : 4'b1111;
									assign node335 = (inp[7]) ? 4'b1101 : node336;
										assign node336 = (inp[9]) ? 4'b1101 : node337;
											assign node337 = (inp[8]) ? 4'b1101 : node338;
												assign node338 = (inp[1]) ? node340 : 4'b1111;
													assign node340 = (inp[3]) ? node342 : 4'b1111;
														assign node342 = (inp[0]) ? 4'b1111 : 4'b1101;
							assign node348 = (inp[13]) ? node350 : 4'b1110;
								assign node350 = (inp[2]) ? 4'b1100 : node351;
									assign node351 = (inp[9]) ? 4'b1100 : node352;
										assign node352 = (inp[8]) ? node354 : 4'b1110;
											assign node354 = (inp[0]) ? 4'b1110 : node355;
												assign node355 = (inp[1]) ? node357 : 4'b1110;
													assign node357 = (inp[11]) ? 4'b1100 : 4'b1110;
				assign node363 = (inp[6]) ? node445 : node364;
					assign node364 = (inp[14]) ? node414 : node365;
						assign node365 = (inp[4]) ? node395 : node366;
							assign node366 = (inp[9]) ? node382 : node367;
								assign node367 = (inp[2]) ? node371 : node368;
									assign node368 = (inp[13]) ? 4'b1110 : 4'b1100;
									assign node371 = (inp[8]) ? node373 : 4'b1110;
										assign node373 = (inp[13]) ? node375 : 4'b1110;
											assign node375 = (inp[7]) ? 4'b1100 : node376;
												assign node376 = (inp[15]) ? node378 : 4'b1110;
													assign node378 = (inp[1]) ? 4'b1100 : 4'b1110;
								assign node382 = (inp[2]) ? node392 : node383;
									assign node383 = (inp[13]) ? 4'b1110 : node384;
										assign node384 = (inp[7]) ? node386 : 4'b1100;
											assign node386 = (inp[8]) ? node388 : 4'b1100;
												assign node388 = (inp[15]) ? 4'b1110 : 4'b1100;
									assign node392 = (inp[13]) ? 4'b1100 : 4'b1110;
							assign node395 = (inp[13]) ? node403 : node396;
								assign node396 = (inp[2]) ? node398 : 4'b1110;
									assign node398 = (inp[8]) ? 4'b1100 : node399;
										assign node399 = (inp[9]) ? 4'b1100 : 4'b1110;
								assign node403 = (inp[2]) ? node405 : 4'b1100;
									assign node405 = (inp[9]) ? 4'b1110 : node406;
										assign node406 = (inp[15]) ? node408 : 4'b1100;
											assign node408 = (inp[7]) ? node410 : 4'b1100;
												assign node410 = (inp[8]) ? 4'b1110 : 4'b1100;
						assign node414 = (inp[13]) ? node436 : node415;
							assign node415 = (inp[4]) ? node423 : node416;
								assign node416 = (inp[9]) ? node418 : 4'b1100;
									assign node418 = (inp[2]) ? node420 : 4'b1100;
										assign node420 = (inp[8]) ? 4'b1010 : 4'b1100;
								assign node423 = (inp[9]) ? node425 : 4'b1110;
									assign node425 = (inp[2]) ? node427 : 4'b1110;
										assign node427 = (inp[8]) ? 4'b1100 : node428;
											assign node428 = (inp[7]) ? 4'b1100 : node429;
												assign node429 = (inp[15]) ? node431 : 4'b1110;
													assign node431 = (inp[11]) ? 4'b1100 : 4'b1110;
							assign node436 = (inp[4]) ? node438 : 4'b1010;
								assign node438 = (inp[9]) ? node440 : 4'b1100;
									assign node440 = (inp[2]) ? node442 : 4'b1100;
										assign node442 = (inp[8]) ? 4'b1010 : 4'b1100;
					assign node445 = (inp[13]) ? node489 : node446;
						assign node446 = (inp[4]) ? node478 : node447;
							assign node447 = (inp[2]) ? 4'b1000 : node448;
								assign node448 = (inp[14]) ? node462 : node449;
									assign node449 = (inp[9]) ? 4'b1000 : node450;
										assign node450 = (inp[8]) ? 4'b1000 : node451;
											assign node451 = (inp[7]) ? 4'b1000 : node452;
												assign node452 = (inp[3]) ? 4'b1010 : node453;
													assign node453 = (inp[0]) ? node455 : 4'b1010;
														assign node455 = (inp[1]) ? 4'b1000 : 4'b1010;
									assign node462 = (inp[8]) ? node474 : node463;
										assign node463 = (inp[15]) ? node465 : 4'b1010;
											assign node465 = (inp[7]) ? node467 : 4'b1010;
												assign node467 = (inp[9]) ? node469 : 4'b1010;
													assign node469 = (inp[1]) ? node471 : 4'b1010;
														assign node471 = (inp[0]) ? 4'b1010 : 4'b1000;
										assign node474 = (inp[9]) ? 4'b1000 : 4'b1010;
							assign node478 = (inp[7]) ? node480 : 4'b1010;
								assign node480 = (inp[14]) ? 4'b1010 : node481;
									assign node481 = (inp[2]) ? node483 : 4'b1010;
										assign node483 = (inp[8]) ? node485 : 4'b1010;
											assign node485 = (inp[9]) ? 4'b1000 : 4'b1010;
						assign node489 = (inp[4]) ? node505 : node490;
							assign node490 = (inp[2]) ? node502 : node491;
								assign node491 = (inp[14]) ? 4'b1000 : node492;
									assign node492 = (inp[9]) ? 4'b1010 : node493;
										assign node493 = (inp[8]) ? node495 : 4'b1000;
											assign node495 = (inp[7]) ? node497 : 4'b1000;
												assign node497 = (inp[1]) ? 4'b1010 : 4'b1000;
								assign node502 = (inp[14]) ? 4'b1110 : 4'b1010;
							assign node505 = (inp[8]) ? node507 : 4'b1000;
								assign node507 = (inp[14]) ? 4'b1000 : node508;
									assign node508 = (inp[9]) ? node510 : 4'b1000;
										assign node510 = (inp[2]) ? node512 : 4'b1000;
											assign node512 = (inp[7]) ? node514 : 4'b1000;
												assign node514 = (inp[15]) ? 4'b1010 : 4'b1000;
		assign node518 = (inp[5]) ? node788 : node519;
			assign node519 = (inp[4]) ? node633 : node520;
				assign node520 = (inp[6]) ? node584 : node521;
					assign node521 = (inp[14]) ? node553 : node522;
						assign node522 = (inp[2]) ? node544 : node523;
							assign node523 = (inp[13]) ? node533 : node524;
								assign node524 = (inp[12]) ? node526 : 4'b1100;
									assign node526 = (inp[9]) ? node528 : 4'b1110;
										assign node528 = (inp[8]) ? 4'b1100 : node529;
											assign node529 = (inp[7]) ? 4'b1100 : 4'b1110;
								assign node533 = (inp[7]) ? node535 : 4'b1100;
									assign node535 = (inp[12]) ? 4'b1100 : node536;
										assign node536 = (inp[9]) ? node538 : 4'b1100;
											assign node538 = (inp[8]) ? node540 : 4'b1100;
												assign node540 = (inp[15]) ? 4'b1110 : 4'b1100;
							assign node544 = (inp[13]) ? node546 : 4'b1100;
								assign node546 = (inp[12]) ? node548 : 4'b1110;
									assign node548 = (inp[8]) ? node550 : 4'b1100;
										assign node550 = (inp[9]) ? 4'b1010 : 4'b1100;
						assign node553 = (inp[12]) ? node569 : node554;
							assign node554 = (inp[13]) ? node556 : 4'b1110;
								assign node556 = (inp[9]) ? 4'b1100 : node557;
									assign node557 = (inp[2]) ? 4'b1100 : node558;
										assign node558 = (inp[8]) ? node560 : 4'b1110;
											assign node560 = (inp[7]) ? 4'b1100 : node561;
												assign node561 = (inp[11]) ? node563 : 4'b1110;
													assign node563 = (inp[1]) ? 4'b1100 : 4'b1110;
							assign node569 = (inp[13]) ? node571 : 4'b1010;
								assign node571 = (inp[2]) ? 4'b1000 : node572;
									assign node572 = (inp[9]) ? node574 : 4'b1010;
										assign node574 = (inp[8]) ? node576 : 4'b1010;
											assign node576 = (inp[7]) ? 4'b1000 : node577;
												assign node577 = (inp[11]) ? node579 : 4'b1010;
													assign node579 = (inp[1]) ? 4'b1000 : 4'b1010;
					assign node584 = (inp[14]) ? node606 : node585;
						assign node585 = (inp[13]) ? 4'b1010 : node586;
							assign node586 = (inp[12]) ? node594 : node587;
								assign node587 = (inp[8]) ? node589 : 4'b1100;
									assign node589 = (inp[9]) ? node591 : 4'b1100;
										assign node591 = (inp[2]) ? 4'b1010 : 4'b1100;
								assign node594 = (inp[2]) ? node596 : 4'b1000;
									assign node596 = (inp[8]) ? node598 : 4'b1000;
										assign node598 = (inp[15]) ? node600 : 4'b1000;
											assign node600 = (inp[9]) ? node602 : 4'b1000;
												assign node602 = (inp[7]) ? 4'b1010 : 4'b1000;
						assign node606 = (inp[13]) ? 4'b1000 : node607;
							assign node607 = (inp[2]) ? node623 : node608;
								assign node608 = (inp[1]) ? node610 : 4'b1010;
									assign node610 = (inp[11]) ? node612 : 4'b1010;
										assign node612 = (inp[15]) ? node614 : 4'b1010;
											assign node614 = (inp[12]) ? node616 : 4'b1010;
												assign node616 = (inp[9]) ? node618 : 4'b1010;
													assign node618 = (inp[8]) ? node620 : 4'b1010;
														assign node620 = (inp[7]) ? 4'b1000 : 4'b1010;
								assign node623 = (inp[12]) ? 4'b1000 : node624;
									assign node624 = (inp[9]) ? 4'b1000 : node625;
										assign node625 = (inp[8]) ? 4'b1000 : node626;
											assign node626 = (inp[7]) ? 4'b1000 : 4'b1010;
				assign node633 = (inp[12]) ? node721 : node634;
					assign node634 = (inp[6]) ? node666 : node635;
						assign node635 = (inp[14]) ? node661 : node636;
							assign node636 = (inp[9]) ? node648 : node637;
								assign node637 = (inp[2]) ? 4'b1010 : node638;
									assign node638 = (inp[13]) ? 4'b1010 : node639;
										assign node639 = (inp[7]) ? node641 : 4'b1000;
											assign node641 = (inp[15]) ? node643 : 4'b1000;
												assign node643 = (inp[8]) ? 4'b1010 : 4'b1000;
								assign node648 = (inp[2]) ? node650 : 4'b1010;
									assign node650 = (inp[13]) ? node652 : 4'b1010;
										assign node652 = (inp[8]) ? 4'b1000 : node653;
											assign node653 = (inp[15]) ? node655 : 4'b1010;
												assign node655 = (inp[11]) ? node657 : 4'b1010;
													assign node657 = (inp[7]) ? 4'b1000 : 4'b1010;
							assign node661 = (inp[13]) ? node663 : 4'b1000;
								assign node663 = (inp[2]) ? 4'b1110 : 4'b1000;
						assign node666 = (inp[3]) ? node692 : node667;
							assign node667 = (inp[2]) ? node679 : node668;
								assign node668 = (inp[13]) ? node672 : node669;
									assign node669 = (inp[14]) ? 4'b1100 : 4'b1110;
									assign node672 = (inp[14]) ? 4'b1110 : node673;
										assign node673 = (inp[8]) ? 4'b1100 : node674;
											assign node674 = (inp[9]) ? 4'b1100 : 4'b1110;
								assign node679 = (inp[14]) ? node683 : node680;
									assign node680 = (inp[13]) ? 4'b1100 : 4'b1110;
									assign node683 = (inp[13]) ? 4'b1110 : node684;
										assign node684 = (inp[9]) ? 4'b1110 : node685;
											assign node685 = (inp[7]) ? node687 : 4'b1100;
												assign node687 = (inp[8]) ? 4'b1110 : 4'b1100;
							assign node692 = (inp[13]) ? node706 : node693;
								assign node693 = (inp[14]) ? node695 : 4'b1110;
									assign node695 = (inp[2]) ? node697 : 4'b1100;
										assign node697 = (inp[9]) ? 4'b1110 : node698;
											assign node698 = (inp[8]) ? node700 : 4'b1100;
												assign node700 = (inp[7]) ? node702 : 4'b1100;
													assign node702 = (inp[15]) ? 4'b1110 : 4'b1100;
								assign node706 = (inp[14]) ? 4'b1110 : node707;
									assign node707 = (inp[8]) ? 4'b1100 : node708;
										assign node708 = (inp[9]) ? 4'b1100 : node709;
											assign node709 = (inp[2]) ? 4'b1100 : node710;
												assign node710 = (inp[11]) ? node712 : 4'b1110;
													assign node712 = (inp[7]) ? node714 : 4'b1110;
														assign node714 = (inp[1]) ? 4'b1100 : 4'b1110;
					assign node721 = (inp[6]) ? node751 : node722;
						assign node722 = (inp[14]) ? node738 : node723;
							assign node723 = (inp[13]) ? node725 : 4'b1111;
								assign node725 = (inp[2]) ? 4'b1101 : node726;
									assign node726 = (inp[1]) ? node728 : 4'b1111;
										assign node728 = (inp[9]) ? node730 : 4'b1111;
											assign node730 = (inp[15]) ? node732 : 4'b1111;
												assign node732 = (inp[11]) ? node734 : 4'b1111;
													assign node734 = (inp[8]) ? 4'b1101 : 4'b1111;
							assign node738 = (inp[13]) ? 4'b1111 : node739;
								assign node739 = (inp[2]) ? node741 : 4'b1101;
									assign node741 = (inp[9]) ? node743 : 4'b1101;
										assign node743 = (inp[8]) ? node745 : 4'b1101;
											assign node745 = (inp[15]) ? node747 : 4'b1101;
												assign node747 = (inp[7]) ? 4'b1111 : 4'b1101;
						assign node751 = (inp[14]) ? node773 : node752;
							assign node752 = (inp[13]) ? node766 : node753;
								assign node753 = (inp[2]) ? 4'b1101 : node754;
									assign node754 = (inp[8]) ? node756 : 4'b1111;
										assign node756 = (inp[9]) ? node758 : 4'b1111;
											assign node758 = (inp[7]) ? 4'b1101 : node759;
												assign node759 = (inp[15]) ? node761 : 4'b1111;
													assign node761 = (inp[11]) ? 4'b1101 : 4'b1111;
								assign node766 = (inp[2]) ? node768 : 4'b1101;
									assign node768 = (inp[8]) ? node770 : 4'b1101;
										assign node770 = (inp[9]) ? 4'b1011 : 4'b1101;
							assign node773 = (inp[13]) ? node775 : 4'b1011;
								assign node775 = (inp[2]) ? 4'b1001 : node776;
									assign node776 = (inp[9]) ? node778 : 4'b1011;
										assign node778 = (inp[7]) ? 4'b1001 : node779;
											assign node779 = (inp[8]) ? 4'b1001 : node780;
												assign node780 = (inp[1]) ? node782 : 4'b1011;
													assign node782 = (inp[11]) ? 4'b1001 : 4'b1011;
			assign node788 = (inp[12]) ? node1018 : node789;
				assign node789 = (inp[6]) ? node877 : node790;
					assign node790 = (inp[13]) ? node836 : node791;
						assign node791 = (inp[4]) ? node809 : node792;
							assign node792 = (inp[14]) ? node794 : 4'b0111;
								assign node794 = (inp[9]) ? node796 : 4'b0111;
									assign node796 = (inp[8]) ? node798 : 4'b0111;
										assign node798 = (inp[2]) ? node800 : 4'b0111;
											assign node800 = (inp[7]) ? 4'b0101 : node801;
												assign node801 = (inp[15]) ? node803 : 4'b0111;
													assign node803 = (inp[11]) ? node805 : 4'b0111;
														assign node805 = (inp[1]) ? 4'b0101 : 4'b0111;
							assign node809 = (inp[2]) ? node829 : node810;
								assign node810 = (inp[14]) ? node816 : node811;
									assign node811 = (inp[9]) ? node813 : 4'b0111;
										assign node813 = (inp[8]) ? 4'b0101 : 4'b0111;
									assign node816 = (inp[9]) ? 4'b0101 : node817;
										assign node817 = (inp[8]) ? 4'b0101 : node818;
											assign node818 = (inp[7]) ? 4'b0101 : node819;
												assign node819 = (inp[1]) ? node821 : 4'b0111;
													assign node821 = (inp[11]) ? node823 : 4'b0111;
														assign node823 = (inp[15]) ? 4'b0101 : 4'b0111;
								assign node829 = (inp[14]) ? node831 : 4'b0101;
									assign node831 = (inp[9]) ? node833 : 4'b0101;
										assign node833 = (inp[8]) ? 4'b0011 : 4'b0101;
						assign node836 = (inp[4]) ? node850 : node837;
							assign node837 = (inp[9]) ? node839 : 4'b0101;
								assign node839 = (inp[2]) ? node841 : 4'b0101;
									assign node841 = (inp[8]) ? node843 : 4'b0101;
										assign node843 = (inp[14]) ? 4'b0011 : node844;
											assign node844 = (inp[15]) ? node846 : 4'b0101;
												assign node846 = (inp[7]) ? 4'b0111 : 4'b0101;
							assign node850 = (inp[14]) ? node862 : node851;
								assign node851 = (inp[2]) ? 4'b0111 : node852;
									assign node852 = (inp[9]) ? 4'b0111 : node853;
										assign node853 = (inp[8]) ? node855 : 4'b0101;
											assign node855 = (inp[7]) ? node857 : 4'b0101;
												assign node857 = (inp[15]) ? 4'b0111 : 4'b0101;
								assign node862 = (inp[2]) ? node864 : 4'b0011;
									assign node864 = (inp[9]) ? 4'b0001 : node865;
										assign node865 = (inp[8]) ? node867 : 4'b0011;
											assign node867 = (inp[7]) ? 4'b0001 : node868;
												assign node868 = (inp[1]) ? node870 : 4'b0011;
													assign node870 = (inp[15]) ? node872 : 4'b0011;
														assign node872 = (inp[11]) ? 4'b0001 : 4'b0011;
					assign node877 = (inp[14]) ? node981 : node878;
						assign node878 = (inp[13]) ? node904 : node879;
							assign node879 = (inp[4]) ? node893 : node880;
								assign node880 = (inp[2]) ? node882 : 4'b0011;
									assign node882 = (inp[9]) ? node884 : 4'b0011;
										assign node884 = (inp[8]) ? 4'b0001 : node885;
											assign node885 = (inp[7]) ? 4'b0001 : node886;
												assign node886 = (inp[1]) ? node888 : 4'b0011;
													assign node888 = (inp[3]) ? 4'b0001 : 4'b0011;
								assign node893 = (inp[2]) ? 4'b0011 : node894;
									assign node894 = (inp[15]) ? node896 : 4'b0001;
										assign node896 = (inp[8]) ? node898 : 4'b0001;
											assign node898 = (inp[9]) ? node900 : 4'b0001;
												assign node900 = (inp[7]) ? 4'b0011 : 4'b0001;
							assign node904 = (inp[11]) ? node920 : node905;
								assign node905 = (inp[4]) ? node915 : node906;
									assign node906 = (inp[2]) ? node908 : 4'b0001;
										assign node908 = (inp[9]) ? 4'b0011 : node909;
											assign node909 = (inp[7]) ? node911 : 4'b0001;
												assign node911 = (inp[8]) ? 4'b0011 : 4'b0001;
									assign node915 = (inp[2]) ? 4'b0001 : node916;
										assign node916 = (inp[9]) ? 4'b0001 : 4'b0011;
								assign node920 = (inp[8]) ? node964 : node921;
									assign node921 = (inp[0]) ? node953 : node922;
										assign node922 = (inp[1]) ? node938 : node923;
											assign node923 = (inp[7]) ? node929 : node924;
												assign node924 = (inp[2]) ? 4'b0011 : node925;
													assign node925 = (inp[9]) ? 4'b0001 : 4'b0011;
												assign node929 = (inp[2]) ? node933 : node930;
													assign node930 = (inp[4]) ? 4'b0011 : 4'b0001;
													assign node933 = (inp[4]) ? 4'b0001 : node934;
														assign node934 = (inp[9]) ? 4'b0011 : 4'b0001;
											assign node938 = (inp[15]) ? node940 : 4'b0001;
												assign node940 = (inp[7]) ? node948 : node941;
													assign node941 = (inp[9]) ? node945 : node942;
														assign node942 = (inp[2]) ? 4'b0001 : 4'b0011;
														assign node945 = (inp[2]) ? 4'b0001 : 4'b0001;
													assign node948 = (inp[9]) ? node950 : 4'b0001;
														assign node950 = (inp[2]) ? 4'b0011 : 4'b0001;
										assign node953 = (inp[9]) ? node959 : node954;
											assign node954 = (inp[4]) ? node956 : 4'b0001;
												assign node956 = (inp[2]) ? 4'b0001 : 4'b0011;
											assign node959 = (inp[2]) ? node961 : 4'b0001;
												assign node961 = (inp[4]) ? 4'b0001 : 4'b0011;
									assign node964 = (inp[2]) ? node976 : node965;
										assign node965 = (inp[4]) ? node967 : 4'b0001;
											assign node967 = (inp[9]) ? 4'b0001 : node968;
												assign node968 = (inp[7]) ? node970 : 4'b0011;
													assign node970 = (inp[15]) ? node972 : 4'b0011;
														assign node972 = (inp[1]) ? 4'b0001 : 4'b0011;
										assign node976 = (inp[4]) ? 4'b0001 : node977;
											assign node977 = (inp[9]) ? 4'b0011 : 4'b0001;
						assign node981 = (inp[4]) ? node993 : node982;
							assign node982 = (inp[13]) ? node990 : node983;
								assign node983 = (inp[2]) ? node985 : 4'b0011;
									assign node985 = (inp[8]) ? 4'b0001 : node986;
										assign node986 = (inp[9]) ? 4'b0001 : 4'b0011;
								assign node990 = (inp[2]) ? 4'b0111 : 4'b0001;
							assign node993 = (inp[13]) ? node1007 : node994;
								assign node994 = (inp[2]) ? node996 : 4'b0110;
									assign node996 = (inp[9]) ? 4'b0100 : node997;
										assign node997 = (inp[7]) ? node999 : 4'b0110;
											assign node999 = (inp[15]) ? node1001 : 4'b0110;
												assign node1001 = (inp[1]) ? node1003 : 4'b0110;
													assign node1003 = (inp[8]) ? 4'b0100 : 4'b0110;
								assign node1007 = (inp[2]) ? 4'b0110 : node1008;
									assign node1008 = (inp[15]) ? node1010 : 4'b0100;
										assign node1010 = (inp[8]) ? node1012 : 4'b0100;
											assign node1012 = (inp[9]) ? node1014 : 4'b0100;
												assign node1014 = (inp[7]) ? 4'b0110 : 4'b0100;
				assign node1018 = (inp[4]) ? node1144 : node1019;
					assign node1019 = (inp[14]) ? node1089 : node1020;
						assign node1020 = (inp[13]) ? node1062 : node1021;
							assign node1021 = (inp[6]) ? node1041 : node1022;
								assign node1022 = (inp[8]) ? node1028 : node1023;
									assign node1023 = (inp[2]) ? 4'b0100 : node1024;
										assign node1024 = (inp[9]) ? 4'b0100 : 4'b0110;
									assign node1028 = (inp[9]) ? node1038 : node1029;
										assign node1029 = (inp[2]) ? 4'b0100 : node1030;
											assign node1030 = (inp[7]) ? 4'b0100 : node1031;
												assign node1031 = (inp[11]) ? node1033 : 4'b0110;
													assign node1033 = (inp[3]) ? 4'b0110 : 4'b0100;
										assign node1038 = (inp[2]) ? 4'b0010 : 4'b0100;
								assign node1041 = (inp[2]) ? node1053 : node1042;
									assign node1042 = (inp[9]) ? 4'b0100 : node1043;
										assign node1043 = (inp[8]) ? 4'b0100 : node1044;
											assign node1044 = (inp[11]) ? node1046 : 4'b0110;
												assign node1046 = (inp[1]) ? node1048 : 4'b0110;
													assign node1048 = (inp[3]) ? 4'b0100 : 4'b0110;
									assign node1053 = (inp[9]) ? 4'b0110 : node1054;
										assign node1054 = (inp[8]) ? node1056 : 4'b0100;
											assign node1056 = (inp[7]) ? node1058 : 4'b0100;
												assign node1058 = (inp[15]) ? 4'b0110 : 4'b0100;
							assign node1062 = (inp[6]) ? node1072 : node1063;
								assign node1063 = (inp[2]) ? node1065 : 4'b0010;
									assign node1065 = (inp[8]) ? 4'b0000 : node1066;
										assign node1066 = (inp[7]) ? 4'b0000 : node1067;
											assign node1067 = (inp[9]) ? 4'b0000 : 4'b0010;
								assign node1072 = (inp[2]) ? node1084 : node1073;
									assign node1073 = (inp[9]) ? node1075 : 4'b0110;
										assign node1075 = (inp[8]) ? 4'b0100 : node1076;
											assign node1076 = (inp[7]) ? 4'b0100 : node1077;
												assign node1077 = (inp[15]) ? node1079 : 4'b0110;
													assign node1079 = (inp[1]) ? 4'b0100 : 4'b0110;
									assign node1084 = (inp[8]) ? node1086 : 4'b0100;
										assign node1086 = (inp[9]) ? 4'b0010 : 4'b0100;
						assign node1089 = (inp[2]) ? node1125 : node1090;
							assign node1090 = (inp[6]) ? node1102 : node1091;
								assign node1091 = (inp[13]) ? 4'b0000 : node1092;
									assign node1092 = (inp[9]) ? 4'b0010 : node1093;
										assign node1093 = (inp[8]) ? node1095 : 4'b0000;
											assign node1095 = (inp[15]) ? node1097 : 4'b0000;
												assign node1097 = (inp[7]) ? 4'b0010 : 4'b0000;
								assign node1102 = (inp[9]) ? node1104 : 4'b0010;
									assign node1104 = (inp[8]) ? node1106 : 4'b0010;
										assign node1106 = (inp[13]) ? node1116 : node1107;
											assign node1107 = (inp[7]) ? 4'b0000 : node1108;
												assign node1108 = (inp[3]) ? node1110 : 4'b0010;
													assign node1110 = (inp[11]) ? node1112 : 4'b0010;
														assign node1112 = (inp[15]) ? 4'b0000 : 4'b0010;
											assign node1116 = (inp[15]) ? node1118 : 4'b0010;
												assign node1118 = (inp[1]) ? node1120 : 4'b0010;
													assign node1120 = (inp[11]) ? node1122 : 4'b0010;
														assign node1122 = (inp[7]) ? 4'b0000 : 4'b0010;
							assign node1125 = (inp[6]) ? node1133 : node1126;
								assign node1126 = (inp[13]) ? 4'b0110 : node1127;
									assign node1127 = (inp[8]) ? node1129 : 4'b0010;
										assign node1129 = (inp[9]) ? 4'b0000 : 4'b0010;
								assign node1133 = (inp[9]) ? node1135 : 4'b0000;
									assign node1135 = (inp[15]) ? node1137 : 4'b0000;
										assign node1137 = (inp[13]) ? 4'b0000 : node1138;
											assign node1138 = (inp[7]) ? node1140 : 4'b0000;
												assign node1140 = (inp[8]) ? 4'b0010 : 4'b0000;
					assign node1144 = (inp[14]) ? node1232 : node1145;
						assign node1145 = (inp[6]) ? node1177 : node1146;
							assign node1146 = (inp[2]) ? node1166 : node1147;
								assign node1147 = (inp[9]) ? node1149 : 4'b0111;
									assign node1149 = (inp[8]) ? node1151 : 4'b0111;
										assign node1151 = (inp[13]) ? node1159 : node1152;
											assign node1152 = (inp[11]) ? node1154 : 4'b0111;
												assign node1154 = (inp[1]) ? node1156 : 4'b0111;
													assign node1156 = (inp[3]) ? 4'b0111 : 4'b0101;
											assign node1159 = (inp[7]) ? 4'b0101 : node1160;
												assign node1160 = (inp[11]) ? node1162 : 4'b0111;
													assign node1162 = (inp[1]) ? 4'b0101 : 4'b0111;
								assign node1166 = (inp[8]) ? node1168 : 4'b0101;
									assign node1168 = (inp[9]) ? node1170 : 4'b0101;
										assign node1170 = (inp[13]) ? 4'b0011 : node1171;
											assign node1171 = (inp[15]) ? node1173 : 4'b0101;
												assign node1173 = (inp[7]) ? 4'b0111 : 4'b0101;
							assign node1177 = (inp[13]) ? node1205 : node1178;
								assign node1178 = (inp[9]) ? node1198 : node1179;
									assign node1179 = (inp[7]) ? node1191 : node1180;
										assign node1180 = (inp[2]) ? node1182 : 4'b0101;
											assign node1182 = (inp[8]) ? 4'b0101 : node1183;
												assign node1183 = (inp[15]) ? node1185 : 4'b0111;
													assign node1185 = (inp[1]) ? node1187 : 4'b0111;
														assign node1187 = (inp[11]) ? 4'b0101 : 4'b0111;
										assign node1191 = (inp[15]) ? node1193 : 4'b0101;
											assign node1193 = (inp[2]) ? 4'b0101 : node1194;
												assign node1194 = (inp[8]) ? 4'b0111 : 4'b0101;
									assign node1198 = (inp[8]) ? node1202 : node1199;
										assign node1199 = (inp[2]) ? 4'b0101 : 4'b0111;
										assign node1202 = (inp[2]) ? 4'b0011 : 4'b0111;
								assign node1205 = (inp[9]) ? node1223 : node1206;
									assign node1206 = (inp[8]) ? node1208 : 4'b0011;
										assign node1208 = (inp[7]) ? node1216 : node1209;
											assign node1209 = (inp[11]) ? node1211 : 4'b0011;
												assign node1211 = (inp[3]) ? node1213 : 4'b0011;
													assign node1213 = (inp[2]) ? 4'b0011 : 4'b0001;
											assign node1216 = (inp[2]) ? node1218 : 4'b0001;
												assign node1218 = (inp[15]) ? node1220 : 4'b0011;
													assign node1220 = (inp[1]) ? 4'b0001 : 4'b0011;
									assign node1223 = (inp[15]) ? node1225 : 4'b0001;
										assign node1225 = (inp[8]) ? node1227 : 4'b0001;
											assign node1227 = (inp[2]) ? 4'b0001 : node1228;
												assign node1228 = (inp[7]) ? 4'b0011 : 4'b0001;
						assign node1232 = (inp[6]) ? node1280 : node1233;
							assign node1233 = (inp[2]) ? node1257 : node1234;
								assign node1234 = (inp[9]) ? node1246 : node1235;
									assign node1235 = (inp[13]) ? node1237 : 4'b0011;
										assign node1237 = (inp[8]) ? 4'b0001 : node1238;
											assign node1238 = (inp[7]) ? node1240 : 4'b0011;
												assign node1240 = (inp[15]) ? node1242 : 4'b0011;
													assign node1242 = (inp[11]) ? 4'b0001 : 4'b0011;
									assign node1246 = (inp[13]) ? 4'b0001 : node1247;
										assign node1247 = (inp[8]) ? 4'b0001 : node1248;
											assign node1248 = (inp[7]) ? 4'b0001 : node1249;
												assign node1249 = (inp[11]) ? node1251 : 4'b0011;
													assign node1251 = (inp[1]) ? 4'b0001 : 4'b0011;
								assign node1257 = (inp[13]) ? node1267 : node1258;
									assign node1258 = (inp[9]) ? 4'b0011 : node1259;
										assign node1259 = (inp[15]) ? node1261 : 4'b0001;
											assign node1261 = (inp[7]) ? node1263 : 4'b0001;
												assign node1263 = (inp[8]) ? 4'b0011 : 4'b0001;
									assign node1267 = (inp[9]) ? node1269 : 4'b0111;
										assign node1269 = (inp[8]) ? 4'b0101 : node1270;
											assign node1270 = (inp[15]) ? node1272 : 4'b0111;
												assign node1272 = (inp[1]) ? node1274 : 4'b0111;
													assign node1274 = (inp[7]) ? node1276 : 4'b0111;
														assign node1276 = (inp[11]) ? 4'b0101 : 4'b0111;
							assign node1280 = (inp[13]) ? node1304 : node1281;
								assign node1281 = (inp[9]) ? node1295 : node1282;
									assign node1282 = (inp[8]) ? node1284 : 4'b0110;
										assign node1284 = (inp[2]) ? node1292 : node1285;
											assign node1285 = (inp[15]) ? node1287 : 4'b0110;
												assign node1287 = (inp[1]) ? node1289 : 4'b0110;
													assign node1289 = (inp[11]) ? 4'b0100 : 4'b0110;
											assign node1292 = (inp[7]) ? 4'b0100 : 4'b0110;
									assign node1295 = (inp[8]) ? node1297 : 4'b0100;
										assign node1297 = (inp[2]) ? 4'b0010 : node1298;
											assign node1298 = (inp[7]) ? node1300 : 4'b0100;
												assign node1300 = (inp[15]) ? 4'b0110 : 4'b0100;
								assign node1304 = (inp[2]) ? node1328 : node1305;
									assign node1305 = (inp[8]) ? node1321 : node1306;
										assign node1306 = (inp[7]) ? node1314 : node1307;
											assign node1307 = (inp[3]) ? node1309 : 4'b0010;
												assign node1309 = (inp[11]) ? node1311 : 4'b0010;
													assign node1311 = (inp[1]) ? 4'b0000 : 4'b0010;
											assign node1314 = (inp[9]) ? node1316 : 4'b0000;
												assign node1316 = (inp[1]) ? node1318 : 4'b0010;
													assign node1318 = (inp[11]) ? 4'b0000 : 4'b0010;
										assign node1321 = (inp[7]) ? node1323 : 4'b0000;
											assign node1323 = (inp[9]) ? 4'b0000 : node1324;
												assign node1324 = (inp[15]) ? 4'b0010 : 4'b0000;
									assign node1328 = (inp[9]) ? node1344 : node1329;
										assign node1329 = (inp[8]) ? node1339 : node1330;
											assign node1330 = (inp[0]) ? 4'b0110 : node1331;
												assign node1331 = (inp[11]) ? node1333 : 4'b0110;
													assign node1333 = (inp[3]) ? node1335 : 4'b0100;
														assign node1335 = (inp[1]) ? 4'b0100 : 4'b0110;
											assign node1339 = (inp[15]) ? node1341 : 4'b0100;
												assign node1341 = (inp[7]) ? 4'b0110 : 4'b0100;
										assign node1344 = (inp[8]) ? node1352 : node1345;
											assign node1345 = (inp[7]) ? 4'b0100 : node1346;
												assign node1346 = (inp[11]) ? node1348 : 4'b0110;
													assign node1348 = (inp[15]) ? 4'b0100 : 4'b0110;
											assign node1352 = (inp[7]) ? node1354 : 4'b0010;
												assign node1354 = (inp[15]) ? node1356 : 4'b0000;
													assign node1356 = (inp[3]) ? node1358 : 4'b0010;
														assign node1358 = (inp[11]) ? 4'b0000 : 4'b0010;

endmodule