module dtc_split33_bm5 (
	input  wire [10-1:0] inp,
	output wire [1-1:0] outp
);

	wire [1-1:0] node1;
	wire [1-1:0] node2;
	wire [1-1:0] node3;
	wire [1-1:0] node4;
	wire [1-1:0] node5;
	wire [1-1:0] node6;
	wire [1-1:0] node9;
	wire [1-1:0] node12;
	wire [1-1:0] node13;
	wire [1-1:0] node16;
	wire [1-1:0] node19;
	wire [1-1:0] node20;
	wire [1-1:0] node22;
	wire [1-1:0] node25;
	wire [1-1:0] node26;
	wire [1-1:0] node29;
	wire [1-1:0] node32;
	wire [1-1:0] node33;
	wire [1-1:0] node35;
	wire [1-1:0] node36;
	wire [1-1:0] node40;
	wire [1-1:0] node41;
	wire [1-1:0] node42;
	wire [1-1:0] node46;
	wire [1-1:0] node47;
	wire [1-1:0] node50;
	wire [1-1:0] node53;
	wire [1-1:0] node54;
	wire [1-1:0] node55;
	wire [1-1:0] node56;
	wire [1-1:0] node57;
	wire [1-1:0] node60;
	wire [1-1:0] node63;
	wire [1-1:0] node64;
	wire [1-1:0] node67;
	wire [1-1:0] node70;
	wire [1-1:0] node71;
	wire [1-1:0] node72;
	wire [1-1:0] node75;
	wire [1-1:0] node78;
	wire [1-1:0] node79;
	wire [1-1:0] node82;
	wire [1-1:0] node85;
	wire [1-1:0] node86;
	wire [1-1:0] node87;
	wire [1-1:0] node88;
	wire [1-1:0] node91;
	wire [1-1:0] node94;
	wire [1-1:0] node96;
	wire [1-1:0] node99;
	wire [1-1:0] node101;
	wire [1-1:0] node104;
	wire [1-1:0] node105;
	wire [1-1:0] node106;
	wire [1-1:0] node107;
	wire [1-1:0] node108;
	wire [1-1:0] node109;
	wire [1-1:0] node113;
	wire [1-1:0] node114;
	wire [1-1:0] node117;
	wire [1-1:0] node120;
	wire [1-1:0] node121;
	wire [1-1:0] node122;
	wire [1-1:0] node126;
	wire [1-1:0] node128;
	wire [1-1:0] node131;
	wire [1-1:0] node132;
	wire [1-1:0] node133;
	wire [1-1:0] node134;
	wire [1-1:0] node138;
	wire [1-1:0] node139;
	wire [1-1:0] node142;
	wire [1-1:0] node145;
	wire [1-1:0] node146;
	wire [1-1:0] node147;
	wire [1-1:0] node150;
	wire [1-1:0] node153;
	wire [1-1:0] node154;
	wire [1-1:0] node157;
	wire [1-1:0] node160;
	wire [1-1:0] node161;
	wire [1-1:0] node162;
	wire [1-1:0] node163;
	wire [1-1:0] node165;
	wire [1-1:0] node168;
	wire [1-1:0] node170;
	wire [1-1:0] node173;
	wire [1-1:0] node174;
	wire [1-1:0] node176;
	wire [1-1:0] node179;
	wire [1-1:0] node180;
	wire [1-1:0] node183;
	wire [1-1:0] node186;
	wire [1-1:0] node187;
	wire [1-1:0] node188;
	wire [1-1:0] node189;
	wire [1-1:0] node194;
	wire [1-1:0] node195;
	wire [1-1:0] node196;
	wire [1-1:0] node199;
	wire [1-1:0] node202;
	wire [1-1:0] node203;
	wire [1-1:0] node206;

	assign outp = (inp[8]) ? node104 : node1;
		assign node1 = (inp[6]) ? node53 : node2;
			assign node2 = (inp[4]) ? node32 : node3;
				assign node3 = (inp[2]) ? node19 : node4;
					assign node4 = (inp[1]) ? node12 : node5;
						assign node5 = (inp[9]) ? node9 : node6;
							assign node6 = (inp[5]) ? 1'b0 : 1'b1;
							assign node9 = (inp[5]) ? 1'b1 : 1'b0;
						assign node12 = (inp[7]) ? node16 : node13;
							assign node13 = (inp[5]) ? 1'b0 : 1'b0;
							assign node16 = (inp[5]) ? 1'b0 : 1'b0;
					assign node19 = (inp[7]) ? node25 : node20;
						assign node20 = (inp[1]) ? node22 : 1'b1;
							assign node22 = (inp[5]) ? 1'b1 : 1'b0;
						assign node25 = (inp[0]) ? node29 : node26;
							assign node26 = (inp[3]) ? 1'b0 : 1'b1;
							assign node29 = (inp[3]) ? 1'b0 : 1'b0;
				assign node32 = (inp[2]) ? node40 : node33;
					assign node33 = (inp[7]) ? node35 : 1'b1;
						assign node35 = (inp[5]) ? 1'b1 : node36;
							assign node36 = (inp[9]) ? 1'b0 : 1'b1;
					assign node40 = (inp[3]) ? node46 : node41;
						assign node41 = (inp[5]) ? 1'b1 : node42;
							assign node42 = (inp[1]) ? 1'b1 : 1'b0;
						assign node46 = (inp[1]) ? node50 : node47;
							assign node47 = (inp[0]) ? 1'b1 : 1'b0;
							assign node50 = (inp[5]) ? 1'b0 : 1'b0;
			assign node53 = (inp[5]) ? node85 : node54;
				assign node54 = (inp[7]) ? node70 : node55;
					assign node55 = (inp[9]) ? node63 : node56;
						assign node56 = (inp[3]) ? node60 : node57;
							assign node57 = (inp[1]) ? 1'b0 : 1'b1;
							assign node60 = (inp[0]) ? 1'b1 : 1'b1;
						assign node63 = (inp[2]) ? node67 : node64;
							assign node64 = (inp[3]) ? 1'b0 : 1'b0;
							assign node67 = (inp[4]) ? 1'b0 : 1'b1;
					assign node70 = (inp[9]) ? node78 : node71;
						assign node71 = (inp[2]) ? node75 : node72;
							assign node72 = (inp[4]) ? 1'b0 : 1'b1;
							assign node75 = (inp[3]) ? 1'b1 : 1'b0;
						assign node78 = (inp[4]) ? node82 : node79;
							assign node79 = (inp[3]) ? 1'b1 : 1'b0;
							assign node82 = (inp[1]) ? 1'b1 : 1'b1;
				assign node85 = (inp[4]) ? node99 : node86;
					assign node86 = (inp[9]) ? node94 : node87;
						assign node87 = (inp[7]) ? node91 : node88;
							assign node88 = (inp[1]) ? 1'b0 : 1'b0;
							assign node91 = (inp[1]) ? 1'b1 : 1'b0;
						assign node94 = (inp[2]) ? node96 : 1'b1;
							assign node96 = (inp[7]) ? 1'b1 : 1'b0;
					assign node99 = (inp[2]) ? node101 : 1'b0;
						assign node101 = (inp[3]) ? 1'b1 : 1'b0;
		assign node104 = (inp[9]) ? node160 : node105;
			assign node105 = (inp[1]) ? node131 : node106;
				assign node106 = (inp[3]) ? node120 : node107;
					assign node107 = (inp[5]) ? node113 : node108;
						assign node108 = (inp[7]) ? 1'b1 : node109;
							assign node109 = (inp[6]) ? 1'b1 : 1'b0;
						assign node113 = (inp[7]) ? node117 : node114;
							assign node114 = (inp[4]) ? 1'b1 : 1'b0;
							assign node117 = (inp[6]) ? 1'b0 : 1'b0;
					assign node120 = (inp[4]) ? node126 : node121;
						assign node121 = (inp[2]) ? 1'b1 : node122;
							assign node122 = (inp[5]) ? 1'b0 : 1'b1;
						assign node126 = (inp[6]) ? node128 : 1'b1;
							assign node128 = (inp[7]) ? 1'b0 : 1'b1;
				assign node131 = (inp[6]) ? node145 : node132;
					assign node132 = (inp[3]) ? node138 : node133;
						assign node133 = (inp[5]) ? 1'b0 : node134;
							assign node134 = (inp[7]) ? 1'b1 : 1'b0;
						assign node138 = (inp[7]) ? node142 : node139;
							assign node139 = (inp[2]) ? 1'b1 : 1'b0;
							assign node142 = (inp[0]) ? 1'b0 : 1'b0;
					assign node145 = (inp[0]) ? node153 : node146;
						assign node146 = (inp[3]) ? node150 : node147;
							assign node147 = (inp[2]) ? 1'b1 : 1'b0;
							assign node150 = (inp[7]) ? 1'b0 : 1'b0;
						assign node153 = (inp[7]) ? node157 : node154;
							assign node154 = (inp[4]) ? 1'b1 : 1'b1;
							assign node157 = (inp[2]) ? 1'b1 : 1'b0;
			assign node160 = (inp[0]) ? node186 : node161;
				assign node161 = (inp[4]) ? node173 : node162;
					assign node162 = (inp[1]) ? node168 : node163;
						assign node163 = (inp[6]) ? node165 : 1'b1;
							assign node165 = (inp[7]) ? 1'b0 : 1'b1;
						assign node168 = (inp[2]) ? node170 : 1'b0;
							assign node170 = (inp[3]) ? 1'b1 : 1'b0;
					assign node173 = (inp[7]) ? node179 : node174;
						assign node174 = (inp[2]) ? node176 : 1'b0;
							assign node176 = (inp[1]) ? 1'b1 : 1'b0;
						assign node179 = (inp[5]) ? node183 : node180;
							assign node180 = (inp[1]) ? 1'b0 : 1'b0;
							assign node183 = (inp[3]) ? 1'b0 : 1'b1;
				assign node186 = (inp[1]) ? node194 : node187;
					assign node187 = (inp[4]) ? 1'b0 : node188;
						assign node188 = (inp[5]) ? 1'b0 : node189;
							assign node189 = (inp[6]) ? 1'b0 : 1'b0;
					assign node194 = (inp[7]) ? node202 : node195;
						assign node195 = (inp[2]) ? node199 : node196;
							assign node196 = (inp[4]) ? 1'b0 : 1'b1;
							assign node199 = (inp[3]) ? 1'b0 : 1'b0;
						assign node202 = (inp[2]) ? node206 : node203;
							assign node203 = (inp[6]) ? 1'b0 : 1'b0;
							assign node206 = (inp[6]) ? 1'b1 : 1'b0;

endmodule