module dtc_split33_bm45 (
	input  wire [16-1:0] inp,
	output wire [46-1:0] outp
);

	wire [46-1:0] node1;
	wire [46-1:0] node2;
	wire [46-1:0] node5;
	wire [46-1:0] node6;
	wire [46-1:0] node7;
	wire [46-1:0] node9;
	wire [46-1:0] node11;
	wire [46-1:0] node13;
	wire [46-1:0] node14;
	wire [46-1:0] node16;
	wire [46-1:0] node18;
	wire [46-1:0] node20;
	wire [46-1:0] node24;
	wire [46-1:0] node26;
	wire [46-1:0] node27;
	wire [46-1:0] node29;
	wire [46-1:0] node31;
	wire [46-1:0] node33;
	wire [46-1:0] node35;
	wire [46-1:0] node37;
	wire [46-1:0] node39;
	wire [46-1:0] node43;
	wire [46-1:0] node44;
	wire [46-1:0] node45;
	wire [46-1:0] node46;
	wire [46-1:0] node47;
	wire [46-1:0] node51;
	wire [46-1:0] node53;
	wire [46-1:0] node55;
	wire [46-1:0] node57;
	wire [46-1:0] node59;
	wire [46-1:0] node60;
	wire [46-1:0] node61;
	wire [46-1:0] node62;
	wire [46-1:0] node65;
	wire [46-1:0] node67;
	wire [46-1:0] node70;
	wire [46-1:0] node71;
	wire [46-1:0] node73;
	wire [46-1:0] node74;
	wire [46-1:0] node80;
	wire [46-1:0] node81;
	wire [46-1:0] node82;
	wire [46-1:0] node86;
	wire [46-1:0] node87;
	wire [46-1:0] node90;
	wire [46-1:0] node93;
	wire [46-1:0] node94;
	wire [46-1:0] node95;
	wire [46-1:0] node96;
	wire [46-1:0] node100;
	wire [46-1:0] node102;
	wire [46-1:0] node104;
	wire [46-1:0] node106;
	wire [46-1:0] node107;
	wire [46-1:0] node109;
	wire [46-1:0] node111;
	wire [46-1:0] node112;
	wire [46-1:0] node113;
	wire [46-1:0] node116;
	wire [46-1:0] node119;
	wire [46-1:0] node122;
	wire [46-1:0] node123;
	wire [46-1:0] node124;
	wire [46-1:0] node125;
	wire [46-1:0] node126;
	wire [46-1:0] node130;
	wire [46-1:0] node133;
	wire [46-1:0] node136;
	wire [46-1:0] node138;
	wire [46-1:0] node139;
	wire [46-1:0] node140;
	wire [46-1:0] node145;
	wire [46-1:0] node146;
	wire [46-1:0] node147;
	wire [46-1:0] node150;
	wire [46-1:0] node152;
	wire [46-1:0] node154;
	wire [46-1:0] node155;
	wire [46-1:0] node157;
	wire [46-1:0] node158;
	wire [46-1:0] node159;
	wire [46-1:0] node162;
	wire [46-1:0] node163;
	wire [46-1:0] node167;
	wire [46-1:0] node169;
	wire [46-1:0] node171;
	wire [46-1:0] node175;
	wire [46-1:0] node177;
	wire [46-1:0] node179;
	wire [46-1:0] node180;
	wire [46-1:0] node182;
	wire [46-1:0] node184;
	wire [46-1:0] node185;
	wire [46-1:0] node189;
	wire [46-1:0] node191;
	wire [46-1:0] node192;
	wire [46-1:0] node194;
	wire [46-1:0] node197;
	wire [46-1:0] node198;
	wire [46-1:0] node199;
	wire [46-1:0] node202;
	wire [46-1:0] node205;
	wire [46-1:0] node206;
	wire [46-1:0] node210;
	wire [46-1:0] node211;
	wire [46-1:0] node212;
	wire [46-1:0] node215;
	wire [46-1:0] node216;
	wire [46-1:0] node217;
	wire [46-1:0] node218;
	wire [46-1:0] node219;
	wire [46-1:0] node222;
	wire [46-1:0] node225;
	wire [46-1:0] node226;
	wire [46-1:0] node229;
	wire [46-1:0] node232;
	wire [46-1:0] node233;
	wire [46-1:0] node234;
	wire [46-1:0] node237;
	wire [46-1:0] node240;
	wire [46-1:0] node241;
	wire [46-1:0] node244;
	wire [46-1:0] node247;
	wire [46-1:0] node248;
	wire [46-1:0] node249;
	wire [46-1:0] node250;
	wire [46-1:0] node253;
	wire [46-1:0] node256;
	wire [46-1:0] node257;
	wire [46-1:0] node260;
	wire [46-1:0] node263;
	wire [46-1:0] node264;
	wire [46-1:0] node265;
	wire [46-1:0] node268;
	wire [46-1:0] node271;
	wire [46-1:0] node272;
	wire [46-1:0] node275;
	wire [46-1:0] node278;
	wire [46-1:0] node279;
	wire [46-1:0] node282;
	wire [46-1:0] node284;
	wire [46-1:0] node285;
	wire [46-1:0] node286;
	wire [46-1:0] node287;
	wire [46-1:0] node288;
	wire [46-1:0] node289;
	wire [46-1:0] node290;
	wire [46-1:0] node291;
	wire [46-1:0] node292;
	wire [46-1:0] node294;
	wire [46-1:0] node296;
	wire [46-1:0] node297;
	wire [46-1:0] node300;
	wire [46-1:0] node303;
	wire [46-1:0] node304;
	wire [46-1:0] node306;
	wire [46-1:0] node307;
	wire [46-1:0] node311;
	wire [46-1:0] node313;
	wire [46-1:0] node316;
	wire [46-1:0] node317;
	wire [46-1:0] node320;
	wire [46-1:0] node321;
	wire [46-1:0] node324;
	wire [46-1:0] node325;
	wire [46-1:0] node327;
	wire [46-1:0] node330;
	wire [46-1:0] node332;
	wire [46-1:0] node335;
	wire [46-1:0] node336;
	wire [46-1:0] node337;
	wire [46-1:0] node339;
	wire [46-1:0] node342;
	wire [46-1:0] node343;
	wire [46-1:0] node344;
	wire [46-1:0] node347;
	wire [46-1:0] node350;
	wire [46-1:0] node351;
	wire [46-1:0] node355;
	wire [46-1:0] node356;
	wire [46-1:0] node357;
	wire [46-1:0] node359;
	wire [46-1:0] node362;
	wire [46-1:0] node363;
	wire [46-1:0] node367;
	wire [46-1:0] node368;
	wire [46-1:0] node371;
	wire [46-1:0] node372;
	wire [46-1:0] node376;
	wire [46-1:0] node377;
	wire [46-1:0] node378;
	wire [46-1:0] node379;
	wire [46-1:0] node380;
	wire [46-1:0] node383;
	wire [46-1:0] node385;
	wire [46-1:0] node388;
	wire [46-1:0] node389;
	wire [46-1:0] node392;
	wire [46-1:0] node395;
	wire [46-1:0] node396;
	wire [46-1:0] node397;
	wire [46-1:0] node398;
	wire [46-1:0] node400;
	wire [46-1:0] node405;
	wire [46-1:0] node406;
	wire [46-1:0] node409;
	wire [46-1:0] node410;
	wire [46-1:0] node414;
	wire [46-1:0] node415;
	wire [46-1:0] node416;
	wire [46-1:0] node417;
	wire [46-1:0] node419;
	wire [46-1:0] node422;
	wire [46-1:0] node424;
	wire [46-1:0] node426;
	wire [46-1:0] node429;
	wire [46-1:0] node430;
	wire [46-1:0] node434;
	wire [46-1:0] node435;
	wire [46-1:0] node436;
	wire [46-1:0] node437;
	wire [46-1:0] node441;
	wire [46-1:0] node442;
	wire [46-1:0] node446;
	wire [46-1:0] node447;
	wire [46-1:0] node449;
	wire [46-1:0] node452;
	wire [46-1:0] node453;
	wire [46-1:0] node457;
	wire [46-1:0] node458;
	wire [46-1:0] node459;
	wire [46-1:0] node460;
	wire [46-1:0] node461;
	wire [46-1:0] node462;
	wire [46-1:0] node463;
	wire [46-1:0] node467;
	wire [46-1:0] node470;
	wire [46-1:0] node471;
	wire [46-1:0] node474;
	wire [46-1:0] node475;
	wire [46-1:0] node476;
	wire [46-1:0] node481;
	wire [46-1:0] node482;
	wire [46-1:0] node483;
	wire [46-1:0] node486;
	wire [46-1:0] node487;
	wire [46-1:0] node490;
	wire [46-1:0] node493;
	wire [46-1:0] node495;
	wire [46-1:0] node498;
	wire [46-1:0] node499;
	wire [46-1:0] node500;
	wire [46-1:0] node501;
	wire [46-1:0] node503;
	wire [46-1:0] node506;
	wire [46-1:0] node507;
	wire [46-1:0] node511;
	wire [46-1:0] node512;
	wire [46-1:0] node515;
	wire [46-1:0] node517;
	wire [46-1:0] node520;
	wire [46-1:0] node521;
	wire [46-1:0] node522;
	wire [46-1:0] node523;
	wire [46-1:0] node528;
	wire [46-1:0] node529;
	wire [46-1:0] node530;
	wire [46-1:0] node534;
	wire [46-1:0] node535;
	wire [46-1:0] node536;
	wire [46-1:0] node541;
	wire [46-1:0] node542;
	wire [46-1:0] node543;
	wire [46-1:0] node544;
	wire [46-1:0] node545;
	wire [46-1:0] node548;
	wire [46-1:0] node549;
	wire [46-1:0] node552;
	wire [46-1:0] node555;
	wire [46-1:0] node557;
	wire [46-1:0] node558;
	wire [46-1:0] node561;
	wire [46-1:0] node563;
	wire [46-1:0] node566;
	wire [46-1:0] node567;
	wire [46-1:0] node568;
	wire [46-1:0] node571;
	wire [46-1:0] node573;
	wire [46-1:0] node574;
	wire [46-1:0] node578;
	wire [46-1:0] node580;
	wire [46-1:0] node583;
	wire [46-1:0] node584;
	wire [46-1:0] node585;
	wire [46-1:0] node586;
	wire [46-1:0] node587;
	wire [46-1:0] node588;
	wire [46-1:0] node592;
	wire [46-1:0] node595;
	wire [46-1:0] node598;
	wire [46-1:0] node599;
	wire [46-1:0] node602;
	wire [46-1:0] node604;
	wire [46-1:0] node607;
	wire [46-1:0] node608;
	wire [46-1:0] node609;
	wire [46-1:0] node612;
	wire [46-1:0] node613;
	wire [46-1:0] node617;
	wire [46-1:0] node618;
	wire [46-1:0] node619;
	wire [46-1:0] node623;
	wire [46-1:0] node624;
	wire [46-1:0] node628;
	wire [46-1:0] node629;
	wire [46-1:0] node630;
	wire [46-1:0] node632;
	wire [46-1:0] node633;
	wire [46-1:0] node634;
	wire [46-1:0] node635;
	wire [46-1:0] node638;
	wire [46-1:0] node639;
	wire [46-1:0] node640;
	wire [46-1:0] node645;
	wire [46-1:0] node646;
	wire [46-1:0] node647;
	wire [46-1:0] node651;
	wire [46-1:0] node654;
	wire [46-1:0] node655;
	wire [46-1:0] node656;
	wire [46-1:0] node658;
	wire [46-1:0] node663;
	wire [46-1:0] node664;
	wire [46-1:0] node665;
	wire [46-1:0] node667;
	wire [46-1:0] node670;
	wire [46-1:0] node671;
	wire [46-1:0] node672;
	wire [46-1:0] node673;
	wire [46-1:0] node677;
	wire [46-1:0] node679;
	wire [46-1:0] node682;
	wire [46-1:0] node683;
	wire [46-1:0] node685;
	wire [46-1:0] node686;
	wire [46-1:0] node689;
	wire [46-1:0] node695;
	wire [46-1:0] node696;
	wire [46-1:0] node697;
	wire [46-1:0] node699;
	wire [46-1:0] node701;
	wire [46-1:0] node702;
	wire [46-1:0] node704;
	wire [46-1:0] node705;
	wire [46-1:0] node706;
	wire [46-1:0] node708;
	wire [46-1:0] node712;
	wire [46-1:0] node713;
	wire [46-1:0] node714;
	wire [46-1:0] node718;
	wire [46-1:0] node719;
	wire [46-1:0] node723;
	wire [46-1:0] node724;
	wire [46-1:0] node725;
	wire [46-1:0] node730;
	wire [46-1:0] node731;
	wire [46-1:0] node732;
	wire [46-1:0] node733;
	wire [46-1:0] node734;
	wire [46-1:0] node735;
	wire [46-1:0] node736;
	wire [46-1:0] node737;
	wire [46-1:0] node742;
	wire [46-1:0] node745;
	wire [46-1:0] node746;
	wire [46-1:0] node748;
	wire [46-1:0] node751;
	wire [46-1:0] node754;
	wire [46-1:0] node755;
	wire [46-1:0] node756;
	wire [46-1:0] node759;
	wire [46-1:0] node762;
	wire [46-1:0] node763;
	wire [46-1:0] node764;
	wire [46-1:0] node767;
	wire [46-1:0] node770;
	wire [46-1:0] node771;
	wire [46-1:0] node775;
	wire [46-1:0] node776;
	wire [46-1:0] node777;
	wire [46-1:0] node779;
	wire [46-1:0] node782;
	wire [46-1:0] node783;
	wire [46-1:0] node786;
	wire [46-1:0] node787;
	wire [46-1:0] node790;
	wire [46-1:0] node793;
	wire [46-1:0] node794;
	wire [46-1:0] node795;
	wire [46-1:0] node797;
	wire [46-1:0] node800;
	wire [46-1:0] node801;
	wire [46-1:0] node802;
	wire [46-1:0] node807;
	wire [46-1:0] node808;
	wire [46-1:0] node809;
	wire [46-1:0] node811;
	wire [46-1:0] node814;
	wire [46-1:0] node817;
	wire [46-1:0] node819;
	wire [46-1:0] node822;
	wire [46-1:0] node823;
	wire [46-1:0] node824;
	wire [46-1:0] node825;
	wire [46-1:0] node826;
	wire [46-1:0] node829;
	wire [46-1:0] node832;
	wire [46-1:0] node835;
	wire [46-1:0] node836;
	wire [46-1:0] node838;
	wire [46-1:0] node839;
	wire [46-1:0] node843;
	wire [46-1:0] node844;
	wire [46-1:0] node846;
	wire [46-1:0] node849;
	wire [46-1:0] node850;
	wire [46-1:0] node852;
	wire [46-1:0] node856;
	wire [46-1:0] node857;
	wire [46-1:0] node859;
	wire [46-1:0] node860;
	wire [46-1:0] node863;
	wire [46-1:0] node864;
	wire [46-1:0] node867;
	wire [46-1:0] node868;
	wire [46-1:0] node872;
	wire [46-1:0] node873;
	wire [46-1:0] node874;
	wire [46-1:0] node875;
	wire [46-1:0] node878;
	wire [46-1:0] node881;
	wire [46-1:0] node882;
	wire [46-1:0] node884;
	wire [46-1:0] node887;
	wire [46-1:0] node890;
	wire [46-1:0] node892;
	wire [46-1:0] node895;
	wire [46-1:0] node896;
	wire [46-1:0] node897;
	wire [46-1:0] node898;
	wire [46-1:0] node899;
	wire [46-1:0] node900;
	wire [46-1:0] node901;
	wire [46-1:0] node905;
	wire [46-1:0] node906;
	wire [46-1:0] node909;
	wire [46-1:0] node910;
	wire [46-1:0] node911;
	wire [46-1:0] node916;
	wire [46-1:0] node917;
	wire [46-1:0] node918;
	wire [46-1:0] node919;
	wire [46-1:0] node923;
	wire [46-1:0] node924;
	wire [46-1:0] node928;
	wire [46-1:0] node930;
	wire [46-1:0] node933;
	wire [46-1:0] node934;
	wire [46-1:0] node935;
	wire [46-1:0] node936;
	wire [46-1:0] node937;
	wire [46-1:0] node940;
	wire [46-1:0] node943;
	wire [46-1:0] node946;
	wire [46-1:0] node947;
	wire [46-1:0] node948;
	wire [46-1:0] node952;
	wire [46-1:0] node955;
	wire [46-1:0] node956;
	wire [46-1:0] node957;
	wire [46-1:0] node960;
	wire [46-1:0] node963;
	wire [46-1:0] node965;
	wire [46-1:0] node966;
	wire [46-1:0] node969;
	wire [46-1:0] node972;
	wire [46-1:0] node973;
	wire [46-1:0] node974;
	wire [46-1:0] node975;
	wire [46-1:0] node976;
	wire [46-1:0] node977;
	wire [46-1:0] node980;
	wire [46-1:0] node984;
	wire [46-1:0] node985;
	wire [46-1:0] node988;
	wire [46-1:0] node990;
	wire [46-1:0] node992;
	wire [46-1:0] node995;
	wire [46-1:0] node996;
	wire [46-1:0] node997;
	wire [46-1:0] node1000;
	wire [46-1:0] node1001;
	wire [46-1:0] node1004;
	wire [46-1:0] node1006;
	wire [46-1:0] node1009;
	wire [46-1:0] node1010;
	wire [46-1:0] node1011;
	wire [46-1:0] node1013;
	wire [46-1:0] node1017;
	wire [46-1:0] node1018;
	wire [46-1:0] node1022;
	wire [46-1:0] node1023;
	wire [46-1:0] node1024;
	wire [46-1:0] node1025;
	wire [46-1:0] node1026;
	wire [46-1:0] node1030;
	wire [46-1:0] node1033;
	wire [46-1:0] node1034;
	wire [46-1:0] node1035;
	wire [46-1:0] node1038;
	wire [46-1:0] node1042;
	wire [46-1:0] node1043;
	wire [46-1:0] node1044;
	wire [46-1:0] node1045;
	wire [46-1:0] node1050;
	wire [46-1:0] node1051;
	wire [46-1:0] node1052;
	wire [46-1:0] node1056;
	wire [46-1:0] node1057;
	wire [46-1:0] node1058;
	wire [46-1:0] node1062;
	wire [46-1:0] node1065;
	wire [46-1:0] node1066;
	wire [46-1:0] node1067;
	wire [46-1:0] node1068;
	wire [46-1:0] node1069;
	wire [46-1:0] node1070;
	wire [46-1:0] node1072;
	wire [46-1:0] node1073;
	wire [46-1:0] node1077;
	wire [46-1:0] node1078;
	wire [46-1:0] node1082;
	wire [46-1:0] node1083;
	wire [46-1:0] node1085;
	wire [46-1:0] node1088;
	wire [46-1:0] node1091;
	wire [46-1:0] node1092;
	wire [46-1:0] node1095;
	wire [46-1:0] node1097;
	wire [46-1:0] node1099;
	wire [46-1:0] node1102;
	wire [46-1:0] node1103;
	wire [46-1:0] node1104;
	wire [46-1:0] node1105;
	wire [46-1:0] node1107;
	wire [46-1:0] node1110;
	wire [46-1:0] node1112;
	wire [46-1:0] node1115;
	wire [46-1:0] node1116;
	wire [46-1:0] node1117;
	wire [46-1:0] node1118;
	wire [46-1:0] node1121;
	wire [46-1:0] node1125;
	wire [46-1:0] node1127;
	wire [46-1:0] node1128;
	wire [46-1:0] node1131;
	wire [46-1:0] node1134;
	wire [46-1:0] node1135;
	wire [46-1:0] node1136;
	wire [46-1:0] node1138;
	wire [46-1:0] node1141;
	wire [46-1:0] node1144;
	wire [46-1:0] node1145;
	wire [46-1:0] node1146;
	wire [46-1:0] node1149;
	wire [46-1:0] node1152;
	wire [46-1:0] node1153;
	wire [46-1:0] node1157;
	wire [46-1:0] node1158;
	wire [46-1:0] node1159;
	wire [46-1:0] node1160;
	wire [46-1:0] node1161;
	wire [46-1:0] node1162;
	wire [46-1:0] node1166;
	wire [46-1:0] node1168;
	wire [46-1:0] node1170;
	wire [46-1:0] node1173;
	wire [46-1:0] node1174;
	wire [46-1:0] node1175;
	wire [46-1:0] node1179;
	wire [46-1:0] node1180;
	wire [46-1:0] node1183;
	wire [46-1:0] node1186;
	wire [46-1:0] node1187;
	wire [46-1:0] node1188;
	wire [46-1:0] node1191;
	wire [46-1:0] node1192;
	wire [46-1:0] node1196;
	wire [46-1:0] node1198;
	wire [46-1:0] node1200;
	wire [46-1:0] node1202;
	wire [46-1:0] node1205;
	wire [46-1:0] node1206;
	wire [46-1:0] node1207;
	wire [46-1:0] node1208;
	wire [46-1:0] node1211;
	wire [46-1:0] node1212;
	wire [46-1:0] node1216;
	wire [46-1:0] node1217;
	wire [46-1:0] node1218;
	wire [46-1:0] node1223;
	wire [46-1:0] node1224;
	wire [46-1:0] node1225;
	wire [46-1:0] node1226;
	wire [46-1:0] node1230;
	wire [46-1:0] node1233;
	wire [46-1:0] node1234;
	wire [46-1:0] node1237;
	wire [46-1:0] node1238;
	wire [46-1:0] node1242;
	wire [46-1:0] node1243;
	wire [46-1:0] node1244;
	wire [46-1:0] node1245;
	wire [46-1:0] node1247;
	wire [46-1:0] node1249;
	wire [46-1:0] node1251;
	wire [46-1:0] node1253;
	wire [46-1:0] node1255;
	wire [46-1:0] node1257;
	wire [46-1:0] node1259;
	wire [46-1:0] node1262;
	wire [46-1:0] node1263;
	wire [46-1:0] node1265;
	wire [46-1:0] node1267;
	wire [46-1:0] node1268;
	wire [46-1:0] node1271;
	wire [46-1:0] node1273;
	wire [46-1:0] node1274;
	wire [46-1:0] node1277;
	wire [46-1:0] node1280;
	wire [46-1:0] node1281;
	wire [46-1:0] node1282;
	wire [46-1:0] node1283;
	wire [46-1:0] node1284;
	wire [46-1:0] node1287;
	wire [46-1:0] node1288;
	wire [46-1:0] node1289;
	wire [46-1:0] node1293;
	wire [46-1:0] node1296;
	wire [46-1:0] node1297;
	wire [46-1:0] node1299;
	wire [46-1:0] node1302;
	wire [46-1:0] node1305;
	wire [46-1:0] node1306;
	wire [46-1:0] node1307;
	wire [46-1:0] node1308;
	wire [46-1:0] node1309;
	wire [46-1:0] node1315;
	wire [46-1:0] node1317;
	wire [46-1:0] node1320;
	wire [46-1:0] node1321;
	wire [46-1:0] node1323;
	wire [46-1:0] node1324;
	wire [46-1:0] node1325;
	wire [46-1:0] node1328;
	wire [46-1:0] node1331;
	wire [46-1:0] node1333;
	wire [46-1:0] node1336;
	wire [46-1:0] node1337;
	wire [46-1:0] node1339;
	wire [46-1:0] node1343;
	wire [46-1:0] node1344;
	wire [46-1:0] node1345;
	wire [46-1:0] node1346;
	wire [46-1:0] node1347;
	wire [46-1:0] node1348;
	wire [46-1:0] node1349;
	wire [46-1:0] node1350;
	wire [46-1:0] node1352;
	wire [46-1:0] node1356;
	wire [46-1:0] node1359;
	wire [46-1:0] node1360;
	wire [46-1:0] node1362;
	wire [46-1:0] node1364;
	wire [46-1:0] node1367;
	wire [46-1:0] node1369;
	wire [46-1:0] node1371;
	wire [46-1:0] node1374;
	wire [46-1:0] node1375;
	wire [46-1:0] node1378;
	wire [46-1:0] node1379;
	wire [46-1:0] node1382;
	wire [46-1:0] node1383;
	wire [46-1:0] node1387;
	wire [46-1:0] node1388;
	wire [46-1:0] node1389;
	wire [46-1:0] node1391;
	wire [46-1:0] node1394;
	wire [46-1:0] node1395;
	wire [46-1:0] node1398;
	wire [46-1:0] node1399;
	wire [46-1:0] node1402;
	wire [46-1:0] node1405;
	wire [46-1:0] node1406;
	wire [46-1:0] node1407;
	wire [46-1:0] node1408;
	wire [46-1:0] node1409;
	wire [46-1:0] node1412;
	wire [46-1:0] node1415;
	wire [46-1:0] node1418;
	wire [46-1:0] node1420;
	wire [46-1:0] node1423;
	wire [46-1:0] node1426;
	wire [46-1:0] node1427;
	wire [46-1:0] node1428;
	wire [46-1:0] node1429;
	wire [46-1:0] node1430;
	wire [46-1:0] node1433;
	wire [46-1:0] node1436;
	wire [46-1:0] node1437;
	wire [46-1:0] node1439;
	wire [46-1:0] node1442;
	wire [46-1:0] node1444;
	wire [46-1:0] node1447;
	wire [46-1:0] node1448;
	wire [46-1:0] node1449;
	wire [46-1:0] node1450;
	wire [46-1:0] node1455;
	wire [46-1:0] node1458;
	wire [46-1:0] node1459;
	wire [46-1:0] node1460;
	wire [46-1:0] node1461;
	wire [46-1:0] node1465;
	wire [46-1:0] node1466;
	wire [46-1:0] node1469;
	wire [46-1:0] node1472;
	wire [46-1:0] node1473;
	wire [46-1:0] node1474;
	wire [46-1:0] node1476;
	wire [46-1:0] node1479;
	wire [46-1:0] node1480;
	wire [46-1:0] node1484;
	wire [46-1:0] node1486;
	wire [46-1:0] node1489;
	wire [46-1:0] node1490;
	wire [46-1:0] node1491;
	wire [46-1:0] node1492;
	wire [46-1:0] node1493;
	wire [46-1:0] node1494;
	wire [46-1:0] node1497;
	wire [46-1:0] node1499;
	wire [46-1:0] node1502;
	wire [46-1:0] node1504;
	wire [46-1:0] node1506;
	wire [46-1:0] node1509;
	wire [46-1:0] node1510;
	wire [46-1:0] node1512;
	wire [46-1:0] node1513;
	wire [46-1:0] node1515;
	wire [46-1:0] node1518;
	wire [46-1:0] node1521;
	wire [46-1:0] node1522;
	wire [46-1:0] node1525;
	wire [46-1:0] node1526;
	wire [46-1:0] node1530;
	wire [46-1:0] node1531;
	wire [46-1:0] node1532;
	wire [46-1:0] node1533;
	wire [46-1:0] node1536;
	wire [46-1:0] node1539;
	wire [46-1:0] node1540;
	wire [46-1:0] node1543;
	wire [46-1:0] node1546;
	wire [46-1:0] node1547;
	wire [46-1:0] node1548;
	wire [46-1:0] node1551;
	wire [46-1:0] node1554;
	wire [46-1:0] node1555;
	wire [46-1:0] node1559;
	wire [46-1:0] node1560;
	wire [46-1:0] node1561;
	wire [46-1:0] node1562;
	wire [46-1:0] node1563;
	wire [46-1:0] node1564;
	wire [46-1:0] node1568;
	wire [46-1:0] node1570;
	wire [46-1:0] node1573;
	wire [46-1:0] node1574;
	wire [46-1:0] node1577;
	wire [46-1:0] node1578;
	wire [46-1:0] node1581;
	wire [46-1:0] node1584;
	wire [46-1:0] node1585;
	wire [46-1:0] node1586;
	wire [46-1:0] node1588;
	wire [46-1:0] node1591;
	wire [46-1:0] node1594;
	wire [46-1:0] node1595;
	wire [46-1:0] node1597;
	wire [46-1:0] node1599;
	wire [46-1:0] node1603;
	wire [46-1:0] node1604;
	wire [46-1:0] node1605;
	wire [46-1:0] node1608;
	wire [46-1:0] node1609;
	wire [46-1:0] node1612;
	wire [46-1:0] node1615;
	wire [46-1:0] node1616;
	wire [46-1:0] node1617;
	wire [46-1:0] node1619;
	wire [46-1:0] node1620;
	wire [46-1:0] node1624;
	wire [46-1:0] node1627;
	wire [46-1:0] node1628;
	wire [46-1:0] node1631;
	wire [46-1:0] node1634;
	wire [46-1:0] node1635;
	wire [46-1:0] node1636;
	wire [46-1:0] node1637;
	wire [46-1:0] node1638;
	wire [46-1:0] node1639;
	wire [46-1:0] node1642;
	wire [46-1:0] node1647;
	wire [46-1:0] node1648;
	wire [46-1:0] node1649;
	wire [46-1:0] node1650;
	wire [46-1:0] node1653;
	wire [46-1:0] node1656;
	wire [46-1:0] node1657;
	wire [46-1:0] node1660;
	wire [46-1:0] node1663;
	wire [46-1:0] node1664;
	wire [46-1:0] node1665;
	wire [46-1:0] node1668;
	wire [46-1:0] node1672;
	wire [46-1:0] node1673;
	wire [46-1:0] node1674;
	wire [46-1:0] node1675;
	wire [46-1:0] node1676;
	wire [46-1:0] node1679;
	wire [46-1:0] node1682;
	wire [46-1:0] node1683;
	wire [46-1:0] node1686;
	wire [46-1:0] node1689;
	wire [46-1:0] node1690;
	wire [46-1:0] node1691;
	wire [46-1:0] node1694;
	wire [46-1:0] node1698;
	wire [46-1:0] node1699;
	wire [46-1:0] node1700;
	wire [46-1:0] node1701;
	wire [46-1:0] node1704;

	assign outp = (inp[1]) ? node210 : node1;
		assign node1 = (inp[3]) ? node5 : node2;
			assign node2 = (inp[15]) ? 46'b0000000000000000000000000000001000000000000000 : 46'b0000000000000000000000000000000000000000000000;
			assign node5 = (inp[15]) ? node43 : node6;
				assign node6 = (inp[0]) ? node24 : node7;
					assign node7 = (inp[12]) ? node9 : 46'b0000000000000000000000000000000000000000000000;
						assign node9 = (inp[7]) ? node11 : 46'b0000000000000000000000000000000000000000000000;
							assign node11 = (inp[13]) ? node13 : 46'b0000000000000000000000000000000000000000000000;
								assign node13 = (inp[11]) ? 46'b0000000000000000000000000000000000000000000000 : node14;
									assign node14 = (inp[6]) ? node16 : 46'b0000000000000000000000000000000000000000000000;
										assign node16 = (inp[5]) ? node18 : 46'b0000000000000000000000000000000000000000000000;
											assign node18 = (inp[2]) ? node20 : 46'b0000000000000000000000000000000000000000000000;
												assign node20 = (inp[9]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0000000000000000000000000000000000000100000000;
					assign node24 = (inp[7]) ? node26 : 46'b0000000000000000000000000000000000000000000000;
						assign node26 = (inp[11]) ? 46'b0000000000000000000000000000000000000000000000 : node27;
							assign node27 = (inp[10]) ? node29 : 46'b0000000000000000000000000000000000000000000000;
								assign node29 = (inp[4]) ? node31 : 46'b0000000000000000000000000000000000000000000000;
									assign node31 = (inp[12]) ? node33 : 46'b0000000000000000000000000000000000000000000000;
										assign node33 = (inp[13]) ? node35 : 46'b0000000000000000000000000000000000000000000000;
											assign node35 = (inp[8]) ? node37 : 46'b0000000000000000000000000000000000000000000000;
												assign node37 = (inp[14]) ? node39 : 46'b0000000000000000000000000000000000000000000000;
													assign node39 = (inp[6]) ? 46'b0000000001000000000000000000001000000000000000 : 46'b0000000000000000000000000000000000000000000000;
				assign node43 = (inp[9]) ? node93 : node44;
					assign node44 = (inp[11]) ? node80 : node45;
						assign node45 = (inp[13]) ? node51 : node46;
							assign node46 = (inp[2]) ? 46'b0000000000000000000000000000000000000000000000 : node47;
								assign node47 = (inp[0]) ? 46'b0000000000001000000000000010000000000000000000 : 46'b0000001000001000000000000000000000000000000000;
							assign node51 = (inp[6]) ? node53 : 46'b0000000000000000000000000000000000000000000000;
								assign node53 = (inp[14]) ? node55 : 46'b0000000000000000000000000000000000000000000000;
									assign node55 = (inp[5]) ? node57 : 46'b0000000000000000000000000000000000000000000000;
										assign node57 = (inp[8]) ? node59 : 46'b0000000000000000000000000000000000000000000000;
											assign node59 = (inp[0]) ? 46'b0000000000000000000000000000000000000000000000 : node60;
												assign node60 = (inp[2]) ? node70 : node61;
													assign node61 = (inp[4]) ? node65 : node62;
														assign node62 = (inp[10]) ? 46'b0000000000001000010100010000000000000000010000 : 46'b0000000000000000000000000000000000000000000000;
														assign node65 = (inp[12]) ? node67 : 46'b0000000000000000000000000000000000000000000000;
															assign node67 = (inp[7]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0000010000000000010100000000000100000000010000;
													assign node70 = (inp[7]) ? 46'b0000000000000000000000000000000000000000000000 : node71;
														assign node71 = (inp[12]) ? node73 : 46'b0000000000000000000000000000000000000000000000;
															assign node73 = (inp[4]) ? 46'b0000010000000000010000000000000101000010000000 : node74;
																assign node74 = (inp[10]) ? 46'b0000010000000000010000010000000001000010000000 : 46'b0000000000000000000000000000000000000000000000;
						assign node80 = (inp[13]) ? node86 : node81;
							assign node81 = (inp[2]) ? 46'b0000000000000000000000000000000000000000000000 : node82;
								assign node82 = (inp[0]) ? 46'b0000010000000000000000000010000000000000000000 : 46'b0000011000000000000000000000000000000000000000;
							assign node86 = (inp[2]) ? node90 : node87;
								assign node87 = (inp[0]) ? 46'b0000001000000000011000000100000000000000010000 : 46'b0000001000000000010000000100000000000000010010;
								assign node90 = (inp[0]) ? 46'b0000001000000000010010000000010000000010000000 : 46'b0000001000000000010010100000000000000010000000;
					assign node93 = (inp[0]) ? node145 : node94;
						assign node94 = (inp[13]) ? node100 : node95;
							assign node95 = (inp[2]) ? 46'b0000000000000000000000000000000000000000000000 : node96;
								assign node96 = (inp[11]) ? 46'b0000010100000000000000000000000000000000000000 : 46'b0000000100001000000000000000000000000000000000;
							assign node100 = (inp[5]) ? node102 : 46'b0000000000000000000000000000000000000000000000;
								assign node102 = (inp[14]) ? node104 : 46'b0000000000000000000000000000000000000000000000;
									assign node104 = (inp[6]) ? node106 : 46'b0000000000000000000000000000000000000000000000;
										assign node106 = (inp[10]) ? node122 : node107;
											assign node107 = (inp[4]) ? node109 : 46'b0000000000000000000000000000000000000000000000;
												assign node109 = (inp[8]) ? node111 : 46'b0000000000000000000000000000000000000000000000;
													assign node111 = (inp[7]) ? node119 : node112;
														assign node112 = (inp[12]) ? node116 : node113;
															assign node113 = (inp[2]) ? 46'b0010000000000000000000000000000100000010000000 : 46'b0010000000000000000000000000000100000000010000;
															assign node116 = (inp[2]) ? 46'b0000010000000000010000000000000100000010000000 : 46'b0000010000000000010000000000000100000000010000;
														assign node119 = (inp[12]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0000000000001000010000000000000100000010000000;
											assign node122 = (inp[2]) ? node136 : node123;
												assign node123 = (inp[12]) ? node133 : node124;
													assign node124 = (inp[11]) ? node130 : node125;
														assign node125 = (inp[7]) ? 46'b0000000000000000000000000000000000000000000000 : node126;
															assign node126 = (inp[8]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0010000000010000000000000000000000000000010000;
														assign node130 = (inp[4]) ? 46'b0000000000011000010000000100000000000000010010 : 46'b0000000000000000000000000000000000000000000000;
													assign node133 = (inp[11]) ? 46'b0000010000000000010000010100000000000000010010 : 46'b0000010000000000010000010000000000000000010000;
												assign node136 = (inp[4]) ? node138 : 46'b0000000000000000000000000000000000000000000000;
													assign node138 = (inp[11]) ? 46'b0000010000010000010010100000000000000010000000 : node139;
														assign node139 = (inp[12]) ? 46'b0000000000000000000000000000000000000000000000 : node140;
															assign node140 = (inp[7]) ? 46'b0000000000011000010000000000000000000010000000 : 46'b0010000000010000000000000000000000000010000000;
						assign node145 = (inp[11]) ? node175 : node146;
							assign node146 = (inp[13]) ? node150 : node147;
								assign node147 = (inp[2]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0010001000000000000000000000000000000000010000;
								assign node150 = (inp[6]) ? node152 : 46'b0000000000000000000000000000000000000000000000;
									assign node152 = (inp[14]) ? node154 : 46'b0000000000000000000000000000000000000000000000;
										assign node154 = (inp[2]) ? 46'b0000000000000000000000000000000000000000000000 : node155;
											assign node155 = (inp[5]) ? node157 : 46'b0000000000000000000000000000000000000000000000;
												assign node157 = (inp[12]) ? node167 : node158;
													assign node158 = (inp[10]) ? node162 : node159;
														assign node159 = (inp[4]) ? 46'b0000000000001000010000000000000100000000010100 : 46'b0000000000000000000000000000000000000000000000;
														assign node162 = (inp[7]) ? 46'b0000000000000000000000000000000000000000000000 : node163;
															assign node163 = (inp[8]) ? 46'b0010000000000000000000010000000000000000010100 : 46'b0010000000010000000000000000000000000000010100;
													assign node167 = (inp[4]) ? node169 : 46'b0000000000000000000000000000000000000000000000;
														assign node169 = (inp[10]) ? node171 : 46'b0000000000000000000000000000000000000000000000;
															assign node171 = (inp[8]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0000010000010000010000000000000000000000010100;
							assign node175 = (inp[14]) ? node177 : 46'b0000000000000000000000000000000000000000000000;
								assign node177 = (inp[5]) ? node179 : 46'b0000000000000000000000000000000000000000000000;
									assign node179 = (inp[6]) ? node189 : node180;
										assign node180 = (inp[10]) ? node182 : 46'b0000000000000000000000000000000000000000000000;
											assign node182 = (inp[12]) ? node184 : 46'b0000000000000000000000000000000000000000000000;
												assign node184 = (inp[7]) ? 46'b0000000000000000000000000000000000000000000000 : node185;
													assign node185 = (inp[8]) ? 46'b0000000000000000000110000000010000000000000000 : 46'b0000000000000000000000000000000000000000000000;
										assign node189 = (inp[13]) ? node191 : 46'b0000000000000000000000000000000000000000000000;
											assign node191 = (inp[10]) ? node197 : node192;
												assign node192 = (inp[4]) ? node194 : 46'b0000000000000000000000000000000000000000000000;
													assign node194 = (inp[8]) ? 46'b0000010000000000011000000100000100000000010000 : 46'b0000000000000000000000000000000000000000000000;
												assign node197 = (inp[2]) ? node205 : node198;
													assign node198 = (inp[4]) ? node202 : node199;
														assign node199 = (inp[12]) ? 46'b0000010000000000011000010100000000000000010000 : 46'b0010000000000000001000010100000000000000010000;
														assign node202 = (inp[12]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0000000000011000011000000100000000000000010000;
													assign node205 = (inp[4]) ? 46'b0000000000000000000000000000000000000000000000 : node206;
														assign node206 = (inp[8]) ? 46'b0000010000000000010010010000010000000010000000 : 46'b0000000000000000000000000000000000000000000000;
		assign node210 = (inp[15]) ? node278 : node211;
			assign node211 = (inp[13]) ? node215 : node212;
				assign node212 = (inp[3]) ? 46'b0000100000000000000000000000001000000000000000 : 46'b0000100000000000000000000000000000000000000000;
				assign node215 = (inp[2]) ? node247 : node216;
					assign node216 = (inp[11]) ? node232 : node217;
						assign node217 = (inp[0]) ? node225 : node218;
							assign node218 = (inp[9]) ? node222 : node219;
								assign node219 = (inp[3]) ? 46'b0000100000001000010000010100001000000000010010 : 46'b0000100000001000010000010100000000000000010010;
								assign node222 = (inp[3]) ? 46'b0000110000000000010000010100001000000000010010 : 46'b0000110000000000010000010100000000000000010010;
							assign node225 = (inp[9]) ? node229 : node226;
								assign node226 = (inp[3]) ? 46'b0000100000001000010000000100001100000000010010 : 46'b0000100000001000010000000100000100000000010010;
								assign node229 = (inp[3]) ? 46'b0000110000000000010000000100001100000000010010 : 46'b0000110000000000010000000100000100000000010010;
						assign node232 = (inp[9]) ? node240 : node233;
							assign node233 = (inp[0]) ? node237 : node234;
								assign node234 = (inp[3]) ? 46'b0000100000001000011000010100001000000000010000 : 46'b0000100000001000011000010100000000000000010000;
								assign node237 = (inp[3]) ? 46'b0000100000001000011000000100001100000000010000 : 46'b0000100000001000011000000100000100000000010000;
							assign node240 = (inp[0]) ? node244 : node241;
								assign node241 = (inp[3]) ? 46'b0000110000000000011000010100001000000000010000 : 46'b0000110000000000011000010100000000000000010000;
								assign node244 = (inp[3]) ? 46'b0000110000000000011000000100001100000000010000 : 46'b0000110000000000011000000100000100000000010000;
					assign node247 = (inp[0]) ? node263 : node248;
						assign node248 = (inp[11]) ? node256 : node249;
							assign node249 = (inp[9]) ? node253 : node250;
								assign node250 = (inp[3]) ? 46'b0000100000001000010010110000001000000010000000 : 46'b0000100000001000010010110000000000000010000000;
								assign node253 = (inp[3]) ? 46'b0000110000000000010010110000001000000010000000 : 46'b0000110000000000010010110000000000000010000000;
							assign node256 = (inp[9]) ? node260 : node257;
								assign node257 = (inp[3]) ? 46'b0000100000001000010010010000011000000010000000 : 46'b0000100000001000010010010000010000000010000000;
								assign node260 = (inp[3]) ? 46'b0000110000000000010010010000011000000010000000 : 46'b0000110000000000010010010000010000000010000000;
						assign node263 = (inp[11]) ? node271 : node264;
							assign node264 = (inp[9]) ? node268 : node265;
								assign node265 = (inp[3]) ? 46'b0000100000001000010010100000001100000010000000 : 46'b0000100000001000010010100000000100000010000000;
								assign node268 = (inp[3]) ? 46'b0000110000000000010010100000001100000010000000 : 46'b0000110000000000010010100000000100000010000000;
							assign node271 = (inp[9]) ? node275 : node272;
								assign node272 = (inp[3]) ? 46'b0000100000001000010010000000011100000010000000 : 46'b0000100000001000010010000000010100000010000000;
								assign node275 = (inp[3]) ? 46'b0000110000000000010010000000011100000010000000 : 46'b0000110000000000010010000000010100000010000000;
			assign node278 = (inp[3]) ? node282 : node279;
				assign node279 = (inp[13]) ? 46'b0000000000000000000000000000001000000000000000 : 46'b0000000000000000000000000000001000000000001000;
				assign node282 = (inp[13]) ? node284 : 46'b0000000000000000000000000000000000000000001000;
					assign node284 = (inp[2]) ? node1242 : node285;
						assign node285 = (inp[11]) ? node695 : node286;
							assign node286 = (inp[9]) ? node628 : node287;
								assign node287 = (inp[0]) ? node457 : node288;
									assign node288 = (inp[7]) ? node376 : node289;
										assign node289 = (inp[5]) ? node335 : node290;
											assign node290 = (inp[14]) ? node316 : node291;
												assign node291 = (inp[8]) ? node303 : node292;
													assign node292 = (inp[12]) ? node294 : 46'b0011000000000100001000010001100010010001010000;
														assign node294 = (inp[6]) ? node296 : 46'b0011000000000100000000010000100000110001010000;
															assign node296 = (inp[10]) ? node300 : node297;
																assign node297 = (inp[4]) ? 46'b0011000000000100001000010001100000010001010000 : 46'b0011000000000100000000010000100000010001010000;
																assign node300 = (inp[4]) ? 46'b0011000000000110000000010000100000010001010000 : 46'b0011000000000100000000010001100000010001010010;
													assign node303 = (inp[4]) ? node311 : node304;
														assign node304 = (inp[12]) ? node306 : 46'b0011000000000100000000010001100010110001010010;
															assign node306 = (inp[6]) ? 46'b0011000000000100000000010001100000010001010010 : node307;
																assign node307 = (inp[10]) ? 46'b0011000000000000000000010001100000110001010010 : 46'b0011000000000100000000010001100000110001010010;
														assign node311 = (inp[6]) ? node313 : 46'b0011000000000000001000010001100000110001010010;
															assign node313 = (inp[12]) ? 46'b0011000000000000001000010001100000010001010010 : 46'b0011000000000000001000010001100010010001010010;
												assign node316 = (inp[8]) ? node320 : node317;
													assign node317 = (inp[10]) ? 46'b0011000000000000001000010001100000110001010010 : 46'b0011000000000000001000010001100010010001010000;
													assign node320 = (inp[4]) ? node324 : node321;
														assign node321 = (inp[6]) ? 46'b0011000000000110000000010000100010010001010000 : 46'b0011000000000110000000010000100010110001010000;
														assign node324 = (inp[10]) ? node330 : node325;
															assign node325 = (inp[12]) ? node327 : 46'b0011000000000010001000010001100010110001010000;
																assign node327 = (inp[6]) ? 46'b0011000000000010001000010001100000010001010000 : 46'b0011000000000010001000010001100000110001010000;
															assign node330 = (inp[6]) ? node332 : 46'b0011000000000010000000010000100000110001010000;
																assign node332 = (inp[12]) ? 46'b0011000000000010000000010000100000010001010000 : 46'b0011000000000010000000010000100010010001010000;
											assign node335 = (inp[6]) ? node355 : node336;
												assign node336 = (inp[14]) ? node342 : node337;
													assign node337 = (inp[12]) ? node339 : 46'b0010000000000000000000010001100010110001010010;
														assign node339 = (inp[4]) ? 46'b0010000000000010000000010001100000110001010010 : 46'b0010000000000000000000010001100000110001010010;
													assign node342 = (inp[12]) ? node350 : node343;
														assign node343 = (inp[4]) ? node347 : node344;
															assign node344 = (inp[10]) ? 46'b0010000000000010000000010001100010110001010010 : 46'b0010000000000110000000010000100010110001010000;
															assign node347 = (inp[10]) ? 46'b0010000000000010000000010000100010110001010000 : 46'b0010000000000010001000010001100010110001010000;
														assign node350 = (inp[10]) ? 46'b0010000000000010000000010000100000110001010000 : node351;
															assign node351 = (inp[8]) ? 46'b0010000000000010001000010001100000110001010000 : 46'b0010000000000000001000010001100000110001010000;
												assign node355 = (inp[12]) ? node367 : node356;
													assign node356 = (inp[14]) ? node362 : node357;
														assign node357 = (inp[8]) ? node359 : 46'b0010000000000110000000010000100010010001010000;
															assign node359 = (inp[4]) ? 46'b0010000000000010000000010001100010010001010010 : 46'b0010000000000100000000010001100010010001010010;
														assign node362 = (inp[10]) ? 46'b0010000000000000001000010001100010010001010010 : node363;
															assign node363 = (inp[4]) ? 46'b0010000000000010001000010001100010010001010000 : 46'b0010000000000110000000010000100010010001010000;
													assign node367 = (inp[10]) ? node371 : node368;
														assign node368 = (inp[8]) ? 46'b0010000000000110000000010000100000010001010000 : 46'b0010000000000100001000010001100000010001010000;
														assign node371 = (inp[8]) ? 46'b0010000000000010000000010001100000010001010010 : node372;
															assign node372 = (inp[4]) ? 46'b0010000000000010001000010001100000010001010000 : 46'b0010000000000000001000010001100000010001010010;
										assign node376 = (inp[12]) ? node414 : node377;
											assign node377 = (inp[6]) ? node395 : node378;
												assign node378 = (inp[5]) ? node388 : node379;
													assign node379 = (inp[8]) ? node383 : node380;
														assign node380 = (inp[10]) ? 46'b0011000000000000001000010001000010110001010010 : 46'b0011000000000100001000010001000010110001010000;
														assign node383 = (inp[14]) ? node385 : 46'b0011000000000000001000010001000010110001010010;
															assign node385 = (inp[4]) ? 46'b0011000000000010001000010001000010110001010000 : 46'b0011000000000010000000010001000010110001010010;
													assign node388 = (inp[14]) ? node392 : node389;
														assign node389 = (inp[10]) ? 46'b0010000000000100000000010001000010110001010010 : 46'b0010000000000000001000010001000010110001010010;
														assign node392 = (inp[4]) ? 46'b0010000000000010001000010001000010110001010000 : 46'b0010000000000000001000010001000010110001010010;
												assign node395 = (inp[5]) ? node405 : node396;
													assign node396 = (inp[8]) ? 46'b0011000000000100000000010001000010010001010010 : node397;
														assign node397 = (inp[10]) ? 46'b0011000000000000001000010001000010010001010010 : node398;
															assign node398 = (inp[4]) ? node400 : 46'b0011000000000100001000010001000010010001010000;
																assign node400 = (inp[14]) ? 46'b0011000000000000001000010001000010010001010000 : 46'b0011000000000100001000010001000010010001010000;
													assign node405 = (inp[8]) ? node409 : node406;
														assign node406 = (inp[10]) ? 46'b0010000000000100000000010001000010010001010010 : 46'b0010000000000100000000010000000010010001010000;
														assign node409 = (inp[10]) ? 46'b0010000000000010000000010001000010010001010010 : node410;
															assign node410 = (inp[14]) ? 46'b0010000000000010001000010001000010010001010000 : 46'b0010000000000000001000010001000010010001010010;
											assign node414 = (inp[6]) ? node434 : node415;
												assign node415 = (inp[5]) ? node429 : node416;
													assign node416 = (inp[10]) ? node422 : node417;
														assign node417 = (inp[4]) ? node419 : 46'b0011000000000100001000010001000000110001010000;
															assign node419 = (inp[8]) ? 46'b0011000000000000001000010001000000110001010010 : 46'b0011000000000000001000010001000000110001010000;
														assign node422 = (inp[4]) ? node424 : 46'b0011000000000010000000010001000000110001010010;
															assign node424 = (inp[14]) ? node426 : 46'b0011000000000110000000010000000000110001010000;
																assign node426 = (inp[8]) ? 46'b0011000000000010000000010000000000110001010000 : 46'b0011000000000010001000010001000000110001010000;
													assign node429 = (inp[10]) ? 46'b0010000000000010000000010001000000110001010010 : node430;
														assign node430 = (inp[14]) ? 46'b0010000000000110000000010000000000110001010000 : 46'b0010000000000100000000010000000000110001010000;
												assign node434 = (inp[5]) ? node446 : node435;
													assign node435 = (inp[8]) ? node441 : node436;
														assign node436 = (inp[14]) ? 46'b0011000000000010001000010001000000010001010000 : node437;
															assign node437 = (inp[10]) ? 46'b0011000000000110000000010000000000010001010000 : 46'b0011000000000100000000010000000000010001010000;
														assign node441 = (inp[10]) ? 46'b0011000000000010000000010001000000010001010010 : node442;
															assign node442 = (inp[4]) ? 46'b0011000000000000001000010001000000010001010010 : 46'b0011000000000100000000010001000000010001010010;
													assign node446 = (inp[14]) ? node452 : node447;
														assign node447 = (inp[10]) ? node449 : 46'b0010000000000000001000010001000000010001010010;
															assign node449 = (inp[4]) ? 46'b0010000000000010000000010001000000010001010010 : 46'b0010000000000000000000010001000000010001010010;
														assign node452 = (inp[4]) ? 46'b0010000000000010001000010001000000010001010000 : node453;
															assign node453 = (inp[10]) ? 46'b0010000000000000001000010001000000010001010010 : 46'b0010000000000100001000010001000000010001010000;
									assign node457 = (inp[5]) ? node541 : node458;
										assign node458 = (inp[6]) ? node498 : node459;
											assign node459 = (inp[12]) ? node481 : node460;
												assign node460 = (inp[7]) ? node470 : node461;
													assign node461 = (inp[10]) ? node467 : node462;
														assign node462 = (inp[8]) ? 46'b0011000000000010001000010001100010110000010000 : node463;
															assign node463 = (inp[4]) ? 46'b0011000000000000001000010001100010110000010000 : 46'b0011000000000100001000010001100010110000010000;
														assign node467 = (inp[14]) ? 46'b0011000000000010000000010000100010110000010000 : 46'b0011000000000010000000010001100010110000010010;
													assign node470 = (inp[10]) ? node474 : node471;
														assign node471 = (inp[8]) ? 46'b0011000000000110000000010000000010110000010000 : 46'b0011000000000100000000010000000010110000010000;
														assign node474 = (inp[4]) ? 46'b0011000000000010001000010001000010110000010000 : node475;
															assign node475 = (inp[14]) ? 46'b0011000000000010000000010001000010110000010010 : node476;
																assign node476 = (inp[8]) ? 46'b0011000000000000000000010001000010110000010010 : 46'b0011000000000100000000010001000010110000010010;
												assign node481 = (inp[8]) ? node493 : node482;
													assign node482 = (inp[14]) ? node486 : node483;
														assign node483 = (inp[10]) ? 46'b0011000000000110000000010000100000110000010000 : 46'b0011000000000100001000010001100000110000010000;
														assign node486 = (inp[4]) ? node490 : node487;
															assign node487 = (inp[7]) ? 46'b0011000000000100001000010001000000110000010000 : 46'b0011000000000000001000010001100000110000010010;
															assign node490 = (inp[7]) ? 46'b0011000000000010001000010001000000110000010000 : 46'b0011000000000010001000010001100000110000010000;
													assign node493 = (inp[10]) ? node495 : 46'b0011000000000110000000010000100000110000010000;
														assign node495 = (inp[7]) ? 46'b0011000000000010000000010000000000110000010000 : 46'b0011000000000010000000010001100000110000010010;
											assign node498 = (inp[7]) ? node520 : node499;
												assign node499 = (inp[14]) ? node511 : node500;
													assign node500 = (inp[4]) ? node506 : node501;
														assign node501 = (inp[12]) ? node503 : 46'b0011000000000100000000010001100010010000010010;
															assign node503 = (inp[8]) ? 46'b0011000000000100000000010001100000010000010010 : 46'b0011000000000100000000010000100000010000010000;
														assign node506 = (inp[8]) ? 46'b0011000000000000001000010001100000010000010010 : node507;
															assign node507 = (inp[12]) ? 46'b0011000000000100001000010001100000010000010000 : 46'b0011000000000100001000010001100010010000010000;
													assign node511 = (inp[12]) ? node515 : node512;
														assign node512 = (inp[4]) ? 46'b0011000000000010001000010001100010010000010000 : 46'b0011000000000110000000010000100010010000010000;
														assign node515 = (inp[10]) ? node517 : 46'b0011000000000110000000010000100000010000010000;
															assign node517 = (inp[4]) ? 46'b0011000000000010000000010000100000010000010000 : 46'b0011000000000010000000010001100000010000010010;
												assign node520 = (inp[14]) ? node528 : node521;
													assign node521 = (inp[8]) ? 46'b0011000000000000001000010001000000010000010010 : node522;
														assign node522 = (inp[4]) ? 46'b0011000000000110000000010000000000010000010000 : node523;
															assign node523 = (inp[10]) ? 46'b0011000000000100000000010001000000010000010010 : 46'b0011000000000100000000010000000000010000010000;
													assign node528 = (inp[8]) ? node534 : node529;
														assign node529 = (inp[10]) ? 46'b0011000000000010001000010001000000010000010000 : node530;
															assign node530 = (inp[12]) ? 46'b0011000000000000001000010001000000010000010000 : 46'b0011000000000000001000010001000010010000010000;
														assign node534 = (inp[12]) ? 46'b0011000000000010000000010000000000010000010000 : node535;
															assign node535 = (inp[10]) ? 46'b0011000000000010000000010001000010010000010010 : node536;
																assign node536 = (inp[4]) ? 46'b0011000000000010001000010001000010010000010000 : 46'b0011000000000110000000010000000010010000010000;
										assign node541 = (inp[7]) ? node583 : node542;
											assign node542 = (inp[6]) ? node566 : node543;
												assign node543 = (inp[12]) ? node555 : node544;
													assign node544 = (inp[4]) ? node548 : node545;
														assign node545 = (inp[10]) ? 46'b0010000000000100000000010001100010110000010010 : 46'b0010000000000100000000010000100010110000010000;
														assign node548 = (inp[10]) ? node552 : node549;
															assign node549 = (inp[8]) ? 46'b0010000000000010001000010001100010110000010000 : 46'b0010000000000000001000010001100010110000010000;
															assign node552 = (inp[14]) ? 46'b0010000000000010000000010000100010110000010000 : 46'b0010000000000010000000010001100010110000010010;
													assign node555 = (inp[10]) ? node557 : 46'b0010000000000110000000010000100000110000010000;
														assign node557 = (inp[4]) ? node561 : node558;
															assign node558 = (inp[8]) ? 46'b0010000000000010000000010001100000110000010010 : 46'b0010000000000000001000010001100000110000010010;
															assign node561 = (inp[8]) ? node563 : 46'b0010000000000110000000010000100000110000010000;
																assign node563 = (inp[14]) ? 46'b0010000000000010000000010000100000110000010000 : 46'b0010000000000010000000010001100000110000010010;
												assign node566 = (inp[12]) ? node578 : node567;
													assign node567 = (inp[10]) ? node571 : node568;
														assign node568 = (inp[4]) ? 46'b0010000000000010001000010001100010010000010000 : 46'b0010000000000110000000010000100010010000010000;
														assign node571 = (inp[8]) ? node573 : 46'b0010000000000100000000010001100010010000010010;
															assign node573 = (inp[14]) ? 46'b0010000000000010000000010001100010010000010010 : node574;
																assign node574 = (inp[4]) ? 46'b0010000000000010000000010001100010010000010010 : 46'b0010000000000000000000010001100010010000010010;
													assign node578 = (inp[8]) ? node580 : 46'b0010000000000110000000010000100000010000010000;
														assign node580 = (inp[4]) ? 46'b0010000000000000001000010001100000010000010010 : 46'b0010000000000000000000010001100000010000010010;
											assign node583 = (inp[6]) ? node607 : node584;
												assign node584 = (inp[10]) ? node598 : node585;
													assign node585 = (inp[12]) ? node595 : node586;
														assign node586 = (inp[8]) ? node592 : node587;
															assign node587 = (inp[4]) ? 46'b0010000000000100001000010001000010110000010000 : node588;
																assign node588 = (inp[14]) ? 46'b0010000000000100001000010001000010110000010000 : 46'b0010000000000100000000010000000010110000010000;
															assign node592 = (inp[14]) ? 46'b0010000000000110000000010000000010110000010000 : 46'b0010000000000100000000010001000010110000010010;
														assign node595 = (inp[14]) ? 46'b0010000000000000001000010001000000110000010000 : 46'b0010000000000100000000010001000000110000010010;
													assign node598 = (inp[4]) ? node602 : node599;
														assign node599 = (inp[12]) ? 46'b0010000000000000000000010001000000110000010010 : 46'b0010000000000010000000010001000010110000010010;
														assign node602 = (inp[8]) ? node604 : 46'b0010000000000010001000010001000010110000010000;
															assign node604 = (inp[12]) ? 46'b0010000000000010000000010000000000110000010000 : 46'b0010000000000010000000010000000010110000010000;
												assign node607 = (inp[12]) ? node617 : node608;
													assign node608 = (inp[8]) ? node612 : node609;
														assign node609 = (inp[10]) ? 46'b0010000000000100000000010001000010010000010010 : 46'b0010000000000100000000010000000010010000010000;
														assign node612 = (inp[14]) ? 46'b0010000000000010001000010001000010010000010000 : node613;
															assign node613 = (inp[10]) ? 46'b0010000000000010000000010001000010010000010010 : 46'b0010000000000000001000010001000010010000010010;
													assign node617 = (inp[10]) ? node623 : node618;
														assign node618 = (inp[4]) ? 46'b0010000000000100001000010001000000010000010000 : node619;
															assign node619 = (inp[14]) ? 46'b0010000000000110000000010000000000010000010000 : 46'b0010000000000100000000010000000000010000010000;
														assign node623 = (inp[4]) ? 46'b0010000000000110000000010000000000010000010000 : node624;
															assign node624 = (inp[8]) ? 46'b0010000000000010000000010001000000010000010010 : 46'b0010000000000100000000010001000000010000010010;
								assign node628 = (inp[0]) ? 46'b0000000000000000000000000000000000000000000000 : node629;
									assign node629 = (inp[5]) ? node663 : node630;
										assign node630 = (inp[7]) ? node632 : 46'b0000000000000000000000000000000000000000000000;
											assign node632 = (inp[8]) ? node654 : node633;
												assign node633 = (inp[12]) ? node645 : node634;
													assign node634 = (inp[6]) ? node638 : node635;
														assign node635 = (inp[14]) ? 46'b0001000000000100001000001001000010100000000000 : 46'b0001000000000100000000001001000010100000000010;
														assign node638 = (inp[10]) ? 46'b0001000000000110000000001000000010000000000000 : node639;
															assign node639 = (inp[4]) ? 46'b0001000000000100001000001001000010000000000000 : node640;
																assign node640 = (inp[14]) ? 46'b0001000000000100001000001001000010000000000000 : 46'b0001000000000100000000001000000010000000000000;
													assign node645 = (inp[10]) ? node651 : node646;
														assign node646 = (inp[14]) ? 46'b0001000000000100001000001001000000100000000000 : node647;
															assign node647 = (inp[4]) ? 46'b0001000000000100001000001001000000100000000000 : 46'b0001000000000100000000001000000000100000000000;
														assign node651 = (inp[14]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0001000000000110000000001000000000100000000000;
												assign node654 = (inp[4]) ? 46'b0000000000000000000000000000000000000000000000 : node655;
													assign node655 = (inp[10]) ? 46'b0000000000000000000000000000000000000000000000 : node656;
														assign node656 = (inp[14]) ? node658 : 46'b0001000000000100000000001001000010100000000010;
															assign node658 = (inp[12]) ? 46'b0001000000000110000000001000000000100000000000 : 46'b0001000000000110000000001000000010100000000000;
										assign node663 = (inp[7]) ? 46'b0000000000000000000000000000000000000000000000 : node664;
											assign node664 = (inp[10]) ? node670 : node665;
												assign node665 = (inp[8]) ? node667 : 46'b0000000000000000000000000000000000000000000000;
													assign node667 = (inp[14]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0000000000000000001000001001100000100000000010;
												assign node670 = (inp[4]) ? node682 : node671;
													assign node671 = (inp[14]) ? node677 : node672;
														assign node672 = (inp[8]) ? 46'b0000000000000000000000001001100010000000000010 : node673;
															assign node673 = (inp[12]) ? 46'b0000000000000100000000001001100000000000000010 : 46'b0000000000000100000000001001100010000000000010;
														assign node677 = (inp[8]) ? node679 : 46'b0000000000000000001000001001100000000000000010;
															assign node679 = (inp[6]) ? 46'b0000000000000010000000001001100000000000000010 : 46'b0000000000000010000000001001100000100000000010;
													assign node682 = (inp[14]) ? 46'b0000000000000000000000000000000000000000000000 : node683;
														assign node683 = (inp[8]) ? node685 : 46'b0000000000000000000000000000000000000000000000;
															assign node685 = (inp[6]) ? node689 : node686;
																assign node686 = (inp[12]) ? 46'b0000000000000010000000001001100000100000000010 : 46'b0000000000000010000000001001100010100000000010;
																assign node689 = (inp[12]) ? 46'b0000000000000010000000001001100000000000000010 : 46'b0000000000000010000000001001100010000000000010;
							assign node695 = (inp[0]) ? node895 : node696;
								assign node696 = (inp[9]) ? node730 : node697;
									assign node697 = (inp[7]) ? node699 : 46'b0000000000000000000000000000000000000000000000;
										assign node699 = (inp[5]) ? node701 : 46'b0000000000000000000000000000000000000000000000;
											assign node701 = (inp[12]) ? node723 : node702;
												assign node702 = (inp[6]) ? node704 : 46'b0000000000000000000000000000000000000000000000;
													assign node704 = (inp[4]) ? node712 : node705;
														assign node705 = (inp[14]) ? 46'b0000000000000110000001000000000010000000000000 : node706;
															assign node706 = (inp[10]) ? node708 : 46'b0000000000000100000001000001000010000000000010;
																assign node708 = (inp[8]) ? 46'b0000000000000000000001000001000010000000000010 : 46'b0000000000000100000001000001000010000000000010;
														assign node712 = (inp[10]) ? node718 : node713;
															assign node713 = (inp[8]) ? 46'b0000000000000000001001000001000010000000000010 : node714;
																assign node714 = (inp[14]) ? 46'b0000000000000000001001000001000010000000000000 : 46'b0000000000000100001001000001000010000000000000;
															assign node718 = (inp[8]) ? 46'b0000000000000010000001000001000010000000000010 : node719;
																assign node719 = (inp[14]) ? 46'b0000000000000010001001000001000010000000000000 : 46'b0000000000000110000001000000000010000000000000;
												assign node723 = (inp[6]) ? 46'b0000000000000000000000000000000000000000000000 : node724;
													assign node724 = (inp[10]) ? 46'b0000000000000100000001000001000000100000000010 : node725;
														assign node725 = (inp[8]) ? 46'b0000000000000100000001000001000000100000000010 : 46'b0000000000000100001001000001000000100000000000;
									assign node730 = (inp[7]) ? node822 : node731;
										assign node731 = (inp[12]) ? node775 : node732;
											assign node732 = (inp[5]) ? node754 : node733;
												assign node733 = (inp[8]) ? node745 : node734;
													assign node734 = (inp[10]) ? node742 : node735;
														assign node735 = (inp[6]) ? 46'b1001000000000100001000000001100010000000000000 : node736;
															assign node736 = (inp[14]) ? 46'b1001000000000100001000000001100010100000000000 : node737;
																assign node737 = (inp[4]) ? 46'b1001000000000100001000000001100010100000000000 : 46'b1001000000000100000000000000100010100000000000;
														assign node742 = (inp[14]) ? 46'b1001000000000010001000000001100010000000000000 : 46'b1001000000000110000000000000100010000000000000;
													assign node745 = (inp[4]) ? node751 : node746;
														assign node746 = (inp[6]) ? node748 : 46'b1001000000000000000000000001100010100000000010;
															assign node748 = (inp[10]) ? 46'b1001000000000000000000000001100010000000000010 : 46'b1001000000000100000000000001100010000000000010;
														assign node751 = (inp[14]) ? 46'b1001000000000010001000000001100010100000000000 : 46'b1001000000000000001000000001100010100000000010;
												assign node754 = (inp[14]) ? node762 : node755;
													assign node755 = (inp[4]) ? node759 : node756;
														assign node756 = (inp[6]) ? 46'b1000000000000100000000000000100010000000000000 : 46'b1000000000000100000000000000100010100000000000;
														assign node759 = (inp[10]) ? 46'b1000000000000110000000000000100010000000000000 : 46'b1000000000000100001000000001100010000000000000;
													assign node762 = (inp[8]) ? node770 : node763;
														assign node763 = (inp[10]) ? node767 : node764;
															assign node764 = (inp[4]) ? 46'b1000000000000000001000000001100010100000000000 : 46'b1000000000000100001000000001100010100000000000;
															assign node767 = (inp[6]) ? 46'b1000000000000000001000000001100010000000000010 : 46'b1000000000000000001000000001100010100000000010;
														assign node770 = (inp[6]) ? 46'b1000000000000010001000000001100010000000000000 : node771;
															assign node771 = (inp[10]) ? 46'b1000000000000010000000000001100010100000000010 : 46'b1000000000000110000000000000100010100000000000;
											assign node775 = (inp[6]) ? node793 : node776;
												assign node776 = (inp[5]) ? node782 : node777;
													assign node777 = (inp[4]) ? node779 : 46'b1001000000000000001000000001100000100000000010;
														assign node779 = (inp[14]) ? 46'b1001000000000010000000000000100000100000000000 : 46'b1001000000000110000000000000100000100000000000;
													assign node782 = (inp[8]) ? node786 : node783;
														assign node783 = (inp[10]) ? 46'b1000000000000010001000000001100000100000000000 : 46'b1000000000000100001000000001100000100000000000;
														assign node786 = (inp[14]) ? node790 : node787;
															assign node787 = (inp[10]) ? 46'b1000000000000000000000000001100000100000000010 : 46'b1000000000000100000000000001100000100000000010;
															assign node790 = (inp[10]) ? 46'b1000000000000010000000000001100000100000000010 : 46'b1000000000000110000000000000100000100000000000;
												assign node793 = (inp[5]) ? node807 : node794;
													assign node794 = (inp[14]) ? node800 : node795;
														assign node795 = (inp[10]) ? node797 : 46'b1001000000000100000000000001100000000000000010;
															assign node797 = (inp[8]) ? 46'b1001000000000000000000000001100000000000000010 : 46'b1001000000000100000000000001100000000000000010;
														assign node800 = (inp[8]) ? 46'b1001000000000010000000000001100000000000000010 : node801;
															assign node801 = (inp[10]) ? 46'b1001000000000010001000000001100000000000000000 : node802;
																assign node802 = (inp[4]) ? 46'b1001000000000000001000000001100000000000000000 : 46'b1001000000000100001000000001100000000000000000;
													assign node807 = (inp[10]) ? node817 : node808;
														assign node808 = (inp[8]) ? node814 : node809;
															assign node809 = (inp[14]) ? node811 : 46'b1000000000000100001000000001100000000000000000;
																assign node811 = (inp[4]) ? 46'b1000000000000000001000000001100000000000000000 : 46'b1000000000000100001000000001100000000000000000;
															assign node814 = (inp[4]) ? 46'b1000000000000000001000000001100000000000000010 : 46'b1000000000000100000000000001100000000000000010;
														assign node817 = (inp[4]) ? node819 : 46'b1000000000000000001000000001100000000000000010;
															assign node819 = (inp[8]) ? 46'b1000000000000010000000000000100000000000000000 : 46'b1000000000000010001000000001100000000000000000;
										assign node822 = (inp[5]) ? node856 : node823;
											assign node823 = (inp[12]) ? node835 : node824;
												assign node824 = (inp[10]) ? node832 : node825;
													assign node825 = (inp[6]) ? node829 : node826;
														assign node826 = (inp[4]) ? 46'b1001000000000000001000000001000010100000000000 : 46'b1001000000000100001000000001000010100000000000;
														assign node829 = (inp[4]) ? 46'b1001000000000010001000000001000010000000000000 : 46'b1001000000000110000000000000000010000000000000;
													assign node832 = (inp[8]) ? 46'b1001000000000010000000000000000010100000000000 : 46'b1001000000000110000000000000000010100000000000;
												assign node835 = (inp[6]) ? node843 : node836;
													assign node836 = (inp[4]) ? node838 : 46'b1001000000000110000000000000000000100000000000;
														assign node838 = (inp[14]) ? 46'b1001000000000000001000000001000000100000000000 : node839;
															assign node839 = (inp[8]) ? 46'b1001000000000010000000000001000000100000000010 : 46'b1001000000000110000000000000000000100000000000;
													assign node843 = (inp[14]) ? node849 : node844;
														assign node844 = (inp[8]) ? node846 : 46'b1001000000000100000000000001000000000000000010;
															assign node846 = (inp[10]) ? 46'b1001000000000000000000000001000000000000000010 : 46'b1001000000000100000000000001000000000000000010;
														assign node849 = (inp[8]) ? 46'b1001000000000110000000000000000000000000000000 : node850;
															assign node850 = (inp[4]) ? node852 : 46'b1001000000000000001000000001000000000000000010;
																assign node852 = (inp[10]) ? 46'b1001000000000010001000000001000000000000000000 : 46'b1001000000000000001000000001000000000000000000;
											assign node856 = (inp[6]) ? node872 : node857;
												assign node857 = (inp[4]) ? node859 : 46'b1000000000000100000000000001000010100000000010;
													assign node859 = (inp[10]) ? node863 : node860;
														assign node860 = (inp[8]) ? 46'b1000000000000010001000000001000010100000000000 : 46'b1000000000000000001000000001000000100000000000;
														assign node863 = (inp[8]) ? node867 : node864;
															assign node864 = (inp[12]) ? 46'b1000000000000110000000000000000000100000000000 : 46'b1000000000000110000000000000000010100000000000;
															assign node867 = (inp[14]) ? 46'b1000000000000010000000000000000000100000000000 : node868;
																assign node868 = (inp[12]) ? 46'b1000000000000010000000000001000000100000000010 : 46'b1000000000000010000000000001000010100000000010;
												assign node872 = (inp[12]) ? node890 : node873;
													assign node873 = (inp[10]) ? node881 : node874;
														assign node874 = (inp[4]) ? node878 : node875;
															assign node875 = (inp[14]) ? 46'b1000000000000110000000000000000010000000000000 : 46'b1000000000000100000000000000000010000000000000;
															assign node878 = (inp[14]) ? 46'b1000000000000000001000000001000010000000000000 : 46'b1000000000000000001000000001000010000000000010;
														assign node881 = (inp[4]) ? node887 : node882;
															assign node882 = (inp[8]) ? node884 : 46'b1000000000000000001000000001000010000000000010;
																assign node884 = (inp[14]) ? 46'b1000000000000010000000000001000010000000000010 : 46'b1000000000000000000000000001000010000000000010;
															assign node887 = (inp[14]) ? 46'b1000000000000010000000000000000010000000000000 : 46'b1000000000000110000000000000000010000000000000;
													assign node890 = (inp[14]) ? node892 : 46'b1000000000000010000000000001000000000000000010;
														assign node892 = (inp[8]) ? 46'b1000000000000010001000000001000000000000000000 : 46'b1000000000000100001000000001000000000000000000;
								assign node895 = (inp[9]) ? node1065 : node896;
									assign node896 = (inp[12]) ? node972 : node897;
										assign node897 = (inp[7]) ? node933 : node898;
											assign node898 = (inp[5]) ? node916 : node899;
												assign node899 = (inp[10]) ? node905 : node900;
													assign node900 = (inp[8]) ? 46'b0101000000000010001000000001100010000000000000 : node901;
														assign node901 = (inp[6]) ? 46'b0101000000000100001000000001100010000000000000 : 46'b0101000000000100001000000001100010100000000000;
													assign node905 = (inp[8]) ? node909 : node906;
														assign node906 = (inp[6]) ? 46'b0101000000000000001000000001100010000000000010 : 46'b0101000000000000001000000001100010100000000010;
														assign node909 = (inp[6]) ? 46'b0101000000000010000000000001100010000000000010 : node910;
															assign node910 = (inp[4]) ? 46'b0101000000000010000000000001100010100000000010 : node911;
																assign node911 = (inp[14]) ? 46'b0101000000000010000000000001100010100000000010 : 46'b0101000000000000000000000001100010100000000010;
												assign node916 = (inp[4]) ? node928 : node917;
													assign node917 = (inp[10]) ? node923 : node918;
														assign node918 = (inp[14]) ? 46'b0100000000000110000000000000100010100000000000 : node919;
															assign node919 = (inp[8]) ? 46'b0100000000000100000000000001100010000000000010 : 46'b0100000000000100000000000000100010000000000000;
														assign node923 = (inp[14]) ? 46'b0100000000000000001000000001100010100000000010 : node924;
															assign node924 = (inp[8]) ? 46'b0100000000000000000000000001100010000000000010 : 46'b0100000000000100000000000001100010100000000010;
													assign node928 = (inp[14]) ? node930 : 46'b0100000000000000001000000001100010100000000010;
														assign node930 = (inp[8]) ? 46'b0100000000000010001000000001100010100000000000 : 46'b0100000000000010001000000001100010000000000000;
											assign node933 = (inp[6]) ? node955 : node934;
												assign node934 = (inp[5]) ? node946 : node935;
													assign node935 = (inp[4]) ? node943 : node936;
														assign node936 = (inp[10]) ? node940 : node937;
															assign node937 = (inp[14]) ? 46'b0101000000000110000000000000000010100000000000 : 46'b0101000000000100000000000000000010100000000000;
															assign node940 = (inp[14]) ? 46'b0101000000000010000000000001000010100000000010 : 46'b0101000000000100000000000001000010100000000010;
														assign node943 = (inp[14]) ? 46'b0101000000000010001000000001000010100000000000 : 46'b0101000000000000001000000001000010100000000010;
													assign node946 = (inp[8]) ? node952 : node947;
														assign node947 = (inp[14]) ? 46'b0100000000000000001000000001000010100000000010 : node948;
															assign node948 = (inp[10]) ? 46'b0100000000000110000000000000000010100000000000 : 46'b0100000000000100001000000001000010100000000000;
														assign node952 = (inp[14]) ? 46'b0100000000000110000000000000000010100000000000 : 46'b0100000000000100000000000001000010100000000010;
												assign node955 = (inp[8]) ? node963 : node956;
													assign node956 = (inp[4]) ? node960 : node957;
														assign node957 = (inp[10]) ? 46'b0100000000000100000000000001000010000000000010 : 46'b0100000000000100000000000000000010000000000000;
														assign node960 = (inp[10]) ? 46'b0101000000000110000000000000000010000000000000 : 46'b0101000000000100001000000001000010000000000000;
													assign node963 = (inp[10]) ? node965 : 46'b0100000000000010001000000001000010000000000000;
														assign node965 = (inp[4]) ? node969 : node966;
															assign node966 = (inp[5]) ? 46'b0100000000000000000000000001000010000000000010 : 46'b0101000000000000000000000001000010000000000010;
															assign node969 = (inp[5]) ? 46'b0100000000000010000000000001000010000000000010 : 46'b0101000000000010000000000001000010000000000010;
										assign node972 = (inp[7]) ? node1022 : node973;
											assign node973 = (inp[5]) ? node995 : node974;
												assign node974 = (inp[8]) ? node984 : node975;
													assign node975 = (inp[14]) ? 46'b0101000000000100001000000001100000000000000000 : node976;
														assign node976 = (inp[6]) ? node980 : node977;
															assign node977 = (inp[4]) ? 46'b0101000000000110000000000000100000100000000000 : 46'b0101000000000100000000000000100000100000000000;
															assign node980 = (inp[10]) ? 46'b0101000000000110000000000000100000000000000000 : 46'b0101000000000100000000000000100000000000000000;
													assign node984 = (inp[6]) ? node988 : node985;
														assign node985 = (inp[14]) ? 46'b0101000000000010001000000001100000100000000000 : 46'b0101000000000000001000000001100000100000000010;
														assign node988 = (inp[14]) ? node990 : 46'b0101000000000010000000000001100000000000000010;
															assign node990 = (inp[4]) ? node992 : 46'b0101000000000110000000000000100000000000000000;
																assign node992 = (inp[10]) ? 46'b0101000000000010000000000000100000000000000000 : 46'b0101000000000010001000000001100000000000000000;
												assign node995 = (inp[6]) ? node1009 : node996;
													assign node996 = (inp[10]) ? node1000 : node997;
														assign node997 = (inp[8]) ? 46'b0100000000000000001000000001100000100000000010 : 46'b0100000000000100001000000001100000100000000000;
														assign node1000 = (inp[4]) ? node1004 : node1001;
															assign node1001 = (inp[8]) ? 46'b0100000000000000000000000001100000100000000010 : 46'b0100000000000100000000000001100000100000000010;
															assign node1004 = (inp[8]) ? node1006 : 46'b0100000000000110000000000000100000100000000000;
																assign node1006 = (inp[14]) ? 46'b0100000000000010000000000000100000100000000000 : 46'b0100000000000010000000000001100000100000000010;
													assign node1009 = (inp[14]) ? node1017 : node1010;
														assign node1010 = (inp[4]) ? 46'b0100000000000000001000000001100000000000000010 : node1011;
															assign node1011 = (inp[8]) ? node1013 : 46'b0100000000000100000000000001100000000000000010;
																assign node1013 = (inp[10]) ? 46'b0100000000000000000000000001100000000000000010 : 46'b0100000000000100000000000001100000000000000010;
														assign node1017 = (inp[10]) ? 46'b0100000000000010001000000001100000000000000000 : node1018;
															assign node1018 = (inp[4]) ? 46'b0100000000000000001000000001100000000000000000 : 46'b0100000000000100001000000001100000000000000000;
											assign node1022 = (inp[6]) ? node1042 : node1023;
												assign node1023 = (inp[8]) ? node1033 : node1024;
													assign node1024 = (inp[10]) ? node1030 : node1025;
														assign node1025 = (inp[14]) ? 46'b0101000000000100001000000001000000100000000000 : node1026;
															assign node1026 = (inp[4]) ? 46'b0100000000000100001000000001000000100000000000 : 46'b0100000000000100000000000000000000100000000000;
														assign node1030 = (inp[14]) ? 46'b0100000000000010001000000001000000100000000000 : 46'b0100000000000110000000000000000000100000000000;
													assign node1033 = (inp[14]) ? 46'b0101000000000010001000000001000000100000000000 : node1034;
														assign node1034 = (inp[5]) ? node1038 : node1035;
															assign node1035 = (inp[10]) ? 46'b0101000000000000000000000001000000100000000010 : 46'b0101000000000100000000000001000000100000000010;
															assign node1038 = (inp[4]) ? 46'b0100000000000010000000000001000000100000000010 : 46'b0100000000000000000000000001000000100000000010;
												assign node1042 = (inp[5]) ? node1050 : node1043;
													assign node1043 = (inp[8]) ? 46'b0101000000000000001000000001000000000000000010 : node1044;
														assign node1044 = (inp[4]) ? 46'b0101000000000100001000000001000000000000000000 : node1045;
															assign node1045 = (inp[14]) ? 46'b0101000000000100001000000001000000000000000000 : 46'b0101000000000100000000000000000000000000000000;
													assign node1050 = (inp[4]) ? node1056 : node1051;
														assign node1051 = (inp[10]) ? 46'b0100000000000100000000000001000000000000000010 : node1052;
															assign node1052 = (inp[14]) ? 46'b0100000000000100001000000001000000000000000000 : 46'b0100000000000100000000000000000000000000000000;
														assign node1056 = (inp[10]) ? node1062 : node1057;
															assign node1057 = (inp[8]) ? 46'b0100000000000000001000000001000000000000000010 : node1058;
																assign node1058 = (inp[14]) ? 46'b0100000000000000001000000001000000000000000000 : 46'b0100000000000100001000000001000000000000000000;
															assign node1062 = (inp[8]) ? 46'b0100000000000010000000000000000000000000000000 : 46'b0100000000000010001000000001000000000000000000;
									assign node1065 = (inp[6]) ? node1157 : node1066;
										assign node1066 = (inp[5]) ? node1102 : node1067;
											assign node1067 = (inp[7]) ? node1091 : node1068;
												assign node1068 = (inp[12]) ? node1082 : node1069;
													assign node1069 = (inp[4]) ? node1077 : node1070;
														assign node1070 = (inp[14]) ? node1072 : 46'b0001000000000100000000000001100010101000000010;
															assign node1072 = (inp[8]) ? 46'b0001000000000010000000000001100010101000000010 : node1073;
																assign node1073 = (inp[10]) ? 46'b0001000000000000001000000001100010101000000010 : 46'b0001000000000100001000000001100010101000000000;
														assign node1077 = (inp[8]) ? 46'b0001000000000000001000000001100010101000000010 : node1078;
															assign node1078 = (inp[10]) ? 46'b0001000000000010001000000001100010101000000000 : 46'b0001000000000000001000000001100010101000000000;
													assign node1082 = (inp[8]) ? node1088 : node1083;
														assign node1083 = (inp[10]) ? node1085 : 46'b0001000000000100001000000001100000101000000000;
															assign node1085 = (inp[14]) ? 46'b0001000000000000001000000001100000101000000010 : 46'b0001000000000100000000000001100000101000000010;
														assign node1088 = (inp[14]) ? 46'b0001000000000010000000000000100000101000000000 : 46'b0001000000000000001000000001100000101000000010;
												assign node1091 = (inp[8]) ? node1095 : node1092;
													assign node1092 = (inp[4]) ? 46'b0001000000000100001000000001000010101000000000 : 46'b0001000000000100000000000000000000101000000000;
													assign node1095 = (inp[10]) ? node1097 : 46'b0001000000000010001000000001000000101000000000;
														assign node1097 = (inp[4]) ? node1099 : 46'b0001000000000010000000000001000010101000000010;
															assign node1099 = (inp[14]) ? 46'b0001000000000010000000000000000000101000000000 : 46'b0001000000000010000000000001000000101000000010;
											assign node1102 = (inp[7]) ? node1134 : node1103;
												assign node1103 = (inp[12]) ? node1115 : node1104;
													assign node1104 = (inp[14]) ? node1110 : node1105;
														assign node1105 = (inp[10]) ? node1107 : 46'b0000000000000000001000000001100010101000000010;
															assign node1107 = (inp[4]) ? 46'b0000000000000010000000000001100010101000000010 : 46'b0000000000000000000000000001100010101000000010;
														assign node1110 = (inp[4]) ? node1112 : 46'b0000000000000110000000000000100010101000000000;
															assign node1112 = (inp[10]) ? 46'b0000000000000010000000000000100010101000000000 : 46'b0000000000000010001000000001100010101000000000;
													assign node1115 = (inp[8]) ? node1125 : node1116;
														assign node1116 = (inp[14]) ? 46'b0000000000000000001000000001100000101000000000 : node1117;
															assign node1117 = (inp[4]) ? node1121 : node1118;
																assign node1118 = (inp[10]) ? 46'b0000000000000100000000000001100000101000000010 : 46'b0000000000000100000000000000100000101000000000;
																assign node1121 = (inp[10]) ? 46'b0000000000000110000000000000100000101000000000 : 46'b0000000000000100001000000001100000101000000000;
														assign node1125 = (inp[10]) ? node1127 : 46'b0000000000000000001000000001100000101000000010;
															assign node1127 = (inp[14]) ? node1131 : node1128;
																assign node1128 = (inp[4]) ? 46'b0000000000000010000000000001100000101000000010 : 46'b0000000000000000000000000001100000101000000010;
																assign node1131 = (inp[4]) ? 46'b0000000000000010000000000000100000101000000000 : 46'b0000000000000010000000000001100000101000000010;
												assign node1134 = (inp[12]) ? node1144 : node1135;
													assign node1135 = (inp[8]) ? node1141 : node1136;
														assign node1136 = (inp[4]) ? node1138 : 46'b0000000000000100000000000000000010101000000000;
															assign node1138 = (inp[14]) ? 46'b0000000000000000001000000001000010101000000000 : 46'b0000000000000100001000000001000010101000000000;
														assign node1141 = (inp[10]) ? 46'b0000000000000010000000000001000010101000000010 : 46'b0000000000000100000000000001000010101000000010;
													assign node1144 = (inp[10]) ? node1152 : node1145;
														assign node1145 = (inp[8]) ? node1149 : node1146;
															assign node1146 = (inp[14]) ? 46'b0000000000000000001000000001000000101000000000 : 46'b0000000000000100001000000001000000101000000000;
															assign node1149 = (inp[14]) ? 46'b0000000000000010001000000001000000101000000000 : 46'b0000000000000000001000000001000000101000000010;
														assign node1152 = (inp[4]) ? 46'b0000000000000010000000000001000000101000000010 : node1153;
															assign node1153 = (inp[14]) ? 46'b0000000000000000001000000001000000101000000010 : 46'b0000000000000100000000000001000000101000000010;
										assign node1157 = (inp[5]) ? node1205 : node1158;
											assign node1158 = (inp[12]) ? node1186 : node1159;
												assign node1159 = (inp[7]) ? node1173 : node1160;
													assign node1160 = (inp[4]) ? node1166 : node1161;
														assign node1161 = (inp[14]) ? 46'b0001000000000100001000000001100010001000000000 : node1162;
															assign node1162 = (inp[8]) ? 46'b0001000000000100000000000001100010001000000010 : 46'b0001000000000100000000000000100010001000000000;
														assign node1166 = (inp[10]) ? node1168 : 46'b0001000000000000001000000001100010001000000010;
															assign node1168 = (inp[14]) ? node1170 : 46'b0001000000000010000000000001100010001000000010;
																assign node1170 = (inp[8]) ? 46'b0001000000000010000000000000100010001000000000 : 46'b0001000000000010001000000001100010001000000000;
													assign node1173 = (inp[10]) ? node1179 : node1174;
														assign node1174 = (inp[8]) ? 46'b0001000000000010001000000001000010001000000000 : node1175;
															assign node1175 = (inp[14]) ? 46'b0001000000000000001000000001000010001000000000 : 46'b0001000000000100001000000001000010001000000000;
														assign node1179 = (inp[4]) ? node1183 : node1180;
															assign node1180 = (inp[14]) ? 46'b0001000000000000001000000001000010001000000010 : 46'b0001000000000000000000000001000010001000000010;
															assign node1183 = (inp[14]) ? 46'b0001000000000010000000000000000010001000000000 : 46'b0001000000000010000000000001000010001000000010;
												assign node1186 = (inp[4]) ? node1196 : node1187;
													assign node1187 = (inp[14]) ? node1191 : node1188;
														assign node1188 = (inp[7]) ? 46'b0001000000000100000000000001000000001000000010 : 46'b0001000000000100000000000001100000001000000010;
														assign node1191 = (inp[8]) ? 46'b0001000000000110000000000000100000001000000000 : node1192;
															assign node1192 = (inp[10]) ? 46'b0001000000000000001000000001100000001000000010 : 46'b0001000000000100001000000001100000001000000000;
													assign node1196 = (inp[10]) ? node1198 : 46'b0001000000000000001000000001000000001000000000;
														assign node1198 = (inp[8]) ? node1200 : 46'b0001000000000110000000000000000000001000000000;
															assign node1200 = (inp[14]) ? node1202 : 46'b0001000000000010000000000001000000001000000010;
																assign node1202 = (inp[7]) ? 46'b0001000000000010000000000000000000001000000000 : 46'b0001000000000010000000000000100000001000000000;
											assign node1205 = (inp[12]) ? node1223 : node1206;
												assign node1206 = (inp[4]) ? node1216 : node1207;
													assign node1207 = (inp[7]) ? node1211 : node1208;
														assign node1208 = (inp[14]) ? 46'b0000000000000000001000000001100010001000000010 : 46'b0000000000000000000000000001100010001000000010;
														assign node1211 = (inp[14]) ? 46'b0000000000000010000000000001000010001000000010 : node1212;
															assign node1212 = (inp[8]) ? 46'b0000000000000000000000000001000010001000000010 : 46'b0000000000000100000000000001000010001000000010;
													assign node1216 = (inp[7]) ? 46'b0000000000000010000000000000000010001000000000 : node1217;
														assign node1217 = (inp[14]) ? 46'b0000000000000010001000000001100010001000000000 : node1218;
															assign node1218 = (inp[8]) ? 46'b0000000000000010000000000001100010001000000010 : 46'b0000000000000110000000000000100010001000000000;
												assign node1223 = (inp[7]) ? node1233 : node1224;
													assign node1224 = (inp[10]) ? node1230 : node1225;
														assign node1225 = (inp[14]) ? 46'b0000000000000010001000000001100000001000000000 : node1226;
															assign node1226 = (inp[8]) ? 46'b0000000000000000001000000001100000001000000010 : 46'b0000000000000100001000000001100000001000000000;
														assign node1230 = (inp[4]) ? 46'b0000000000000010000000000001100000001000000010 : 46'b0000000000000000000000000001100000001000000010;
													assign node1233 = (inp[14]) ? node1237 : node1234;
														assign node1234 = (inp[8]) ? 46'b0000000000000100000000000001000000001000000010 : 46'b0000000000000110000000000000000000001000000000;
														assign node1237 = (inp[10]) ? 46'b0000000000000000001000000001000000001000000010 : node1238;
															assign node1238 = (inp[8]) ? 46'b0000000000000010001000000001000000001000000000 : 46'b0000000000000000001000000001000000001000000000;
						assign node1242 = (inp[11]) ? node1634 : node1243;
							assign node1243 = (inp[9]) ? node1343 : node1244;
								assign node1244 = (inp[7]) ? node1262 : node1245;
									assign node1245 = (inp[12]) ? node1247 : 46'b0000000000000000000000000000000000000000000000;
										assign node1247 = (inp[6]) ? node1249 : 46'b0000000000000000000000000000000000000000000000;
											assign node1249 = (inp[0]) ? node1251 : 46'b0000000000000000000000000000000000000000000000;
												assign node1251 = (inp[5]) ? node1253 : 46'b0000000000000000000000000000000000000000000000;
													assign node1253 = (inp[14]) ? node1255 : 46'b0000000000000111000000000000100000000000100000;
														assign node1255 = (inp[8]) ? node1257 : 46'b0000000000000001001000000001100000000000100010;
															assign node1257 = (inp[4]) ? node1259 : 46'b0000000000000111000000000000100000000000100000;
																assign node1259 = (inp[10]) ? 46'b0000000000000011000000000000100000000000100000 : 46'b0000000000000011001000000001100000000000100000;
									assign node1262 = (inp[5]) ? node1280 : node1263;
										assign node1263 = (inp[6]) ? node1265 : 46'b0000000000000000000000000000000000000000000000;
											assign node1265 = (inp[0]) ? node1267 : 46'b0000000000000000000000000000000000000000000000;
												assign node1267 = (inp[8]) ? node1271 : node1268;
													assign node1268 = (inp[10]) ? 46'b0001000000000001001000000001000000000000100010 : 46'b0001000000000101001000000001000000000000100000;
													assign node1271 = (inp[10]) ? node1273 : 46'b0001000000000001001000000001000000000000100010;
														assign node1273 = (inp[4]) ? node1277 : node1274;
															assign node1274 = (inp[14]) ? 46'b0001000000000011000000000001000000000000100010 : 46'b0001000000000001000000000001000000000000100010;
															assign node1277 = (inp[14]) ? 46'b0001000000000011000000000000000000000000100000 : 46'b0001000000000011000000000001000000000000100010;
										assign node1280 = (inp[0]) ? node1320 : node1281;
											assign node1281 = (inp[12]) ? node1305 : node1282;
												assign node1282 = (inp[6]) ? node1296 : node1283;
													assign node1283 = (inp[10]) ? node1287 : node1284;
														assign node1284 = (inp[8]) ? 46'b0000000000100000001001000001000010100000000010 : 46'b0000000000100100001001000001000010100000000000;
														assign node1287 = (inp[4]) ? node1293 : node1288;
															assign node1288 = (inp[14]) ? 46'b0000000000100000001001000001000010100000000010 : node1289;
																assign node1289 = (inp[8]) ? 46'b0000000000100000000001000001000010100000000010 : 46'b0000000000100100000001000001000010100000000010;
															assign node1293 = (inp[8]) ? 46'b0000000000100010000001000000000010100000000000 : 46'b0000000000100110000001000000000010100000000000;
													assign node1296 = (inp[10]) ? node1302 : node1297;
														assign node1297 = (inp[4]) ? node1299 : 46'b0000000000100100001001000001000010000000000000;
															assign node1299 = (inp[14]) ? 46'b0000000000100000001001000001000010000000000000 : 46'b0000000000100000001001000001000010000000000010;
														assign node1302 = (inp[8]) ? 46'b0000000000100000000001000001000010000000000010 : 46'b0000000000100100000001000001000010000000000010;
												assign node1305 = (inp[10]) ? node1315 : node1306;
													assign node1306 = (inp[4]) ? 46'b0000000000100000001001000001000000000000000000 : node1307;
														assign node1307 = (inp[8]) ? 46'b0000000000100110000001000000000000000000000000 : node1308;
															assign node1308 = (inp[14]) ? 46'b0000000000100100001001000001000000000000000000 : node1309;
																assign node1309 = (inp[6]) ? 46'b0000000000100100000001000000000000000000000000 : 46'b0000000000100100000001000000000000100000000000;
													assign node1315 = (inp[6]) ? node1317 : 46'b0000000000100000001001000001000000100000000010;
														assign node1317 = (inp[8]) ? 46'b0000000000100010000001000001000000000000000010 : 46'b0000000000100100000001000001000000000000000010;
											assign node1320 = (inp[12]) ? node1336 : node1321;
												assign node1321 = (inp[6]) ? node1323 : 46'b0000000000000000000000000000000000000000000000;
													assign node1323 = (inp[14]) ? node1331 : node1324;
														assign node1324 = (inp[4]) ? node1328 : node1325;
															assign node1325 = (inp[8]) ? 46'b0000000000000001000000000001000010000000100010 : 46'b0000000000000101000000000001000010000000100010;
															assign node1328 = (inp[8]) ? 46'b0000000000000001001000000001000010000000100010 : 46'b0000000000000101001000000001000010000000100000;
														assign node1331 = (inp[10]) ? node1333 : 46'b0000000000000111000000000000000010000000100000;
															assign node1333 = (inp[4]) ? 46'b0000000000000011000000000000000010000000100000 : 46'b0000000000000011000000000001000010000000100010;
												assign node1336 = (inp[6]) ? 46'b0000000000000000000000000000000000000000000000 : node1337;
													assign node1337 = (inp[4]) ? node1339 : 46'b0000000000000001000000000001000000100000100010;
														assign node1339 = (inp[8]) ? 46'b0000000000000001001000000001000000100000100010 : 46'b0000000000000001001000000001000000100000100000;
								assign node1343 = (inp[7]) ? node1489 : node1344;
									assign node1344 = (inp[5]) ? node1426 : node1345;
										assign node1345 = (inp[6]) ? node1387 : node1346;
											assign node1346 = (inp[12]) ? node1374 : node1347;
												assign node1347 = (inp[0]) ? node1359 : node1348;
													assign node1348 = (inp[8]) ? node1356 : node1349;
														assign node1349 = (inp[10]) ? 46'b0001000000100110000000000000100010100000100000 : node1350;
															assign node1350 = (inp[4]) ? node1352 : 46'b0001000000100100000000000000100010100000100000;
																assign node1352 = (inp[14]) ? 46'b0001000000100000001000000001100010100000100000 : 46'b0001000000100100001000000001100010100000100000;
														assign node1356 = (inp[4]) ? 46'b0001000000100010000000000001100010100000100010 : 46'b0001000000100000000000000001100010100000100010;
													assign node1359 = (inp[14]) ? node1367 : node1360;
														assign node1360 = (inp[8]) ? node1362 : 46'b0001000000000100000000000000100010100000100000;
															assign node1362 = (inp[10]) ? node1364 : 46'b0001000000000000001000000001100010100000100010;
																assign node1364 = (inp[4]) ? 46'b0001000000000010000000000001100010100000100010 : 46'b0001000000000000000000000001100010100000100010;
														assign node1367 = (inp[4]) ? node1369 : 46'b0001000000000110000000000000100010100000100000;
															assign node1369 = (inp[8]) ? node1371 : 46'b0001000000000010001000000001100010100000100000;
																assign node1371 = (inp[10]) ? 46'b0001000000000010000000000000100010100000100000 : 46'b0001000000000010001000000001100010100000100000;
												assign node1374 = (inp[0]) ? node1378 : node1375;
													assign node1375 = (inp[14]) ? 46'b0001000000100010001000000001100000100000100000 : 46'b0001000000100010000000000001100000100000100010;
													assign node1378 = (inp[8]) ? node1382 : node1379;
														assign node1379 = (inp[10]) ? 46'b0001000000000000001000000001100000100000100010 : 46'b0001000000000000001000000001100000100000100000;
														assign node1382 = (inp[10]) ? 46'b0001000000000010000000000000100000100000100000 : node1383;
															assign node1383 = (inp[14]) ? 46'b0001000000000010001000000001100000100000100000 : 46'b0001000000000000001000000001100000100000100010;
											assign node1387 = (inp[0]) ? node1405 : node1388;
												assign node1388 = (inp[10]) ? node1394 : node1389;
													assign node1389 = (inp[4]) ? node1391 : 46'b0001000000100100001000000001100000000000100000;
														assign node1391 = (inp[8]) ? 46'b0001000000100010001000000001100010000000100000 : 46'b0001000000100000001000000001100010000000100000;
													assign node1394 = (inp[4]) ? node1398 : node1395;
														assign node1395 = (inp[14]) ? 46'b0001000000100010000000000001100010000000100010 : 46'b0001000000100000000000000001100010000000100010;
														assign node1398 = (inp[14]) ? node1402 : node1399;
															assign node1399 = (inp[12]) ? 46'b0001000000100110000000000000100000000000100000 : 46'b0001000000100110000000000000100010000000100000;
															assign node1402 = (inp[12]) ? 46'b0001000000100010000000000000100000000000100000 : 46'b0001000000100010000000000000100010000000100000;
												assign node1405 = (inp[12]) ? node1423 : node1406;
													assign node1406 = (inp[14]) ? node1418 : node1407;
														assign node1407 = (inp[8]) ? node1415 : node1408;
															assign node1408 = (inp[4]) ? node1412 : node1409;
																assign node1409 = (inp[10]) ? 46'b0001000000000100000000000001100010000000100010 : 46'b0001000000000100000000000000100010000000100000;
																assign node1412 = (inp[10]) ? 46'b0001000000000110000000000000100010000000100000 : 46'b0001000000000100001000000001100010000000100000;
															assign node1415 = (inp[4]) ? 46'b0001000000000000001000000001100010000000100010 : 46'b0001000000000100000000000001100010000000100010;
														assign node1418 = (inp[4]) ? node1420 : 46'b0001000000000100001000000001100010000000100000;
															assign node1420 = (inp[10]) ? 46'b0001000000000010001000000001100010000000100000 : 46'b0001000000000000001000000001100010000000100000;
													assign node1423 = (inp[10]) ? 46'b0001000000000010000000000001100000000000100010 : 46'b0001000000000110000000000000100000000000100000;
										assign node1426 = (inp[6]) ? node1458 : node1427;
											assign node1427 = (inp[12]) ? node1447 : node1428;
												assign node1428 = (inp[8]) ? node1436 : node1429;
													assign node1429 = (inp[0]) ? node1433 : node1430;
														assign node1430 = (inp[10]) ? 46'b0000000000100000001000000001100010100000100010 : 46'b0000000000100100001000000001100010100000100000;
														assign node1433 = (inp[10]) ? 46'b0000000000000010001000000001100010100000100000 : 46'b0000000000000000001000000001100010100000100000;
													assign node1436 = (inp[0]) ? node1442 : node1437;
														assign node1437 = (inp[4]) ? node1439 : 46'b0000000000100010000000000001100010100000100010;
															assign node1439 = (inp[10]) ? 46'b0000000000100010000000000000100010100000100000 : 46'b0000000000100010001000000001100010100000100000;
														assign node1442 = (inp[14]) ? node1444 : 46'b0000000000000100000000000001100010100000100010;
															assign node1444 = (inp[4]) ? 46'b0000000000000010000000000000100010100000100000 : 46'b0000000000000110000000000000100010100000100000;
												assign node1447 = (inp[4]) ? node1455 : node1448;
													assign node1448 = (inp[10]) ? 46'b0000000000000100000000000001100000100000100010 : node1449;
														assign node1449 = (inp[0]) ? 46'b0000000000000100000000000000100000100000100000 : node1450;
															assign node1450 = (inp[8]) ? 46'b0000000000100110000000000000100000100000100000 : 46'b0000000000100100000000000000100000100000100000;
													assign node1455 = (inp[0]) ? 46'b0000000000000000001000000001100000100000100000 : 46'b0000000000100000001000000001100000100000100010;
											assign node1458 = (inp[12]) ? node1472 : node1459;
												assign node1459 = (inp[0]) ? node1465 : node1460;
													assign node1460 = (inp[8]) ? 46'b0000000000100010000000000001100010000000100010 : node1461;
														assign node1461 = (inp[4]) ? 46'b0000000000100000001000000001100010000000100000 : 46'b0000000000100000001000000001100010000000100010;
													assign node1465 = (inp[4]) ? node1469 : node1466;
														assign node1466 = (inp[8]) ? 46'b0000000000000100000000000001100010000000100010 : 46'b0000000000000000001000000001100010000000100010;
														assign node1469 = (inp[14]) ? 46'b0000000000000010000000000000100010000000100000 : 46'b0000000000000110000000000000100010000000100000;
												assign node1472 = (inp[0]) ? node1484 : node1473;
													assign node1473 = (inp[14]) ? node1479 : node1474;
														assign node1474 = (inp[8]) ? node1476 : 46'b0000000000100100001000000001100000000000100000;
															assign node1476 = (inp[10]) ? 46'b0000000000100000000000000001100000000000100010 : 46'b0000000000100000001000000001100000000000100010;
														assign node1479 = (inp[8]) ? 46'b0000000000100010001000000001100000000000100000 : node1480;
															assign node1480 = (inp[10]) ? 46'b0000000000100010001000000001100000000000100000 : 46'b0000000000100000001000000001100000000000100000;
													assign node1484 = (inp[4]) ? node1486 : 46'b0000000000000000001000000001100000000000100010;
														assign node1486 = (inp[10]) ? 46'b0000000000000010001000000001100000000000100000 : 46'b0000000000000000001000000001100000000000100000;
									assign node1489 = (inp[6]) ? node1559 : node1490;
										assign node1490 = (inp[0]) ? node1530 : node1491;
											assign node1491 = (inp[5]) ? node1509 : node1492;
												assign node1492 = (inp[4]) ? node1502 : node1493;
													assign node1493 = (inp[14]) ? node1497 : node1494;
														assign node1494 = (inp[8]) ? 46'b0001000000100000000000000001000010100000100010 : 46'b0001000000100100000000000001000010100000100010;
														assign node1497 = (inp[10]) ? node1499 : 46'b0001000000100100001000000001000010100000100000;
															assign node1499 = (inp[12]) ? 46'b0001000000100000001000000001000000100000100010 : 46'b0001000000100000001000000001000010100000100010;
													assign node1502 = (inp[14]) ? node1504 : 46'b0001000000100000001000000001000000100000100010;
														assign node1504 = (inp[8]) ? node1506 : 46'b0001000000100010001000000001000000100000100000;
															assign node1506 = (inp[12]) ? 46'b0001000000100010000000000000000000100000100000 : 46'b0001000000100010000000000000000010100000100000;
												assign node1509 = (inp[14]) ? node1521 : node1510;
													assign node1510 = (inp[8]) ? node1512 : 46'b0000000000100100000000000000000010100000100000;
														assign node1512 = (inp[4]) ? node1518 : node1513;
															assign node1513 = (inp[10]) ? node1515 : 46'b0000000000100100000000000001000010100000100010;
																assign node1515 = (inp[12]) ? 46'b0000000000100000000000000001000000100000100010 : 46'b0000000000100000000000000001000010100000100010;
															assign node1518 = (inp[12]) ? 46'b0000000000100000001000000001000000100000100010 : 46'b0000000000100000001000000001000010100000100010;
													assign node1521 = (inp[8]) ? node1525 : node1522;
														assign node1522 = (inp[10]) ? 46'b0000000000100000001000000001000010100000100010 : 46'b0000000000100100001000000001000010100000100000;
														assign node1525 = (inp[4]) ? 46'b0000000000100010001000000001000010100000100000 : node1526;
															assign node1526 = (inp[12]) ? 46'b0000000000100110000000000000000000100000100000 : 46'b0000000000100110000000000000000010100000100000;
											assign node1530 = (inp[12]) ? node1546 : node1531;
												assign node1531 = (inp[14]) ? node1539 : node1532;
													assign node1532 = (inp[10]) ? node1536 : node1533;
														assign node1533 = (inp[5]) ? 46'b0000000000000100000000000000000010100000100000 : 46'b0001000000000100000000000000000010100000100000;
														assign node1536 = (inp[5]) ? 46'b0000000000000000000000000001000010100000100010 : 46'b0001000000000100000000000001000010100000100010;
													assign node1539 = (inp[5]) ? node1543 : node1540;
														assign node1540 = (inp[10]) ? 46'b0001000000000010001000000001000010100000100000 : 46'b0001000000000000001000000001000010100000100000;
														assign node1543 = (inp[10]) ? 46'b0000000000000000001000000001000010100000100010 : 46'b0000000000000000001000000001000010100000100000;
												assign node1546 = (inp[10]) ? node1554 : node1547;
													assign node1547 = (inp[8]) ? node1551 : node1548;
														assign node1548 = (inp[14]) ? 46'b0000000000000100001000000001000000100000100000 : 46'b0001000000000100001000000001000000100000100000;
														assign node1551 = (inp[4]) ? 46'b0000000000000010001000000001000000100000100000 : 46'b0000000000000110000000000000000000100000100000;
													assign node1554 = (inp[4]) ? 46'b0001000000000110000000000000000000100000100000 : node1555;
														assign node1555 = (inp[5]) ? 46'b0000000000000000000000000001000000100000100010 : 46'b0001000000000000000000000001000000100000100010;
										assign node1559 = (inp[12]) ? node1603 : node1560;
											assign node1560 = (inp[0]) ? node1584 : node1561;
												assign node1561 = (inp[5]) ? node1573 : node1562;
													assign node1562 = (inp[14]) ? node1568 : node1563;
														assign node1563 = (inp[10]) ? 46'b0001000000100010000000000001000010000000100010 : node1564;
															assign node1564 = (inp[8]) ? 46'b0001000000100000001000000001000010000000100010 : 46'b0001000000100100001000000001000010000000100000;
														assign node1568 = (inp[8]) ? node1570 : 46'b0001000000100010001000000001000010000000100000;
															assign node1570 = (inp[4]) ? 46'b0001000000100010000000000000000010000000100000 : 46'b0001000000100110000000000000000010000000100000;
													assign node1573 = (inp[8]) ? node1577 : node1574;
														assign node1574 = (inp[10]) ? 46'b0000000000100110000000000000000010000000100000 : 46'b0000000000100100000000000000000010000000100000;
														assign node1577 = (inp[10]) ? node1581 : node1578;
															assign node1578 = (inp[4]) ? 46'b0000000000100010001000000001000010000000100000 : 46'b0000000000100110000000000000000010000000100000;
															assign node1581 = (inp[4]) ? 46'b0000000000100010000000000000000010000000100000 : 46'b0000000000100010000000000001000010000000100010;
												assign node1584 = (inp[14]) ? node1594 : node1585;
													assign node1585 = (inp[4]) ? node1591 : node1586;
														assign node1586 = (inp[5]) ? node1588 : 46'b0001000000000100000000000001000010000000100010;
															assign node1588 = (inp[8]) ? 46'b0000000000000100000000000001000010000000100010 : 46'b0000000000000100000000000000000010000000100000;
														assign node1591 = (inp[8]) ? 46'b0001000000000010000000000001000010000000100010 : 46'b0001000000000110000000000000000010000000100000;
													assign node1594 = (inp[8]) ? 46'b0001000000000010000000000000000010000000100000 : node1595;
														assign node1595 = (inp[5]) ? node1597 : 46'b0001000000000000001000000001000010000000100000;
															assign node1597 = (inp[4]) ? node1599 : 46'b0000000000000000001000000001000010000000100010;
																assign node1599 = (inp[10]) ? 46'b0000000000000010001000000001000010000000100000 : 46'b0000000000000000001000000001000010000000100000;
											assign node1603 = (inp[10]) ? node1615 : node1604;
												assign node1604 = (inp[8]) ? node1608 : node1605;
													assign node1605 = (inp[0]) ? 46'b0001000000000100001000000001000000000000100000 : 46'b0001000000100100001000000001000000000000100000;
													assign node1608 = (inp[14]) ? node1612 : node1609;
														assign node1609 = (inp[0]) ? 46'b0001000000000100000000000001000000000000100010 : 46'b0001000000100100000000000001000000000000100010;
														assign node1612 = (inp[0]) ? 46'b0001000000000010001000000001000000000000100000 : 46'b0001000000100110000000000000000000000000100000;
												assign node1615 = (inp[8]) ? node1627 : node1616;
													assign node1616 = (inp[4]) ? node1624 : node1617;
														assign node1617 = (inp[14]) ? node1619 : 46'b0000000000000100000000000001000000000000100010;
															assign node1619 = (inp[5]) ? 46'b0000000000000000001000000001000000000000100010 : node1620;
																assign node1620 = (inp[0]) ? 46'b0001000000000000001000000001000000000000100010 : 46'b0001000000100000001000000001000000000000100010;
														assign node1624 = (inp[5]) ? 46'b0000000000000010001000000001000000000000100000 : 46'b0001000000000010001000000001000000000000100000;
													assign node1627 = (inp[0]) ? node1631 : node1628;
														assign node1628 = (inp[5]) ? 46'b0000000000100010000000000001000000000000100010 : 46'b0001000000100010000000000001000000000000100010;
														assign node1631 = (inp[4]) ? 46'b0000000000000010000000000000000000000000100000 : 46'b0001000000000010000000000001000000000000100010;
							assign node1634 = (inp[7]) ? node1672 : node1635;
								assign node1635 = (inp[5]) ? node1647 : node1636;
									assign node1636 = (inp[9]) ? 46'b0000000000000000000000000000000000000000000000 : node1637;
										assign node1637 = (inp[0]) ? 46'b0000000000000000000000000000000000000000000000 : node1638;
											assign node1638 = (inp[6]) ? node1642 : node1639;
												assign node1639 = (inp[12]) ? 46'b0001000000100000001000000001100000100000100000 : 46'b0000000000000000000000000000000000000000000000;
												assign node1642 = (inp[12]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0001000000100010000000000000100010000000100000;
									assign node1647 = (inp[9]) ? node1663 : node1648;
										assign node1648 = (inp[0]) ? node1656 : node1649;
											assign node1649 = (inp[12]) ? node1653 : node1650;
												assign node1650 = (inp[6]) ? 46'b0000000000100010000000000000100010000000100000 : 46'b0000000000000000000000000000000000000000000000;
												assign node1653 = (inp[6]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0000000000100000001000000001100000100000100000;
											assign node1656 = (inp[12]) ? node1660 : node1657;
												assign node1657 = (inp[6]) ? 46'b0000000010000000000000000001100010000000000010 : 46'b0000000010000000000000000001100010100000000010;
												assign node1660 = (inp[6]) ? 46'b0000000010000000000000000001100000000000000010 : 46'b0000000010000000000000000001100000100000000010;
										assign node1663 = (inp[0]) ? 46'b0000000000000000000000000000000000000000000000 : node1664;
											assign node1664 = (inp[6]) ? node1668 : node1665;
												assign node1665 = (inp[12]) ? 46'b0000000010000000000000000001100000100001000010 : 46'b0000000010000000000000000001100010100001000010;
												assign node1668 = (inp[12]) ? 46'b0000000010000000000000000001100000000001000010 : 46'b0000000010000000000000000001100010000001000010;
								assign node1672 = (inp[5]) ? node1698 : node1673;
									assign node1673 = (inp[0]) ? node1689 : node1674;
										assign node1674 = (inp[9]) ? node1682 : node1675;
											assign node1675 = (inp[12]) ? node1679 : node1676;
												assign node1676 = (inp[6]) ? 46'b0001000000100010000000000000000010000000100000 : 46'b0000000000000000000000000000000000000000000000;
												assign node1679 = (inp[6]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0001000000100000001000000001000000100000100000;
											assign node1682 = (inp[12]) ? node1686 : node1683;
												assign node1683 = (inp[6]) ? 46'b0001000010000100000000000000000010000001000000 : 46'b0001000010000100000000000000000010100001000000;
												assign node1686 = (inp[6]) ? 46'b0001000010000100000000000000000000000001000000 : 46'b0001000010000100000000000000000000100001000000;
										assign node1689 = (inp[9]) ? 46'b0000000000000000000000000000000000000000000000 : node1690;
											assign node1690 = (inp[6]) ? node1694 : node1691;
												assign node1691 = (inp[12]) ? 46'b0001000010000100000000000000000000100000000000 : 46'b0001000010000100000000000000000010100000000000;
												assign node1694 = (inp[12]) ? 46'b0001000010000100000000000000000000000000000000 : 46'b0001000010000100000000000000000010000000000000;
									assign node1698 = (inp[9]) ? 46'b0000000000000000000000000000000000000000000000 : node1699;
										assign node1699 = (inp[0]) ? 46'b0000000000000000000000000000000000000000000000 : node1700;
											assign node1700 = (inp[12]) ? node1704 : node1701;
												assign node1701 = (inp[6]) ? 46'b0000000000100010000000000000000010000000100000 : 46'b0000000000000000000000000000000000000000000000;
												assign node1704 = (inp[6]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0000000000100000001000000001000000100000100000;

endmodule