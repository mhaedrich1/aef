module dtc_split25_bm27 (
	input  wire [16-1:0] inp,
	output wire [16-1:0] outp
);

	wire [16-1:0] node1;
	wire [16-1:0] node2;
	wire [16-1:0] node3;
	wire [16-1:0] node4;
	wire [16-1:0] node5;
	wire [16-1:0] node6;
	wire [16-1:0] node7;
	wire [16-1:0] node8;
	wire [16-1:0] node9;
	wire [16-1:0] node10;
	wire [16-1:0] node11;
	wire [16-1:0] node12;
	wire [16-1:0] node13;
	wire [16-1:0] node16;
	wire [16-1:0] node19;
	wire [16-1:0] node20;
	wire [16-1:0] node22;
	wire [16-1:0] node23;
	wire [16-1:0] node28;
	wire [16-1:0] node29;
	wire [16-1:0] node30;
	wire [16-1:0] node34;
	wire [16-1:0] node35;
	wire [16-1:0] node39;
	wire [16-1:0] node40;
	wire [16-1:0] node41;
	wire [16-1:0] node42;
	wire [16-1:0] node45;
	wire [16-1:0] node48;
	wire [16-1:0] node51;
	wire [16-1:0] node53;
	wire [16-1:0] node54;
	wire [16-1:0] node55;
	wire [16-1:0] node56;
	wire [16-1:0] node62;
	wire [16-1:0] node63;
	wire [16-1:0] node64;
	wire [16-1:0] node65;
	wire [16-1:0] node66;
	wire [16-1:0] node69;
	wire [16-1:0] node71;
	wire [16-1:0] node74;
	wire [16-1:0] node76;
	wire [16-1:0] node79;
	wire [16-1:0] node80;
	wire [16-1:0] node81;
	wire [16-1:0] node82;
	wire [16-1:0] node86;
	wire [16-1:0] node90;
	wire [16-1:0] node91;
	wire [16-1:0] node92;
	wire [16-1:0] node94;
	wire [16-1:0] node98;
	wire [16-1:0] node99;
	wire [16-1:0] node101;
	wire [16-1:0] node104;
	wire [16-1:0] node107;
	wire [16-1:0] node108;
	wire [16-1:0] node109;
	wire [16-1:0] node110;
	wire [16-1:0] node111;
	wire [16-1:0] node112;
	wire [16-1:0] node115;
	wire [16-1:0] node119;
	wire [16-1:0] node120;
	wire [16-1:0] node123;
	wire [16-1:0] node124;
	wire [16-1:0] node125;
	wire [16-1:0] node127;
	wire [16-1:0] node131;
	wire [16-1:0] node133;
	wire [16-1:0] node136;
	wire [16-1:0] node137;
	wire [16-1:0] node138;
	wire [16-1:0] node140;
	wire [16-1:0] node142;
	wire [16-1:0] node145;
	wire [16-1:0] node146;
	wire [16-1:0] node147;
	wire [16-1:0] node149;
	wire [16-1:0] node154;
	wire [16-1:0] node155;
	wire [16-1:0] node156;
	wire [16-1:0] node157;
	wire [16-1:0] node163;
	wire [16-1:0] node164;
	wire [16-1:0] node165;
	wire [16-1:0] node166;
	wire [16-1:0] node169;
	wire [16-1:0] node171;
	wire [16-1:0] node174;
	wire [16-1:0] node175;
	wire [16-1:0] node176;
	wire [16-1:0] node179;
	wire [16-1:0] node182;
	wire [16-1:0] node184;
	wire [16-1:0] node187;
	wire [16-1:0] node188;
	wire [16-1:0] node190;
	wire [16-1:0] node191;
	wire [16-1:0] node193;
	wire [16-1:0] node197;
	wire [16-1:0] node198;
	wire [16-1:0] node201;
	wire [16-1:0] node202;
	wire [16-1:0] node205;
	wire [16-1:0] node207;
	wire [16-1:0] node208;
	wire [16-1:0] node212;
	wire [16-1:0] node213;
	wire [16-1:0] node214;
	wire [16-1:0] node215;
	wire [16-1:0] node216;
	wire [16-1:0] node217;
	wire [16-1:0] node219;
	wire [16-1:0] node222;
	wire [16-1:0] node223;
	wire [16-1:0] node227;
	wire [16-1:0] node228;
	wire [16-1:0] node229;
	wire [16-1:0] node233;
	wire [16-1:0] node234;
	wire [16-1:0] node236;
	wire [16-1:0] node237;
	wire [16-1:0] node241;
	wire [16-1:0] node244;
	wire [16-1:0] node245;
	wire [16-1:0] node246;
	wire [16-1:0] node248;
	wire [16-1:0] node251;
	wire [16-1:0] node252;
	wire [16-1:0] node256;
	wire [16-1:0] node257;
	wire [16-1:0] node258;
	wire [16-1:0] node263;
	wire [16-1:0] node264;
	wire [16-1:0] node265;
	wire [16-1:0] node266;
	wire [16-1:0] node267;
	wire [16-1:0] node270;
	wire [16-1:0] node273;
	wire [16-1:0] node275;
	wire [16-1:0] node278;
	wire [16-1:0] node280;
	wire [16-1:0] node281;
	wire [16-1:0] node283;
	wire [16-1:0] node287;
	wire [16-1:0] node288;
	wire [16-1:0] node289;
	wire [16-1:0] node290;
	wire [16-1:0] node291;
	wire [16-1:0] node296;
	wire [16-1:0] node297;
	wire [16-1:0] node298;
	wire [16-1:0] node300;
	wire [16-1:0] node303;
	wire [16-1:0] node304;
	wire [16-1:0] node308;
	wire [16-1:0] node310;
	wire [16-1:0] node313;
	wire [16-1:0] node314;
	wire [16-1:0] node315;
	wire [16-1:0] node316;
	wire [16-1:0] node320;
	wire [16-1:0] node322;
	wire [16-1:0] node326;
	wire [16-1:0] node327;
	wire [16-1:0] node328;
	wire [16-1:0] node329;
	wire [16-1:0] node330;
	wire [16-1:0] node331;
	wire [16-1:0] node336;
	wire [16-1:0] node337;
	wire [16-1:0] node339;
	wire [16-1:0] node342;
	wire [16-1:0] node343;
	wire [16-1:0] node347;
	wire [16-1:0] node348;
	wire [16-1:0] node350;
	wire [16-1:0] node351;
	wire [16-1:0] node355;
	wire [16-1:0] node356;
	wire [16-1:0] node357;
	wire [16-1:0] node360;
	wire [16-1:0] node363;
	wire [16-1:0] node365;
	wire [16-1:0] node368;
	wire [16-1:0] node369;
	wire [16-1:0] node370;
	wire [16-1:0] node371;
	wire [16-1:0] node372;
	wire [16-1:0] node375;
	wire [16-1:0] node377;
	wire [16-1:0] node380;
	wire [16-1:0] node381;
	wire [16-1:0] node384;
	wire [16-1:0] node385;
	wire [16-1:0] node389;
	wire [16-1:0] node390;
	wire [16-1:0] node393;
	wire [16-1:0] node394;
	wire [16-1:0] node397;
	wire [16-1:0] node400;
	wire [16-1:0] node401;
	wire [16-1:0] node403;
	wire [16-1:0] node405;
	wire [16-1:0] node406;
	wire [16-1:0] node410;
	wire [16-1:0] node411;
	wire [16-1:0] node414;
	wire [16-1:0] node416;
	wire [16-1:0] node418;
	wire [16-1:0] node421;
	wire [16-1:0] node422;
	wire [16-1:0] node423;
	wire [16-1:0] node424;
	wire [16-1:0] node425;
	wire [16-1:0] node426;
	wire [16-1:0] node427;
	wire [16-1:0] node428;
	wire [16-1:0] node432;
	wire [16-1:0] node435;
	wire [16-1:0] node436;
	wire [16-1:0] node438;
	wire [16-1:0] node442;
	wire [16-1:0] node443;
	wire [16-1:0] node444;
	wire [16-1:0] node445;
	wire [16-1:0] node449;
	wire [16-1:0] node452;
	wire [16-1:0] node455;
	wire [16-1:0] node456;
	wire [16-1:0] node457;
	wire [16-1:0] node458;
	wire [16-1:0] node459;
	wire [16-1:0] node460;
	wire [16-1:0] node464;
	wire [16-1:0] node466;
	wire [16-1:0] node470;
	wire [16-1:0] node471;
	wire [16-1:0] node473;
	wire [16-1:0] node475;
	wire [16-1:0] node476;
	wire [16-1:0] node481;
	wire [16-1:0] node482;
	wire [16-1:0] node484;
	wire [16-1:0] node486;
	wire [16-1:0] node489;
	wire [16-1:0] node490;
	wire [16-1:0] node491;
	wire [16-1:0] node494;
	wire [16-1:0] node495;
	wire [16-1:0] node499;
	wire [16-1:0] node501;
	wire [16-1:0] node504;
	wire [16-1:0] node505;
	wire [16-1:0] node506;
	wire [16-1:0] node507;
	wire [16-1:0] node509;
	wire [16-1:0] node512;
	wire [16-1:0] node513;
	wire [16-1:0] node516;
	wire [16-1:0] node518;
	wire [16-1:0] node521;
	wire [16-1:0] node522;
	wire [16-1:0] node524;
	wire [16-1:0] node525;
	wire [16-1:0] node528;
	wire [16-1:0] node531;
	wire [16-1:0] node532;
	wire [16-1:0] node533;
	wire [16-1:0] node535;
	wire [16-1:0] node537;
	wire [16-1:0] node540;
	wire [16-1:0] node543;
	wire [16-1:0] node545;
	wire [16-1:0] node548;
	wire [16-1:0] node549;
	wire [16-1:0] node550;
	wire [16-1:0] node551;
	wire [16-1:0] node552;
	wire [16-1:0] node556;
	wire [16-1:0] node557;
	wire [16-1:0] node561;
	wire [16-1:0] node563;
	wire [16-1:0] node564;
	wire [16-1:0] node567;
	wire [16-1:0] node570;
	wire [16-1:0] node571;
	wire [16-1:0] node574;
	wire [16-1:0] node575;
	wire [16-1:0] node576;
	wire [16-1:0] node578;
	wire [16-1:0] node582;
	wire [16-1:0] node583;
	wire [16-1:0] node584;
	wire [16-1:0] node586;
	wire [16-1:0] node591;
	wire [16-1:0] node592;
	wire [16-1:0] node593;
	wire [16-1:0] node594;
	wire [16-1:0] node595;
	wire [16-1:0] node596;
	wire [16-1:0] node597;
	wire [16-1:0] node601;
	wire [16-1:0] node602;
	wire [16-1:0] node606;
	wire [16-1:0] node608;
	wire [16-1:0] node611;
	wire [16-1:0] node612;
	wire [16-1:0] node614;
	wire [16-1:0] node615;
	wire [16-1:0] node619;
	wire [16-1:0] node620;
	wire [16-1:0] node621;
	wire [16-1:0] node622;
	wire [16-1:0] node626;
	wire [16-1:0] node629;
	wire [16-1:0] node631;
	wire [16-1:0] node634;
	wire [16-1:0] node635;
	wire [16-1:0] node636;
	wire [16-1:0] node637;
	wire [16-1:0] node638;
	wire [16-1:0] node640;
	wire [16-1:0] node645;
	wire [16-1:0] node646;
	wire [16-1:0] node649;
	wire [16-1:0] node650;
	wire [16-1:0] node654;
	wire [16-1:0] node655;
	wire [16-1:0] node656;
	wire [16-1:0] node658;
	wire [16-1:0] node661;
	wire [16-1:0] node662;
	wire [16-1:0] node666;
	wire [16-1:0] node667;
	wire [16-1:0] node668;
	wire [16-1:0] node671;
	wire [16-1:0] node674;
	wire [16-1:0] node676;
	wire [16-1:0] node679;
	wire [16-1:0] node680;
	wire [16-1:0] node681;
	wire [16-1:0] node682;
	wire [16-1:0] node683;
	wire [16-1:0] node684;
	wire [16-1:0] node685;
	wire [16-1:0] node687;
	wire [16-1:0] node693;
	wire [16-1:0] node695;
	wire [16-1:0] node696;
	wire [16-1:0] node699;
	wire [16-1:0] node702;
	wire [16-1:0] node703;
	wire [16-1:0] node704;
	wire [16-1:0] node705;
	wire [16-1:0] node709;
	wire [16-1:0] node710;
	wire [16-1:0] node712;
	wire [16-1:0] node713;
	wire [16-1:0] node718;
	wire [16-1:0] node719;
	wire [16-1:0] node722;
	wire [16-1:0] node723;
	wire [16-1:0] node727;
	wire [16-1:0] node728;
	wire [16-1:0] node729;
	wire [16-1:0] node731;
	wire [16-1:0] node734;
	wire [16-1:0] node735;
	wire [16-1:0] node737;
	wire [16-1:0] node739;
	wire [16-1:0] node741;
	wire [16-1:0] node745;
	wire [16-1:0] node746;
	wire [16-1:0] node747;
	wire [16-1:0] node749;
	wire [16-1:0] node753;
	wire [16-1:0] node755;
	wire [16-1:0] node758;
	wire [16-1:0] node759;
	wire [16-1:0] node760;
	wire [16-1:0] node761;
	wire [16-1:0] node762;
	wire [16-1:0] node763;
	wire [16-1:0] node764;
	wire [16-1:0] node765;
	wire [16-1:0] node767;
	wire [16-1:0] node770;
	wire [16-1:0] node771;
	wire [16-1:0] node774;
	wire [16-1:0] node776;
	wire [16-1:0] node779;
	wire [16-1:0] node780;
	wire [16-1:0] node781;
	wire [16-1:0] node784;
	wire [16-1:0] node787;
	wire [16-1:0] node788;
	wire [16-1:0] node792;
	wire [16-1:0] node793;
	wire [16-1:0] node794;
	wire [16-1:0] node796;
	wire [16-1:0] node797;
	wire [16-1:0] node802;
	wire [16-1:0] node803;
	wire [16-1:0] node805;
	wire [16-1:0] node808;
	wire [16-1:0] node809;
	wire [16-1:0] node813;
	wire [16-1:0] node814;
	wire [16-1:0] node815;
	wire [16-1:0] node816;
	wire [16-1:0] node817;
	wire [16-1:0] node822;
	wire [16-1:0] node823;
	wire [16-1:0] node824;
	wire [16-1:0] node827;
	wire [16-1:0] node830;
	wire [16-1:0] node831;
	wire [16-1:0] node832;
	wire [16-1:0] node837;
	wire [16-1:0] node838;
	wire [16-1:0] node840;
	wire [16-1:0] node843;
	wire [16-1:0] node844;
	wire [16-1:0] node846;
	wire [16-1:0] node849;
	wire [16-1:0] node850;
	wire [16-1:0] node851;
	wire [16-1:0] node855;
	wire [16-1:0] node858;
	wire [16-1:0] node859;
	wire [16-1:0] node860;
	wire [16-1:0] node861;
	wire [16-1:0] node863;
	wire [16-1:0] node865;
	wire [16-1:0] node867;
	wire [16-1:0] node870;
	wire [16-1:0] node872;
	wire [16-1:0] node875;
	wire [16-1:0] node876;
	wire [16-1:0] node877;
	wire [16-1:0] node879;
	wire [16-1:0] node882;
	wire [16-1:0] node883;
	wire [16-1:0] node886;
	wire [16-1:0] node887;
	wire [16-1:0] node892;
	wire [16-1:0] node893;
	wire [16-1:0] node894;
	wire [16-1:0] node895;
	wire [16-1:0] node897;
	wire [16-1:0] node899;
	wire [16-1:0] node903;
	wire [16-1:0] node905;
	wire [16-1:0] node908;
	wire [16-1:0] node909;
	wire [16-1:0] node910;
	wire [16-1:0] node914;
	wire [16-1:0] node915;
	wire [16-1:0] node918;
	wire [16-1:0] node920;
	wire [16-1:0] node922;
	wire [16-1:0] node925;
	wire [16-1:0] node926;
	wire [16-1:0] node927;
	wire [16-1:0] node928;
	wire [16-1:0] node929;
	wire [16-1:0] node930;
	wire [16-1:0] node931;
	wire [16-1:0] node934;
	wire [16-1:0] node937;
	wire [16-1:0] node938;
	wire [16-1:0] node942;
	wire [16-1:0] node943;
	wire [16-1:0] node945;
	wire [16-1:0] node947;
	wire [16-1:0] node950;
	wire [16-1:0] node951;
	wire [16-1:0] node955;
	wire [16-1:0] node956;
	wire [16-1:0] node957;
	wire [16-1:0] node958;
	wire [16-1:0] node959;
	wire [16-1:0] node964;
	wire [16-1:0] node965;
	wire [16-1:0] node968;
	wire [16-1:0] node971;
	wire [16-1:0] node973;
	wire [16-1:0] node975;
	wire [16-1:0] node978;
	wire [16-1:0] node979;
	wire [16-1:0] node980;
	wire [16-1:0] node981;
	wire [16-1:0] node983;
	wire [16-1:0] node987;
	wire [16-1:0] node990;
	wire [16-1:0] node991;
	wire [16-1:0] node992;
	wire [16-1:0] node994;
	wire [16-1:0] node997;
	wire [16-1:0] node998;
	wire [16-1:0] node1001;
	wire [16-1:0] node1003;
	wire [16-1:0] node1006;
	wire [16-1:0] node1008;
	wire [16-1:0] node1009;
	wire [16-1:0] node1013;
	wire [16-1:0] node1014;
	wire [16-1:0] node1015;
	wire [16-1:0] node1016;
	wire [16-1:0] node1017;
	wire [16-1:0] node1020;
	wire [16-1:0] node1021;
	wire [16-1:0] node1025;
	wire [16-1:0] node1026;
	wire [16-1:0] node1027;
	wire [16-1:0] node1030;
	wire [16-1:0] node1034;
	wire [16-1:0] node1035;
	wire [16-1:0] node1036;
	wire [16-1:0] node1038;
	wire [16-1:0] node1041;
	wire [16-1:0] node1042;
	wire [16-1:0] node1046;
	wire [16-1:0] node1047;
	wire [16-1:0] node1048;
	wire [16-1:0] node1050;
	wire [16-1:0] node1053;
	wire [16-1:0] node1055;
	wire [16-1:0] node1058;
	wire [16-1:0] node1060;
	wire [16-1:0] node1063;
	wire [16-1:0] node1064;
	wire [16-1:0] node1065;
	wire [16-1:0] node1066;
	wire [16-1:0] node1067;
	wire [16-1:0] node1070;
	wire [16-1:0] node1073;
	wire [16-1:0] node1074;
	wire [16-1:0] node1075;
	wire [16-1:0] node1077;
	wire [16-1:0] node1082;
	wire [16-1:0] node1083;
	wire [16-1:0] node1085;
	wire [16-1:0] node1088;
	wire [16-1:0] node1089;
	wire [16-1:0] node1092;
	wire [16-1:0] node1094;
	wire [16-1:0] node1095;
	wire [16-1:0] node1099;
	wire [16-1:0] node1100;
	wire [16-1:0] node1101;
	wire [16-1:0] node1103;
	wire [16-1:0] node1104;
	wire [16-1:0] node1108;
	wire [16-1:0] node1111;
	wire [16-1:0] node1112;
	wire [16-1:0] node1116;
	wire [16-1:0] node1117;
	wire [16-1:0] node1118;
	wire [16-1:0] node1119;
	wire [16-1:0] node1120;
	wire [16-1:0] node1121;
	wire [16-1:0] node1123;
	wire [16-1:0] node1126;
	wire [16-1:0] node1127;
	wire [16-1:0] node1128;
	wire [16-1:0] node1133;
	wire [16-1:0] node1134;
	wire [16-1:0] node1135;
	wire [16-1:0] node1136;
	wire [16-1:0] node1140;
	wire [16-1:0] node1141;
	wire [16-1:0] node1142;
	wire [16-1:0] node1146;
	wire [16-1:0] node1149;
	wire [16-1:0] node1152;
	wire [16-1:0] node1153;
	wire [16-1:0] node1154;
	wire [16-1:0] node1155;
	wire [16-1:0] node1158;
	wire [16-1:0] node1159;
	wire [16-1:0] node1160;
	wire [16-1:0] node1165;
	wire [16-1:0] node1166;
	wire [16-1:0] node1167;
	wire [16-1:0] node1168;
	wire [16-1:0] node1173;
	wire [16-1:0] node1176;
	wire [16-1:0] node1177;
	wire [16-1:0] node1179;
	wire [16-1:0] node1180;
	wire [16-1:0] node1184;
	wire [16-1:0] node1185;
	wire [16-1:0] node1187;
	wire [16-1:0] node1190;
	wire [16-1:0] node1191;
	wire [16-1:0] node1195;
	wire [16-1:0] node1196;
	wire [16-1:0] node1197;
	wire [16-1:0] node1198;
	wire [16-1:0] node1199;
	wire [16-1:0] node1202;
	wire [16-1:0] node1204;
	wire [16-1:0] node1207;
	wire [16-1:0] node1208;
	wire [16-1:0] node1209;
	wire [16-1:0] node1213;
	wire [16-1:0] node1214;
	wire [16-1:0] node1218;
	wire [16-1:0] node1219;
	wire [16-1:0] node1220;
	wire [16-1:0] node1223;
	wire [16-1:0] node1224;
	wire [16-1:0] node1228;
	wire [16-1:0] node1230;
	wire [16-1:0] node1232;
	wire [16-1:0] node1235;
	wire [16-1:0] node1236;
	wire [16-1:0] node1237;
	wire [16-1:0] node1238;
	wire [16-1:0] node1240;
	wire [16-1:0] node1241;
	wire [16-1:0] node1243;
	wire [16-1:0] node1247;
	wire [16-1:0] node1249;
	wire [16-1:0] node1252;
	wire [16-1:0] node1253;
	wire [16-1:0] node1254;
	wire [16-1:0] node1258;
	wire [16-1:0] node1260;
	wire [16-1:0] node1261;
	wire [16-1:0] node1265;
	wire [16-1:0] node1266;
	wire [16-1:0] node1267;
	wire [16-1:0] node1269;
	wire [16-1:0] node1272;
	wire [16-1:0] node1273;
	wire [16-1:0] node1277;
	wire [16-1:0] node1278;
	wire [16-1:0] node1280;
	wire [16-1:0] node1283;
	wire [16-1:0] node1285;
	wire [16-1:0] node1288;
	wire [16-1:0] node1289;
	wire [16-1:0] node1290;
	wire [16-1:0] node1291;
	wire [16-1:0] node1292;
	wire [16-1:0] node1293;
	wire [16-1:0] node1294;
	wire [16-1:0] node1297;
	wire [16-1:0] node1301;
	wire [16-1:0] node1302;
	wire [16-1:0] node1305;
	wire [16-1:0] node1307;
	wire [16-1:0] node1310;
	wire [16-1:0] node1311;
	wire [16-1:0] node1312;
	wire [16-1:0] node1313;
	wire [16-1:0] node1316;
	wire [16-1:0] node1319;
	wire [16-1:0] node1320;
	wire [16-1:0] node1322;
	wire [16-1:0] node1326;
	wire [16-1:0] node1327;
	wire [16-1:0] node1329;
	wire [16-1:0] node1330;
	wire [16-1:0] node1334;
	wire [16-1:0] node1336;
	wire [16-1:0] node1338;
	wire [16-1:0] node1341;
	wire [16-1:0] node1342;
	wire [16-1:0] node1343;
	wire [16-1:0] node1344;
	wire [16-1:0] node1346;
	wire [16-1:0] node1349;
	wire [16-1:0] node1350;
	wire [16-1:0] node1353;
	wire [16-1:0] node1355;
	wire [16-1:0] node1358;
	wire [16-1:0] node1359;
	wire [16-1:0] node1363;
	wire [16-1:0] node1364;
	wire [16-1:0] node1366;
	wire [16-1:0] node1367;
	wire [16-1:0] node1371;
	wire [16-1:0] node1373;
	wire [16-1:0] node1374;
	wire [16-1:0] node1376;
	wire [16-1:0] node1377;
	wire [16-1:0] node1382;
	wire [16-1:0] node1383;
	wire [16-1:0] node1384;
	wire [16-1:0] node1385;
	wire [16-1:0] node1386;
	wire [16-1:0] node1387;
	wire [16-1:0] node1390;
	wire [16-1:0] node1391;
	wire [16-1:0] node1396;
	wire [16-1:0] node1397;
	wire [16-1:0] node1398;
	wire [16-1:0] node1401;
	wire [16-1:0] node1404;
	wire [16-1:0] node1405;
	wire [16-1:0] node1407;
	wire [16-1:0] node1408;
	wire [16-1:0] node1413;
	wire [16-1:0] node1414;
	wire [16-1:0] node1415;
	wire [16-1:0] node1416;
	wire [16-1:0] node1419;
	wire [16-1:0] node1422;
	wire [16-1:0] node1423;
	wire [16-1:0] node1425;
	wire [16-1:0] node1428;
	wire [16-1:0] node1431;
	wire [16-1:0] node1432;
	wire [16-1:0] node1434;
	wire [16-1:0] node1437;
	wire [16-1:0] node1439;
	wire [16-1:0] node1442;
	wire [16-1:0] node1443;
	wire [16-1:0] node1444;
	wire [16-1:0] node1445;
	wire [16-1:0] node1449;
	wire [16-1:0] node1450;
	wire [16-1:0] node1451;
	wire [16-1:0] node1452;
	wire [16-1:0] node1456;
	wire [16-1:0] node1460;
	wire [16-1:0] node1461;
	wire [16-1:0] node1462;
	wire [16-1:0] node1464;
	wire [16-1:0] node1465;
	wire [16-1:0] node1467;
	wire [16-1:0] node1472;
	wire [16-1:0] node1474;
	wire [16-1:0] node1475;
	wire [16-1:0] node1479;
	wire [16-1:0] node1480;
	wire [16-1:0] node1481;
	wire [16-1:0] node1482;
	wire [16-1:0] node1483;
	wire [16-1:0] node1484;
	wire [16-1:0] node1485;
	wire [16-1:0] node1486;
	wire [16-1:0] node1487;
	wire [16-1:0] node1489;
	wire [16-1:0] node1490;
	wire [16-1:0] node1494;
	wire [16-1:0] node1495;
	wire [16-1:0] node1499;
	wire [16-1:0] node1500;
	wire [16-1:0] node1502;
	wire [16-1:0] node1504;
	wire [16-1:0] node1508;
	wire [16-1:0] node1509;
	wire [16-1:0] node1510;
	wire [16-1:0] node1511;
	wire [16-1:0] node1516;
	wire [16-1:0] node1519;
	wire [16-1:0] node1520;
	wire [16-1:0] node1521;
	wire [16-1:0] node1522;
	wire [16-1:0] node1523;
	wire [16-1:0] node1527;
	wire [16-1:0] node1528;
	wire [16-1:0] node1529;
	wire [16-1:0] node1530;
	wire [16-1:0] node1535;
	wire [16-1:0] node1538;
	wire [16-1:0] node1539;
	wire [16-1:0] node1543;
	wire [16-1:0] node1544;
	wire [16-1:0] node1545;
	wire [16-1:0] node1546;
	wire [16-1:0] node1551;
	wire [16-1:0] node1552;
	wire [16-1:0] node1553;
	wire [16-1:0] node1557;
	wire [16-1:0] node1559;
	wire [16-1:0] node1562;
	wire [16-1:0] node1563;
	wire [16-1:0] node1564;
	wire [16-1:0] node1565;
	wire [16-1:0] node1567;
	wire [16-1:0] node1568;
	wire [16-1:0] node1569;
	wire [16-1:0] node1571;
	wire [16-1:0] node1576;
	wire [16-1:0] node1577;
	wire [16-1:0] node1580;
	wire [16-1:0] node1583;
	wire [16-1:0] node1584;
	wire [16-1:0] node1586;
	wire [16-1:0] node1588;
	wire [16-1:0] node1591;
	wire [16-1:0] node1592;
	wire [16-1:0] node1593;
	wire [16-1:0] node1595;
	wire [16-1:0] node1596;
	wire [16-1:0] node1599;
	wire [16-1:0] node1603;
	wire [16-1:0] node1604;
	wire [16-1:0] node1607;
	wire [16-1:0] node1610;
	wire [16-1:0] node1611;
	wire [16-1:0] node1612;
	wire [16-1:0] node1613;
	wire [16-1:0] node1615;
	wire [16-1:0] node1617;
	wire [16-1:0] node1621;
	wire [16-1:0] node1622;
	wire [16-1:0] node1623;
	wire [16-1:0] node1625;
	wire [16-1:0] node1628;
	wire [16-1:0] node1631;
	wire [16-1:0] node1632;
	wire [16-1:0] node1634;
	wire [16-1:0] node1637;
	wire [16-1:0] node1640;
	wire [16-1:0] node1641;
	wire [16-1:0] node1643;
	wire [16-1:0] node1647;
	wire [16-1:0] node1648;
	wire [16-1:0] node1649;
	wire [16-1:0] node1650;
	wire [16-1:0] node1651;
	wire [16-1:0] node1652;
	wire [16-1:0] node1653;
	wire [16-1:0] node1656;
	wire [16-1:0] node1658;
	wire [16-1:0] node1661;
	wire [16-1:0] node1662;
	wire [16-1:0] node1664;
	wire [16-1:0] node1665;
	wire [16-1:0] node1669;
	wire [16-1:0] node1671;
	wire [16-1:0] node1674;
	wire [16-1:0] node1676;
	wire [16-1:0] node1679;
	wire [16-1:0] node1680;
	wire [16-1:0] node1681;
	wire [16-1:0] node1682;
	wire [16-1:0] node1686;
	wire [16-1:0] node1687;
	wire [16-1:0] node1690;
	wire [16-1:0] node1692;
	wire [16-1:0] node1695;
	wire [16-1:0] node1696;
	wire [16-1:0] node1698;
	wire [16-1:0] node1699;
	wire [16-1:0] node1704;
	wire [16-1:0] node1705;
	wire [16-1:0] node1706;
	wire [16-1:0] node1708;
	wire [16-1:0] node1709;
	wire [16-1:0] node1710;
	wire [16-1:0] node1714;
	wire [16-1:0] node1717;
	wire [16-1:0] node1718;
	wire [16-1:0] node1719;
	wire [16-1:0] node1723;
	wire [16-1:0] node1725;
	wire [16-1:0] node1728;
	wire [16-1:0] node1729;
	wire [16-1:0] node1731;
	wire [16-1:0] node1734;
	wire [16-1:0] node1735;
	wire [16-1:0] node1736;
	wire [16-1:0] node1740;
	wire [16-1:0] node1742;
	wire [16-1:0] node1743;
	wire [16-1:0] node1745;
	wire [16-1:0] node1749;
	wire [16-1:0] node1750;
	wire [16-1:0] node1751;
	wire [16-1:0] node1752;
	wire [16-1:0] node1753;
	wire [16-1:0] node1755;
	wire [16-1:0] node1756;
	wire [16-1:0] node1760;
	wire [16-1:0] node1762;
	wire [16-1:0] node1763;
	wire [16-1:0] node1767;
	wire [16-1:0] node1768;
	wire [16-1:0] node1769;
	wire [16-1:0] node1773;
	wire [16-1:0] node1774;
	wire [16-1:0] node1777;
	wire [16-1:0] node1780;
	wire [16-1:0] node1781;
	wire [16-1:0] node1782;
	wire [16-1:0] node1783;
	wire [16-1:0] node1787;
	wire [16-1:0] node1789;
	wire [16-1:0] node1792;
	wire [16-1:0] node1793;
	wire [16-1:0] node1794;
	wire [16-1:0] node1797;
	wire [16-1:0] node1800;
	wire [16-1:0] node1801;
	wire [16-1:0] node1805;
	wire [16-1:0] node1806;
	wire [16-1:0] node1807;
	wire [16-1:0] node1808;
	wire [16-1:0] node1810;
	wire [16-1:0] node1813;
	wire [16-1:0] node1815;
	wire [16-1:0] node1818;
	wire [16-1:0] node1819;
	wire [16-1:0] node1820;
	wire [16-1:0] node1823;
	wire [16-1:0] node1827;
	wire [16-1:0] node1828;
	wire [16-1:0] node1829;
	wire [16-1:0] node1831;
	wire [16-1:0] node1834;
	wire [16-1:0] node1836;
	wire [16-1:0] node1838;
	wire [16-1:0] node1841;
	wire [16-1:0] node1842;
	wire [16-1:0] node1843;
	wire [16-1:0] node1846;
	wire [16-1:0] node1849;
	wire [16-1:0] node1850;
	wire [16-1:0] node1851;
	wire [16-1:0] node1855;
	wire [16-1:0] node1858;
	wire [16-1:0] node1859;
	wire [16-1:0] node1860;
	wire [16-1:0] node1861;
	wire [16-1:0] node1862;
	wire [16-1:0] node1863;
	wire [16-1:0] node1864;
	wire [16-1:0] node1865;
	wire [16-1:0] node1866;
	wire [16-1:0] node1869;
	wire [16-1:0] node1873;
	wire [16-1:0] node1876;
	wire [16-1:0] node1877;
	wire [16-1:0] node1878;
	wire [16-1:0] node1882;
	wire [16-1:0] node1884;
	wire [16-1:0] node1887;
	wire [16-1:0] node1888;
	wire [16-1:0] node1889;
	wire [16-1:0] node1891;
	wire [16-1:0] node1892;
	wire [16-1:0] node1896;
	wire [16-1:0] node1897;
	wire [16-1:0] node1901;
	wire [16-1:0] node1903;
	wire [16-1:0] node1904;
	wire [16-1:0] node1908;
	wire [16-1:0] node1909;
	wire [16-1:0] node1910;
	wire [16-1:0] node1911;
	wire [16-1:0] node1913;
	wire [16-1:0] node1916;
	wire [16-1:0] node1917;
	wire [16-1:0] node1921;
	wire [16-1:0] node1922;
	wire [16-1:0] node1925;
	wire [16-1:0] node1927;
	wire [16-1:0] node1930;
	wire [16-1:0] node1931;
	wire [16-1:0] node1933;
	wire [16-1:0] node1934;
	wire [16-1:0] node1936;
	wire [16-1:0] node1939;
	wire [16-1:0] node1941;
	wire [16-1:0] node1942;
	wire [16-1:0] node1946;
	wire [16-1:0] node1947;
	wire [16-1:0] node1948;
	wire [16-1:0] node1951;
	wire [16-1:0] node1953;
	wire [16-1:0] node1956;
	wire [16-1:0] node1958;
	wire [16-1:0] node1960;
	wire [16-1:0] node1963;
	wire [16-1:0] node1964;
	wire [16-1:0] node1965;
	wire [16-1:0] node1966;
	wire [16-1:0] node1967;
	wire [16-1:0] node1970;
	wire [16-1:0] node1971;
	wire [16-1:0] node1975;
	wire [16-1:0] node1977;
	wire [16-1:0] node1978;
	wire [16-1:0] node1982;
	wire [16-1:0] node1983;
	wire [16-1:0] node1984;
	wire [16-1:0] node1986;
	wire [16-1:0] node1989;
	wire [16-1:0] node1990;
	wire [16-1:0] node1994;
	wire [16-1:0] node1995;
	wire [16-1:0] node1997;
	wire [16-1:0] node1999;
	wire [16-1:0] node2000;
	wire [16-1:0] node2005;
	wire [16-1:0] node2006;
	wire [16-1:0] node2007;
	wire [16-1:0] node2008;
	wire [16-1:0] node2009;
	wire [16-1:0] node2011;
	wire [16-1:0] node2013;
	wire [16-1:0] node2017;
	wire [16-1:0] node2020;
	wire [16-1:0] node2022;
	wire [16-1:0] node2023;
	wire [16-1:0] node2025;
	wire [16-1:0] node2029;
	wire [16-1:0] node2030;
	wire [16-1:0] node2031;
	wire [16-1:0] node2032;
	wire [16-1:0] node2036;
	wire [16-1:0] node2037;
	wire [16-1:0] node2039;
	wire [16-1:0] node2040;
	wire [16-1:0] node2045;
	wire [16-1:0] node2047;
	wire [16-1:0] node2050;
	wire [16-1:0] node2051;
	wire [16-1:0] node2052;
	wire [16-1:0] node2053;
	wire [16-1:0] node2054;
	wire [16-1:0] node2055;
	wire [16-1:0] node2056;
	wire [16-1:0] node2057;
	wire [16-1:0] node2062;
	wire [16-1:0] node2063;
	wire [16-1:0] node2067;
	wire [16-1:0] node2068;
	wire [16-1:0] node2069;
	wire [16-1:0] node2073;
	wire [16-1:0] node2074;
	wire [16-1:0] node2078;
	wire [16-1:0] node2079;
	wire [16-1:0] node2080;
	wire [16-1:0] node2083;
	wire [16-1:0] node2084;
	wire [16-1:0] node2088;
	wire [16-1:0] node2089;
	wire [16-1:0] node2091;
	wire [16-1:0] node2094;
	wire [16-1:0] node2095;
	wire [16-1:0] node2099;
	wire [16-1:0] node2100;
	wire [16-1:0] node2101;
	wire [16-1:0] node2102;
	wire [16-1:0] node2103;
	wire [16-1:0] node2106;
	wire [16-1:0] node2109;
	wire [16-1:0] node2110;
	wire [16-1:0] node2113;
	wire [16-1:0] node2116;
	wire [16-1:0] node2117;
	wire [16-1:0] node2118;
	wire [16-1:0] node2121;
	wire [16-1:0] node2124;
	wire [16-1:0] node2125;
	wire [16-1:0] node2127;
	wire [16-1:0] node2130;
	wire [16-1:0] node2133;
	wire [16-1:0] node2134;
	wire [16-1:0] node2135;
	wire [16-1:0] node2136;
	wire [16-1:0] node2139;
	wire [16-1:0] node2142;
	wire [16-1:0] node2143;
	wire [16-1:0] node2146;
	wire [16-1:0] node2148;
	wire [16-1:0] node2151;
	wire [16-1:0] node2152;
	wire [16-1:0] node2156;
	wire [16-1:0] node2157;
	wire [16-1:0] node2158;
	wire [16-1:0] node2159;
	wire [16-1:0] node2160;
	wire [16-1:0] node2161;
	wire [16-1:0] node2162;
	wire [16-1:0] node2165;
	wire [16-1:0] node2170;
	wire [16-1:0] node2171;
	wire [16-1:0] node2172;
	wire [16-1:0] node2173;
	wire [16-1:0] node2177;
	wire [16-1:0] node2180;
	wire [16-1:0] node2181;
	wire [16-1:0] node2185;
	wire [16-1:0] node2186;
	wire [16-1:0] node2187;
	wire [16-1:0] node2191;
	wire [16-1:0] node2192;
	wire [16-1:0] node2194;
	wire [16-1:0] node2197;
	wire [16-1:0] node2198;
	wire [16-1:0] node2202;
	wire [16-1:0] node2203;
	wire [16-1:0] node2204;
	wire [16-1:0] node2205;
	wire [16-1:0] node2207;
	wire [16-1:0] node2210;
	wire [16-1:0] node2211;
	wire [16-1:0] node2213;
	wire [16-1:0] node2216;
	wire [16-1:0] node2217;
	wire [16-1:0] node2221;
	wire [16-1:0] node2222;
	wire [16-1:0] node2224;
	wire [16-1:0] node2227;
	wire [16-1:0] node2229;
	wire [16-1:0] node2230;
	wire [16-1:0] node2234;
	wire [16-1:0] node2235;
	wire [16-1:0] node2236;
	wire [16-1:0] node2238;
	wire [16-1:0] node2240;
	wire [16-1:0] node2243;
	wire [16-1:0] node2246;
	wire [16-1:0] node2247;
	wire [16-1:0] node2249;
	wire [16-1:0] node2252;
	wire [16-1:0] node2254;
	wire [16-1:0] node2255;
	wire [16-1:0] node2259;
	wire [16-1:0] node2260;
	wire [16-1:0] node2261;
	wire [16-1:0] node2262;
	wire [16-1:0] node2263;
	wire [16-1:0] node2264;
	wire [16-1:0] node2265;
	wire [16-1:0] node2266;
	wire [16-1:0] node2269;
	wire [16-1:0] node2270;
	wire [16-1:0] node2272;
	wire [16-1:0] node2275;
	wire [16-1:0] node2278;
	wire [16-1:0] node2280;
	wire [16-1:0] node2281;
	wire [16-1:0] node2285;
	wire [16-1:0] node2286;
	wire [16-1:0] node2287;
	wire [16-1:0] node2291;
	wire [16-1:0] node2293;
	wire [16-1:0] node2296;
	wire [16-1:0] node2297;
	wire [16-1:0] node2298;
	wire [16-1:0] node2300;
	wire [16-1:0] node2301;
	wire [16-1:0] node2302;
	wire [16-1:0] node2307;
	wire [16-1:0] node2308;
	wire [16-1:0] node2310;
	wire [16-1:0] node2313;
	wire [16-1:0] node2314;
	wire [16-1:0] node2315;
	wire [16-1:0] node2320;
	wire [16-1:0] node2321;
	wire [16-1:0] node2322;
	wire [16-1:0] node2323;
	wire [16-1:0] node2324;
	wire [16-1:0] node2328;
	wire [16-1:0] node2329;
	wire [16-1:0] node2333;
	wire [16-1:0] node2334;
	wire [16-1:0] node2335;
	wire [16-1:0] node2339;
	wire [16-1:0] node2342;
	wire [16-1:0] node2344;
	wire [16-1:0] node2347;
	wire [16-1:0] node2348;
	wire [16-1:0] node2349;
	wire [16-1:0] node2350;
	wire [16-1:0] node2351;
	wire [16-1:0] node2355;
	wire [16-1:0] node2356;
	wire [16-1:0] node2357;
	wire [16-1:0] node2360;
	wire [16-1:0] node2363;
	wire [16-1:0] node2364;
	wire [16-1:0] node2365;
	wire [16-1:0] node2370;
	wire [16-1:0] node2371;
	wire [16-1:0] node2373;
	wire [16-1:0] node2374;
	wire [16-1:0] node2378;
	wire [16-1:0] node2379;
	wire [16-1:0] node2381;
	wire [16-1:0] node2384;
	wire [16-1:0] node2387;
	wire [16-1:0] node2388;
	wire [16-1:0] node2389;
	wire [16-1:0] node2391;
	wire [16-1:0] node2392;
	wire [16-1:0] node2395;
	wire [16-1:0] node2397;
	wire [16-1:0] node2400;
	wire [16-1:0] node2401;
	wire [16-1:0] node2403;
	wire [16-1:0] node2406;
	wire [16-1:0] node2408;
	wire [16-1:0] node2411;
	wire [16-1:0] node2412;
	wire [16-1:0] node2413;
	wire [16-1:0] node2416;
	wire [16-1:0] node2419;
	wire [16-1:0] node2420;
	wire [16-1:0] node2424;
	wire [16-1:0] node2425;
	wire [16-1:0] node2426;
	wire [16-1:0] node2427;
	wire [16-1:0] node2428;
	wire [16-1:0] node2429;
	wire [16-1:0] node2430;
	wire [16-1:0] node2434;
	wire [16-1:0] node2437;
	wire [16-1:0] node2439;
	wire [16-1:0] node2440;
	wire [16-1:0] node2441;
	wire [16-1:0] node2442;
	wire [16-1:0] node2448;
	wire [16-1:0] node2449;
	wire [16-1:0] node2450;
	wire [16-1:0] node2451;
	wire [16-1:0] node2455;
	wire [16-1:0] node2456;
	wire [16-1:0] node2460;
	wire [16-1:0] node2462;
	wire [16-1:0] node2464;
	wire [16-1:0] node2467;
	wire [16-1:0] node2468;
	wire [16-1:0] node2469;
	wire [16-1:0] node2470;
	wire [16-1:0] node2471;
	wire [16-1:0] node2472;
	wire [16-1:0] node2476;
	wire [16-1:0] node2479;
	wire [16-1:0] node2482;
	wire [16-1:0] node2483;
	wire [16-1:0] node2484;
	wire [16-1:0] node2487;
	wire [16-1:0] node2490;
	wire [16-1:0] node2491;
	wire [16-1:0] node2495;
	wire [16-1:0] node2496;
	wire [16-1:0] node2497;
	wire [16-1:0] node2501;
	wire [16-1:0] node2502;
	wire [16-1:0] node2504;
	wire [16-1:0] node2508;
	wire [16-1:0] node2509;
	wire [16-1:0] node2510;
	wire [16-1:0] node2511;
	wire [16-1:0] node2512;
	wire [16-1:0] node2514;
	wire [16-1:0] node2516;
	wire [16-1:0] node2520;
	wire [16-1:0] node2522;
	wire [16-1:0] node2523;
	wire [16-1:0] node2527;
	wire [16-1:0] node2528;
	wire [16-1:0] node2529;
	wire [16-1:0] node2530;
	wire [16-1:0] node2533;
	wire [16-1:0] node2536;
	wire [16-1:0] node2537;
	wire [16-1:0] node2539;
	wire [16-1:0] node2540;
	wire [16-1:0] node2545;
	wire [16-1:0] node2546;
	wire [16-1:0] node2547;
	wire [16-1:0] node2550;
	wire [16-1:0] node2553;
	wire [16-1:0] node2554;
	wire [16-1:0] node2557;
	wire [16-1:0] node2560;
	wire [16-1:0] node2561;
	wire [16-1:0] node2562;
	wire [16-1:0] node2564;
	wire [16-1:0] node2565;
	wire [16-1:0] node2566;
	wire [16-1:0] node2571;
	wire [16-1:0] node2573;
	wire [16-1:0] node2574;
	wire [16-1:0] node2577;
	wire [16-1:0] node2579;
	wire [16-1:0] node2582;
	wire [16-1:0] node2583;
	wire [16-1:0] node2584;
	wire [16-1:0] node2586;
	wire [16-1:0] node2590;
	wire [16-1:0] node2591;
	wire [16-1:0] node2593;
	wire [16-1:0] node2596;
	wire [16-1:0] node2597;
	wire [16-1:0] node2601;
	wire [16-1:0] node2602;
	wire [16-1:0] node2603;
	wire [16-1:0] node2604;
	wire [16-1:0] node2605;
	wire [16-1:0] node2606;
	wire [16-1:0] node2607;
	wire [16-1:0] node2608;
	wire [16-1:0] node2609;
	wire [16-1:0] node2614;
	wire [16-1:0] node2617;
	wire [16-1:0] node2619;
	wire [16-1:0] node2620;
	wire [16-1:0] node2621;
	wire [16-1:0] node2622;
	wire [16-1:0] node2628;
	wire [16-1:0] node2629;
	wire [16-1:0] node2630;
	wire [16-1:0] node2633;
	wire [16-1:0] node2634;
	wire [16-1:0] node2638;
	wire [16-1:0] node2639;
	wire [16-1:0] node2640;
	wire [16-1:0] node2644;
	wire [16-1:0] node2645;
	wire [16-1:0] node2649;
	wire [16-1:0] node2650;
	wire [16-1:0] node2651;
	wire [16-1:0] node2652;
	wire [16-1:0] node2653;
	wire [16-1:0] node2657;
	wire [16-1:0] node2659;
	wire [16-1:0] node2662;
	wire [16-1:0] node2663;
	wire [16-1:0] node2667;
	wire [16-1:0] node2668;
	wire [16-1:0] node2669;
	wire [16-1:0] node2671;
	wire [16-1:0] node2673;
	wire [16-1:0] node2676;
	wire [16-1:0] node2677;
	wire [16-1:0] node2678;
	wire [16-1:0] node2683;
	wire [16-1:0] node2684;
	wire [16-1:0] node2686;
	wire [16-1:0] node2690;
	wire [16-1:0] node2691;
	wire [16-1:0] node2692;
	wire [16-1:0] node2693;
	wire [16-1:0] node2695;
	wire [16-1:0] node2696;
	wire [16-1:0] node2700;
	wire [16-1:0] node2701;
	wire [16-1:0] node2702;
	wire [16-1:0] node2707;
	wire [16-1:0] node2708;
	wire [16-1:0] node2709;
	wire [16-1:0] node2711;
	wire [16-1:0] node2715;
	wire [16-1:0] node2717;
	wire [16-1:0] node2718;
	wire [16-1:0] node2722;
	wire [16-1:0] node2723;
	wire [16-1:0] node2724;
	wire [16-1:0] node2725;
	wire [16-1:0] node2726;
	wire [16-1:0] node2730;
	wire [16-1:0] node2732;
	wire [16-1:0] node2735;
	wire [16-1:0] node2736;
	wire [16-1:0] node2737;
	wire [16-1:0] node2738;
	wire [16-1:0] node2740;
	wire [16-1:0] node2745;
	wire [16-1:0] node2746;
	wire [16-1:0] node2748;
	wire [16-1:0] node2749;
	wire [16-1:0] node2753;
	wire [16-1:0] node2756;
	wire [16-1:0] node2757;
	wire [16-1:0] node2758;
	wire [16-1:0] node2760;
	wire [16-1:0] node2764;
	wire [16-1:0] node2765;
	wire [16-1:0] node2766;
	wire [16-1:0] node2769;
	wire [16-1:0] node2771;
	wire [16-1:0] node2772;
	wire [16-1:0] node2776;
	wire [16-1:0] node2777;
	wire [16-1:0] node2778;
	wire [16-1:0] node2783;
	wire [16-1:0] node2784;
	wire [16-1:0] node2785;
	wire [16-1:0] node2786;
	wire [16-1:0] node2787;
	wire [16-1:0] node2788;
	wire [16-1:0] node2791;
	wire [16-1:0] node2794;
	wire [16-1:0] node2795;
	wire [16-1:0] node2797;
	wire [16-1:0] node2800;
	wire [16-1:0] node2803;
	wire [16-1:0] node2804;
	wire [16-1:0] node2805;
	wire [16-1:0] node2808;
	wire [16-1:0] node2810;
	wire [16-1:0] node2813;
	wire [16-1:0] node2815;
	wire [16-1:0] node2818;
	wire [16-1:0] node2819;
	wire [16-1:0] node2820;
	wire [16-1:0] node2821;
	wire [16-1:0] node2822;
	wire [16-1:0] node2826;
	wire [16-1:0] node2827;
	wire [16-1:0] node2831;
	wire [16-1:0] node2832;
	wire [16-1:0] node2833;
	wire [16-1:0] node2836;
	wire [16-1:0] node2838;
	wire [16-1:0] node2841;
	wire [16-1:0] node2843;
	wire [16-1:0] node2846;
	wire [16-1:0] node2847;
	wire [16-1:0] node2849;
	wire [16-1:0] node2850;
	wire [16-1:0] node2851;
	wire [16-1:0] node2855;
	wire [16-1:0] node2858;
	wire [16-1:0] node2859;
	wire [16-1:0] node2861;
	wire [16-1:0] node2865;
	wire [16-1:0] node2866;
	wire [16-1:0] node2867;
	wire [16-1:0] node2868;
	wire [16-1:0] node2869;
	wire [16-1:0] node2871;
	wire [16-1:0] node2874;
	wire [16-1:0] node2876;
	wire [16-1:0] node2879;
	wire [16-1:0] node2882;
	wire [16-1:0] node2883;
	wire [16-1:0] node2884;
	wire [16-1:0] node2886;
	wire [16-1:0] node2887;
	wire [16-1:0] node2889;
	wire [16-1:0] node2894;
	wire [16-1:0] node2895;
	wire [16-1:0] node2898;
	wire [16-1:0] node2899;
	wire [16-1:0] node2903;
	wire [16-1:0] node2904;
	wire [16-1:0] node2905;
	wire [16-1:0] node2906;
	wire [16-1:0] node2907;
	wire [16-1:0] node2911;
	wire [16-1:0] node2913;
	wire [16-1:0] node2914;
	wire [16-1:0] node2918;
	wire [16-1:0] node2919;
	wire [16-1:0] node2921;
	wire [16-1:0] node2922;
	wire [16-1:0] node2926;
	wire [16-1:0] node2928;
	wire [16-1:0] node2930;
	wire [16-1:0] node2933;
	wire [16-1:0] node2934;
	wire [16-1:0] node2935;
	wire [16-1:0] node2936;
	wire [16-1:0] node2941;
	wire [16-1:0] node2942;
	wire [16-1:0] node2943;
	wire [16-1:0] node2944;
	wire [16-1:0] node2947;
	wire [16-1:0] node2949;
	wire [16-1:0] node2952;
	wire [16-1:0] node2956;
	wire [16-1:0] node2957;
	wire [16-1:0] node2958;
	wire [16-1:0] node2959;
	wire [16-1:0] node2960;
	wire [16-1:0] node2961;
	wire [16-1:0] node2962;
	wire [16-1:0] node2963;
	wire [16-1:0] node2964;
	wire [16-1:0] node2965;
	wire [16-1:0] node2966;
	wire [16-1:0] node2971;
	wire [16-1:0] node2972;
	wire [16-1:0] node2973;
	wire [16-1:0] node2977;
	wire [16-1:0] node2979;
	wire [16-1:0] node2982;
	wire [16-1:0] node2983;
	wire [16-1:0] node2984;
	wire [16-1:0] node2985;
	wire [16-1:0] node2986;
	wire [16-1:0] node2990;
	wire [16-1:0] node2994;
	wire [16-1:0] node2995;
	wire [16-1:0] node2996;
	wire [16-1:0] node2998;
	wire [16-1:0] node3002;
	wire [16-1:0] node3004;
	wire [16-1:0] node3007;
	wire [16-1:0] node3008;
	wire [16-1:0] node3009;
	wire [16-1:0] node3010;
	wire [16-1:0] node3011;
	wire [16-1:0] node3013;
	wire [16-1:0] node3014;
	wire [16-1:0] node3018;
	wire [16-1:0] node3021;
	wire [16-1:0] node3022;
	wire [16-1:0] node3026;
	wire [16-1:0] node3028;
	wire [16-1:0] node3030;
	wire [16-1:0] node3033;
	wire [16-1:0] node3034;
	wire [16-1:0] node3036;
	wire [16-1:0] node3037;
	wire [16-1:0] node3041;
	wire [16-1:0] node3042;
	wire [16-1:0] node3044;
	wire [16-1:0] node3047;
	wire [16-1:0] node3048;
	wire [16-1:0] node3052;
	wire [16-1:0] node3053;
	wire [16-1:0] node3054;
	wire [16-1:0] node3055;
	wire [16-1:0] node3056;
	wire [16-1:0] node3057;
	wire [16-1:0] node3058;
	wire [16-1:0] node3062;
	wire [16-1:0] node3065;
	wire [16-1:0] node3066;
	wire [16-1:0] node3070;
	wire [16-1:0] node3071;
	wire [16-1:0] node3073;
	wire [16-1:0] node3076;
	wire [16-1:0] node3077;
	wire [16-1:0] node3079;
	wire [16-1:0] node3082;
	wire [16-1:0] node3083;
	wire [16-1:0] node3084;
	wire [16-1:0] node3089;
	wire [16-1:0] node3090;
	wire [16-1:0] node3091;
	wire [16-1:0] node3095;
	wire [16-1:0] node3097;
	wire [16-1:0] node3100;
	wire [16-1:0] node3101;
	wire [16-1:0] node3102;
	wire [16-1:0] node3103;
	wire [16-1:0] node3104;
	wire [16-1:0] node3108;
	wire [16-1:0] node3110;
	wire [16-1:0] node3113;
	wire [16-1:0] node3114;
	wire [16-1:0] node3116;
	wire [16-1:0] node3120;
	wire [16-1:0] node3121;
	wire [16-1:0] node3122;
	wire [16-1:0] node3123;
	wire [16-1:0] node3125;
	wire [16-1:0] node3129;
	wire [16-1:0] node3131;
	wire [16-1:0] node3132;
	wire [16-1:0] node3134;
	wire [16-1:0] node3138;
	wire [16-1:0] node3140;
	wire [16-1:0] node3141;
	wire [16-1:0] node3143;
	wire [16-1:0] node3147;
	wire [16-1:0] node3148;
	wire [16-1:0] node3149;
	wire [16-1:0] node3150;
	wire [16-1:0] node3151;
	wire [16-1:0] node3152;
	wire [16-1:0] node3154;
	wire [16-1:0] node3156;
	wire [16-1:0] node3157;
	wire [16-1:0] node3161;
	wire [16-1:0] node3162;
	wire [16-1:0] node3166;
	wire [16-1:0] node3167;
	wire [16-1:0] node3169;
	wire [16-1:0] node3172;
	wire [16-1:0] node3175;
	wire [16-1:0] node3176;
	wire [16-1:0] node3177;
	wire [16-1:0] node3179;
	wire [16-1:0] node3183;
	wire [16-1:0] node3185;
	wire [16-1:0] node3186;
	wire [16-1:0] node3187;
	wire [16-1:0] node3192;
	wire [16-1:0] node3193;
	wire [16-1:0] node3194;
	wire [16-1:0] node3195;
	wire [16-1:0] node3198;
	wire [16-1:0] node3199;
	wire [16-1:0] node3201;
	wire [16-1:0] node3205;
	wire [16-1:0] node3207;
	wire [16-1:0] node3208;
	wire [16-1:0] node3212;
	wire [16-1:0] node3213;
	wire [16-1:0] node3214;
	wire [16-1:0] node3216;
	wire [16-1:0] node3219;
	wire [16-1:0] node3220;
	wire [16-1:0] node3224;
	wire [16-1:0] node3225;
	wire [16-1:0] node3226;
	wire [16-1:0] node3227;
	wire [16-1:0] node3229;
	wire [16-1:0] node3232;
	wire [16-1:0] node3236;
	wire [16-1:0] node3237;
	wire [16-1:0] node3241;
	wire [16-1:0] node3242;
	wire [16-1:0] node3243;
	wire [16-1:0] node3244;
	wire [16-1:0] node3245;
	wire [16-1:0] node3246;
	wire [16-1:0] node3249;
	wire [16-1:0] node3252;
	wire [16-1:0] node3255;
	wire [16-1:0] node3256;
	wire [16-1:0] node3257;
	wire [16-1:0] node3260;
	wire [16-1:0] node3261;
	wire [16-1:0] node3266;
	wire [16-1:0] node3267;
	wire [16-1:0] node3268;
	wire [16-1:0] node3271;
	wire [16-1:0] node3273;
	wire [16-1:0] node3276;
	wire [16-1:0] node3278;
	wire [16-1:0] node3279;
	wire [16-1:0] node3282;
	wire [16-1:0] node3285;
	wire [16-1:0] node3286;
	wire [16-1:0] node3287;
	wire [16-1:0] node3288;
	wire [16-1:0] node3291;
	wire [16-1:0] node3292;
	wire [16-1:0] node3294;
	wire [16-1:0] node3298;
	wire [16-1:0] node3299;
	wire [16-1:0] node3300;
	wire [16-1:0] node3301;
	wire [16-1:0] node3303;
	wire [16-1:0] node3306;
	wire [16-1:0] node3307;
	wire [16-1:0] node3311;
	wire [16-1:0] node3314;
	wire [16-1:0] node3315;
	wire [16-1:0] node3318;
	wire [16-1:0] node3321;
	wire [16-1:0] node3322;
	wire [16-1:0] node3323;
	wire [16-1:0] node3327;
	wire [16-1:0] node3328;
	wire [16-1:0] node3330;
	wire [16-1:0] node3333;
	wire [16-1:0] node3335;
	wire [16-1:0] node3336;
	wire [16-1:0] node3340;
	wire [16-1:0] node3341;
	wire [16-1:0] node3342;
	wire [16-1:0] node3343;
	wire [16-1:0] node3344;
	wire [16-1:0] node3345;
	wire [16-1:0] node3347;
	wire [16-1:0] node3348;
	wire [16-1:0] node3350;
	wire [16-1:0] node3352;
	wire [16-1:0] node3356;
	wire [16-1:0] node3357;
	wire [16-1:0] node3358;
	wire [16-1:0] node3359;
	wire [16-1:0] node3365;
	wire [16-1:0] node3366;
	wire [16-1:0] node3368;
	wire [16-1:0] node3369;
	wire [16-1:0] node3373;
	wire [16-1:0] node3374;
	wire [16-1:0] node3376;
	wire [16-1:0] node3379;
	wire [16-1:0] node3382;
	wire [16-1:0] node3383;
	wire [16-1:0] node3384;
	wire [16-1:0] node3387;
	wire [16-1:0] node3388;
	wire [16-1:0] node3389;
	wire [16-1:0] node3393;
	wire [16-1:0] node3394;
	wire [16-1:0] node3398;
	wire [16-1:0] node3399;
	wire [16-1:0] node3400;
	wire [16-1:0] node3401;
	wire [16-1:0] node3404;
	wire [16-1:0] node3407;
	wire [16-1:0] node3408;
	wire [16-1:0] node3411;
	wire [16-1:0] node3414;
	wire [16-1:0] node3415;
	wire [16-1:0] node3416;
	wire [16-1:0] node3420;
	wire [16-1:0] node3422;
	wire [16-1:0] node3425;
	wire [16-1:0] node3426;
	wire [16-1:0] node3427;
	wire [16-1:0] node3428;
	wire [16-1:0] node3429;
	wire [16-1:0] node3430;
	wire [16-1:0] node3434;
	wire [16-1:0] node3436;
	wire [16-1:0] node3439;
	wire [16-1:0] node3441;
	wire [16-1:0] node3444;
	wire [16-1:0] node3445;
	wire [16-1:0] node3446;
	wire [16-1:0] node3448;
	wire [16-1:0] node3449;
	wire [16-1:0] node3450;
	wire [16-1:0] node3455;
	wire [16-1:0] node3457;
	wire [16-1:0] node3459;
	wire [16-1:0] node3460;
	wire [16-1:0] node3464;
	wire [16-1:0] node3466;
	wire [16-1:0] node3469;
	wire [16-1:0] node3470;
	wire [16-1:0] node3471;
	wire [16-1:0] node3472;
	wire [16-1:0] node3473;
	wire [16-1:0] node3475;
	wire [16-1:0] node3480;
	wire [16-1:0] node3482;
	wire [16-1:0] node3483;
	wire [16-1:0] node3487;
	wire [16-1:0] node3488;
	wire [16-1:0] node3489;
	wire [16-1:0] node3491;
	wire [16-1:0] node3493;
	wire [16-1:0] node3497;
	wire [16-1:0] node3499;
	wire [16-1:0] node3500;
	wire [16-1:0] node3502;
	wire [16-1:0] node3506;
	wire [16-1:0] node3507;
	wire [16-1:0] node3508;
	wire [16-1:0] node3509;
	wire [16-1:0] node3510;
	wire [16-1:0] node3511;
	wire [16-1:0] node3512;
	wire [16-1:0] node3516;
	wire [16-1:0] node3518;
	wire [16-1:0] node3519;
	wire [16-1:0] node3521;
	wire [16-1:0] node3525;
	wire [16-1:0] node3526;
	wire [16-1:0] node3527;
	wire [16-1:0] node3532;
	wire [16-1:0] node3533;
	wire [16-1:0] node3534;
	wire [16-1:0] node3536;
	wire [16-1:0] node3539;
	wire [16-1:0] node3540;
	wire [16-1:0] node3542;
	wire [16-1:0] node3545;
	wire [16-1:0] node3547;
	wire [16-1:0] node3550;
	wire [16-1:0] node3551;
	wire [16-1:0] node3553;
	wire [16-1:0] node3555;
	wire [16-1:0] node3558;
	wire [16-1:0] node3560;
	wire [16-1:0] node3563;
	wire [16-1:0] node3564;
	wire [16-1:0] node3565;
	wire [16-1:0] node3568;
	wire [16-1:0] node3569;
	wire [16-1:0] node3571;
	wire [16-1:0] node3575;
	wire [16-1:0] node3576;
	wire [16-1:0] node3577;
	wire [16-1:0] node3578;
	wire [16-1:0] node3582;
	wire [16-1:0] node3584;
	wire [16-1:0] node3585;
	wire [16-1:0] node3589;
	wire [16-1:0] node3590;
	wire [16-1:0] node3594;
	wire [16-1:0] node3595;
	wire [16-1:0] node3596;
	wire [16-1:0] node3597;
	wire [16-1:0] node3598;
	wire [16-1:0] node3601;
	wire [16-1:0] node3602;
	wire [16-1:0] node3604;
	wire [16-1:0] node3608;
	wire [16-1:0] node3610;
	wire [16-1:0] node3611;
	wire [16-1:0] node3614;
	wire [16-1:0] node3617;
	wire [16-1:0] node3618;
	wire [16-1:0] node3619;
	wire [16-1:0] node3620;
	wire [16-1:0] node3622;
	wire [16-1:0] node3626;
	wire [16-1:0] node3628;
	wire [16-1:0] node3631;
	wire [16-1:0] node3632;
	wire [16-1:0] node3634;
	wire [16-1:0] node3635;
	wire [16-1:0] node3637;
	wire [16-1:0] node3642;
	wire [16-1:0] node3643;
	wire [16-1:0] node3644;
	wire [16-1:0] node3647;
	wire [16-1:0] node3648;
	wire [16-1:0] node3650;
	wire [16-1:0] node3653;
	wire [16-1:0] node3654;
	wire [16-1:0] node3655;
	wire [16-1:0] node3660;
	wire [16-1:0] node3661;
	wire [16-1:0] node3662;
	wire [16-1:0] node3664;
	wire [16-1:0] node3667;
	wire [16-1:0] node3670;
	wire [16-1:0] node3671;
	wire [16-1:0] node3673;
	wire [16-1:0] node3675;
	wire [16-1:0] node3678;
	wire [16-1:0] node3681;
	wire [16-1:0] node3682;
	wire [16-1:0] node3683;
	wire [16-1:0] node3684;
	wire [16-1:0] node3685;
	wire [16-1:0] node3686;
	wire [16-1:0] node3687;
	wire [16-1:0] node3688;
	wire [16-1:0] node3689;
	wire [16-1:0] node3691;
	wire [16-1:0] node3695;
	wire [16-1:0] node3696;
	wire [16-1:0] node3698;
	wire [16-1:0] node3699;
	wire [16-1:0] node3704;
	wire [16-1:0] node3705;
	wire [16-1:0] node3706;
	wire [16-1:0] node3709;
	wire [16-1:0] node3712;
	wire [16-1:0] node3713;
	wire [16-1:0] node3717;
	wire [16-1:0] node3718;
	wire [16-1:0] node3719;
	wire [16-1:0] node3722;
	wire [16-1:0] node3724;
	wire [16-1:0] node3727;
	wire [16-1:0] node3728;
	wire [16-1:0] node3729;
	wire [16-1:0] node3733;
	wire [16-1:0] node3734;
	wire [16-1:0] node3736;
	wire [16-1:0] node3737;
	wire [16-1:0] node3742;
	wire [16-1:0] node3743;
	wire [16-1:0] node3744;
	wire [16-1:0] node3745;
	wire [16-1:0] node3748;
	wire [16-1:0] node3751;
	wire [16-1:0] node3752;
	wire [16-1:0] node3753;
	wire [16-1:0] node3758;
	wire [16-1:0] node3759;
	wire [16-1:0] node3761;
	wire [16-1:0] node3764;
	wire [16-1:0] node3765;
	wire [16-1:0] node3766;
	wire [16-1:0] node3770;
	wire [16-1:0] node3771;
	wire [16-1:0] node3775;
	wire [16-1:0] node3776;
	wire [16-1:0] node3777;
	wire [16-1:0] node3778;
	wire [16-1:0] node3780;
	wire [16-1:0] node3781;
	wire [16-1:0] node3783;
	wire [16-1:0] node3787;
	wire [16-1:0] node3788;
	wire [16-1:0] node3790;
	wire [16-1:0] node3792;
	wire [16-1:0] node3795;
	wire [16-1:0] node3798;
	wire [16-1:0] node3799;
	wire [16-1:0] node3800;
	wire [16-1:0] node3803;
	wire [16-1:0] node3805;
	wire [16-1:0] node3808;
	wire [16-1:0] node3810;
	wire [16-1:0] node3812;
	wire [16-1:0] node3815;
	wire [16-1:0] node3816;
	wire [16-1:0] node3817;
	wire [16-1:0] node3818;
	wire [16-1:0] node3820;
	wire [16-1:0] node3824;
	wire [16-1:0] node3825;
	wire [16-1:0] node3827;
	wire [16-1:0] node3831;
	wire [16-1:0] node3832;
	wire [16-1:0] node3833;
	wire [16-1:0] node3834;
	wire [16-1:0] node3839;
	wire [16-1:0] node3840;
	wire [16-1:0] node3842;
	wire [16-1:0] node3845;
	wire [16-1:0] node3847;
	wire [16-1:0] node3850;
	wire [16-1:0] node3851;
	wire [16-1:0] node3852;
	wire [16-1:0] node3853;
	wire [16-1:0] node3854;
	wire [16-1:0] node3855;
	wire [16-1:0] node3856;
	wire [16-1:0] node3857;
	wire [16-1:0] node3859;
	wire [16-1:0] node3864;
	wire [16-1:0] node3867;
	wire [16-1:0] node3868;
	wire [16-1:0] node3869;
	wire [16-1:0] node3871;
	wire [16-1:0] node3875;
	wire [16-1:0] node3876;
	wire [16-1:0] node3880;
	wire [16-1:0] node3881;
	wire [16-1:0] node3882;
	wire [16-1:0] node3885;
	wire [16-1:0] node3887;
	wire [16-1:0] node3889;
	wire [16-1:0] node3892;
	wire [16-1:0] node3894;
	wire [16-1:0] node3896;
	wire [16-1:0] node3899;
	wire [16-1:0] node3900;
	wire [16-1:0] node3901;
	wire [16-1:0] node3902;
	wire [16-1:0] node3904;
	wire [16-1:0] node3907;
	wire [16-1:0] node3910;
	wire [16-1:0] node3911;
	wire [16-1:0] node3913;
	wire [16-1:0] node3916;
	wire [16-1:0] node3919;
	wire [16-1:0] node3920;
	wire [16-1:0] node3921;
	wire [16-1:0] node3924;
	wire [16-1:0] node3926;
	wire [16-1:0] node3929;
	wire [16-1:0] node3930;
	wire [16-1:0] node3931;
	wire [16-1:0] node3933;
	wire [16-1:0] node3936;
	wire [16-1:0] node3937;
	wire [16-1:0] node3941;
	wire [16-1:0] node3943;
	wire [16-1:0] node3944;
	wire [16-1:0] node3948;
	wire [16-1:0] node3949;
	wire [16-1:0] node3950;
	wire [16-1:0] node3951;
	wire [16-1:0] node3952;
	wire [16-1:0] node3953;
	wire [16-1:0] node3955;
	wire [16-1:0] node3960;
	wire [16-1:0] node3961;
	wire [16-1:0] node3965;
	wire [16-1:0] node3966;
	wire [16-1:0] node3968;
	wire [16-1:0] node3970;
	wire [16-1:0] node3973;
	wire [16-1:0] node3975;
	wire [16-1:0] node3978;
	wire [16-1:0] node3979;
	wire [16-1:0] node3980;
	wire [16-1:0] node3981;
	wire [16-1:0] node3983;
	wire [16-1:0] node3986;
	wire [16-1:0] node3989;
	wire [16-1:0] node3990;
	wire [16-1:0] node3992;
	wire [16-1:0] node3995;
	wire [16-1:0] node3996;
	wire [16-1:0] node3997;
	wire [16-1:0] node4001;
	wire [16-1:0] node4003;
	wire [16-1:0] node4006;
	wire [16-1:0] node4007;
	wire [16-1:0] node4008;
	wire [16-1:0] node4011;
	wire [16-1:0] node4012;
	wire [16-1:0] node4013;
	wire [16-1:0] node4017;
	wire [16-1:0] node4020;
	wire [16-1:0] node4021;
	wire [16-1:0] node4023;
	wire [16-1:0] node4024;
	wire [16-1:0] node4026;
	wire [16-1:0] node4029;
	wire [16-1:0] node4032;
	wire [16-1:0] node4035;
	wire [16-1:0] node4036;
	wire [16-1:0] node4037;
	wire [16-1:0] node4038;
	wire [16-1:0] node4039;
	wire [16-1:0] node4040;
	wire [16-1:0] node4041;
	wire [16-1:0] node4043;
	wire [16-1:0] node4046;
	wire [16-1:0] node4047;
	wire [16-1:0] node4051;
	wire [16-1:0] node4052;
	wire [16-1:0] node4054;
	wire [16-1:0] node4057;
	wire [16-1:0] node4060;
	wire [16-1:0] node4061;
	wire [16-1:0] node4062;
	wire [16-1:0] node4064;
	wire [16-1:0] node4067;
	wire [16-1:0] node4070;
	wire [16-1:0] node4071;
	wire [16-1:0] node4072;
	wire [16-1:0] node4076;
	wire [16-1:0] node4079;
	wire [16-1:0] node4080;
	wire [16-1:0] node4081;
	wire [16-1:0] node4083;
	wire [16-1:0] node4085;
	wire [16-1:0] node4088;
	wire [16-1:0] node4089;
	wire [16-1:0] node4092;
	wire [16-1:0] node4093;
	wire [16-1:0] node4097;
	wire [16-1:0] node4098;
	wire [16-1:0] node4100;
	wire [16-1:0] node4102;
	wire [16-1:0] node4105;
	wire [16-1:0] node4107;
	wire [16-1:0] node4108;
	wire [16-1:0] node4109;
	wire [16-1:0] node4113;
	wire [16-1:0] node4116;
	wire [16-1:0] node4117;
	wire [16-1:0] node4118;
	wire [16-1:0] node4119;
	wire [16-1:0] node4120;
	wire [16-1:0] node4122;
	wire [16-1:0] node4126;
	wire [16-1:0] node4129;
	wire [16-1:0] node4130;
	wire [16-1:0] node4132;
	wire [16-1:0] node4133;
	wire [16-1:0] node4136;
	wire [16-1:0] node4139;
	wire [16-1:0] node4140;
	wire [16-1:0] node4141;
	wire [16-1:0] node4145;
	wire [16-1:0] node4146;
	wire [16-1:0] node4150;
	wire [16-1:0] node4151;
	wire [16-1:0] node4152;
	wire [16-1:0] node4154;
	wire [16-1:0] node4156;
	wire [16-1:0] node4159;
	wire [16-1:0] node4160;
	wire [16-1:0] node4162;
	wire [16-1:0] node4166;
	wire [16-1:0] node4167;
	wire [16-1:0] node4169;
	wire [16-1:0] node4171;
	wire [16-1:0] node4172;
	wire [16-1:0] node4176;
	wire [16-1:0] node4178;
	wire [16-1:0] node4180;
	wire [16-1:0] node4183;
	wire [16-1:0] node4184;
	wire [16-1:0] node4185;
	wire [16-1:0] node4186;
	wire [16-1:0] node4187;
	wire [16-1:0] node4188;
	wire [16-1:0] node4190;
	wire [16-1:0] node4194;
	wire [16-1:0] node4195;
	wire [16-1:0] node4197;
	wire [16-1:0] node4201;
	wire [16-1:0] node4202;
	wire [16-1:0] node4203;
	wire [16-1:0] node4205;
	wire [16-1:0] node4207;
	wire [16-1:0] node4210;
	wire [16-1:0] node4213;
	wire [16-1:0] node4214;
	wire [16-1:0] node4215;
	wire [16-1:0] node4219;
	wire [16-1:0] node4221;
	wire [16-1:0] node4224;
	wire [16-1:0] node4225;
	wire [16-1:0] node4226;
	wire [16-1:0] node4227;
	wire [16-1:0] node4228;
	wire [16-1:0] node4232;
	wire [16-1:0] node4233;
	wire [16-1:0] node4237;
	wire [16-1:0] node4238;
	wire [16-1:0] node4239;
	wire [16-1:0] node4240;
	wire [16-1:0] node4245;
	wire [16-1:0] node4246;
	wire [16-1:0] node4250;
	wire [16-1:0] node4251;
	wire [16-1:0] node4252;
	wire [16-1:0] node4253;
	wire [16-1:0] node4258;
	wire [16-1:0] node4259;
	wire [16-1:0] node4262;
	wire [16-1:0] node4263;
	wire [16-1:0] node4267;
	wire [16-1:0] node4268;
	wire [16-1:0] node4269;
	wire [16-1:0] node4270;
	wire [16-1:0] node4271;
	wire [16-1:0] node4274;
	wire [16-1:0] node4275;
	wire [16-1:0] node4278;
	wire [16-1:0] node4281;
	wire [16-1:0] node4283;
	wire [16-1:0] node4284;
	wire [16-1:0] node4288;
	wire [16-1:0] node4289;
	wire [16-1:0] node4290;
	wire [16-1:0] node4291;
	wire [16-1:0] node4295;
	wire [16-1:0] node4296;
	wire [16-1:0] node4299;
	wire [16-1:0] node4302;
	wire [16-1:0] node4304;
	wire [16-1:0] node4307;
	wire [16-1:0] node4308;
	wire [16-1:0] node4309;
	wire [16-1:0] node4310;
	wire [16-1:0] node4312;
	wire [16-1:0] node4316;
	wire [16-1:0] node4317;
	wire [16-1:0] node4320;
	wire [16-1:0] node4321;
	wire [16-1:0] node4322;
	wire [16-1:0] node4324;
	wire [16-1:0] node4328;
	wire [16-1:0] node4331;
	wire [16-1:0] node4332;
	wire [16-1:0] node4333;
	wire [16-1:0] node4334;
	wire [16-1:0] node4338;
	wire [16-1:0] node4341;
	wire [16-1:0] node4343;
	wire [16-1:0] node4344;
	wire [16-1:0] node4347;
	wire [16-1:0] node4348;
	wire [16-1:0] node4352;
	wire [16-1:0] node4353;
	wire [16-1:0] node4354;
	wire [16-1:0] node4355;
	wire [16-1:0] node4356;
	wire [16-1:0] node4357;
	wire [16-1:0] node4358;
	wire [16-1:0] node4359;
	wire [16-1:0] node4360;
	wire [16-1:0] node4361;
	wire [16-1:0] node4365;
	wire [16-1:0] node4366;
	wire [16-1:0] node4367;
	wire [16-1:0] node4372;
	wire [16-1:0] node4374;
	wire [16-1:0] node4375;
	wire [16-1:0] node4379;
	wire [16-1:0] node4380;
	wire [16-1:0] node4381;
	wire [16-1:0] node4384;
	wire [16-1:0] node4385;
	wire [16-1:0] node4389;
	wire [16-1:0] node4390;
	wire [16-1:0] node4391;
	wire [16-1:0] node4394;
	wire [16-1:0] node4397;
	wire [16-1:0] node4398;
	wire [16-1:0] node4401;
	wire [16-1:0] node4403;
	wire [16-1:0] node4406;
	wire [16-1:0] node4407;
	wire [16-1:0] node4408;
	wire [16-1:0] node4409;
	wire [16-1:0] node4410;
	wire [16-1:0] node4413;
	wire [16-1:0] node4416;
	wire [16-1:0] node4418;
	wire [16-1:0] node4420;
	wire [16-1:0] node4423;
	wire [16-1:0] node4424;
	wire [16-1:0] node4426;
	wire [16-1:0] node4429;
	wire [16-1:0] node4430;
	wire [16-1:0] node4433;
	wire [16-1:0] node4434;
	wire [16-1:0] node4437;
	wire [16-1:0] node4438;
	wire [16-1:0] node4442;
	wire [16-1:0] node4443;
	wire [16-1:0] node4444;
	wire [16-1:0] node4445;
	wire [16-1:0] node4450;
	wire [16-1:0] node4453;
	wire [16-1:0] node4454;
	wire [16-1:0] node4455;
	wire [16-1:0] node4456;
	wire [16-1:0] node4457;
	wire [16-1:0] node4460;
	wire [16-1:0] node4461;
	wire [16-1:0] node4462;
	wire [16-1:0] node4466;
	wire [16-1:0] node4469;
	wire [16-1:0] node4470;
	wire [16-1:0] node4471;
	wire [16-1:0] node4474;
	wire [16-1:0] node4477;
	wire [16-1:0] node4478;
	wire [16-1:0] node4482;
	wire [16-1:0] node4483;
	wire [16-1:0] node4485;
	wire [16-1:0] node4486;
	wire [16-1:0] node4490;
	wire [16-1:0] node4492;
	wire [16-1:0] node4493;
	wire [16-1:0] node4495;
	wire [16-1:0] node4496;
	wire [16-1:0] node4501;
	wire [16-1:0] node4502;
	wire [16-1:0] node4503;
	wire [16-1:0] node4504;
	wire [16-1:0] node4507;
	wire [16-1:0] node4508;
	wire [16-1:0] node4512;
	wire [16-1:0] node4513;
	wire [16-1:0] node4515;
	wire [16-1:0] node4517;
	wire [16-1:0] node4518;
	wire [16-1:0] node4522;
	wire [16-1:0] node4523;
	wire [16-1:0] node4524;
	wire [16-1:0] node4529;
	wire [16-1:0] node4530;
	wire [16-1:0] node4532;
	wire [16-1:0] node4533;
	wire [16-1:0] node4535;
	wire [16-1:0] node4536;
	wire [16-1:0] node4541;
	wire [16-1:0] node4542;
	wire [16-1:0] node4544;
	wire [16-1:0] node4546;
	wire [16-1:0] node4548;
	wire [16-1:0] node4552;
	wire [16-1:0] node4553;
	wire [16-1:0] node4554;
	wire [16-1:0] node4555;
	wire [16-1:0] node4556;
	wire [16-1:0] node4557;
	wire [16-1:0] node4558;
	wire [16-1:0] node4559;
	wire [16-1:0] node4561;
	wire [16-1:0] node4566;
	wire [16-1:0] node4567;
	wire [16-1:0] node4571;
	wire [16-1:0] node4572;
	wire [16-1:0] node4573;
	wire [16-1:0] node4574;
	wire [16-1:0] node4579;
	wire [16-1:0] node4581;
	wire [16-1:0] node4584;
	wire [16-1:0] node4585;
	wire [16-1:0] node4587;
	wire [16-1:0] node4588;
	wire [16-1:0] node4592;
	wire [16-1:0] node4594;
	wire [16-1:0] node4596;
	wire [16-1:0] node4599;
	wire [16-1:0] node4600;
	wire [16-1:0] node4601;
	wire [16-1:0] node4603;
	wire [16-1:0] node4604;
	wire [16-1:0] node4605;
	wire [16-1:0] node4606;
	wire [16-1:0] node4612;
	wire [16-1:0] node4613;
	wire [16-1:0] node4614;
	wire [16-1:0] node4617;
	wire [16-1:0] node4618;
	wire [16-1:0] node4622;
	wire [16-1:0] node4625;
	wire [16-1:0] node4626;
	wire [16-1:0] node4628;
	wire [16-1:0] node4630;
	wire [16-1:0] node4633;
	wire [16-1:0] node4634;
	wire [16-1:0] node4637;
	wire [16-1:0] node4639;
	wire [16-1:0] node4641;
	wire [16-1:0] node4644;
	wire [16-1:0] node4645;
	wire [16-1:0] node4646;
	wire [16-1:0] node4647;
	wire [16-1:0] node4649;
	wire [16-1:0] node4650;
	wire [16-1:0] node4651;
	wire [16-1:0] node4653;
	wire [16-1:0] node4656;
	wire [16-1:0] node4657;
	wire [16-1:0] node4660;
	wire [16-1:0] node4664;
	wire [16-1:0] node4665;
	wire [16-1:0] node4667;
	wire [16-1:0] node4670;
	wire [16-1:0] node4672;
	wire [16-1:0] node4673;
	wire [16-1:0] node4677;
	wire [16-1:0] node4678;
	wire [16-1:0] node4680;
	wire [16-1:0] node4681;
	wire [16-1:0] node4685;
	wire [16-1:0] node4687;
	wire [16-1:0] node4688;
	wire [16-1:0] node4692;
	wire [16-1:0] node4693;
	wire [16-1:0] node4694;
	wire [16-1:0] node4695;
	wire [16-1:0] node4699;
	wire [16-1:0] node4700;
	wire [16-1:0] node4701;
	wire [16-1:0] node4703;
	wire [16-1:0] node4706;
	wire [16-1:0] node4709;
	wire [16-1:0] node4711;
	wire [16-1:0] node4714;
	wire [16-1:0] node4715;
	wire [16-1:0] node4717;
	wire [16-1:0] node4718;
	wire [16-1:0] node4721;
	wire [16-1:0] node4724;
	wire [16-1:0] node4725;
	wire [16-1:0] node4728;
	wire [16-1:0] node4729;
	wire [16-1:0] node4733;
	wire [16-1:0] node4734;
	wire [16-1:0] node4735;
	wire [16-1:0] node4736;
	wire [16-1:0] node4737;
	wire [16-1:0] node4738;
	wire [16-1:0] node4741;
	wire [16-1:0] node4743;
	wire [16-1:0] node4744;
	wire [16-1:0] node4748;
	wire [16-1:0] node4749;
	wire [16-1:0] node4750;
	wire [16-1:0] node4751;
	wire [16-1:0] node4754;
	wire [16-1:0] node4757;
	wire [16-1:0] node4758;
	wire [16-1:0] node4760;
	wire [16-1:0] node4763;
	wire [16-1:0] node4766;
	wire [16-1:0] node4767;
	wire [16-1:0] node4768;
	wire [16-1:0] node4770;
	wire [16-1:0] node4771;
	wire [16-1:0] node4775;
	wire [16-1:0] node4778;
	wire [16-1:0] node4779;
	wire [16-1:0] node4780;
	wire [16-1:0] node4782;
	wire [16-1:0] node4786;
	wire [16-1:0] node4789;
	wire [16-1:0] node4790;
	wire [16-1:0] node4791;
	wire [16-1:0] node4792;
	wire [16-1:0] node4793;
	wire [16-1:0] node4795;
	wire [16-1:0] node4800;
	wire [16-1:0] node4801;
	wire [16-1:0] node4802;
	wire [16-1:0] node4804;
	wire [16-1:0] node4805;
	wire [16-1:0] node4809;
	wire [16-1:0] node4811;
	wire [16-1:0] node4814;
	wire [16-1:0] node4815;
	wire [16-1:0] node4816;
	wire [16-1:0] node4820;
	wire [16-1:0] node4823;
	wire [16-1:0] node4824;
	wire [16-1:0] node4825;
	wire [16-1:0] node4827;
	wire [16-1:0] node4828;
	wire [16-1:0] node4832;
	wire [16-1:0] node4833;
	wire [16-1:0] node4837;
	wire [16-1:0] node4838;
	wire [16-1:0] node4839;
	wire [16-1:0] node4844;
	wire [16-1:0] node4845;
	wire [16-1:0] node4846;
	wire [16-1:0] node4847;
	wire [16-1:0] node4848;
	wire [16-1:0] node4851;
	wire [16-1:0] node4852;
	wire [16-1:0] node4856;
	wire [16-1:0] node4857;
	wire [16-1:0] node4858;
	wire [16-1:0] node4860;
	wire [16-1:0] node4861;
	wire [16-1:0] node4865;
	wire [16-1:0] node4868;
	wire [16-1:0] node4869;
	wire [16-1:0] node4873;
	wire [16-1:0] node4874;
	wire [16-1:0] node4875;
	wire [16-1:0] node4876;
	wire [16-1:0] node4880;
	wire [16-1:0] node4881;
	wire [16-1:0] node4885;
	wire [16-1:0] node4886;
	wire [16-1:0] node4887;
	wire [16-1:0] node4890;
	wire [16-1:0] node4892;
	wire [16-1:0] node4895;
	wire [16-1:0] node4897;
	wire [16-1:0] node4900;
	wire [16-1:0] node4901;
	wire [16-1:0] node4902;
	wire [16-1:0] node4903;
	wire [16-1:0] node4905;
	wire [16-1:0] node4908;
	wire [16-1:0] node4910;
	wire [16-1:0] node4913;
	wire [16-1:0] node4914;
	wire [16-1:0] node4917;
	wire [16-1:0] node4918;
	wire [16-1:0] node4922;
	wire [16-1:0] node4923;
	wire [16-1:0] node4924;
	wire [16-1:0] node4927;
	wire [16-1:0] node4928;
	wire [16-1:0] node4931;
	wire [16-1:0] node4933;
	wire [16-1:0] node4936;
	wire [16-1:0] node4937;
	wire [16-1:0] node4939;
	wire [16-1:0] node4940;
	wire [16-1:0] node4944;
	wire [16-1:0] node4946;
	wire [16-1:0] node4949;
	wire [16-1:0] node4950;
	wire [16-1:0] node4951;
	wire [16-1:0] node4952;
	wire [16-1:0] node4953;
	wire [16-1:0] node4954;
	wire [16-1:0] node4955;
	wire [16-1:0] node4958;
	wire [16-1:0] node4959;
	wire [16-1:0] node4961;
	wire [16-1:0] node4966;
	wire [16-1:0] node4967;
	wire [16-1:0] node4968;
	wire [16-1:0] node4969;
	wire [16-1:0] node4973;
	wire [16-1:0] node4975;
	wire [16-1:0] node4978;
	wire [16-1:0] node4979;
	wire [16-1:0] node4983;
	wire [16-1:0] node4984;
	wire [16-1:0] node4985;
	wire [16-1:0] node4986;
	wire [16-1:0] node4991;
	wire [16-1:0] node4992;
	wire [16-1:0] node4995;
	wire [16-1:0] node4996;
	wire [16-1:0] node5000;
	wire [16-1:0] node5001;
	wire [16-1:0] node5002;
	wire [16-1:0] node5003;
	wire [16-1:0] node5004;
	wire [16-1:0] node5008;
	wire [16-1:0] node5009;
	wire [16-1:0] node5013;
	wire [16-1:0] node5016;
	wire [16-1:0] node5017;
	wire [16-1:0] node5018;
	wire [16-1:0] node5021;
	wire [16-1:0] node5023;
	wire [16-1:0] node5026;
	wire [16-1:0] node5027;
	wire [16-1:0] node5029;
	wire [16-1:0] node5032;
	wire [16-1:0] node5033;
	wire [16-1:0] node5035;
	wire [16-1:0] node5038;
	wire [16-1:0] node5041;
	wire [16-1:0] node5042;
	wire [16-1:0] node5043;
	wire [16-1:0] node5044;
	wire [16-1:0] node5046;
	wire [16-1:0] node5049;
	wire [16-1:0] node5051;
	wire [16-1:0] node5052;
	wire [16-1:0] node5055;
	wire [16-1:0] node5058;
	wire [16-1:0] node5059;
	wire [16-1:0] node5060;
	wire [16-1:0] node5062;
	wire [16-1:0] node5065;
	wire [16-1:0] node5066;
	wire [16-1:0] node5067;
	wire [16-1:0] node5071;
	wire [16-1:0] node5072;
	wire [16-1:0] node5074;
	wire [16-1:0] node5078;
	wire [16-1:0] node5079;
	wire [16-1:0] node5081;
	wire [16-1:0] node5083;
	wire [16-1:0] node5084;
	wire [16-1:0] node5088;
	wire [16-1:0] node5089;
	wire [16-1:0] node5093;
	wire [16-1:0] node5094;
	wire [16-1:0] node5095;
	wire [16-1:0] node5096;
	wire [16-1:0] node5097;
	wire [16-1:0] node5100;
	wire [16-1:0] node5103;
	wire [16-1:0] node5104;
	wire [16-1:0] node5105;
	wire [16-1:0] node5109;
	wire [16-1:0] node5111;
	wire [16-1:0] node5114;
	wire [16-1:0] node5115;
	wire [16-1:0] node5117;
	wire [16-1:0] node5120;
	wire [16-1:0] node5121;
	wire [16-1:0] node5125;
	wire [16-1:0] node5126;
	wire [16-1:0] node5127;
	wire [16-1:0] node5128;
	wire [16-1:0] node5129;
	wire [16-1:0] node5130;
	wire [16-1:0] node5135;
	wire [16-1:0] node5137;
	wire [16-1:0] node5140;
	wire [16-1:0] node5141;
	wire [16-1:0] node5144;
	wire [16-1:0] node5146;
	wire [16-1:0] node5149;
	wire [16-1:0] node5150;
	wire [16-1:0] node5152;
	wire [16-1:0] node5156;
	wire [16-1:0] node5157;
	wire [16-1:0] node5158;
	wire [16-1:0] node5159;
	wire [16-1:0] node5160;
	wire [16-1:0] node5161;
	wire [16-1:0] node5162;
	wire [16-1:0] node5164;
	wire [16-1:0] node5167;
	wire [16-1:0] node5168;
	wire [16-1:0] node5171;
	wire [16-1:0] node5172;
	wire [16-1:0] node5173;
	wire [16-1:0] node5178;
	wire [16-1:0] node5179;
	wire [16-1:0] node5181;
	wire [16-1:0] node5184;
	wire [16-1:0] node5185;
	wire [16-1:0] node5186;
	wire [16-1:0] node5190;
	wire [16-1:0] node5191;
	wire [16-1:0] node5194;
	wire [16-1:0] node5197;
	wire [16-1:0] node5198;
	wire [16-1:0] node5199;
	wire [16-1:0] node5200;
	wire [16-1:0] node5202;
	wire [16-1:0] node5203;
	wire [16-1:0] node5205;
	wire [16-1:0] node5209;
	wire [16-1:0] node5210;
	wire [16-1:0] node5211;
	wire [16-1:0] node5216;
	wire [16-1:0] node5218;
	wire [16-1:0] node5219;
	wire [16-1:0] node5221;
	wire [16-1:0] node5222;
	wire [16-1:0] node5227;
	wire [16-1:0] node5228;
	wire [16-1:0] node5230;
	wire [16-1:0] node5231;
	wire [16-1:0] node5235;
	wire [16-1:0] node5236;
	wire [16-1:0] node5237;
	wire [16-1:0] node5239;
	wire [16-1:0] node5244;
	wire [16-1:0] node5245;
	wire [16-1:0] node5246;
	wire [16-1:0] node5247;
	wire [16-1:0] node5248;
	wire [16-1:0] node5251;
	wire [16-1:0] node5254;
	wire [16-1:0] node5256;
	wire [16-1:0] node5257;
	wire [16-1:0] node5259;
	wire [16-1:0] node5263;
	wire [16-1:0] node5264;
	wire [16-1:0] node5266;
	wire [16-1:0] node5267;
	wire [16-1:0] node5269;
	wire [16-1:0] node5272;
	wire [16-1:0] node5275;
	wire [16-1:0] node5277;
	wire [16-1:0] node5280;
	wire [16-1:0] node5281;
	wire [16-1:0] node5282;
	wire [16-1:0] node5283;
	wire [16-1:0] node5284;
	wire [16-1:0] node5288;
	wire [16-1:0] node5289;
	wire [16-1:0] node5290;
	wire [16-1:0] node5295;
	wire [16-1:0] node5296;
	wire [16-1:0] node5297;
	wire [16-1:0] node5301;
	wire [16-1:0] node5303;
	wire [16-1:0] node5306;
	wire [16-1:0] node5307;
	wire [16-1:0] node5310;
	wire [16-1:0] node5311;
	wire [16-1:0] node5313;
	wire [16-1:0] node5317;
	wire [16-1:0] node5318;
	wire [16-1:0] node5319;
	wire [16-1:0] node5320;
	wire [16-1:0] node5321;
	wire [16-1:0] node5322;
	wire [16-1:0] node5323;
	wire [16-1:0] node5324;
	wire [16-1:0] node5326;
	wire [16-1:0] node5331;
	wire [16-1:0] node5332;
	wire [16-1:0] node5334;
	wire [16-1:0] node5337;
	wire [16-1:0] node5340;
	wire [16-1:0] node5341;
	wire [16-1:0] node5343;
	wire [16-1:0] node5344;
	wire [16-1:0] node5348;
	wire [16-1:0] node5350;
	wire [16-1:0] node5353;
	wire [16-1:0] node5354;
	wire [16-1:0] node5355;
	wire [16-1:0] node5358;
	wire [16-1:0] node5359;
	wire [16-1:0] node5363;
	wire [16-1:0] node5364;
	wire [16-1:0] node5366;
	wire [16-1:0] node5369;
	wire [16-1:0] node5370;
	wire [16-1:0] node5373;
	wire [16-1:0] node5376;
	wire [16-1:0] node5377;
	wire [16-1:0] node5378;
	wire [16-1:0] node5379;
	wire [16-1:0] node5380;
	wire [16-1:0] node5385;
	wire [16-1:0] node5386;
	wire [16-1:0] node5387;
	wire [16-1:0] node5391;
	wire [16-1:0] node5392;
	wire [16-1:0] node5393;
	wire [16-1:0] node5398;
	wire [16-1:0] node5399;
	wire [16-1:0] node5400;
	wire [16-1:0] node5404;
	wire [16-1:0] node5405;
	wire [16-1:0] node5406;
	wire [16-1:0] node5407;
	wire [16-1:0] node5411;
	wire [16-1:0] node5412;
	wire [16-1:0] node5416;
	wire [16-1:0] node5418;
	wire [16-1:0] node5420;
	wire [16-1:0] node5422;
	wire [16-1:0] node5425;
	wire [16-1:0] node5426;
	wire [16-1:0] node5427;
	wire [16-1:0] node5428;
	wire [16-1:0] node5431;
	wire [16-1:0] node5432;
	wire [16-1:0] node5433;
	wire [16-1:0] node5434;
	wire [16-1:0] node5436;
	wire [16-1:0] node5440;
	wire [16-1:0] node5443;
	wire [16-1:0] node5444;
	wire [16-1:0] node5445;
	wire [16-1:0] node5449;
	wire [16-1:0] node5450;
	wire [16-1:0] node5452;
	wire [16-1:0] node5456;
	wire [16-1:0] node5457;
	wire [16-1:0] node5458;
	wire [16-1:0] node5462;
	wire [16-1:0] node5463;
	wire [16-1:0] node5466;
	wire [16-1:0] node5469;
	wire [16-1:0] node5470;
	wire [16-1:0] node5471;
	wire [16-1:0] node5472;
	wire [16-1:0] node5474;
	wire [16-1:0] node5476;
	wire [16-1:0] node5480;
	wire [16-1:0] node5481;
	wire [16-1:0] node5482;
	wire [16-1:0] node5484;
	wire [16-1:0] node5488;
	wire [16-1:0] node5491;
	wire [16-1:0] node5492;
	wire [16-1:0] node5493;
	wire [16-1:0] node5495;
	wire [16-1:0] node5496;
	wire [16-1:0] node5500;
	wire [16-1:0] node5501;
	wire [16-1:0] node5503;
	wire [16-1:0] node5508;
	wire [16-1:0] node5509;
	wire [16-1:0] node5510;
	wire [16-1:0] node5511;
	wire [16-1:0] node5512;
	wire [16-1:0] node5513;
	wire [16-1:0] node5514;
	wire [16-1:0] node5516;
	wire [16-1:0] node5518;
	wire [16-1:0] node5521;
	wire [16-1:0] node5522;
	wire [16-1:0] node5526;
	wire [16-1:0] node5527;
	wire [16-1:0] node5529;
	wire [16-1:0] node5530;
	wire [16-1:0] node5532;
	wire [16-1:0] node5537;
	wire [16-1:0] node5538;
	wire [16-1:0] node5539;
	wire [16-1:0] node5540;
	wire [16-1:0] node5541;
	wire [16-1:0] node5545;
	wire [16-1:0] node5547;
	wire [16-1:0] node5550;
	wire [16-1:0] node5552;
	wire [16-1:0] node5555;
	wire [16-1:0] node5556;
	wire [16-1:0] node5559;
	wire [16-1:0] node5561;
	wire [16-1:0] node5563;
	wire [16-1:0] node5566;
	wire [16-1:0] node5567;
	wire [16-1:0] node5568;
	wire [16-1:0] node5569;
	wire [16-1:0] node5573;
	wire [16-1:0] node5574;
	wire [16-1:0] node5578;
	wire [16-1:0] node5579;
	wire [16-1:0] node5580;
	wire [16-1:0] node5581;
	wire [16-1:0] node5584;
	wire [16-1:0] node5587;
	wire [16-1:0] node5590;
	wire [16-1:0] node5592;
	wire [16-1:0] node5593;
	wire [16-1:0] node5595;
	wire [16-1:0] node5599;
	wire [16-1:0] node5600;
	wire [16-1:0] node5601;
	wire [16-1:0] node5602;
	wire [16-1:0] node5603;
	wire [16-1:0] node5604;
	wire [16-1:0] node5607;
	wire [16-1:0] node5610;
	wire [16-1:0] node5611;
	wire [16-1:0] node5613;
	wire [16-1:0] node5614;
	wire [16-1:0] node5619;
	wire [16-1:0] node5621;
	wire [16-1:0] node5622;
	wire [16-1:0] node5626;
	wire [16-1:0] node5627;
	wire [16-1:0] node5628;
	wire [16-1:0] node5629;
	wire [16-1:0] node5632;
	wire [16-1:0] node5635;
	wire [16-1:0] node5636;
	wire [16-1:0] node5639;
	wire [16-1:0] node5642;
	wire [16-1:0] node5643;
	wire [16-1:0] node5645;
	wire [16-1:0] node5649;
	wire [16-1:0] node5650;
	wire [16-1:0] node5651;
	wire [16-1:0] node5652;
	wire [16-1:0] node5654;
	wire [16-1:0] node5655;
	wire [16-1:0] node5657;
	wire [16-1:0] node5660;
	wire [16-1:0] node5664;
	wire [16-1:0] node5666;
	wire [16-1:0] node5667;
	wire [16-1:0] node5669;
	wire [16-1:0] node5671;
	wire [16-1:0] node5675;
	wire [16-1:0] node5676;
	wire [16-1:0] node5679;
	wire [16-1:0] node5680;
	wire [16-1:0] node5682;
	wire [16-1:0] node5685;
	wire [16-1:0] node5687;
	wire [16-1:0] node5690;
	wire [16-1:0] node5691;
	wire [16-1:0] node5692;
	wire [16-1:0] node5693;
	wire [16-1:0] node5694;
	wire [16-1:0] node5697;
	wire [16-1:0] node5698;
	wire [16-1:0] node5700;
	wire [16-1:0] node5702;
	wire [16-1:0] node5703;
	wire [16-1:0] node5707;
	wire [16-1:0] node5708;
	wire [16-1:0] node5709;
	wire [16-1:0] node5714;
	wire [16-1:0] node5715;
	wire [16-1:0] node5716;
	wire [16-1:0] node5718;
	wire [16-1:0] node5721;
	wire [16-1:0] node5722;
	wire [16-1:0] node5723;
	wire [16-1:0] node5727;
	wire [16-1:0] node5730;
	wire [16-1:0] node5733;
	wire [16-1:0] node5734;
	wire [16-1:0] node5735;
	wire [16-1:0] node5736;
	wire [16-1:0] node5739;
	wire [16-1:0] node5740;
	wire [16-1:0] node5743;
	wire [16-1:0] node5746;
	wire [16-1:0] node5749;
	wire [16-1:0] node5750;
	wire [16-1:0] node5751;
	wire [16-1:0] node5752;
	wire [16-1:0] node5754;
	wire [16-1:0] node5758;
	wire [16-1:0] node5759;
	wire [16-1:0] node5760;
	wire [16-1:0] node5764;
	wire [16-1:0] node5767;
	wire [16-1:0] node5768;
	wire [16-1:0] node5770;
	wire [16-1:0] node5773;
	wire [16-1:0] node5776;
	wire [16-1:0] node5777;
	wire [16-1:0] node5778;
	wire [16-1:0] node5779;
	wire [16-1:0] node5780;
	wire [16-1:0] node5781;
	wire [16-1:0] node5785;
	wire [16-1:0] node5788;
	wire [16-1:0] node5790;
	wire [16-1:0] node5793;
	wire [16-1:0] node5794;
	wire [16-1:0] node5795;
	wire [16-1:0] node5796;
	wire [16-1:0] node5797;
	wire [16-1:0] node5799;
	wire [16-1:0] node5802;
	wire [16-1:0] node5807;
	wire [16-1:0] node5809;
	wire [16-1:0] node5810;
	wire [16-1:0] node5812;
	wire [16-1:0] node5815;
	wire [16-1:0] node5818;
	wire [16-1:0] node5819;
	wire [16-1:0] node5820;
	wire [16-1:0] node5821;
	wire [16-1:0] node5824;
	wire [16-1:0] node5825;
	wire [16-1:0] node5827;
	wire [16-1:0] node5828;
	wire [16-1:0] node5832;
	wire [16-1:0] node5835;
	wire [16-1:0] node5836;
	wire [16-1:0] node5837;
	wire [16-1:0] node5841;
	wire [16-1:0] node5842;
	wire [16-1:0] node5846;
	wire [16-1:0] node5847;
	wire [16-1:0] node5848;
	wire [16-1:0] node5850;
	wire [16-1:0] node5853;
	wire [16-1:0] node5854;
	wire [16-1:0] node5858;
	wire [16-1:0] node5859;
	wire [16-1:0] node5861;
	wire [16-1:0] node5864;
	wire [16-1:0] node5865;
	wire [16-1:0] node5866;
	wire [16-1:0] node5868;
	wire [16-1:0] node5872;
	wire [16-1:0] node5873;
	wire [16-1:0] node5877;
	wire [16-1:0] node5878;
	wire [16-1:0] node5879;
	wire [16-1:0] node5880;
	wire [16-1:0] node5881;
	wire [16-1:0] node5882;
	wire [16-1:0] node5883;
	wire [16-1:0] node5884;
	wire [16-1:0] node5885;
	wire [16-1:0] node5886;
	wire [16-1:0] node5887;
	wire [16-1:0] node5890;
	wire [16-1:0] node5892;
	wire [16-1:0] node5894;
	wire [16-1:0] node5897;
	wire [16-1:0] node5898;
	wire [16-1:0] node5899;
	wire [16-1:0] node5902;
	wire [16-1:0] node5904;
	wire [16-1:0] node5907;
	wire [16-1:0] node5908;
	wire [16-1:0] node5910;
	wire [16-1:0] node5914;
	wire [16-1:0] node5915;
	wire [16-1:0] node5916;
	wire [16-1:0] node5917;
	wire [16-1:0] node5921;
	wire [16-1:0] node5923;
	wire [16-1:0] node5924;
	wire [16-1:0] node5928;
	wire [16-1:0] node5929;
	wire [16-1:0] node5930;
	wire [16-1:0] node5934;
	wire [16-1:0] node5935;
	wire [16-1:0] node5939;
	wire [16-1:0] node5940;
	wire [16-1:0] node5941;
	wire [16-1:0] node5942;
	wire [16-1:0] node5943;
	wire [16-1:0] node5944;
	wire [16-1:0] node5950;
	wire [16-1:0] node5951;
	wire [16-1:0] node5954;
	wire [16-1:0] node5955;
	wire [16-1:0] node5957;
	wire [16-1:0] node5958;
	wire [16-1:0] node5963;
	wire [16-1:0] node5964;
	wire [16-1:0] node5965;
	wire [16-1:0] node5967;
	wire [16-1:0] node5968;
	wire [16-1:0] node5972;
	wire [16-1:0] node5974;
	wire [16-1:0] node5977;
	wire [16-1:0] node5978;
	wire [16-1:0] node5979;
	wire [16-1:0] node5982;
	wire [16-1:0] node5985;
	wire [16-1:0] node5986;
	wire [16-1:0] node5989;
	wire [16-1:0] node5991;
	wire [16-1:0] node5994;
	wire [16-1:0] node5995;
	wire [16-1:0] node5996;
	wire [16-1:0] node5997;
	wire [16-1:0] node5998;
	wire [16-1:0] node5999;
	wire [16-1:0] node6002;
	wire [16-1:0] node6005;
	wire [16-1:0] node6007;
	wire [16-1:0] node6010;
	wire [16-1:0] node6012;
	wire [16-1:0] node6015;
	wire [16-1:0] node6016;
	wire [16-1:0] node6017;
	wire [16-1:0] node6019;
	wire [16-1:0] node6022;
	wire [16-1:0] node6023;
	wire [16-1:0] node6027;
	wire [16-1:0] node6028;
	wire [16-1:0] node6029;
	wire [16-1:0] node6032;
	wire [16-1:0] node6035;
	wire [16-1:0] node6036;
	wire [16-1:0] node6039;
	wire [16-1:0] node6042;
	wire [16-1:0] node6043;
	wire [16-1:0] node6044;
	wire [16-1:0] node6045;
	wire [16-1:0] node6046;
	wire [16-1:0] node6047;
	wire [16-1:0] node6053;
	wire [16-1:0] node6054;
	wire [16-1:0] node6055;
	wire [16-1:0] node6058;
	wire [16-1:0] node6061;
	wire [16-1:0] node6064;
	wire [16-1:0] node6065;
	wire [16-1:0] node6066;
	wire [16-1:0] node6069;
	wire [16-1:0] node6072;
	wire [16-1:0] node6075;
	wire [16-1:0] node6076;
	wire [16-1:0] node6077;
	wire [16-1:0] node6078;
	wire [16-1:0] node6079;
	wire [16-1:0] node6080;
	wire [16-1:0] node6083;
	wire [16-1:0] node6084;
	wire [16-1:0] node6086;
	wire [16-1:0] node6087;
	wire [16-1:0] node6092;
	wire [16-1:0] node6093;
	wire [16-1:0] node6095;
	wire [16-1:0] node6098;
	wire [16-1:0] node6100;
	wire [16-1:0] node6101;
	wire [16-1:0] node6105;
	wire [16-1:0] node6106;
	wire [16-1:0] node6108;
	wire [16-1:0] node6109;
	wire [16-1:0] node6113;
	wire [16-1:0] node6114;
	wire [16-1:0] node6115;
	wire [16-1:0] node6118;
	wire [16-1:0] node6121;
	wire [16-1:0] node6124;
	wire [16-1:0] node6125;
	wire [16-1:0] node6126;
	wire [16-1:0] node6127;
	wire [16-1:0] node6128;
	wire [16-1:0] node6132;
	wire [16-1:0] node6135;
	wire [16-1:0] node6136;
	wire [16-1:0] node6138;
	wire [16-1:0] node6140;
	wire [16-1:0] node6143;
	wire [16-1:0] node6144;
	wire [16-1:0] node6148;
	wire [16-1:0] node6149;
	wire [16-1:0] node6150;
	wire [16-1:0] node6151;
	wire [16-1:0] node6154;
	wire [16-1:0] node6157;
	wire [16-1:0] node6159;
	wire [16-1:0] node6162;
	wire [16-1:0] node6163;
	wire [16-1:0] node6166;
	wire [16-1:0] node6169;
	wire [16-1:0] node6170;
	wire [16-1:0] node6171;
	wire [16-1:0] node6172;
	wire [16-1:0] node6173;
	wire [16-1:0] node6174;
	wire [16-1:0] node6177;
	wire [16-1:0] node6180;
	wire [16-1:0] node6181;
	wire [16-1:0] node6182;
	wire [16-1:0] node6186;
	wire [16-1:0] node6189;
	wire [16-1:0] node6192;
	wire [16-1:0] node6193;
	wire [16-1:0] node6194;
	wire [16-1:0] node6195;
	wire [16-1:0] node6198;
	wire [16-1:0] node6201;
	wire [16-1:0] node6202;
	wire [16-1:0] node6205;
	wire [16-1:0] node6208;
	wire [16-1:0] node6209;
	wire [16-1:0] node6210;
	wire [16-1:0] node6214;
	wire [16-1:0] node6217;
	wire [16-1:0] node6218;
	wire [16-1:0] node6219;
	wire [16-1:0] node6222;
	wire [16-1:0] node6224;
	wire [16-1:0] node6225;
	wire [16-1:0] node6229;
	wire [16-1:0] node6230;
	wire [16-1:0] node6231;
	wire [16-1:0] node6233;
	wire [16-1:0] node6236;
	wire [16-1:0] node6237;
	wire [16-1:0] node6241;
	wire [16-1:0] node6242;
	wire [16-1:0] node6243;
	wire [16-1:0] node6246;
	wire [16-1:0] node6249;
	wire [16-1:0] node6250;
	wire [16-1:0] node6254;
	wire [16-1:0] node6255;
	wire [16-1:0] node6256;
	wire [16-1:0] node6257;
	wire [16-1:0] node6258;
	wire [16-1:0] node6259;
	wire [16-1:0] node6260;
	wire [16-1:0] node6263;
	wire [16-1:0] node6264;
	wire [16-1:0] node6267;
	wire [16-1:0] node6270;
	wire [16-1:0] node6271;
	wire [16-1:0] node6272;
	wire [16-1:0] node6273;
	wire [16-1:0] node6278;
	wire [16-1:0] node6279;
	wire [16-1:0] node6283;
	wire [16-1:0] node6284;
	wire [16-1:0] node6285;
	wire [16-1:0] node6288;
	wire [16-1:0] node6291;
	wire [16-1:0] node6292;
	wire [16-1:0] node6293;
	wire [16-1:0] node6296;
	wire [16-1:0] node6297;
	wire [16-1:0] node6301;
	wire [16-1:0] node6304;
	wire [16-1:0] node6305;
	wire [16-1:0] node6306;
	wire [16-1:0] node6307;
	wire [16-1:0] node6308;
	wire [16-1:0] node6310;
	wire [16-1:0] node6313;
	wire [16-1:0] node6315;
	wire [16-1:0] node6318;
	wire [16-1:0] node6319;
	wire [16-1:0] node6322;
	wire [16-1:0] node6325;
	wire [16-1:0] node6326;
	wire [16-1:0] node6327;
	wire [16-1:0] node6328;
	wire [16-1:0] node6332;
	wire [16-1:0] node6333;
	wire [16-1:0] node6334;
	wire [16-1:0] node6337;
	wire [16-1:0] node6341;
	wire [16-1:0] node6344;
	wire [16-1:0] node6345;
	wire [16-1:0] node6346;
	wire [16-1:0] node6348;
	wire [16-1:0] node6350;
	wire [16-1:0] node6353;
	wire [16-1:0] node6354;
	wire [16-1:0] node6357;
	wire [16-1:0] node6359;
	wire [16-1:0] node6362;
	wire [16-1:0] node6363;
	wire [16-1:0] node6364;
	wire [16-1:0] node6368;
	wire [16-1:0] node6369;
	wire [16-1:0] node6373;
	wire [16-1:0] node6374;
	wire [16-1:0] node6375;
	wire [16-1:0] node6376;
	wire [16-1:0] node6377;
	wire [16-1:0] node6380;
	wire [16-1:0] node6383;
	wire [16-1:0] node6384;
	wire [16-1:0] node6385;
	wire [16-1:0] node6388;
	wire [16-1:0] node6391;
	wire [16-1:0] node6393;
	wire [16-1:0] node6396;
	wire [16-1:0] node6397;
	wire [16-1:0] node6398;
	wire [16-1:0] node6402;
	wire [16-1:0] node6405;
	wire [16-1:0] node6406;
	wire [16-1:0] node6408;
	wire [16-1:0] node6410;
	wire [16-1:0] node6411;
	wire [16-1:0] node6415;
	wire [16-1:0] node6416;
	wire [16-1:0] node6417;
	wire [16-1:0] node6418;
	wire [16-1:0] node6421;
	wire [16-1:0] node6423;
	wire [16-1:0] node6426;
	wire [16-1:0] node6427;
	wire [16-1:0] node6428;
	wire [16-1:0] node6433;
	wire [16-1:0] node6434;
	wire [16-1:0] node6435;
	wire [16-1:0] node6437;
	wire [16-1:0] node6440;
	wire [16-1:0] node6442;
	wire [16-1:0] node6445;
	wire [16-1:0] node6446;
	wire [16-1:0] node6450;
	wire [16-1:0] node6451;
	wire [16-1:0] node6452;
	wire [16-1:0] node6453;
	wire [16-1:0] node6454;
	wire [16-1:0] node6456;
	wire [16-1:0] node6458;
	wire [16-1:0] node6459;
	wire [16-1:0] node6463;
	wire [16-1:0] node6464;
	wire [16-1:0] node6466;
	wire [16-1:0] node6467;
	wire [16-1:0] node6468;
	wire [16-1:0] node6473;
	wire [16-1:0] node6475;
	wire [16-1:0] node6476;
	wire [16-1:0] node6477;
	wire [16-1:0] node6482;
	wire [16-1:0] node6484;
	wire [16-1:0] node6485;
	wire [16-1:0] node6489;
	wire [16-1:0] node6490;
	wire [16-1:0] node6491;
	wire [16-1:0] node6493;
	wire [16-1:0] node6494;
	wire [16-1:0] node6499;
	wire [16-1:0] node6500;
	wire [16-1:0] node6501;
	wire [16-1:0] node6504;
	wire [16-1:0] node6505;
	wire [16-1:0] node6509;
	wire [16-1:0] node6510;
	wire [16-1:0] node6513;
	wire [16-1:0] node6516;
	wire [16-1:0] node6517;
	wire [16-1:0] node6518;
	wire [16-1:0] node6519;
	wire [16-1:0] node6521;
	wire [16-1:0] node6523;
	wire [16-1:0] node6526;
	wire [16-1:0] node6527;
	wire [16-1:0] node6529;
	wire [16-1:0] node6530;
	wire [16-1:0] node6531;
	wire [16-1:0] node6536;
	wire [16-1:0] node6537;
	wire [16-1:0] node6541;
	wire [16-1:0] node6542;
	wire [16-1:0] node6543;
	wire [16-1:0] node6544;
	wire [16-1:0] node6548;
	wire [16-1:0] node6551;
	wire [16-1:0] node6552;
	wire [16-1:0] node6554;
	wire [16-1:0] node6557;
	wire [16-1:0] node6559;
	wire [16-1:0] node6561;
	wire [16-1:0] node6564;
	wire [16-1:0] node6565;
	wire [16-1:0] node6566;
	wire [16-1:0] node6567;
	wire [16-1:0] node6570;
	wire [16-1:0] node6572;
	wire [16-1:0] node6574;
	wire [16-1:0] node6577;
	wire [16-1:0] node6578;
	wire [16-1:0] node6580;
	wire [16-1:0] node6582;
	wire [16-1:0] node6585;
	wire [16-1:0] node6588;
	wire [16-1:0] node6589;
	wire [16-1:0] node6590;
	wire [16-1:0] node6593;
	wire [16-1:0] node6595;
	wire [16-1:0] node6598;
	wire [16-1:0] node6600;
	wire [16-1:0] node6601;
	wire [16-1:0] node6604;
	wire [16-1:0] node6607;
	wire [16-1:0] node6608;
	wire [16-1:0] node6609;
	wire [16-1:0] node6610;
	wire [16-1:0] node6611;
	wire [16-1:0] node6612;
	wire [16-1:0] node6613;
	wire [16-1:0] node6614;
	wire [16-1:0] node6615;
	wire [16-1:0] node6616;
	wire [16-1:0] node6617;
	wire [16-1:0] node6621;
	wire [16-1:0] node6623;
	wire [16-1:0] node6627;
	wire [16-1:0] node6630;
	wire [16-1:0] node6631;
	wire [16-1:0] node6632;
	wire [16-1:0] node6635;
	wire [16-1:0] node6637;
	wire [16-1:0] node6640;
	wire [16-1:0] node6641;
	wire [16-1:0] node6642;
	wire [16-1:0] node6646;
	wire [16-1:0] node6649;
	wire [16-1:0] node6650;
	wire [16-1:0] node6651;
	wire [16-1:0] node6653;
	wire [16-1:0] node6654;
	wire [16-1:0] node6656;
	wire [16-1:0] node6659;
	wire [16-1:0] node6663;
	wire [16-1:0] node6664;
	wire [16-1:0] node6665;
	wire [16-1:0] node6668;
	wire [16-1:0] node6669;
	wire [16-1:0] node6671;
	wire [16-1:0] node6675;
	wire [16-1:0] node6678;
	wire [16-1:0] node6679;
	wire [16-1:0] node6680;
	wire [16-1:0] node6681;
	wire [16-1:0] node6682;
	wire [16-1:0] node6683;
	wire [16-1:0] node6687;
	wire [16-1:0] node6690;
	wire [16-1:0] node6691;
	wire [16-1:0] node6695;
	wire [16-1:0] node6696;
	wire [16-1:0] node6697;
	wire [16-1:0] node6701;
	wire [16-1:0] node6702;
	wire [16-1:0] node6704;
	wire [16-1:0] node6707;
	wire [16-1:0] node6710;
	wire [16-1:0] node6711;
	wire [16-1:0] node6712;
	wire [16-1:0] node6713;
	wire [16-1:0] node6717;
	wire [16-1:0] node6718;
	wire [16-1:0] node6720;
	wire [16-1:0] node6721;
	wire [16-1:0] node6725;
	wire [16-1:0] node6728;
	wire [16-1:0] node6729;
	wire [16-1:0] node6730;
	wire [16-1:0] node6731;
	wire [16-1:0] node6736;
	wire [16-1:0] node6737;
	wire [16-1:0] node6740;
	wire [16-1:0] node6743;
	wire [16-1:0] node6744;
	wire [16-1:0] node6745;
	wire [16-1:0] node6746;
	wire [16-1:0] node6748;
	wire [16-1:0] node6749;
	wire [16-1:0] node6753;
	wire [16-1:0] node6755;
	wire [16-1:0] node6756;
	wire [16-1:0] node6760;
	wire [16-1:0] node6761;
	wire [16-1:0] node6762;
	wire [16-1:0] node6765;
	wire [16-1:0] node6767;
	wire [16-1:0] node6769;
	wire [16-1:0] node6772;
	wire [16-1:0] node6774;
	wire [16-1:0] node6777;
	wire [16-1:0] node6778;
	wire [16-1:0] node6779;
	wire [16-1:0] node6780;
	wire [16-1:0] node6781;
	wire [16-1:0] node6785;
	wire [16-1:0] node6788;
	wire [16-1:0] node6790;
	wire [16-1:0] node6792;
	wire [16-1:0] node6794;
	wire [16-1:0] node6795;
	wire [16-1:0] node6799;
	wire [16-1:0] node6800;
	wire [16-1:0] node6801;
	wire [16-1:0] node6803;
	wire [16-1:0] node6806;
	wire [16-1:0] node6809;
	wire [16-1:0] node6812;
	wire [16-1:0] node6813;
	wire [16-1:0] node6814;
	wire [16-1:0] node6815;
	wire [16-1:0] node6816;
	wire [16-1:0] node6817;
	wire [16-1:0] node6818;
	wire [16-1:0] node6822;
	wire [16-1:0] node6823;
	wire [16-1:0] node6827;
	wire [16-1:0] node6828;
	wire [16-1:0] node6829;
	wire [16-1:0] node6834;
	wire [16-1:0] node6835;
	wire [16-1:0] node6836;
	wire [16-1:0] node6837;
	wire [16-1:0] node6838;
	wire [16-1:0] node6842;
	wire [16-1:0] node6845;
	wire [16-1:0] node6846;
	wire [16-1:0] node6849;
	wire [16-1:0] node6850;
	wire [16-1:0] node6854;
	wire [16-1:0] node6855;
	wire [16-1:0] node6856;
	wire [16-1:0] node6857;
	wire [16-1:0] node6861;
	wire [16-1:0] node6864;
	wire [16-1:0] node6865;
	wire [16-1:0] node6869;
	wire [16-1:0] node6870;
	wire [16-1:0] node6871;
	wire [16-1:0] node6872;
	wire [16-1:0] node6875;
	wire [16-1:0] node6876;
	wire [16-1:0] node6880;
	wire [16-1:0] node6881;
	wire [16-1:0] node6882;
	wire [16-1:0] node6885;
	wire [16-1:0] node6888;
	wire [16-1:0] node6890;
	wire [16-1:0] node6892;
	wire [16-1:0] node6895;
	wire [16-1:0] node6896;
	wire [16-1:0] node6898;
	wire [16-1:0] node6899;
	wire [16-1:0] node6902;
	wire [16-1:0] node6903;
	wire [16-1:0] node6905;
	wire [16-1:0] node6909;
	wire [16-1:0] node6910;
	wire [16-1:0] node6913;
	wire [16-1:0] node6916;
	wire [16-1:0] node6917;
	wire [16-1:0] node6918;
	wire [16-1:0] node6919;
	wire [16-1:0] node6920;
	wire [16-1:0] node6922;
	wire [16-1:0] node6925;
	wire [16-1:0] node6926;
	wire [16-1:0] node6930;
	wire [16-1:0] node6931;
	wire [16-1:0] node6932;
	wire [16-1:0] node6936;
	wire [16-1:0] node6938;
	wire [16-1:0] node6941;
	wire [16-1:0] node6942;
	wire [16-1:0] node6943;
	wire [16-1:0] node6946;
	wire [16-1:0] node6947;
	wire [16-1:0] node6950;
	wire [16-1:0] node6953;
	wire [16-1:0] node6954;
	wire [16-1:0] node6955;
	wire [16-1:0] node6956;
	wire [16-1:0] node6961;
	wire [16-1:0] node6962;
	wire [16-1:0] node6965;
	wire [16-1:0] node6966;
	wire [16-1:0] node6968;
	wire [16-1:0] node6972;
	wire [16-1:0] node6973;
	wire [16-1:0] node6974;
	wire [16-1:0] node6976;
	wire [16-1:0] node6977;
	wire [16-1:0] node6978;
	wire [16-1:0] node6982;
	wire [16-1:0] node6985;
	wire [16-1:0] node6986;
	wire [16-1:0] node6988;
	wire [16-1:0] node6991;
	wire [16-1:0] node6992;
	wire [16-1:0] node6995;
	wire [16-1:0] node6997;
	wire [16-1:0] node7000;
	wire [16-1:0] node7001;
	wire [16-1:0] node7002;
	wire [16-1:0] node7004;
	wire [16-1:0] node7006;
	wire [16-1:0] node7009;
	wire [16-1:0] node7011;
	wire [16-1:0] node7012;
	wire [16-1:0] node7014;
	wire [16-1:0] node7018;
	wire [16-1:0] node7019;
	wire [16-1:0] node7021;
	wire [16-1:0] node7024;
	wire [16-1:0] node7025;
	wire [16-1:0] node7028;
	wire [16-1:0] node7031;
	wire [16-1:0] node7032;
	wire [16-1:0] node7033;
	wire [16-1:0] node7034;
	wire [16-1:0] node7035;
	wire [16-1:0] node7036;
	wire [16-1:0] node7037;
	wire [16-1:0] node7038;
	wire [16-1:0] node7041;
	wire [16-1:0] node7044;
	wire [16-1:0] node7045;
	wire [16-1:0] node7046;
	wire [16-1:0] node7050;
	wire [16-1:0] node7053;
	wire [16-1:0] node7056;
	wire [16-1:0] node7057;
	wire [16-1:0] node7058;
	wire [16-1:0] node7059;
	wire [16-1:0] node7060;
	wire [16-1:0] node7064;
	wire [16-1:0] node7067;
	wire [16-1:0] node7069;
	wire [16-1:0] node7073;
	wire [16-1:0] node7074;
	wire [16-1:0] node7075;
	wire [16-1:0] node7076;
	wire [16-1:0] node7078;
	wire [16-1:0] node7081;
	wire [16-1:0] node7082;
	wire [16-1:0] node7083;
	wire [16-1:0] node7088;
	wire [16-1:0] node7090;
	wire [16-1:0] node7091;
	wire [16-1:0] node7092;
	wire [16-1:0] node7097;
	wire [16-1:0] node7098;
	wire [16-1:0] node7100;
	wire [16-1:0] node7101;
	wire [16-1:0] node7105;
	wire [16-1:0] node7107;
	wire [16-1:0] node7108;
	wire [16-1:0] node7109;
	wire [16-1:0] node7111;
	wire [16-1:0] node7116;
	wire [16-1:0] node7117;
	wire [16-1:0] node7118;
	wire [16-1:0] node7119;
	wire [16-1:0] node7121;
	wire [16-1:0] node7122;
	wire [16-1:0] node7126;
	wire [16-1:0] node7127;
	wire [16-1:0] node7128;
	wire [16-1:0] node7132;
	wire [16-1:0] node7133;
	wire [16-1:0] node7137;
	wire [16-1:0] node7138;
	wire [16-1:0] node7139;
	wire [16-1:0] node7140;
	wire [16-1:0] node7144;
	wire [16-1:0] node7145;
	wire [16-1:0] node7146;
	wire [16-1:0] node7148;
	wire [16-1:0] node7152;
	wire [16-1:0] node7155;
	wire [16-1:0] node7156;
	wire [16-1:0] node7158;
	wire [16-1:0] node7160;
	wire [16-1:0] node7163;
	wire [16-1:0] node7164;
	wire [16-1:0] node7168;
	wire [16-1:0] node7169;
	wire [16-1:0] node7170;
	wire [16-1:0] node7171;
	wire [16-1:0] node7175;
	wire [16-1:0] node7176;
	wire [16-1:0] node7177;
	wire [16-1:0] node7181;
	wire [16-1:0] node7182;
	wire [16-1:0] node7186;
	wire [16-1:0] node7187;
	wire [16-1:0] node7189;
	wire [16-1:0] node7190;
	wire [16-1:0] node7191;
	wire [16-1:0] node7196;
	wire [16-1:0] node7197;
	wire [16-1:0] node7199;
	wire [16-1:0] node7202;
	wire [16-1:0] node7203;
	wire [16-1:0] node7204;
	wire [16-1:0] node7208;
	wire [16-1:0] node7211;
	wire [16-1:0] node7212;
	wire [16-1:0] node7213;
	wire [16-1:0] node7214;
	wire [16-1:0] node7215;
	wire [16-1:0] node7216;
	wire [16-1:0] node7217;
	wire [16-1:0] node7220;
	wire [16-1:0] node7221;
	wire [16-1:0] node7223;
	wire [16-1:0] node7226;
	wire [16-1:0] node7230;
	wire [16-1:0] node7232;
	wire [16-1:0] node7235;
	wire [16-1:0] node7236;
	wire [16-1:0] node7237;
	wire [16-1:0] node7238;
	wire [16-1:0] node7242;
	wire [16-1:0] node7243;
	wire [16-1:0] node7244;
	wire [16-1:0] node7249;
	wire [16-1:0] node7250;
	wire [16-1:0] node7251;
	wire [16-1:0] node7252;
	wire [16-1:0] node7254;
	wire [16-1:0] node7258;
	wire [16-1:0] node7261;
	wire [16-1:0] node7264;
	wire [16-1:0] node7265;
	wire [16-1:0] node7266;
	wire [16-1:0] node7267;
	wire [16-1:0] node7268;
	wire [16-1:0] node7269;
	wire [16-1:0] node7273;
	wire [16-1:0] node7276;
	wire [16-1:0] node7277;
	wire [16-1:0] node7280;
	wire [16-1:0] node7282;
	wire [16-1:0] node7285;
	wire [16-1:0] node7286;
	wire [16-1:0] node7288;
	wire [16-1:0] node7291;
	wire [16-1:0] node7294;
	wire [16-1:0] node7295;
	wire [16-1:0] node7296;
	wire [16-1:0] node7299;
	wire [16-1:0] node7301;
	wire [16-1:0] node7304;
	wire [16-1:0] node7305;
	wire [16-1:0] node7306;
	wire [16-1:0] node7310;
	wire [16-1:0] node7311;
	wire [16-1:0] node7312;
	wire [16-1:0] node7317;
	wire [16-1:0] node7318;
	wire [16-1:0] node7319;
	wire [16-1:0] node7320;
	wire [16-1:0] node7321;
	wire [16-1:0] node7322;
	wire [16-1:0] node7323;
	wire [16-1:0] node7327;
	wire [16-1:0] node7330;
	wire [16-1:0] node7332;
	wire [16-1:0] node7335;
	wire [16-1:0] node7337;
	wire [16-1:0] node7338;
	wire [16-1:0] node7342;
	wire [16-1:0] node7343;
	wire [16-1:0] node7344;
	wire [16-1:0] node7345;
	wire [16-1:0] node7349;
	wire [16-1:0] node7351;
	wire [16-1:0] node7354;
	wire [16-1:0] node7355;
	wire [16-1:0] node7356;
	wire [16-1:0] node7360;
	wire [16-1:0] node7362;
	wire [16-1:0] node7364;
	wire [16-1:0] node7366;
	wire [16-1:0] node7369;
	wire [16-1:0] node7370;
	wire [16-1:0] node7371;
	wire [16-1:0] node7372;
	wire [16-1:0] node7374;
	wire [16-1:0] node7377;
	wire [16-1:0] node7379;
	wire [16-1:0] node7382;
	wire [16-1:0] node7383;
	wire [16-1:0] node7384;
	wire [16-1:0] node7387;
	wire [16-1:0] node7390;
	wire [16-1:0] node7393;
	wire [16-1:0] node7394;
	wire [16-1:0] node7395;
	wire [16-1:0] node7399;
	wire [16-1:0] node7400;
	wire [16-1:0] node7403;
	wire [16-1:0] node7404;
	wire [16-1:0] node7407;
	wire [16-1:0] node7409;
	wire [16-1:0] node7412;
	wire [16-1:0] node7413;
	wire [16-1:0] node7414;
	wire [16-1:0] node7415;
	wire [16-1:0] node7416;
	wire [16-1:0] node7417;
	wire [16-1:0] node7418;
	wire [16-1:0] node7419;
	wire [16-1:0] node7420;
	wire [16-1:0] node7422;
	wire [16-1:0] node7424;
	wire [16-1:0] node7427;
	wire [16-1:0] node7428;
	wire [16-1:0] node7432;
	wire [16-1:0] node7433;
	wire [16-1:0] node7434;
	wire [16-1:0] node7435;
	wire [16-1:0] node7441;
	wire [16-1:0] node7442;
	wire [16-1:0] node7445;
	wire [16-1:0] node7447;
	wire [16-1:0] node7448;
	wire [16-1:0] node7452;
	wire [16-1:0] node7453;
	wire [16-1:0] node7454;
	wire [16-1:0] node7455;
	wire [16-1:0] node7456;
	wire [16-1:0] node7461;
	wire [16-1:0] node7463;
	wire [16-1:0] node7464;
	wire [16-1:0] node7468;
	wire [16-1:0] node7469;
	wire [16-1:0] node7470;
	wire [16-1:0] node7471;
	wire [16-1:0] node7475;
	wire [16-1:0] node7477;
	wire [16-1:0] node7479;
	wire [16-1:0] node7482;
	wire [16-1:0] node7483;
	wire [16-1:0] node7485;
	wire [16-1:0] node7488;
	wire [16-1:0] node7490;
	wire [16-1:0] node7493;
	wire [16-1:0] node7494;
	wire [16-1:0] node7495;
	wire [16-1:0] node7496;
	wire [16-1:0] node7497;
	wire [16-1:0] node7499;
	wire [16-1:0] node7502;
	wire [16-1:0] node7504;
	wire [16-1:0] node7506;
	wire [16-1:0] node7507;
	wire [16-1:0] node7511;
	wire [16-1:0] node7512;
	wire [16-1:0] node7514;
	wire [16-1:0] node7518;
	wire [16-1:0] node7519;
	wire [16-1:0] node7520;
	wire [16-1:0] node7523;
	wire [16-1:0] node7526;
	wire [16-1:0] node7527;
	wire [16-1:0] node7528;
	wire [16-1:0] node7531;
	wire [16-1:0] node7535;
	wire [16-1:0] node7536;
	wire [16-1:0] node7537;
	wire [16-1:0] node7538;
	wire [16-1:0] node7540;
	wire [16-1:0] node7542;
	wire [16-1:0] node7544;
	wire [16-1:0] node7548;
	wire [16-1:0] node7549;
	wire [16-1:0] node7550;
	wire [16-1:0] node7551;
	wire [16-1:0] node7553;
	wire [16-1:0] node7558;
	wire [16-1:0] node7561;
	wire [16-1:0] node7562;
	wire [16-1:0] node7565;
	wire [16-1:0] node7566;
	wire [16-1:0] node7569;
	wire [16-1:0] node7570;
	wire [16-1:0] node7573;
	wire [16-1:0] node7576;
	wire [16-1:0] node7577;
	wire [16-1:0] node7578;
	wire [16-1:0] node7579;
	wire [16-1:0] node7580;
	wire [16-1:0] node7581;
	wire [16-1:0] node7582;
	wire [16-1:0] node7586;
	wire [16-1:0] node7589;
	wire [16-1:0] node7590;
	wire [16-1:0] node7591;
	wire [16-1:0] node7593;
	wire [16-1:0] node7596;
	wire [16-1:0] node7599;
	wire [16-1:0] node7602;
	wire [16-1:0] node7603;
	wire [16-1:0] node7604;
	wire [16-1:0] node7606;
	wire [16-1:0] node7609;
	wire [16-1:0] node7610;
	wire [16-1:0] node7614;
	wire [16-1:0] node7615;
	wire [16-1:0] node7617;
	wire [16-1:0] node7619;
	wire [16-1:0] node7620;
	wire [16-1:0] node7624;
	wire [16-1:0] node7626;
	wire [16-1:0] node7629;
	wire [16-1:0] node7630;
	wire [16-1:0] node7631;
	wire [16-1:0] node7633;
	wire [16-1:0] node7636;
	wire [16-1:0] node7638;
	wire [16-1:0] node7640;
	wire [16-1:0] node7643;
	wire [16-1:0] node7644;
	wire [16-1:0] node7645;
	wire [16-1:0] node7646;
	wire [16-1:0] node7650;
	wire [16-1:0] node7651;
	wire [16-1:0] node7654;
	wire [16-1:0] node7656;
	wire [16-1:0] node7659;
	wire [16-1:0] node7660;
	wire [16-1:0] node7663;
	wire [16-1:0] node7666;
	wire [16-1:0] node7667;
	wire [16-1:0] node7668;
	wire [16-1:0] node7669;
	wire [16-1:0] node7670;
	wire [16-1:0] node7671;
	wire [16-1:0] node7675;
	wire [16-1:0] node7676;
	wire [16-1:0] node7677;
	wire [16-1:0] node7679;
	wire [16-1:0] node7684;
	wire [16-1:0] node7685;
	wire [16-1:0] node7686;
	wire [16-1:0] node7687;
	wire [16-1:0] node7693;
	wire [16-1:0] node7694;
	wire [16-1:0] node7696;
	wire [16-1:0] node7699;
	wire [16-1:0] node7701;
	wire [16-1:0] node7703;
	wire [16-1:0] node7704;
	wire [16-1:0] node7708;
	wire [16-1:0] node7709;
	wire [16-1:0] node7710;
	wire [16-1:0] node7712;
	wire [16-1:0] node7713;
	wire [16-1:0] node7716;
	wire [16-1:0] node7717;
	wire [16-1:0] node7721;
	wire [16-1:0] node7722;
	wire [16-1:0] node7723;
	wire [16-1:0] node7724;
	wire [16-1:0] node7729;
	wire [16-1:0] node7730;
	wire [16-1:0] node7732;
	wire [16-1:0] node7736;
	wire [16-1:0] node7737;
	wire [16-1:0] node7740;
	wire [16-1:0] node7741;
	wire [16-1:0] node7742;
	wire [16-1:0] node7743;
	wire [16-1:0] node7745;
	wire [16-1:0] node7750;
	wire [16-1:0] node7751;
	wire [16-1:0] node7753;
	wire [16-1:0] node7756;
	wire [16-1:0] node7759;
	wire [16-1:0] node7760;
	wire [16-1:0] node7761;
	wire [16-1:0] node7762;
	wire [16-1:0] node7763;
	wire [16-1:0] node7764;
	wire [16-1:0] node7765;
	wire [16-1:0] node7768;
	wire [16-1:0] node7769;
	wire [16-1:0] node7770;
	wire [16-1:0] node7772;
	wire [16-1:0] node7777;
	wire [16-1:0] node7780;
	wire [16-1:0] node7781;
	wire [16-1:0] node7782;
	wire [16-1:0] node7783;
	wire [16-1:0] node7787;
	wire [16-1:0] node7788;
	wire [16-1:0] node7789;
	wire [16-1:0] node7794;
	wire [16-1:0] node7795;
	wire [16-1:0] node7796;
	wire [16-1:0] node7800;
	wire [16-1:0] node7801;
	wire [16-1:0] node7805;
	wire [16-1:0] node7806;
	wire [16-1:0] node7807;
	wire [16-1:0] node7808;
	wire [16-1:0] node7810;
	wire [16-1:0] node7811;
	wire [16-1:0] node7813;
	wire [16-1:0] node7816;
	wire [16-1:0] node7817;
	wire [16-1:0] node7821;
	wire [16-1:0] node7822;
	wire [16-1:0] node7826;
	wire [16-1:0] node7828;
	wire [16-1:0] node7829;
	wire [16-1:0] node7832;
	wire [16-1:0] node7834;
	wire [16-1:0] node7837;
	wire [16-1:0] node7838;
	wire [16-1:0] node7840;
	wire [16-1:0] node7841;
	wire [16-1:0] node7844;
	wire [16-1:0] node7846;
	wire [16-1:0] node7849;
	wire [16-1:0] node7850;
	wire [16-1:0] node7852;
	wire [16-1:0] node7855;
	wire [16-1:0] node7856;
	wire [16-1:0] node7857;
	wire [16-1:0] node7861;
	wire [16-1:0] node7864;
	wire [16-1:0] node7865;
	wire [16-1:0] node7866;
	wire [16-1:0] node7867;
	wire [16-1:0] node7868;
	wire [16-1:0] node7871;
	wire [16-1:0] node7874;
	wire [16-1:0] node7875;
	wire [16-1:0] node7876;
	wire [16-1:0] node7880;
	wire [16-1:0] node7882;
	wire [16-1:0] node7885;
	wire [16-1:0] node7886;
	wire [16-1:0] node7887;
	wire [16-1:0] node7888;
	wire [16-1:0] node7890;
	wire [16-1:0] node7895;
	wire [16-1:0] node7896;
	wire [16-1:0] node7897;
	wire [16-1:0] node7899;
	wire [16-1:0] node7902;
	wire [16-1:0] node7905;
	wire [16-1:0] node7908;
	wire [16-1:0] node7909;
	wire [16-1:0] node7910;
	wire [16-1:0] node7911;
	wire [16-1:0] node7915;
	wire [16-1:0] node7917;
	wire [16-1:0] node7919;
	wire [16-1:0] node7921;
	wire [16-1:0] node7924;
	wire [16-1:0] node7925;
	wire [16-1:0] node7926;
	wire [16-1:0] node7930;
	wire [16-1:0] node7931;
	wire [16-1:0] node7934;
	wire [16-1:0] node7936;
	wire [16-1:0] node7939;
	wire [16-1:0] node7940;
	wire [16-1:0] node7941;
	wire [16-1:0] node7942;
	wire [16-1:0] node7943;
	wire [16-1:0] node7944;
	wire [16-1:0] node7946;
	wire [16-1:0] node7947;
	wire [16-1:0] node7951;
	wire [16-1:0] node7952;
	wire [16-1:0] node7953;
	wire [16-1:0] node7958;
	wire [16-1:0] node7959;
	wire [16-1:0] node7960;
	wire [16-1:0] node7964;
	wire [16-1:0] node7965;
	wire [16-1:0] node7968;
	wire [16-1:0] node7971;
	wire [16-1:0] node7972;
	wire [16-1:0] node7973;
	wire [16-1:0] node7975;
	wire [16-1:0] node7978;
	wire [16-1:0] node7979;
	wire [16-1:0] node7980;
	wire [16-1:0] node7982;
	wire [16-1:0] node7987;
	wire [16-1:0] node7988;
	wire [16-1:0] node7990;
	wire [16-1:0] node7993;
	wire [16-1:0] node7995;
	wire [16-1:0] node7997;
	wire [16-1:0] node7998;
	wire [16-1:0] node8002;
	wire [16-1:0] node8003;
	wire [16-1:0] node8004;
	wire [16-1:0] node8005;
	wire [16-1:0] node8006;
	wire [16-1:0] node8009;
	wire [16-1:0] node8011;
	wire [16-1:0] node8014;
	wire [16-1:0] node8016;
	wire [16-1:0] node8019;
	wire [16-1:0] node8020;
	wire [16-1:0] node8021;
	wire [16-1:0] node8023;
	wire [16-1:0] node8025;
	wire [16-1:0] node8029;
	wire [16-1:0] node8031;
	wire [16-1:0] node8034;
	wire [16-1:0] node8035;
	wire [16-1:0] node8036;
	wire [16-1:0] node8038;
	wire [16-1:0] node8041;
	wire [16-1:0] node8042;
	wire [16-1:0] node8045;
	wire [16-1:0] node8048;
	wire [16-1:0] node8049;
	wire [16-1:0] node8050;
	wire [16-1:0] node8053;
	wire [16-1:0] node8056;
	wire [16-1:0] node8057;
	wire [16-1:0] node8059;
	wire [16-1:0] node8063;
	wire [16-1:0] node8064;
	wire [16-1:0] node8065;
	wire [16-1:0] node8066;
	wire [16-1:0] node8067;
	wire [16-1:0] node8071;
	wire [16-1:0] node8072;
	wire [16-1:0] node8076;
	wire [16-1:0] node8077;
	wire [16-1:0] node8078;
	wire [16-1:0] node8080;
	wire [16-1:0] node8083;
	wire [16-1:0] node8084;
	wire [16-1:0] node8087;
	wire [16-1:0] node8089;
	wire [16-1:0] node8092;
	wire [16-1:0] node8093;
	wire [16-1:0] node8095;
	wire [16-1:0] node8096;
	wire [16-1:0] node8098;
	wire [16-1:0] node8103;
	wire [16-1:0] node8104;
	wire [16-1:0] node8105;
	wire [16-1:0] node8106;
	wire [16-1:0] node8109;
	wire [16-1:0] node8110;
	wire [16-1:0] node8114;
	wire [16-1:0] node8115;
	wire [16-1:0] node8117;
	wire [16-1:0] node8120;
	wire [16-1:0] node8123;
	wire [16-1:0] node8124;
	wire [16-1:0] node8125;
	wire [16-1:0] node8127;
	wire [16-1:0] node8129;
	wire [16-1:0] node8133;
	wire [16-1:0] node8135;
	wire [16-1:0] node8137;
	wire [16-1:0] node8139;
	wire [16-1:0] node8142;
	wire [16-1:0] node8143;
	wire [16-1:0] node8144;
	wire [16-1:0] node8145;
	wire [16-1:0] node8146;
	wire [16-1:0] node8147;
	wire [16-1:0] node8148;
	wire [16-1:0] node8149;
	wire [16-1:0] node8150;
	wire [16-1:0] node8154;
	wire [16-1:0] node8157;
	wire [16-1:0] node8158;
	wire [16-1:0] node8159;
	wire [16-1:0] node8161;
	wire [16-1:0] node8165;
	wire [16-1:0] node8168;
	wire [16-1:0] node8169;
	wire [16-1:0] node8170;
	wire [16-1:0] node8171;
	wire [16-1:0] node8174;
	wire [16-1:0] node8178;
	wire [16-1:0] node8179;
	wire [16-1:0] node8181;
	wire [16-1:0] node8185;
	wire [16-1:0] node8186;
	wire [16-1:0] node8187;
	wire [16-1:0] node8188;
	wire [16-1:0] node8189;
	wire [16-1:0] node8193;
	wire [16-1:0] node8196;
	wire [16-1:0] node8197;
	wire [16-1:0] node8200;
	wire [16-1:0] node8201;
	wire [16-1:0] node8204;
	wire [16-1:0] node8207;
	wire [16-1:0] node8208;
	wire [16-1:0] node8209;
	wire [16-1:0] node8210;
	wire [16-1:0] node8211;
	wire [16-1:0] node8215;
	wire [16-1:0] node8217;
	wire [16-1:0] node8221;
	wire [16-1:0] node8222;
	wire [16-1:0] node8223;
	wire [16-1:0] node8225;
	wire [16-1:0] node8228;
	wire [16-1:0] node8230;
	wire [16-1:0] node8233;
	wire [16-1:0] node8235;
	wire [16-1:0] node8238;
	wire [16-1:0] node8239;
	wire [16-1:0] node8240;
	wire [16-1:0] node8241;
	wire [16-1:0] node8242;
	wire [16-1:0] node8243;
	wire [16-1:0] node8244;
	wire [16-1:0] node8247;
	wire [16-1:0] node8248;
	wire [16-1:0] node8252;
	wire [16-1:0] node8256;
	wire [16-1:0] node8257;
	wire [16-1:0] node8258;
	wire [16-1:0] node8259;
	wire [16-1:0] node8263;
	wire [16-1:0] node8265;
	wire [16-1:0] node8266;
	wire [16-1:0] node8270;
	wire [16-1:0] node8272;
	wire [16-1:0] node8275;
	wire [16-1:0] node8276;
	wire [16-1:0] node8277;
	wire [16-1:0] node8278;
	wire [16-1:0] node8280;
	wire [16-1:0] node8282;
	wire [16-1:0] node8285;
	wire [16-1:0] node8286;
	wire [16-1:0] node8290;
	wire [16-1:0] node8291;
	wire [16-1:0] node8294;
	wire [16-1:0] node8297;
	wire [16-1:0] node8298;
	wire [16-1:0] node8302;
	wire [16-1:0] node8303;
	wire [16-1:0] node8304;
	wire [16-1:0] node8306;
	wire [16-1:0] node8307;
	wire [16-1:0] node8309;
	wire [16-1:0] node8312;
	wire [16-1:0] node8315;
	wire [16-1:0] node8316;
	wire [16-1:0] node8318;
	wire [16-1:0] node8321;
	wire [16-1:0] node8322;
	wire [16-1:0] node8326;
	wire [16-1:0] node8327;
	wire [16-1:0] node8328;
	wire [16-1:0] node8329;
	wire [16-1:0] node8332;
	wire [16-1:0] node8333;
	wire [16-1:0] node8335;
	wire [16-1:0] node8339;
	wire [16-1:0] node8340;
	wire [16-1:0] node8341;
	wire [16-1:0] node8346;
	wire [16-1:0] node8347;
	wire [16-1:0] node8349;
	wire [16-1:0] node8352;
	wire [16-1:0] node8353;
	wire [16-1:0] node8357;
	wire [16-1:0] node8358;
	wire [16-1:0] node8359;
	wire [16-1:0] node8360;
	wire [16-1:0] node8361;
	wire [16-1:0] node8362;
	wire [16-1:0] node8364;
	wire [16-1:0] node8366;
	wire [16-1:0] node8370;
	wire [16-1:0] node8371;
	wire [16-1:0] node8372;
	wire [16-1:0] node8373;
	wire [16-1:0] node8377;
	wire [16-1:0] node8380;
	wire [16-1:0] node8383;
	wire [16-1:0] node8384;
	wire [16-1:0] node8385;
	wire [16-1:0] node8386;
	wire [16-1:0] node8389;
	wire [16-1:0] node8390;
	wire [16-1:0] node8395;
	wire [16-1:0] node8398;
	wire [16-1:0] node8399;
	wire [16-1:0] node8400;
	wire [16-1:0] node8401;
	wire [16-1:0] node8402;
	wire [16-1:0] node8404;
	wire [16-1:0] node8408;
	wire [16-1:0] node8409;
	wire [16-1:0] node8411;
	wire [16-1:0] node8414;
	wire [16-1:0] node8417;
	wire [16-1:0] node8419;
	wire [16-1:0] node8420;
	wire [16-1:0] node8423;
	wire [16-1:0] node8426;
	wire [16-1:0] node8427;
	wire [16-1:0] node8428;
	wire [16-1:0] node8429;
	wire [16-1:0] node8432;
	wire [16-1:0] node8435;
	wire [16-1:0] node8436;
	wire [16-1:0] node8437;
	wire [16-1:0] node8439;
	wire [16-1:0] node8443;
	wire [16-1:0] node8446;
	wire [16-1:0] node8447;
	wire [16-1:0] node8448;
	wire [16-1:0] node8450;
	wire [16-1:0] node8451;
	wire [16-1:0] node8456;
	wire [16-1:0] node8458;
	wire [16-1:0] node8461;
	wire [16-1:0] node8462;
	wire [16-1:0] node8463;
	wire [16-1:0] node8464;
	wire [16-1:0] node8466;
	wire [16-1:0] node8467;
	wire [16-1:0] node8470;
	wire [16-1:0] node8472;
	wire [16-1:0] node8475;
	wire [16-1:0] node8477;
	wire [16-1:0] node8478;
	wire [16-1:0] node8480;
	wire [16-1:0] node8484;
	wire [16-1:0] node8485;
	wire [16-1:0] node8487;
	wire [16-1:0] node8488;
	wire [16-1:0] node8490;
	wire [16-1:0] node8494;
	wire [16-1:0] node8495;
	wire [16-1:0] node8497;
	wire [16-1:0] node8501;
	wire [16-1:0] node8502;
	wire [16-1:0] node8503;
	wire [16-1:0] node8504;
	wire [16-1:0] node8505;
	wire [16-1:0] node8509;
	wire [16-1:0] node8510;
	wire [16-1:0] node8514;
	wire [16-1:0] node8515;
	wire [16-1:0] node8516;
	wire [16-1:0] node8517;
	wire [16-1:0] node8522;
	wire [16-1:0] node8525;
	wire [16-1:0] node8526;
	wire [16-1:0] node8527;
	wire [16-1:0] node8529;
	wire [16-1:0] node8531;
	wire [16-1:0] node8534;
	wire [16-1:0] node8535;
	wire [16-1:0] node8536;
	wire [16-1:0] node8538;
	wire [16-1:0] node8543;
	wire [16-1:0] node8544;
	wire [16-1:0] node8546;
	wire [16-1:0] node8548;
	wire [16-1:0] node8552;
	wire [16-1:0] node8553;
	wire [16-1:0] node8554;
	wire [16-1:0] node8555;
	wire [16-1:0] node8556;
	wire [16-1:0] node8557;
	wire [16-1:0] node8558;
	wire [16-1:0] node8559;
	wire [16-1:0] node8562;
	wire [16-1:0] node8565;
	wire [16-1:0] node8566;
	wire [16-1:0] node8567;
	wire [16-1:0] node8571;
	wire [16-1:0] node8574;
	wire [16-1:0] node8575;
	wire [16-1:0] node8577;
	wire [16-1:0] node8580;
	wire [16-1:0] node8581;
	wire [16-1:0] node8585;
	wire [16-1:0] node8586;
	wire [16-1:0] node8587;
	wire [16-1:0] node8588;
	wire [16-1:0] node8589;
	wire [16-1:0] node8591;
	wire [16-1:0] node8595;
	wire [16-1:0] node8598;
	wire [16-1:0] node8599;
	wire [16-1:0] node8603;
	wire [16-1:0] node8604;
	wire [16-1:0] node8606;
	wire [16-1:0] node8609;
	wire [16-1:0] node8611;
	wire [16-1:0] node8613;
	wire [16-1:0] node8615;
	wire [16-1:0] node8618;
	wire [16-1:0] node8619;
	wire [16-1:0] node8620;
	wire [16-1:0] node8621;
	wire [16-1:0] node8623;
	wire [16-1:0] node8625;
	wire [16-1:0] node8626;
	wire [16-1:0] node8630;
	wire [16-1:0] node8631;
	wire [16-1:0] node8635;
	wire [16-1:0] node8637;
	wire [16-1:0] node8639;
	wire [16-1:0] node8641;
	wire [16-1:0] node8644;
	wire [16-1:0] node8645;
	wire [16-1:0] node8647;
	wire [16-1:0] node8648;
	wire [16-1:0] node8652;
	wire [16-1:0] node8653;
	wire [16-1:0] node8654;
	wire [16-1:0] node8658;
	wire [16-1:0] node8659;
	wire [16-1:0] node8661;
	wire [16-1:0] node8664;
	wire [16-1:0] node8667;
	wire [16-1:0] node8668;
	wire [16-1:0] node8669;
	wire [16-1:0] node8670;
	wire [16-1:0] node8671;
	wire [16-1:0] node8674;
	wire [16-1:0] node8677;
	wire [16-1:0] node8678;
	wire [16-1:0] node8679;
	wire [16-1:0] node8681;
	wire [16-1:0] node8684;
	wire [16-1:0] node8686;
	wire [16-1:0] node8689;
	wire [16-1:0] node8692;
	wire [16-1:0] node8693;
	wire [16-1:0] node8694;
	wire [16-1:0] node8696;
	wire [16-1:0] node8697;
	wire [16-1:0] node8702;
	wire [16-1:0] node8703;
	wire [16-1:0] node8704;
	wire [16-1:0] node8709;
	wire [16-1:0] node8710;
	wire [16-1:0] node8711;
	wire [16-1:0] node8712;
	wire [16-1:0] node8713;
	wire [16-1:0] node8716;
	wire [16-1:0] node8718;
	wire [16-1:0] node8721;
	wire [16-1:0] node8722;
	wire [16-1:0] node8725;
	wire [16-1:0] node8728;
	wire [16-1:0] node8729;
	wire [16-1:0] node8732;
	wire [16-1:0] node8733;
	wire [16-1:0] node8737;
	wire [16-1:0] node8738;
	wire [16-1:0] node8739;
	wire [16-1:0] node8740;
	wire [16-1:0] node8742;
	wire [16-1:0] node8745;
	wire [16-1:0] node8748;
	wire [16-1:0] node8749;
	wire [16-1:0] node8752;
	wire [16-1:0] node8753;
	wire [16-1:0] node8755;
	wire [16-1:0] node8759;
	wire [16-1:0] node8760;
	wire [16-1:0] node8761;
	wire [16-1:0] node8764;
	wire [16-1:0] node8766;
	wire [16-1:0] node8768;
	wire [16-1:0] node8771;
	wire [16-1:0] node8773;
	wire [16-1:0] node8775;
	wire [16-1:0] node8778;
	wire [16-1:0] node8779;
	wire [16-1:0] node8780;
	wire [16-1:0] node8781;
	wire [16-1:0] node8782;
	wire [16-1:0] node8784;
	wire [16-1:0] node8785;
	wire [16-1:0] node8789;
	wire [16-1:0] node8790;
	wire [16-1:0] node8791;
	wire [16-1:0] node8795;
	wire [16-1:0] node8796;
	wire [16-1:0] node8800;
	wire [16-1:0] node8801;
	wire [16-1:0] node8803;
	wire [16-1:0] node8805;
	wire [16-1:0] node8807;
	wire [16-1:0] node8810;
	wire [16-1:0] node8811;
	wire [16-1:0] node8814;
	wire [16-1:0] node8815;
	wire [16-1:0] node8819;
	wire [16-1:0] node8820;
	wire [16-1:0] node8821;
	wire [16-1:0] node8822;
	wire [16-1:0] node8823;
	wire [16-1:0] node8827;
	wire [16-1:0] node8829;
	wire [16-1:0] node8832;
	wire [16-1:0] node8834;
	wire [16-1:0] node8835;
	wire [16-1:0] node8837;
	wire [16-1:0] node8841;
	wire [16-1:0] node8842;
	wire [16-1:0] node8843;
	wire [16-1:0] node8844;
	wire [16-1:0] node8849;
	wire [16-1:0] node8850;
	wire [16-1:0] node8852;
	wire [16-1:0] node8853;
	wire [16-1:0] node8856;
	wire [16-1:0] node8859;
	wire [16-1:0] node8861;
	wire [16-1:0] node8862;
	wire [16-1:0] node8863;
	wire [16-1:0] node8866;
	wire [16-1:0] node8869;
	wire [16-1:0] node8871;
	wire [16-1:0] node8874;
	wire [16-1:0] node8875;
	wire [16-1:0] node8876;
	wire [16-1:0] node8877;
	wire [16-1:0] node8880;
	wire [16-1:0] node8881;
	wire [16-1:0] node8883;
	wire [16-1:0] node8885;
	wire [16-1:0] node8887;
	wire [16-1:0] node8890;
	wire [16-1:0] node8891;
	wire [16-1:0] node8895;
	wire [16-1:0] node8896;
	wire [16-1:0] node8897;
	wire [16-1:0] node8901;
	wire [16-1:0] node8903;
	wire [16-1:0] node8905;
	wire [16-1:0] node8908;
	wire [16-1:0] node8909;
	wire [16-1:0] node8910;
	wire [16-1:0] node8911;
	wire [16-1:0] node8912;
	wire [16-1:0] node8915;
	wire [16-1:0] node8918;
	wire [16-1:0] node8921;
	wire [16-1:0] node8924;
	wire [16-1:0] node8925;
	wire [16-1:0] node8926;
	wire [16-1:0] node8928;
	wire [16-1:0] node8931;
	wire [16-1:0] node8934;
	wire [16-1:0] node8935;
	wire [16-1:0] node8937;
	wire [16-1:0] node8940;
	wire [16-1:0] node8941;
	wire [16-1:0] node8943;
	wire [16-1:0] node8944;
	wire [16-1:0] node8948;
	wire [16-1:0] node8951;
	wire [16-1:0] node8952;
	wire [16-1:0] node8953;
	wire [16-1:0] node8954;
	wire [16-1:0] node8955;
	wire [16-1:0] node8956;
	wire [16-1:0] node8957;
	wire [16-1:0] node8958;
	wire [16-1:0] node8959;
	wire [16-1:0] node8960;
	wire [16-1:0] node8961;
	wire [16-1:0] node8965;
	wire [16-1:0] node8966;
	wire [16-1:0] node8968;
	wire [16-1:0] node8971;
	wire [16-1:0] node8974;
	wire [16-1:0] node8975;
	wire [16-1:0] node8976;
	wire [16-1:0] node8979;
	wire [16-1:0] node8981;
	wire [16-1:0] node8984;
	wire [16-1:0] node8987;
	wire [16-1:0] node8988;
	wire [16-1:0] node8990;
	wire [16-1:0] node8991;
	wire [16-1:0] node8993;
	wire [16-1:0] node8997;
	wire [16-1:0] node8999;
	wire [16-1:0] node9001;
	wire [16-1:0] node9004;
	wire [16-1:0] node9005;
	wire [16-1:0] node9006;
	wire [16-1:0] node9007;
	wire [16-1:0] node9010;
	wire [16-1:0] node9012;
	wire [16-1:0] node9015;
	wire [16-1:0] node9016;
	wire [16-1:0] node9019;
	wire [16-1:0] node9021;
	wire [16-1:0] node9023;
	wire [16-1:0] node9026;
	wire [16-1:0] node9027;
	wire [16-1:0] node9028;
	wire [16-1:0] node9030;
	wire [16-1:0] node9033;
	wire [16-1:0] node9034;
	wire [16-1:0] node9038;
	wire [16-1:0] node9040;
	wire [16-1:0] node9041;
	wire [16-1:0] node9043;
	wire [16-1:0] node9047;
	wire [16-1:0] node9048;
	wire [16-1:0] node9049;
	wire [16-1:0] node9050;
	wire [16-1:0] node9051;
	wire [16-1:0] node9053;
	wire [16-1:0] node9056;
	wire [16-1:0] node9057;
	wire [16-1:0] node9058;
	wire [16-1:0] node9060;
	wire [16-1:0] node9065;
	wire [16-1:0] node9066;
	wire [16-1:0] node9067;
	wire [16-1:0] node9071;
	wire [16-1:0] node9072;
	wire [16-1:0] node9074;
	wire [16-1:0] node9075;
	wire [16-1:0] node9080;
	wire [16-1:0] node9081;
	wire [16-1:0] node9083;
	wire [16-1:0] node9084;
	wire [16-1:0] node9086;
	wire [16-1:0] node9090;
	wire [16-1:0] node9091;
	wire [16-1:0] node9092;
	wire [16-1:0] node9095;
	wire [16-1:0] node9098;
	wire [16-1:0] node9100;
	wire [16-1:0] node9103;
	wire [16-1:0] node9104;
	wire [16-1:0] node9105;
	wire [16-1:0] node9106;
	wire [16-1:0] node9107;
	wire [16-1:0] node9112;
	wire [16-1:0] node9114;
	wire [16-1:0] node9115;
	wire [16-1:0] node9116;
	wire [16-1:0] node9118;
	wire [16-1:0] node9122;
	wire [16-1:0] node9125;
	wire [16-1:0] node9126;
	wire [16-1:0] node9127;
	wire [16-1:0] node9128;
	wire [16-1:0] node9131;
	wire [16-1:0] node9134;
	wire [16-1:0] node9135;
	wire [16-1:0] node9136;
	wire [16-1:0] node9138;
	wire [16-1:0] node9143;
	wire [16-1:0] node9144;
	wire [16-1:0] node9145;
	wire [16-1:0] node9150;
	wire [16-1:0] node9151;
	wire [16-1:0] node9152;
	wire [16-1:0] node9153;
	wire [16-1:0] node9154;
	wire [16-1:0] node9155;
	wire [16-1:0] node9156;
	wire [16-1:0] node9158;
	wire [16-1:0] node9159;
	wire [16-1:0] node9163;
	wire [16-1:0] node9167;
	wire [16-1:0] node9168;
	wire [16-1:0] node9171;
	wire [16-1:0] node9174;
	wire [16-1:0] node9175;
	wire [16-1:0] node9176;
	wire [16-1:0] node9178;
	wire [16-1:0] node9181;
	wire [16-1:0] node9184;
	wire [16-1:0] node9185;
	wire [16-1:0] node9187;
	wire [16-1:0] node9190;
	wire [16-1:0] node9193;
	wire [16-1:0] node9194;
	wire [16-1:0] node9195;
	wire [16-1:0] node9196;
	wire [16-1:0] node9197;
	wire [16-1:0] node9201;
	wire [16-1:0] node9202;
	wire [16-1:0] node9203;
	wire [16-1:0] node9207;
	wire [16-1:0] node9208;
	wire [16-1:0] node9212;
	wire [16-1:0] node9213;
	wire [16-1:0] node9214;
	wire [16-1:0] node9217;
	wire [16-1:0] node9220;
	wire [16-1:0] node9221;
	wire [16-1:0] node9223;
	wire [16-1:0] node9224;
	wire [16-1:0] node9229;
	wire [16-1:0] node9230;
	wire [16-1:0] node9231;
	wire [16-1:0] node9234;
	wire [16-1:0] node9236;
	wire [16-1:0] node9239;
	wire [16-1:0] node9240;
	wire [16-1:0] node9241;
	wire [16-1:0] node9246;
	wire [16-1:0] node9247;
	wire [16-1:0] node9248;
	wire [16-1:0] node9249;
	wire [16-1:0] node9250;
	wire [16-1:0] node9252;
	wire [16-1:0] node9255;
	wire [16-1:0] node9256;
	wire [16-1:0] node9259;
	wire [16-1:0] node9262;
	wire [16-1:0] node9263;
	wire [16-1:0] node9265;
	wire [16-1:0] node9266;
	wire [16-1:0] node9268;
	wire [16-1:0] node9272;
	wire [16-1:0] node9273;
	wire [16-1:0] node9276;
	wire [16-1:0] node9279;
	wire [16-1:0] node9280;
	wire [16-1:0] node9281;
	wire [16-1:0] node9285;
	wire [16-1:0] node9286;
	wire [16-1:0] node9287;
	wire [16-1:0] node9288;
	wire [16-1:0] node9292;
	wire [16-1:0] node9295;
	wire [16-1:0] node9298;
	wire [16-1:0] node9299;
	wire [16-1:0] node9300;
	wire [16-1:0] node9301;
	wire [16-1:0] node9304;
	wire [16-1:0] node9305;
	wire [16-1:0] node9309;
	wire [16-1:0] node9310;
	wire [16-1:0] node9311;
	wire [16-1:0] node9314;
	wire [16-1:0] node9317;
	wire [16-1:0] node9318;
	wire [16-1:0] node9321;
	wire [16-1:0] node9324;
	wire [16-1:0] node9325;
	wire [16-1:0] node9326;
	wire [16-1:0] node9327;
	wire [16-1:0] node9332;
	wire [16-1:0] node9333;
	wire [16-1:0] node9335;
	wire [16-1:0] node9339;
	wire [16-1:0] node9340;
	wire [16-1:0] node9341;
	wire [16-1:0] node9342;
	wire [16-1:0] node9343;
	wire [16-1:0] node9344;
	wire [16-1:0] node9345;
	wire [16-1:0] node9348;
	wire [16-1:0] node9350;
	wire [16-1:0] node9353;
	wire [16-1:0] node9355;
	wire [16-1:0] node9356;
	wire [16-1:0] node9359;
	wire [16-1:0] node9362;
	wire [16-1:0] node9363;
	wire [16-1:0] node9364;
	wire [16-1:0] node9366;
	wire [16-1:0] node9369;
	wire [16-1:0] node9372;
	wire [16-1:0] node9373;
	wire [16-1:0] node9374;
	wire [16-1:0] node9376;
	wire [16-1:0] node9381;
	wire [16-1:0] node9382;
	wire [16-1:0] node9383;
	wire [16-1:0] node9384;
	wire [16-1:0] node9387;
	wire [16-1:0] node9388;
	wire [16-1:0] node9390;
	wire [16-1:0] node9391;
	wire [16-1:0] node9395;
	wire [16-1:0] node9398;
	wire [16-1:0] node9400;
	wire [16-1:0] node9402;
	wire [16-1:0] node9405;
	wire [16-1:0] node9406;
	wire [16-1:0] node9407;
	wire [16-1:0] node9409;
	wire [16-1:0] node9412;
	wire [16-1:0] node9413;
	wire [16-1:0] node9417;
	wire [16-1:0] node9418;
	wire [16-1:0] node9419;
	wire [16-1:0] node9423;
	wire [16-1:0] node9426;
	wire [16-1:0] node9427;
	wire [16-1:0] node9428;
	wire [16-1:0] node9429;
	wire [16-1:0] node9430;
	wire [16-1:0] node9432;
	wire [16-1:0] node9433;
	wire [16-1:0] node9437;
	wire [16-1:0] node9438;
	wire [16-1:0] node9440;
	wire [16-1:0] node9443;
	wire [16-1:0] node9445;
	wire [16-1:0] node9448;
	wire [16-1:0] node9449;
	wire [16-1:0] node9450;
	wire [16-1:0] node9453;
	wire [16-1:0] node9456;
	wire [16-1:0] node9459;
	wire [16-1:0] node9460;
	wire [16-1:0] node9461;
	wire [16-1:0] node9462;
	wire [16-1:0] node9466;
	wire [16-1:0] node9468;
	wire [16-1:0] node9470;
	wire [16-1:0] node9473;
	wire [16-1:0] node9474;
	wire [16-1:0] node9477;
	wire [16-1:0] node9479;
	wire [16-1:0] node9482;
	wire [16-1:0] node9483;
	wire [16-1:0] node9484;
	wire [16-1:0] node9485;
	wire [16-1:0] node9489;
	wire [16-1:0] node9490;
	wire [16-1:0] node9493;
	wire [16-1:0] node9494;
	wire [16-1:0] node9498;
	wire [16-1:0] node9499;
	wire [16-1:0] node9501;
	wire [16-1:0] node9504;
	wire [16-1:0] node9506;
	wire [16-1:0] node9508;
	wire [16-1:0] node9511;
	wire [16-1:0] node9512;
	wire [16-1:0] node9513;
	wire [16-1:0] node9514;
	wire [16-1:0] node9515;
	wire [16-1:0] node9516;
	wire [16-1:0] node9517;
	wire [16-1:0] node9522;
	wire [16-1:0] node9523;
	wire [16-1:0] node9524;
	wire [16-1:0] node9525;
	wire [16-1:0] node9527;
	wire [16-1:0] node9532;
	wire [16-1:0] node9534;
	wire [16-1:0] node9537;
	wire [16-1:0] node9538;
	wire [16-1:0] node9540;
	wire [16-1:0] node9541;
	wire [16-1:0] node9544;
	wire [16-1:0] node9546;
	wire [16-1:0] node9549;
	wire [16-1:0] node9550;
	wire [16-1:0] node9554;
	wire [16-1:0] node9555;
	wire [16-1:0] node9556;
	wire [16-1:0] node9557;
	wire [16-1:0] node9560;
	wire [16-1:0] node9561;
	wire [16-1:0] node9565;
	wire [16-1:0] node9566;
	wire [16-1:0] node9567;
	wire [16-1:0] node9570;
	wire [16-1:0] node9573;
	wire [16-1:0] node9575;
	wire [16-1:0] node9578;
	wire [16-1:0] node9579;
	wire [16-1:0] node9580;
	wire [16-1:0] node9581;
	wire [16-1:0] node9585;
	wire [16-1:0] node9587;
	wire [16-1:0] node9590;
	wire [16-1:0] node9591;
	wire [16-1:0] node9594;
	wire [16-1:0] node9596;
	wire [16-1:0] node9599;
	wire [16-1:0] node9600;
	wire [16-1:0] node9601;
	wire [16-1:0] node9602;
	wire [16-1:0] node9603;
	wire [16-1:0] node9604;
	wire [16-1:0] node9608;
	wire [16-1:0] node9610;
	wire [16-1:0] node9613;
	wire [16-1:0] node9614;
	wire [16-1:0] node9616;
	wire [16-1:0] node9617;
	wire [16-1:0] node9619;
	wire [16-1:0] node9623;
	wire [16-1:0] node9626;
	wire [16-1:0] node9627;
	wire [16-1:0] node9629;
	wire [16-1:0] node9630;
	wire [16-1:0] node9634;
	wire [16-1:0] node9635;
	wire [16-1:0] node9637;
	wire [16-1:0] node9640;
	wire [16-1:0] node9641;
	wire [16-1:0] node9645;
	wire [16-1:0] node9646;
	wire [16-1:0] node9647;
	wire [16-1:0] node9648;
	wire [16-1:0] node9651;
	wire [16-1:0] node9652;
	wire [16-1:0] node9656;
	wire [16-1:0] node9657;
	wire [16-1:0] node9658;
	wire [16-1:0] node9661;
	wire [16-1:0] node9664;
	wire [16-1:0] node9666;
	wire [16-1:0] node9667;
	wire [16-1:0] node9671;
	wire [16-1:0] node9672;
	wire [16-1:0] node9674;
	wire [16-1:0] node9675;
	wire [16-1:0] node9678;
	wire [16-1:0] node9681;
	wire [16-1:0] node9682;
	wire [16-1:0] node9683;
	wire [16-1:0] node9686;
	wire [16-1:0] node9689;
	wire [16-1:0] node9691;
	wire [16-1:0] node9694;
	wire [16-1:0] node9695;
	wire [16-1:0] node9696;
	wire [16-1:0] node9697;
	wire [16-1:0] node9698;
	wire [16-1:0] node9699;
	wire [16-1:0] node9700;
	wire [16-1:0] node9701;
	wire [16-1:0] node9705;
	wire [16-1:0] node9706;
	wire [16-1:0] node9707;
	wire [16-1:0] node9711;
	wire [16-1:0] node9713;
	wire [16-1:0] node9716;
	wire [16-1:0] node9717;
	wire [16-1:0] node9718;
	wire [16-1:0] node9719;
	wire [16-1:0] node9720;
	wire [16-1:0] node9722;
	wire [16-1:0] node9726;
	wire [16-1:0] node9729;
	wire [16-1:0] node9731;
	wire [16-1:0] node9734;
	wire [16-1:0] node9736;
	wire [16-1:0] node9737;
	wire [16-1:0] node9738;
	wire [16-1:0] node9739;
	wire [16-1:0] node9743;
	wire [16-1:0] node9744;
	wire [16-1:0] node9749;
	wire [16-1:0] node9750;
	wire [16-1:0] node9751;
	wire [16-1:0] node9752;
	wire [16-1:0] node9754;
	wire [16-1:0] node9759;
	wire [16-1:0] node9760;
	wire [16-1:0] node9762;
	wire [16-1:0] node9763;
	wire [16-1:0] node9765;
	wire [16-1:0] node9768;
	wire [16-1:0] node9771;
	wire [16-1:0] node9772;
	wire [16-1:0] node9774;
	wire [16-1:0] node9776;
	wire [16-1:0] node9779;
	wire [16-1:0] node9780;
	wire [16-1:0] node9784;
	wire [16-1:0] node9785;
	wire [16-1:0] node9786;
	wire [16-1:0] node9787;
	wire [16-1:0] node9788;
	wire [16-1:0] node9792;
	wire [16-1:0] node9793;
	wire [16-1:0] node9794;
	wire [16-1:0] node9795;
	wire [16-1:0] node9800;
	wire [16-1:0] node9803;
	wire [16-1:0] node9804;
	wire [16-1:0] node9805;
	wire [16-1:0] node9807;
	wire [16-1:0] node9808;
	wire [16-1:0] node9812;
	wire [16-1:0] node9813;
	wire [16-1:0] node9816;
	wire [16-1:0] node9819;
	wire [16-1:0] node9822;
	wire [16-1:0] node9823;
	wire [16-1:0] node9824;
	wire [16-1:0] node9825;
	wire [16-1:0] node9829;
	wire [16-1:0] node9830;
	wire [16-1:0] node9833;
	wire [16-1:0] node9834;
	wire [16-1:0] node9838;
	wire [16-1:0] node9839;
	wire [16-1:0] node9840;
	wire [16-1:0] node9843;
	wire [16-1:0] node9846;
	wire [16-1:0] node9847;
	wire [16-1:0] node9850;
	wire [16-1:0] node9853;
	wire [16-1:0] node9854;
	wire [16-1:0] node9855;
	wire [16-1:0] node9856;
	wire [16-1:0] node9857;
	wire [16-1:0] node9859;
	wire [16-1:0] node9860;
	wire [16-1:0] node9864;
	wire [16-1:0] node9865;
	wire [16-1:0] node9866;
	wire [16-1:0] node9869;
	wire [16-1:0] node9872;
	wire [16-1:0] node9873;
	wire [16-1:0] node9877;
	wire [16-1:0] node9878;
	wire [16-1:0] node9879;
	wire [16-1:0] node9881;
	wire [16-1:0] node9885;
	wire [16-1:0] node9887;
	wire [16-1:0] node9888;
	wire [16-1:0] node9892;
	wire [16-1:0] node9893;
	wire [16-1:0] node9894;
	wire [16-1:0] node9895;
	wire [16-1:0] node9896;
	wire [16-1:0] node9899;
	wire [16-1:0] node9902;
	wire [16-1:0] node9905;
	wire [16-1:0] node9907;
	wire [16-1:0] node9908;
	wire [16-1:0] node9912;
	wire [16-1:0] node9913;
	wire [16-1:0] node9914;
	wire [16-1:0] node9915;
	wire [16-1:0] node9919;
	wire [16-1:0] node9921;
	wire [16-1:0] node9924;
	wire [16-1:0] node9925;
	wire [16-1:0] node9929;
	wire [16-1:0] node9930;
	wire [16-1:0] node9931;
	wire [16-1:0] node9932;
	wire [16-1:0] node9934;
	wire [16-1:0] node9937;
	wire [16-1:0] node9938;
	wire [16-1:0] node9939;
	wire [16-1:0] node9942;
	wire [16-1:0] node9945;
	wire [16-1:0] node9946;
	wire [16-1:0] node9950;
	wire [16-1:0] node9951;
	wire [16-1:0] node9952;
	wire [16-1:0] node9953;
	wire [16-1:0] node9956;
	wire [16-1:0] node9959;
	wire [16-1:0] node9960;
	wire [16-1:0] node9963;
	wire [16-1:0] node9966;
	wire [16-1:0] node9968;
	wire [16-1:0] node9969;
	wire [16-1:0] node9972;
	wire [16-1:0] node9973;
	wire [16-1:0] node9977;
	wire [16-1:0] node9978;
	wire [16-1:0] node9979;
	wire [16-1:0] node9980;
	wire [16-1:0] node9984;
	wire [16-1:0] node9985;
	wire [16-1:0] node9988;
	wire [16-1:0] node9991;
	wire [16-1:0] node9992;
	wire [16-1:0] node9993;
	wire [16-1:0] node9996;
	wire [16-1:0] node9998;
	wire [16-1:0] node10001;
	wire [16-1:0] node10002;
	wire [16-1:0] node10004;
	wire [16-1:0] node10007;
	wire [16-1:0] node10008;
	wire [16-1:0] node10012;
	wire [16-1:0] node10013;
	wire [16-1:0] node10014;
	wire [16-1:0] node10015;
	wire [16-1:0] node10016;
	wire [16-1:0] node10017;
	wire [16-1:0] node10018;
	wire [16-1:0] node10020;
	wire [16-1:0] node10023;
	wire [16-1:0] node10024;
	wire [16-1:0] node10027;
	wire [16-1:0] node10030;
	wire [16-1:0] node10032;
	wire [16-1:0] node10033;
	wire [16-1:0] node10034;
	wire [16-1:0] node10036;
	wire [16-1:0] node10040;
	wire [16-1:0] node10043;
	wire [16-1:0] node10044;
	wire [16-1:0] node10046;
	wire [16-1:0] node10047;
	wire [16-1:0] node10050;
	wire [16-1:0] node10052;
	wire [16-1:0] node10055;
	wire [16-1:0] node10056;
	wire [16-1:0] node10059;
	wire [16-1:0] node10062;
	wire [16-1:0] node10063;
	wire [16-1:0] node10064;
	wire [16-1:0] node10065;
	wire [16-1:0] node10069;
	wire [16-1:0] node10070;
	wire [16-1:0] node10072;
	wire [16-1:0] node10076;
	wire [16-1:0] node10077;
	wire [16-1:0] node10078;
	wire [16-1:0] node10079;
	wire [16-1:0] node10084;
	wire [16-1:0] node10085;
	wire [16-1:0] node10087;
	wire [16-1:0] node10091;
	wire [16-1:0] node10092;
	wire [16-1:0] node10093;
	wire [16-1:0] node10094;
	wire [16-1:0] node10095;
	wire [16-1:0] node10096;
	wire [16-1:0] node10101;
	wire [16-1:0] node10102;
	wire [16-1:0] node10104;
	wire [16-1:0] node10106;
	wire [16-1:0] node10109;
	wire [16-1:0] node10110;
	wire [16-1:0] node10113;
	wire [16-1:0] node10114;
	wire [16-1:0] node10118;
	wire [16-1:0] node10119;
	wire [16-1:0] node10120;
	wire [16-1:0] node10122;
	wire [16-1:0] node10125;
	wire [16-1:0] node10126;
	wire [16-1:0] node10127;
	wire [16-1:0] node10130;
	wire [16-1:0] node10132;
	wire [16-1:0] node10136;
	wire [16-1:0] node10139;
	wire [16-1:0] node10140;
	wire [16-1:0] node10141;
	wire [16-1:0] node10142;
	wire [16-1:0] node10145;
	wire [16-1:0] node10146;
	wire [16-1:0] node10150;
	wire [16-1:0] node10151;
	wire [16-1:0] node10152;
	wire [16-1:0] node10156;
	wire [16-1:0] node10158;
	wire [16-1:0] node10160;
	wire [16-1:0] node10163;
	wire [16-1:0] node10164;
	wire [16-1:0] node10166;
	wire [16-1:0] node10167;
	wire [16-1:0] node10171;
	wire [16-1:0] node10172;
	wire [16-1:0] node10175;
	wire [16-1:0] node10177;
	wire [16-1:0] node10180;
	wire [16-1:0] node10181;
	wire [16-1:0] node10182;
	wire [16-1:0] node10183;
	wire [16-1:0] node10184;
	wire [16-1:0] node10186;
	wire [16-1:0] node10187;
	wire [16-1:0] node10190;
	wire [16-1:0] node10192;
	wire [16-1:0] node10195;
	wire [16-1:0] node10196;
	wire [16-1:0] node10199;
	wire [16-1:0] node10200;
	wire [16-1:0] node10204;
	wire [16-1:0] node10205;
	wire [16-1:0] node10207;
	wire [16-1:0] node10208;
	wire [16-1:0] node10212;
	wire [16-1:0] node10213;
	wire [16-1:0] node10214;
	wire [16-1:0] node10217;
	wire [16-1:0] node10220;
	wire [16-1:0] node10221;
	wire [16-1:0] node10224;
	wire [16-1:0] node10227;
	wire [16-1:0] node10228;
	wire [16-1:0] node10229;
	wire [16-1:0] node10231;
	wire [16-1:0] node10233;
	wire [16-1:0] node10234;
	wire [16-1:0] node10238;
	wire [16-1:0] node10239;
	wire [16-1:0] node10241;
	wire [16-1:0] node10242;
	wire [16-1:0] node10244;
	wire [16-1:0] node10248;
	wire [16-1:0] node10249;
	wire [16-1:0] node10252;
	wire [16-1:0] node10254;
	wire [16-1:0] node10257;
	wire [16-1:0] node10258;
	wire [16-1:0] node10260;
	wire [16-1:0] node10261;
	wire [16-1:0] node10264;
	wire [16-1:0] node10267;
	wire [16-1:0] node10268;
	wire [16-1:0] node10270;
	wire [16-1:0] node10273;
	wire [16-1:0] node10275;
	wire [16-1:0] node10276;
	wire [16-1:0] node10280;
	wire [16-1:0] node10281;
	wire [16-1:0] node10282;
	wire [16-1:0] node10283;
	wire [16-1:0] node10284;
	wire [16-1:0] node10285;
	wire [16-1:0] node10288;
	wire [16-1:0] node10289;
	wire [16-1:0] node10293;
	wire [16-1:0] node10295;
	wire [16-1:0] node10298;
	wire [16-1:0] node10299;
	wire [16-1:0] node10300;
	wire [16-1:0] node10303;
	wire [16-1:0] node10307;
	wire [16-1:0] node10308;
	wire [16-1:0] node10310;
	wire [16-1:0] node10313;
	wire [16-1:0] node10314;
	wire [16-1:0] node10315;
	wire [16-1:0] node10318;
	wire [16-1:0] node10320;
	wire [16-1:0] node10323;
	wire [16-1:0] node10324;
	wire [16-1:0] node10327;
	wire [16-1:0] node10330;
	wire [16-1:0] node10331;
	wire [16-1:0] node10332;
	wire [16-1:0] node10333;
	wire [16-1:0] node10334;
	wire [16-1:0] node10337;
	wire [16-1:0] node10339;
	wire [16-1:0] node10342;
	wire [16-1:0] node10344;
	wire [16-1:0] node10347;
	wire [16-1:0] node10348;
	wire [16-1:0] node10350;
	wire [16-1:0] node10353;
	wire [16-1:0] node10356;
	wire [16-1:0] node10357;
	wire [16-1:0] node10358;
	wire [16-1:0] node10360;
	wire [16-1:0] node10363;
	wire [16-1:0] node10364;
	wire [16-1:0] node10366;
	wire [16-1:0] node10367;
	wire [16-1:0] node10372;
	wire [16-1:0] node10373;
	wire [16-1:0] node10374;
	wire [16-1:0] node10375;
	wire [16-1:0] node10380;
	wire [16-1:0] node10381;
	wire [16-1:0] node10382;
	wire [16-1:0] node10386;
	wire [16-1:0] node10389;
	wire [16-1:0] node10390;
	wire [16-1:0] node10391;
	wire [16-1:0] node10392;
	wire [16-1:0] node10393;
	wire [16-1:0] node10394;
	wire [16-1:0] node10395;
	wire [16-1:0] node10396;
	wire [16-1:0] node10398;
	wire [16-1:0] node10399;
	wire [16-1:0] node10403;
	wire [16-1:0] node10404;
	wire [16-1:0] node10405;
	wire [16-1:0] node10408;
	wire [16-1:0] node10411;
	wire [16-1:0] node10412;
	wire [16-1:0] node10416;
	wire [16-1:0] node10417;
	wire [16-1:0] node10418;
	wire [16-1:0] node10419;
	wire [16-1:0] node10422;
	wire [16-1:0] node10423;
	wire [16-1:0] node10425;
	wire [16-1:0] node10430;
	wire [16-1:0] node10431;
	wire [16-1:0] node10432;
	wire [16-1:0] node10435;
	wire [16-1:0] node10439;
	wire [16-1:0] node10440;
	wire [16-1:0] node10441;
	wire [16-1:0] node10442;
	wire [16-1:0] node10444;
	wire [16-1:0] node10447;
	wire [16-1:0] node10448;
	wire [16-1:0] node10452;
	wire [16-1:0] node10453;
	wire [16-1:0] node10455;
	wire [16-1:0] node10458;
	wire [16-1:0] node10459;
	wire [16-1:0] node10462;
	wire [16-1:0] node10465;
	wire [16-1:0] node10466;
	wire [16-1:0] node10467;
	wire [16-1:0] node10470;
	wire [16-1:0] node10471;
	wire [16-1:0] node10473;
	wire [16-1:0] node10474;
	wire [16-1:0] node10478;
	wire [16-1:0] node10480;
	wire [16-1:0] node10483;
	wire [16-1:0] node10484;
	wire [16-1:0] node10486;
	wire [16-1:0] node10489;
	wire [16-1:0] node10490;
	wire [16-1:0] node10493;
	wire [16-1:0] node10495;
	wire [16-1:0] node10498;
	wire [16-1:0] node10499;
	wire [16-1:0] node10500;
	wire [16-1:0] node10501;
	wire [16-1:0] node10503;
	wire [16-1:0] node10506;
	wire [16-1:0] node10507;
	wire [16-1:0] node10509;
	wire [16-1:0] node10512;
	wire [16-1:0] node10513;
	wire [16-1:0] node10516;
	wire [16-1:0] node10518;
	wire [16-1:0] node10520;
	wire [16-1:0] node10523;
	wire [16-1:0] node10524;
	wire [16-1:0] node10525;
	wire [16-1:0] node10527;
	wire [16-1:0] node10531;
	wire [16-1:0] node10533;
	wire [16-1:0] node10534;
	wire [16-1:0] node10536;
	wire [16-1:0] node10540;
	wire [16-1:0] node10541;
	wire [16-1:0] node10542;
	wire [16-1:0] node10543;
	wire [16-1:0] node10546;
	wire [16-1:0] node10547;
	wire [16-1:0] node10550;
	wire [16-1:0] node10553;
	wire [16-1:0] node10554;
	wire [16-1:0] node10556;
	wire [16-1:0] node10559;
	wire [16-1:0] node10562;
	wire [16-1:0] node10563;
	wire [16-1:0] node10565;
	wire [16-1:0] node10568;
	wire [16-1:0] node10570;
	wire [16-1:0] node10571;
	wire [16-1:0] node10575;
	wire [16-1:0] node10576;
	wire [16-1:0] node10577;
	wire [16-1:0] node10578;
	wire [16-1:0] node10579;
	wire [16-1:0] node10582;
	wire [16-1:0] node10584;
	wire [16-1:0] node10585;
	wire [16-1:0] node10589;
	wire [16-1:0] node10590;
	wire [16-1:0] node10591;
	wire [16-1:0] node10594;
	wire [16-1:0] node10595;
	wire [16-1:0] node10599;
	wire [16-1:0] node10601;
	wire [16-1:0] node10604;
	wire [16-1:0] node10605;
	wire [16-1:0] node10606;
	wire [16-1:0] node10607;
	wire [16-1:0] node10608;
	wire [16-1:0] node10610;
	wire [16-1:0] node10613;
	wire [16-1:0] node10615;
	wire [16-1:0] node10618;
	wire [16-1:0] node10619;
	wire [16-1:0] node10623;
	wire [16-1:0] node10624;
	wire [16-1:0] node10625;
	wire [16-1:0] node10628;
	wire [16-1:0] node10631;
	wire [16-1:0] node10632;
	wire [16-1:0] node10635;
	wire [16-1:0] node10638;
	wire [16-1:0] node10639;
	wire [16-1:0] node10641;
	wire [16-1:0] node10644;
	wire [16-1:0] node10646;
	wire [16-1:0] node10648;
	wire [16-1:0] node10649;
	wire [16-1:0] node10653;
	wire [16-1:0] node10654;
	wire [16-1:0] node10655;
	wire [16-1:0] node10656;
	wire [16-1:0] node10657;
	wire [16-1:0] node10659;
	wire [16-1:0] node10663;
	wire [16-1:0] node10664;
	wire [16-1:0] node10665;
	wire [16-1:0] node10667;
	wire [16-1:0] node10670;
	wire [16-1:0] node10671;
	wire [16-1:0] node10676;
	wire [16-1:0] node10677;
	wire [16-1:0] node10679;
	wire [16-1:0] node10682;
	wire [16-1:0] node10684;
	wire [16-1:0] node10686;
	wire [16-1:0] node10689;
	wire [16-1:0] node10690;
	wire [16-1:0] node10691;
	wire [16-1:0] node10692;
	wire [16-1:0] node10694;
	wire [16-1:0] node10697;
	wire [16-1:0] node10698;
	wire [16-1:0] node10701;
	wire [16-1:0] node10704;
	wire [16-1:0] node10705;
	wire [16-1:0] node10706;
	wire [16-1:0] node10708;
	wire [16-1:0] node10712;
	wire [16-1:0] node10713;
	wire [16-1:0] node10717;
	wire [16-1:0] node10718;
	wire [16-1:0] node10720;
	wire [16-1:0] node10721;
	wire [16-1:0] node10724;
	wire [16-1:0] node10727;
	wire [16-1:0] node10728;
	wire [16-1:0] node10729;
	wire [16-1:0] node10730;
	wire [16-1:0] node10734;
	wire [16-1:0] node10737;
	wire [16-1:0] node10739;
	wire [16-1:0] node10741;
	wire [16-1:0] node10744;
	wire [16-1:0] node10745;
	wire [16-1:0] node10746;
	wire [16-1:0] node10747;
	wire [16-1:0] node10748;
	wire [16-1:0] node10749;
	wire [16-1:0] node10750;
	wire [16-1:0] node10751;
	wire [16-1:0] node10754;
	wire [16-1:0] node10757;
	wire [16-1:0] node10760;
	wire [16-1:0] node10761;
	wire [16-1:0] node10764;
	wire [16-1:0] node10767;
	wire [16-1:0] node10768;
	wire [16-1:0] node10769;
	wire [16-1:0] node10771;
	wire [16-1:0] node10774;
	wire [16-1:0] node10775;
	wire [16-1:0] node10779;
	wire [16-1:0] node10781;
	wire [16-1:0] node10783;
	wire [16-1:0] node10786;
	wire [16-1:0] node10787;
	wire [16-1:0] node10788;
	wire [16-1:0] node10789;
	wire [16-1:0] node10791;
	wire [16-1:0] node10794;
	wire [16-1:0] node10795;
	wire [16-1:0] node10796;
	wire [16-1:0] node10800;
	wire [16-1:0] node10803;
	wire [16-1:0] node10804;
	wire [16-1:0] node10805;
	wire [16-1:0] node10806;
	wire [16-1:0] node10810;
	wire [16-1:0] node10813;
	wire [16-1:0] node10815;
	wire [16-1:0] node10818;
	wire [16-1:0] node10819;
	wire [16-1:0] node10821;
	wire [16-1:0] node10823;
	wire [16-1:0] node10826;
	wire [16-1:0] node10827;
	wire [16-1:0] node10829;
	wire [16-1:0] node10832;
	wire [16-1:0] node10835;
	wire [16-1:0] node10836;
	wire [16-1:0] node10837;
	wire [16-1:0] node10838;
	wire [16-1:0] node10839;
	wire [16-1:0] node10842;
	wire [16-1:0] node10843;
	wire [16-1:0] node10844;
	wire [16-1:0] node10848;
	wire [16-1:0] node10850;
	wire [16-1:0] node10853;
	wire [16-1:0] node10855;
	wire [16-1:0] node10858;
	wire [16-1:0] node10859;
	wire [16-1:0] node10860;
	wire [16-1:0] node10863;
	wire [16-1:0] node10866;
	wire [16-1:0] node10867;
	wire [16-1:0] node10868;
	wire [16-1:0] node10871;
	wire [16-1:0] node10874;
	wire [16-1:0] node10876;
	wire [16-1:0] node10879;
	wire [16-1:0] node10880;
	wire [16-1:0] node10881;
	wire [16-1:0] node10882;
	wire [16-1:0] node10884;
	wire [16-1:0] node10887;
	wire [16-1:0] node10888;
	wire [16-1:0] node10891;
	wire [16-1:0] node10893;
	wire [16-1:0] node10896;
	wire [16-1:0] node10897;
	wire [16-1:0] node10899;
	wire [16-1:0] node10902;
	wire [16-1:0] node10904;
	wire [16-1:0] node10905;
	wire [16-1:0] node10907;
	wire [16-1:0] node10911;
	wire [16-1:0] node10912;
	wire [16-1:0] node10913;
	wire [16-1:0] node10914;
	wire [16-1:0] node10916;
	wire [16-1:0] node10920;
	wire [16-1:0] node10922;
	wire [16-1:0] node10925;
	wire [16-1:0] node10926;
	wire [16-1:0] node10928;
	wire [16-1:0] node10929;
	wire [16-1:0] node10933;
	wire [16-1:0] node10935;
	wire [16-1:0] node10938;
	wire [16-1:0] node10939;
	wire [16-1:0] node10940;
	wire [16-1:0] node10941;
	wire [16-1:0] node10942;
	wire [16-1:0] node10943;
	wire [16-1:0] node10944;
	wire [16-1:0] node10948;
	wire [16-1:0] node10950;
	wire [16-1:0] node10953;
	wire [16-1:0] node10954;
	wire [16-1:0] node10955;
	wire [16-1:0] node10958;
	wire [16-1:0] node10962;
	wire [16-1:0] node10963;
	wire [16-1:0] node10964;
	wire [16-1:0] node10966;
	wire [16-1:0] node10967;
	wire [16-1:0] node10969;
	wire [16-1:0] node10973;
	wire [16-1:0] node10974;
	wire [16-1:0] node10978;
	wire [16-1:0] node10980;
	wire [16-1:0] node10983;
	wire [16-1:0] node10984;
	wire [16-1:0] node10985;
	wire [16-1:0] node10986;
	wire [16-1:0] node10987;
	wire [16-1:0] node10990;
	wire [16-1:0] node10991;
	wire [16-1:0] node10994;
	wire [16-1:0] node10998;
	wire [16-1:0] node10999;
	wire [16-1:0] node11001;
	wire [16-1:0] node11003;
	wire [16-1:0] node11007;
	wire [16-1:0] node11008;
	wire [16-1:0] node11009;
	wire [16-1:0] node11011;
	wire [16-1:0] node11014;
	wire [16-1:0] node11016;
	wire [16-1:0] node11018;
	wire [16-1:0] node11021;
	wire [16-1:0] node11022;
	wire [16-1:0] node11024;
	wire [16-1:0] node11027;
	wire [16-1:0] node11029;
	wire [16-1:0] node11030;
	wire [16-1:0] node11034;
	wire [16-1:0] node11035;
	wire [16-1:0] node11036;
	wire [16-1:0] node11037;
	wire [16-1:0] node11038;
	wire [16-1:0] node11040;
	wire [16-1:0] node11043;
	wire [16-1:0] node11046;
	wire [16-1:0] node11047;
	wire [16-1:0] node11049;
	wire [16-1:0] node11052;
	wire [16-1:0] node11053;
	wire [16-1:0] node11054;
	wire [16-1:0] node11058;
	wire [16-1:0] node11061;
	wire [16-1:0] node11062;
	wire [16-1:0] node11063;
	wire [16-1:0] node11066;
	wire [16-1:0] node11068;
	wire [16-1:0] node11071;
	wire [16-1:0] node11074;
	wire [16-1:0] node11075;
	wire [16-1:0] node11076;
	wire [16-1:0] node11077;
	wire [16-1:0] node11079;
	wire [16-1:0] node11082;
	wire [16-1:0] node11083;
	wire [16-1:0] node11084;
	wire [16-1:0] node11089;
	wire [16-1:0] node11090;
	wire [16-1:0] node11093;
	wire [16-1:0] node11096;
	wire [16-1:0] node11097;
	wire [16-1:0] node11098;
	wire [16-1:0] node11101;
	wire [16-1:0] node11103;
	wire [16-1:0] node11106;
	wire [16-1:0] node11107;
	wire [16-1:0] node11108;
	wire [16-1:0] node11112;
	wire [16-1:0] node11114;
	wire [16-1:0] node11117;
	wire [16-1:0] node11118;
	wire [16-1:0] node11119;
	wire [16-1:0] node11120;
	wire [16-1:0] node11121;
	wire [16-1:0] node11122;
	wire [16-1:0] node11123;
	wire [16-1:0] node11124;
	wire [16-1:0] node11126;
	wire [16-1:0] node11129;
	wire [16-1:0] node11131;
	wire [16-1:0] node11134;
	wire [16-1:0] node11136;
	wire [16-1:0] node11137;
	wire [16-1:0] node11141;
	wire [16-1:0] node11142;
	wire [16-1:0] node11143;
	wire [16-1:0] node11145;
	wire [16-1:0] node11147;
	wire [16-1:0] node11148;
	wire [16-1:0] node11153;
	wire [16-1:0] node11154;
	wire [16-1:0] node11155;
	wire [16-1:0] node11158;
	wire [16-1:0] node11160;
	wire [16-1:0] node11163;
	wire [16-1:0] node11165;
	wire [16-1:0] node11168;
	wire [16-1:0] node11169;
	wire [16-1:0] node11170;
	wire [16-1:0] node11171;
	wire [16-1:0] node11173;
	wire [16-1:0] node11174;
	wire [16-1:0] node11175;
	wire [16-1:0] node11180;
	wire [16-1:0] node11182;
	wire [16-1:0] node11184;
	wire [16-1:0] node11187;
	wire [16-1:0] node11188;
	wire [16-1:0] node11190;
	wire [16-1:0] node11193;
	wire [16-1:0] node11196;
	wire [16-1:0] node11197;
	wire [16-1:0] node11199;
	wire [16-1:0] node11200;
	wire [16-1:0] node11201;
	wire [16-1:0] node11206;
	wire [16-1:0] node11208;
	wire [16-1:0] node11209;
	wire [16-1:0] node11211;
	wire [16-1:0] node11215;
	wire [16-1:0] node11216;
	wire [16-1:0] node11217;
	wire [16-1:0] node11218;
	wire [16-1:0] node11219;
	wire [16-1:0] node11221;
	wire [16-1:0] node11224;
	wire [16-1:0] node11226;
	wire [16-1:0] node11227;
	wire [16-1:0] node11228;
	wire [16-1:0] node11233;
	wire [16-1:0] node11234;
	wire [16-1:0] node11235;
	wire [16-1:0] node11240;
	wire [16-1:0] node11241;
	wire [16-1:0] node11242;
	wire [16-1:0] node11244;
	wire [16-1:0] node11247;
	wire [16-1:0] node11248;
	wire [16-1:0] node11249;
	wire [16-1:0] node11253;
	wire [16-1:0] node11256;
	wire [16-1:0] node11257;
	wire [16-1:0] node11259;
	wire [16-1:0] node11260;
	wire [16-1:0] node11265;
	wire [16-1:0] node11266;
	wire [16-1:0] node11268;
	wire [16-1:0] node11269;
	wire [16-1:0] node11270;
	wire [16-1:0] node11273;
	wire [16-1:0] node11276;
	wire [16-1:0] node11277;
	wire [16-1:0] node11280;
	wire [16-1:0] node11283;
	wire [16-1:0] node11284;
	wire [16-1:0] node11285;
	wire [16-1:0] node11286;
	wire [16-1:0] node11289;
	wire [16-1:0] node11291;
	wire [16-1:0] node11294;
	wire [16-1:0] node11295;
	wire [16-1:0] node11296;
	wire [16-1:0] node11298;
	wire [16-1:0] node11302;
	wire [16-1:0] node11305;
	wire [16-1:0] node11306;
	wire [16-1:0] node11307;
	wire [16-1:0] node11310;
	wire [16-1:0] node11312;
	wire [16-1:0] node11316;
	wire [16-1:0] node11317;
	wire [16-1:0] node11318;
	wire [16-1:0] node11319;
	wire [16-1:0] node11320;
	wire [16-1:0] node11321;
	wire [16-1:0] node11325;
	wire [16-1:0] node11326;
	wire [16-1:0] node11327;
	wire [16-1:0] node11330;
	wire [16-1:0] node11334;
	wire [16-1:0] node11335;
	wire [16-1:0] node11336;
	wire [16-1:0] node11339;
	wire [16-1:0] node11340;
	wire [16-1:0] node11344;
	wire [16-1:0] node11346;
	wire [16-1:0] node11349;
	wire [16-1:0] node11350;
	wire [16-1:0] node11351;
	wire [16-1:0] node11352;
	wire [16-1:0] node11353;
	wire [16-1:0] node11356;
	wire [16-1:0] node11359;
	wire [16-1:0] node11360;
	wire [16-1:0] node11363;
	wire [16-1:0] node11365;
	wire [16-1:0] node11368;
	wire [16-1:0] node11369;
	wire [16-1:0] node11371;
	wire [16-1:0] node11374;
	wire [16-1:0] node11375;
	wire [16-1:0] node11379;
	wire [16-1:0] node11380;
	wire [16-1:0] node11381;
	wire [16-1:0] node11382;
	wire [16-1:0] node11384;
	wire [16-1:0] node11389;
	wire [16-1:0] node11391;
	wire [16-1:0] node11392;
	wire [16-1:0] node11396;
	wire [16-1:0] node11397;
	wire [16-1:0] node11398;
	wire [16-1:0] node11399;
	wire [16-1:0] node11400;
	wire [16-1:0] node11402;
	wire [16-1:0] node11405;
	wire [16-1:0] node11409;
	wire [16-1:0] node11410;
	wire [16-1:0] node11411;
	wire [16-1:0] node11412;
	wire [16-1:0] node11414;
	wire [16-1:0] node11418;
	wire [16-1:0] node11419;
	wire [16-1:0] node11420;
	wire [16-1:0] node11424;
	wire [16-1:0] node11427;
	wire [16-1:0] node11428;
	wire [16-1:0] node11431;
	wire [16-1:0] node11433;
	wire [16-1:0] node11436;
	wire [16-1:0] node11437;
	wire [16-1:0] node11438;
	wire [16-1:0] node11439;
	wire [16-1:0] node11441;
	wire [16-1:0] node11443;
	wire [16-1:0] node11446;
	wire [16-1:0] node11448;
	wire [16-1:0] node11451;
	wire [16-1:0] node11452;
	wire [16-1:0] node11455;
	wire [16-1:0] node11457;
	wire [16-1:0] node11459;
	wire [16-1:0] node11462;
	wire [16-1:0] node11463;
	wire [16-1:0] node11464;
	wire [16-1:0] node11465;
	wire [16-1:0] node11468;
	wire [16-1:0] node11470;
	wire [16-1:0] node11473;
	wire [16-1:0] node11474;
	wire [16-1:0] node11475;
	wire [16-1:0] node11480;
	wire [16-1:0] node11481;
	wire [16-1:0] node11483;
	wire [16-1:0] node11485;
	wire [16-1:0] node11486;
	wire [16-1:0] node11490;
	wire [16-1:0] node11491;
	wire [16-1:0] node11492;
	wire [16-1:0] node11496;
	wire [16-1:0] node11498;
	wire [16-1:0] node11499;
	wire [16-1:0] node11503;
	wire [16-1:0] node11504;
	wire [16-1:0] node11505;
	wire [16-1:0] node11506;
	wire [16-1:0] node11507;
	wire [16-1:0] node11508;
	wire [16-1:0] node11509;
	wire [16-1:0] node11512;
	wire [16-1:0] node11513;
	wire [16-1:0] node11514;
	wire [16-1:0] node11519;
	wire [16-1:0] node11521;
	wire [16-1:0] node11522;
	wire [16-1:0] node11523;
	wire [16-1:0] node11528;
	wire [16-1:0] node11529;
	wire [16-1:0] node11530;
	wire [16-1:0] node11534;
	wire [16-1:0] node11535;
	wire [16-1:0] node11536;
	wire [16-1:0] node11539;
	wire [16-1:0] node11541;
	wire [16-1:0] node11544;
	wire [16-1:0] node11545;
	wire [16-1:0] node11548;
	wire [16-1:0] node11551;
	wire [16-1:0] node11552;
	wire [16-1:0] node11553;
	wire [16-1:0] node11555;
	wire [16-1:0] node11556;
	wire [16-1:0] node11559;
	wire [16-1:0] node11560;
	wire [16-1:0] node11561;
	wire [16-1:0] node11566;
	wire [16-1:0] node11567;
	wire [16-1:0] node11568;
	wire [16-1:0] node11571;
	wire [16-1:0] node11574;
	wire [16-1:0] node11575;
	wire [16-1:0] node11578;
	wire [16-1:0] node11580;
	wire [16-1:0] node11583;
	wire [16-1:0] node11584;
	wire [16-1:0] node11585;
	wire [16-1:0] node11586;
	wire [16-1:0] node11590;
	wire [16-1:0] node11592;
	wire [16-1:0] node11595;
	wire [16-1:0] node11596;
	wire [16-1:0] node11598;
	wire [16-1:0] node11599;
	wire [16-1:0] node11601;
	wire [16-1:0] node11605;
	wire [16-1:0] node11606;
	wire [16-1:0] node11610;
	wire [16-1:0] node11611;
	wire [16-1:0] node11612;
	wire [16-1:0] node11613;
	wire [16-1:0] node11614;
	wire [16-1:0] node11617;
	wire [16-1:0] node11618;
	wire [16-1:0] node11621;
	wire [16-1:0] node11624;
	wire [16-1:0] node11625;
	wire [16-1:0] node11626;
	wire [16-1:0] node11629;
	wire [16-1:0] node11632;
	wire [16-1:0] node11635;
	wire [16-1:0] node11636;
	wire [16-1:0] node11637;
	wire [16-1:0] node11639;
	wire [16-1:0] node11643;
	wire [16-1:0] node11644;
	wire [16-1:0] node11646;
	wire [16-1:0] node11649;
	wire [16-1:0] node11650;
	wire [16-1:0] node11654;
	wire [16-1:0] node11655;
	wire [16-1:0] node11656;
	wire [16-1:0] node11657;
	wire [16-1:0] node11658;
	wire [16-1:0] node11660;
	wire [16-1:0] node11663;
	wire [16-1:0] node11666;
	wire [16-1:0] node11667;
	wire [16-1:0] node11668;
	wire [16-1:0] node11672;
	wire [16-1:0] node11674;
	wire [16-1:0] node11677;
	wire [16-1:0] node11678;
	wire [16-1:0] node11679;
	wire [16-1:0] node11683;
	wire [16-1:0] node11684;
	wire [16-1:0] node11686;
	wire [16-1:0] node11690;
	wire [16-1:0] node11691;
	wire [16-1:0] node11692;
	wire [16-1:0] node11695;
	wire [16-1:0] node11697;
	wire [16-1:0] node11700;
	wire [16-1:0] node11701;
	wire [16-1:0] node11703;
	wire [16-1:0] node11705;
	wire [16-1:0] node11708;
	wire [16-1:0] node11710;
	wire [16-1:0] node11713;
	wire [16-1:0] node11714;
	wire [16-1:0] node11715;
	wire [16-1:0] node11716;
	wire [16-1:0] node11717;
	wire [16-1:0] node11718;
	wire [16-1:0] node11721;
	wire [16-1:0] node11722;
	wire [16-1:0] node11724;
	wire [16-1:0] node11725;
	wire [16-1:0] node11730;
	wire [16-1:0] node11731;
	wire [16-1:0] node11733;
	wire [16-1:0] node11736;
	wire [16-1:0] node11738;
	wire [16-1:0] node11741;
	wire [16-1:0] node11742;
	wire [16-1:0] node11743;
	wire [16-1:0] node11746;
	wire [16-1:0] node11748;
	wire [16-1:0] node11749;
	wire [16-1:0] node11750;
	wire [16-1:0] node11755;
	wire [16-1:0] node11756;
	wire [16-1:0] node11757;
	wire [16-1:0] node11758;
	wire [16-1:0] node11763;
	wire [16-1:0] node11765;
	wire [16-1:0] node11768;
	wire [16-1:0] node11769;
	wire [16-1:0] node11770;
	wire [16-1:0] node11772;
	wire [16-1:0] node11773;
	wire [16-1:0] node11777;
	wire [16-1:0] node11778;
	wire [16-1:0] node11780;
	wire [16-1:0] node11782;
	wire [16-1:0] node11783;
	wire [16-1:0] node11787;
	wire [16-1:0] node11790;
	wire [16-1:0] node11791;
	wire [16-1:0] node11792;
	wire [16-1:0] node11794;
	wire [16-1:0] node11795;
	wire [16-1:0] node11799;
	wire [16-1:0] node11800;
	wire [16-1:0] node11803;
	wire [16-1:0] node11806;
	wire [16-1:0] node11808;
	wire [16-1:0] node11809;
	wire [16-1:0] node11813;
	wire [16-1:0] node11814;
	wire [16-1:0] node11815;
	wire [16-1:0] node11816;
	wire [16-1:0] node11818;
	wire [16-1:0] node11821;
	wire [16-1:0] node11822;
	wire [16-1:0] node11823;
	wire [16-1:0] node11825;
	wire [16-1:0] node11828;
	wire [16-1:0] node11832;
	wire [16-1:0] node11833;
	wire [16-1:0] node11835;
	wire [16-1:0] node11836;
	wire [16-1:0] node11840;
	wire [16-1:0] node11841;
	wire [16-1:0] node11842;
	wire [16-1:0] node11846;
	wire [16-1:0] node11848;
	wire [16-1:0] node11849;
	wire [16-1:0] node11851;
	wire [16-1:0] node11855;
	wire [16-1:0] node11856;
	wire [16-1:0] node11857;
	wire [16-1:0] node11858;
	wire [16-1:0] node11859;
	wire [16-1:0] node11862;
	wire [16-1:0] node11865;
	wire [16-1:0] node11867;
	wire [16-1:0] node11869;
	wire [16-1:0] node11872;
	wire [16-1:0] node11873;
	wire [16-1:0] node11874;
	wire [16-1:0] node11878;
	wire [16-1:0] node11880;
	wire [16-1:0] node11882;
	wire [16-1:0] node11885;
	wire [16-1:0] node11886;
	wire [16-1:0] node11887;
	wire [16-1:0] node11889;
	wire [16-1:0] node11892;
	wire [16-1:0] node11894;
	wire [16-1:0] node11897;
	wire [16-1:0] node11898;
	wire [16-1:0] node11899;
	wire [16-1:0] node11902;
	wire [16-1:0] node11903;
	wire [16-1:0] node11905;
	wire [16-1:0] node11908;
	wire [16-1:0] node11911;
	wire [16-1:0] node11913;
	wire [16-1:0] node11916;
	wire [16-1:0] node11917;
	wire [16-1:0] node11918;
	wire [16-1:0] node11919;
	wire [16-1:0] node11920;
	wire [16-1:0] node11921;
	wire [16-1:0] node11922;
	wire [16-1:0] node11923;
	wire [16-1:0] node11924;
	wire [16-1:0] node11925;
	wire [16-1:0] node11926;
	wire [16-1:0] node11927;
	wire [16-1:0] node11928;
	wire [16-1:0] node11932;
	wire [16-1:0] node11933;
	wire [16-1:0] node11937;
	wire [16-1:0] node11938;
	wire [16-1:0] node11939;
	wire [16-1:0] node11943;
	wire [16-1:0] node11944;
	wire [16-1:0] node11945;
	wire [16-1:0] node11948;
	wire [16-1:0] node11952;
	wire [16-1:0] node11953;
	wire [16-1:0] node11955;
	wire [16-1:0] node11956;
	wire [16-1:0] node11957;
	wire [16-1:0] node11960;
	wire [16-1:0] node11961;
	wire [16-1:0] node11966;
	wire [16-1:0] node11969;
	wire [16-1:0] node11970;
	wire [16-1:0] node11971;
	wire [16-1:0] node11973;
	wire [16-1:0] node11974;
	wire [16-1:0] node11975;
	wire [16-1:0] node11976;
	wire [16-1:0] node11981;
	wire [16-1:0] node11984;
	wire [16-1:0] node11985;
	wire [16-1:0] node11987;
	wire [16-1:0] node11991;
	wire [16-1:0] node11992;
	wire [16-1:0] node11993;
	wire [16-1:0] node11996;
	wire [16-1:0] node11998;
	wire [16-1:0] node11999;
	wire [16-1:0] node12001;
	wire [16-1:0] node12005;
	wire [16-1:0] node12006;
	wire [16-1:0] node12007;
	wire [16-1:0] node12011;
	wire [16-1:0] node12012;
	wire [16-1:0] node12016;
	wire [16-1:0] node12017;
	wire [16-1:0] node12018;
	wire [16-1:0] node12019;
	wire [16-1:0] node12020;
	wire [16-1:0] node12021;
	wire [16-1:0] node12025;
	wire [16-1:0] node12026;
	wire [16-1:0] node12030;
	wire [16-1:0] node12032;
	wire [16-1:0] node12033;
	wire [16-1:0] node12034;
	wire [16-1:0] node12035;
	wire [16-1:0] node12039;
	wire [16-1:0] node12043;
	wire [16-1:0] node12044;
	wire [16-1:0] node12045;
	wire [16-1:0] node12046;
	wire [16-1:0] node12047;
	wire [16-1:0] node12049;
	wire [16-1:0] node12054;
	wire [16-1:0] node12055;
	wire [16-1:0] node12058;
	wire [16-1:0] node12061;
	wire [16-1:0] node12062;
	wire [16-1:0] node12064;
	wire [16-1:0] node12067;
	wire [16-1:0] node12068;
	wire [16-1:0] node12070;
	wire [16-1:0] node12074;
	wire [16-1:0] node12075;
	wire [16-1:0] node12076;
	wire [16-1:0] node12077;
	wire [16-1:0] node12078;
	wire [16-1:0] node12083;
	wire [16-1:0] node12084;
	wire [16-1:0] node12085;
	wire [16-1:0] node12090;
	wire [16-1:0] node12091;
	wire [16-1:0] node12092;
	wire [16-1:0] node12093;
	wire [16-1:0] node12095;
	wire [16-1:0] node12099;
	wire [16-1:0] node12101;
	wire [16-1:0] node12104;
	wire [16-1:0] node12105;
	wire [16-1:0] node12108;
	wire [16-1:0] node12109;
	wire [16-1:0] node12112;
	wire [16-1:0] node12115;
	wire [16-1:0] node12116;
	wire [16-1:0] node12117;
	wire [16-1:0] node12118;
	wire [16-1:0] node12119;
	wire [16-1:0] node12120;
	wire [16-1:0] node12121;
	wire [16-1:0] node12124;
	wire [16-1:0] node12126;
	wire [16-1:0] node12130;
	wire [16-1:0] node12131;
	wire [16-1:0] node12132;
	wire [16-1:0] node12133;
	wire [16-1:0] node12138;
	wire [16-1:0] node12139;
	wire [16-1:0] node12143;
	wire [16-1:0] node12144;
	wire [16-1:0] node12145;
	wire [16-1:0] node12146;
	wire [16-1:0] node12150;
	wire [16-1:0] node12151;
	wire [16-1:0] node12154;
	wire [16-1:0] node12157;
	wire [16-1:0] node12158;
	wire [16-1:0] node12159;
	wire [16-1:0] node12160;
	wire [16-1:0] node12164;
	wire [16-1:0] node12167;
	wire [16-1:0] node12168;
	wire [16-1:0] node12169;
	wire [16-1:0] node12171;
	wire [16-1:0] node12176;
	wire [16-1:0] node12177;
	wire [16-1:0] node12178;
	wire [16-1:0] node12179;
	wire [16-1:0] node12182;
	wire [16-1:0] node12183;
	wire [16-1:0] node12187;
	wire [16-1:0] node12188;
	wire [16-1:0] node12190;
	wire [16-1:0] node12194;
	wire [16-1:0] node12195;
	wire [16-1:0] node12196;
	wire [16-1:0] node12198;
	wire [16-1:0] node12199;
	wire [16-1:0] node12203;
	wire [16-1:0] node12204;
	wire [16-1:0] node12207;
	wire [16-1:0] node12210;
	wire [16-1:0] node12211;
	wire [16-1:0] node12213;
	wire [16-1:0] node12217;
	wire [16-1:0] node12218;
	wire [16-1:0] node12219;
	wire [16-1:0] node12220;
	wire [16-1:0] node12221;
	wire [16-1:0] node12224;
	wire [16-1:0] node12225;
	wire [16-1:0] node12227;
	wire [16-1:0] node12231;
	wire [16-1:0] node12232;
	wire [16-1:0] node12233;
	wire [16-1:0] node12236;
	wire [16-1:0] node12239;
	wire [16-1:0] node12242;
	wire [16-1:0] node12243;
	wire [16-1:0] node12245;
	wire [16-1:0] node12246;
	wire [16-1:0] node12249;
	wire [16-1:0] node12250;
	wire [16-1:0] node12254;
	wire [16-1:0] node12255;
	wire [16-1:0] node12259;
	wire [16-1:0] node12260;
	wire [16-1:0] node12261;
	wire [16-1:0] node12262;
	wire [16-1:0] node12266;
	wire [16-1:0] node12267;
	wire [16-1:0] node12271;
	wire [16-1:0] node12272;
	wire [16-1:0] node12274;
	wire [16-1:0] node12275;
	wire [16-1:0] node12277;
	wire [16-1:0] node12281;
	wire [16-1:0] node12282;
	wire [16-1:0] node12283;
	wire [16-1:0] node12286;
	wire [16-1:0] node12287;
	wire [16-1:0] node12289;
	wire [16-1:0] node12293;
	wire [16-1:0] node12295;
	wire [16-1:0] node12298;
	wire [16-1:0] node12299;
	wire [16-1:0] node12300;
	wire [16-1:0] node12301;
	wire [16-1:0] node12302;
	wire [16-1:0] node12303;
	wire [16-1:0] node12304;
	wire [16-1:0] node12306;
	wire [16-1:0] node12308;
	wire [16-1:0] node12309;
	wire [16-1:0] node12315;
	wire [16-1:0] node12316;
	wire [16-1:0] node12317;
	wire [16-1:0] node12318;
	wire [16-1:0] node12321;
	wire [16-1:0] node12323;
	wire [16-1:0] node12326;
	wire [16-1:0] node12327;
	wire [16-1:0] node12331;
	wire [16-1:0] node12333;
	wire [16-1:0] node12335;
	wire [16-1:0] node12338;
	wire [16-1:0] node12339;
	wire [16-1:0] node12340;
	wire [16-1:0] node12341;
	wire [16-1:0] node12342;
	wire [16-1:0] node12347;
	wire [16-1:0] node12349;
	wire [16-1:0] node12350;
	wire [16-1:0] node12352;
	wire [16-1:0] node12356;
	wire [16-1:0] node12357;
	wire [16-1:0] node12359;
	wire [16-1:0] node12362;
	wire [16-1:0] node12363;
	wire [16-1:0] node12365;
	wire [16-1:0] node12368;
	wire [16-1:0] node12369;
	wire [16-1:0] node12372;
	wire [16-1:0] node12375;
	wire [16-1:0] node12376;
	wire [16-1:0] node12377;
	wire [16-1:0] node12378;
	wire [16-1:0] node12380;
	wire [16-1:0] node12382;
	wire [16-1:0] node12385;
	wire [16-1:0] node12386;
	wire [16-1:0] node12387;
	wire [16-1:0] node12391;
	wire [16-1:0] node12392;
	wire [16-1:0] node12395;
	wire [16-1:0] node12398;
	wire [16-1:0] node12399;
	wire [16-1:0] node12401;
	wire [16-1:0] node12403;
	wire [16-1:0] node12404;
	wire [16-1:0] node12408;
	wire [16-1:0] node12410;
	wire [16-1:0] node12412;
	wire [16-1:0] node12415;
	wire [16-1:0] node12416;
	wire [16-1:0] node12417;
	wire [16-1:0] node12418;
	wire [16-1:0] node12419;
	wire [16-1:0] node12421;
	wire [16-1:0] node12424;
	wire [16-1:0] node12426;
	wire [16-1:0] node12429;
	wire [16-1:0] node12430;
	wire [16-1:0] node12432;
	wire [16-1:0] node12435;
	wire [16-1:0] node12437;
	wire [16-1:0] node12438;
	wire [16-1:0] node12442;
	wire [16-1:0] node12444;
	wire [16-1:0] node12446;
	wire [16-1:0] node12449;
	wire [16-1:0] node12450;
	wire [16-1:0] node12452;
	wire [16-1:0] node12453;
	wire [16-1:0] node12455;
	wire [16-1:0] node12458;
	wire [16-1:0] node12461;
	wire [16-1:0] node12462;
	wire [16-1:0] node12464;
	wire [16-1:0] node12468;
	wire [16-1:0] node12469;
	wire [16-1:0] node12470;
	wire [16-1:0] node12471;
	wire [16-1:0] node12472;
	wire [16-1:0] node12474;
	wire [16-1:0] node12477;
	wire [16-1:0] node12478;
	wire [16-1:0] node12479;
	wire [16-1:0] node12480;
	wire [16-1:0] node12485;
	wire [16-1:0] node12486;
	wire [16-1:0] node12489;
	wire [16-1:0] node12492;
	wire [16-1:0] node12493;
	wire [16-1:0] node12494;
	wire [16-1:0] node12496;
	wire [16-1:0] node12498;
	wire [16-1:0] node12501;
	wire [16-1:0] node12502;
	wire [16-1:0] node12504;
	wire [16-1:0] node12505;
	wire [16-1:0] node12510;
	wire [16-1:0] node12511;
	wire [16-1:0] node12512;
	wire [16-1:0] node12516;
	wire [16-1:0] node12517;
	wire [16-1:0] node12519;
	wire [16-1:0] node12523;
	wire [16-1:0] node12524;
	wire [16-1:0] node12525;
	wire [16-1:0] node12526;
	wire [16-1:0] node12527;
	wire [16-1:0] node12529;
	wire [16-1:0] node12532;
	wire [16-1:0] node12535;
	wire [16-1:0] node12536;
	wire [16-1:0] node12540;
	wire [16-1:0] node12541;
	wire [16-1:0] node12543;
	wire [16-1:0] node12545;
	wire [16-1:0] node12546;
	wire [16-1:0] node12550;
	wire [16-1:0] node12551;
	wire [16-1:0] node12552;
	wire [16-1:0] node12554;
	wire [16-1:0] node12558;
	wire [16-1:0] node12561;
	wire [16-1:0] node12562;
	wire [16-1:0] node12563;
	wire [16-1:0] node12564;
	wire [16-1:0] node12568;
	wire [16-1:0] node12570;
	wire [16-1:0] node12572;
	wire [16-1:0] node12575;
	wire [16-1:0] node12576;
	wire [16-1:0] node12578;
	wire [16-1:0] node12579;
	wire [16-1:0] node12583;
	wire [16-1:0] node12585;
	wire [16-1:0] node12586;
	wire [16-1:0] node12590;
	wire [16-1:0] node12591;
	wire [16-1:0] node12592;
	wire [16-1:0] node12593;
	wire [16-1:0] node12594;
	wire [16-1:0] node12595;
	wire [16-1:0] node12597;
	wire [16-1:0] node12601;
	wire [16-1:0] node12602;
	wire [16-1:0] node12604;
	wire [16-1:0] node12607;
	wire [16-1:0] node12610;
	wire [16-1:0] node12611;
	wire [16-1:0] node12612;
	wire [16-1:0] node12615;
	wire [16-1:0] node12618;
	wire [16-1:0] node12619;
	wire [16-1:0] node12620;
	wire [16-1:0] node12625;
	wire [16-1:0] node12626;
	wire [16-1:0] node12627;
	wire [16-1:0] node12629;
	wire [16-1:0] node12630;
	wire [16-1:0] node12634;
	wire [16-1:0] node12635;
	wire [16-1:0] node12638;
	wire [16-1:0] node12641;
	wire [16-1:0] node12642;
	wire [16-1:0] node12644;
	wire [16-1:0] node12647;
	wire [16-1:0] node12650;
	wire [16-1:0] node12651;
	wire [16-1:0] node12652;
	wire [16-1:0] node12653;
	wire [16-1:0] node12654;
	wire [16-1:0] node12657;
	wire [16-1:0] node12660;
	wire [16-1:0] node12661;
	wire [16-1:0] node12664;
	wire [16-1:0] node12667;
	wire [16-1:0] node12668;
	wire [16-1:0] node12670;
	wire [16-1:0] node12672;
	wire [16-1:0] node12673;
	wire [16-1:0] node12677;
	wire [16-1:0] node12678;
	wire [16-1:0] node12682;
	wire [16-1:0] node12683;
	wire [16-1:0] node12684;
	wire [16-1:0] node12686;
	wire [16-1:0] node12687;
	wire [16-1:0] node12689;
	wire [16-1:0] node12693;
	wire [16-1:0] node12695;
	wire [16-1:0] node12696;
	wire [16-1:0] node12698;
	wire [16-1:0] node12702;
	wire [16-1:0] node12703;
	wire [16-1:0] node12706;
	wire [16-1:0] node12709;
	wire [16-1:0] node12710;
	wire [16-1:0] node12711;
	wire [16-1:0] node12712;
	wire [16-1:0] node12713;
	wire [16-1:0] node12714;
	wire [16-1:0] node12715;
	wire [16-1:0] node12716;
	wire [16-1:0] node12717;
	wire [16-1:0] node12721;
	wire [16-1:0] node12722;
	wire [16-1:0] node12723;
	wire [16-1:0] node12724;
	wire [16-1:0] node12730;
	wire [16-1:0] node12731;
	wire [16-1:0] node12732;
	wire [16-1:0] node12734;
	wire [16-1:0] node12735;
	wire [16-1:0] node12739;
	wire [16-1:0] node12740;
	wire [16-1:0] node12742;
	wire [16-1:0] node12745;
	wire [16-1:0] node12748;
	wire [16-1:0] node12750;
	wire [16-1:0] node12753;
	wire [16-1:0] node12754;
	wire [16-1:0] node12756;
	wire [16-1:0] node12757;
	wire [16-1:0] node12760;
	wire [16-1:0] node12763;
	wire [16-1:0] node12765;
	wire [16-1:0] node12766;
	wire [16-1:0] node12770;
	wire [16-1:0] node12771;
	wire [16-1:0] node12772;
	wire [16-1:0] node12773;
	wire [16-1:0] node12774;
	wire [16-1:0] node12775;
	wire [16-1:0] node12779;
	wire [16-1:0] node12782;
	wire [16-1:0] node12783;
	wire [16-1:0] node12784;
	wire [16-1:0] node12789;
	wire [16-1:0] node12791;
	wire [16-1:0] node12792;
	wire [16-1:0] node12795;
	wire [16-1:0] node12798;
	wire [16-1:0] node12799;
	wire [16-1:0] node12802;
	wire [16-1:0] node12804;
	wire [16-1:0] node12805;
	wire [16-1:0] node12808;
	wire [16-1:0] node12810;
	wire [16-1:0] node12813;
	wire [16-1:0] node12814;
	wire [16-1:0] node12815;
	wire [16-1:0] node12816;
	wire [16-1:0] node12817;
	wire [16-1:0] node12820;
	wire [16-1:0] node12823;
	wire [16-1:0] node12825;
	wire [16-1:0] node12827;
	wire [16-1:0] node12830;
	wire [16-1:0] node12831;
	wire [16-1:0] node12832;
	wire [16-1:0] node12834;
	wire [16-1:0] node12835;
	wire [16-1:0] node12840;
	wire [16-1:0] node12841;
	wire [16-1:0] node12842;
	wire [16-1:0] node12843;
	wire [16-1:0] node12847;
	wire [16-1:0] node12850;
	wire [16-1:0] node12851;
	wire [16-1:0] node12854;
	wire [16-1:0] node12857;
	wire [16-1:0] node12858;
	wire [16-1:0] node12859;
	wire [16-1:0] node12860;
	wire [16-1:0] node12862;
	wire [16-1:0] node12865;
	wire [16-1:0] node12866;
	wire [16-1:0] node12870;
	wire [16-1:0] node12872;
	wire [16-1:0] node12873;
	wire [16-1:0] node12876;
	wire [16-1:0] node12879;
	wire [16-1:0] node12880;
	wire [16-1:0] node12881;
	wire [16-1:0] node12883;
	wire [16-1:0] node12885;
	wire [16-1:0] node12886;
	wire [16-1:0] node12891;
	wire [16-1:0] node12893;
	wire [16-1:0] node12894;
	wire [16-1:0] node12898;
	wire [16-1:0] node12899;
	wire [16-1:0] node12900;
	wire [16-1:0] node12901;
	wire [16-1:0] node12902;
	wire [16-1:0] node12903;
	wire [16-1:0] node12906;
	wire [16-1:0] node12909;
	wire [16-1:0] node12910;
	wire [16-1:0] node12911;
	wire [16-1:0] node12913;
	wire [16-1:0] node12917;
	wire [16-1:0] node12919;
	wire [16-1:0] node12922;
	wire [16-1:0] node12923;
	wire [16-1:0] node12924;
	wire [16-1:0] node12926;
	wire [16-1:0] node12929;
	wire [16-1:0] node12930;
	wire [16-1:0] node12934;
	wire [16-1:0] node12936;
	wire [16-1:0] node12937;
	wire [16-1:0] node12941;
	wire [16-1:0] node12942;
	wire [16-1:0] node12943;
	wire [16-1:0] node12944;
	wire [16-1:0] node12945;
	wire [16-1:0] node12948;
	wire [16-1:0] node12951;
	wire [16-1:0] node12952;
	wire [16-1:0] node12955;
	wire [16-1:0] node12956;
	wire [16-1:0] node12960;
	wire [16-1:0] node12961;
	wire [16-1:0] node12964;
	wire [16-1:0] node12965;
	wire [16-1:0] node12969;
	wire [16-1:0] node12970;
	wire [16-1:0] node12971;
	wire [16-1:0] node12973;
	wire [16-1:0] node12977;
	wire [16-1:0] node12978;
	wire [16-1:0] node12979;
	wire [16-1:0] node12982;
	wire [16-1:0] node12985;
	wire [16-1:0] node12986;
	wire [16-1:0] node12987;
	wire [16-1:0] node12992;
	wire [16-1:0] node12993;
	wire [16-1:0] node12994;
	wire [16-1:0] node12995;
	wire [16-1:0] node12996;
	wire [16-1:0] node12999;
	wire [16-1:0] node13000;
	wire [16-1:0] node13004;
	wire [16-1:0] node13005;
	wire [16-1:0] node13006;
	wire [16-1:0] node13009;
	wire [16-1:0] node13012;
	wire [16-1:0] node13013;
	wire [16-1:0] node13017;
	wire [16-1:0] node13018;
	wire [16-1:0] node13019;
	wire [16-1:0] node13020;
	wire [16-1:0] node13023;
	wire [16-1:0] node13026;
	wire [16-1:0] node13029;
	wire [16-1:0] node13030;
	wire [16-1:0] node13032;
	wire [16-1:0] node13033;
	wire [16-1:0] node13035;
	wire [16-1:0] node13039;
	wire [16-1:0] node13040;
	wire [16-1:0] node13041;
	wire [16-1:0] node13045;
	wire [16-1:0] node13046;
	wire [16-1:0] node13048;
	wire [16-1:0] node13052;
	wire [16-1:0] node13053;
	wire [16-1:0] node13054;
	wire [16-1:0] node13056;
	wire [16-1:0] node13060;
	wire [16-1:0] node13062;
	wire [16-1:0] node13063;
	wire [16-1:0] node13066;
	wire [16-1:0] node13068;
	wire [16-1:0] node13071;
	wire [16-1:0] node13072;
	wire [16-1:0] node13073;
	wire [16-1:0] node13074;
	wire [16-1:0] node13075;
	wire [16-1:0] node13076;
	wire [16-1:0] node13077;
	wire [16-1:0] node13078;
	wire [16-1:0] node13079;
	wire [16-1:0] node13081;
	wire [16-1:0] node13085;
	wire [16-1:0] node13089;
	wire [16-1:0] node13090;
	wire [16-1:0] node13091;
	wire [16-1:0] node13095;
	wire [16-1:0] node13096;
	wire [16-1:0] node13100;
	wire [16-1:0] node13101;
	wire [16-1:0] node13102;
	wire [16-1:0] node13103;
	wire [16-1:0] node13108;
	wire [16-1:0] node13109;
	wire [16-1:0] node13111;
	wire [16-1:0] node13113;
	wire [16-1:0] node13116;
	wire [16-1:0] node13117;
	wire [16-1:0] node13118;
	wire [16-1:0] node13122;
	wire [16-1:0] node13125;
	wire [16-1:0] node13126;
	wire [16-1:0] node13127;
	wire [16-1:0] node13129;
	wire [16-1:0] node13131;
	wire [16-1:0] node13134;
	wire [16-1:0] node13136;
	wire [16-1:0] node13137;
	wire [16-1:0] node13138;
	wire [16-1:0] node13143;
	wire [16-1:0] node13144;
	wire [16-1:0] node13146;
	wire [16-1:0] node13149;
	wire [16-1:0] node13150;
	wire [16-1:0] node13151;
	wire [16-1:0] node13152;
	wire [16-1:0] node13157;
	wire [16-1:0] node13158;
	wire [16-1:0] node13162;
	wire [16-1:0] node13163;
	wire [16-1:0] node13164;
	wire [16-1:0] node13165;
	wire [16-1:0] node13166;
	wire [16-1:0] node13168;
	wire [16-1:0] node13169;
	wire [16-1:0] node13174;
	wire [16-1:0] node13175;
	wire [16-1:0] node13176;
	wire [16-1:0] node13180;
	wire [16-1:0] node13182;
	wire [16-1:0] node13185;
	wire [16-1:0] node13186;
	wire [16-1:0] node13187;
	wire [16-1:0] node13189;
	wire [16-1:0] node13191;
	wire [16-1:0] node13194;
	wire [16-1:0] node13195;
	wire [16-1:0] node13198;
	wire [16-1:0] node13200;
	wire [16-1:0] node13203;
	wire [16-1:0] node13204;
	wire [16-1:0] node13205;
	wire [16-1:0] node13209;
	wire [16-1:0] node13211;
	wire [16-1:0] node13213;
	wire [16-1:0] node13216;
	wire [16-1:0] node13217;
	wire [16-1:0] node13218;
	wire [16-1:0] node13219;
	wire [16-1:0] node13222;
	wire [16-1:0] node13224;
	wire [16-1:0] node13227;
	wire [16-1:0] node13228;
	wire [16-1:0] node13230;
	wire [16-1:0] node13233;
	wire [16-1:0] node13235;
	wire [16-1:0] node13238;
	wire [16-1:0] node13239;
	wire [16-1:0] node13240;
	wire [16-1:0] node13241;
	wire [16-1:0] node13246;
	wire [16-1:0] node13247;
	wire [16-1:0] node13248;
	wire [16-1:0] node13249;
	wire [16-1:0] node13253;
	wire [16-1:0] node13256;
	wire [16-1:0] node13258;
	wire [16-1:0] node13261;
	wire [16-1:0] node13262;
	wire [16-1:0] node13263;
	wire [16-1:0] node13264;
	wire [16-1:0] node13265;
	wire [16-1:0] node13268;
	wire [16-1:0] node13270;
	wire [16-1:0] node13271;
	wire [16-1:0] node13272;
	wire [16-1:0] node13273;
	wire [16-1:0] node13279;
	wire [16-1:0] node13280;
	wire [16-1:0] node13282;
	wire [16-1:0] node13284;
	wire [16-1:0] node13287;
	wire [16-1:0] node13288;
	wire [16-1:0] node13289;
	wire [16-1:0] node13290;
	wire [16-1:0] node13295;
	wire [16-1:0] node13298;
	wire [16-1:0] node13299;
	wire [16-1:0] node13300;
	wire [16-1:0] node13301;
	wire [16-1:0] node13302;
	wire [16-1:0] node13305;
	wire [16-1:0] node13306;
	wire [16-1:0] node13310;
	wire [16-1:0] node13311;
	wire [16-1:0] node13312;
	wire [16-1:0] node13316;
	wire [16-1:0] node13319;
	wire [16-1:0] node13321;
	wire [16-1:0] node13322;
	wire [16-1:0] node13325;
	wire [16-1:0] node13328;
	wire [16-1:0] node13329;
	wire [16-1:0] node13330;
	wire [16-1:0] node13331;
	wire [16-1:0] node13334;
	wire [16-1:0] node13336;
	wire [16-1:0] node13337;
	wire [16-1:0] node13342;
	wire [16-1:0] node13343;
	wire [16-1:0] node13344;
	wire [16-1:0] node13348;
	wire [16-1:0] node13349;
	wire [16-1:0] node13352;
	wire [16-1:0] node13354;
	wire [16-1:0] node13357;
	wire [16-1:0] node13358;
	wire [16-1:0] node13359;
	wire [16-1:0] node13360;
	wire [16-1:0] node13361;
	wire [16-1:0] node13362;
	wire [16-1:0] node13364;
	wire [16-1:0] node13365;
	wire [16-1:0] node13371;
	wire [16-1:0] node13372;
	wire [16-1:0] node13373;
	wire [16-1:0] node13377;
	wire [16-1:0] node13379;
	wire [16-1:0] node13382;
	wire [16-1:0] node13383;
	wire [16-1:0] node13384;
	wire [16-1:0] node13386;
	wire [16-1:0] node13389;
	wire [16-1:0] node13390;
	wire [16-1:0] node13394;
	wire [16-1:0] node13395;
	wire [16-1:0] node13397;
	wire [16-1:0] node13399;
	wire [16-1:0] node13402;
	wire [16-1:0] node13403;
	wire [16-1:0] node13407;
	wire [16-1:0] node13408;
	wire [16-1:0] node13409;
	wire [16-1:0] node13410;
	wire [16-1:0] node13413;
	wire [16-1:0] node13415;
	wire [16-1:0] node13416;
	wire [16-1:0] node13417;
	wire [16-1:0] node13422;
	wire [16-1:0] node13423;
	wire [16-1:0] node13425;
	wire [16-1:0] node13426;
	wire [16-1:0] node13428;
	wire [16-1:0] node13432;
	wire [16-1:0] node13433;
	wire [16-1:0] node13436;
	wire [16-1:0] node13439;
	wire [16-1:0] node13440;
	wire [16-1:0] node13441;
	wire [16-1:0] node13443;
	wire [16-1:0] node13447;
	wire [16-1:0] node13448;
	wire [16-1:0] node13450;
	wire [16-1:0] node13451;
	wire [16-1:0] node13453;
	wire [16-1:0] node13456;
	wire [16-1:0] node13458;
	wire [16-1:0] node13461;
	wire [16-1:0] node13464;
	wire [16-1:0] node13465;
	wire [16-1:0] node13466;
	wire [16-1:0] node13467;
	wire [16-1:0] node13468;
	wire [16-1:0] node13469;
	wire [16-1:0] node13470;
	wire [16-1:0] node13471;
	wire [16-1:0] node13472;
	wire [16-1:0] node13473;
	wire [16-1:0] node13474;
	wire [16-1:0] node13478;
	wire [16-1:0] node13479;
	wire [16-1:0] node13483;
	wire [16-1:0] node13484;
	wire [16-1:0] node13485;
	wire [16-1:0] node13490;
	wire [16-1:0] node13491;
	wire [16-1:0] node13492;
	wire [16-1:0] node13495;
	wire [16-1:0] node13497;
	wire [16-1:0] node13500;
	wire [16-1:0] node13501;
	wire [16-1:0] node13502;
	wire [16-1:0] node13506;
	wire [16-1:0] node13509;
	wire [16-1:0] node13510;
	wire [16-1:0] node13511;
	wire [16-1:0] node13512;
	wire [16-1:0] node13515;
	wire [16-1:0] node13518;
	wire [16-1:0] node13521;
	wire [16-1:0] node13522;
	wire [16-1:0] node13524;
	wire [16-1:0] node13525;
	wire [16-1:0] node13530;
	wire [16-1:0] node13531;
	wire [16-1:0] node13532;
	wire [16-1:0] node13533;
	wire [16-1:0] node13535;
	wire [16-1:0] node13537;
	wire [16-1:0] node13540;
	wire [16-1:0] node13541;
	wire [16-1:0] node13545;
	wire [16-1:0] node13546;
	wire [16-1:0] node13547;
	wire [16-1:0] node13550;
	wire [16-1:0] node13552;
	wire [16-1:0] node13554;
	wire [16-1:0] node13558;
	wire [16-1:0] node13559;
	wire [16-1:0] node13560;
	wire [16-1:0] node13561;
	wire [16-1:0] node13566;
	wire [16-1:0] node13567;
	wire [16-1:0] node13568;
	wire [16-1:0] node13571;
	wire [16-1:0] node13573;
	wire [16-1:0] node13576;
	wire [16-1:0] node13577;
	wire [16-1:0] node13580;
	wire [16-1:0] node13583;
	wire [16-1:0] node13584;
	wire [16-1:0] node13585;
	wire [16-1:0] node13586;
	wire [16-1:0] node13587;
	wire [16-1:0] node13588;
	wire [16-1:0] node13589;
	wire [16-1:0] node13594;
	wire [16-1:0] node13597;
	wire [16-1:0] node13600;
	wire [16-1:0] node13601;
	wire [16-1:0] node13603;
	wire [16-1:0] node13604;
	wire [16-1:0] node13608;
	wire [16-1:0] node13609;
	wire [16-1:0] node13612;
	wire [16-1:0] node13615;
	wire [16-1:0] node13616;
	wire [16-1:0] node13617;
	wire [16-1:0] node13618;
	wire [16-1:0] node13620;
	wire [16-1:0] node13622;
	wire [16-1:0] node13624;
	wire [16-1:0] node13628;
	wire [16-1:0] node13629;
	wire [16-1:0] node13630;
	wire [16-1:0] node13631;
	wire [16-1:0] node13635;
	wire [16-1:0] node13638;
	wire [16-1:0] node13639;
	wire [16-1:0] node13643;
	wire [16-1:0] node13644;
	wire [16-1:0] node13645;
	wire [16-1:0] node13649;
	wire [16-1:0] node13650;
	wire [16-1:0] node13652;
	wire [16-1:0] node13655;
	wire [16-1:0] node13657;
	wire [16-1:0] node13660;
	wire [16-1:0] node13661;
	wire [16-1:0] node13662;
	wire [16-1:0] node13663;
	wire [16-1:0] node13664;
	wire [16-1:0] node13665;
	wire [16-1:0] node13666;
	wire [16-1:0] node13669;
	wire [16-1:0] node13671;
	wire [16-1:0] node13674;
	wire [16-1:0] node13675;
	wire [16-1:0] node13679;
	wire [16-1:0] node13680;
	wire [16-1:0] node13683;
	wire [16-1:0] node13686;
	wire [16-1:0] node13687;
	wire [16-1:0] node13688;
	wire [16-1:0] node13689;
	wire [16-1:0] node13692;
	wire [16-1:0] node13695;
	wire [16-1:0] node13696;
	wire [16-1:0] node13699;
	wire [16-1:0] node13702;
	wire [16-1:0] node13704;
	wire [16-1:0] node13705;
	wire [16-1:0] node13709;
	wire [16-1:0] node13710;
	wire [16-1:0] node13711;
	wire [16-1:0] node13712;
	wire [16-1:0] node13713;
	wire [16-1:0] node13717;
	wire [16-1:0] node13718;
	wire [16-1:0] node13720;
	wire [16-1:0] node13721;
	wire [16-1:0] node13725;
	wire [16-1:0] node13728;
	wire [16-1:0] node13729;
	wire [16-1:0] node13731;
	wire [16-1:0] node13733;
	wire [16-1:0] node13736;
	wire [16-1:0] node13738;
	wire [16-1:0] node13741;
	wire [16-1:0] node13742;
	wire [16-1:0] node13743;
	wire [16-1:0] node13744;
	wire [16-1:0] node13747;
	wire [16-1:0] node13751;
	wire [16-1:0] node13753;
	wire [16-1:0] node13754;
	wire [16-1:0] node13757;
	wire [16-1:0] node13759;
	wire [16-1:0] node13762;
	wire [16-1:0] node13763;
	wire [16-1:0] node13764;
	wire [16-1:0] node13765;
	wire [16-1:0] node13766;
	wire [16-1:0] node13768;
	wire [16-1:0] node13769;
	wire [16-1:0] node13772;
	wire [16-1:0] node13776;
	wire [16-1:0] node13777;
	wire [16-1:0] node13779;
	wire [16-1:0] node13782;
	wire [16-1:0] node13783;
	wire [16-1:0] node13787;
	wire [16-1:0] node13788;
	wire [16-1:0] node13789;
	wire [16-1:0] node13790;
	wire [16-1:0] node13794;
	wire [16-1:0] node13795;
	wire [16-1:0] node13798;
	wire [16-1:0] node13801;
	wire [16-1:0] node13803;
	wire [16-1:0] node13805;
	wire [16-1:0] node13808;
	wire [16-1:0] node13809;
	wire [16-1:0] node13810;
	wire [16-1:0] node13811;
	wire [16-1:0] node13813;
	wire [16-1:0] node13816;
	wire [16-1:0] node13817;
	wire [16-1:0] node13821;
	wire [16-1:0] node13822;
	wire [16-1:0] node13823;
	wire [16-1:0] node13826;
	wire [16-1:0] node13828;
	wire [16-1:0] node13829;
	wire [16-1:0] node13833;
	wire [16-1:0] node13834;
	wire [16-1:0] node13838;
	wire [16-1:0] node13839;
	wire [16-1:0] node13840;
	wire [16-1:0] node13842;
	wire [16-1:0] node13845;
	wire [16-1:0] node13846;
	wire [16-1:0] node13849;
	wire [16-1:0] node13852;
	wire [16-1:0] node13853;
	wire [16-1:0] node13854;
	wire [16-1:0] node13856;
	wire [16-1:0] node13860;
	wire [16-1:0] node13862;
	wire [16-1:0] node13864;
	wire [16-1:0] node13867;
	wire [16-1:0] node13868;
	wire [16-1:0] node13869;
	wire [16-1:0] node13870;
	wire [16-1:0] node13871;
	wire [16-1:0] node13872;
	wire [16-1:0] node13873;
	wire [16-1:0] node13874;
	wire [16-1:0] node13875;
	wire [16-1:0] node13878;
	wire [16-1:0] node13882;
	wire [16-1:0] node13883;
	wire [16-1:0] node13885;
	wire [16-1:0] node13886;
	wire [16-1:0] node13890;
	wire [16-1:0] node13893;
	wire [16-1:0] node13894;
	wire [16-1:0] node13895;
	wire [16-1:0] node13899;
	wire [16-1:0] node13900;
	wire [16-1:0] node13903;
	wire [16-1:0] node13906;
	wire [16-1:0] node13907;
	wire [16-1:0] node13908;
	wire [16-1:0] node13909;
	wire [16-1:0] node13912;
	wire [16-1:0] node13915;
	wire [16-1:0] node13918;
	wire [16-1:0] node13919;
	wire [16-1:0] node13922;
	wire [16-1:0] node13923;
	wire [16-1:0] node13925;
	wire [16-1:0] node13929;
	wire [16-1:0] node13930;
	wire [16-1:0] node13931;
	wire [16-1:0] node13933;
	wire [16-1:0] node13934;
	wire [16-1:0] node13937;
	wire [16-1:0] node13940;
	wire [16-1:0] node13942;
	wire [16-1:0] node13943;
	wire [16-1:0] node13947;
	wire [16-1:0] node13948;
	wire [16-1:0] node13949;
	wire [16-1:0] node13951;
	wire [16-1:0] node13952;
	wire [16-1:0] node13953;
	wire [16-1:0] node13958;
	wire [16-1:0] node13959;
	wire [16-1:0] node13961;
	wire [16-1:0] node13963;
	wire [16-1:0] node13967;
	wire [16-1:0] node13968;
	wire [16-1:0] node13969;
	wire [16-1:0] node13971;
	wire [16-1:0] node13975;
	wire [16-1:0] node13977;
	wire [16-1:0] node13980;
	wire [16-1:0] node13981;
	wire [16-1:0] node13982;
	wire [16-1:0] node13983;
	wire [16-1:0] node13984;
	wire [16-1:0] node13985;
	wire [16-1:0] node13986;
	wire [16-1:0] node13991;
	wire [16-1:0] node13993;
	wire [16-1:0] node13996;
	wire [16-1:0] node13997;
	wire [16-1:0] node14000;
	wire [16-1:0] node14001;
	wire [16-1:0] node14005;
	wire [16-1:0] node14006;
	wire [16-1:0] node14009;
	wire [16-1:0] node14010;
	wire [16-1:0] node14011;
	wire [16-1:0] node14014;
	wire [16-1:0] node14015;
	wire [16-1:0] node14017;
	wire [16-1:0] node14021;
	wire [16-1:0] node14022;
	wire [16-1:0] node14025;
	wire [16-1:0] node14028;
	wire [16-1:0] node14029;
	wire [16-1:0] node14030;
	wire [16-1:0] node14031;
	wire [16-1:0] node14033;
	wire [16-1:0] node14034;
	wire [16-1:0] node14039;
	wire [16-1:0] node14041;
	wire [16-1:0] node14043;
	wire [16-1:0] node14046;
	wire [16-1:0] node14047;
	wire [16-1:0] node14048;
	wire [16-1:0] node14049;
	wire [16-1:0] node14054;
	wire [16-1:0] node14055;
	wire [16-1:0] node14056;
	wire [16-1:0] node14059;
	wire [16-1:0] node14062;
	wire [16-1:0] node14063;
	wire [16-1:0] node14067;
	wire [16-1:0] node14068;
	wire [16-1:0] node14069;
	wire [16-1:0] node14070;
	wire [16-1:0] node14071;
	wire [16-1:0] node14073;
	wire [16-1:0] node14076;
	wire [16-1:0] node14077;
	wire [16-1:0] node14081;
	wire [16-1:0] node14082;
	wire [16-1:0] node14083;
	wire [16-1:0] node14084;
	wire [16-1:0] node14085;
	wire [16-1:0] node14087;
	wire [16-1:0] node14091;
	wire [16-1:0] node14094;
	wire [16-1:0] node14096;
	wire [16-1:0] node14098;
	wire [16-1:0] node14100;
	wire [16-1:0] node14103;
	wire [16-1:0] node14104;
	wire [16-1:0] node14107;
	wire [16-1:0] node14108;
	wire [16-1:0] node14111;
	wire [16-1:0] node14113;
	wire [16-1:0] node14116;
	wire [16-1:0] node14117;
	wire [16-1:0] node14118;
	wire [16-1:0] node14121;
	wire [16-1:0] node14122;
	wire [16-1:0] node14123;
	wire [16-1:0] node14126;
	wire [16-1:0] node14128;
	wire [16-1:0] node14132;
	wire [16-1:0] node14133;
	wire [16-1:0] node14134;
	wire [16-1:0] node14135;
	wire [16-1:0] node14136;
	wire [16-1:0] node14141;
	wire [16-1:0] node14143;
	wire [16-1:0] node14144;
	wire [16-1:0] node14148;
	wire [16-1:0] node14149;
	wire [16-1:0] node14151;
	wire [16-1:0] node14155;
	wire [16-1:0] node14156;
	wire [16-1:0] node14157;
	wire [16-1:0] node14158;
	wire [16-1:0] node14159;
	wire [16-1:0] node14162;
	wire [16-1:0] node14163;
	wire [16-1:0] node14164;
	wire [16-1:0] node14169;
	wire [16-1:0] node14170;
	wire [16-1:0] node14172;
	wire [16-1:0] node14175;
	wire [16-1:0] node14177;
	wire [16-1:0] node14178;
	wire [16-1:0] node14182;
	wire [16-1:0] node14183;
	wire [16-1:0] node14184;
	wire [16-1:0] node14186;
	wire [16-1:0] node14189;
	wire [16-1:0] node14190;
	wire [16-1:0] node14191;
	wire [16-1:0] node14195;
	wire [16-1:0] node14196;
	wire [16-1:0] node14200;
	wire [16-1:0] node14201;
	wire [16-1:0] node14203;
	wire [16-1:0] node14204;
	wire [16-1:0] node14208;
	wire [16-1:0] node14210;
	wire [16-1:0] node14213;
	wire [16-1:0] node14214;
	wire [16-1:0] node14215;
	wire [16-1:0] node14216;
	wire [16-1:0] node14220;
	wire [16-1:0] node14222;
	wire [16-1:0] node14223;
	wire [16-1:0] node14224;
	wire [16-1:0] node14228;
	wire [16-1:0] node14230;
	wire [16-1:0] node14233;
	wire [16-1:0] node14234;
	wire [16-1:0] node14235;
	wire [16-1:0] node14236;
	wire [16-1:0] node14239;
	wire [16-1:0] node14242;
	wire [16-1:0] node14243;
	wire [16-1:0] node14246;
	wire [16-1:0] node14249;
	wire [16-1:0] node14250;
	wire [16-1:0] node14252;
	wire [16-1:0] node14255;
	wire [16-1:0] node14256;
	wire [16-1:0] node14259;
	wire [16-1:0] node14262;
	wire [16-1:0] node14263;
	wire [16-1:0] node14264;
	wire [16-1:0] node14265;
	wire [16-1:0] node14266;
	wire [16-1:0] node14267;
	wire [16-1:0] node14268;
	wire [16-1:0] node14269;
	wire [16-1:0] node14270;
	wire [16-1:0] node14271;
	wire [16-1:0] node14272;
	wire [16-1:0] node14277;
	wire [16-1:0] node14281;
	wire [16-1:0] node14282;
	wire [16-1:0] node14283;
	wire [16-1:0] node14287;
	wire [16-1:0] node14288;
	wire [16-1:0] node14292;
	wire [16-1:0] node14293;
	wire [16-1:0] node14294;
	wire [16-1:0] node14295;
	wire [16-1:0] node14296;
	wire [16-1:0] node14300;
	wire [16-1:0] node14302;
	wire [16-1:0] node14303;
	wire [16-1:0] node14307;
	wire [16-1:0] node14310;
	wire [16-1:0] node14311;
	wire [16-1:0] node14312;
	wire [16-1:0] node14315;
	wire [16-1:0] node14318;
	wire [16-1:0] node14319;
	wire [16-1:0] node14320;
	wire [16-1:0] node14325;
	wire [16-1:0] node14326;
	wire [16-1:0] node14327;
	wire [16-1:0] node14328;
	wire [16-1:0] node14329;
	wire [16-1:0] node14334;
	wire [16-1:0] node14335;
	wire [16-1:0] node14338;
	wire [16-1:0] node14340;
	wire [16-1:0] node14343;
	wire [16-1:0] node14344;
	wire [16-1:0] node14345;
	wire [16-1:0] node14346;
	wire [16-1:0] node14349;
	wire [16-1:0] node14350;
	wire [16-1:0] node14352;
	wire [16-1:0] node14356;
	wire [16-1:0] node14359;
	wire [16-1:0] node14360;
	wire [16-1:0] node14361;
	wire [16-1:0] node14364;
	wire [16-1:0] node14367;
	wire [16-1:0] node14368;
	wire [16-1:0] node14372;
	wire [16-1:0] node14373;
	wire [16-1:0] node14374;
	wire [16-1:0] node14375;
	wire [16-1:0] node14376;
	wire [16-1:0] node14377;
	wire [16-1:0] node14381;
	wire [16-1:0] node14384;
	wire [16-1:0] node14386;
	wire [16-1:0] node14387;
	wire [16-1:0] node14388;
	wire [16-1:0] node14393;
	wire [16-1:0] node14394;
	wire [16-1:0] node14395;
	wire [16-1:0] node14396;
	wire [16-1:0] node14397;
	wire [16-1:0] node14403;
	wire [16-1:0] node14405;
	wire [16-1:0] node14407;
	wire [16-1:0] node14409;
	wire [16-1:0] node14412;
	wire [16-1:0] node14413;
	wire [16-1:0] node14414;
	wire [16-1:0] node14415;
	wire [16-1:0] node14419;
	wire [16-1:0] node14420;
	wire [16-1:0] node14421;
	wire [16-1:0] node14422;
	wire [16-1:0] node14424;
	wire [16-1:0] node14428;
	wire [16-1:0] node14431;
	wire [16-1:0] node14432;
	wire [16-1:0] node14436;
	wire [16-1:0] node14437;
	wire [16-1:0] node14438;
	wire [16-1:0] node14440;
	wire [16-1:0] node14443;
	wire [16-1:0] node14446;
	wire [16-1:0] node14447;
	wire [16-1:0] node14448;
	wire [16-1:0] node14451;
	wire [16-1:0] node14452;
	wire [16-1:0] node14456;
	wire [16-1:0] node14457;
	wire [16-1:0] node14460;
	wire [16-1:0] node14462;
	wire [16-1:0] node14465;
	wire [16-1:0] node14466;
	wire [16-1:0] node14467;
	wire [16-1:0] node14468;
	wire [16-1:0] node14469;
	wire [16-1:0] node14470;
	wire [16-1:0] node14473;
	wire [16-1:0] node14476;
	wire [16-1:0] node14477;
	wire [16-1:0] node14479;
	wire [16-1:0] node14482;
	wire [16-1:0] node14483;
	wire [16-1:0] node14487;
	wire [16-1:0] node14488;
	wire [16-1:0] node14489;
	wire [16-1:0] node14490;
	wire [16-1:0] node14491;
	wire [16-1:0] node14493;
	wire [16-1:0] node14498;
	wire [16-1:0] node14499;
	wire [16-1:0] node14503;
	wire [16-1:0] node14505;
	wire [16-1:0] node14506;
	wire [16-1:0] node14509;
	wire [16-1:0] node14510;
	wire [16-1:0] node14514;
	wire [16-1:0] node14515;
	wire [16-1:0] node14516;
	wire [16-1:0] node14517;
	wire [16-1:0] node14518;
	wire [16-1:0] node14522;
	wire [16-1:0] node14523;
	wire [16-1:0] node14527;
	wire [16-1:0] node14528;
	wire [16-1:0] node14530;
	wire [16-1:0] node14533;
	wire [16-1:0] node14536;
	wire [16-1:0] node14537;
	wire [16-1:0] node14538;
	wire [16-1:0] node14539;
	wire [16-1:0] node14540;
	wire [16-1:0] node14545;
	wire [16-1:0] node14547;
	wire [16-1:0] node14550;
	wire [16-1:0] node14551;
	wire [16-1:0] node14555;
	wire [16-1:0] node14556;
	wire [16-1:0] node14557;
	wire [16-1:0] node14558;
	wire [16-1:0] node14559;
	wire [16-1:0] node14560;
	wire [16-1:0] node14563;
	wire [16-1:0] node14565;
	wire [16-1:0] node14566;
	wire [16-1:0] node14570;
	wire [16-1:0] node14572;
	wire [16-1:0] node14573;
	wire [16-1:0] node14577;
	wire [16-1:0] node14579;
	wire [16-1:0] node14580;
	wire [16-1:0] node14581;
	wire [16-1:0] node14583;
	wire [16-1:0] node14588;
	wire [16-1:0] node14589;
	wire [16-1:0] node14590;
	wire [16-1:0] node14593;
	wire [16-1:0] node14596;
	wire [16-1:0] node14598;
	wire [16-1:0] node14599;
	wire [16-1:0] node14601;
	wire [16-1:0] node14602;
	wire [16-1:0] node14606;
	wire [16-1:0] node14609;
	wire [16-1:0] node14610;
	wire [16-1:0] node14611;
	wire [16-1:0] node14614;
	wire [16-1:0] node14615;
	wire [16-1:0] node14616;
	wire [16-1:0] node14618;
	wire [16-1:0] node14621;
	wire [16-1:0] node14622;
	wire [16-1:0] node14626;
	wire [16-1:0] node14627;
	wire [16-1:0] node14631;
	wire [16-1:0] node14632;
	wire [16-1:0] node14633;
	wire [16-1:0] node14635;
	wire [16-1:0] node14638;
	wire [16-1:0] node14641;
	wire [16-1:0] node14642;
	wire [16-1:0] node14645;
	wire [16-1:0] node14648;
	wire [16-1:0] node14649;
	wire [16-1:0] node14650;
	wire [16-1:0] node14651;
	wire [16-1:0] node14652;
	wire [16-1:0] node14653;
	wire [16-1:0] node14654;
	wire [16-1:0] node14655;
	wire [16-1:0] node14660;
	wire [16-1:0] node14663;
	wire [16-1:0] node14664;
	wire [16-1:0] node14666;
	wire [16-1:0] node14667;
	wire [16-1:0] node14669;
	wire [16-1:0] node14673;
	wire [16-1:0] node14675;
	wire [16-1:0] node14676;
	wire [16-1:0] node14678;
	wire [16-1:0] node14682;
	wire [16-1:0] node14683;
	wire [16-1:0] node14684;
	wire [16-1:0] node14685;
	wire [16-1:0] node14686;
	wire [16-1:0] node14690;
	wire [16-1:0] node14691;
	wire [16-1:0] node14692;
	wire [16-1:0] node14694;
	wire [16-1:0] node14699;
	wire [16-1:0] node14700;
	wire [16-1:0] node14703;
	wire [16-1:0] node14706;
	wire [16-1:0] node14707;
	wire [16-1:0] node14708;
	wire [16-1:0] node14711;
	wire [16-1:0] node14712;
	wire [16-1:0] node14713;
	wire [16-1:0] node14715;
	wire [16-1:0] node14720;
	wire [16-1:0] node14721;
	wire [16-1:0] node14722;
	wire [16-1:0] node14724;
	wire [16-1:0] node14729;
	wire [16-1:0] node14730;
	wire [16-1:0] node14731;
	wire [16-1:0] node14732;
	wire [16-1:0] node14734;
	wire [16-1:0] node14737;
	wire [16-1:0] node14738;
	wire [16-1:0] node14739;
	wire [16-1:0] node14741;
	wire [16-1:0] node14742;
	wire [16-1:0] node14747;
	wire [16-1:0] node14748;
	wire [16-1:0] node14750;
	wire [16-1:0] node14753;
	wire [16-1:0] node14756;
	wire [16-1:0] node14757;
	wire [16-1:0] node14759;
	wire [16-1:0] node14760;
	wire [16-1:0] node14761;
	wire [16-1:0] node14766;
	wire [16-1:0] node14767;
	wire [16-1:0] node14769;
	wire [16-1:0] node14771;
	wire [16-1:0] node14774;
	wire [16-1:0] node14775;
	wire [16-1:0] node14779;
	wire [16-1:0] node14780;
	wire [16-1:0] node14781;
	wire [16-1:0] node14782;
	wire [16-1:0] node14785;
	wire [16-1:0] node14786;
	wire [16-1:0] node14790;
	wire [16-1:0] node14792;
	wire [16-1:0] node14795;
	wire [16-1:0] node14796;
	wire [16-1:0] node14797;
	wire [16-1:0] node14799;
	wire [16-1:0] node14800;
	wire [16-1:0] node14802;
	wire [16-1:0] node14807;
	wire [16-1:0] node14808;
	wire [16-1:0] node14811;
	wire [16-1:0] node14812;
	wire [16-1:0] node14814;
	wire [16-1:0] node14818;
	wire [16-1:0] node14819;
	wire [16-1:0] node14820;
	wire [16-1:0] node14821;
	wire [16-1:0] node14822;
	wire [16-1:0] node14824;
	wire [16-1:0] node14825;
	wire [16-1:0] node14827;
	wire [16-1:0] node14830;
	wire [16-1:0] node14833;
	wire [16-1:0] node14834;
	wire [16-1:0] node14836;
	wire [16-1:0] node14840;
	wire [16-1:0] node14841;
	wire [16-1:0] node14842;
	wire [16-1:0] node14843;
	wire [16-1:0] node14846;
	wire [16-1:0] node14849;
	wire [16-1:0] node14850;
	wire [16-1:0] node14851;
	wire [16-1:0] node14855;
	wire [16-1:0] node14858;
	wire [16-1:0] node14859;
	wire [16-1:0] node14862;
	wire [16-1:0] node14864;
	wire [16-1:0] node14866;
	wire [16-1:0] node14869;
	wire [16-1:0] node14870;
	wire [16-1:0] node14871;
	wire [16-1:0] node14872;
	wire [16-1:0] node14874;
	wire [16-1:0] node14876;
	wire [16-1:0] node14879;
	wire [16-1:0] node14880;
	wire [16-1:0] node14881;
	wire [16-1:0] node14885;
	wire [16-1:0] node14887;
	wire [16-1:0] node14888;
	wire [16-1:0] node14892;
	wire [16-1:0] node14893;
	wire [16-1:0] node14896;
	wire [16-1:0] node14897;
	wire [16-1:0] node14899;
	wire [16-1:0] node14903;
	wire [16-1:0] node14904;
	wire [16-1:0] node14906;
	wire [16-1:0] node14909;
	wire [16-1:0] node14910;
	wire [16-1:0] node14912;
	wire [16-1:0] node14915;
	wire [16-1:0] node14917;
	wire [16-1:0] node14920;
	wire [16-1:0] node14921;
	wire [16-1:0] node14922;
	wire [16-1:0] node14923;
	wire [16-1:0] node14924;
	wire [16-1:0] node14925;
	wire [16-1:0] node14928;
	wire [16-1:0] node14930;
	wire [16-1:0] node14931;
	wire [16-1:0] node14935;
	wire [16-1:0] node14936;
	wire [16-1:0] node14937;
	wire [16-1:0] node14941;
	wire [16-1:0] node14942;
	wire [16-1:0] node14947;
	wire [16-1:0] node14948;
	wire [16-1:0] node14949;
	wire [16-1:0] node14950;
	wire [16-1:0] node14952;
	wire [16-1:0] node14954;
	wire [16-1:0] node14959;
	wire [16-1:0] node14960;
	wire [16-1:0] node14963;
	wire [16-1:0] node14964;
	wire [16-1:0] node14966;
	wire [16-1:0] node14968;
	wire [16-1:0] node14971;
	wire [16-1:0] node14972;
	wire [16-1:0] node14975;
	wire [16-1:0] node14978;
	wire [16-1:0] node14979;
	wire [16-1:0] node14980;
	wire [16-1:0] node14981;
	wire [16-1:0] node14985;
	wire [16-1:0] node14986;
	wire [16-1:0] node14987;
	wire [16-1:0] node14990;
	wire [16-1:0] node14993;
	wire [16-1:0] node14994;
	wire [16-1:0] node14997;
	wire [16-1:0] node15000;
	wire [16-1:0] node15001;
	wire [16-1:0] node15002;
	wire [16-1:0] node15004;
	wire [16-1:0] node15005;
	wire [16-1:0] node15007;
	wire [16-1:0] node15012;
	wire [16-1:0] node15013;
	wire [16-1:0] node15014;
	wire [16-1:0] node15015;
	wire [16-1:0] node15019;
	wire [16-1:0] node15022;
	wire [16-1:0] node15024;
	wire [16-1:0] node15025;
	wire [16-1:0] node15027;
	wire [16-1:0] node15031;
	wire [16-1:0] node15032;
	wire [16-1:0] node15033;
	wire [16-1:0] node15034;
	wire [16-1:0] node15035;
	wire [16-1:0] node15036;
	wire [16-1:0] node15037;
	wire [16-1:0] node15038;
	wire [16-1:0] node15039;
	wire [16-1:0] node15040;
	wire [16-1:0] node15044;
	wire [16-1:0] node15045;
	wire [16-1:0] node15049;
	wire [16-1:0] node15050;
	wire [16-1:0] node15051;
	wire [16-1:0] node15053;
	wire [16-1:0] node15056;
	wire [16-1:0] node15058;
	wire [16-1:0] node15061;
	wire [16-1:0] node15062;
	wire [16-1:0] node15064;
	wire [16-1:0] node15067;
	wire [16-1:0] node15068;
	wire [16-1:0] node15069;
	wire [16-1:0] node15071;
	wire [16-1:0] node15076;
	wire [16-1:0] node15077;
	wire [16-1:0] node15078;
	wire [16-1:0] node15079;
	wire [16-1:0] node15082;
	wire [16-1:0] node15083;
	wire [16-1:0] node15087;
	wire [16-1:0] node15088;
	wire [16-1:0] node15089;
	wire [16-1:0] node15090;
	wire [16-1:0] node15094;
	wire [16-1:0] node15097;
	wire [16-1:0] node15098;
	wire [16-1:0] node15101;
	wire [16-1:0] node15104;
	wire [16-1:0] node15105;
	wire [16-1:0] node15106;
	wire [16-1:0] node15107;
	wire [16-1:0] node15110;
	wire [16-1:0] node15113;
	wire [16-1:0] node15114;
	wire [16-1:0] node15117;
	wire [16-1:0] node15119;
	wire [16-1:0] node15122;
	wire [16-1:0] node15124;
	wire [16-1:0] node15127;
	wire [16-1:0] node15128;
	wire [16-1:0] node15129;
	wire [16-1:0] node15130;
	wire [16-1:0] node15132;
	wire [16-1:0] node15133;
	wire [16-1:0] node15137;
	wire [16-1:0] node15139;
	wire [16-1:0] node15140;
	wire [16-1:0] node15142;
	wire [16-1:0] node15146;
	wire [16-1:0] node15147;
	wire [16-1:0] node15148;
	wire [16-1:0] node15149;
	wire [16-1:0] node15152;
	wire [16-1:0] node15155;
	wire [16-1:0] node15158;
	wire [16-1:0] node15159;
	wire [16-1:0] node15161;
	wire [16-1:0] node15164;
	wire [16-1:0] node15165;
	wire [16-1:0] node15169;
	wire [16-1:0] node15170;
	wire [16-1:0] node15171;
	wire [16-1:0] node15172;
	wire [16-1:0] node15175;
	wire [16-1:0] node15178;
	wire [16-1:0] node15180;
	wire [16-1:0] node15181;
	wire [16-1:0] node15184;
	wire [16-1:0] node15187;
	wire [16-1:0] node15188;
	wire [16-1:0] node15189;
	wire [16-1:0] node15192;
	wire [16-1:0] node15194;
	wire [16-1:0] node15197;
	wire [16-1:0] node15198;
	wire [16-1:0] node15200;
	wire [16-1:0] node15202;
	wire [16-1:0] node15206;
	wire [16-1:0] node15207;
	wire [16-1:0] node15208;
	wire [16-1:0] node15209;
	wire [16-1:0] node15210;
	wire [16-1:0] node15211;
	wire [16-1:0] node15212;
	wire [16-1:0] node15215;
	wire [16-1:0] node15218;
	wire [16-1:0] node15220;
	wire [16-1:0] node15223;
	wire [16-1:0] node15225;
	wire [16-1:0] node15226;
	wire [16-1:0] node15227;
	wire [16-1:0] node15232;
	wire [16-1:0] node15233;
	wire [16-1:0] node15234;
	wire [16-1:0] node15237;
	wire [16-1:0] node15238;
	wire [16-1:0] node15239;
	wire [16-1:0] node15241;
	wire [16-1:0] node15246;
	wire [16-1:0] node15247;
	wire [16-1:0] node15249;
	wire [16-1:0] node15253;
	wire [16-1:0] node15254;
	wire [16-1:0] node15255;
	wire [16-1:0] node15256;
	wire [16-1:0] node15260;
	wire [16-1:0] node15261;
	wire [16-1:0] node15262;
	wire [16-1:0] node15263;
	wire [16-1:0] node15267;
	wire [16-1:0] node15270;
	wire [16-1:0] node15272;
	wire [16-1:0] node15275;
	wire [16-1:0] node15276;
	wire [16-1:0] node15277;
	wire [16-1:0] node15280;
	wire [16-1:0] node15283;
	wire [16-1:0] node15285;
	wire [16-1:0] node15287;
	wire [16-1:0] node15289;
	wire [16-1:0] node15292;
	wire [16-1:0] node15293;
	wire [16-1:0] node15294;
	wire [16-1:0] node15295;
	wire [16-1:0] node15296;
	wire [16-1:0] node15299;
	wire [16-1:0] node15301;
	wire [16-1:0] node15304;
	wire [16-1:0] node15305;
	wire [16-1:0] node15307;
	wire [16-1:0] node15309;
	wire [16-1:0] node15310;
	wire [16-1:0] node15314;
	wire [16-1:0] node15317;
	wire [16-1:0] node15318;
	wire [16-1:0] node15319;
	wire [16-1:0] node15322;
	wire [16-1:0] node15323;
	wire [16-1:0] node15326;
	wire [16-1:0] node15328;
	wire [16-1:0] node15331;
	wire [16-1:0] node15332;
	wire [16-1:0] node15335;
	wire [16-1:0] node15336;
	wire [16-1:0] node15340;
	wire [16-1:0] node15341;
	wire [16-1:0] node15342;
	wire [16-1:0] node15343;
	wire [16-1:0] node15345;
	wire [16-1:0] node15348;
	wire [16-1:0] node15349;
	wire [16-1:0] node15352;
	wire [16-1:0] node15354;
	wire [16-1:0] node15357;
	wire [16-1:0] node15359;
	wire [16-1:0] node15360;
	wire [16-1:0] node15364;
	wire [16-1:0] node15365;
	wire [16-1:0] node15367;
	wire [16-1:0] node15368;
	wire [16-1:0] node15369;
	wire [16-1:0] node15373;
	wire [16-1:0] node15376;
	wire [16-1:0] node15378;
	wire [16-1:0] node15380;
	wire [16-1:0] node15383;
	wire [16-1:0] node15384;
	wire [16-1:0] node15385;
	wire [16-1:0] node15386;
	wire [16-1:0] node15387;
	wire [16-1:0] node15388;
	wire [16-1:0] node15389;
	wire [16-1:0] node15392;
	wire [16-1:0] node15393;
	wire [16-1:0] node15397;
	wire [16-1:0] node15398;
	wire [16-1:0] node15399;
	wire [16-1:0] node15403;
	wire [16-1:0] node15404;
	wire [16-1:0] node15406;
	wire [16-1:0] node15410;
	wire [16-1:0] node15411;
	wire [16-1:0] node15412;
	wire [16-1:0] node15413;
	wire [16-1:0] node15416;
	wire [16-1:0] node15420;
	wire [16-1:0] node15421;
	wire [16-1:0] node15422;
	wire [16-1:0] node15424;
	wire [16-1:0] node15428;
	wire [16-1:0] node15429;
	wire [16-1:0] node15432;
	wire [16-1:0] node15434;
	wire [16-1:0] node15437;
	wire [16-1:0] node15438;
	wire [16-1:0] node15439;
	wire [16-1:0] node15440;
	wire [16-1:0] node15442;
	wire [16-1:0] node15445;
	wire [16-1:0] node15448;
	wire [16-1:0] node15449;
	wire [16-1:0] node15450;
	wire [16-1:0] node15455;
	wire [16-1:0] node15456;
	wire [16-1:0] node15457;
	wire [16-1:0] node15458;
	wire [16-1:0] node15461;
	wire [16-1:0] node15463;
	wire [16-1:0] node15464;
	wire [16-1:0] node15468;
	wire [16-1:0] node15470;
	wire [16-1:0] node15473;
	wire [16-1:0] node15474;
	wire [16-1:0] node15475;
	wire [16-1:0] node15480;
	wire [16-1:0] node15481;
	wire [16-1:0] node15482;
	wire [16-1:0] node15483;
	wire [16-1:0] node15484;
	wire [16-1:0] node15487;
	wire [16-1:0] node15488;
	wire [16-1:0] node15492;
	wire [16-1:0] node15494;
	wire [16-1:0] node15495;
	wire [16-1:0] node15496;
	wire [16-1:0] node15498;
	wire [16-1:0] node15503;
	wire [16-1:0] node15504;
	wire [16-1:0] node15506;
	wire [16-1:0] node15507;
	wire [16-1:0] node15511;
	wire [16-1:0] node15512;
	wire [16-1:0] node15513;
	wire [16-1:0] node15515;
	wire [16-1:0] node15516;
	wire [16-1:0] node15521;
	wire [16-1:0] node15522;
	wire [16-1:0] node15523;
	wire [16-1:0] node15525;
	wire [16-1:0] node15529;
	wire [16-1:0] node15532;
	wire [16-1:0] node15533;
	wire [16-1:0] node15534;
	wire [16-1:0] node15536;
	wire [16-1:0] node15538;
	wire [16-1:0] node15540;
	wire [16-1:0] node15543;
	wire [16-1:0] node15544;
	wire [16-1:0] node15546;
	wire [16-1:0] node15548;
	wire [16-1:0] node15551;
	wire [16-1:0] node15553;
	wire [16-1:0] node15556;
	wire [16-1:0] node15557;
	wire [16-1:0] node15559;
	wire [16-1:0] node15561;
	wire [16-1:0] node15563;
	wire [16-1:0] node15567;
	wire [16-1:0] node15568;
	wire [16-1:0] node15569;
	wire [16-1:0] node15570;
	wire [16-1:0] node15571;
	wire [16-1:0] node15572;
	wire [16-1:0] node15575;
	wire [16-1:0] node15576;
	wire [16-1:0] node15580;
	wire [16-1:0] node15581;
	wire [16-1:0] node15582;
	wire [16-1:0] node15586;
	wire [16-1:0] node15587;
	wire [16-1:0] node15591;
	wire [16-1:0] node15592;
	wire [16-1:0] node15593;
	wire [16-1:0] node15594;
	wire [16-1:0] node15598;
	wire [16-1:0] node15599;
	wire [16-1:0] node15603;
	wire [16-1:0] node15605;
	wire [16-1:0] node15606;
	wire [16-1:0] node15610;
	wire [16-1:0] node15611;
	wire [16-1:0] node15612;
	wire [16-1:0] node15613;
	wire [16-1:0] node15615;
	wire [16-1:0] node15616;
	wire [16-1:0] node15621;
	wire [16-1:0] node15622;
	wire [16-1:0] node15625;
	wire [16-1:0] node15628;
	wire [16-1:0] node15629;
	wire [16-1:0] node15630;
	wire [16-1:0] node15632;
	wire [16-1:0] node15635;
	wire [16-1:0] node15638;
	wire [16-1:0] node15639;
	wire [16-1:0] node15641;
	wire [16-1:0] node15644;
	wire [16-1:0] node15646;
	wire [16-1:0] node15649;
	wire [16-1:0] node15650;
	wire [16-1:0] node15651;
	wire [16-1:0] node15652;
	wire [16-1:0] node15653;
	wire [16-1:0] node15654;
	wire [16-1:0] node15657;
	wire [16-1:0] node15660;
	wire [16-1:0] node15661;
	wire [16-1:0] node15664;
	wire [16-1:0] node15665;
	wire [16-1:0] node15669;
	wire [16-1:0] node15670;
	wire [16-1:0] node15671;
	wire [16-1:0] node15674;
	wire [16-1:0] node15676;
	wire [16-1:0] node15679;
	wire [16-1:0] node15681;
	wire [16-1:0] node15684;
	wire [16-1:0] node15685;
	wire [16-1:0] node15686;
	wire [16-1:0] node15687;
	wire [16-1:0] node15689;
	wire [16-1:0] node15693;
	wire [16-1:0] node15695;
	wire [16-1:0] node15698;
	wire [16-1:0] node15699;
	wire [16-1:0] node15700;
	wire [16-1:0] node15704;
	wire [16-1:0] node15705;
	wire [16-1:0] node15709;
	wire [16-1:0] node15710;
	wire [16-1:0] node15711;
	wire [16-1:0] node15714;
	wire [16-1:0] node15715;
	wire [16-1:0] node15719;
	wire [16-1:0] node15720;
	wire [16-1:0] node15721;
	wire [16-1:0] node15724;
	wire [16-1:0] node15725;
	wire [16-1:0] node15727;
	wire [16-1:0] node15730;
	wire [16-1:0] node15731;
	wire [16-1:0] node15733;
	wire [16-1:0] node15737;
	wire [16-1:0] node15738;
	wire [16-1:0] node15740;
	wire [16-1:0] node15743;
	wire [16-1:0] node15746;
	wire [16-1:0] node15747;
	wire [16-1:0] node15748;
	wire [16-1:0] node15749;
	wire [16-1:0] node15750;
	wire [16-1:0] node15751;
	wire [16-1:0] node15752;
	wire [16-1:0] node15754;
	wire [16-1:0] node15755;
	wire [16-1:0] node15759;
	wire [16-1:0] node15760;
	wire [16-1:0] node15762;
	wire [16-1:0] node15766;
	wire [16-1:0] node15767;
	wire [16-1:0] node15768;
	wire [16-1:0] node15771;
	wire [16-1:0] node15772;
	wire [16-1:0] node15774;
	wire [16-1:0] node15777;
	wire [16-1:0] node15779;
	wire [16-1:0] node15780;
	wire [16-1:0] node15784;
	wire [16-1:0] node15785;
	wire [16-1:0] node15788;
	wire [16-1:0] node15791;
	wire [16-1:0] node15792;
	wire [16-1:0] node15793;
	wire [16-1:0] node15794;
	wire [16-1:0] node15795;
	wire [16-1:0] node15798;
	wire [16-1:0] node15799;
	wire [16-1:0] node15801;
	wire [16-1:0] node15805;
	wire [16-1:0] node15806;
	wire [16-1:0] node15809;
	wire [16-1:0] node15812;
	wire [16-1:0] node15814;
	wire [16-1:0] node15815;
	wire [16-1:0] node15817;
	wire [16-1:0] node15820;
	wire [16-1:0] node15823;
	wire [16-1:0] node15824;
	wire [16-1:0] node15825;
	wire [16-1:0] node15827;
	wire [16-1:0] node15828;
	wire [16-1:0] node15832;
	wire [16-1:0] node15834;
	wire [16-1:0] node15837;
	wire [16-1:0] node15838;
	wire [16-1:0] node15840;
	wire [16-1:0] node15843;
	wire [16-1:0] node15845;
	wire [16-1:0] node15848;
	wire [16-1:0] node15849;
	wire [16-1:0] node15850;
	wire [16-1:0] node15851;
	wire [16-1:0] node15853;
	wire [16-1:0] node15856;
	wire [16-1:0] node15857;
	wire [16-1:0] node15858;
	wire [16-1:0] node15861;
	wire [16-1:0] node15865;
	wire [16-1:0] node15866;
	wire [16-1:0] node15867;
	wire [16-1:0] node15868;
	wire [16-1:0] node15871;
	wire [16-1:0] node15875;
	wire [16-1:0] node15876;
	wire [16-1:0] node15877;
	wire [16-1:0] node15882;
	wire [16-1:0] node15883;
	wire [16-1:0] node15884;
	wire [16-1:0] node15885;
	wire [16-1:0] node15887;
	wire [16-1:0] node15890;
	wire [16-1:0] node15892;
	wire [16-1:0] node15895;
	wire [16-1:0] node15896;
	wire [16-1:0] node15897;
	wire [16-1:0] node15898;
	wire [16-1:0] node15902;
	wire [16-1:0] node15905;
	wire [16-1:0] node15907;
	wire [16-1:0] node15910;
	wire [16-1:0] node15911;
	wire [16-1:0] node15912;
	wire [16-1:0] node15913;
	wire [16-1:0] node15917;
	wire [16-1:0] node15920;
	wire [16-1:0] node15921;
	wire [16-1:0] node15924;
	wire [16-1:0] node15927;
	wire [16-1:0] node15928;
	wire [16-1:0] node15929;
	wire [16-1:0] node15930;
	wire [16-1:0] node15931;
	wire [16-1:0] node15932;
	wire [16-1:0] node15934;
	wire [16-1:0] node15936;
	wire [16-1:0] node15939;
	wire [16-1:0] node15940;
	wire [16-1:0] node15941;
	wire [16-1:0] node15943;
	wire [16-1:0] node15948;
	wire [16-1:0] node15951;
	wire [16-1:0] node15952;
	wire [16-1:0] node15953;
	wire [16-1:0] node15954;
	wire [16-1:0] node15958;
	wire [16-1:0] node15959;
	wire [16-1:0] node15961;
	wire [16-1:0] node15962;
	wire [16-1:0] node15966;
	wire [16-1:0] node15969;
	wire [16-1:0] node15970;
	wire [16-1:0] node15973;
	wire [16-1:0] node15975;
	wire [16-1:0] node15978;
	wire [16-1:0] node15979;
	wire [16-1:0] node15980;
	wire [16-1:0] node15982;
	wire [16-1:0] node15983;
	wire [16-1:0] node15987;
	wire [16-1:0] node15989;
	wire [16-1:0] node15990;
	wire [16-1:0] node15992;
	wire [16-1:0] node15996;
	wire [16-1:0] node15997;
	wire [16-1:0] node15998;
	wire [16-1:0] node16000;
	wire [16-1:0] node16001;
	wire [16-1:0] node16004;
	wire [16-1:0] node16005;
	wire [16-1:0] node16009;
	wire [16-1:0] node16011;
	wire [16-1:0] node16014;
	wire [16-1:0] node16015;
	wire [16-1:0] node16017;
	wire [16-1:0] node16021;
	wire [16-1:0] node16022;
	wire [16-1:0] node16023;
	wire [16-1:0] node16024;
	wire [16-1:0] node16025;
	wire [16-1:0] node16027;
	wire [16-1:0] node16030;
	wire [16-1:0] node16031;
	wire [16-1:0] node16034;
	wire [16-1:0] node16037;
	wire [16-1:0] node16039;
	wire [16-1:0] node16040;
	wire [16-1:0] node16043;
	wire [16-1:0] node16046;
	wire [16-1:0] node16047;
	wire [16-1:0] node16048;
	wire [16-1:0] node16050;
	wire [16-1:0] node16053;
	wire [16-1:0] node16054;
	wire [16-1:0] node16057;
	wire [16-1:0] node16058;
	wire [16-1:0] node16062;
	wire [16-1:0] node16063;
	wire [16-1:0] node16065;
	wire [16-1:0] node16067;
	wire [16-1:0] node16070;
	wire [16-1:0] node16071;
	wire [16-1:0] node16074;
	wire [16-1:0] node16077;
	wire [16-1:0] node16078;
	wire [16-1:0] node16079;
	wire [16-1:0] node16080;
	wire [16-1:0] node16081;
	wire [16-1:0] node16084;
	wire [16-1:0] node16085;
	wire [16-1:0] node16086;
	wire [16-1:0] node16091;
	wire [16-1:0] node16092;
	wire [16-1:0] node16095;
	wire [16-1:0] node16098;
	wire [16-1:0] node16099;
	wire [16-1:0] node16101;
	wire [16-1:0] node16104;
	wire [16-1:0] node16105;
	wire [16-1:0] node16108;
	wire [16-1:0] node16110;
	wire [16-1:0] node16112;
	wire [16-1:0] node16115;
	wire [16-1:0] node16116;
	wire [16-1:0] node16117;
	wire [16-1:0] node16119;
	wire [16-1:0] node16122;
	wire [16-1:0] node16124;
	wire [16-1:0] node16125;
	wire [16-1:0] node16127;
	wire [16-1:0] node16130;
	wire [16-1:0] node16133;
	wire [16-1:0] node16134;
	wire [16-1:0] node16137;
	wire [16-1:0] node16138;
	wire [16-1:0] node16140;
	wire [16-1:0] node16144;
	wire [16-1:0] node16145;
	wire [16-1:0] node16146;
	wire [16-1:0] node16147;
	wire [16-1:0] node16148;
	wire [16-1:0] node16149;
	wire [16-1:0] node16150;
	wire [16-1:0] node16151;
	wire [16-1:0] node16155;
	wire [16-1:0] node16156;
	wire [16-1:0] node16158;
	wire [16-1:0] node16162;
	wire [16-1:0] node16163;
	wire [16-1:0] node16166;
	wire [16-1:0] node16167;
	wire [16-1:0] node16168;
	wire [16-1:0] node16172;
	wire [16-1:0] node16173;
	wire [16-1:0] node16175;
	wire [16-1:0] node16179;
	wire [16-1:0] node16180;
	wire [16-1:0] node16181;
	wire [16-1:0] node16184;
	wire [16-1:0] node16187;
	wire [16-1:0] node16188;
	wire [16-1:0] node16190;
	wire [16-1:0] node16193;
	wire [16-1:0] node16194;
	wire [16-1:0] node16198;
	wire [16-1:0] node16199;
	wire [16-1:0] node16200;
	wire [16-1:0] node16201;
	wire [16-1:0] node16202;
	wire [16-1:0] node16203;
	wire [16-1:0] node16207;
	wire [16-1:0] node16210;
	wire [16-1:0] node16211;
	wire [16-1:0] node16215;
	wire [16-1:0] node16216;
	wire [16-1:0] node16218;
	wire [16-1:0] node16219;
	wire [16-1:0] node16222;
	wire [16-1:0] node16226;
	wire [16-1:0] node16227;
	wire [16-1:0] node16228;
	wire [16-1:0] node16229;
	wire [16-1:0] node16230;
	wire [16-1:0] node16234;
	wire [16-1:0] node16237;
	wire [16-1:0] node16240;
	wire [16-1:0] node16241;
	wire [16-1:0] node16243;
	wire [16-1:0] node16246;
	wire [16-1:0] node16247;
	wire [16-1:0] node16248;
	wire [16-1:0] node16252;
	wire [16-1:0] node16255;
	wire [16-1:0] node16256;
	wire [16-1:0] node16257;
	wire [16-1:0] node16258;
	wire [16-1:0] node16259;
	wire [16-1:0] node16260;
	wire [16-1:0] node16264;
	wire [16-1:0] node16265;
	wire [16-1:0] node16269;
	wire [16-1:0] node16271;
	wire [16-1:0] node16272;
	wire [16-1:0] node16273;
	wire [16-1:0] node16275;
	wire [16-1:0] node16280;
	wire [16-1:0] node16281;
	wire [16-1:0] node16282;
	wire [16-1:0] node16283;
	wire [16-1:0] node16286;
	wire [16-1:0] node16289;
	wire [16-1:0] node16290;
	wire [16-1:0] node16293;
	wire [16-1:0] node16294;
	wire [16-1:0] node16296;
	wire [16-1:0] node16300;
	wire [16-1:0] node16301;
	wire [16-1:0] node16303;
	wire [16-1:0] node16306;
	wire [16-1:0] node16307;
	wire [16-1:0] node16310;
	wire [16-1:0] node16313;
	wire [16-1:0] node16314;
	wire [16-1:0] node16315;
	wire [16-1:0] node16316;
	wire [16-1:0] node16319;
	wire [16-1:0] node16320;
	wire [16-1:0] node16323;
	wire [16-1:0] node16324;
	wire [16-1:0] node16328;
	wire [16-1:0] node16329;
	wire [16-1:0] node16331;
	wire [16-1:0] node16333;
	wire [16-1:0] node16336;
	wire [16-1:0] node16338;
	wire [16-1:0] node16341;
	wire [16-1:0] node16342;
	wire [16-1:0] node16343;
	wire [16-1:0] node16346;
	wire [16-1:0] node16347;
	wire [16-1:0] node16348;
	wire [16-1:0] node16352;
	wire [16-1:0] node16355;
	wire [16-1:0] node16356;
	wire [16-1:0] node16357;
	wire [16-1:0] node16361;
	wire [16-1:0] node16363;
	wire [16-1:0] node16366;
	wire [16-1:0] node16367;
	wire [16-1:0] node16368;
	wire [16-1:0] node16369;
	wire [16-1:0] node16370;
	wire [16-1:0] node16371;
	wire [16-1:0] node16374;
	wire [16-1:0] node16375;
	wire [16-1:0] node16376;
	wire [16-1:0] node16378;
	wire [16-1:0] node16383;
	wire [16-1:0] node16384;
	wire [16-1:0] node16385;
	wire [16-1:0] node16388;
	wire [16-1:0] node16390;
	wire [16-1:0] node16394;
	wire [16-1:0] node16395;
	wire [16-1:0] node16396;
	wire [16-1:0] node16398;
	wire [16-1:0] node16401;
	wire [16-1:0] node16402;
	wire [16-1:0] node16405;
	wire [16-1:0] node16408;
	wire [16-1:0] node16409;
	wire [16-1:0] node16410;
	wire [16-1:0] node16411;
	wire [16-1:0] node16415;
	wire [16-1:0] node16416;
	wire [16-1:0] node16420;
	wire [16-1:0] node16421;
	wire [16-1:0] node16424;
	wire [16-1:0] node16427;
	wire [16-1:0] node16428;
	wire [16-1:0] node16429;
	wire [16-1:0] node16430;
	wire [16-1:0] node16432;
	wire [16-1:0] node16434;
	wire [16-1:0] node16437;
	wire [16-1:0] node16439;
	wire [16-1:0] node16442;
	wire [16-1:0] node16444;
	wire [16-1:0] node16445;
	wire [16-1:0] node16449;
	wire [16-1:0] node16450;
	wire [16-1:0] node16452;
	wire [16-1:0] node16454;
	wire [16-1:0] node16455;
	wire [16-1:0] node16456;
	wire [16-1:0] node16461;
	wire [16-1:0] node16462;
	wire [16-1:0] node16464;
	wire [16-1:0] node16465;
	wire [16-1:0] node16469;
	wire [16-1:0] node16470;
	wire [16-1:0] node16473;
	wire [16-1:0] node16475;
	wire [16-1:0] node16478;
	wire [16-1:0] node16479;
	wire [16-1:0] node16480;
	wire [16-1:0] node16481;
	wire [16-1:0] node16482;
	wire [16-1:0] node16485;
	wire [16-1:0] node16487;
	wire [16-1:0] node16490;
	wire [16-1:0] node16491;
	wire [16-1:0] node16493;
	wire [16-1:0] node16494;
	wire [16-1:0] node16498;
	wire [16-1:0] node16500;
	wire [16-1:0] node16502;
	wire [16-1:0] node16505;
	wire [16-1:0] node16506;
	wire [16-1:0] node16507;
	wire [16-1:0] node16509;
	wire [16-1:0] node16510;
	wire [16-1:0] node16514;
	wire [16-1:0] node16517;
	wire [16-1:0] node16519;
	wire [16-1:0] node16520;
	wire [16-1:0] node16523;
	wire [16-1:0] node16526;
	wire [16-1:0] node16527;
	wire [16-1:0] node16528;
	wire [16-1:0] node16529;
	wire [16-1:0] node16530;
	wire [16-1:0] node16534;
	wire [16-1:0] node16537;
	wire [16-1:0] node16540;
	wire [16-1:0] node16541;
	wire [16-1:0] node16542;
	wire [16-1:0] node16543;
	wire [16-1:0] node16545;
	wire [16-1:0] node16549;
	wire [16-1:0] node16551;
	wire [16-1:0] node16552;
	wire [16-1:0] node16556;
	wire [16-1:0] node16559;
	wire [16-1:0] node16560;
	wire [16-1:0] node16561;
	wire [16-1:0] node16562;
	wire [16-1:0] node16563;
	wire [16-1:0] node16564;
	wire [16-1:0] node16565;
	wire [16-1:0] node16566;
	wire [16-1:0] node16567;
	wire [16-1:0] node16568;
	wire [16-1:0] node16570;
	wire [16-1:0] node16571;
	wire [16-1:0] node16576;
	wire [16-1:0] node16579;
	wire [16-1:0] node16580;
	wire [16-1:0] node16581;
	wire [16-1:0] node16585;
	wire [16-1:0] node16587;
	wire [16-1:0] node16589;
	wire [16-1:0] node16592;
	wire [16-1:0] node16593;
	wire [16-1:0] node16594;
	wire [16-1:0] node16596;
	wire [16-1:0] node16597;
	wire [16-1:0] node16602;
	wire [16-1:0] node16603;
	wire [16-1:0] node16604;
	wire [16-1:0] node16605;
	wire [16-1:0] node16609;
	wire [16-1:0] node16612;
	wire [16-1:0] node16613;
	wire [16-1:0] node16617;
	wire [16-1:0] node16618;
	wire [16-1:0] node16619;
	wire [16-1:0] node16620;
	wire [16-1:0] node16621;
	wire [16-1:0] node16624;
	wire [16-1:0] node16626;
	wire [16-1:0] node16627;
	wire [16-1:0] node16631;
	wire [16-1:0] node16632;
	wire [16-1:0] node16636;
	wire [16-1:0] node16637;
	wire [16-1:0] node16639;
	wire [16-1:0] node16640;
	wire [16-1:0] node16642;
	wire [16-1:0] node16646;
	wire [16-1:0] node16649;
	wire [16-1:0] node16650;
	wire [16-1:0] node16651;
	wire [16-1:0] node16655;
	wire [16-1:0] node16656;
	wire [16-1:0] node16658;
	wire [16-1:0] node16659;
	wire [16-1:0] node16661;
	wire [16-1:0] node16666;
	wire [16-1:0] node16667;
	wire [16-1:0] node16668;
	wire [16-1:0] node16669;
	wire [16-1:0] node16670;
	wire [16-1:0] node16673;
	wire [16-1:0] node16674;
	wire [16-1:0] node16679;
	wire [16-1:0] node16680;
	wire [16-1:0] node16683;
	wire [16-1:0] node16684;
	wire [16-1:0] node16685;
	wire [16-1:0] node16686;
	wire [16-1:0] node16688;
	wire [16-1:0] node16692;
	wire [16-1:0] node16693;
	wire [16-1:0] node16697;
	wire [16-1:0] node16700;
	wire [16-1:0] node16701;
	wire [16-1:0] node16702;
	wire [16-1:0] node16703;
	wire [16-1:0] node16704;
	wire [16-1:0] node16707;
	wire [16-1:0] node16711;
	wire [16-1:0] node16712;
	wire [16-1:0] node16713;
	wire [16-1:0] node16716;
	wire [16-1:0] node16719;
	wire [16-1:0] node16720;
	wire [16-1:0] node16724;
	wire [16-1:0] node16725;
	wire [16-1:0] node16726;
	wire [16-1:0] node16728;
	wire [16-1:0] node16732;
	wire [16-1:0] node16733;
	wire [16-1:0] node16736;
	wire [16-1:0] node16739;
	wire [16-1:0] node16740;
	wire [16-1:0] node16741;
	wire [16-1:0] node16742;
	wire [16-1:0] node16743;
	wire [16-1:0] node16744;
	wire [16-1:0] node16745;
	wire [16-1:0] node16747;
	wire [16-1:0] node16750;
	wire [16-1:0] node16752;
	wire [16-1:0] node16756;
	wire [16-1:0] node16757;
	wire [16-1:0] node16759;
	wire [16-1:0] node16762;
	wire [16-1:0] node16764;
	wire [16-1:0] node16767;
	wire [16-1:0] node16768;
	wire [16-1:0] node16769;
	wire [16-1:0] node16770;
	wire [16-1:0] node16773;
	wire [16-1:0] node16776;
	wire [16-1:0] node16777;
	wire [16-1:0] node16780;
	wire [16-1:0] node16783;
	wire [16-1:0] node16784;
	wire [16-1:0] node16785;
	wire [16-1:0] node16790;
	wire [16-1:0] node16791;
	wire [16-1:0] node16792;
	wire [16-1:0] node16793;
	wire [16-1:0] node16794;
	wire [16-1:0] node16798;
	wire [16-1:0] node16801;
	wire [16-1:0] node16802;
	wire [16-1:0] node16804;
	wire [16-1:0] node16807;
	wire [16-1:0] node16808;
	wire [16-1:0] node16811;
	wire [16-1:0] node16814;
	wire [16-1:0] node16815;
	wire [16-1:0] node16816;
	wire [16-1:0] node16818;
	wire [16-1:0] node16820;
	wire [16-1:0] node16821;
	wire [16-1:0] node16825;
	wire [16-1:0] node16828;
	wire [16-1:0] node16830;
	wire [16-1:0] node16831;
	wire [16-1:0] node16835;
	wire [16-1:0] node16836;
	wire [16-1:0] node16837;
	wire [16-1:0] node16838;
	wire [16-1:0] node16839;
	wire [16-1:0] node16841;
	wire [16-1:0] node16844;
	wire [16-1:0] node16845;
	wire [16-1:0] node16849;
	wire [16-1:0] node16850;
	wire [16-1:0] node16851;
	wire [16-1:0] node16854;
	wire [16-1:0] node16856;
	wire [16-1:0] node16859;
	wire [16-1:0] node16860;
	wire [16-1:0] node16864;
	wire [16-1:0] node16865;
	wire [16-1:0] node16868;
	wire [16-1:0] node16869;
	wire [16-1:0] node16871;
	wire [16-1:0] node16873;
	wire [16-1:0] node16876;
	wire [16-1:0] node16877;
	wire [16-1:0] node16881;
	wire [16-1:0] node16882;
	wire [16-1:0] node16883;
	wire [16-1:0] node16884;
	wire [16-1:0] node16885;
	wire [16-1:0] node16890;
	wire [16-1:0] node16891;
	wire [16-1:0] node16892;
	wire [16-1:0] node16895;
	wire [16-1:0] node16897;
	wire [16-1:0] node16898;
	wire [16-1:0] node16902;
	wire [16-1:0] node16904;
	wire [16-1:0] node16905;
	wire [16-1:0] node16909;
	wire [16-1:0] node16910;
	wire [16-1:0] node16911;
	wire [16-1:0] node16912;
	wire [16-1:0] node16916;
	wire [16-1:0] node16917;
	wire [16-1:0] node16918;
	wire [16-1:0] node16923;
	wire [16-1:0] node16924;
	wire [16-1:0] node16926;
	wire [16-1:0] node16929;
	wire [16-1:0] node16931;
	wire [16-1:0] node16932;
	wire [16-1:0] node16934;
	wire [16-1:0] node16938;
	wire [16-1:0] node16939;
	wire [16-1:0] node16940;
	wire [16-1:0] node16941;
	wire [16-1:0] node16942;
	wire [16-1:0] node16943;
	wire [16-1:0] node16944;
	wire [16-1:0] node16945;
	wire [16-1:0] node16950;
	wire [16-1:0] node16951;
	wire [16-1:0] node16952;
	wire [16-1:0] node16956;
	wire [16-1:0] node16957;
	wire [16-1:0] node16961;
	wire [16-1:0] node16962;
	wire [16-1:0] node16963;
	wire [16-1:0] node16965;
	wire [16-1:0] node16968;
	wire [16-1:0] node16969;
	wire [16-1:0] node16973;
	wire [16-1:0] node16974;
	wire [16-1:0] node16975;
	wire [16-1:0] node16978;
	wire [16-1:0] node16981;
	wire [16-1:0] node16984;
	wire [16-1:0] node16985;
	wire [16-1:0] node16986;
	wire [16-1:0] node16987;
	wire [16-1:0] node16990;
	wire [16-1:0] node16991;
	wire [16-1:0] node16992;
	wire [16-1:0] node16994;
	wire [16-1:0] node16998;
	wire [16-1:0] node17001;
	wire [16-1:0] node17002;
	wire [16-1:0] node17005;
	wire [16-1:0] node17006;
	wire [16-1:0] node17010;
	wire [16-1:0] node17011;
	wire [16-1:0] node17012;
	wire [16-1:0] node17013;
	wire [16-1:0] node17014;
	wire [16-1:0] node17018;
	wire [16-1:0] node17020;
	wire [16-1:0] node17021;
	wire [16-1:0] node17025;
	wire [16-1:0] node17026;
	wire [16-1:0] node17029;
	wire [16-1:0] node17031;
	wire [16-1:0] node17034;
	wire [16-1:0] node17035;
	wire [16-1:0] node17036;
	wire [16-1:0] node17039;
	wire [16-1:0] node17040;
	wire [16-1:0] node17044;
	wire [16-1:0] node17047;
	wire [16-1:0] node17048;
	wire [16-1:0] node17049;
	wire [16-1:0] node17050;
	wire [16-1:0] node17051;
	wire [16-1:0] node17052;
	wire [16-1:0] node17056;
	wire [16-1:0] node17058;
	wire [16-1:0] node17059;
	wire [16-1:0] node17061;
	wire [16-1:0] node17065;
	wire [16-1:0] node17066;
	wire [16-1:0] node17068;
	wire [16-1:0] node17072;
	wire [16-1:0] node17073;
	wire [16-1:0] node17074;
	wire [16-1:0] node17075;
	wire [16-1:0] node17078;
	wire [16-1:0] node17081;
	wire [16-1:0] node17082;
	wire [16-1:0] node17083;
	wire [16-1:0] node17087;
	wire [16-1:0] node17090;
	wire [16-1:0] node17091;
	wire [16-1:0] node17093;
	wire [16-1:0] node17097;
	wire [16-1:0] node17098;
	wire [16-1:0] node17099;
	wire [16-1:0] node17100;
	wire [16-1:0] node17101;
	wire [16-1:0] node17104;
	wire [16-1:0] node17107;
	wire [16-1:0] node17108;
	wire [16-1:0] node17110;
	wire [16-1:0] node17114;
	wire [16-1:0] node17115;
	wire [16-1:0] node17118;
	wire [16-1:0] node17120;
	wire [16-1:0] node17123;
	wire [16-1:0] node17124;
	wire [16-1:0] node17125;
	wire [16-1:0] node17127;
	wire [16-1:0] node17130;
	wire [16-1:0] node17131;
	wire [16-1:0] node17135;
	wire [16-1:0] node17136;
	wire [16-1:0] node17139;
	wire [16-1:0] node17140;
	wire [16-1:0] node17141;
	wire [16-1:0] node17145;
	wire [16-1:0] node17147;
	wire [16-1:0] node17150;
	wire [16-1:0] node17151;
	wire [16-1:0] node17152;
	wire [16-1:0] node17153;
	wire [16-1:0] node17154;
	wire [16-1:0] node17155;
	wire [16-1:0] node17157;
	wire [16-1:0] node17160;
	wire [16-1:0] node17161;
	wire [16-1:0] node17165;
	wire [16-1:0] node17166;
	wire [16-1:0] node17168;
	wire [16-1:0] node17172;
	wire [16-1:0] node17173;
	wire [16-1:0] node17175;
	wire [16-1:0] node17178;
	wire [16-1:0] node17179;
	wire [16-1:0] node17183;
	wire [16-1:0] node17184;
	wire [16-1:0] node17185;
	wire [16-1:0] node17186;
	wire [16-1:0] node17187;
	wire [16-1:0] node17192;
	wire [16-1:0] node17193;
	wire [16-1:0] node17195;
	wire [16-1:0] node17198;
	wire [16-1:0] node17199;
	wire [16-1:0] node17203;
	wire [16-1:0] node17204;
	wire [16-1:0] node17205;
	wire [16-1:0] node17208;
	wire [16-1:0] node17209;
	wire [16-1:0] node17212;
	wire [16-1:0] node17215;
	wire [16-1:0] node17216;
	wire [16-1:0] node17218;
	wire [16-1:0] node17221;
	wire [16-1:0] node17222;
	wire [16-1:0] node17226;
	wire [16-1:0] node17227;
	wire [16-1:0] node17228;
	wire [16-1:0] node17229;
	wire [16-1:0] node17230;
	wire [16-1:0] node17231;
	wire [16-1:0] node17234;
	wire [16-1:0] node17236;
	wire [16-1:0] node17239;
	wire [16-1:0] node17242;
	wire [16-1:0] node17243;
	wire [16-1:0] node17245;
	wire [16-1:0] node17248;
	wire [16-1:0] node17250;
	wire [16-1:0] node17252;
	wire [16-1:0] node17255;
	wire [16-1:0] node17256;
	wire [16-1:0] node17258;
	wire [16-1:0] node17259;
	wire [16-1:0] node17262;
	wire [16-1:0] node17265;
	wire [16-1:0] node17266;
	wire [16-1:0] node17268;
	wire [16-1:0] node17271;
	wire [16-1:0] node17272;
	wire [16-1:0] node17274;
	wire [16-1:0] node17277;
	wire [16-1:0] node17280;
	wire [16-1:0] node17281;
	wire [16-1:0] node17282;
	wire [16-1:0] node17283;
	wire [16-1:0] node17285;
	wire [16-1:0] node17286;
	wire [16-1:0] node17290;
	wire [16-1:0] node17292;
	wire [16-1:0] node17295;
	wire [16-1:0] node17296;
	wire [16-1:0] node17297;
	wire [16-1:0] node17299;
	wire [16-1:0] node17301;
	wire [16-1:0] node17305;
	wire [16-1:0] node17306;
	wire [16-1:0] node17310;
	wire [16-1:0] node17311;
	wire [16-1:0] node17312;
	wire [16-1:0] node17316;
	wire [16-1:0] node17318;
	wire [16-1:0] node17319;
	wire [16-1:0] node17320;
	wire [16-1:0] node17324;
	wire [16-1:0] node17326;
	wire [16-1:0] node17327;
	wire [16-1:0] node17331;
	wire [16-1:0] node17332;
	wire [16-1:0] node17333;
	wire [16-1:0] node17334;
	wire [16-1:0] node17335;
	wire [16-1:0] node17336;
	wire [16-1:0] node17337;
	wire [16-1:0] node17338;
	wire [16-1:0] node17339;
	wire [16-1:0] node17343;
	wire [16-1:0] node17345;
	wire [16-1:0] node17346;
	wire [16-1:0] node17350;
	wire [16-1:0] node17353;
	wire [16-1:0] node17354;
	wire [16-1:0] node17355;
	wire [16-1:0] node17356;
	wire [16-1:0] node17359;
	wire [16-1:0] node17362;
	wire [16-1:0] node17363;
	wire [16-1:0] node17367;
	wire [16-1:0] node17368;
	wire [16-1:0] node17370;
	wire [16-1:0] node17374;
	wire [16-1:0] node17375;
	wire [16-1:0] node17376;
	wire [16-1:0] node17377;
	wire [16-1:0] node17378;
	wire [16-1:0] node17381;
	wire [16-1:0] node17384;
	wire [16-1:0] node17385;
	wire [16-1:0] node17388;
	wire [16-1:0] node17390;
	wire [16-1:0] node17393;
	wire [16-1:0] node17394;
	wire [16-1:0] node17396;
	wire [16-1:0] node17399;
	wire [16-1:0] node17401;
	wire [16-1:0] node17404;
	wire [16-1:0] node17405;
	wire [16-1:0] node17408;
	wire [16-1:0] node17410;
	wire [16-1:0] node17412;
	wire [16-1:0] node17414;
	wire [16-1:0] node17417;
	wire [16-1:0] node17418;
	wire [16-1:0] node17419;
	wire [16-1:0] node17420;
	wire [16-1:0] node17421;
	wire [16-1:0] node17424;
	wire [16-1:0] node17427;
	wire [16-1:0] node17428;
	wire [16-1:0] node17431;
	wire [16-1:0] node17433;
	wire [16-1:0] node17434;
	wire [16-1:0] node17438;
	wire [16-1:0] node17439;
	wire [16-1:0] node17441;
	wire [16-1:0] node17442;
	wire [16-1:0] node17445;
	wire [16-1:0] node17448;
	wire [16-1:0] node17449;
	wire [16-1:0] node17452;
	wire [16-1:0] node17455;
	wire [16-1:0] node17456;
	wire [16-1:0] node17457;
	wire [16-1:0] node17458;
	wire [16-1:0] node17460;
	wire [16-1:0] node17463;
	wire [16-1:0] node17464;
	wire [16-1:0] node17465;
	wire [16-1:0] node17470;
	wire [16-1:0] node17471;
	wire [16-1:0] node17472;
	wire [16-1:0] node17473;
	wire [16-1:0] node17475;
	wire [16-1:0] node17481;
	wire [16-1:0] node17482;
	wire [16-1:0] node17483;
	wire [16-1:0] node17484;
	wire [16-1:0] node17488;
	wire [16-1:0] node17490;
	wire [16-1:0] node17493;
	wire [16-1:0] node17495;
	wire [16-1:0] node17496;
	wire [16-1:0] node17499;
	wire [16-1:0] node17501;
	wire [16-1:0] node17504;
	wire [16-1:0] node17505;
	wire [16-1:0] node17506;
	wire [16-1:0] node17507;
	wire [16-1:0] node17508;
	wire [16-1:0] node17509;
	wire [16-1:0] node17511;
	wire [16-1:0] node17514;
	wire [16-1:0] node17515;
	wire [16-1:0] node17519;
	wire [16-1:0] node17520;
	wire [16-1:0] node17521;
	wire [16-1:0] node17525;
	wire [16-1:0] node17527;
	wire [16-1:0] node17530;
	wire [16-1:0] node17531;
	wire [16-1:0] node17532;
	wire [16-1:0] node17533;
	wire [16-1:0] node17536;
	wire [16-1:0] node17539;
	wire [16-1:0] node17540;
	wire [16-1:0] node17541;
	wire [16-1:0] node17543;
	wire [16-1:0] node17548;
	wire [16-1:0] node17549;
	wire [16-1:0] node17551;
	wire [16-1:0] node17552;
	wire [16-1:0] node17554;
	wire [16-1:0] node17558;
	wire [16-1:0] node17561;
	wire [16-1:0] node17562;
	wire [16-1:0] node17563;
	wire [16-1:0] node17564;
	wire [16-1:0] node17566;
	wire [16-1:0] node17567;
	wire [16-1:0] node17572;
	wire [16-1:0] node17573;
	wire [16-1:0] node17574;
	wire [16-1:0] node17577;
	wire [16-1:0] node17580;
	wire [16-1:0] node17583;
	wire [16-1:0] node17584;
	wire [16-1:0] node17585;
	wire [16-1:0] node17587;
	wire [16-1:0] node17590;
	wire [16-1:0] node17593;
	wire [16-1:0] node17594;
	wire [16-1:0] node17597;
	wire [16-1:0] node17599;
	wire [16-1:0] node17601;
	wire [16-1:0] node17604;
	wire [16-1:0] node17605;
	wire [16-1:0] node17606;
	wire [16-1:0] node17607;
	wire [16-1:0] node17608;
	wire [16-1:0] node17609;
	wire [16-1:0] node17613;
	wire [16-1:0] node17614;
	wire [16-1:0] node17617;
	wire [16-1:0] node17620;
	wire [16-1:0] node17621;
	wire [16-1:0] node17623;
	wire [16-1:0] node17625;
	wire [16-1:0] node17629;
	wire [16-1:0] node17630;
	wire [16-1:0] node17631;
	wire [16-1:0] node17632;
	wire [16-1:0] node17633;
	wire [16-1:0] node17638;
	wire [16-1:0] node17639;
	wire [16-1:0] node17643;
	wire [16-1:0] node17644;
	wire [16-1:0] node17646;
	wire [16-1:0] node17649;
	wire [16-1:0] node17651;
	wire [16-1:0] node17654;
	wire [16-1:0] node17655;
	wire [16-1:0] node17656;
	wire [16-1:0] node17657;
	wire [16-1:0] node17658;
	wire [16-1:0] node17663;
	wire [16-1:0] node17664;
	wire [16-1:0] node17665;
	wire [16-1:0] node17668;
	wire [16-1:0] node17671;
	wire [16-1:0] node17672;
	wire [16-1:0] node17675;
	wire [16-1:0] node17678;
	wire [16-1:0] node17679;
	wire [16-1:0] node17680;
	wire [16-1:0] node17681;
	wire [16-1:0] node17684;
	wire [16-1:0] node17687;
	wire [16-1:0] node17688;
	wire [16-1:0] node17691;
	wire [16-1:0] node17692;
	wire [16-1:0] node17694;
	wire [16-1:0] node17698;
	wire [16-1:0] node17699;
	wire [16-1:0] node17701;
	wire [16-1:0] node17704;
	wire [16-1:0] node17706;
	wire [16-1:0] node17709;
	wire [16-1:0] node17710;
	wire [16-1:0] node17711;
	wire [16-1:0] node17712;
	wire [16-1:0] node17713;
	wire [16-1:0] node17714;
	wire [16-1:0] node17715;
	wire [16-1:0] node17717;
	wire [16-1:0] node17720;
	wire [16-1:0] node17721;
	wire [16-1:0] node17724;
	wire [16-1:0] node17726;
	wire [16-1:0] node17729;
	wire [16-1:0] node17730;
	wire [16-1:0] node17731;
	wire [16-1:0] node17735;
	wire [16-1:0] node17737;
	wire [16-1:0] node17740;
	wire [16-1:0] node17741;
	wire [16-1:0] node17742;
	wire [16-1:0] node17746;
	wire [16-1:0] node17747;
	wire [16-1:0] node17748;
	wire [16-1:0] node17751;
	wire [16-1:0] node17753;
	wire [16-1:0] node17754;
	wire [16-1:0] node17759;
	wire [16-1:0] node17760;
	wire [16-1:0] node17761;
	wire [16-1:0] node17762;
	wire [16-1:0] node17765;
	wire [16-1:0] node17767;
	wire [16-1:0] node17770;
	wire [16-1:0] node17771;
	wire [16-1:0] node17773;
	wire [16-1:0] node17776;
	wire [16-1:0] node17777;
	wire [16-1:0] node17780;
	wire [16-1:0] node17781;
	wire [16-1:0] node17785;
	wire [16-1:0] node17787;
	wire [16-1:0] node17788;
	wire [16-1:0] node17791;
	wire [16-1:0] node17794;
	wire [16-1:0] node17795;
	wire [16-1:0] node17796;
	wire [16-1:0] node17797;
	wire [16-1:0] node17798;
	wire [16-1:0] node17801;
	wire [16-1:0] node17802;
	wire [16-1:0] node17806;
	wire [16-1:0] node17807;
	wire [16-1:0] node17810;
	wire [16-1:0] node17811;
	wire [16-1:0] node17813;
	wire [16-1:0] node17817;
	wire [16-1:0] node17818;
	wire [16-1:0] node17819;
	wire [16-1:0] node17820;
	wire [16-1:0] node17823;
	wire [16-1:0] node17825;
	wire [16-1:0] node17828;
	wire [16-1:0] node17830;
	wire [16-1:0] node17833;
	wire [16-1:0] node17834;
	wire [16-1:0] node17835;
	wire [16-1:0] node17836;
	wire [16-1:0] node17840;
	wire [16-1:0] node17844;
	wire [16-1:0] node17845;
	wire [16-1:0] node17846;
	wire [16-1:0] node17848;
	wire [16-1:0] node17849;
	wire [16-1:0] node17850;
	wire [16-1:0] node17851;
	wire [16-1:0] node17856;
	wire [16-1:0] node17859;
	wire [16-1:0] node17861;
	wire [16-1:0] node17863;
	wire [16-1:0] node17864;
	wire [16-1:0] node17868;
	wire [16-1:0] node17869;
	wire [16-1:0] node17870;
	wire [16-1:0] node17872;
	wire [16-1:0] node17875;
	wire [16-1:0] node17876;
	wire [16-1:0] node17879;
	wire [16-1:0] node17881;
	wire [16-1:0] node17882;
	wire [16-1:0] node17886;
	wire [16-1:0] node17887;
	wire [16-1:0] node17888;
	wire [16-1:0] node17889;
	wire [16-1:0] node17892;
	wire [16-1:0] node17894;
	wire [16-1:0] node17897;
	wire [16-1:0] node17900;
	wire [16-1:0] node17903;
	wire [16-1:0] node17904;
	wire [16-1:0] node17905;
	wire [16-1:0] node17906;
	wire [16-1:0] node17907;
	wire [16-1:0] node17908;
	wire [16-1:0] node17909;
	wire [16-1:0] node17910;
	wire [16-1:0] node17915;
	wire [16-1:0] node17916;
	wire [16-1:0] node17919;
	wire [16-1:0] node17920;
	wire [16-1:0] node17924;
	wire [16-1:0] node17926;
	wire [16-1:0] node17929;
	wire [16-1:0] node17930;
	wire [16-1:0] node17931;
	wire [16-1:0] node17932;
	wire [16-1:0] node17936;
	wire [16-1:0] node17937;
	wire [16-1:0] node17940;
	wire [16-1:0] node17943;
	wire [16-1:0] node17944;
	wire [16-1:0] node17946;
	wire [16-1:0] node17949;
	wire [16-1:0] node17952;
	wire [16-1:0] node17953;
	wire [16-1:0] node17954;
	wire [16-1:0] node17955;
	wire [16-1:0] node17957;
	wire [16-1:0] node17960;
	wire [16-1:0] node17963;
	wire [16-1:0] node17964;
	wire [16-1:0] node17965;
	wire [16-1:0] node17968;
	wire [16-1:0] node17971;
	wire [16-1:0] node17972;
	wire [16-1:0] node17975;
	wire [16-1:0] node17978;
	wire [16-1:0] node17979;
	wire [16-1:0] node17980;
	wire [16-1:0] node17982;
	wire [16-1:0] node17985;
	wire [16-1:0] node17987;
	wire [16-1:0] node17989;
	wire [16-1:0] node17992;
	wire [16-1:0] node17993;
	wire [16-1:0] node17995;
	wire [16-1:0] node17999;
	wire [16-1:0] node18000;
	wire [16-1:0] node18001;
	wire [16-1:0] node18002;
	wire [16-1:0] node18004;
	wire [16-1:0] node18005;
	wire [16-1:0] node18009;
	wire [16-1:0] node18010;
	wire [16-1:0] node18011;
	wire [16-1:0] node18012;
	wire [16-1:0] node18017;
	wire [16-1:0] node18018;
	wire [16-1:0] node18022;
	wire [16-1:0] node18023;
	wire [16-1:0] node18024;
	wire [16-1:0] node18025;
	wire [16-1:0] node18026;
	wire [16-1:0] node18030;
	wire [16-1:0] node18033;
	wire [16-1:0] node18036;
	wire [16-1:0] node18037;
	wire [16-1:0] node18039;
	wire [16-1:0] node18042;
	wire [16-1:0] node18044;
	wire [16-1:0] node18045;
	wire [16-1:0] node18049;
	wire [16-1:0] node18050;
	wire [16-1:0] node18051;
	wire [16-1:0] node18052;
	wire [16-1:0] node18053;
	wire [16-1:0] node18057;
	wire [16-1:0] node18058;
	wire [16-1:0] node18061;
	wire [16-1:0] node18064;
	wire [16-1:0] node18065;
	wire [16-1:0] node18066;
	wire [16-1:0] node18069;
	wire [16-1:0] node18070;
	wire [16-1:0] node18072;
	wire [16-1:0] node18075;
	wire [16-1:0] node18076;
	wire [16-1:0] node18080;
	wire [16-1:0] node18081;
	wire [16-1:0] node18084;
	wire [16-1:0] node18086;
	wire [16-1:0] node18089;
	wire [16-1:0] node18090;
	wire [16-1:0] node18091;
	wire [16-1:0] node18092;
	wire [16-1:0] node18095;
	wire [16-1:0] node18098;
	wire [16-1:0] node18099;
	wire [16-1:0] node18102;
	wire [16-1:0] node18105;
	wire [16-1:0] node18106;
	wire [16-1:0] node18108;
	wire [16-1:0] node18111;
	wire [16-1:0] node18112;
	wire [16-1:0] node18113;
	wire [16-1:0] node18117;
	wire [16-1:0] node18118;
	wire [16-1:0] node18121;
	wire [16-1:0] node18124;
	wire [16-1:0] node18125;
	wire [16-1:0] node18126;
	wire [16-1:0] node18127;
	wire [16-1:0] node18128;
	wire [16-1:0] node18129;
	wire [16-1:0] node18130;
	wire [16-1:0] node18131;
	wire [16-1:0] node18132;
	wire [16-1:0] node18133;
	wire [16-1:0] node18134;
	wire [16-1:0] node18135;
	wire [16-1:0] node18139;
	wire [16-1:0] node18142;
	wire [16-1:0] node18143;
	wire [16-1:0] node18144;
	wire [16-1:0] node18145;
	wire [16-1:0] node18146;
	wire [16-1:0] node18152;
	wire [16-1:0] node18153;
	wire [16-1:0] node18155;
	wire [16-1:0] node18159;
	wire [16-1:0] node18160;
	wire [16-1:0] node18161;
	wire [16-1:0] node18163;
	wire [16-1:0] node18166;
	wire [16-1:0] node18169;
	wire [16-1:0] node18171;
	wire [16-1:0] node18172;
	wire [16-1:0] node18176;
	wire [16-1:0] node18177;
	wire [16-1:0] node18178;
	wire [16-1:0] node18179;
	wire [16-1:0] node18180;
	wire [16-1:0] node18181;
	wire [16-1:0] node18182;
	wire [16-1:0] node18188;
	wire [16-1:0] node18189;
	wire [16-1:0] node18192;
	wire [16-1:0] node18195;
	wire [16-1:0] node18197;
	wire [16-1:0] node18200;
	wire [16-1:0] node18201;
	wire [16-1:0] node18202;
	wire [16-1:0] node18205;
	wire [16-1:0] node18206;
	wire [16-1:0] node18209;
	wire [16-1:0] node18212;
	wire [16-1:0] node18214;
	wire [16-1:0] node18215;
	wire [16-1:0] node18219;
	wire [16-1:0] node18220;
	wire [16-1:0] node18221;
	wire [16-1:0] node18222;
	wire [16-1:0] node18223;
	wire [16-1:0] node18224;
	wire [16-1:0] node18227;
	wire [16-1:0] node18230;
	wire [16-1:0] node18232;
	wire [16-1:0] node18235;
	wire [16-1:0] node18236;
	wire [16-1:0] node18237;
	wire [16-1:0] node18241;
	wire [16-1:0] node18242;
	wire [16-1:0] node18246;
	wire [16-1:0] node18247;
	wire [16-1:0] node18248;
	wire [16-1:0] node18249;
	wire [16-1:0] node18252;
	wire [16-1:0] node18255;
	wire [16-1:0] node18256;
	wire [16-1:0] node18259;
	wire [16-1:0] node18262;
	wire [16-1:0] node18263;
	wire [16-1:0] node18266;
	wire [16-1:0] node18268;
	wire [16-1:0] node18271;
	wire [16-1:0] node18272;
	wire [16-1:0] node18273;
	wire [16-1:0] node18274;
	wire [16-1:0] node18276;
	wire [16-1:0] node18277;
	wire [16-1:0] node18280;
	wire [16-1:0] node18284;
	wire [16-1:0] node18286;
	wire [16-1:0] node18288;
	wire [16-1:0] node18291;
	wire [16-1:0] node18292;
	wire [16-1:0] node18293;
	wire [16-1:0] node18294;
	wire [16-1:0] node18297;
	wire [16-1:0] node18300;
	wire [16-1:0] node18301;
	wire [16-1:0] node18302;
	wire [16-1:0] node18307;
	wire [16-1:0] node18308;
	wire [16-1:0] node18312;
	wire [16-1:0] node18313;
	wire [16-1:0] node18314;
	wire [16-1:0] node18315;
	wire [16-1:0] node18316;
	wire [16-1:0] node18317;
	wire [16-1:0] node18319;
	wire [16-1:0] node18321;
	wire [16-1:0] node18324;
	wire [16-1:0] node18325;
	wire [16-1:0] node18327;
	wire [16-1:0] node18330;
	wire [16-1:0] node18331;
	wire [16-1:0] node18332;
	wire [16-1:0] node18336;
	wire [16-1:0] node18339;
	wire [16-1:0] node18340;
	wire [16-1:0] node18341;
	wire [16-1:0] node18344;
	wire [16-1:0] node18346;
	wire [16-1:0] node18349;
	wire [16-1:0] node18350;
	wire [16-1:0] node18353;
	wire [16-1:0] node18356;
	wire [16-1:0] node18357;
	wire [16-1:0] node18358;
	wire [16-1:0] node18360;
	wire [16-1:0] node18361;
	wire [16-1:0] node18363;
	wire [16-1:0] node18367;
	wire [16-1:0] node18368;
	wire [16-1:0] node18371;
	wire [16-1:0] node18374;
	wire [16-1:0] node18375;
	wire [16-1:0] node18376;
	wire [16-1:0] node18378;
	wire [16-1:0] node18380;
	wire [16-1:0] node18385;
	wire [16-1:0] node18386;
	wire [16-1:0] node18387;
	wire [16-1:0] node18388;
	wire [16-1:0] node18389;
	wire [16-1:0] node18394;
	wire [16-1:0] node18395;
	wire [16-1:0] node18396;
	wire [16-1:0] node18399;
	wire [16-1:0] node18401;
	wire [16-1:0] node18404;
	wire [16-1:0] node18405;
	wire [16-1:0] node18409;
	wire [16-1:0] node18410;
	wire [16-1:0] node18411;
	wire [16-1:0] node18414;
	wire [16-1:0] node18415;
	wire [16-1:0] node18417;
	wire [16-1:0] node18420;
	wire [16-1:0] node18422;
	wire [16-1:0] node18425;
	wire [16-1:0] node18427;
	wire [16-1:0] node18428;
	wire [16-1:0] node18429;
	wire [16-1:0] node18433;
	wire [16-1:0] node18436;
	wire [16-1:0] node18437;
	wire [16-1:0] node18438;
	wire [16-1:0] node18439;
	wire [16-1:0] node18440;
	wire [16-1:0] node18441;
	wire [16-1:0] node18443;
	wire [16-1:0] node18448;
	wire [16-1:0] node18449;
	wire [16-1:0] node18450;
	wire [16-1:0] node18454;
	wire [16-1:0] node18455;
	wire [16-1:0] node18459;
	wire [16-1:0] node18460;
	wire [16-1:0] node18461;
	wire [16-1:0] node18462;
	wire [16-1:0] node18466;
	wire [16-1:0] node18468;
	wire [16-1:0] node18471;
	wire [16-1:0] node18472;
	wire [16-1:0] node18473;
	wire [16-1:0] node18478;
	wire [16-1:0] node18479;
	wire [16-1:0] node18480;
	wire [16-1:0] node18482;
	wire [16-1:0] node18483;
	wire [16-1:0] node18486;
	wire [16-1:0] node18489;
	wire [16-1:0] node18490;
	wire [16-1:0] node18491;
	wire [16-1:0] node18492;
	wire [16-1:0] node18497;
	wire [16-1:0] node18498;
	wire [16-1:0] node18499;
	wire [16-1:0] node18504;
	wire [16-1:0] node18505;
	wire [16-1:0] node18506;
	wire [16-1:0] node18507;
	wire [16-1:0] node18509;
	wire [16-1:0] node18514;
	wire [16-1:0] node18515;
	wire [16-1:0] node18518;
	wire [16-1:0] node18519;
	wire [16-1:0] node18521;
	wire [16-1:0] node18524;
	wire [16-1:0] node18527;
	wire [16-1:0] node18528;
	wire [16-1:0] node18529;
	wire [16-1:0] node18530;
	wire [16-1:0] node18531;
	wire [16-1:0] node18533;
	wire [16-1:0] node18534;
	wire [16-1:0] node18537;
	wire [16-1:0] node18538;
	wire [16-1:0] node18539;
	wire [16-1:0] node18540;
	wire [16-1:0] node18545;
	wire [16-1:0] node18548;
	wire [16-1:0] node18549;
	wire [16-1:0] node18551;
	wire [16-1:0] node18552;
	wire [16-1:0] node18554;
	wire [16-1:0] node18557;
	wire [16-1:0] node18559;
	wire [16-1:0] node18562;
	wire [16-1:0] node18563;
	wire [16-1:0] node18565;
	wire [16-1:0] node18569;
	wire [16-1:0] node18570;
	wire [16-1:0] node18571;
	wire [16-1:0] node18573;
	wire [16-1:0] node18576;
	wire [16-1:0] node18578;
	wire [16-1:0] node18579;
	wire [16-1:0] node18583;
	wire [16-1:0] node18584;
	wire [16-1:0] node18585;
	wire [16-1:0] node18587;
	wire [16-1:0] node18591;
	wire [16-1:0] node18593;
	wire [16-1:0] node18596;
	wire [16-1:0] node18597;
	wire [16-1:0] node18598;
	wire [16-1:0] node18599;
	wire [16-1:0] node18600;
	wire [16-1:0] node18603;
	wire [16-1:0] node18605;
	wire [16-1:0] node18608;
	wire [16-1:0] node18609;
	wire [16-1:0] node18610;
	wire [16-1:0] node18614;
	wire [16-1:0] node18615;
	wire [16-1:0] node18619;
	wire [16-1:0] node18620;
	wire [16-1:0] node18621;
	wire [16-1:0] node18622;
	wire [16-1:0] node18626;
	wire [16-1:0] node18628;
	wire [16-1:0] node18630;
	wire [16-1:0] node18632;
	wire [16-1:0] node18635;
	wire [16-1:0] node18636;
	wire [16-1:0] node18638;
	wire [16-1:0] node18641;
	wire [16-1:0] node18642;
	wire [16-1:0] node18646;
	wire [16-1:0] node18647;
	wire [16-1:0] node18648;
	wire [16-1:0] node18649;
	wire [16-1:0] node18651;
	wire [16-1:0] node18655;
	wire [16-1:0] node18656;
	wire [16-1:0] node18657;
	wire [16-1:0] node18660;
	wire [16-1:0] node18663;
	wire [16-1:0] node18665;
	wire [16-1:0] node18668;
	wire [16-1:0] node18669;
	wire [16-1:0] node18670;
	wire [16-1:0] node18673;
	wire [16-1:0] node18674;
	wire [16-1:0] node18677;
	wire [16-1:0] node18679;
	wire [16-1:0] node18682;
	wire [16-1:0] node18683;
	wire [16-1:0] node18685;
	wire [16-1:0] node18688;
	wire [16-1:0] node18691;
	wire [16-1:0] node18692;
	wire [16-1:0] node18693;
	wire [16-1:0] node18694;
	wire [16-1:0] node18695;
	wire [16-1:0] node18696;
	wire [16-1:0] node18697;
	wire [16-1:0] node18701;
	wire [16-1:0] node18702;
	wire [16-1:0] node18705;
	wire [16-1:0] node18707;
	wire [16-1:0] node18710;
	wire [16-1:0] node18711;
	wire [16-1:0] node18712;
	wire [16-1:0] node18714;
	wire [16-1:0] node18718;
	wire [16-1:0] node18720;
	wire [16-1:0] node18721;
	wire [16-1:0] node18725;
	wire [16-1:0] node18726;
	wire [16-1:0] node18727;
	wire [16-1:0] node18729;
	wire [16-1:0] node18733;
	wire [16-1:0] node18734;
	wire [16-1:0] node18735;
	wire [16-1:0] node18739;
	wire [16-1:0] node18740;
	wire [16-1:0] node18742;
	wire [16-1:0] node18745;
	wire [16-1:0] node18748;
	wire [16-1:0] node18749;
	wire [16-1:0] node18750;
	wire [16-1:0] node18752;
	wire [16-1:0] node18754;
	wire [16-1:0] node18757;
	wire [16-1:0] node18758;
	wire [16-1:0] node18760;
	wire [16-1:0] node18761;
	wire [16-1:0] node18765;
	wire [16-1:0] node18767;
	wire [16-1:0] node18770;
	wire [16-1:0] node18771;
	wire [16-1:0] node18772;
	wire [16-1:0] node18774;
	wire [16-1:0] node18779;
	wire [16-1:0] node18780;
	wire [16-1:0] node18781;
	wire [16-1:0] node18782;
	wire [16-1:0] node18784;
	wire [16-1:0] node18787;
	wire [16-1:0] node18788;
	wire [16-1:0] node18789;
	wire [16-1:0] node18791;
	wire [16-1:0] node18794;
	wire [16-1:0] node18797;
	wire [16-1:0] node18798;
	wire [16-1:0] node18802;
	wire [16-1:0] node18803;
	wire [16-1:0] node18804;
	wire [16-1:0] node18806;
	wire [16-1:0] node18809;
	wire [16-1:0] node18810;
	wire [16-1:0] node18813;
	wire [16-1:0] node18816;
	wire [16-1:0] node18817;
	wire [16-1:0] node18819;
	wire [16-1:0] node18820;
	wire [16-1:0] node18825;
	wire [16-1:0] node18826;
	wire [16-1:0] node18827;
	wire [16-1:0] node18828;
	wire [16-1:0] node18831;
	wire [16-1:0] node18832;
	wire [16-1:0] node18836;
	wire [16-1:0] node18837;
	wire [16-1:0] node18839;
	wire [16-1:0] node18842;
	wire [16-1:0] node18844;
	wire [16-1:0] node18846;
	wire [16-1:0] node18849;
	wire [16-1:0] node18850;
	wire [16-1:0] node18852;
	wire [16-1:0] node18853;
	wire [16-1:0] node18856;
	wire [16-1:0] node18859;
	wire [16-1:0] node18860;
	wire [16-1:0] node18862;
	wire [16-1:0] node18866;
	wire [16-1:0] node18867;
	wire [16-1:0] node18868;
	wire [16-1:0] node18869;
	wire [16-1:0] node18870;
	wire [16-1:0] node18871;
	wire [16-1:0] node18872;
	wire [16-1:0] node18873;
	wire [16-1:0] node18874;
	wire [16-1:0] node18875;
	wire [16-1:0] node18877;
	wire [16-1:0] node18881;
	wire [16-1:0] node18884;
	wire [16-1:0] node18886;
	wire [16-1:0] node18889;
	wire [16-1:0] node18890;
	wire [16-1:0] node18893;
	wire [16-1:0] node18894;
	wire [16-1:0] node18895;
	wire [16-1:0] node18899;
	wire [16-1:0] node18902;
	wire [16-1:0] node18903;
	wire [16-1:0] node18904;
	wire [16-1:0] node18905;
	wire [16-1:0] node18908;
	wire [16-1:0] node18909;
	wire [16-1:0] node18913;
	wire [16-1:0] node18915;
	wire [16-1:0] node18918;
	wire [16-1:0] node18919;
	wire [16-1:0] node18920;
	wire [16-1:0] node18923;
	wire [16-1:0] node18925;
	wire [16-1:0] node18926;
	wire [16-1:0] node18931;
	wire [16-1:0] node18932;
	wire [16-1:0] node18933;
	wire [16-1:0] node18935;
	wire [16-1:0] node18936;
	wire [16-1:0] node18940;
	wire [16-1:0] node18942;
	wire [16-1:0] node18943;
	wire [16-1:0] node18947;
	wire [16-1:0] node18948;
	wire [16-1:0] node18949;
	wire [16-1:0] node18950;
	wire [16-1:0] node18954;
	wire [16-1:0] node18955;
	wire [16-1:0] node18956;
	wire [16-1:0] node18961;
	wire [16-1:0] node18962;
	wire [16-1:0] node18964;
	wire [16-1:0] node18967;
	wire [16-1:0] node18970;
	wire [16-1:0] node18971;
	wire [16-1:0] node18972;
	wire [16-1:0] node18973;
	wire [16-1:0] node18975;
	wire [16-1:0] node18976;
	wire [16-1:0] node18979;
	wire [16-1:0] node18982;
	wire [16-1:0] node18983;
	wire [16-1:0] node18984;
	wire [16-1:0] node18988;
	wire [16-1:0] node18990;
	wire [16-1:0] node18993;
	wire [16-1:0] node18994;
	wire [16-1:0] node18996;
	wire [16-1:0] node18997;
	wire [16-1:0] node19001;
	wire [16-1:0] node19002;
	wire [16-1:0] node19003;
	wire [16-1:0] node19004;
	wire [16-1:0] node19006;
	wire [16-1:0] node19011;
	wire [16-1:0] node19013;
	wire [16-1:0] node19016;
	wire [16-1:0] node19017;
	wire [16-1:0] node19018;
	wire [16-1:0] node19021;
	wire [16-1:0] node19022;
	wire [16-1:0] node19023;
	wire [16-1:0] node19028;
	wire [16-1:0] node19029;
	wire [16-1:0] node19030;
	wire [16-1:0] node19031;
	wire [16-1:0] node19035;
	wire [16-1:0] node19036;
	wire [16-1:0] node19039;
	wire [16-1:0] node19040;
	wire [16-1:0] node19044;
	wire [16-1:0] node19045;
	wire [16-1:0] node19047;
	wire [16-1:0] node19050;
	wire [16-1:0] node19051;
	wire [16-1:0] node19053;
	wire [16-1:0] node19057;
	wire [16-1:0] node19058;
	wire [16-1:0] node19059;
	wire [16-1:0] node19060;
	wire [16-1:0] node19061;
	wire [16-1:0] node19062;
	wire [16-1:0] node19063;
	wire [16-1:0] node19066;
	wire [16-1:0] node19070;
	wire [16-1:0] node19071;
	wire [16-1:0] node19072;
	wire [16-1:0] node19075;
	wire [16-1:0] node19079;
	wire [16-1:0] node19080;
	wire [16-1:0] node19081;
	wire [16-1:0] node19082;
	wire [16-1:0] node19084;
	wire [16-1:0] node19087;
	wire [16-1:0] node19088;
	wire [16-1:0] node19091;
	wire [16-1:0] node19092;
	wire [16-1:0] node19096;
	wire [16-1:0] node19099;
	wire [16-1:0] node19101;
	wire [16-1:0] node19102;
	wire [16-1:0] node19105;
	wire [16-1:0] node19107;
	wire [16-1:0] node19110;
	wire [16-1:0] node19111;
	wire [16-1:0] node19112;
	wire [16-1:0] node19113;
	wire [16-1:0] node19115;
	wire [16-1:0] node19116;
	wire [16-1:0] node19121;
	wire [16-1:0] node19122;
	wire [16-1:0] node19123;
	wire [16-1:0] node19124;
	wire [16-1:0] node19126;
	wire [16-1:0] node19130;
	wire [16-1:0] node19131;
	wire [16-1:0] node19135;
	wire [16-1:0] node19136;
	wire [16-1:0] node19140;
	wire [16-1:0] node19141;
	wire [16-1:0] node19142;
	wire [16-1:0] node19145;
	wire [16-1:0] node19148;
	wire [16-1:0] node19149;
	wire [16-1:0] node19150;
	wire [16-1:0] node19153;
	wire [16-1:0] node19156;
	wire [16-1:0] node19157;
	wire [16-1:0] node19160;
	wire [16-1:0] node19163;
	wire [16-1:0] node19164;
	wire [16-1:0] node19165;
	wire [16-1:0] node19166;
	wire [16-1:0] node19168;
	wire [16-1:0] node19169;
	wire [16-1:0] node19172;
	wire [16-1:0] node19175;
	wire [16-1:0] node19176;
	wire [16-1:0] node19178;
	wire [16-1:0] node19179;
	wire [16-1:0] node19183;
	wire [16-1:0] node19184;
	wire [16-1:0] node19188;
	wire [16-1:0] node19189;
	wire [16-1:0] node19190;
	wire [16-1:0] node19194;
	wire [16-1:0] node19195;
	wire [16-1:0] node19197;
	wire [16-1:0] node19200;
	wire [16-1:0] node19203;
	wire [16-1:0] node19204;
	wire [16-1:0] node19205;
	wire [16-1:0] node19206;
	wire [16-1:0] node19207;
	wire [16-1:0] node19209;
	wire [16-1:0] node19212;
	wire [16-1:0] node19213;
	wire [16-1:0] node19217;
	wire [16-1:0] node19220;
	wire [16-1:0] node19221;
	wire [16-1:0] node19222;
	wire [16-1:0] node19225;
	wire [16-1:0] node19228;
	wire [16-1:0] node19230;
	wire [16-1:0] node19233;
	wire [16-1:0] node19234;
	wire [16-1:0] node19235;
	wire [16-1:0] node19237;
	wire [16-1:0] node19239;
	wire [16-1:0] node19243;
	wire [16-1:0] node19244;
	wire [16-1:0] node19248;
	wire [16-1:0] node19249;
	wire [16-1:0] node19250;
	wire [16-1:0] node19251;
	wire [16-1:0] node19252;
	wire [16-1:0] node19253;
	wire [16-1:0] node19254;
	wire [16-1:0] node19255;
	wire [16-1:0] node19260;
	wire [16-1:0] node19261;
	wire [16-1:0] node19263;
	wire [16-1:0] node19267;
	wire [16-1:0] node19268;
	wire [16-1:0] node19270;
	wire [16-1:0] node19273;
	wire [16-1:0] node19275;
	wire [16-1:0] node19276;
	wire [16-1:0] node19280;
	wire [16-1:0] node19281;
	wire [16-1:0] node19282;
	wire [16-1:0] node19283;
	wire [16-1:0] node19284;
	wire [16-1:0] node19285;
	wire [16-1:0] node19289;
	wire [16-1:0] node19292;
	wire [16-1:0] node19293;
	wire [16-1:0] node19296;
	wire [16-1:0] node19299;
	wire [16-1:0] node19300;
	wire [16-1:0] node19301;
	wire [16-1:0] node19304;
	wire [16-1:0] node19307;
	wire [16-1:0] node19309;
	wire [16-1:0] node19312;
	wire [16-1:0] node19313;
	wire [16-1:0] node19314;
	wire [16-1:0] node19315;
	wire [16-1:0] node19319;
	wire [16-1:0] node19320;
	wire [16-1:0] node19324;
	wire [16-1:0] node19325;
	wire [16-1:0] node19326;
	wire [16-1:0] node19328;
	wire [16-1:0] node19331;
	wire [16-1:0] node19334;
	wire [16-1:0] node19336;
	wire [16-1:0] node19337;
	wire [16-1:0] node19341;
	wire [16-1:0] node19342;
	wire [16-1:0] node19343;
	wire [16-1:0] node19344;
	wire [16-1:0] node19345;
	wire [16-1:0] node19346;
	wire [16-1:0] node19349;
	wire [16-1:0] node19351;
	wire [16-1:0] node19354;
	wire [16-1:0] node19355;
	wire [16-1:0] node19359;
	wire [16-1:0] node19360;
	wire [16-1:0] node19361;
	wire [16-1:0] node19365;
	wire [16-1:0] node19367;
	wire [16-1:0] node19370;
	wire [16-1:0] node19371;
	wire [16-1:0] node19372;
	wire [16-1:0] node19373;
	wire [16-1:0] node19377;
	wire [16-1:0] node19378;
	wire [16-1:0] node19379;
	wire [16-1:0] node19383;
	wire [16-1:0] node19386;
	wire [16-1:0] node19387;
	wire [16-1:0] node19389;
	wire [16-1:0] node19392;
	wire [16-1:0] node19395;
	wire [16-1:0] node19396;
	wire [16-1:0] node19397;
	wire [16-1:0] node19398;
	wire [16-1:0] node19401;
	wire [16-1:0] node19403;
	wire [16-1:0] node19404;
	wire [16-1:0] node19408;
	wire [16-1:0] node19409;
	wire [16-1:0] node19412;
	wire [16-1:0] node19413;
	wire [16-1:0] node19415;
	wire [16-1:0] node19416;
	wire [16-1:0] node19420;
	wire [16-1:0] node19421;
	wire [16-1:0] node19422;
	wire [16-1:0] node19427;
	wire [16-1:0] node19428;
	wire [16-1:0] node19429;
	wire [16-1:0] node19431;
	wire [16-1:0] node19435;
	wire [16-1:0] node19436;
	wire [16-1:0] node19438;
	wire [16-1:0] node19440;
	wire [16-1:0] node19443;
	wire [16-1:0] node19444;
	wire [16-1:0] node19447;
	wire [16-1:0] node19448;
	wire [16-1:0] node19450;
	wire [16-1:0] node19454;
	wire [16-1:0] node19455;
	wire [16-1:0] node19456;
	wire [16-1:0] node19457;
	wire [16-1:0] node19458;
	wire [16-1:0] node19459;
	wire [16-1:0] node19460;
	wire [16-1:0] node19462;
	wire [16-1:0] node19463;
	wire [16-1:0] node19468;
	wire [16-1:0] node19469;
	wire [16-1:0] node19473;
	wire [16-1:0] node19474;
	wire [16-1:0] node19475;
	wire [16-1:0] node19479;
	wire [16-1:0] node19480;
	wire [16-1:0] node19483;
	wire [16-1:0] node19486;
	wire [16-1:0] node19487;
	wire [16-1:0] node19490;
	wire [16-1:0] node19491;
	wire [16-1:0] node19492;
	wire [16-1:0] node19494;
	wire [16-1:0] node19495;
	wire [16-1:0] node19499;
	wire [16-1:0] node19501;
	wire [16-1:0] node19505;
	wire [16-1:0] node19506;
	wire [16-1:0] node19507;
	wire [16-1:0] node19509;
	wire [16-1:0] node19510;
	wire [16-1:0] node19514;
	wire [16-1:0] node19515;
	wire [16-1:0] node19517;
	wire [16-1:0] node19520;
	wire [16-1:0] node19523;
	wire [16-1:0] node19524;
	wire [16-1:0] node19525;
	wire [16-1:0] node19529;
	wire [16-1:0] node19530;
	wire [16-1:0] node19531;
	wire [16-1:0] node19532;
	wire [16-1:0] node19536;
	wire [16-1:0] node19539;
	wire [16-1:0] node19541;
	wire [16-1:0] node19543;
	wire [16-1:0] node19546;
	wire [16-1:0] node19547;
	wire [16-1:0] node19548;
	wire [16-1:0] node19549;
	wire [16-1:0] node19550;
	wire [16-1:0] node19552;
	wire [16-1:0] node19555;
	wire [16-1:0] node19556;
	wire [16-1:0] node19559;
	wire [16-1:0] node19562;
	wire [16-1:0] node19564;
	wire [16-1:0] node19565;
	wire [16-1:0] node19569;
	wire [16-1:0] node19570;
	wire [16-1:0] node19571;
	wire [16-1:0] node19572;
	wire [16-1:0] node19576;
	wire [16-1:0] node19577;
	wire [16-1:0] node19581;
	wire [16-1:0] node19582;
	wire [16-1:0] node19583;
	wire [16-1:0] node19585;
	wire [16-1:0] node19586;
	wire [16-1:0] node19590;
	wire [16-1:0] node19593;
	wire [16-1:0] node19596;
	wire [16-1:0] node19597;
	wire [16-1:0] node19598;
	wire [16-1:0] node19599;
	wire [16-1:0] node19600;
	wire [16-1:0] node19605;
	wire [16-1:0] node19606;
	wire [16-1:0] node19607;
	wire [16-1:0] node19612;
	wire [16-1:0] node19613;
	wire [16-1:0] node19614;
	wire [16-1:0] node19615;
	wire [16-1:0] node19619;
	wire [16-1:0] node19621;
	wire [16-1:0] node19623;
	wire [16-1:0] node19626;
	wire [16-1:0] node19628;
	wire [16-1:0] node19629;
	wire [16-1:0] node19630;
	wire [16-1:0] node19632;
	wire [16-1:0] node19636;
	wire [16-1:0] node19638;
	wire [16-1:0] node19639;
	wire [16-1:0] node19643;
	wire [16-1:0] node19644;
	wire [16-1:0] node19645;
	wire [16-1:0] node19646;
	wire [16-1:0] node19647;
	wire [16-1:0] node19648;
	wire [16-1:0] node19649;
	wire [16-1:0] node19650;
	wire [16-1:0] node19651;
	wire [16-1:0] node19652;
	wire [16-1:0] node19655;
	wire [16-1:0] node19658;
	wire [16-1:0] node19659;
	wire [16-1:0] node19660;
	wire [16-1:0] node19662;
	wire [16-1:0] node19667;
	wire [16-1:0] node19668;
	wire [16-1:0] node19670;
	wire [16-1:0] node19672;
	wire [16-1:0] node19675;
	wire [16-1:0] node19678;
	wire [16-1:0] node19679;
	wire [16-1:0] node19680;
	wire [16-1:0] node19681;
	wire [16-1:0] node19685;
	wire [16-1:0] node19686;
	wire [16-1:0] node19688;
	wire [16-1:0] node19689;
	wire [16-1:0] node19694;
	wire [16-1:0] node19695;
	wire [16-1:0] node19696;
	wire [16-1:0] node19699;
	wire [16-1:0] node19703;
	wire [16-1:0] node19704;
	wire [16-1:0] node19705;
	wire [16-1:0] node19706;
	wire [16-1:0] node19707;
	wire [16-1:0] node19711;
	wire [16-1:0] node19714;
	wire [16-1:0] node19716;
	wire [16-1:0] node19719;
	wire [16-1:0] node19720;
	wire [16-1:0] node19721;
	wire [16-1:0] node19723;
	wire [16-1:0] node19725;
	wire [16-1:0] node19728;
	wire [16-1:0] node19731;
	wire [16-1:0] node19733;
	wire [16-1:0] node19734;
	wire [16-1:0] node19738;
	wire [16-1:0] node19739;
	wire [16-1:0] node19740;
	wire [16-1:0] node19741;
	wire [16-1:0] node19742;
	wire [16-1:0] node19743;
	wire [16-1:0] node19744;
	wire [16-1:0] node19749;
	wire [16-1:0] node19750;
	wire [16-1:0] node19754;
	wire [16-1:0] node19755;
	wire [16-1:0] node19756;
	wire [16-1:0] node19759;
	wire [16-1:0] node19762;
	wire [16-1:0] node19764;
	wire [16-1:0] node19765;
	wire [16-1:0] node19767;
	wire [16-1:0] node19771;
	wire [16-1:0] node19772;
	wire [16-1:0] node19775;
	wire [16-1:0] node19776;
	wire [16-1:0] node19777;
	wire [16-1:0] node19780;
	wire [16-1:0] node19783;
	wire [16-1:0] node19784;
	wire [16-1:0] node19785;
	wire [16-1:0] node19790;
	wire [16-1:0] node19791;
	wire [16-1:0] node19792;
	wire [16-1:0] node19793;
	wire [16-1:0] node19797;
	wire [16-1:0] node19798;
	wire [16-1:0] node19800;
	wire [16-1:0] node19803;
	wire [16-1:0] node19804;
	wire [16-1:0] node19805;
	wire [16-1:0] node19809;
	wire [16-1:0] node19812;
	wire [16-1:0] node19813;
	wire [16-1:0] node19814;
	wire [16-1:0] node19817;
	wire [16-1:0] node19818;
	wire [16-1:0] node19822;
	wire [16-1:0] node19823;
	wire [16-1:0] node19826;
	wire [16-1:0] node19828;
	wire [16-1:0] node19831;
	wire [16-1:0] node19832;
	wire [16-1:0] node19833;
	wire [16-1:0] node19834;
	wire [16-1:0] node19835;
	wire [16-1:0] node19836;
	wire [16-1:0] node19837;
	wire [16-1:0] node19838;
	wire [16-1:0] node19839;
	wire [16-1:0] node19845;
	wire [16-1:0] node19846;
	wire [16-1:0] node19849;
	wire [16-1:0] node19852;
	wire [16-1:0] node19853;
	wire [16-1:0] node19854;
	wire [16-1:0] node19857;
	wire [16-1:0] node19861;
	wire [16-1:0] node19862;
	wire [16-1:0] node19863;
	wire [16-1:0] node19864;
	wire [16-1:0] node19867;
	wire [16-1:0] node19870;
	wire [16-1:0] node19871;
	wire [16-1:0] node19875;
	wire [16-1:0] node19876;
	wire [16-1:0] node19879;
	wire [16-1:0] node19882;
	wire [16-1:0] node19883;
	wire [16-1:0] node19884;
	wire [16-1:0] node19885;
	wire [16-1:0] node19886;
	wire [16-1:0] node19890;
	wire [16-1:0] node19891;
	wire [16-1:0] node19894;
	wire [16-1:0] node19896;
	wire [16-1:0] node19899;
	wire [16-1:0] node19900;
	wire [16-1:0] node19904;
	wire [16-1:0] node19905;
	wire [16-1:0] node19907;
	wire [16-1:0] node19908;
	wire [16-1:0] node19912;
	wire [16-1:0] node19913;
	wire [16-1:0] node19915;
	wire [16-1:0] node19917;
	wire [16-1:0] node19918;
	wire [16-1:0] node19923;
	wire [16-1:0] node19924;
	wire [16-1:0] node19925;
	wire [16-1:0] node19926;
	wire [16-1:0] node19927;
	wire [16-1:0] node19928;
	wire [16-1:0] node19933;
	wire [16-1:0] node19934;
	wire [16-1:0] node19935;
	wire [16-1:0] node19938;
	wire [16-1:0] node19941;
	wire [16-1:0] node19942;
	wire [16-1:0] node19944;
	wire [16-1:0] node19947;
	wire [16-1:0] node19948;
	wire [16-1:0] node19949;
	wire [16-1:0] node19954;
	wire [16-1:0] node19955;
	wire [16-1:0] node19956;
	wire [16-1:0] node19958;
	wire [16-1:0] node19962;
	wire [16-1:0] node19964;
	wire [16-1:0] node19966;
	wire [16-1:0] node19969;
	wire [16-1:0] node19970;
	wire [16-1:0] node19971;
	wire [16-1:0] node19972;
	wire [16-1:0] node19973;
	wire [16-1:0] node19978;
	wire [16-1:0] node19979;
	wire [16-1:0] node19980;
	wire [16-1:0] node19984;
	wire [16-1:0] node19985;
	wire [16-1:0] node19989;
	wire [16-1:0] node19990;
	wire [16-1:0] node19991;
	wire [16-1:0] node19992;
	wire [16-1:0] node19996;
	wire [16-1:0] node19999;
	wire [16-1:0] node20000;
	wire [16-1:0] node20002;
	wire [16-1:0] node20003;
	wire [16-1:0] node20005;
	wire [16-1:0] node20009;
	wire [16-1:0] node20010;
	wire [16-1:0] node20013;
	wire [16-1:0] node20016;
	wire [16-1:0] node20017;
	wire [16-1:0] node20018;
	wire [16-1:0] node20019;
	wire [16-1:0] node20020;
	wire [16-1:0] node20021;
	wire [16-1:0] node20022;
	wire [16-1:0] node20024;
	wire [16-1:0] node20026;
	wire [16-1:0] node20028;
	wire [16-1:0] node20031;
	wire [16-1:0] node20033;
	wire [16-1:0] node20034;
	wire [16-1:0] node20038;
	wire [16-1:0] node20039;
	wire [16-1:0] node20041;
	wire [16-1:0] node20044;
	wire [16-1:0] node20046;
	wire [16-1:0] node20049;
	wire [16-1:0] node20050;
	wire [16-1:0] node20051;
	wire [16-1:0] node20055;
	wire [16-1:0] node20058;
	wire [16-1:0] node20059;
	wire [16-1:0] node20060;
	wire [16-1:0] node20062;
	wire [16-1:0] node20063;
	wire [16-1:0] node20067;
	wire [16-1:0] node20068;
	wire [16-1:0] node20069;
	wire [16-1:0] node20071;
	wire [16-1:0] node20076;
	wire [16-1:0] node20077;
	wire [16-1:0] node20078;
	wire [16-1:0] node20082;
	wire [16-1:0] node20083;
	wire [16-1:0] node20084;
	wire [16-1:0] node20088;
	wire [16-1:0] node20090;
	wire [16-1:0] node20092;
	wire [16-1:0] node20095;
	wire [16-1:0] node20096;
	wire [16-1:0] node20097;
	wire [16-1:0] node20098;
	wire [16-1:0] node20099;
	wire [16-1:0] node20100;
	wire [16-1:0] node20104;
	wire [16-1:0] node20107;
	wire [16-1:0] node20109;
	wire [16-1:0] node20111;
	wire [16-1:0] node20114;
	wire [16-1:0] node20115;
	wire [16-1:0] node20116;
	wire [16-1:0] node20117;
	wire [16-1:0] node20118;
	wire [16-1:0] node20122;
	wire [16-1:0] node20126;
	wire [16-1:0] node20127;
	wire [16-1:0] node20129;
	wire [16-1:0] node20132;
	wire [16-1:0] node20133;
	wire [16-1:0] node20137;
	wire [16-1:0] node20138;
	wire [16-1:0] node20139;
	wire [16-1:0] node20140;
	wire [16-1:0] node20141;
	wire [16-1:0] node20144;
	wire [16-1:0] node20147;
	wire [16-1:0] node20149;
	wire [16-1:0] node20152;
	wire [16-1:0] node20153;
	wire [16-1:0] node20155;
	wire [16-1:0] node20158;
	wire [16-1:0] node20159;
	wire [16-1:0] node20163;
	wire [16-1:0] node20164;
	wire [16-1:0] node20167;
	wire [16-1:0] node20168;
	wire [16-1:0] node20169;
	wire [16-1:0] node20171;
	wire [16-1:0] node20176;
	wire [16-1:0] node20177;
	wire [16-1:0] node20178;
	wire [16-1:0] node20179;
	wire [16-1:0] node20180;
	wire [16-1:0] node20181;
	wire [16-1:0] node20183;
	wire [16-1:0] node20186;
	wire [16-1:0] node20187;
	wire [16-1:0] node20191;
	wire [16-1:0] node20193;
	wire [16-1:0] node20194;
	wire [16-1:0] node20195;
	wire [16-1:0] node20197;
	wire [16-1:0] node20202;
	wire [16-1:0] node20203;
	wire [16-1:0] node20204;
	wire [16-1:0] node20205;
	wire [16-1:0] node20209;
	wire [16-1:0] node20210;
	wire [16-1:0] node20213;
	wire [16-1:0] node20216;
	wire [16-1:0] node20217;
	wire [16-1:0] node20219;
	wire [16-1:0] node20220;
	wire [16-1:0] node20221;
	wire [16-1:0] node20226;
	wire [16-1:0] node20228;
	wire [16-1:0] node20231;
	wire [16-1:0] node20232;
	wire [16-1:0] node20233;
	wire [16-1:0] node20235;
	wire [16-1:0] node20237;
	wire [16-1:0] node20240;
	wire [16-1:0] node20241;
	wire [16-1:0] node20242;
	wire [16-1:0] node20246;
	wire [16-1:0] node20247;
	wire [16-1:0] node20251;
	wire [16-1:0] node20252;
	wire [16-1:0] node20253;
	wire [16-1:0] node20255;
	wire [16-1:0] node20259;
	wire [16-1:0] node20260;
	wire [16-1:0] node20261;
	wire [16-1:0] node20262;
	wire [16-1:0] node20266;
	wire [16-1:0] node20269;
	wire [16-1:0] node20271;
	wire [16-1:0] node20274;
	wire [16-1:0] node20275;
	wire [16-1:0] node20276;
	wire [16-1:0] node20277;
	wire [16-1:0] node20278;
	wire [16-1:0] node20279;
	wire [16-1:0] node20283;
	wire [16-1:0] node20284;
	wire [16-1:0] node20288;
	wire [16-1:0] node20290;
	wire [16-1:0] node20293;
	wire [16-1:0] node20294;
	wire [16-1:0] node20295;
	wire [16-1:0] node20297;
	wire [16-1:0] node20298;
	wire [16-1:0] node20303;
	wire [16-1:0] node20304;
	wire [16-1:0] node20306;
	wire [16-1:0] node20309;
	wire [16-1:0] node20312;
	wire [16-1:0] node20313;
	wire [16-1:0] node20314;
	wire [16-1:0] node20315;
	wire [16-1:0] node20316;
	wire [16-1:0] node20319;
	wire [16-1:0] node20323;
	wire [16-1:0] node20324;
	wire [16-1:0] node20325;
	wire [16-1:0] node20328;
	wire [16-1:0] node20331;
	wire [16-1:0] node20332;
	wire [16-1:0] node20335;
	wire [16-1:0] node20337;
	wire [16-1:0] node20340;
	wire [16-1:0] node20341;
	wire [16-1:0] node20342;
	wire [16-1:0] node20343;
	wire [16-1:0] node20347;
	wire [16-1:0] node20348;
	wire [16-1:0] node20351;
	wire [16-1:0] node20352;
	wire [16-1:0] node20356;
	wire [16-1:0] node20357;
	wire [16-1:0] node20359;
	wire [16-1:0] node20360;
	wire [16-1:0] node20364;
	wire [16-1:0] node20366;
	wire [16-1:0] node20368;
	wire [16-1:0] node20370;
	wire [16-1:0] node20373;
	wire [16-1:0] node20374;
	wire [16-1:0] node20375;
	wire [16-1:0] node20376;
	wire [16-1:0] node20377;
	wire [16-1:0] node20378;
	wire [16-1:0] node20379;
	wire [16-1:0] node20380;
	wire [16-1:0] node20382;
	wire [16-1:0] node20383;
	wire [16-1:0] node20388;
	wire [16-1:0] node20389;
	wire [16-1:0] node20390;
	wire [16-1:0] node20391;
	wire [16-1:0] node20395;
	wire [16-1:0] node20399;
	wire [16-1:0] node20400;
	wire [16-1:0] node20401;
	wire [16-1:0] node20403;
	wire [16-1:0] node20405;
	wire [16-1:0] node20406;
	wire [16-1:0] node20411;
	wire [16-1:0] node20413;
	wire [16-1:0] node20414;
	wire [16-1:0] node20416;
	wire [16-1:0] node20419;
	wire [16-1:0] node20422;
	wire [16-1:0] node20423;
	wire [16-1:0] node20424;
	wire [16-1:0] node20426;
	wire [16-1:0] node20427;
	wire [16-1:0] node20431;
	wire [16-1:0] node20432;
	wire [16-1:0] node20434;
	wire [16-1:0] node20436;
	wire [16-1:0] node20437;
	wire [16-1:0] node20442;
	wire [16-1:0] node20443;
	wire [16-1:0] node20444;
	wire [16-1:0] node20447;
	wire [16-1:0] node20448;
	wire [16-1:0] node20452;
	wire [16-1:0] node20453;
	wire [16-1:0] node20456;
	wire [16-1:0] node20458;
	wire [16-1:0] node20459;
	wire [16-1:0] node20461;
	wire [16-1:0] node20464;
	wire [16-1:0] node20467;
	wire [16-1:0] node20468;
	wire [16-1:0] node20469;
	wire [16-1:0] node20470;
	wire [16-1:0] node20472;
	wire [16-1:0] node20473;
	wire [16-1:0] node20477;
	wire [16-1:0] node20478;
	wire [16-1:0] node20479;
	wire [16-1:0] node20482;
	wire [16-1:0] node20485;
	wire [16-1:0] node20488;
	wire [16-1:0] node20489;
	wire [16-1:0] node20490;
	wire [16-1:0] node20491;
	wire [16-1:0] node20494;
	wire [16-1:0] node20495;
	wire [16-1:0] node20499;
	wire [16-1:0] node20500;
	wire [16-1:0] node20501;
	wire [16-1:0] node20505;
	wire [16-1:0] node20507;
	wire [16-1:0] node20510;
	wire [16-1:0] node20511;
	wire [16-1:0] node20514;
	wire [16-1:0] node20517;
	wire [16-1:0] node20518;
	wire [16-1:0] node20519;
	wire [16-1:0] node20520;
	wire [16-1:0] node20522;
	wire [16-1:0] node20525;
	wire [16-1:0] node20527;
	wire [16-1:0] node20530;
	wire [16-1:0] node20531;
	wire [16-1:0] node20532;
	wire [16-1:0] node20535;
	wire [16-1:0] node20539;
	wire [16-1:0] node20540;
	wire [16-1:0] node20541;
	wire [16-1:0] node20543;
	wire [16-1:0] node20546;
	wire [16-1:0] node20547;
	wire [16-1:0] node20548;
	wire [16-1:0] node20553;
	wire [16-1:0] node20554;
	wire [16-1:0] node20556;
	wire [16-1:0] node20559;
	wire [16-1:0] node20560;
	wire [16-1:0] node20561;
	wire [16-1:0] node20565;
	wire [16-1:0] node20568;
	wire [16-1:0] node20569;
	wire [16-1:0] node20570;
	wire [16-1:0] node20571;
	wire [16-1:0] node20572;
	wire [16-1:0] node20573;
	wire [16-1:0] node20575;
	wire [16-1:0] node20579;
	wire [16-1:0] node20580;
	wire [16-1:0] node20582;
	wire [16-1:0] node20585;
	wire [16-1:0] node20586;
	wire [16-1:0] node20587;
	wire [16-1:0] node20592;
	wire [16-1:0] node20593;
	wire [16-1:0] node20594;
	wire [16-1:0] node20595;
	wire [16-1:0] node20598;
	wire [16-1:0] node20600;
	wire [16-1:0] node20601;
	wire [16-1:0] node20605;
	wire [16-1:0] node20606;
	wire [16-1:0] node20607;
	wire [16-1:0] node20612;
	wire [16-1:0] node20613;
	wire [16-1:0] node20615;
	wire [16-1:0] node20616;
	wire [16-1:0] node20618;
	wire [16-1:0] node20622;
	wire [16-1:0] node20623;
	wire [16-1:0] node20627;
	wire [16-1:0] node20628;
	wire [16-1:0] node20629;
	wire [16-1:0] node20630;
	wire [16-1:0] node20631;
	wire [16-1:0] node20633;
	wire [16-1:0] node20638;
	wire [16-1:0] node20639;
	wire [16-1:0] node20641;
	wire [16-1:0] node20644;
	wire [16-1:0] node20647;
	wire [16-1:0] node20648;
	wire [16-1:0] node20649;
	wire [16-1:0] node20651;
	wire [16-1:0] node20653;
	wire [16-1:0] node20654;
	wire [16-1:0] node20658;
	wire [16-1:0] node20659;
	wire [16-1:0] node20663;
	wire [16-1:0] node20664;
	wire [16-1:0] node20665;
	wire [16-1:0] node20666;
	wire [16-1:0] node20671;
	wire [16-1:0] node20674;
	wire [16-1:0] node20675;
	wire [16-1:0] node20676;
	wire [16-1:0] node20677;
	wire [16-1:0] node20678;
	wire [16-1:0] node20680;
	wire [16-1:0] node20683;
	wire [16-1:0] node20684;
	wire [16-1:0] node20685;
	wire [16-1:0] node20690;
	wire [16-1:0] node20691;
	wire [16-1:0] node20692;
	wire [16-1:0] node20696;
	wire [16-1:0] node20697;
	wire [16-1:0] node20698;
	wire [16-1:0] node20703;
	wire [16-1:0] node20704;
	wire [16-1:0] node20705;
	wire [16-1:0] node20707;
	wire [16-1:0] node20710;
	wire [16-1:0] node20713;
	wire [16-1:0] node20714;
	wire [16-1:0] node20715;
	wire [16-1:0] node20716;
	wire [16-1:0] node20720;
	wire [16-1:0] node20723;
	wire [16-1:0] node20724;
	wire [16-1:0] node20727;
	wire [16-1:0] node20730;
	wire [16-1:0] node20731;
	wire [16-1:0] node20732;
	wire [16-1:0] node20733;
	wire [16-1:0] node20735;
	wire [16-1:0] node20739;
	wire [16-1:0] node20740;
	wire [16-1:0] node20741;
	wire [16-1:0] node20745;
	wire [16-1:0] node20747;
	wire [16-1:0] node20750;
	wire [16-1:0] node20751;
	wire [16-1:0] node20752;
	wire [16-1:0] node20754;
	wire [16-1:0] node20755;
	wire [16-1:0] node20760;
	wire [16-1:0] node20761;
	wire [16-1:0] node20764;
	wire [16-1:0] node20767;
	wire [16-1:0] node20768;
	wire [16-1:0] node20769;
	wire [16-1:0] node20770;
	wire [16-1:0] node20771;
	wire [16-1:0] node20772;
	wire [16-1:0] node20773;
	wire [16-1:0] node20777;
	wire [16-1:0] node20778;
	wire [16-1:0] node20780;
	wire [16-1:0] node20782;
	wire [16-1:0] node20785;
	wire [16-1:0] node20786;
	wire [16-1:0] node20788;
	wire [16-1:0] node20789;
	wire [16-1:0] node20794;
	wire [16-1:0] node20795;
	wire [16-1:0] node20797;
	wire [16-1:0] node20798;
	wire [16-1:0] node20802;
	wire [16-1:0] node20803;
	wire [16-1:0] node20805;
	wire [16-1:0] node20808;
	wire [16-1:0] node20810;
	wire [16-1:0] node20811;
	wire [16-1:0] node20815;
	wire [16-1:0] node20816;
	wire [16-1:0] node20817;
	wire [16-1:0] node20819;
	wire [16-1:0] node20820;
	wire [16-1:0] node20824;
	wire [16-1:0] node20825;
	wire [16-1:0] node20827;
	wire [16-1:0] node20828;
	wire [16-1:0] node20829;
	wire [16-1:0] node20835;
	wire [16-1:0] node20836;
	wire [16-1:0] node20837;
	wire [16-1:0] node20840;
	wire [16-1:0] node20841;
	wire [16-1:0] node20844;
	wire [16-1:0] node20847;
	wire [16-1:0] node20849;
	wire [16-1:0] node20850;
	wire [16-1:0] node20853;
	wire [16-1:0] node20854;
	wire [16-1:0] node20857;
	wire [16-1:0] node20858;
	wire [16-1:0] node20862;
	wire [16-1:0] node20863;
	wire [16-1:0] node20864;
	wire [16-1:0] node20865;
	wire [16-1:0] node20866;
	wire [16-1:0] node20869;
	wire [16-1:0] node20872;
	wire [16-1:0] node20873;
	wire [16-1:0] node20874;
	wire [16-1:0] node20877;
	wire [16-1:0] node20881;
	wire [16-1:0] node20882;
	wire [16-1:0] node20884;
	wire [16-1:0] node20885;
	wire [16-1:0] node20887;
	wire [16-1:0] node20891;
	wire [16-1:0] node20892;
	wire [16-1:0] node20893;
	wire [16-1:0] node20895;
	wire [16-1:0] node20900;
	wire [16-1:0] node20901;
	wire [16-1:0] node20902;
	wire [16-1:0] node20903;
	wire [16-1:0] node20906;
	wire [16-1:0] node20907;
	wire [16-1:0] node20909;
	wire [16-1:0] node20913;
	wire [16-1:0] node20914;
	wire [16-1:0] node20915;
	wire [16-1:0] node20917;
	wire [16-1:0] node20922;
	wire [16-1:0] node20923;
	wire [16-1:0] node20924;
	wire [16-1:0] node20926;
	wire [16-1:0] node20928;
	wire [16-1:0] node20929;
	wire [16-1:0] node20934;
	wire [16-1:0] node20935;
	wire [16-1:0] node20936;
	wire [16-1:0] node20939;
	wire [16-1:0] node20941;
	wire [16-1:0] node20944;
	wire [16-1:0] node20945;
	wire [16-1:0] node20949;
	wire [16-1:0] node20950;
	wire [16-1:0] node20951;
	wire [16-1:0] node20952;
	wire [16-1:0] node20953;
	wire [16-1:0] node20955;
	wire [16-1:0] node20958;
	wire [16-1:0] node20959;
	wire [16-1:0] node20962;
	wire [16-1:0] node20963;
	wire [16-1:0] node20967;
	wire [16-1:0] node20968;
	wire [16-1:0] node20969;
	wire [16-1:0] node20971;
	wire [16-1:0] node20973;
	wire [16-1:0] node20977;
	wire [16-1:0] node20978;
	wire [16-1:0] node20980;
	wire [16-1:0] node20981;
	wire [16-1:0] node20986;
	wire [16-1:0] node20987;
	wire [16-1:0] node20988;
	wire [16-1:0] node20989;
	wire [16-1:0] node20991;
	wire [16-1:0] node20993;
	wire [16-1:0] node20996;
	wire [16-1:0] node20997;
	wire [16-1:0] node20999;
	wire [16-1:0] node21002;
	wire [16-1:0] node21005;
	wire [16-1:0] node21007;
	wire [16-1:0] node21009;
	wire [16-1:0] node21010;
	wire [16-1:0] node21014;
	wire [16-1:0] node21015;
	wire [16-1:0] node21017;
	wire [16-1:0] node21018;
	wire [16-1:0] node21019;
	wire [16-1:0] node21024;
	wire [16-1:0] node21025;
	wire [16-1:0] node21027;
	wire [16-1:0] node21030;
	wire [16-1:0] node21033;
	wire [16-1:0] node21034;
	wire [16-1:0] node21035;
	wire [16-1:0] node21036;
	wire [16-1:0] node21038;
	wire [16-1:0] node21039;
	wire [16-1:0] node21043;
	wire [16-1:0] node21045;
	wire [16-1:0] node21048;
	wire [16-1:0] node21049;
	wire [16-1:0] node21050;
	wire [16-1:0] node21051;
	wire [16-1:0] node21054;
	wire [16-1:0] node21057;
	wire [16-1:0] node21059;
	wire [16-1:0] node21062;
	wire [16-1:0] node21063;
	wire [16-1:0] node21064;
	wire [16-1:0] node21067;
	wire [16-1:0] node21068;
	wire [16-1:0] node21070;
	wire [16-1:0] node21074;
	wire [16-1:0] node21077;
	wire [16-1:0] node21078;
	wire [16-1:0] node21079;
	wire [16-1:0] node21080;
	wire [16-1:0] node21082;
	wire [16-1:0] node21085;
	wire [16-1:0] node21087;
	wire [16-1:0] node21088;
	wire [16-1:0] node21090;
	wire [16-1:0] node21094;
	wire [16-1:0] node21095;
	wire [16-1:0] node21097;
	wire [16-1:0] node21100;
	wire [16-1:0] node21101;
	wire [16-1:0] node21102;
	wire [16-1:0] node21107;
	wire [16-1:0] node21108;
	wire [16-1:0] node21109;
	wire [16-1:0] node21110;
	wire [16-1:0] node21113;
	wire [16-1:0] node21116;
	wire [16-1:0] node21117;
	wire [16-1:0] node21118;
	wire [16-1:0] node21123;
	wire [16-1:0] node21124;
	wire [16-1:0] node21127;
	wire [16-1:0] node21129;
	wire [16-1:0] node21132;
	wire [16-1:0] node21133;
	wire [16-1:0] node21134;
	wire [16-1:0] node21135;
	wire [16-1:0] node21136;
	wire [16-1:0] node21137;
	wire [16-1:0] node21138;
	wire [16-1:0] node21139;
	wire [16-1:0] node21140;
	wire [16-1:0] node21142;
	wire [16-1:0] node21144;
	wire [16-1:0] node21145;
	wire [16-1:0] node21146;
	wire [16-1:0] node21151;
	wire [16-1:0] node21152;
	wire [16-1:0] node21153;
	wire [16-1:0] node21156;
	wire [16-1:0] node21159;
	wire [16-1:0] node21160;
	wire [16-1:0] node21164;
	wire [16-1:0] node21165;
	wire [16-1:0] node21166;
	wire [16-1:0] node21168;
	wire [16-1:0] node21172;
	wire [16-1:0] node21173;
	wire [16-1:0] node21174;
	wire [16-1:0] node21177;
	wire [16-1:0] node21179;
	wire [16-1:0] node21183;
	wire [16-1:0] node21184;
	wire [16-1:0] node21186;
	wire [16-1:0] node21187;
	wire [16-1:0] node21188;
	wire [16-1:0] node21189;
	wire [16-1:0] node21193;
	wire [16-1:0] node21196;
	wire [16-1:0] node21197;
	wire [16-1:0] node21199;
	wire [16-1:0] node21202;
	wire [16-1:0] node21205;
	wire [16-1:0] node21206;
	wire [16-1:0] node21207;
	wire [16-1:0] node21208;
	wire [16-1:0] node21213;
	wire [16-1:0] node21215;
	wire [16-1:0] node21216;
	wire [16-1:0] node21219;
	wire [16-1:0] node21222;
	wire [16-1:0] node21223;
	wire [16-1:0] node21224;
	wire [16-1:0] node21225;
	wire [16-1:0] node21226;
	wire [16-1:0] node21227;
	wire [16-1:0] node21232;
	wire [16-1:0] node21233;
	wire [16-1:0] node21236;
	wire [16-1:0] node21237;
	wire [16-1:0] node21239;
	wire [16-1:0] node21242;
	wire [16-1:0] node21244;
	wire [16-1:0] node21247;
	wire [16-1:0] node21248;
	wire [16-1:0] node21249;
	wire [16-1:0] node21251;
	wire [16-1:0] node21255;
	wire [16-1:0] node21256;
	wire [16-1:0] node21259;
	wire [16-1:0] node21261;
	wire [16-1:0] node21263;
	wire [16-1:0] node21266;
	wire [16-1:0] node21267;
	wire [16-1:0] node21268;
	wire [16-1:0] node21269;
	wire [16-1:0] node21271;
	wire [16-1:0] node21272;
	wire [16-1:0] node21276;
	wire [16-1:0] node21278;
	wire [16-1:0] node21280;
	wire [16-1:0] node21283;
	wire [16-1:0] node21285;
	wire [16-1:0] node21287;
	wire [16-1:0] node21288;
	wire [16-1:0] node21292;
	wire [16-1:0] node21293;
	wire [16-1:0] node21294;
	wire [16-1:0] node21296;
	wire [16-1:0] node21299;
	wire [16-1:0] node21300;
	wire [16-1:0] node21304;
	wire [16-1:0] node21305;
	wire [16-1:0] node21306;
	wire [16-1:0] node21309;
	wire [16-1:0] node21313;
	wire [16-1:0] node21314;
	wire [16-1:0] node21315;
	wire [16-1:0] node21316;
	wire [16-1:0] node21317;
	wire [16-1:0] node21318;
	wire [16-1:0] node21319;
	wire [16-1:0] node21323;
	wire [16-1:0] node21324;
	wire [16-1:0] node21325;
	wire [16-1:0] node21330;
	wire [16-1:0] node21331;
	wire [16-1:0] node21333;
	wire [16-1:0] node21334;
	wire [16-1:0] node21336;
	wire [16-1:0] node21341;
	wire [16-1:0] node21342;
	wire [16-1:0] node21343;
	wire [16-1:0] node21345;
	wire [16-1:0] node21349;
	wire [16-1:0] node21350;
	wire [16-1:0] node21351;
	wire [16-1:0] node21352;
	wire [16-1:0] node21356;
	wire [16-1:0] node21358;
	wire [16-1:0] node21361;
	wire [16-1:0] node21363;
	wire [16-1:0] node21366;
	wire [16-1:0] node21367;
	wire [16-1:0] node21368;
	wire [16-1:0] node21369;
	wire [16-1:0] node21370;
	wire [16-1:0] node21374;
	wire [16-1:0] node21376;
	wire [16-1:0] node21377;
	wire [16-1:0] node21381;
	wire [16-1:0] node21382;
	wire [16-1:0] node21384;
	wire [16-1:0] node21385;
	wire [16-1:0] node21388;
	wire [16-1:0] node21389;
	wire [16-1:0] node21393;
	wire [16-1:0] node21394;
	wire [16-1:0] node21398;
	wire [16-1:0] node21399;
	wire [16-1:0] node21400;
	wire [16-1:0] node21401;
	wire [16-1:0] node21404;
	wire [16-1:0] node21407;
	wire [16-1:0] node21408;
	wire [16-1:0] node21410;
	wire [16-1:0] node21413;
	wire [16-1:0] node21416;
	wire [16-1:0] node21417;
	wire [16-1:0] node21418;
	wire [16-1:0] node21421;
	wire [16-1:0] node21423;
	wire [16-1:0] node21426;
	wire [16-1:0] node21429;
	wire [16-1:0] node21430;
	wire [16-1:0] node21431;
	wire [16-1:0] node21432;
	wire [16-1:0] node21435;
	wire [16-1:0] node21436;
	wire [16-1:0] node21437;
	wire [16-1:0] node21441;
	wire [16-1:0] node21443;
	wire [16-1:0] node21444;
	wire [16-1:0] node21448;
	wire [16-1:0] node21449;
	wire [16-1:0] node21450;
	wire [16-1:0] node21451;
	wire [16-1:0] node21456;
	wire [16-1:0] node21457;
	wire [16-1:0] node21459;
	wire [16-1:0] node21462;
	wire [16-1:0] node21465;
	wire [16-1:0] node21466;
	wire [16-1:0] node21467;
	wire [16-1:0] node21468;
	wire [16-1:0] node21469;
	wire [16-1:0] node21472;
	wire [16-1:0] node21475;
	wire [16-1:0] node21478;
	wire [16-1:0] node21479;
	wire [16-1:0] node21480;
	wire [16-1:0] node21484;
	wire [16-1:0] node21487;
	wire [16-1:0] node21488;
	wire [16-1:0] node21489;
	wire [16-1:0] node21491;
	wire [16-1:0] node21492;
	wire [16-1:0] node21495;
	wire [16-1:0] node21499;
	wire [16-1:0] node21501;
	wire [16-1:0] node21503;
	wire [16-1:0] node21506;
	wire [16-1:0] node21507;
	wire [16-1:0] node21508;
	wire [16-1:0] node21509;
	wire [16-1:0] node21510;
	wire [16-1:0] node21511;
	wire [16-1:0] node21513;
	wire [16-1:0] node21514;
	wire [16-1:0] node21518;
	wire [16-1:0] node21520;
	wire [16-1:0] node21522;
	wire [16-1:0] node21525;
	wire [16-1:0] node21526;
	wire [16-1:0] node21527;
	wire [16-1:0] node21528;
	wire [16-1:0] node21529;
	wire [16-1:0] node21533;
	wire [16-1:0] node21536;
	wire [16-1:0] node21537;
	wire [16-1:0] node21539;
	wire [16-1:0] node21540;
	wire [16-1:0] node21544;
	wire [16-1:0] node21547;
	wire [16-1:0] node21549;
	wire [16-1:0] node21550;
	wire [16-1:0] node21554;
	wire [16-1:0] node21555;
	wire [16-1:0] node21556;
	wire [16-1:0] node21558;
	wire [16-1:0] node21559;
	wire [16-1:0] node21561;
	wire [16-1:0] node21562;
	wire [16-1:0] node21566;
	wire [16-1:0] node21569;
	wire [16-1:0] node21570;
	wire [16-1:0] node21572;
	wire [16-1:0] node21576;
	wire [16-1:0] node21577;
	wire [16-1:0] node21578;
	wire [16-1:0] node21580;
	wire [16-1:0] node21583;
	wire [16-1:0] node21584;
	wire [16-1:0] node21587;
	wire [16-1:0] node21590;
	wire [16-1:0] node21592;
	wire [16-1:0] node21593;
	wire [16-1:0] node21597;
	wire [16-1:0] node21598;
	wire [16-1:0] node21599;
	wire [16-1:0] node21600;
	wire [16-1:0] node21601;
	wire [16-1:0] node21604;
	wire [16-1:0] node21607;
	wire [16-1:0] node21608;
	wire [16-1:0] node21609;
	wire [16-1:0] node21610;
	wire [16-1:0] node21615;
	wire [16-1:0] node21616;
	wire [16-1:0] node21620;
	wire [16-1:0] node21621;
	wire [16-1:0] node21622;
	wire [16-1:0] node21623;
	wire [16-1:0] node21625;
	wire [16-1:0] node21626;
	wire [16-1:0] node21631;
	wire [16-1:0] node21634;
	wire [16-1:0] node21635;
	wire [16-1:0] node21636;
	wire [16-1:0] node21639;
	wire [16-1:0] node21642;
	wire [16-1:0] node21644;
	wire [16-1:0] node21645;
	wire [16-1:0] node21649;
	wire [16-1:0] node21650;
	wire [16-1:0] node21651;
	wire [16-1:0] node21652;
	wire [16-1:0] node21653;
	wire [16-1:0] node21657;
	wire [16-1:0] node21658;
	wire [16-1:0] node21662;
	wire [16-1:0] node21663;
	wire [16-1:0] node21665;
	wire [16-1:0] node21667;
	wire [16-1:0] node21670;
	wire [16-1:0] node21671;
	wire [16-1:0] node21673;
	wire [16-1:0] node21676;
	wire [16-1:0] node21679;
	wire [16-1:0] node21680;
	wire [16-1:0] node21681;
	wire [16-1:0] node21682;
	wire [16-1:0] node21685;
	wire [16-1:0] node21688;
	wire [16-1:0] node21689;
	wire [16-1:0] node21692;
	wire [16-1:0] node21693;
	wire [16-1:0] node21697;
	wire [16-1:0] node21699;
	wire [16-1:0] node21700;
	wire [16-1:0] node21703;
	wire [16-1:0] node21704;
	wire [16-1:0] node21706;
	wire [16-1:0] node21710;
	wire [16-1:0] node21711;
	wire [16-1:0] node21712;
	wire [16-1:0] node21713;
	wire [16-1:0] node21714;
	wire [16-1:0] node21716;
	wire [16-1:0] node21717;
	wire [16-1:0] node21719;
	wire [16-1:0] node21720;
	wire [16-1:0] node21725;
	wire [16-1:0] node21726;
	wire [16-1:0] node21729;
	wire [16-1:0] node21730;
	wire [16-1:0] node21733;
	wire [16-1:0] node21736;
	wire [16-1:0] node21738;
	wire [16-1:0] node21739;
	wire [16-1:0] node21740;
	wire [16-1:0] node21743;
	wire [16-1:0] node21746;
	wire [16-1:0] node21747;
	wire [16-1:0] node21750;
	wire [16-1:0] node21753;
	wire [16-1:0] node21754;
	wire [16-1:0] node21755;
	wire [16-1:0] node21756;
	wire [16-1:0] node21757;
	wire [16-1:0] node21758;
	wire [16-1:0] node21760;
	wire [16-1:0] node21764;
	wire [16-1:0] node21767;
	wire [16-1:0] node21768;
	wire [16-1:0] node21771;
	wire [16-1:0] node21773;
	wire [16-1:0] node21776;
	wire [16-1:0] node21778;
	wire [16-1:0] node21779;
	wire [16-1:0] node21780;
	wire [16-1:0] node21783;
	wire [16-1:0] node21784;
	wire [16-1:0] node21788;
	wire [16-1:0] node21790;
	wire [16-1:0] node21793;
	wire [16-1:0] node21794;
	wire [16-1:0] node21795;
	wire [16-1:0] node21796;
	wire [16-1:0] node21799;
	wire [16-1:0] node21803;
	wire [16-1:0] node21804;
	wire [16-1:0] node21805;
	wire [16-1:0] node21808;
	wire [16-1:0] node21811;
	wire [16-1:0] node21812;
	wire [16-1:0] node21814;
	wire [16-1:0] node21817;
	wire [16-1:0] node21818;
	wire [16-1:0] node21822;
	wire [16-1:0] node21823;
	wire [16-1:0] node21824;
	wire [16-1:0] node21825;
	wire [16-1:0] node21826;
	wire [16-1:0] node21828;
	wire [16-1:0] node21829;
	wire [16-1:0] node21830;
	wire [16-1:0] node21835;
	wire [16-1:0] node21837;
	wire [16-1:0] node21840;
	wire [16-1:0] node21841;
	wire [16-1:0] node21843;
	wire [16-1:0] node21846;
	wire [16-1:0] node21847;
	wire [16-1:0] node21850;
	wire [16-1:0] node21851;
	wire [16-1:0] node21855;
	wire [16-1:0] node21856;
	wire [16-1:0] node21857;
	wire [16-1:0] node21859;
	wire [16-1:0] node21860;
	wire [16-1:0] node21863;
	wire [16-1:0] node21866;
	wire [16-1:0] node21867;
	wire [16-1:0] node21872;
	wire [16-1:0] node21873;
	wire [16-1:0] node21874;
	wire [16-1:0] node21875;
	wire [16-1:0] node21877;
	wire [16-1:0] node21881;
	wire [16-1:0] node21883;
	wire [16-1:0] node21885;
	wire [16-1:0] node21888;
	wire [16-1:0] node21889;
	wire [16-1:0] node21890;
	wire [16-1:0] node21891;
	wire [16-1:0] node21895;
	wire [16-1:0] node21896;
	wire [16-1:0] node21897;
	wire [16-1:0] node21901;
	wire [16-1:0] node21904;
	wire [16-1:0] node21905;
	wire [16-1:0] node21907;
	wire [16-1:0] node21910;
	wire [16-1:0] node21913;
	wire [16-1:0] node21914;
	wire [16-1:0] node21915;
	wire [16-1:0] node21916;
	wire [16-1:0] node21917;
	wire [16-1:0] node21918;
	wire [16-1:0] node21919;
	wire [16-1:0] node21920;
	wire [16-1:0] node21921;
	wire [16-1:0] node21923;
	wire [16-1:0] node21927;
	wire [16-1:0] node21929;
	wire [16-1:0] node21931;
	wire [16-1:0] node21934;
	wire [16-1:0] node21935;
	wire [16-1:0] node21938;
	wire [16-1:0] node21939;
	wire [16-1:0] node21943;
	wire [16-1:0] node21944;
	wire [16-1:0] node21945;
	wire [16-1:0] node21946;
	wire [16-1:0] node21949;
	wire [16-1:0] node21950;
	wire [16-1:0] node21952;
	wire [16-1:0] node21955;
	wire [16-1:0] node21956;
	wire [16-1:0] node21960;
	wire [16-1:0] node21961;
	wire [16-1:0] node21964;
	wire [16-1:0] node21967;
	wire [16-1:0] node21968;
	wire [16-1:0] node21970;
	wire [16-1:0] node21974;
	wire [16-1:0] node21975;
	wire [16-1:0] node21976;
	wire [16-1:0] node21977;
	wire [16-1:0] node21978;
	wire [16-1:0] node21981;
	wire [16-1:0] node21984;
	wire [16-1:0] node21985;
	wire [16-1:0] node21988;
	wire [16-1:0] node21990;
	wire [16-1:0] node21993;
	wire [16-1:0] node21994;
	wire [16-1:0] node21996;
	wire [16-1:0] node22000;
	wire [16-1:0] node22001;
	wire [16-1:0] node22003;
	wire [16-1:0] node22004;
	wire [16-1:0] node22005;
	wire [16-1:0] node22007;
	wire [16-1:0] node22011;
	wire [16-1:0] node22014;
	wire [16-1:0] node22016;
	wire [16-1:0] node22019;
	wire [16-1:0] node22020;
	wire [16-1:0] node22021;
	wire [16-1:0] node22022;
	wire [16-1:0] node22023;
	wire [16-1:0] node22024;
	wire [16-1:0] node22026;
	wire [16-1:0] node22030;
	wire [16-1:0] node22031;
	wire [16-1:0] node22033;
	wire [16-1:0] node22036;
	wire [16-1:0] node22039;
	wire [16-1:0] node22040;
	wire [16-1:0] node22041;
	wire [16-1:0] node22044;
	wire [16-1:0] node22047;
	wire [16-1:0] node22050;
	wire [16-1:0] node22051;
	wire [16-1:0] node22052;
	wire [16-1:0] node22054;
	wire [16-1:0] node22057;
	wire [16-1:0] node22058;
	wire [16-1:0] node22061;
	wire [16-1:0] node22064;
	wire [16-1:0] node22065;
	wire [16-1:0] node22066;
	wire [16-1:0] node22069;
	wire [16-1:0] node22072;
	wire [16-1:0] node22075;
	wire [16-1:0] node22076;
	wire [16-1:0] node22077;
	wire [16-1:0] node22078;
	wire [16-1:0] node22079;
	wire [16-1:0] node22082;
	wire [16-1:0] node22085;
	wire [16-1:0] node22087;
	wire [16-1:0] node22090;
	wire [16-1:0] node22091;
	wire [16-1:0] node22094;
	wire [16-1:0] node22095;
	wire [16-1:0] node22096;
	wire [16-1:0] node22100;
	wire [16-1:0] node22102;
	wire [16-1:0] node22103;
	wire [16-1:0] node22107;
	wire [16-1:0] node22108;
	wire [16-1:0] node22111;
	wire [16-1:0] node22112;
	wire [16-1:0] node22113;
	wire [16-1:0] node22114;
	wire [16-1:0] node22118;
	wire [16-1:0] node22119;
	wire [16-1:0] node22121;
	wire [16-1:0] node22125;
	wire [16-1:0] node22127;
	wire [16-1:0] node22130;
	wire [16-1:0] node22131;
	wire [16-1:0] node22132;
	wire [16-1:0] node22133;
	wire [16-1:0] node22134;
	wire [16-1:0] node22135;
	wire [16-1:0] node22137;
	wire [16-1:0] node22138;
	wire [16-1:0] node22142;
	wire [16-1:0] node22143;
	wire [16-1:0] node22147;
	wire [16-1:0] node22148;
	wire [16-1:0] node22150;
	wire [16-1:0] node22153;
	wire [16-1:0] node22154;
	wire [16-1:0] node22157;
	wire [16-1:0] node22160;
	wire [16-1:0] node22161;
	wire [16-1:0] node22162;
	wire [16-1:0] node22164;
	wire [16-1:0] node22165;
	wire [16-1:0] node22167;
	wire [16-1:0] node22171;
	wire [16-1:0] node22172;
	wire [16-1:0] node22173;
	wire [16-1:0] node22177;
	wire [16-1:0] node22179;
	wire [16-1:0] node22182;
	wire [16-1:0] node22183;
	wire [16-1:0] node22186;
	wire [16-1:0] node22187;
	wire [16-1:0] node22188;
	wire [16-1:0] node22190;
	wire [16-1:0] node22194;
	wire [16-1:0] node22197;
	wire [16-1:0] node22198;
	wire [16-1:0] node22199;
	wire [16-1:0] node22201;
	wire [16-1:0] node22204;
	wire [16-1:0] node22205;
	wire [16-1:0] node22206;
	wire [16-1:0] node22209;
	wire [16-1:0] node22210;
	wire [16-1:0] node22214;
	wire [16-1:0] node22215;
	wire [16-1:0] node22216;
	wire [16-1:0] node22218;
	wire [16-1:0] node22222;
	wire [16-1:0] node22225;
	wire [16-1:0] node22226;
	wire [16-1:0] node22229;
	wire [16-1:0] node22230;
	wire [16-1:0] node22232;
	wire [16-1:0] node22233;
	wire [16-1:0] node22238;
	wire [16-1:0] node22239;
	wire [16-1:0] node22240;
	wire [16-1:0] node22241;
	wire [16-1:0] node22242;
	wire [16-1:0] node22244;
	wire [16-1:0] node22246;
	wire [16-1:0] node22248;
	wire [16-1:0] node22251;
	wire [16-1:0] node22252;
	wire [16-1:0] node22255;
	wire [16-1:0] node22258;
	wire [16-1:0] node22259;
	wire [16-1:0] node22261;
	wire [16-1:0] node22264;
	wire [16-1:0] node22265;
	wire [16-1:0] node22268;
	wire [16-1:0] node22271;
	wire [16-1:0] node22272;
	wire [16-1:0] node22273;
	wire [16-1:0] node22277;
	wire [16-1:0] node22278;
	wire [16-1:0] node22280;
	wire [16-1:0] node22282;
	wire [16-1:0] node22285;
	wire [16-1:0] node22286;
	wire [16-1:0] node22289;
	wire [16-1:0] node22291;
	wire [16-1:0] node22294;
	wire [16-1:0] node22295;
	wire [16-1:0] node22296;
	wire [16-1:0] node22297;
	wire [16-1:0] node22300;
	wire [16-1:0] node22301;
	wire [16-1:0] node22305;
	wire [16-1:0] node22306;
	wire [16-1:0] node22308;
	wire [16-1:0] node22309;
	wire [16-1:0] node22313;
	wire [16-1:0] node22316;
	wire [16-1:0] node22317;
	wire [16-1:0] node22318;
	wire [16-1:0] node22320;
	wire [16-1:0] node22321;
	wire [16-1:0] node22324;
	wire [16-1:0] node22327;
	wire [16-1:0] node22329;
	wire [16-1:0] node22331;
	wire [16-1:0] node22334;
	wire [16-1:0] node22336;
	wire [16-1:0] node22337;
	wire [16-1:0] node22340;
	wire [16-1:0] node22341;
	wire [16-1:0] node22343;
	wire [16-1:0] node22347;
	wire [16-1:0] node22348;
	wire [16-1:0] node22349;
	wire [16-1:0] node22350;
	wire [16-1:0] node22351;
	wire [16-1:0] node22352;
	wire [16-1:0] node22353;
	wire [16-1:0] node22354;
	wire [16-1:0] node22358;
	wire [16-1:0] node22359;
	wire [16-1:0] node22361;
	wire [16-1:0] node22364;
	wire [16-1:0] node22365;
	wire [16-1:0] node22366;
	wire [16-1:0] node22371;
	wire [16-1:0] node22372;
	wire [16-1:0] node22374;
	wire [16-1:0] node22377;
	wire [16-1:0] node22378;
	wire [16-1:0] node22382;
	wire [16-1:0] node22383;
	wire [16-1:0] node22384;
	wire [16-1:0] node22385;
	wire [16-1:0] node22389;
	wire [16-1:0] node22390;
	wire [16-1:0] node22393;
	wire [16-1:0] node22394;
	wire [16-1:0] node22398;
	wire [16-1:0] node22399;
	wire [16-1:0] node22402;
	wire [16-1:0] node22403;
	wire [16-1:0] node22404;
	wire [16-1:0] node22408;
	wire [16-1:0] node22411;
	wire [16-1:0] node22412;
	wire [16-1:0] node22413;
	wire [16-1:0] node22414;
	wire [16-1:0] node22416;
	wire [16-1:0] node22419;
	wire [16-1:0] node22420;
	wire [16-1:0] node22421;
	wire [16-1:0] node22426;
	wire [16-1:0] node22427;
	wire [16-1:0] node22431;
	wire [16-1:0] node22432;
	wire [16-1:0] node22433;
	wire [16-1:0] node22434;
	wire [16-1:0] node22438;
	wire [16-1:0] node22439;
	wire [16-1:0] node22442;
	wire [16-1:0] node22445;
	wire [16-1:0] node22447;
	wire [16-1:0] node22448;
	wire [16-1:0] node22452;
	wire [16-1:0] node22453;
	wire [16-1:0] node22454;
	wire [16-1:0] node22455;
	wire [16-1:0] node22457;
	wire [16-1:0] node22458;
	wire [16-1:0] node22462;
	wire [16-1:0] node22463;
	wire [16-1:0] node22467;
	wire [16-1:0] node22468;
	wire [16-1:0] node22469;
	wire [16-1:0] node22471;
	wire [16-1:0] node22472;
	wire [16-1:0] node22476;
	wire [16-1:0] node22478;
	wire [16-1:0] node22480;
	wire [16-1:0] node22483;
	wire [16-1:0] node22486;
	wire [16-1:0] node22487;
	wire [16-1:0] node22488;
	wire [16-1:0] node22490;
	wire [16-1:0] node22491;
	wire [16-1:0] node22493;
	wire [16-1:0] node22496;
	wire [16-1:0] node22497;
	wire [16-1:0] node22501;
	wire [16-1:0] node22503;
	wire [16-1:0] node22504;
	wire [16-1:0] node22508;
	wire [16-1:0] node22509;
	wire [16-1:0] node22511;
	wire [16-1:0] node22512;
	wire [16-1:0] node22514;
	wire [16-1:0] node22515;
	wire [16-1:0] node22520;
	wire [16-1:0] node22521;
	wire [16-1:0] node22523;
	wire [16-1:0] node22526;
	wire [16-1:0] node22527;
	wire [16-1:0] node22528;
	wire [16-1:0] node22532;
	wire [16-1:0] node22535;
	wire [16-1:0] node22536;
	wire [16-1:0] node22537;
	wire [16-1:0] node22538;
	wire [16-1:0] node22539;
	wire [16-1:0] node22540;
	wire [16-1:0] node22543;
	wire [16-1:0] node22544;
	wire [16-1:0] node22545;
	wire [16-1:0] node22550;
	wire [16-1:0] node22551;
	wire [16-1:0] node22553;
	wire [16-1:0] node22555;
	wire [16-1:0] node22558;
	wire [16-1:0] node22559;
	wire [16-1:0] node22560;
	wire [16-1:0] node22562;
	wire [16-1:0] node22567;
	wire [16-1:0] node22568;
	wire [16-1:0] node22570;
	wire [16-1:0] node22571;
	wire [16-1:0] node22575;
	wire [16-1:0] node22576;
	wire [16-1:0] node22579;
	wire [16-1:0] node22581;
	wire [16-1:0] node22584;
	wire [16-1:0] node22585;
	wire [16-1:0] node22586;
	wire [16-1:0] node22587;
	wire [16-1:0] node22589;
	wire [16-1:0] node22591;
	wire [16-1:0] node22594;
	wire [16-1:0] node22595;
	wire [16-1:0] node22596;
	wire [16-1:0] node22600;
	wire [16-1:0] node22603;
	wire [16-1:0] node22605;
	wire [16-1:0] node22606;
	wire [16-1:0] node22610;
	wire [16-1:0] node22611;
	wire [16-1:0] node22613;
	wire [16-1:0] node22614;
	wire [16-1:0] node22618;
	wire [16-1:0] node22619;
	wire [16-1:0] node22621;
	wire [16-1:0] node22624;
	wire [16-1:0] node22625;
	wire [16-1:0] node22626;
	wire [16-1:0] node22630;
	wire [16-1:0] node22633;
	wire [16-1:0] node22634;
	wire [16-1:0] node22635;
	wire [16-1:0] node22636;
	wire [16-1:0] node22637;
	wire [16-1:0] node22638;
	wire [16-1:0] node22641;
	wire [16-1:0] node22644;
	wire [16-1:0] node22647;
	wire [16-1:0] node22649;
	wire [16-1:0] node22650;
	wire [16-1:0] node22652;
	wire [16-1:0] node22656;
	wire [16-1:0] node22657;
	wire [16-1:0] node22658;
	wire [16-1:0] node22660;
	wire [16-1:0] node22661;
	wire [16-1:0] node22665;
	wire [16-1:0] node22666;
	wire [16-1:0] node22668;
	wire [16-1:0] node22672;
	wire [16-1:0] node22673;
	wire [16-1:0] node22676;
	wire [16-1:0] node22677;
	wire [16-1:0] node22678;
	wire [16-1:0] node22680;
	wire [16-1:0] node22685;
	wire [16-1:0] node22686;
	wire [16-1:0] node22687;
	wire [16-1:0] node22688;
	wire [16-1:0] node22689;
	wire [16-1:0] node22691;
	wire [16-1:0] node22695;
	wire [16-1:0] node22697;
	wire [16-1:0] node22698;
	wire [16-1:0] node22700;
	wire [16-1:0] node22704;
	wire [16-1:0] node22706;
	wire [16-1:0] node22707;
	wire [16-1:0] node22711;
	wire [16-1:0] node22712;
	wire [16-1:0] node22713;
	wire [16-1:0] node22714;
	wire [16-1:0] node22717;
	wire [16-1:0] node22720;
	wire [16-1:0] node22722;
	wire [16-1:0] node22724;
	wire [16-1:0] node22725;
	wire [16-1:0] node22729;
	wire [16-1:0] node22731;
	wire [16-1:0] node22732;
	wire [16-1:0] node22734;
	wire [16-1:0] node22738;
	wire [16-1:0] node22739;
	wire [16-1:0] node22740;
	wire [16-1:0] node22741;
	wire [16-1:0] node22742;
	wire [16-1:0] node22743;
	wire [16-1:0] node22744;
	wire [16-1:0] node22745;
	wire [16-1:0] node22746;
	wire [16-1:0] node22747;
	wire [16-1:0] node22750;
	wire [16-1:0] node22753;
	wire [16-1:0] node22754;
	wire [16-1:0] node22757;
	wire [16-1:0] node22760;
	wire [16-1:0] node22761;
	wire [16-1:0] node22762;
	wire [16-1:0] node22763;
	wire [16-1:0] node22767;
	wire [16-1:0] node22769;
	wire [16-1:0] node22772;
	wire [16-1:0] node22774;
	wire [16-1:0] node22777;
	wire [16-1:0] node22778;
	wire [16-1:0] node22779;
	wire [16-1:0] node22780;
	wire [16-1:0] node22784;
	wire [16-1:0] node22785;
	wire [16-1:0] node22789;
	wire [16-1:0] node22790;
	wire [16-1:0] node22793;
	wire [16-1:0] node22795;
	wire [16-1:0] node22798;
	wire [16-1:0] node22799;
	wire [16-1:0] node22800;
	wire [16-1:0] node22801;
	wire [16-1:0] node22804;
	wire [16-1:0] node22807;
	wire [16-1:0] node22809;
	wire [16-1:0] node22812;
	wire [16-1:0] node22813;
	wire [16-1:0] node22814;
	wire [16-1:0] node22816;
	wire [16-1:0] node22819;
	wire [16-1:0] node22820;
	wire [16-1:0] node22824;
	wire [16-1:0] node22825;
	wire [16-1:0] node22827;
	wire [16-1:0] node22829;
	wire [16-1:0] node22832;
	wire [16-1:0] node22833;
	wire [16-1:0] node22837;
	wire [16-1:0] node22838;
	wire [16-1:0] node22839;
	wire [16-1:0] node22840;
	wire [16-1:0] node22841;
	wire [16-1:0] node22843;
	wire [16-1:0] node22844;
	wire [16-1:0] node22846;
	wire [16-1:0] node22850;
	wire [16-1:0] node22853;
	wire [16-1:0] node22856;
	wire [16-1:0] node22857;
	wire [16-1:0] node22858;
	wire [16-1:0] node22859;
	wire [16-1:0] node22863;
	wire [16-1:0] node22865;
	wire [16-1:0] node22868;
	wire [16-1:0] node22869;
	wire [16-1:0] node22871;
	wire [16-1:0] node22875;
	wire [16-1:0] node22876;
	wire [16-1:0] node22877;
	wire [16-1:0] node22878;
	wire [16-1:0] node22880;
	wire [16-1:0] node22884;
	wire [16-1:0] node22885;
	wire [16-1:0] node22886;
	wire [16-1:0] node22889;
	wire [16-1:0] node22893;
	wire [16-1:0] node22894;
	wire [16-1:0] node22895;
	wire [16-1:0] node22897;
	wire [16-1:0] node22900;
	wire [16-1:0] node22901;
	wire [16-1:0] node22905;
	wire [16-1:0] node22906;
	wire [16-1:0] node22907;
	wire [16-1:0] node22911;
	wire [16-1:0] node22913;
	wire [16-1:0] node22914;
	wire [16-1:0] node22918;
	wire [16-1:0] node22919;
	wire [16-1:0] node22920;
	wire [16-1:0] node22921;
	wire [16-1:0] node22922;
	wire [16-1:0] node22923;
	wire [16-1:0] node22926;
	wire [16-1:0] node22927;
	wire [16-1:0] node22930;
	wire [16-1:0] node22932;
	wire [16-1:0] node22935;
	wire [16-1:0] node22936;
	wire [16-1:0] node22937;
	wire [16-1:0] node22941;
	wire [16-1:0] node22944;
	wire [16-1:0] node22945;
	wire [16-1:0] node22946;
	wire [16-1:0] node22948;
	wire [16-1:0] node22952;
	wire [16-1:0] node22953;
	wire [16-1:0] node22955;
	wire [16-1:0] node22957;
	wire [16-1:0] node22961;
	wire [16-1:0] node22962;
	wire [16-1:0] node22963;
	wire [16-1:0] node22966;
	wire [16-1:0] node22967;
	wire [16-1:0] node22969;
	wire [16-1:0] node22971;
	wire [16-1:0] node22972;
	wire [16-1:0] node22976;
	wire [16-1:0] node22978;
	wire [16-1:0] node22981;
	wire [16-1:0] node22982;
	wire [16-1:0] node22983;
	wire [16-1:0] node22985;
	wire [16-1:0] node22988;
	wire [16-1:0] node22989;
	wire [16-1:0] node22991;
	wire [16-1:0] node22995;
	wire [16-1:0] node22996;
	wire [16-1:0] node22998;
	wire [16-1:0] node22999;
	wire [16-1:0] node23004;
	wire [16-1:0] node23005;
	wire [16-1:0] node23006;
	wire [16-1:0] node23007;
	wire [16-1:0] node23008;
	wire [16-1:0] node23011;
	wire [16-1:0] node23012;
	wire [16-1:0] node23014;
	wire [16-1:0] node23015;
	wire [16-1:0] node23020;
	wire [16-1:0] node23021;
	wire [16-1:0] node23024;
	wire [16-1:0] node23027;
	wire [16-1:0] node23028;
	wire [16-1:0] node23029;
	wire [16-1:0] node23031;
	wire [16-1:0] node23034;
	wire [16-1:0] node23035;
	wire [16-1:0] node23038;
	wire [16-1:0] node23041;
	wire [16-1:0] node23042;
	wire [16-1:0] node23044;
	wire [16-1:0] node23045;
	wire [16-1:0] node23050;
	wire [16-1:0] node23051;
	wire [16-1:0] node23053;
	wire [16-1:0] node23056;
	wire [16-1:0] node23057;
	wire [16-1:0] node23058;
	wire [16-1:0] node23060;
	wire [16-1:0] node23062;
	wire [16-1:0] node23065;
	wire [16-1:0] node23068;
	wire [16-1:0] node23069;
	wire [16-1:0] node23070;
	wire [16-1:0] node23074;
	wire [16-1:0] node23075;
	wire [16-1:0] node23077;
	wire [16-1:0] node23081;
	wire [16-1:0] node23082;
	wire [16-1:0] node23083;
	wire [16-1:0] node23084;
	wire [16-1:0] node23085;
	wire [16-1:0] node23086;
	wire [16-1:0] node23087;
	wire [16-1:0] node23088;
	wire [16-1:0] node23092;
	wire [16-1:0] node23093;
	wire [16-1:0] node23095;
	wire [16-1:0] node23099;
	wire [16-1:0] node23100;
	wire [16-1:0] node23101;
	wire [16-1:0] node23106;
	wire [16-1:0] node23107;
	wire [16-1:0] node23108;
	wire [16-1:0] node23109;
	wire [16-1:0] node23113;
	wire [16-1:0] node23116;
	wire [16-1:0] node23118;
	wire [16-1:0] node23119;
	wire [16-1:0] node23122;
	wire [16-1:0] node23125;
	wire [16-1:0] node23126;
	wire [16-1:0] node23127;
	wire [16-1:0] node23128;
	wire [16-1:0] node23129;
	wire [16-1:0] node23132;
	wire [16-1:0] node23134;
	wire [16-1:0] node23138;
	wire [16-1:0] node23141;
	wire [16-1:0] node23142;
	wire [16-1:0] node23143;
	wire [16-1:0] node23144;
	wire [16-1:0] node23147;
	wire [16-1:0] node23150;
	wire [16-1:0] node23151;
	wire [16-1:0] node23155;
	wire [16-1:0] node23156;
	wire [16-1:0] node23157;
	wire [16-1:0] node23159;
	wire [16-1:0] node23163;
	wire [16-1:0] node23164;
	wire [16-1:0] node23168;
	wire [16-1:0] node23169;
	wire [16-1:0] node23170;
	wire [16-1:0] node23171;
	wire [16-1:0] node23172;
	wire [16-1:0] node23174;
	wire [16-1:0] node23177;
	wire [16-1:0] node23178;
	wire [16-1:0] node23180;
	wire [16-1:0] node23184;
	wire [16-1:0] node23185;
	wire [16-1:0] node23187;
	wire [16-1:0] node23190;
	wire [16-1:0] node23193;
	wire [16-1:0] node23194;
	wire [16-1:0] node23195;
	wire [16-1:0] node23196;
	wire [16-1:0] node23199;
	wire [16-1:0] node23202;
	wire [16-1:0] node23203;
	wire [16-1:0] node23204;
	wire [16-1:0] node23209;
	wire [16-1:0] node23210;
	wire [16-1:0] node23212;
	wire [16-1:0] node23214;
	wire [16-1:0] node23217;
	wire [16-1:0] node23218;
	wire [16-1:0] node23222;
	wire [16-1:0] node23223;
	wire [16-1:0] node23224;
	wire [16-1:0] node23225;
	wire [16-1:0] node23227;
	wire [16-1:0] node23230;
	wire [16-1:0] node23231;
	wire [16-1:0] node23233;
	wire [16-1:0] node23236;
	wire [16-1:0] node23239;
	wire [16-1:0] node23240;
	wire [16-1:0] node23241;
	wire [16-1:0] node23245;
	wire [16-1:0] node23246;
	wire [16-1:0] node23248;
	wire [16-1:0] node23252;
	wire [16-1:0] node23253;
	wire [16-1:0] node23254;
	wire [16-1:0] node23255;
	wire [16-1:0] node23256;
	wire [16-1:0] node23261;
	wire [16-1:0] node23262;
	wire [16-1:0] node23266;
	wire [16-1:0] node23267;
	wire [16-1:0] node23268;
	wire [16-1:0] node23272;
	wire [16-1:0] node23274;
	wire [16-1:0] node23277;
	wire [16-1:0] node23278;
	wire [16-1:0] node23279;
	wire [16-1:0] node23280;
	wire [16-1:0] node23281;
	wire [16-1:0] node23282;
	wire [16-1:0] node23284;
	wire [16-1:0] node23288;
	wire [16-1:0] node23289;
	wire [16-1:0] node23291;
	wire [16-1:0] node23294;
	wire [16-1:0] node23297;
	wire [16-1:0] node23298;
	wire [16-1:0] node23299;
	wire [16-1:0] node23300;
	wire [16-1:0] node23302;
	wire [16-1:0] node23305;
	wire [16-1:0] node23306;
	wire [16-1:0] node23307;
	wire [16-1:0] node23312;
	wire [16-1:0] node23314;
	wire [16-1:0] node23316;
	wire [16-1:0] node23319;
	wire [16-1:0] node23321;
	wire [16-1:0] node23322;
	wire [16-1:0] node23324;
	wire [16-1:0] node23327;
	wire [16-1:0] node23329;
	wire [16-1:0] node23332;
	wire [16-1:0] node23333;
	wire [16-1:0] node23334;
	wire [16-1:0] node23335;
	wire [16-1:0] node23336;
	wire [16-1:0] node23339;
	wire [16-1:0] node23340;
	wire [16-1:0] node23342;
	wire [16-1:0] node23346;
	wire [16-1:0] node23347;
	wire [16-1:0] node23350;
	wire [16-1:0] node23353;
	wire [16-1:0] node23354;
	wire [16-1:0] node23356;
	wire [16-1:0] node23357;
	wire [16-1:0] node23359;
	wire [16-1:0] node23363;
	wire [16-1:0] node23364;
	wire [16-1:0] node23368;
	wire [16-1:0] node23369;
	wire [16-1:0] node23370;
	wire [16-1:0] node23372;
	wire [16-1:0] node23376;
	wire [16-1:0] node23377;
	wire [16-1:0] node23378;
	wire [16-1:0] node23379;
	wire [16-1:0] node23384;
	wire [16-1:0] node23385;
	wire [16-1:0] node23388;
	wire [16-1:0] node23389;
	wire [16-1:0] node23392;
	wire [16-1:0] node23394;
	wire [16-1:0] node23397;
	wire [16-1:0] node23398;
	wire [16-1:0] node23399;
	wire [16-1:0] node23400;
	wire [16-1:0] node23401;
	wire [16-1:0] node23404;
	wire [16-1:0] node23406;
	wire [16-1:0] node23408;
	wire [16-1:0] node23411;
	wire [16-1:0] node23412;
	wire [16-1:0] node23414;
	wire [16-1:0] node23415;
	wire [16-1:0] node23419;
	wire [16-1:0] node23421;
	wire [16-1:0] node23424;
	wire [16-1:0] node23425;
	wire [16-1:0] node23426;
	wire [16-1:0] node23428;
	wire [16-1:0] node23431;
	wire [16-1:0] node23432;
	wire [16-1:0] node23436;
	wire [16-1:0] node23437;
	wire [16-1:0] node23438;
	wire [16-1:0] node23441;
	wire [16-1:0] node23442;
	wire [16-1:0] node23444;
	wire [16-1:0] node23448;
	wire [16-1:0] node23450;
	wire [16-1:0] node23452;
	wire [16-1:0] node23455;
	wire [16-1:0] node23456;
	wire [16-1:0] node23457;
	wire [16-1:0] node23458;
	wire [16-1:0] node23461;
	wire [16-1:0] node23462;
	wire [16-1:0] node23466;
	wire [16-1:0] node23468;
	wire [16-1:0] node23469;
	wire [16-1:0] node23473;
	wire [16-1:0] node23474;
	wire [16-1:0] node23475;
	wire [16-1:0] node23478;
	wire [16-1:0] node23481;
	wire [16-1:0] node23482;
	wire [16-1:0] node23485;
	wire [16-1:0] node23487;
	wire [16-1:0] node23489;
	wire [16-1:0] node23490;
	wire [16-1:0] node23494;
	wire [16-1:0] node23495;
	wire [16-1:0] node23496;
	wire [16-1:0] node23497;
	wire [16-1:0] node23498;
	wire [16-1:0] node23499;
	wire [16-1:0] node23500;
	wire [16-1:0] node23501;
	wire [16-1:0] node23504;
	wire [16-1:0] node23505;
	wire [16-1:0] node23509;
	wire [16-1:0] node23511;
	wire [16-1:0] node23514;
	wire [16-1:0] node23515;
	wire [16-1:0] node23516;
	wire [16-1:0] node23518;
	wire [16-1:0] node23519;
	wire [16-1:0] node23523;
	wire [16-1:0] node23524;
	wire [16-1:0] node23528;
	wire [16-1:0] node23529;
	wire [16-1:0] node23530;
	wire [16-1:0] node23533;
	wire [16-1:0] node23535;
	wire [16-1:0] node23538;
	wire [16-1:0] node23541;
	wire [16-1:0] node23542;
	wire [16-1:0] node23543;
	wire [16-1:0] node23545;
	wire [16-1:0] node23548;
	wire [16-1:0] node23550;
	wire [16-1:0] node23551;
	wire [16-1:0] node23555;
	wire [16-1:0] node23556;
	wire [16-1:0] node23557;
	wire [16-1:0] node23558;
	wire [16-1:0] node23560;
	wire [16-1:0] node23565;
	wire [16-1:0] node23567;
	wire [16-1:0] node23568;
	wire [16-1:0] node23572;
	wire [16-1:0] node23573;
	wire [16-1:0] node23574;
	wire [16-1:0] node23575;
	wire [16-1:0] node23576;
	wire [16-1:0] node23577;
	wire [16-1:0] node23581;
	wire [16-1:0] node23582;
	wire [16-1:0] node23583;
	wire [16-1:0] node23586;
	wire [16-1:0] node23587;
	wire [16-1:0] node23591;
	wire [16-1:0] node23594;
	wire [16-1:0] node23595;
	wire [16-1:0] node23598;
	wire [16-1:0] node23599;
	wire [16-1:0] node23600;
	wire [16-1:0] node23602;
	wire [16-1:0] node23607;
	wire [16-1:0] node23608;
	wire [16-1:0] node23609;
	wire [16-1:0] node23612;
	wire [16-1:0] node23613;
	wire [16-1:0] node23615;
	wire [16-1:0] node23616;
	wire [16-1:0] node23620;
	wire [16-1:0] node23623;
	wire [16-1:0] node23624;
	wire [16-1:0] node23626;
	wire [16-1:0] node23629;
	wire [16-1:0] node23631;
	wire [16-1:0] node23632;
	wire [16-1:0] node23636;
	wire [16-1:0] node23637;
	wire [16-1:0] node23638;
	wire [16-1:0] node23639;
	wire [16-1:0] node23643;
	wire [16-1:0] node23644;
	wire [16-1:0] node23647;
	wire [16-1:0] node23649;
	wire [16-1:0] node23652;
	wire [16-1:0] node23653;
	wire [16-1:0] node23654;
	wire [16-1:0] node23655;
	wire [16-1:0] node23660;
	wire [16-1:0] node23662;
	wire [16-1:0] node23663;
	wire [16-1:0] node23666;
	wire [16-1:0] node23669;
	wire [16-1:0] node23670;
	wire [16-1:0] node23671;
	wire [16-1:0] node23672;
	wire [16-1:0] node23673;
	wire [16-1:0] node23674;
	wire [16-1:0] node23676;
	wire [16-1:0] node23678;
	wire [16-1:0] node23681;
	wire [16-1:0] node23683;
	wire [16-1:0] node23686;
	wire [16-1:0] node23687;
	wire [16-1:0] node23689;
	wire [16-1:0] node23693;
	wire [16-1:0] node23694;
	wire [16-1:0] node23695;
	wire [16-1:0] node23697;
	wire [16-1:0] node23701;
	wire [16-1:0] node23702;
	wire [16-1:0] node23704;
	wire [16-1:0] node23708;
	wire [16-1:0] node23709;
	wire [16-1:0] node23710;
	wire [16-1:0] node23711;
	wire [16-1:0] node23712;
	wire [16-1:0] node23716;
	wire [16-1:0] node23717;
	wire [16-1:0] node23719;
	wire [16-1:0] node23720;
	wire [16-1:0] node23725;
	wire [16-1:0] node23726;
	wire [16-1:0] node23727;
	wire [16-1:0] node23731;
	wire [16-1:0] node23733;
	wire [16-1:0] node23736;
	wire [16-1:0] node23737;
	wire [16-1:0] node23738;
	wire [16-1:0] node23739;
	wire [16-1:0] node23740;
	wire [16-1:0] node23744;
	wire [16-1:0] node23747;
	wire [16-1:0] node23748;
	wire [16-1:0] node23751;
	wire [16-1:0] node23753;
	wire [16-1:0] node23756;
	wire [16-1:0] node23757;
	wire [16-1:0] node23758;
	wire [16-1:0] node23761;
	wire [16-1:0] node23762;
	wire [16-1:0] node23767;
	wire [16-1:0] node23768;
	wire [16-1:0] node23769;
	wire [16-1:0] node23770;
	wire [16-1:0] node23771;
	wire [16-1:0] node23773;
	wire [16-1:0] node23774;
	wire [16-1:0] node23779;
	wire [16-1:0] node23780;
	wire [16-1:0] node23781;
	wire [16-1:0] node23784;
	wire [16-1:0] node23787;
	wire [16-1:0] node23789;
	wire [16-1:0] node23792;
	wire [16-1:0] node23793;
	wire [16-1:0] node23794;
	wire [16-1:0] node23795;
	wire [16-1:0] node23798;
	wire [16-1:0] node23799;
	wire [16-1:0] node23803;
	wire [16-1:0] node23804;
	wire [16-1:0] node23807;
	wire [16-1:0] node23809;
	wire [16-1:0] node23810;
	wire [16-1:0] node23814;
	wire [16-1:0] node23815;
	wire [16-1:0] node23817;
	wire [16-1:0] node23819;
	wire [16-1:0] node23820;
	wire [16-1:0] node23824;
	wire [16-1:0] node23825;
	wire [16-1:0] node23828;
	wire [16-1:0] node23829;
	wire [16-1:0] node23830;
	wire [16-1:0] node23835;
	wire [16-1:0] node23836;
	wire [16-1:0] node23837;
	wire [16-1:0] node23838;
	wire [16-1:0] node23842;
	wire [16-1:0] node23843;
	wire [16-1:0] node23847;
	wire [16-1:0] node23848;
	wire [16-1:0] node23849;
	wire [16-1:0] node23851;
	wire [16-1:0] node23854;
	wire [16-1:0] node23857;
	wire [16-1:0] node23858;
	wire [16-1:0] node23861;
	wire [16-1:0] node23862;
	wire [16-1:0] node23865;
	wire [16-1:0] node23866;
	wire [16-1:0] node23868;
	wire [16-1:0] node23871;
	wire [16-1:0] node23873;
	wire [16-1:0] node23876;
	wire [16-1:0] node23877;
	wire [16-1:0] node23878;
	wire [16-1:0] node23879;
	wire [16-1:0] node23880;
	wire [16-1:0] node23881;
	wire [16-1:0] node23882;
	wire [16-1:0] node23884;
	wire [16-1:0] node23885;
	wire [16-1:0] node23890;
	wire [16-1:0] node23893;
	wire [16-1:0] node23894;
	wire [16-1:0] node23895;
	wire [16-1:0] node23897;
	wire [16-1:0] node23900;
	wire [16-1:0] node23901;
	wire [16-1:0] node23904;
	wire [16-1:0] node23906;
	wire [16-1:0] node23907;
	wire [16-1:0] node23911;
	wire [16-1:0] node23913;
	wire [16-1:0] node23916;
	wire [16-1:0] node23917;
	wire [16-1:0] node23918;
	wire [16-1:0] node23919;
	wire [16-1:0] node23921;
	wire [16-1:0] node23922;
	wire [16-1:0] node23927;
	wire [16-1:0] node23928;
	wire [16-1:0] node23929;
	wire [16-1:0] node23933;
	wire [16-1:0] node23934;
	wire [16-1:0] node23938;
	wire [16-1:0] node23939;
	wire [16-1:0] node23940;
	wire [16-1:0] node23943;
	wire [16-1:0] node23946;
	wire [16-1:0] node23947;
	wire [16-1:0] node23949;
	wire [16-1:0] node23951;
	wire [16-1:0] node23955;
	wire [16-1:0] node23956;
	wire [16-1:0] node23957;
	wire [16-1:0] node23958;
	wire [16-1:0] node23960;
	wire [16-1:0] node23961;
	wire [16-1:0] node23962;
	wire [16-1:0] node23967;
	wire [16-1:0] node23968;
	wire [16-1:0] node23970;
	wire [16-1:0] node23974;
	wire [16-1:0] node23975;
	wire [16-1:0] node23976;
	wire [16-1:0] node23978;
	wire [16-1:0] node23982;
	wire [16-1:0] node23983;
	wire [16-1:0] node23984;
	wire [16-1:0] node23985;
	wire [16-1:0] node23987;
	wire [16-1:0] node23991;
	wire [16-1:0] node23994;
	wire [16-1:0] node23997;
	wire [16-1:0] node23998;
	wire [16-1:0] node23999;
	wire [16-1:0] node24000;
	wire [16-1:0] node24001;
	wire [16-1:0] node24005;
	wire [16-1:0] node24006;
	wire [16-1:0] node24008;
	wire [16-1:0] node24011;
	wire [16-1:0] node24014;
	wire [16-1:0] node24015;
	wire [16-1:0] node24016;
	wire [16-1:0] node24019;
	wire [16-1:0] node24022;
	wire [16-1:0] node24023;
	wire [16-1:0] node24025;
	wire [16-1:0] node24026;
	wire [16-1:0] node24031;
	wire [16-1:0] node24032;
	wire [16-1:0] node24033;
	wire [16-1:0] node24035;
	wire [16-1:0] node24038;
	wire [16-1:0] node24039;
	wire [16-1:0] node24041;
	wire [16-1:0] node24045;
	wire [16-1:0] node24046;
	wire [16-1:0] node24047;
	wire [16-1:0] node24050;
	wire [16-1:0] node24052;
	wire [16-1:0] node24053;
	wire [16-1:0] node24058;
	wire [16-1:0] node24059;
	wire [16-1:0] node24060;
	wire [16-1:0] node24061;
	wire [16-1:0] node24062;
	wire [16-1:0] node24063;
	wire [16-1:0] node24064;
	wire [16-1:0] node24065;
	wire [16-1:0] node24070;
	wire [16-1:0] node24073;
	wire [16-1:0] node24074;
	wire [16-1:0] node24077;
	wire [16-1:0] node24078;
	wire [16-1:0] node24082;
	wire [16-1:0] node24083;
	wire [16-1:0] node24084;
	wire [16-1:0] node24085;
	wire [16-1:0] node24086;
	wire [16-1:0] node24090;
	wire [16-1:0] node24092;
	wire [16-1:0] node24095;
	wire [16-1:0] node24097;
	wire [16-1:0] node24100;
	wire [16-1:0] node24101;
	wire [16-1:0] node24104;
	wire [16-1:0] node24105;
	wire [16-1:0] node24106;
	wire [16-1:0] node24110;
	wire [16-1:0] node24112;
	wire [16-1:0] node24115;
	wire [16-1:0] node24116;
	wire [16-1:0] node24117;
	wire [16-1:0] node24118;
	wire [16-1:0] node24120;
	wire [16-1:0] node24122;
	wire [16-1:0] node24125;
	wire [16-1:0] node24126;
	wire [16-1:0] node24130;
	wire [16-1:0] node24131;
	wire [16-1:0] node24133;
	wire [16-1:0] node24136;
	wire [16-1:0] node24138;
	wire [16-1:0] node24140;
	wire [16-1:0] node24143;
	wire [16-1:0] node24144;
	wire [16-1:0] node24145;
	wire [16-1:0] node24147;
	wire [16-1:0] node24150;
	wire [16-1:0] node24152;
	wire [16-1:0] node24155;
	wire [16-1:0] node24156;
	wire [16-1:0] node24157;
	wire [16-1:0] node24161;
	wire [16-1:0] node24162;
	wire [16-1:0] node24166;
	wire [16-1:0] node24167;
	wire [16-1:0] node24168;
	wire [16-1:0] node24169;
	wire [16-1:0] node24170;
	wire [16-1:0] node24171;
	wire [16-1:0] node24174;
	wire [16-1:0] node24177;
	wire [16-1:0] node24178;
	wire [16-1:0] node24179;
	wire [16-1:0] node24184;
	wire [16-1:0] node24186;
	wire [16-1:0] node24189;
	wire [16-1:0] node24190;
	wire [16-1:0] node24191;
	wire [16-1:0] node24193;
	wire [16-1:0] node24195;
	wire [16-1:0] node24198;
	wire [16-1:0] node24199;
	wire [16-1:0] node24203;
	wire [16-1:0] node24204;
	wire [16-1:0] node24205;
	wire [16-1:0] node24206;
	wire [16-1:0] node24210;
	wire [16-1:0] node24213;
	wire [16-1:0] node24214;
	wire [16-1:0] node24218;
	wire [16-1:0] node24219;
	wire [16-1:0] node24220;
	wire [16-1:0] node24221;
	wire [16-1:0] node24222;
	wire [16-1:0] node24223;
	wire [16-1:0] node24228;
	wire [16-1:0] node24229;
	wire [16-1:0] node24233;
	wire [16-1:0] node24234;
	wire [16-1:0] node24235;
	wire [16-1:0] node24238;
	wire [16-1:0] node24241;
	wire [16-1:0] node24242;
	wire [16-1:0] node24245;
	wire [16-1:0] node24248;
	wire [16-1:0] node24249;
	wire [16-1:0] node24250;
	wire [16-1:0] node24251;
	wire [16-1:0] node24254;
	wire [16-1:0] node24258;
	wire [16-1:0] node24259;
	wire [16-1:0] node24260;
	wire [16-1:0] node24263;
	wire [16-1:0] node24265;
	wire [16-1:0] node24268;
	wire [16-1:0] node24269;
	wire [16-1:0] node24271;
	wire [16-1:0] node24273;
	wire [16-1:0] node24276;
	wire [16-1:0] node24278;

	assign outp = (inp[7]) ? node11916 : node1;
		assign node1 = (inp[11]) ? node5877 : node2;
			assign node2 = (inp[3]) ? node2956 : node3;
				assign node3 = (inp[10]) ? node1479 : node4;
					assign node4 = (inp[9]) ? node758 : node5;
						assign node5 = (inp[8]) ? node421 : node6;
							assign node6 = (inp[5]) ? node212 : node7;
								assign node7 = (inp[15]) ? node107 : node8;
									assign node8 = (inp[2]) ? node62 : node9;
										assign node9 = (inp[1]) ? node39 : node10;
											assign node10 = (inp[6]) ? node28 : node11;
												assign node11 = (inp[14]) ? node19 : node12;
													assign node12 = (inp[12]) ? node16 : node13;
														assign node13 = (inp[4]) ? 16'b0011111111111111 : 16'b0111111111111111;
														assign node16 = (inp[0]) ? 16'b0000111111111111 : 16'b0011111111111111;
													assign node19 = (inp[4]) ? 16'b0001111111111111 : node20;
														assign node20 = (inp[13]) ? node22 : 16'b0011111111111111;
															assign node22 = (inp[12]) ? 16'b0001111111111111 : node23;
																assign node23 = (inp[0]) ? 16'b0001111111111111 : 16'b0011111111111111;
												assign node28 = (inp[0]) ? node34 : node29;
													assign node29 = (inp[13]) ? 16'b0001111111111111 : node30;
														assign node30 = (inp[4]) ? 16'b0000111111111111 : 16'b0001111111111111;
													assign node34 = (inp[14]) ? 16'b0000011111111111 : node35;
														assign node35 = (inp[12]) ? 16'b0000111111111111 : 16'b0011111111111111;
											assign node39 = (inp[0]) ? node51 : node40;
												assign node40 = (inp[12]) ? node48 : node41;
													assign node41 = (inp[14]) ? node45 : node42;
														assign node42 = (inp[6]) ? 16'b0001111111111111 : 16'b0011111111111111;
														assign node45 = (inp[4]) ? 16'b0000111111111111 : 16'b0001111111111111;
													assign node48 = (inp[13]) ? 16'b0000111111111111 : 16'b0001111111111111;
												assign node51 = (inp[14]) ? node53 : 16'b0000111111111111;
													assign node53 = (inp[6]) ? 16'b0000011111111111 : node54;
														assign node54 = (inp[12]) ? 16'b0000011111111111 : node55;
															assign node55 = (inp[4]) ? 16'b0000111111111111 : node56;
																assign node56 = (inp[13]) ? 16'b0000111111111111 : 16'b0001111111111111;
										assign node62 = (inp[13]) ? node90 : node63;
											assign node63 = (inp[0]) ? node79 : node64;
												assign node64 = (inp[6]) ? node74 : node65;
													assign node65 = (inp[4]) ? node69 : node66;
														assign node66 = (inp[12]) ? 16'b0001111111111111 : 16'b0011111111111111;
														assign node69 = (inp[14]) ? node71 : 16'b0001111111111111;
															assign node71 = (inp[12]) ? 16'b0000111111111111 : 16'b0001111111111111;
													assign node74 = (inp[14]) ? node76 : 16'b0001111111111111;
														assign node76 = (inp[12]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node79 = (inp[12]) ? 16'b0000011111111111 : node80;
													assign node80 = (inp[14]) ? node86 : node81;
														assign node81 = (inp[6]) ? 16'b0000111111111111 : node82;
															assign node82 = (inp[4]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node86 = (inp[1]) ? 16'b0000011111111111 : 16'b0000111111111111;
											assign node90 = (inp[6]) ? node98 : node91;
												assign node91 = (inp[0]) ? 16'b0000011111111111 : node92;
													assign node92 = (inp[1]) ? node94 : 16'b0000111111111111;
														assign node94 = (inp[14]) ? 16'b0000001111111111 : 16'b0000111111111111;
												assign node98 = (inp[0]) ? node104 : node99;
													assign node99 = (inp[1]) ? node101 : 16'b0000111111111111;
														assign node101 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node104 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
									assign node107 = (inp[0]) ? node163 : node108;
										assign node108 = (inp[14]) ? node136 : node109;
											assign node109 = (inp[4]) ? node119 : node110;
												assign node110 = (inp[12]) ? 16'b0000111111111111 : node111;
													assign node111 = (inp[6]) ? node115 : node112;
														assign node112 = (inp[2]) ? 16'b0001111111111111 : 16'b0011111111111111;
														assign node115 = (inp[13]) ? 16'b0000111111111111 : 16'b0001111111111111;
												assign node119 = (inp[6]) ? node123 : node120;
													assign node120 = (inp[1]) ? 16'b0000111111111111 : 16'b0001111111111111;
													assign node123 = (inp[12]) ? node131 : node124;
														assign node124 = (inp[2]) ? 16'b0000011111111111 : node125;
															assign node125 = (inp[1]) ? node127 : 16'b0000111111111111;
																assign node127 = (inp[13]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node131 = (inp[1]) ? node133 : 16'b0000011111111111;
															assign node133 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node136 = (inp[13]) ? node154 : node137;
												assign node137 = (inp[4]) ? node145 : node138;
													assign node138 = (inp[2]) ? node140 : 16'b0000111111111111;
														assign node140 = (inp[1]) ? node142 : 16'b0000111111111111;
															assign node142 = (inp[6]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node145 = (inp[12]) ? 16'b0000011111111111 : node146;
														assign node146 = (inp[1]) ? 16'b0000011111111111 : node147;
															assign node147 = (inp[6]) ? node149 : 16'b0000111111111111;
																assign node149 = (inp[2]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node154 = (inp[4]) ? 16'b0000001111111111 : node155;
													assign node155 = (inp[6]) ? 16'b0000011111111111 : node156;
														assign node156 = (inp[1]) ? 16'b0000011111111111 : node157;
															assign node157 = (inp[2]) ? 16'b0000011111111111 : 16'b0000111111111111;
										assign node163 = (inp[6]) ? node187 : node164;
											assign node164 = (inp[4]) ? node174 : node165;
												assign node165 = (inp[2]) ? node169 : node166;
													assign node166 = (inp[1]) ? 16'b0000111111111111 : 16'b0001111111111111;
													assign node169 = (inp[1]) ? node171 : 16'b0000111111111111;
														assign node171 = (inp[14]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node174 = (inp[14]) ? node182 : node175;
													assign node175 = (inp[1]) ? node179 : node176;
														assign node176 = (inp[12]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node179 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node182 = (inp[13]) ? node184 : 16'b0000001111111111;
														assign node184 = (inp[2]) ? 16'b0000000011111111 : 16'b0000001111111111;
											assign node187 = (inp[14]) ? node197 : node188;
												assign node188 = (inp[4]) ? node190 : 16'b0000111111111111;
													assign node190 = (inp[12]) ? 16'b0000001111111111 : node191;
														assign node191 = (inp[2]) ? node193 : 16'b0000011111111111;
															assign node193 = (inp[1]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node197 = (inp[1]) ? node201 : node198;
													assign node198 = (inp[2]) ? 16'b0000011111111111 : 16'b0000001111111111;
													assign node201 = (inp[4]) ? node205 : node202;
														assign node202 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node205 = (inp[2]) ? node207 : 16'b0000000111111111;
															assign node207 = (inp[12]) ? 16'b0000000011111111 : node208;
																assign node208 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
								assign node212 = (inp[13]) ? node326 : node213;
									assign node213 = (inp[15]) ? node263 : node214;
										assign node214 = (inp[2]) ? node244 : node215;
											assign node215 = (inp[1]) ? node227 : node216;
												assign node216 = (inp[0]) ? node222 : node217;
													assign node217 = (inp[12]) ? node219 : 16'b0011111111111111;
														assign node219 = (inp[6]) ? 16'b0000111111111111 : 16'b0011111111111111;
													assign node222 = (inp[14]) ? 16'b0000111111111111 : node223;
														assign node223 = (inp[4]) ? 16'b0000111111111111 : 16'b0001111111111111;
												assign node227 = (inp[12]) ? node233 : node228;
													assign node228 = (inp[14]) ? 16'b0000111111111111 : node229;
														assign node229 = (inp[0]) ? 16'b0000111111111111 : 16'b0011111111111111;
													assign node233 = (inp[14]) ? node241 : node234;
														assign node234 = (inp[4]) ? node236 : 16'b0000111111111111;
															assign node236 = (inp[0]) ? 16'b0000011111111111 : node237;
																assign node237 = (inp[6]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node241 = (inp[6]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node244 = (inp[6]) ? node256 : node245;
												assign node245 = (inp[12]) ? node251 : node246;
													assign node246 = (inp[0]) ? node248 : 16'b0000111111111111;
														assign node248 = (inp[14]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node251 = (inp[4]) ? 16'b0000011111111111 : node252;
														assign node252 = (inp[0]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node256 = (inp[12]) ? 16'b0000000111111111 : node257;
													assign node257 = (inp[4]) ? 16'b0000001111111111 : node258;
														assign node258 = (inp[0]) ? 16'b0000011111111111 : 16'b0000111111111111;
										assign node263 = (inp[12]) ? node287 : node264;
											assign node264 = (inp[14]) ? node278 : node265;
												assign node265 = (inp[6]) ? node273 : node266;
													assign node266 = (inp[0]) ? node270 : node267;
														assign node267 = (inp[2]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node270 = (inp[4]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node273 = (inp[1]) ? node275 : 16'b0000011111111111;
														assign node275 = (inp[4]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node278 = (inp[4]) ? node280 : 16'b0000011111111111;
													assign node280 = (inp[2]) ? 16'b0000000111111111 : node281;
														assign node281 = (inp[0]) ? node283 : 16'b0000011111111111;
															assign node283 = (inp[1]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node287 = (inp[4]) ? node313 : node288;
												assign node288 = (inp[6]) ? node296 : node289;
													assign node289 = (inp[1]) ? 16'b0000011111111111 : node290;
														assign node290 = (inp[14]) ? 16'b0000111111111111 : node291;
															assign node291 = (inp[0]) ? 16'b0000111111111111 : 16'b0001111111111111;
													assign node296 = (inp[14]) ? node308 : node297;
														assign node297 = (inp[0]) ? node303 : node298;
															assign node298 = (inp[2]) ? node300 : 16'b0000011111111111;
																assign node300 = (inp[1]) ? 16'b0000001111111111 : 16'b0000011111111111;
															assign node303 = (inp[1]) ? 16'b0000001111111111 : node304;
																assign node304 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node308 = (inp[2]) ? node310 : 16'b0000001111111111;
															assign node310 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node313 = (inp[2]) ? 16'b0000000111111111 : node314;
													assign node314 = (inp[1]) ? node320 : node315;
														assign node315 = (inp[0]) ? 16'b0000001111111111 : node316;
															assign node316 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node320 = (inp[14]) ? node322 : 16'b0000001111111111;
															assign node322 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
									assign node326 = (inp[6]) ? node368 : node327;
										assign node327 = (inp[12]) ? node347 : node328;
											assign node328 = (inp[14]) ? node336 : node329;
												assign node329 = (inp[1]) ? 16'b0000011111111111 : node330;
													assign node330 = (inp[0]) ? 16'b0000111111111111 : node331;
														assign node331 = (inp[15]) ? 16'b0001111111111111 : 16'b0011111111111111;
												assign node336 = (inp[15]) ? node342 : node337;
													assign node337 = (inp[2]) ? node339 : 16'b0000011111111111;
														assign node339 = (inp[1]) ? 16'b0000000111111111 : 16'b0000011111111111;
													assign node342 = (inp[4]) ? 16'b0000001111111111 : node343;
														assign node343 = (inp[0]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node347 = (inp[0]) ? node355 : node348;
												assign node348 = (inp[2]) ? node350 : 16'b0000011111111111;
													assign node350 = (inp[4]) ? 16'b0000001111111111 : node351;
														assign node351 = (inp[1]) ? 16'b0000001111111111 : 16'b0000111111111111;
												assign node355 = (inp[2]) ? node363 : node356;
													assign node356 = (inp[14]) ? node360 : node357;
														assign node357 = (inp[1]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node360 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node363 = (inp[1]) ? node365 : 16'b0000001111111111;
														assign node365 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node368 = (inp[15]) ? node400 : node369;
											assign node369 = (inp[4]) ? node389 : node370;
												assign node370 = (inp[2]) ? node380 : node371;
													assign node371 = (inp[12]) ? node375 : node372;
														assign node372 = (inp[1]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node375 = (inp[14]) ? node377 : 16'b0000011111111111;
															assign node377 = (inp[0]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node380 = (inp[1]) ? node384 : node381;
														assign node381 = (inp[0]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node384 = (inp[0]) ? 16'b0000000111111111 : node385;
															assign node385 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node389 = (inp[2]) ? node393 : node390;
													assign node390 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node393 = (inp[14]) ? node397 : node394;
														assign node394 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node397 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node400 = (inp[2]) ? node410 : node401;
												assign node401 = (inp[12]) ? node403 : 16'b0000001111111111;
													assign node403 = (inp[4]) ? node405 : 16'b0000001111111111;
														assign node405 = (inp[14]) ? 16'b0000000011111111 : node406;
															assign node406 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node410 = (inp[1]) ? node414 : node411;
													assign node411 = (inp[4]) ? 16'b0000000111111111 : 16'b0000000011111111;
													assign node414 = (inp[4]) ? node416 : 16'b0000000011111111;
														assign node416 = (inp[0]) ? node418 : 16'b0000000011111111;
															assign node418 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
							assign node421 = (inp[2]) ? node591 : node422;
								assign node422 = (inp[0]) ? node504 : node423;
									assign node423 = (inp[14]) ? node455 : node424;
										assign node424 = (inp[15]) ? node442 : node425;
											assign node425 = (inp[4]) ? node435 : node426;
												assign node426 = (inp[12]) ? node432 : node427;
													assign node427 = (inp[1]) ? 16'b0001111111111111 : node428;
														assign node428 = (inp[5]) ? 16'b0001111111111111 : 16'b0011111111111111;
													assign node432 = (inp[5]) ? 16'b0000011111111111 : 16'b0001111111111111;
												assign node435 = (inp[12]) ? 16'b0001111111111111 : node436;
													assign node436 = (inp[1]) ? node438 : 16'b0000111111111111;
														assign node438 = (inp[13]) ? 16'b0000011111111111 : 16'b0000111111111111;
											assign node442 = (inp[6]) ? node452 : node443;
												assign node443 = (inp[12]) ? node449 : node444;
													assign node444 = (inp[1]) ? 16'b0000111111111111 : node445;
														assign node445 = (inp[5]) ? 16'b0000111111111111 : 16'b0011111111111111;
													assign node449 = (inp[1]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node452 = (inp[1]) ? 16'b0000001111111111 : 16'b0000011111111111;
										assign node455 = (inp[5]) ? node481 : node456;
											assign node456 = (inp[1]) ? node470 : node457;
												assign node457 = (inp[6]) ? 16'b0000011111111111 : node458;
													assign node458 = (inp[15]) ? node464 : node459;
														assign node459 = (inp[12]) ? 16'b0000111111111111 : node460;
															assign node460 = (inp[13]) ? 16'b0001111111111111 : 16'b0011111111111111;
														assign node464 = (inp[12]) ? node466 : 16'b0000111111111111;
															assign node466 = (inp[4]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node470 = (inp[4]) ? 16'b0000001111111111 : node471;
													assign node471 = (inp[12]) ? node473 : 16'b0000111111111111;
														assign node473 = (inp[6]) ? node475 : 16'b0000011111111111;
															assign node475 = (inp[13]) ? 16'b0000001111111111 : node476;
																assign node476 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node481 = (inp[15]) ? node489 : node482;
												assign node482 = (inp[13]) ? node484 : 16'b0000011111111111;
													assign node484 = (inp[6]) ? node486 : 16'b0000000111111111;
														assign node486 = (inp[4]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node489 = (inp[13]) ? node499 : node490;
													assign node490 = (inp[6]) ? node494 : node491;
														assign node491 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node494 = (inp[4]) ? 16'b0000000111111111 : node495;
															assign node495 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node499 = (inp[6]) ? node501 : 16'b0000000111111111;
														assign node501 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node504 = (inp[4]) ? node548 : node505;
										assign node505 = (inp[1]) ? node521 : node506;
											assign node506 = (inp[12]) ? node512 : node507;
												assign node507 = (inp[6]) ? node509 : 16'b0001111111111111;
													assign node509 = (inp[5]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node512 = (inp[5]) ? node516 : node513;
													assign node513 = (inp[14]) ? 16'b0000111111111111 : 16'b0000011111111111;
													assign node516 = (inp[6]) ? node518 : 16'b0000011111111111;
														assign node518 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node521 = (inp[5]) ? node531 : node522;
												assign node522 = (inp[12]) ? node524 : 16'b0000011111111111;
													assign node524 = (inp[15]) ? node528 : node525;
														assign node525 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node528 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node531 = (inp[15]) ? node543 : node532;
													assign node532 = (inp[12]) ? node540 : node533;
														assign node533 = (inp[6]) ? node535 : 16'b0000001111111111;
															assign node535 = (inp[13]) ? node537 : 16'b0000001111111111;
																assign node537 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node540 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node543 = (inp[14]) ? node545 : 16'b0000001111111111;
														assign node545 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node548 = (inp[12]) ? node570 : node549;
											assign node549 = (inp[13]) ? node561 : node550;
												assign node550 = (inp[6]) ? node556 : node551;
													assign node551 = (inp[1]) ? 16'b0000011111111111 : node552;
														assign node552 = (inp[5]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node556 = (inp[15]) ? 16'b0000000111111111 : node557;
														assign node557 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node561 = (inp[14]) ? node563 : 16'b0000001111111111;
													assign node563 = (inp[1]) ? node567 : node564;
														assign node564 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node567 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node570 = (inp[6]) ? node574 : node571;
												assign node571 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node574 = (inp[14]) ? node582 : node575;
													assign node575 = (inp[15]) ? 16'b0000000111111111 : node576;
														assign node576 = (inp[1]) ? node578 : 16'b0000000111111111;
															assign node578 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node582 = (inp[1]) ? 16'b0000000011111111 : node583;
														assign node583 = (inp[15]) ? 16'b0000000011111111 : node584;
															assign node584 = (inp[13]) ? node586 : 16'b0000000111111111;
																assign node586 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
								assign node591 = (inp[12]) ? node679 : node592;
									assign node592 = (inp[5]) ? node634 : node593;
										assign node593 = (inp[15]) ? node611 : node594;
											assign node594 = (inp[1]) ? node606 : node595;
												assign node595 = (inp[13]) ? node601 : node596;
													assign node596 = (inp[6]) ? 16'b0000111111111111 : node597;
														assign node597 = (inp[4]) ? 16'b0000111111111111 : 16'b0001111111111111;
													assign node601 = (inp[4]) ? 16'b0000001111111111 : node602;
														assign node602 = (inp[0]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node606 = (inp[6]) ? node608 : 16'b0000011111111111;
													assign node608 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node611 = (inp[13]) ? node619 : node612;
												assign node612 = (inp[1]) ? node614 : 16'b0000011111111111;
													assign node614 = (inp[6]) ? 16'b0000001111111111 : node615;
														assign node615 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node619 = (inp[14]) ? node629 : node620;
													assign node620 = (inp[0]) ? node626 : node621;
														assign node621 = (inp[1]) ? 16'b0000001111111111 : node622;
															assign node622 = (inp[4]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node626 = (inp[6]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node629 = (inp[6]) ? node631 : 16'b0000001111111111;
														assign node631 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node634 = (inp[6]) ? node654 : node635;
											assign node635 = (inp[0]) ? node645 : node636;
												assign node636 = (inp[13]) ? 16'b0000001111111111 : node637;
													assign node637 = (inp[14]) ? 16'b0000001111111111 : node638;
														assign node638 = (inp[1]) ? node640 : 16'b0000011111111111;
															assign node640 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node645 = (inp[4]) ? node649 : node646;
													assign node646 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node649 = (inp[14]) ? 16'b0000000111111111 : node650;
														assign node650 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node654 = (inp[15]) ? node666 : node655;
												assign node655 = (inp[0]) ? node661 : node656;
													assign node656 = (inp[4]) ? node658 : 16'b0000001111111111;
														assign node658 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node661 = (inp[13]) ? 16'b0000000111111111 : node662;
														assign node662 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node666 = (inp[1]) ? node674 : node667;
													assign node667 = (inp[0]) ? node671 : node668;
														assign node668 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node671 = (inp[14]) ? 16'b0000000111111111 : 16'b0000000011111111;
													assign node674 = (inp[4]) ? node676 : 16'b0000000011111111;
														assign node676 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node679 = (inp[13]) ? node727 : node680;
										assign node680 = (inp[0]) ? node702 : node681;
											assign node681 = (inp[5]) ? node693 : node682;
												assign node682 = (inp[14]) ? 16'b0000001111111111 : node683;
													assign node683 = (inp[4]) ? 16'b0000001111111111 : node684;
														assign node684 = (inp[1]) ? 16'b0000011111111111 : node685;
															assign node685 = (inp[6]) ? node687 : 16'b0000111111111111;
																assign node687 = (inp[15]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node693 = (inp[1]) ? node695 : 16'b0000001111111111;
													assign node695 = (inp[15]) ? node699 : node696;
														assign node696 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node699 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node702 = (inp[14]) ? node718 : node703;
												assign node703 = (inp[6]) ? node709 : node704;
													assign node704 = (inp[5]) ? 16'b0000001111111111 : node705;
														assign node705 = (inp[15]) ? 16'b0000011111111111 : 16'b0000001111111111;
													assign node709 = (inp[1]) ? 16'b0000000011111111 : node710;
														assign node710 = (inp[4]) ? node712 : 16'b0000001111111111;
															assign node712 = (inp[5]) ? 16'b0000000111111111 : node713;
																assign node713 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node718 = (inp[4]) ? node722 : node719;
													assign node719 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node722 = (inp[6]) ? 16'b0000000001111111 : node723;
														assign node723 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node727 = (inp[1]) ? node745 : node728;
											assign node728 = (inp[4]) ? node734 : node729;
												assign node729 = (inp[5]) ? node731 : 16'b0000001111111111;
													assign node731 = (inp[6]) ? 16'b0000000111111111 : 16'b0000011111111111;
												assign node734 = (inp[0]) ? 16'b0000000011111111 : node735;
													assign node735 = (inp[6]) ? node737 : 16'b0000000111111111;
														assign node737 = (inp[15]) ? node739 : 16'b0000000111111111;
															assign node739 = (inp[5]) ? node741 : 16'b0000000011111111;
																assign node741 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node745 = (inp[4]) ? node753 : node746;
												assign node746 = (inp[5]) ? 16'b0000000011111111 : node747;
													assign node747 = (inp[0]) ? node749 : 16'b0000000111111111;
														assign node749 = (inp[14]) ? 16'b0000000111111111 : 16'b0000000011111111;
												assign node753 = (inp[5]) ? node755 : 16'b0000000011111111;
													assign node755 = (inp[6]) ? 16'b0000000000011111 : 16'b0000000011111111;
						assign node758 = (inp[0]) ? node1116 : node759;
							assign node759 = (inp[13]) ? node925 : node760;
								assign node760 = (inp[6]) ? node858 : node761;
									assign node761 = (inp[4]) ? node813 : node762;
										assign node762 = (inp[12]) ? node792 : node763;
											assign node763 = (inp[5]) ? node779 : node764;
												assign node764 = (inp[1]) ? node770 : node765;
													assign node765 = (inp[15]) ? node767 : 16'b0011111111111111;
														assign node767 = (inp[8]) ? 16'b0000111111111111 : 16'b0001111111111111;
													assign node770 = (inp[8]) ? node774 : node771;
														assign node771 = (inp[14]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node774 = (inp[14]) ? node776 : 16'b0000111111111111;
															assign node776 = (inp[15]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node779 = (inp[14]) ? node787 : node780;
													assign node780 = (inp[15]) ? node784 : node781;
														assign node781 = (inp[1]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node784 = (inp[1]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node787 = (inp[2]) ? 16'b0000011111111111 : node788;
														assign node788 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node792 = (inp[2]) ? node802 : node793;
												assign node793 = (inp[14]) ? 16'b0000011111111111 : node794;
													assign node794 = (inp[1]) ? node796 : 16'b0000111111111111;
														assign node796 = (inp[8]) ? 16'b0000011111111111 : node797;
															assign node797 = (inp[15]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node802 = (inp[5]) ? node808 : node803;
													assign node803 = (inp[14]) ? node805 : 16'b0000011111111111;
														assign node805 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node808 = (inp[14]) ? 16'b0000000111111111 : node809;
														assign node809 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
										assign node813 = (inp[5]) ? node837 : node814;
											assign node814 = (inp[12]) ? node822 : node815;
												assign node815 = (inp[15]) ? 16'b0000011111111111 : node816;
													assign node816 = (inp[14]) ? 16'b0000111111111111 : node817;
														assign node817 = (inp[8]) ? 16'b0000111111111111 : 16'b0001111111111111;
												assign node822 = (inp[2]) ? node830 : node823;
													assign node823 = (inp[15]) ? node827 : node824;
														assign node824 = (inp[1]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node827 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node830 = (inp[15]) ? 16'b0000001111111111 : node831;
														assign node831 = (inp[14]) ? 16'b0000001111111111 : node832;
															assign node832 = (inp[1]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node837 = (inp[1]) ? node843 : node838;
												assign node838 = (inp[8]) ? node840 : 16'b0000011111111111;
													assign node840 = (inp[15]) ? 16'b0000001111111111 : 16'b0000000111111111;
												assign node843 = (inp[8]) ? node849 : node844;
													assign node844 = (inp[15]) ? node846 : 16'b0000001111111111;
														assign node846 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node849 = (inp[15]) ? node855 : node850;
														assign node850 = (inp[12]) ? 16'b0000000111111111 : node851;
															assign node851 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node855 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node858 = (inp[8]) ? node892 : node859;
										assign node859 = (inp[1]) ? node875 : node860;
											assign node860 = (inp[12]) ? node870 : node861;
												assign node861 = (inp[14]) ? node863 : 16'b0000111111111111;
													assign node863 = (inp[2]) ? node865 : 16'b0000111111111111;
														assign node865 = (inp[15]) ? node867 : 16'b0000011111111111;
															assign node867 = (inp[4]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node870 = (inp[14]) ? node872 : 16'b0000011111111111;
													assign node872 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node875 = (inp[14]) ? 16'b0000001111111111 : node876;
												assign node876 = (inp[2]) ? node882 : node877;
													assign node877 = (inp[15]) ? node879 : 16'b0000011111111111;
														assign node879 = (inp[12]) ? 16'b0000011111111111 : 16'b0000001111111111;
													assign node882 = (inp[4]) ? node886 : node883;
														assign node883 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node886 = (inp[5]) ? 16'b0000001111111111 : node887;
															assign node887 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
										assign node892 = (inp[15]) ? node908 : node893;
											assign node893 = (inp[1]) ? node903 : node894;
												assign node894 = (inp[4]) ? 16'b0000001111111111 : node895;
													assign node895 = (inp[5]) ? node897 : 16'b0000111111111111;
														assign node897 = (inp[2]) ? node899 : 16'b0000011111111111;
															assign node899 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node903 = (inp[4]) ? node905 : 16'b0000001111111111;
													assign node905 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node908 = (inp[12]) ? node914 : node909;
												assign node909 = (inp[4]) ? 16'b0000000001111111 : node910;
													assign node910 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node914 = (inp[1]) ? node918 : node915;
													assign node915 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node918 = (inp[14]) ? node920 : 16'b0000000011111111;
														assign node920 = (inp[5]) ? node922 : 16'b0000000011111111;
															assign node922 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
								assign node925 = (inp[15]) ? node1013 : node926;
									assign node926 = (inp[2]) ? node978 : node927;
										assign node927 = (inp[5]) ? node955 : node928;
											assign node928 = (inp[1]) ? node942 : node929;
												assign node929 = (inp[12]) ? node937 : node930;
													assign node930 = (inp[14]) ? node934 : node931;
														assign node931 = (inp[6]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node934 = (inp[4]) ? 16'b0000001111111111 : 16'b0000111111111111;
													assign node937 = (inp[4]) ? 16'b0000011111111111 : node938;
														assign node938 = (inp[8]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node942 = (inp[4]) ? node950 : node943;
													assign node943 = (inp[12]) ? node945 : 16'b0000111111111111;
														assign node945 = (inp[14]) ? node947 : 16'b0000011111111111;
															assign node947 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node950 = (inp[12]) ? 16'b0000001111111111 : node951;
														assign node951 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node955 = (inp[12]) ? node971 : node956;
												assign node956 = (inp[6]) ? node964 : node957;
													assign node957 = (inp[1]) ? 16'b0000011111111111 : node958;
														assign node958 = (inp[14]) ? 16'b0000011111111111 : node959;
															assign node959 = (inp[4]) ? 16'b0000111111111111 : 16'b0001111111111111;
													assign node964 = (inp[4]) ? node968 : node965;
														assign node965 = (inp[1]) ? 16'b0000011111111111 : 16'b0000001111111111;
														assign node968 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node971 = (inp[8]) ? node973 : 16'b0000001111111111;
													assign node973 = (inp[6]) ? node975 : 16'b0000000111111111;
														assign node975 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000111111111;
										assign node978 = (inp[12]) ? node990 : node979;
											assign node979 = (inp[8]) ? node987 : node980;
												assign node980 = (inp[6]) ? 16'b0000001111111111 : node981;
													assign node981 = (inp[1]) ? node983 : 16'b0000011111111111;
														assign node983 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node987 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node990 = (inp[5]) ? node1006 : node991;
												assign node991 = (inp[1]) ? node997 : node992;
													assign node992 = (inp[4]) ? node994 : 16'b0000111111111111;
														assign node994 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node997 = (inp[14]) ? node1001 : node998;
														assign node998 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node1001 = (inp[4]) ? node1003 : 16'b0000000111111111;
															assign node1003 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node1006 = (inp[8]) ? node1008 : 16'b0000000111111111;
													assign node1008 = (inp[6]) ? 16'b0000000001111111 : node1009;
														assign node1009 = (inp[14]) ? 16'b0000000111111111 : 16'b0000000011111111;
									assign node1013 = (inp[6]) ? node1063 : node1014;
										assign node1014 = (inp[14]) ? node1034 : node1015;
											assign node1015 = (inp[8]) ? node1025 : node1016;
												assign node1016 = (inp[12]) ? node1020 : node1017;
													assign node1017 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node1020 = (inp[4]) ? 16'b0000001111111111 : node1021;
														assign node1021 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node1025 = (inp[5]) ? 16'b0000000111111111 : node1026;
													assign node1026 = (inp[1]) ? node1030 : node1027;
														assign node1027 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node1030 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node1034 = (inp[2]) ? node1046 : node1035;
												assign node1035 = (inp[4]) ? node1041 : node1036;
													assign node1036 = (inp[1]) ? node1038 : 16'b0000011111111111;
														assign node1038 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node1041 = (inp[5]) ? 16'b0000000011111111 : node1042;
														assign node1042 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node1046 = (inp[8]) ? node1058 : node1047;
													assign node1047 = (inp[4]) ? node1053 : node1048;
														assign node1048 = (inp[12]) ? node1050 : 16'b0000001111111111;
															assign node1050 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node1053 = (inp[5]) ? node1055 : 16'b0000000111111111;
															assign node1055 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node1058 = (inp[1]) ? node1060 : 16'b0000000011111111;
														assign node1060 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node1063 = (inp[14]) ? node1099 : node1064;
											assign node1064 = (inp[2]) ? node1082 : node1065;
												assign node1065 = (inp[1]) ? node1073 : node1066;
													assign node1066 = (inp[12]) ? node1070 : node1067;
														assign node1067 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node1070 = (inp[4]) ? 16'b0000000111111111 : 16'b0000011111111111;
													assign node1073 = (inp[5]) ? 16'b0000000111111111 : node1074;
														assign node1074 = (inp[4]) ? 16'b0000000111111111 : node1075;
															assign node1075 = (inp[12]) ? node1077 : 16'b0000001111111111;
																assign node1077 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node1082 = (inp[12]) ? node1088 : node1083;
													assign node1083 = (inp[8]) ? node1085 : 16'b0000000111111111;
														assign node1085 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node1088 = (inp[4]) ? node1092 : node1089;
														assign node1089 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node1092 = (inp[1]) ? node1094 : 16'b0000000011111111;
															assign node1094 = (inp[8]) ? 16'b0000000001111111 : node1095;
																assign node1095 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node1099 = (inp[4]) ? node1111 : node1100;
												assign node1100 = (inp[8]) ? node1108 : node1101;
													assign node1101 = (inp[5]) ? node1103 : 16'b0000001111111111;
														assign node1103 = (inp[1]) ? 16'b0000000011111111 : node1104;
															assign node1104 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node1108 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node1111 = (inp[5]) ? 16'b0000000001111111 : node1112;
													assign node1112 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
							assign node1116 = (inp[2]) ? node1288 : node1117;
								assign node1117 = (inp[4]) ? node1195 : node1118;
									assign node1118 = (inp[12]) ? node1152 : node1119;
										assign node1119 = (inp[5]) ? node1133 : node1120;
											assign node1120 = (inp[14]) ? node1126 : node1121;
												assign node1121 = (inp[8]) ? node1123 : 16'b0000111111111111;
													assign node1123 = (inp[13]) ? 16'b0000001111111111 : 16'b0000111111111111;
												assign node1126 = (inp[13]) ? 16'b0000001111111111 : node1127;
													assign node1127 = (inp[1]) ? 16'b0000011111111111 : node1128;
														assign node1128 = (inp[6]) ? 16'b0000011111111111 : 16'b0000111111111111;
											assign node1133 = (inp[6]) ? node1149 : node1134;
												assign node1134 = (inp[8]) ? node1140 : node1135;
													assign node1135 = (inp[15]) ? 16'b0000011111111111 : node1136;
														assign node1136 = (inp[13]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node1140 = (inp[13]) ? node1146 : node1141;
														assign node1141 = (inp[1]) ? 16'b0000001111111111 : node1142;
															assign node1142 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node1146 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node1149 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node1152 = (inp[5]) ? node1176 : node1153;
											assign node1153 = (inp[14]) ? node1165 : node1154;
												assign node1154 = (inp[13]) ? node1158 : node1155;
													assign node1155 = (inp[1]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node1158 = (inp[8]) ? 16'b0000000111111111 : node1159;
														assign node1159 = (inp[6]) ? 16'b0000001111111111 : node1160;
															assign node1160 = (inp[1]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node1165 = (inp[13]) ? node1173 : node1166;
													assign node1166 = (inp[15]) ? 16'b0000000111111111 : node1167;
														assign node1167 = (inp[8]) ? 16'b0000001111111111 : node1168;
															assign node1168 = (inp[1]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node1173 = (inp[15]) ? 16'b0000001111111111 : 16'b0000000111111111;
											assign node1176 = (inp[14]) ? node1184 : node1177;
												assign node1177 = (inp[1]) ? node1179 : 16'b0000011111111111;
													assign node1179 = (inp[13]) ? 16'b0000000111111111 : node1180;
														assign node1180 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node1184 = (inp[13]) ? node1190 : node1185;
													assign node1185 = (inp[15]) ? node1187 : 16'b0000001111111111;
														assign node1187 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node1190 = (inp[8]) ? 16'b0000000011111111 : node1191;
														assign node1191 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node1195 = (inp[6]) ? node1235 : node1196;
										assign node1196 = (inp[8]) ? node1218 : node1197;
											assign node1197 = (inp[12]) ? node1207 : node1198;
												assign node1198 = (inp[14]) ? node1202 : node1199;
													assign node1199 = (inp[15]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node1202 = (inp[1]) ? node1204 : 16'b0000011111111111;
														assign node1204 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node1207 = (inp[15]) ? node1213 : node1208;
													assign node1208 = (inp[5]) ? 16'b0000001111111111 : node1209;
														assign node1209 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node1213 = (inp[5]) ? 16'b0000000011111111 : node1214;
														assign node1214 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node1218 = (inp[1]) ? node1228 : node1219;
												assign node1219 = (inp[14]) ? node1223 : node1220;
													assign node1220 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node1223 = (inp[15]) ? 16'b0000000011111111 : node1224;
														assign node1224 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node1228 = (inp[5]) ? node1230 : 16'b0000000111111111;
													assign node1230 = (inp[15]) ? node1232 : 16'b0000000011111111;
														assign node1232 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000011111111;
										assign node1235 = (inp[5]) ? node1265 : node1236;
											assign node1236 = (inp[13]) ? node1252 : node1237;
												assign node1237 = (inp[15]) ? node1247 : node1238;
													assign node1238 = (inp[1]) ? node1240 : 16'b0000001111111111;
														assign node1240 = (inp[14]) ? 16'b0000000111111111 : node1241;
															assign node1241 = (inp[8]) ? node1243 : 16'b0000001111111111;
																assign node1243 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node1247 = (inp[8]) ? node1249 : 16'b0000001111111111;
														assign node1249 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node1252 = (inp[12]) ? node1258 : node1253;
													assign node1253 = (inp[1]) ? 16'b0000000111111111 : node1254;
														assign node1254 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node1258 = (inp[14]) ? node1260 : 16'b0000000111111111;
														assign node1260 = (inp[8]) ? 16'b0000000001111111 : node1261;
															assign node1261 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node1265 = (inp[1]) ? node1277 : node1266;
												assign node1266 = (inp[8]) ? node1272 : node1267;
													assign node1267 = (inp[13]) ? node1269 : 16'b0000001111111111;
														assign node1269 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node1272 = (inp[13]) ? 16'b0000000011111111 : node1273;
														assign node1273 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node1277 = (inp[14]) ? node1283 : node1278;
													assign node1278 = (inp[15]) ? node1280 : 16'b0000000011111111;
														assign node1280 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node1283 = (inp[13]) ? node1285 : 16'b0000000001111111;
														assign node1285 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
								assign node1288 = (inp[1]) ? node1382 : node1289;
									assign node1289 = (inp[4]) ? node1341 : node1290;
										assign node1290 = (inp[14]) ? node1310 : node1291;
											assign node1291 = (inp[6]) ? node1301 : node1292;
												assign node1292 = (inp[8]) ? 16'b0000001111111111 : node1293;
													assign node1293 = (inp[15]) ? node1297 : node1294;
														assign node1294 = (inp[12]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node1297 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node1301 = (inp[13]) ? node1305 : node1302;
													assign node1302 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node1305 = (inp[5]) ? node1307 : 16'b0000000111111111;
														assign node1307 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node1310 = (inp[13]) ? node1326 : node1311;
												assign node1311 = (inp[6]) ? node1319 : node1312;
													assign node1312 = (inp[12]) ? node1316 : node1313;
														assign node1313 = (inp[5]) ? 16'b0000001111111111 : 16'b0000111111111111;
														assign node1316 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node1319 = (inp[5]) ? 16'b0000000111111111 : node1320;
														assign node1320 = (inp[8]) ? node1322 : 16'b0000001111111111;
															assign node1322 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node1326 = (inp[6]) ? node1334 : node1327;
													assign node1327 = (inp[15]) ? node1329 : 16'b0000000111111111;
														assign node1329 = (inp[5]) ? 16'b0000000111111111 : node1330;
															assign node1330 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node1334 = (inp[8]) ? node1336 : 16'b0000000011111111;
														assign node1336 = (inp[5]) ? node1338 : 16'b0000000011111111;
															assign node1338 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node1341 = (inp[15]) ? node1363 : node1342;
											assign node1342 = (inp[12]) ? node1358 : node1343;
												assign node1343 = (inp[5]) ? node1349 : node1344;
													assign node1344 = (inp[8]) ? node1346 : 16'b0000001111111111;
														assign node1346 = (inp[6]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node1349 = (inp[8]) ? node1353 : node1350;
														assign node1350 = (inp[6]) ? 16'b0000001111111111 : 16'b0000000111111111;
														assign node1353 = (inp[6]) ? node1355 : 16'b0000000111111111;
															assign node1355 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000111111111;
												assign node1358 = (inp[13]) ? 16'b0000000011111111 : node1359;
													assign node1359 = (inp[14]) ? 16'b0000000011111111 : 16'b0000001111111111;
											assign node1363 = (inp[5]) ? node1371 : node1364;
												assign node1364 = (inp[6]) ? node1366 : 16'b0000000111111111;
													assign node1366 = (inp[8]) ? 16'b0000000011111111 : node1367;
														assign node1367 = (inp[13]) ? 16'b0000000111111111 : 16'b0000000011111111;
												assign node1371 = (inp[14]) ? node1373 : 16'b0000000000111111;
													assign node1373 = (inp[8]) ? 16'b0000000001111111 : node1374;
														assign node1374 = (inp[6]) ? node1376 : 16'b0000000011111111;
															assign node1376 = (inp[12]) ? 16'b0000000001111111 : node1377;
																assign node1377 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node1382 = (inp[13]) ? node1442 : node1383;
										assign node1383 = (inp[5]) ? node1413 : node1384;
											assign node1384 = (inp[12]) ? node1396 : node1385;
												assign node1385 = (inp[8]) ? 16'b0000000111111111 : node1386;
													assign node1386 = (inp[6]) ? node1390 : node1387;
														assign node1387 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node1390 = (inp[14]) ? 16'b0000000111111111 : node1391;
															assign node1391 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node1396 = (inp[8]) ? node1404 : node1397;
													assign node1397 = (inp[15]) ? node1401 : node1398;
														assign node1398 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node1401 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node1404 = (inp[14]) ? 16'b0000000011111111 : node1405;
														assign node1405 = (inp[4]) ? node1407 : 16'b0000000111111111;
															assign node1407 = (inp[6]) ? 16'b0000000011111111 : node1408;
																assign node1408 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node1413 = (inp[4]) ? node1431 : node1414;
												assign node1414 = (inp[6]) ? node1422 : node1415;
													assign node1415 = (inp[12]) ? node1419 : node1416;
														assign node1416 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node1419 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node1422 = (inp[12]) ? node1428 : node1423;
														assign node1423 = (inp[14]) ? node1425 : 16'b0000000011111111;
															assign node1425 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node1428 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node1431 = (inp[15]) ? node1437 : node1432;
													assign node1432 = (inp[12]) ? node1434 : 16'b0000001111111111;
														assign node1434 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node1437 = (inp[12]) ? node1439 : 16'b0000000001111111;
														assign node1439 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node1442 = (inp[15]) ? node1460 : node1443;
											assign node1443 = (inp[8]) ? node1449 : node1444;
												assign node1444 = (inp[6]) ? 16'b0000000011111111 : node1445;
													assign node1445 = (inp[4]) ? 16'b0000000011111111 : 16'b0000001111111111;
												assign node1449 = (inp[14]) ? 16'b0000000001111111 : node1450;
													assign node1450 = (inp[6]) ? node1456 : node1451;
														assign node1451 = (inp[12]) ? 16'b0000000011111111 : node1452;
															assign node1452 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node1456 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000001111111;
											assign node1460 = (inp[6]) ? node1472 : node1461;
												assign node1461 = (inp[5]) ? 16'b0000000001111111 : node1462;
													assign node1462 = (inp[14]) ? node1464 : 16'b0000000111111111;
														assign node1464 = (inp[12]) ? 16'b0000000001111111 : node1465;
															assign node1465 = (inp[8]) ? node1467 : 16'b0000000011111111;
																assign node1467 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node1472 = (inp[14]) ? node1474 : 16'b0000000001111111;
													assign node1474 = (inp[4]) ? 16'b0000000000111111 : node1475;
														assign node1475 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
					assign node1479 = (inp[0]) ? node2259 : node1480;
						assign node1480 = (inp[4]) ? node1858 : node1481;
							assign node1481 = (inp[2]) ? node1647 : node1482;
								assign node1482 = (inp[6]) ? node1562 : node1483;
									assign node1483 = (inp[1]) ? node1519 : node1484;
										assign node1484 = (inp[8]) ? node1508 : node1485;
											assign node1485 = (inp[13]) ? node1499 : node1486;
												assign node1486 = (inp[5]) ? node1494 : node1487;
													assign node1487 = (inp[14]) ? node1489 : 16'b0011111111111111;
														assign node1489 = (inp[9]) ? 16'b0001111111111111 : node1490;
															assign node1490 = (inp[12]) ? 16'b0001111111111111 : 16'b0011111111111111;
													assign node1494 = (inp[12]) ? 16'b0000111111111111 : node1495;
														assign node1495 = (inp[14]) ? 16'b0000111111111111 : 16'b0011111111111111;
												assign node1499 = (inp[14]) ? 16'b0000111111111111 : node1500;
													assign node1500 = (inp[9]) ? node1502 : 16'b0001111111111111;
														assign node1502 = (inp[15]) ? node1504 : 16'b0001111111111111;
															assign node1504 = (inp[12]) ? 16'b0000011111111111 : 16'b0000111111111111;
											assign node1508 = (inp[5]) ? node1516 : node1509;
												assign node1509 = (inp[14]) ? 16'b0000111111111111 : node1510;
													assign node1510 = (inp[13]) ? 16'b0000111111111111 : node1511;
														assign node1511 = (inp[15]) ? 16'b0000111111111111 : 16'b0001111111111111;
												assign node1516 = (inp[12]) ? 16'b0000011111111111 : 16'b0000001111111111;
										assign node1519 = (inp[14]) ? node1543 : node1520;
											assign node1520 = (inp[8]) ? node1538 : node1521;
												assign node1521 = (inp[13]) ? node1527 : node1522;
													assign node1522 = (inp[9]) ? 16'b0000111111111111 : node1523;
														assign node1523 = (inp[12]) ? 16'b0000111111111111 : 16'b0001111111111111;
													assign node1527 = (inp[15]) ? node1535 : node1528;
														assign node1528 = (inp[12]) ? 16'b0000011111111111 : node1529;
															assign node1529 = (inp[9]) ? 16'b0000111111111111 : node1530;
																assign node1530 = (inp[5]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node1535 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node1538 = (inp[9]) ? 16'b0000001111111111 : node1539;
													assign node1539 = (inp[15]) ? 16'b0000111111111111 : 16'b0000011111111111;
											assign node1543 = (inp[9]) ? node1551 : node1544;
												assign node1544 = (inp[5]) ? 16'b0000001111111111 : node1545;
													assign node1545 = (inp[8]) ? 16'b0000011111111111 : node1546;
														assign node1546 = (inp[13]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node1551 = (inp[15]) ? node1557 : node1552;
													assign node1552 = (inp[5]) ? 16'b0000000111111111 : node1553;
														assign node1553 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node1557 = (inp[5]) ? node1559 : 16'b0000000111111111;
														assign node1559 = (inp[8]) ? 16'b0000000111111111 : 16'b0000000011111111;
									assign node1562 = (inp[9]) ? node1610 : node1563;
										assign node1563 = (inp[13]) ? node1583 : node1564;
											assign node1564 = (inp[5]) ? node1576 : node1565;
												assign node1565 = (inp[8]) ? node1567 : 16'b0001111111111111;
													assign node1567 = (inp[14]) ? 16'b0000011111111111 : node1568;
														assign node1568 = (inp[1]) ? 16'b0000011111111111 : node1569;
															assign node1569 = (inp[15]) ? node1571 : 16'b0000111111111111;
																assign node1571 = (inp[12]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node1576 = (inp[1]) ? node1580 : node1577;
													assign node1577 = (inp[15]) ? 16'b0000011111111111 : 16'b0000001111111111;
													assign node1580 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node1583 = (inp[8]) ? node1591 : node1584;
												assign node1584 = (inp[14]) ? node1586 : 16'b0000011111111111;
													assign node1586 = (inp[1]) ? node1588 : 16'b0000001111111111;
														assign node1588 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node1591 = (inp[5]) ? node1603 : node1592;
													assign node1592 = (inp[14]) ? 16'b0000000111111111 : node1593;
														assign node1593 = (inp[15]) ? node1595 : 16'b0000011111111111;
															assign node1595 = (inp[1]) ? node1599 : node1596;
																assign node1596 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
																assign node1599 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node1603 = (inp[1]) ? node1607 : node1604;
														assign node1604 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node1607 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node1610 = (inp[5]) ? node1640 : node1611;
											assign node1611 = (inp[12]) ? node1621 : node1612;
												assign node1612 = (inp[14]) ? 16'b0000001111111111 : node1613;
													assign node1613 = (inp[1]) ? node1615 : 16'b0000001111111111;
														assign node1615 = (inp[13]) ? node1617 : 16'b0000011111111111;
															assign node1617 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node1621 = (inp[15]) ? node1631 : node1622;
													assign node1622 = (inp[13]) ? node1628 : node1623;
														assign node1623 = (inp[1]) ? node1625 : 16'b0000011111111111;
															assign node1625 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node1628 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node1631 = (inp[1]) ? node1637 : node1632;
														assign node1632 = (inp[8]) ? node1634 : 16'b0000001111111111;
															assign node1634 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node1637 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node1640 = (inp[13]) ? 16'b0000000111111111 : node1641;
												assign node1641 = (inp[15]) ? node1643 : 16'b0000000111111111;
													assign node1643 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
								assign node1647 = (inp[8]) ? node1749 : node1648;
									assign node1648 = (inp[12]) ? node1704 : node1649;
										assign node1649 = (inp[9]) ? node1679 : node1650;
											assign node1650 = (inp[6]) ? node1674 : node1651;
												assign node1651 = (inp[1]) ? node1661 : node1652;
													assign node1652 = (inp[5]) ? node1656 : node1653;
														assign node1653 = (inp[13]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node1656 = (inp[13]) ? node1658 : 16'b0000111111111111;
															assign node1658 = (inp[15]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node1661 = (inp[14]) ? node1669 : node1662;
														assign node1662 = (inp[5]) ? node1664 : 16'b0000111111111111;
															assign node1664 = (inp[15]) ? 16'b0000011111111111 : node1665;
																assign node1665 = (inp[13]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node1669 = (inp[13]) ? node1671 : 16'b0000011111111111;
															assign node1671 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node1674 = (inp[5]) ? node1676 : 16'b0000011111111111;
													assign node1676 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node1679 = (inp[15]) ? node1695 : node1680;
												assign node1680 = (inp[14]) ? node1686 : node1681;
													assign node1681 = (inp[13]) ? 16'b0000001111111111 : node1682;
														assign node1682 = (inp[1]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node1686 = (inp[6]) ? node1690 : node1687;
														assign node1687 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node1690 = (inp[5]) ? node1692 : 16'b0000001111111111;
															assign node1692 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node1695 = (inp[14]) ? 16'b0000000111111111 : node1696;
													assign node1696 = (inp[13]) ? node1698 : 16'b0000001111111111;
														assign node1698 = (inp[1]) ? 16'b0000000011111111 : node1699;
															assign node1699 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node1704 = (inp[15]) ? node1728 : node1705;
											assign node1705 = (inp[13]) ? node1717 : node1706;
												assign node1706 = (inp[1]) ? node1708 : 16'b0000011111111111;
													assign node1708 = (inp[6]) ? node1714 : node1709;
														assign node1709 = (inp[14]) ? 16'b0000001111111111 : node1710;
															assign node1710 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node1714 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node1717 = (inp[5]) ? node1723 : node1718;
													assign node1718 = (inp[9]) ? 16'b0000001111111111 : node1719;
														assign node1719 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node1723 = (inp[14]) ? node1725 : 16'b0000000111111111;
														assign node1725 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node1728 = (inp[6]) ? node1734 : node1729;
												assign node1729 = (inp[13]) ? node1731 : 16'b0000001111111111;
													assign node1731 = (inp[5]) ? 16'b0000001111111111 : 16'b0000000111111111;
												assign node1734 = (inp[14]) ? node1740 : node1735;
													assign node1735 = (inp[1]) ? 16'b0000000111111111 : node1736;
														assign node1736 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node1740 = (inp[5]) ? node1742 : 16'b0000000111111111;
														assign node1742 = (inp[13]) ? 16'b0000000001111111 : node1743;
															assign node1743 = (inp[9]) ? node1745 : 16'b0000000011111111;
																assign node1745 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node1749 = (inp[5]) ? node1805 : node1750;
										assign node1750 = (inp[14]) ? node1780 : node1751;
											assign node1751 = (inp[9]) ? node1767 : node1752;
												assign node1752 = (inp[6]) ? node1760 : node1753;
													assign node1753 = (inp[13]) ? node1755 : 16'b0000111111111111;
														assign node1755 = (inp[15]) ? 16'b0000001111111111 : node1756;
															assign node1756 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node1760 = (inp[1]) ? node1762 : 16'b0000001111111111;
														assign node1762 = (inp[12]) ? 16'b0000001111111111 : node1763;
															assign node1763 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node1767 = (inp[12]) ? node1773 : node1768;
													assign node1768 = (inp[6]) ? 16'b0000001111111111 : node1769;
														assign node1769 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node1773 = (inp[1]) ? node1777 : node1774;
														assign node1774 = (inp[15]) ? 16'b0000001111111111 : 16'b0000000111111111;
														assign node1777 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node1780 = (inp[13]) ? node1792 : node1781;
												assign node1781 = (inp[6]) ? node1787 : node1782;
													assign node1782 = (inp[15]) ? 16'b0000001111111111 : node1783;
														assign node1783 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node1787 = (inp[9]) ? node1789 : 16'b0000000111111111;
														assign node1789 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node1792 = (inp[12]) ? node1800 : node1793;
													assign node1793 = (inp[6]) ? node1797 : node1794;
														assign node1794 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node1797 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node1800 = (inp[6]) ? 16'b0000000001111111 : node1801;
														assign node1801 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node1805 = (inp[1]) ? node1827 : node1806;
											assign node1806 = (inp[12]) ? node1818 : node1807;
												assign node1807 = (inp[13]) ? node1813 : node1808;
													assign node1808 = (inp[9]) ? node1810 : 16'b0000001111111111;
														assign node1810 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node1813 = (inp[15]) ? node1815 : 16'b0000000111111111;
														assign node1815 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node1818 = (inp[9]) ? 16'b0000000011111111 : node1819;
													assign node1819 = (inp[15]) ? node1823 : node1820;
														assign node1820 = (inp[13]) ? 16'b0000000111111111 : 16'b0000011111111111;
														assign node1823 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node1827 = (inp[13]) ? node1841 : node1828;
												assign node1828 = (inp[14]) ? node1834 : node1829;
													assign node1829 = (inp[12]) ? node1831 : 16'b0000000111111111;
														assign node1831 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node1834 = (inp[15]) ? node1836 : 16'b0000000111111111;
														assign node1836 = (inp[9]) ? node1838 : 16'b0000000011111111;
															assign node1838 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node1841 = (inp[6]) ? node1849 : node1842;
													assign node1842 = (inp[15]) ? node1846 : node1843;
														assign node1843 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node1846 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node1849 = (inp[14]) ? node1855 : node1850;
														assign node1850 = (inp[9]) ? 16'b0000000001111111 : node1851;
															assign node1851 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node1855 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000001111111;
							assign node1858 = (inp[1]) ? node2050 : node1859;
								assign node1859 = (inp[8]) ? node1963 : node1860;
									assign node1860 = (inp[13]) ? node1908 : node1861;
										assign node1861 = (inp[6]) ? node1887 : node1862;
											assign node1862 = (inp[2]) ? node1876 : node1863;
												assign node1863 = (inp[5]) ? node1873 : node1864;
													assign node1864 = (inp[12]) ? 16'b0000111111111111 : node1865;
														assign node1865 = (inp[14]) ? node1869 : node1866;
															assign node1866 = (inp[15]) ? 16'b0001111111111111 : 16'b0011111111111111;
															assign node1869 = (inp[15]) ? 16'b0000111111111111 : 16'b0001111111111111;
													assign node1873 = (inp[14]) ? 16'b0000001111111111 : 16'b0000111111111111;
												assign node1876 = (inp[14]) ? node1882 : node1877;
													assign node1877 = (inp[5]) ? 16'b0000001111111111 : node1878;
														assign node1878 = (inp[12]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node1882 = (inp[12]) ? node1884 : 16'b0000001111111111;
														assign node1884 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node1887 = (inp[15]) ? node1901 : node1888;
												assign node1888 = (inp[5]) ? node1896 : node1889;
													assign node1889 = (inp[2]) ? node1891 : 16'b0000011111111111;
														assign node1891 = (inp[12]) ? 16'b0000001111111111 : node1892;
															assign node1892 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node1896 = (inp[12]) ? 16'b0000001111111111 : node1897;
														assign node1897 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node1901 = (inp[14]) ? node1903 : 16'b0000001111111111;
													assign node1903 = (inp[5]) ? 16'b0000000011111111 : node1904;
														assign node1904 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node1908 = (inp[15]) ? node1930 : node1909;
											assign node1909 = (inp[2]) ? node1921 : node1910;
												assign node1910 = (inp[5]) ? node1916 : node1911;
													assign node1911 = (inp[14]) ? node1913 : 16'b0000011111111111;
														assign node1913 = (inp[12]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node1916 = (inp[6]) ? 16'b0000000111111111 : node1917;
														assign node1917 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node1921 = (inp[12]) ? node1925 : node1922;
													assign node1922 = (inp[6]) ? 16'b0000000111111111 : 16'b0000011111111111;
													assign node1925 = (inp[6]) ? node1927 : 16'b0000000111111111;
														assign node1927 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node1930 = (inp[9]) ? node1946 : node1931;
												assign node1931 = (inp[14]) ? node1933 : 16'b0000001111111111;
													assign node1933 = (inp[5]) ? node1939 : node1934;
														assign node1934 = (inp[6]) ? node1936 : 16'b0000001111111111;
															assign node1936 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node1939 = (inp[2]) ? node1941 : 16'b0000001111111111;
															assign node1941 = (inp[6]) ? 16'b0000000011111111 : node1942;
																assign node1942 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node1946 = (inp[5]) ? node1956 : node1947;
													assign node1947 = (inp[2]) ? node1951 : node1948;
														assign node1948 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node1951 = (inp[12]) ? node1953 : 16'b0000000111111111;
															assign node1953 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node1956 = (inp[6]) ? node1958 : 16'b0000000011111111;
														assign node1958 = (inp[14]) ? node1960 : 16'b0000000011111111;
															assign node1960 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node1963 = (inp[6]) ? node2005 : node1964;
										assign node1964 = (inp[15]) ? node1982 : node1965;
											assign node1965 = (inp[2]) ? node1975 : node1966;
												assign node1966 = (inp[9]) ? node1970 : node1967;
													assign node1967 = (inp[14]) ? 16'b0000011111111111 : 16'b0001111111111111;
													assign node1970 = (inp[14]) ? 16'b0000000111111111 : node1971;
														assign node1971 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node1975 = (inp[9]) ? node1977 : 16'b0000001111111111;
													assign node1977 = (inp[5]) ? 16'b0000000111111111 : node1978;
														assign node1978 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node1982 = (inp[2]) ? node1994 : node1983;
												assign node1983 = (inp[14]) ? node1989 : node1984;
													assign node1984 = (inp[12]) ? node1986 : 16'b0000011111111111;
														assign node1986 = (inp[13]) ? 16'b0000000011111111 : 16'b0000001111111111;
													assign node1989 = (inp[9]) ? 16'b0000000111111111 : node1990;
														assign node1990 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node1994 = (inp[9]) ? 16'b0000000011111111 : node1995;
													assign node1995 = (inp[12]) ? node1997 : 16'b0000001111111111;
														assign node1997 = (inp[14]) ? node1999 : 16'b0000000111111111;
															assign node1999 = (inp[13]) ? 16'b0000000011111111 : node2000;
																assign node2000 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node2005 = (inp[14]) ? node2029 : node2006;
											assign node2006 = (inp[5]) ? node2020 : node2007;
												assign node2007 = (inp[9]) ? node2017 : node2008;
													assign node2008 = (inp[13]) ? 16'b0000000111111111 : node2009;
														assign node2009 = (inp[2]) ? node2011 : 16'b0000001111111111;
															assign node2011 = (inp[12]) ? node2013 : 16'b0000001111111111;
																assign node2013 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node2017 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node2020 = (inp[15]) ? node2022 : 16'b0000000111111111;
													assign node2022 = (inp[2]) ? 16'b0000000011111111 : node2023;
														assign node2023 = (inp[13]) ? node2025 : 16'b0000000111111111;
															assign node2025 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000111111111;
											assign node2029 = (inp[13]) ? node2045 : node2030;
												assign node2030 = (inp[5]) ? node2036 : node2031;
													assign node2031 = (inp[9]) ? 16'b0000000011111111 : node2032;
														assign node2032 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node2036 = (inp[12]) ? 16'b0000000011111111 : node2037;
														assign node2037 = (inp[9]) ? node2039 : 16'b0000000111111111;
															assign node2039 = (inp[2]) ? 16'b0000000011111111 : node2040;
																assign node2040 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node2045 = (inp[9]) ? node2047 : 16'b0000000011111111;
													assign node2047 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
								assign node2050 = (inp[9]) ? node2156 : node2051;
									assign node2051 = (inp[6]) ? node2099 : node2052;
										assign node2052 = (inp[2]) ? node2078 : node2053;
											assign node2053 = (inp[5]) ? node2067 : node2054;
												assign node2054 = (inp[8]) ? node2062 : node2055;
													assign node2055 = (inp[14]) ? 16'b0000111111111111 : node2056;
														assign node2056 = (inp[13]) ? 16'b0000111111111111 : node2057;
															assign node2057 = (inp[15]) ? 16'b0000111111111111 : 16'b0001111111111111;
													assign node2062 = (inp[15]) ? 16'b0000000111111111 : node2063;
														assign node2063 = (inp[12]) ? 16'b0000011111111111 : 16'b0000001111111111;
												assign node2067 = (inp[13]) ? node2073 : node2068;
													assign node2068 = (inp[14]) ? 16'b0000001111111111 : node2069;
														assign node2069 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node2073 = (inp[12]) ? 16'b0000000111111111 : node2074;
														assign node2074 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node2078 = (inp[5]) ? node2088 : node2079;
												assign node2079 = (inp[14]) ? node2083 : node2080;
													assign node2080 = (inp[12]) ? 16'b0000001111111111 : 16'b0000111111111111;
													assign node2083 = (inp[15]) ? 16'b0000000111111111 : node2084;
														assign node2084 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node2088 = (inp[12]) ? node2094 : node2089;
													assign node2089 = (inp[13]) ? node2091 : 16'b0000001111111111;
														assign node2091 = (inp[8]) ? 16'b0000000111111111 : 16'b0000000011111111;
													assign node2094 = (inp[8]) ? 16'b0000000011111111 : node2095;
														assign node2095 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node2099 = (inp[8]) ? node2133 : node2100;
											assign node2100 = (inp[13]) ? node2116 : node2101;
												assign node2101 = (inp[2]) ? node2109 : node2102;
													assign node2102 = (inp[15]) ? node2106 : node2103;
														assign node2103 = (inp[12]) ? 16'b0000001111111111 : 16'b0000111111111111;
														assign node2106 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node2109 = (inp[15]) ? node2113 : node2110;
														assign node2110 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node2113 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node2116 = (inp[5]) ? node2124 : node2117;
													assign node2117 = (inp[14]) ? node2121 : node2118;
														assign node2118 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node2121 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node2124 = (inp[2]) ? node2130 : node2125;
														assign node2125 = (inp[15]) ? node2127 : 16'b0000000111111111;
															assign node2127 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node2130 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node2133 = (inp[13]) ? node2151 : node2134;
												assign node2134 = (inp[2]) ? node2142 : node2135;
													assign node2135 = (inp[14]) ? node2139 : node2136;
														assign node2136 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node2139 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node2142 = (inp[5]) ? node2146 : node2143;
														assign node2143 = (inp[12]) ? 16'b0000000111111111 : 16'b0000000011111111;
														assign node2146 = (inp[15]) ? node2148 : 16'b0000000001111111;
															assign node2148 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node2151 = (inp[14]) ? 16'b0000000001111111 : node2152;
													assign node2152 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node2156 = (inp[14]) ? node2202 : node2157;
										assign node2157 = (inp[12]) ? node2185 : node2158;
											assign node2158 = (inp[13]) ? node2170 : node2159;
												assign node2159 = (inp[15]) ? 16'b0000000111111111 : node2160;
													assign node2160 = (inp[6]) ? 16'b0000000111111111 : node2161;
														assign node2161 = (inp[5]) ? node2165 : node2162;
															assign node2162 = (inp[2]) ? 16'b0000011111111111 : 16'b0000111111111111;
															assign node2165 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node2170 = (inp[8]) ? node2180 : node2171;
													assign node2171 = (inp[5]) ? node2177 : node2172;
														assign node2172 = (inp[15]) ? 16'b0000000111111111 : node2173;
															assign node2173 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node2177 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node2180 = (inp[6]) ? 16'b0000000011111111 : node2181;
														assign node2181 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000111111111;
											assign node2185 = (inp[15]) ? node2191 : node2186;
												assign node2186 = (inp[8]) ? 16'b0000000011111111 : node2187;
													assign node2187 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node2191 = (inp[6]) ? node2197 : node2192;
													assign node2192 = (inp[8]) ? node2194 : 16'b0000000011111111;
														assign node2194 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000111111111;
													assign node2197 = (inp[5]) ? 16'b0000000000111111 : node2198;
														assign node2198 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node2202 = (inp[5]) ? node2234 : node2203;
											assign node2203 = (inp[2]) ? node2221 : node2204;
												assign node2204 = (inp[6]) ? node2210 : node2205;
													assign node2205 = (inp[12]) ? node2207 : 16'b0000000011111111;
														assign node2207 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node2210 = (inp[15]) ? node2216 : node2211;
														assign node2211 = (inp[13]) ? node2213 : 16'b0000000111111111;
															assign node2213 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node2216 = (inp[8]) ? 16'b0000000011111111 : node2217;
															assign node2217 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node2221 = (inp[6]) ? node2227 : node2222;
													assign node2222 = (inp[13]) ? node2224 : 16'b0000000011111111;
														assign node2224 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node2227 = (inp[15]) ? node2229 : 16'b0000000001111111;
														assign node2229 = (inp[12]) ? 16'b0000000000111111 : node2230;
															assign node2230 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node2234 = (inp[15]) ? node2246 : node2235;
												assign node2235 = (inp[6]) ? node2243 : node2236;
													assign node2236 = (inp[2]) ? node2238 : 16'b0000000111111111;
														assign node2238 = (inp[12]) ? node2240 : 16'b0000000011111111;
															assign node2240 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node2243 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000000111111;
												assign node2246 = (inp[8]) ? node2252 : node2247;
													assign node2247 = (inp[2]) ? node2249 : 16'b0000000001111111;
														assign node2249 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node2252 = (inp[12]) ? node2254 : 16'b0000000001111111;
														assign node2254 = (inp[2]) ? 16'b0000000000011111 : node2255;
															assign node2255 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
						assign node2259 = (inp[1]) ? node2601 : node2260;
							assign node2260 = (inp[12]) ? node2424 : node2261;
								assign node2261 = (inp[9]) ? node2347 : node2262;
									assign node2262 = (inp[8]) ? node2296 : node2263;
										assign node2263 = (inp[6]) ? node2285 : node2264;
											assign node2264 = (inp[2]) ? node2278 : node2265;
												assign node2265 = (inp[4]) ? node2269 : node2266;
													assign node2266 = (inp[14]) ? 16'b0000111111111111 : 16'b0001111111111111;
													assign node2269 = (inp[15]) ? node2275 : node2270;
														assign node2270 = (inp[13]) ? node2272 : 16'b0000111111111111;
															assign node2272 = (inp[14]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node2275 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node2278 = (inp[13]) ? node2280 : 16'b0000011111111111;
													assign node2280 = (inp[14]) ? 16'b0000001111111111 : node2281;
														assign node2281 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node2285 = (inp[4]) ? node2291 : node2286;
												assign node2286 = (inp[5]) ? 16'b0000011111111111 : node2287;
													assign node2287 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node2291 = (inp[5]) ? node2293 : 16'b0000001111111111;
													assign node2293 = (inp[15]) ? 16'b0000000011111111 : 16'b0000001111111111;
										assign node2296 = (inp[15]) ? node2320 : node2297;
											assign node2297 = (inp[14]) ? node2307 : node2298;
												assign node2298 = (inp[5]) ? node2300 : 16'b0000011111111111;
													assign node2300 = (inp[4]) ? 16'b0000001111111111 : node2301;
														assign node2301 = (inp[2]) ? 16'b0000001111111111 : node2302;
															assign node2302 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node2307 = (inp[6]) ? node2313 : node2308;
													assign node2308 = (inp[5]) ? node2310 : 16'b0000001111111111;
														assign node2310 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node2313 = (inp[4]) ? 16'b0000000011111111 : node2314;
														assign node2314 = (inp[13]) ? 16'b0000000111111111 : node2315;
															assign node2315 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node2320 = (inp[6]) ? node2342 : node2321;
												assign node2321 = (inp[2]) ? node2333 : node2322;
													assign node2322 = (inp[5]) ? node2328 : node2323;
														assign node2323 = (inp[4]) ? 16'b0000001111111111 : node2324;
															assign node2324 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node2328 = (inp[14]) ? 16'b0000000111111111 : node2329;
															assign node2329 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node2333 = (inp[13]) ? node2339 : node2334;
														assign node2334 = (inp[14]) ? 16'b0000000111111111 : node2335;
															assign node2335 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node2339 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node2342 = (inp[14]) ? node2344 : 16'b0000000111111111;
													assign node2344 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node2347 = (inp[4]) ? node2387 : node2348;
										assign node2348 = (inp[13]) ? node2370 : node2349;
											assign node2349 = (inp[6]) ? node2355 : node2350;
												assign node2350 = (inp[5]) ? 16'b0000001111111111 : node2351;
													assign node2351 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node2355 = (inp[2]) ? node2363 : node2356;
													assign node2356 = (inp[8]) ? node2360 : node2357;
														assign node2357 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node2360 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node2363 = (inp[8]) ? 16'b0000000011111111 : node2364;
														assign node2364 = (inp[14]) ? 16'b0000000111111111 : node2365;
															assign node2365 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node2370 = (inp[8]) ? node2378 : node2371;
												assign node2371 = (inp[14]) ? node2373 : 16'b0000001111111111;
													assign node2373 = (inp[15]) ? 16'b0000000111111111 : node2374;
														assign node2374 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node2378 = (inp[15]) ? node2384 : node2379;
													assign node2379 = (inp[6]) ? node2381 : 16'b0000000111111111;
														assign node2381 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node2384 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node2387 = (inp[13]) ? node2411 : node2388;
											assign node2388 = (inp[14]) ? node2400 : node2389;
												assign node2389 = (inp[2]) ? node2391 : 16'b0000001111111111;
													assign node2391 = (inp[5]) ? node2395 : node2392;
														assign node2392 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node2395 = (inp[15]) ? node2397 : 16'b0000000111111111;
															assign node2397 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node2400 = (inp[6]) ? node2406 : node2401;
													assign node2401 = (inp[8]) ? node2403 : 16'b0000001111111111;
														assign node2403 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node2406 = (inp[2]) ? node2408 : 16'b0000000011111111;
														assign node2408 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node2411 = (inp[15]) ? node2419 : node2412;
												assign node2412 = (inp[6]) ? node2416 : node2413;
													assign node2413 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node2416 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node2419 = (inp[14]) ? 16'b0000000001111111 : node2420;
													assign node2420 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
								assign node2424 = (inp[4]) ? node2508 : node2425;
									assign node2425 = (inp[6]) ? node2467 : node2426;
										assign node2426 = (inp[13]) ? node2448 : node2427;
											assign node2427 = (inp[14]) ? node2437 : node2428;
												assign node2428 = (inp[2]) ? node2434 : node2429;
													assign node2429 = (inp[9]) ? 16'b0000011111111111 : node2430;
														assign node2430 = (inp[5]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node2434 = (inp[15]) ? 16'b0000000111111111 : 16'b0000011111111111;
												assign node2437 = (inp[9]) ? node2439 : 16'b0000001111111111;
													assign node2439 = (inp[8]) ? 16'b0000000111111111 : node2440;
														assign node2440 = (inp[15]) ? 16'b0000000111111111 : node2441;
															assign node2441 = (inp[5]) ? 16'b0000001111111111 : node2442;
																assign node2442 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node2448 = (inp[5]) ? node2460 : node2449;
												assign node2449 = (inp[8]) ? node2455 : node2450;
													assign node2450 = (inp[9]) ? 16'b0000001111111111 : node2451;
														assign node2451 = (inp[15]) ? 16'b0000000111111111 : 16'b0000011111111111;
													assign node2455 = (inp[2]) ? 16'b0000000011111111 : node2456;
														assign node2456 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node2460 = (inp[9]) ? node2462 : 16'b0000000111111111;
													assign node2462 = (inp[15]) ? node2464 : 16'b0000000011111111;
														assign node2464 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node2467 = (inp[14]) ? node2495 : node2468;
											assign node2468 = (inp[8]) ? node2482 : node2469;
												assign node2469 = (inp[2]) ? node2479 : node2470;
													assign node2470 = (inp[13]) ? node2476 : node2471;
														assign node2471 = (inp[5]) ? 16'b0000001111111111 : node2472;
															assign node2472 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node2476 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node2479 = (inp[13]) ? 16'b0000000111111111 : 16'b0000000011111111;
												assign node2482 = (inp[5]) ? node2490 : node2483;
													assign node2483 = (inp[13]) ? node2487 : node2484;
														assign node2484 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node2487 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node2490 = (inp[2]) ? 16'b0000000011111111 : node2491;
														assign node2491 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node2495 = (inp[15]) ? node2501 : node2496;
												assign node2496 = (inp[2]) ? 16'b0000000011111111 : node2497;
													assign node2497 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node2501 = (inp[2]) ? 16'b0000000001111111 : node2502;
													assign node2502 = (inp[13]) ? node2504 : 16'b0000000011111111;
														assign node2504 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node2508 = (inp[8]) ? node2560 : node2509;
										assign node2509 = (inp[13]) ? node2527 : node2510;
											assign node2510 = (inp[2]) ? node2520 : node2511;
												assign node2511 = (inp[5]) ? 16'b0000000111111111 : node2512;
													assign node2512 = (inp[9]) ? node2514 : 16'b0000001111111111;
														assign node2514 = (inp[6]) ? node2516 : 16'b0000001111111111;
															assign node2516 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node2520 = (inp[5]) ? node2522 : 16'b0000000111111111;
													assign node2522 = (inp[6]) ? 16'b0000000011111111 : node2523;
														assign node2523 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node2527 = (inp[15]) ? node2545 : node2528;
												assign node2528 = (inp[6]) ? node2536 : node2529;
													assign node2529 = (inp[9]) ? node2533 : node2530;
														assign node2530 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node2533 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node2536 = (inp[9]) ? 16'b0000000011111111 : node2537;
														assign node2537 = (inp[14]) ? node2539 : 16'b0000000111111111;
															assign node2539 = (inp[2]) ? 16'b0000000011111111 : node2540;
																assign node2540 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node2545 = (inp[2]) ? node2553 : node2546;
													assign node2546 = (inp[6]) ? node2550 : node2547;
														assign node2547 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node2550 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node2553 = (inp[6]) ? node2557 : node2554;
														assign node2554 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node2557 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node2560 = (inp[15]) ? node2582 : node2561;
											assign node2561 = (inp[13]) ? node2571 : node2562;
												assign node2562 = (inp[9]) ? node2564 : 16'b0000000111111111;
													assign node2564 = (inp[6]) ? 16'b0000000011111111 : node2565;
														assign node2565 = (inp[5]) ? 16'b0000000011111111 : node2566;
															assign node2566 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node2571 = (inp[2]) ? node2573 : 16'b0000000011111111;
													assign node2573 = (inp[14]) ? node2577 : node2574;
														assign node2574 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node2577 = (inp[6]) ? node2579 : 16'b0000000001111111;
															assign node2579 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node2582 = (inp[9]) ? node2590 : node2583;
												assign node2583 = (inp[5]) ? 16'b0000000001111111 : node2584;
													assign node2584 = (inp[6]) ? node2586 : 16'b0000000011111111;
														assign node2586 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node2590 = (inp[6]) ? node2596 : node2591;
													assign node2591 = (inp[14]) ? node2593 : 16'b0000000001111111;
														assign node2593 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node2596 = (inp[13]) ? 16'b0000000000011111 : node2597;
														assign node2597 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000011111111;
							assign node2601 = (inp[4]) ? node2783 : node2602;
								assign node2602 = (inp[12]) ? node2690 : node2603;
									assign node2603 = (inp[9]) ? node2649 : node2604;
										assign node2604 = (inp[8]) ? node2628 : node2605;
											assign node2605 = (inp[6]) ? node2617 : node2606;
												assign node2606 = (inp[14]) ? node2614 : node2607;
													assign node2607 = (inp[5]) ? 16'b0000011111111111 : node2608;
														assign node2608 = (inp[2]) ? 16'b0000111111111111 : node2609;
															assign node2609 = (inp[13]) ? 16'b0000111111111111 : 16'b0001111111111111;
													assign node2614 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node2617 = (inp[13]) ? node2619 : 16'b0000011111111111;
													assign node2619 = (inp[15]) ? 16'b0000000111111111 : node2620;
														assign node2620 = (inp[5]) ? 16'b0000000111111111 : node2621;
															assign node2621 = (inp[2]) ? 16'b0000001111111111 : node2622;
																assign node2622 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node2628 = (inp[2]) ? node2638 : node2629;
												assign node2629 = (inp[5]) ? node2633 : node2630;
													assign node2630 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node2633 = (inp[14]) ? 16'b0000000111111111 : node2634;
														assign node2634 = (inp[15]) ? 16'b0000000111111111 : 16'b0000011111111111;
												assign node2638 = (inp[5]) ? node2644 : node2639;
													assign node2639 = (inp[6]) ? 16'b0000000011111111 : node2640;
														assign node2640 = (inp[13]) ? 16'b0000001111111111 : 16'b0000000111111111;
													assign node2644 = (inp[14]) ? 16'b0000000011111111 : node2645;
														assign node2645 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node2649 = (inp[6]) ? node2667 : node2650;
											assign node2650 = (inp[8]) ? node2662 : node2651;
												assign node2651 = (inp[15]) ? node2657 : node2652;
													assign node2652 = (inp[5]) ? 16'b0000001111111111 : node2653;
														assign node2653 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node2657 = (inp[14]) ? node2659 : 16'b0000000011111111;
														assign node2659 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node2662 = (inp[2]) ? 16'b0000000011111111 : node2663;
													assign node2663 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node2667 = (inp[13]) ? node2683 : node2668;
												assign node2668 = (inp[5]) ? node2676 : node2669;
													assign node2669 = (inp[8]) ? node2671 : 16'b0000000111111111;
														assign node2671 = (inp[2]) ? node2673 : 16'b0000000111111111;
															assign node2673 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node2676 = (inp[14]) ? 16'b0000000001111111 : node2677;
														assign node2677 = (inp[8]) ? 16'b0000000011111111 : node2678;
															assign node2678 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node2683 = (inp[5]) ? 16'b0000000001111111 : node2684;
													assign node2684 = (inp[2]) ? node2686 : 16'b0000000011111111;
														assign node2686 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node2690 = (inp[15]) ? node2722 : node2691;
										assign node2691 = (inp[5]) ? node2707 : node2692;
											assign node2692 = (inp[8]) ? node2700 : node2693;
												assign node2693 = (inp[13]) ? node2695 : 16'b0000001111111111;
													assign node2695 = (inp[14]) ? 16'b0000000111111111 : node2696;
														assign node2696 = (inp[2]) ? 16'b0000001111111111 : 16'b0000000111111111;
												assign node2700 = (inp[13]) ? 16'b0000000011111111 : node2701;
													assign node2701 = (inp[2]) ? 16'b0000000011111111 : node2702;
														assign node2702 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node2707 = (inp[2]) ? node2715 : node2708;
												assign node2708 = (inp[13]) ? 16'b0000000011111111 : node2709;
													assign node2709 = (inp[6]) ? node2711 : 16'b0000000111111111;
														assign node2711 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node2715 = (inp[9]) ? node2717 : 16'b0000000011111111;
													assign node2717 = (inp[8]) ? 16'b0000000001111111 : node2718;
														assign node2718 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node2722 = (inp[5]) ? node2756 : node2723;
											assign node2723 = (inp[2]) ? node2735 : node2724;
												assign node2724 = (inp[8]) ? node2730 : node2725;
													assign node2725 = (inp[13]) ? 16'b0000000111111111 : node2726;
														assign node2726 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node2730 = (inp[9]) ? node2732 : 16'b0000000011111111;
														assign node2732 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node2735 = (inp[6]) ? node2745 : node2736;
													assign node2736 = (inp[9]) ? 16'b0000000001111111 : node2737;
														assign node2737 = (inp[14]) ? 16'b0000000011111111 : node2738;
															assign node2738 = (inp[8]) ? node2740 : 16'b0000000111111111;
																assign node2740 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node2745 = (inp[8]) ? node2753 : node2746;
														assign node2746 = (inp[9]) ? node2748 : 16'b0000000011111111;
															assign node2748 = (inp[14]) ? 16'b0000000001111111 : node2749;
																assign node2749 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node2753 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node2756 = (inp[9]) ? node2764 : node2757;
												assign node2757 = (inp[6]) ? 16'b0000000001111111 : node2758;
													assign node2758 = (inp[13]) ? node2760 : 16'b0000000011111111;
														assign node2760 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node2764 = (inp[6]) ? node2776 : node2765;
													assign node2765 = (inp[2]) ? node2769 : node2766;
														assign node2766 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node2769 = (inp[13]) ? node2771 : 16'b0000000001111111;
															assign node2771 = (inp[14]) ? 16'b0000000000111111 : node2772;
																assign node2772 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node2776 = (inp[8]) ? 16'b0000000000011111 : node2777;
														assign node2777 = (inp[13]) ? 16'b0000000000111111 : node2778;
															assign node2778 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
								assign node2783 = (inp[6]) ? node2865 : node2784;
									assign node2784 = (inp[13]) ? node2818 : node2785;
										assign node2785 = (inp[8]) ? node2803 : node2786;
											assign node2786 = (inp[12]) ? node2794 : node2787;
												assign node2787 = (inp[5]) ? node2791 : node2788;
													assign node2788 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node2791 = (inp[2]) ? 16'b0000000011111111 : 16'b0000001111111111;
												assign node2794 = (inp[14]) ? node2800 : node2795;
													assign node2795 = (inp[5]) ? node2797 : 16'b0000000111111111;
														assign node2797 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node2800 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node2803 = (inp[14]) ? node2813 : node2804;
												assign node2804 = (inp[2]) ? node2808 : node2805;
													assign node2805 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node2808 = (inp[5]) ? node2810 : 16'b0000000011111111;
														assign node2810 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node2813 = (inp[2]) ? node2815 : 16'b0000000011111111;
													assign node2815 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node2818 = (inp[5]) ? node2846 : node2819;
											assign node2819 = (inp[14]) ? node2831 : node2820;
												assign node2820 = (inp[12]) ? node2826 : node2821;
													assign node2821 = (inp[15]) ? 16'b0000000111111111 : node2822;
														assign node2822 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node2826 = (inp[15]) ? 16'b0000000011111111 : node2827;
														assign node2827 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node2831 = (inp[8]) ? node2841 : node2832;
													assign node2832 = (inp[15]) ? node2836 : node2833;
														assign node2833 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node2836 = (inp[12]) ? node2838 : 16'b0000000011111111;
															assign node2838 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node2841 = (inp[9]) ? node2843 : 16'b0000000001111111;
														assign node2843 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000001111111;
											assign node2846 = (inp[12]) ? node2858 : node2847;
												assign node2847 = (inp[9]) ? node2849 : 16'b0000000011111111;
													assign node2849 = (inp[14]) ? node2855 : node2850;
														assign node2850 = (inp[2]) ? 16'b0000000001111111 : node2851;
															assign node2851 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000111111111;
														assign node2855 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node2858 = (inp[9]) ? 16'b0000000000111111 : node2859;
													assign node2859 = (inp[14]) ? node2861 : 16'b0000000001111111;
														assign node2861 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000000111111;
									assign node2865 = (inp[2]) ? node2903 : node2866;
										assign node2866 = (inp[13]) ? node2882 : node2867;
											assign node2867 = (inp[8]) ? node2879 : node2868;
												assign node2868 = (inp[5]) ? node2874 : node2869;
													assign node2869 = (inp[12]) ? node2871 : 16'b0000000111111111;
														assign node2871 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node2874 = (inp[15]) ? node2876 : 16'b0000000011111111;
														assign node2876 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node2879 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node2882 = (inp[8]) ? node2894 : node2883;
												assign node2883 = (inp[12]) ? 16'b0000000001111111 : node2884;
													assign node2884 = (inp[14]) ? node2886 : 16'b0000000111111111;
														assign node2886 = (inp[9]) ? 16'b0000000001111111 : node2887;
															assign node2887 = (inp[15]) ? node2889 : 16'b0000000011111111;
																assign node2889 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node2894 = (inp[14]) ? node2898 : node2895;
													assign node2895 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node2898 = (inp[5]) ? 16'b0000000000111111 : node2899;
														assign node2899 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node2903 = (inp[13]) ? node2933 : node2904;
											assign node2904 = (inp[14]) ? node2918 : node2905;
												assign node2905 = (inp[12]) ? node2911 : node2906;
													assign node2906 = (inp[9]) ? 16'b0000000011111111 : node2907;
														assign node2907 = (inp[15]) ? 16'b0000000011111111 : 16'b0000001111111111;
													assign node2911 = (inp[5]) ? node2913 : 16'b0000000011111111;
														assign node2913 = (inp[9]) ? 16'b0000000000111111 : node2914;
															assign node2914 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node2918 = (inp[8]) ? node2926 : node2919;
													assign node2919 = (inp[12]) ? node2921 : 16'b0000000001111111;
														assign node2921 = (inp[5]) ? 16'b0000000000011111 : node2922;
															assign node2922 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node2926 = (inp[9]) ? node2928 : 16'b0000000000111111;
														assign node2928 = (inp[15]) ? node2930 : 16'b0000000000011111;
															assign node2930 = (inp[12]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node2933 = (inp[15]) ? node2941 : node2934;
												assign node2934 = (inp[14]) ? 16'b0000000000111111 : node2935;
													assign node2935 = (inp[8]) ? 16'b0000000000111111 : node2936;
														assign node2936 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node2941 = (inp[12]) ? 16'b0000000000011111 : node2942;
													assign node2942 = (inp[5]) ? node2952 : node2943;
														assign node2943 = (inp[9]) ? node2947 : node2944;
															assign node2944 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
															assign node2947 = (inp[14]) ? node2949 : 16'b0000000000111111;
																assign node2949 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node2952 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
				assign node2956 = (inp[10]) ? node4352 : node2957;
					assign node2957 = (inp[13]) ? node3681 : node2958;
						assign node2958 = (inp[14]) ? node3340 : node2959;
							assign node2959 = (inp[6]) ? node3147 : node2960;
								assign node2960 = (inp[5]) ? node3052 : node2961;
									assign node2961 = (inp[0]) ? node3007 : node2962;
										assign node2962 = (inp[8]) ? node2982 : node2963;
											assign node2963 = (inp[9]) ? node2971 : node2964;
												assign node2964 = (inp[2]) ? 16'b0000111111111111 : node2965;
													assign node2965 = (inp[15]) ? 16'b0001111111111111 : node2966;
														assign node2966 = (inp[12]) ? 16'b0001111111111111 : 16'b0011111111111111;
												assign node2971 = (inp[1]) ? node2977 : node2972;
													assign node2972 = (inp[12]) ? 16'b0000111111111111 : node2973;
														assign node2973 = (inp[4]) ? 16'b0000111111111111 : 16'b0001111111111111;
													assign node2977 = (inp[12]) ? node2979 : 16'b0000111111111111;
														assign node2979 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node2982 = (inp[4]) ? node2994 : node2983;
												assign node2983 = (inp[12]) ? 16'b0000011111111111 : node2984;
													assign node2984 = (inp[15]) ? node2990 : node2985;
														assign node2985 = (inp[9]) ? 16'b0000111111111111 : node2986;
															assign node2986 = (inp[2]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node2990 = (inp[2]) ? 16'b0000111111111111 : 16'b0000011111111111;
												assign node2994 = (inp[9]) ? node3002 : node2995;
													assign node2995 = (inp[1]) ? 16'b0000011111111111 : node2996;
														assign node2996 = (inp[15]) ? node2998 : 16'b0000111111111111;
															assign node2998 = (inp[12]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node3002 = (inp[15]) ? node3004 : 16'b0000011111111111;
														assign node3004 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node3007 = (inp[8]) ? node3033 : node3008;
											assign node3008 = (inp[9]) ? node3026 : node3009;
												assign node3009 = (inp[4]) ? node3021 : node3010;
													assign node3010 = (inp[12]) ? node3018 : node3011;
														assign node3011 = (inp[2]) ? node3013 : 16'b0001111111111111;
															assign node3013 = (inp[15]) ? 16'b0000111111111111 : node3014;
																assign node3014 = (inp[1]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node3018 = (inp[15]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node3021 = (inp[2]) ? 16'b0000001111111111 : node3022;
														assign node3022 = (inp[15]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node3026 = (inp[1]) ? node3028 : 16'b0000011111111111;
													assign node3028 = (inp[15]) ? node3030 : 16'b0000001111111111;
														assign node3030 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node3033 = (inp[2]) ? node3041 : node3034;
												assign node3034 = (inp[4]) ? node3036 : 16'b0000011111111111;
													assign node3036 = (inp[9]) ? 16'b0000000111111111 : node3037;
														assign node3037 = (inp[1]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node3041 = (inp[1]) ? node3047 : node3042;
													assign node3042 = (inp[12]) ? node3044 : 16'b0000111111111111;
														assign node3044 = (inp[15]) ? 16'b0000001111111111 : 16'b0000000111111111;
													assign node3047 = (inp[12]) ? 16'b0000000011111111 : node3048;
														assign node3048 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
									assign node3052 = (inp[15]) ? node3100 : node3053;
										assign node3053 = (inp[2]) ? node3089 : node3054;
											assign node3054 = (inp[4]) ? node3070 : node3055;
												assign node3055 = (inp[0]) ? node3065 : node3056;
													assign node3056 = (inp[9]) ? node3062 : node3057;
														assign node3057 = (inp[12]) ? 16'b0000111111111111 : node3058;
															assign node3058 = (inp[1]) ? 16'b0001111111111111 : 16'b0011111111111111;
														assign node3062 = (inp[8]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node3065 = (inp[9]) ? 16'b0000011111111111 : node3066;
														assign node3066 = (inp[1]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node3070 = (inp[8]) ? node3076 : node3071;
													assign node3071 = (inp[9]) ? node3073 : 16'b0000011111111111;
														assign node3073 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node3076 = (inp[0]) ? node3082 : node3077;
														assign node3077 = (inp[12]) ? node3079 : 16'b0000011111111111;
															assign node3079 = (inp[1]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node3082 = (inp[1]) ? 16'b0000001111111111 : node3083;
															assign node3083 = (inp[9]) ? 16'b0000001111111111 : node3084;
																assign node3084 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node3089 = (inp[0]) ? node3095 : node3090;
												assign node3090 = (inp[12]) ? 16'b0000001111111111 : node3091;
													assign node3091 = (inp[1]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node3095 = (inp[4]) ? node3097 : 16'b0000001111111111;
													assign node3097 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000111111111;
										assign node3100 = (inp[1]) ? node3120 : node3101;
											assign node3101 = (inp[9]) ? node3113 : node3102;
												assign node3102 = (inp[4]) ? node3108 : node3103;
													assign node3103 = (inp[0]) ? 16'b0000011111111111 : node3104;
														assign node3104 = (inp[12]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node3108 = (inp[2]) ? node3110 : 16'b0000011111111111;
														assign node3110 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node3113 = (inp[4]) ? 16'b0000000111111111 : node3114;
													assign node3114 = (inp[2]) ? node3116 : 16'b0000011111111111;
														assign node3116 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node3120 = (inp[0]) ? node3138 : node3121;
												assign node3121 = (inp[4]) ? node3129 : node3122;
													assign node3122 = (inp[12]) ? 16'b0000000111111111 : node3123;
														assign node3123 = (inp[9]) ? node3125 : 16'b0000011111111111;
															assign node3125 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node3129 = (inp[9]) ? node3131 : 16'b0000001111111111;
														assign node3131 = (inp[12]) ? 16'b0000000011111111 : node3132;
															assign node3132 = (inp[8]) ? node3134 : 16'b0000000111111111;
																assign node3134 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node3138 = (inp[2]) ? node3140 : 16'b0000000111111111;
													assign node3140 = (inp[8]) ? 16'b0000000011111111 : node3141;
														assign node3141 = (inp[12]) ? node3143 : 16'b0000000111111111;
															assign node3143 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
								assign node3147 = (inp[2]) ? node3241 : node3148;
									assign node3148 = (inp[12]) ? node3192 : node3149;
										assign node3149 = (inp[4]) ? node3175 : node3150;
											assign node3150 = (inp[1]) ? node3166 : node3151;
												assign node3151 = (inp[5]) ? node3161 : node3152;
													assign node3152 = (inp[8]) ? node3154 : 16'b0000111111111111;
														assign node3154 = (inp[15]) ? node3156 : 16'b0000111111111111;
															assign node3156 = (inp[9]) ? 16'b0000011111111111 : node3157;
																assign node3157 = (inp[0]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node3161 = (inp[8]) ? 16'b0000001111111111 : node3162;
														assign node3162 = (inp[0]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node3166 = (inp[15]) ? node3172 : node3167;
													assign node3167 = (inp[9]) ? node3169 : 16'b0000011111111111;
														assign node3169 = (inp[0]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node3172 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node3175 = (inp[0]) ? node3183 : node3176;
												assign node3176 = (inp[9]) ? 16'b0000001111111111 : node3177;
													assign node3177 = (inp[15]) ? node3179 : 16'b0000011111111111;
														assign node3179 = (inp[1]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node3183 = (inp[9]) ? node3185 : 16'b0000001111111111;
													assign node3185 = (inp[15]) ? 16'b0000000111111111 : node3186;
														assign node3186 = (inp[1]) ? 16'b0000000111111111 : node3187;
															assign node3187 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
										assign node3192 = (inp[15]) ? node3212 : node3193;
											assign node3193 = (inp[5]) ? node3205 : node3194;
												assign node3194 = (inp[0]) ? node3198 : node3195;
													assign node3195 = (inp[9]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node3198 = (inp[1]) ? 16'b0000001111111111 : node3199;
														assign node3199 = (inp[9]) ? node3201 : 16'b0000011111111111;
															assign node3201 = (inp[4]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node3205 = (inp[9]) ? node3207 : 16'b0000001111111111;
													assign node3207 = (inp[0]) ? 16'b0000000111111111 : node3208;
														assign node3208 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node3212 = (inp[0]) ? node3224 : node3213;
												assign node3213 = (inp[4]) ? node3219 : node3214;
													assign node3214 = (inp[1]) ? node3216 : 16'b0000011111111111;
														assign node3216 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node3219 = (inp[8]) ? 16'b0000000111111111 : node3220;
														assign node3220 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node3224 = (inp[4]) ? node3236 : node3225;
													assign node3225 = (inp[8]) ? 16'b0000000011111111 : node3226;
														assign node3226 = (inp[1]) ? node3232 : node3227;
															assign node3227 = (inp[9]) ? node3229 : 16'b0000001111111111;
																assign node3229 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
															assign node3232 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node3236 = (inp[1]) ? 16'b0000000011111111 : node3237;
														assign node3237 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node3241 = (inp[1]) ? node3285 : node3242;
										assign node3242 = (inp[4]) ? node3266 : node3243;
											assign node3243 = (inp[8]) ? node3255 : node3244;
												assign node3244 = (inp[5]) ? node3252 : node3245;
													assign node3245 = (inp[12]) ? node3249 : node3246;
														assign node3246 = (inp[15]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node3249 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node3252 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node3255 = (inp[0]) ? 16'b0000000111111111 : node3256;
													assign node3256 = (inp[9]) ? node3260 : node3257;
														assign node3257 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node3260 = (inp[5]) ? 16'b0000000111111111 : node3261;
															assign node3261 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node3266 = (inp[9]) ? node3276 : node3267;
												assign node3267 = (inp[15]) ? node3271 : node3268;
													assign node3268 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node3271 = (inp[12]) ? node3273 : 16'b0000001111111111;
														assign node3273 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node3276 = (inp[12]) ? node3278 : 16'b0000000111111111;
													assign node3278 = (inp[0]) ? node3282 : node3279;
														assign node3279 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node3282 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node3285 = (inp[12]) ? node3321 : node3286;
											assign node3286 = (inp[8]) ? node3298 : node3287;
												assign node3287 = (inp[4]) ? node3291 : node3288;
													assign node3288 = (inp[0]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node3291 = (inp[0]) ? 16'b0000000111111111 : node3292;
														assign node3292 = (inp[15]) ? node3294 : 16'b0000001111111111;
															assign node3294 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node3298 = (inp[4]) ? node3314 : node3299;
													assign node3299 = (inp[5]) ? node3311 : node3300;
														assign node3300 = (inp[9]) ? node3306 : node3301;
															assign node3301 = (inp[0]) ? node3303 : 16'b0000001111111111;
																assign node3303 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
															assign node3306 = (inp[15]) ? 16'b0000000111111111 : node3307;
																assign node3307 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node3311 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node3314 = (inp[15]) ? node3318 : node3315;
														assign node3315 = (inp[5]) ? 16'b0000000111111111 : 16'b0000000011111111;
														assign node3318 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node3321 = (inp[8]) ? node3327 : node3322;
												assign node3322 = (inp[5]) ? 16'b0000000011111111 : node3323;
													assign node3323 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node3327 = (inp[9]) ? node3333 : node3328;
													assign node3328 = (inp[15]) ? node3330 : 16'b0000000111111111;
														assign node3330 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node3333 = (inp[5]) ? node3335 : 16'b0000000001111111;
														assign node3335 = (inp[15]) ? 16'b0000000000111111 : node3336;
															assign node3336 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
							assign node3340 = (inp[5]) ? node3506 : node3341;
								assign node3341 = (inp[9]) ? node3425 : node3342;
									assign node3342 = (inp[12]) ? node3382 : node3343;
										assign node3343 = (inp[0]) ? node3365 : node3344;
											assign node3344 = (inp[1]) ? node3356 : node3345;
												assign node3345 = (inp[6]) ? node3347 : 16'b0000111111111111;
													assign node3347 = (inp[4]) ? 16'b0000011111111111 : node3348;
														assign node3348 = (inp[15]) ? node3350 : 16'b0000111111111111;
															assign node3350 = (inp[2]) ? node3352 : 16'b0000111111111111;
																assign node3352 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node3356 = (inp[8]) ? 16'b0000001111111111 : node3357;
													assign node3357 = (inp[6]) ? 16'b0000001111111111 : node3358;
														assign node3358 = (inp[15]) ? 16'b0000011111111111 : node3359;
															assign node3359 = (inp[2]) ? 16'b0000011111111111 : 16'b0000111111111111;
											assign node3365 = (inp[15]) ? node3373 : node3366;
												assign node3366 = (inp[8]) ? node3368 : 16'b0000011111111111;
													assign node3368 = (inp[2]) ? 16'b0000011111111111 : node3369;
														assign node3369 = (inp[4]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node3373 = (inp[1]) ? node3379 : node3374;
													assign node3374 = (inp[2]) ? node3376 : 16'b0000001111111111;
														assign node3376 = (inp[6]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node3379 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node3382 = (inp[2]) ? node3398 : node3383;
											assign node3383 = (inp[8]) ? node3387 : node3384;
												assign node3384 = (inp[4]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node3387 = (inp[15]) ? node3393 : node3388;
													assign node3388 = (inp[6]) ? 16'b0000001111111111 : node3389;
														assign node3389 = (inp[0]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node3393 = (inp[6]) ? 16'b0000000111111111 : node3394;
														assign node3394 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node3398 = (inp[8]) ? node3414 : node3399;
												assign node3399 = (inp[1]) ? node3407 : node3400;
													assign node3400 = (inp[0]) ? node3404 : node3401;
														assign node3401 = (inp[15]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node3404 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node3407 = (inp[15]) ? node3411 : node3408;
														assign node3408 = (inp[6]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node3411 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node3414 = (inp[6]) ? node3420 : node3415;
													assign node3415 = (inp[4]) ? 16'b0000000111111111 : node3416;
														assign node3416 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node3420 = (inp[1]) ? node3422 : 16'b0000000011111111;
														assign node3422 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node3425 = (inp[15]) ? node3469 : node3426;
										assign node3426 = (inp[0]) ? node3444 : node3427;
											assign node3427 = (inp[6]) ? node3439 : node3428;
												assign node3428 = (inp[2]) ? node3434 : node3429;
													assign node3429 = (inp[4]) ? 16'b0000011111111111 : node3430;
														assign node3430 = (inp[8]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node3434 = (inp[4]) ? node3436 : 16'b0000011111111111;
														assign node3436 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node3439 = (inp[8]) ? node3441 : 16'b0000001111111111;
													assign node3441 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node3444 = (inp[1]) ? node3464 : node3445;
												assign node3445 = (inp[2]) ? node3455 : node3446;
													assign node3446 = (inp[8]) ? node3448 : 16'b0000011111111111;
														assign node3448 = (inp[12]) ? 16'b0000001111111111 : node3449;
															assign node3449 = (inp[4]) ? 16'b0000001111111111 : node3450;
																assign node3450 = (inp[6]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node3455 = (inp[4]) ? node3457 : 16'b0000000111111111;
														assign node3457 = (inp[6]) ? node3459 : 16'b0000000111111111;
															assign node3459 = (inp[8]) ? 16'b0000000011111111 : node3460;
																assign node3460 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node3464 = (inp[4]) ? node3466 : 16'b0000000011111111;
													assign node3466 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node3469 = (inp[4]) ? node3487 : node3470;
											assign node3470 = (inp[6]) ? node3480 : node3471;
												assign node3471 = (inp[2]) ? 16'b0000000011111111 : node3472;
													assign node3472 = (inp[0]) ? 16'b0000001111111111 : node3473;
														assign node3473 = (inp[8]) ? node3475 : 16'b0000001111111111;
															assign node3475 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node3480 = (inp[12]) ? node3482 : 16'b0000000111111111;
													assign node3482 = (inp[1]) ? 16'b0000000011111111 : node3483;
														assign node3483 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node3487 = (inp[8]) ? node3497 : node3488;
												assign node3488 = (inp[1]) ? 16'b0000000001111111 : node3489;
													assign node3489 = (inp[6]) ? node3491 : 16'b0000000111111111;
														assign node3491 = (inp[0]) ? node3493 : 16'b0000000111111111;
															assign node3493 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node3497 = (inp[2]) ? node3499 : 16'b0000000001111111;
													assign node3499 = (inp[6]) ? 16'b0000000000111111 : node3500;
														assign node3500 = (inp[0]) ? node3502 : 16'b0000000011111111;
															assign node3502 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
								assign node3506 = (inp[2]) ? node3594 : node3507;
									assign node3507 = (inp[8]) ? node3563 : node3508;
										assign node3508 = (inp[0]) ? node3532 : node3509;
											assign node3509 = (inp[1]) ? node3525 : node3510;
												assign node3510 = (inp[4]) ? node3516 : node3511;
													assign node3511 = (inp[15]) ? 16'b0000001111111111 : node3512;
														assign node3512 = (inp[6]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node3516 = (inp[12]) ? node3518 : 16'b0000001111111111;
														assign node3518 = (inp[9]) ? 16'b0000000111111111 : node3519;
															assign node3519 = (inp[15]) ? node3521 : 16'b0000001111111111;
																assign node3521 = (inp[6]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node3525 = (inp[9]) ? 16'b0000000111111111 : node3526;
													assign node3526 = (inp[12]) ? 16'b0000000111111111 : node3527;
														assign node3527 = (inp[6]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node3532 = (inp[6]) ? node3550 : node3533;
												assign node3533 = (inp[4]) ? node3539 : node3534;
													assign node3534 = (inp[15]) ? node3536 : 16'b0000111111111111;
														assign node3536 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node3539 = (inp[15]) ? node3545 : node3540;
														assign node3540 = (inp[12]) ? node3542 : 16'b0000001111111111;
															assign node3542 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node3545 = (inp[1]) ? node3547 : 16'b0000000111111111;
															assign node3547 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node3550 = (inp[1]) ? node3558 : node3551;
													assign node3551 = (inp[4]) ? node3553 : 16'b0000000111111111;
														assign node3553 = (inp[9]) ? node3555 : 16'b0000000111111111;
															assign node3555 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node3558 = (inp[12]) ? node3560 : 16'b0000000011111111;
														assign node3560 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node3563 = (inp[4]) ? node3575 : node3564;
											assign node3564 = (inp[15]) ? node3568 : node3565;
												assign node3565 = (inp[6]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node3568 = (inp[1]) ? 16'b0000000011111111 : node3569;
													assign node3569 = (inp[6]) ? node3571 : 16'b0000000111111111;
														assign node3571 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000111111111;
											assign node3575 = (inp[15]) ? node3589 : node3576;
												assign node3576 = (inp[6]) ? node3582 : node3577;
													assign node3577 = (inp[12]) ? 16'b0000000011111111 : node3578;
														assign node3578 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node3582 = (inp[1]) ? node3584 : 16'b0000000011111111;
														assign node3584 = (inp[12]) ? 16'b0000000001111111 : node3585;
															assign node3585 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node3589 = (inp[12]) ? 16'b0000000001111111 : node3590;
													assign node3590 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node3594 = (inp[1]) ? node3642 : node3595;
										assign node3595 = (inp[12]) ? node3617 : node3596;
											assign node3596 = (inp[8]) ? node3608 : node3597;
												assign node3597 = (inp[4]) ? node3601 : node3598;
													assign node3598 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node3601 = (inp[9]) ? 16'b0000000111111111 : node3602;
														assign node3602 = (inp[6]) ? node3604 : 16'b0000001111111111;
															assign node3604 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node3608 = (inp[15]) ? node3610 : 16'b0000000111111111;
													assign node3610 = (inp[6]) ? node3614 : node3611;
														assign node3611 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node3614 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node3617 = (inp[15]) ? node3631 : node3618;
												assign node3618 = (inp[8]) ? node3626 : node3619;
													assign node3619 = (inp[6]) ? 16'b0000000011111111 : node3620;
														assign node3620 = (inp[4]) ? node3622 : 16'b0000000111111111;
															assign node3622 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node3626 = (inp[4]) ? node3628 : 16'b0000000011111111;
														assign node3628 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node3631 = (inp[6]) ? 16'b0000000001111111 : node3632;
													assign node3632 = (inp[9]) ? node3634 : 16'b0000000111111111;
														assign node3634 = (inp[0]) ? 16'b0000000001111111 : node3635;
															assign node3635 = (inp[8]) ? node3637 : 16'b0000000011111111;
																assign node3637 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node3642 = (inp[6]) ? node3660 : node3643;
											assign node3643 = (inp[12]) ? node3647 : node3644;
												assign node3644 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node3647 = (inp[4]) ? node3653 : node3648;
													assign node3648 = (inp[15]) ? node3650 : 16'b0000000011111111;
														assign node3650 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node3653 = (inp[9]) ? 16'b0000000000111111 : node3654;
														assign node3654 = (inp[15]) ? 16'b0000000001111111 : node3655;
															assign node3655 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node3660 = (inp[12]) ? node3670 : node3661;
												assign node3661 = (inp[0]) ? node3667 : node3662;
													assign node3662 = (inp[15]) ? node3664 : 16'b0000000111111111;
														assign node3664 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node3667 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node3670 = (inp[15]) ? node3678 : node3671;
													assign node3671 = (inp[8]) ? node3673 : 16'b0000000001111111;
														assign node3673 = (inp[0]) ? node3675 : 16'b0000000001111111;
															assign node3675 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node3678 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000000011111;
						assign node3681 = (inp[15]) ? node4035 : node3682;
							assign node3682 = (inp[9]) ? node3850 : node3683;
								assign node3683 = (inp[0]) ? node3775 : node3684;
									assign node3684 = (inp[1]) ? node3742 : node3685;
										assign node3685 = (inp[6]) ? node3717 : node3686;
											assign node3686 = (inp[12]) ? node3704 : node3687;
												assign node3687 = (inp[8]) ? node3695 : node3688;
													assign node3688 = (inp[5]) ? 16'b0000111111111111 : node3689;
														assign node3689 = (inp[14]) ? node3691 : 16'b0001111111111111;
															assign node3691 = (inp[2]) ? 16'b0000111111111111 : 16'b0001111111111111;
													assign node3695 = (inp[14]) ? 16'b0000001111111111 : node3696;
														assign node3696 = (inp[2]) ? node3698 : 16'b0000111111111111;
															assign node3698 = (inp[5]) ? 16'b0000011111111111 : node3699;
																assign node3699 = (inp[4]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node3704 = (inp[5]) ? node3712 : node3705;
													assign node3705 = (inp[4]) ? node3709 : node3706;
														assign node3706 = (inp[8]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node3709 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node3712 = (inp[4]) ? 16'b0000000111111111 : node3713;
														assign node3713 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node3717 = (inp[8]) ? node3727 : node3718;
												assign node3718 = (inp[2]) ? node3722 : node3719;
													assign node3719 = (inp[14]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node3722 = (inp[14]) ? node3724 : 16'b0000011111111111;
														assign node3724 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node3727 = (inp[12]) ? node3733 : node3728;
													assign node3728 = (inp[14]) ? 16'b0000001111111111 : node3729;
														assign node3729 = (inp[4]) ? 16'b0000011111111111 : 16'b0000001111111111;
													assign node3733 = (inp[5]) ? 16'b0000000111111111 : node3734;
														assign node3734 = (inp[4]) ? node3736 : 16'b0000001111111111;
															assign node3736 = (inp[14]) ? 16'b0000000111111111 : node3737;
																assign node3737 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node3742 = (inp[4]) ? node3758 : node3743;
											assign node3743 = (inp[5]) ? node3751 : node3744;
												assign node3744 = (inp[2]) ? node3748 : node3745;
													assign node3745 = (inp[8]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node3748 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node3751 = (inp[8]) ? 16'b0000000111111111 : node3752;
													assign node3752 = (inp[6]) ? 16'b0000001111111111 : node3753;
														assign node3753 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node3758 = (inp[12]) ? node3764 : node3759;
												assign node3759 = (inp[8]) ? node3761 : 16'b0000001111111111;
													assign node3761 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node3764 = (inp[6]) ? node3770 : node3765;
													assign node3765 = (inp[5]) ? 16'b0000000001111111 : node3766;
														assign node3766 = (inp[2]) ? 16'b0000001111111111 : 16'b0000000111111111;
													assign node3770 = (inp[2]) ? 16'b0000000011111111 : node3771;
														assign node3771 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node3775 = (inp[14]) ? node3815 : node3776;
										assign node3776 = (inp[5]) ? node3798 : node3777;
											assign node3777 = (inp[4]) ? node3787 : node3778;
												assign node3778 = (inp[2]) ? node3780 : 16'b0000111111111111;
													assign node3780 = (inp[8]) ? 16'b0000000111111111 : node3781;
														assign node3781 = (inp[1]) ? node3783 : 16'b0000011111111111;
															assign node3783 = (inp[6]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node3787 = (inp[2]) ? node3795 : node3788;
													assign node3788 = (inp[8]) ? node3790 : 16'b0000011111111111;
														assign node3790 = (inp[6]) ? node3792 : 16'b0000001111111111;
															assign node3792 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node3795 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node3798 = (inp[8]) ? node3808 : node3799;
												assign node3799 = (inp[12]) ? node3803 : node3800;
													assign node3800 = (inp[4]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node3803 = (inp[4]) ? node3805 : 16'b0000000111111111;
														assign node3805 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node3808 = (inp[1]) ? node3810 : 16'b0000000111111111;
													assign node3810 = (inp[4]) ? node3812 : 16'b0000000011111111;
														assign node3812 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node3815 = (inp[6]) ? node3831 : node3816;
											assign node3816 = (inp[1]) ? node3824 : node3817;
												assign node3817 = (inp[12]) ? 16'b0000000111111111 : node3818;
													assign node3818 = (inp[4]) ? node3820 : 16'b0000011111111111;
														assign node3820 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node3824 = (inp[5]) ? 16'b0000000011111111 : node3825;
													assign node3825 = (inp[4]) ? node3827 : 16'b0000000111111111;
														assign node3827 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node3831 = (inp[12]) ? node3839 : node3832;
												assign node3832 = (inp[2]) ? 16'b0000000011111111 : node3833;
													assign node3833 = (inp[4]) ? 16'b0000000011111111 : node3834;
														assign node3834 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node3839 = (inp[2]) ? node3845 : node3840;
													assign node3840 = (inp[5]) ? node3842 : 16'b0000000011111111;
														assign node3842 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node3845 = (inp[1]) ? node3847 : 16'b0000000001111111;
														assign node3847 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
								assign node3850 = (inp[4]) ? node3948 : node3851;
									assign node3851 = (inp[5]) ? node3899 : node3852;
										assign node3852 = (inp[2]) ? node3880 : node3853;
											assign node3853 = (inp[1]) ? node3867 : node3854;
												assign node3854 = (inp[8]) ? node3864 : node3855;
													assign node3855 = (inp[6]) ? 16'b0000011111111111 : node3856;
														assign node3856 = (inp[14]) ? 16'b0000011111111111 : node3857;
															assign node3857 = (inp[0]) ? node3859 : 16'b0000111111111111;
																assign node3859 = (inp[12]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node3864 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node3867 = (inp[0]) ? node3875 : node3868;
													assign node3868 = (inp[12]) ? 16'b0000001111111111 : node3869;
														assign node3869 = (inp[8]) ? node3871 : 16'b0000011111111111;
															assign node3871 = (inp[6]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node3875 = (inp[8]) ? 16'b0000000011111111 : node3876;
														assign node3876 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node3880 = (inp[1]) ? node3892 : node3881;
												assign node3881 = (inp[6]) ? node3885 : node3882;
													assign node3882 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node3885 = (inp[8]) ? node3887 : 16'b0000000111111111;
														assign node3887 = (inp[14]) ? node3889 : 16'b0000000111111111;
															assign node3889 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node3892 = (inp[8]) ? node3894 : 16'b0000000111111111;
													assign node3894 = (inp[0]) ? node3896 : 16'b0000000111111111;
														assign node3896 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node3899 = (inp[0]) ? node3919 : node3900;
											assign node3900 = (inp[1]) ? node3910 : node3901;
												assign node3901 = (inp[6]) ? node3907 : node3902;
													assign node3902 = (inp[14]) ? node3904 : 16'b0000001111111111;
														assign node3904 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node3907 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node3910 = (inp[8]) ? node3916 : node3911;
													assign node3911 = (inp[6]) ? node3913 : 16'b0000000111111111;
														assign node3913 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node3916 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000111111111;
											assign node3919 = (inp[6]) ? node3929 : node3920;
												assign node3920 = (inp[1]) ? node3924 : node3921;
													assign node3921 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node3924 = (inp[12]) ? node3926 : 16'b0000000011111111;
														assign node3926 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000011111111;
												assign node3929 = (inp[14]) ? node3941 : node3930;
													assign node3930 = (inp[2]) ? node3936 : node3931;
														assign node3931 = (inp[1]) ? node3933 : 16'b0000000011111111;
															assign node3933 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node3936 = (inp[8]) ? 16'b0000000001111111 : node3937;
															assign node3937 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node3941 = (inp[2]) ? node3943 : 16'b0000000001111111;
														assign node3943 = (inp[1]) ? 16'b0000000000111111 : node3944;
															assign node3944 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node3948 = (inp[2]) ? node3978 : node3949;
										assign node3949 = (inp[1]) ? node3965 : node3950;
											assign node3950 = (inp[14]) ? node3960 : node3951;
												assign node3951 = (inp[12]) ? 16'b0000000111111111 : node3952;
													assign node3952 = (inp[8]) ? 16'b0000000011111111 : node3953;
														assign node3953 = (inp[6]) ? node3955 : 16'b0000011111111111;
															assign node3955 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node3960 = (inp[5]) ? 16'b0000000011111111 : node3961;
													assign node3961 = (inp[12]) ? 16'b0000000111111111 : 16'b0000000011111111;
											assign node3965 = (inp[0]) ? node3973 : node3966;
												assign node3966 = (inp[6]) ? node3968 : 16'b0000000111111111;
													assign node3968 = (inp[5]) ? node3970 : 16'b0000000111111111;
														assign node3970 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node3973 = (inp[14]) ? node3975 : 16'b0000000001111111;
													assign node3975 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000001111111;
										assign node3978 = (inp[12]) ? node4006 : node3979;
											assign node3979 = (inp[5]) ? node3989 : node3980;
												assign node3980 = (inp[0]) ? node3986 : node3981;
													assign node3981 = (inp[1]) ? node3983 : 16'b0000000111111111;
														assign node3983 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node3986 = (inp[8]) ? 16'b0000000111111111 : 16'b0000000011111111;
												assign node3989 = (inp[6]) ? node3995 : node3990;
													assign node3990 = (inp[8]) ? node3992 : 16'b0000000111111111;
														assign node3992 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000001111111;
													assign node3995 = (inp[14]) ? node4001 : node3996;
														assign node3996 = (inp[0]) ? 16'b0000000001111111 : node3997;
															assign node3997 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000111111111;
														assign node4001 = (inp[0]) ? node4003 : 16'b0000000001111111;
															assign node4003 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node4006 = (inp[1]) ? node4020 : node4007;
												assign node4007 = (inp[5]) ? node4011 : node4008;
													assign node4008 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node4011 = (inp[8]) ? node4017 : node4012;
														assign node4012 = (inp[0]) ? 16'b0000000001111111 : node4013;
															assign node4013 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node4017 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node4020 = (inp[5]) ? node4032 : node4021;
													assign node4021 = (inp[0]) ? node4023 : 16'b0000000001111111;
														assign node4023 = (inp[14]) ? node4029 : node4024;
															assign node4024 = (inp[8]) ? node4026 : 16'b0000000001111111;
																assign node4026 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
															assign node4029 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node4032 = (inp[6]) ? 16'b0000000000011111 : 16'b0000000000111111;
							assign node4035 = (inp[2]) ? node4183 : node4036;
								assign node4036 = (inp[14]) ? node4116 : node4037;
									assign node4037 = (inp[4]) ? node4079 : node4038;
										assign node4038 = (inp[0]) ? node4060 : node4039;
											assign node4039 = (inp[8]) ? node4051 : node4040;
												assign node4040 = (inp[5]) ? node4046 : node4041;
													assign node4041 = (inp[1]) ? node4043 : 16'b0000011111111111;
														assign node4043 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node4046 = (inp[9]) ? 16'b0000000111111111 : node4047;
														assign node4047 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node4051 = (inp[5]) ? node4057 : node4052;
													assign node4052 = (inp[9]) ? node4054 : 16'b0000001111111111;
														assign node4054 = (inp[6]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node4057 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node4060 = (inp[9]) ? node4070 : node4061;
												assign node4061 = (inp[5]) ? node4067 : node4062;
													assign node4062 = (inp[1]) ? node4064 : 16'b0000001111111111;
														assign node4064 = (inp[6]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node4067 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node4070 = (inp[6]) ? node4076 : node4071;
													assign node4071 = (inp[1]) ? 16'b0000000011111111 : node4072;
														assign node4072 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node4076 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node4079 = (inp[1]) ? node4097 : node4080;
											assign node4080 = (inp[12]) ? node4088 : node4081;
												assign node4081 = (inp[0]) ? node4083 : 16'b0000001111111111;
													assign node4083 = (inp[9]) ? node4085 : 16'b0000000111111111;
														assign node4085 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node4088 = (inp[5]) ? node4092 : node4089;
													assign node4089 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node4092 = (inp[9]) ? 16'b0000000011111111 : node4093;
														assign node4093 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node4097 = (inp[5]) ? node4105 : node4098;
												assign node4098 = (inp[12]) ? node4100 : 16'b0000000111111111;
													assign node4100 = (inp[9]) ? node4102 : 16'b0000000111111111;
														assign node4102 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node4105 = (inp[6]) ? node4107 : 16'b0000000011111111;
													assign node4107 = (inp[12]) ? node4113 : node4108;
														assign node4108 = (inp[0]) ? 16'b0000000001111111 : node4109;
															assign node4109 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node4113 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node4116 = (inp[6]) ? node4150 : node4117;
										assign node4117 = (inp[12]) ? node4129 : node4118;
											assign node4118 = (inp[0]) ? node4126 : node4119;
												assign node4119 = (inp[1]) ? 16'b0000000111111111 : node4120;
													assign node4120 = (inp[4]) ? node4122 : 16'b0000011111111111;
														assign node4122 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node4126 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node4129 = (inp[9]) ? node4139 : node4130;
												assign node4130 = (inp[5]) ? node4132 : 16'b0000000111111111;
													assign node4132 = (inp[0]) ? node4136 : node4133;
														assign node4133 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node4136 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node4139 = (inp[8]) ? node4145 : node4140;
													assign node4140 = (inp[4]) ? 16'b0000000011111111 : node4141;
														assign node4141 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node4145 = (inp[4]) ? 16'b0000000000111111 : node4146;
														assign node4146 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node4150 = (inp[4]) ? node4166 : node4151;
											assign node4151 = (inp[9]) ? node4159 : node4152;
												assign node4152 = (inp[5]) ? node4154 : 16'b0000000111111111;
													assign node4154 = (inp[8]) ? node4156 : 16'b0000001111111111;
														assign node4156 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node4159 = (inp[12]) ? 16'b0000000001111111 : node4160;
													assign node4160 = (inp[0]) ? node4162 : 16'b0000000011111111;
														assign node4162 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node4166 = (inp[0]) ? node4176 : node4167;
												assign node4167 = (inp[12]) ? node4169 : 16'b0000000011111111;
													assign node4169 = (inp[8]) ? node4171 : 16'b0000000011111111;
														assign node4171 = (inp[5]) ? 16'b0000000000111111 : node4172;
															assign node4172 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node4176 = (inp[8]) ? node4178 : 16'b0000000001111111;
													assign node4178 = (inp[12]) ? node4180 : 16'b0000000001111111;
														assign node4180 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
								assign node4183 = (inp[6]) ? node4267 : node4184;
									assign node4184 = (inp[4]) ? node4224 : node4185;
										assign node4185 = (inp[5]) ? node4201 : node4186;
											assign node4186 = (inp[9]) ? node4194 : node4187;
												assign node4187 = (inp[0]) ? 16'b0000000111111111 : node4188;
													assign node4188 = (inp[1]) ? node4190 : 16'b0000011111111111;
														assign node4190 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node4194 = (inp[14]) ? 16'b0000000011111111 : node4195;
													assign node4195 = (inp[1]) ? node4197 : 16'b0000000111111111;
														assign node4197 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000111111111;
											assign node4201 = (inp[14]) ? node4213 : node4202;
												assign node4202 = (inp[9]) ? node4210 : node4203;
													assign node4203 = (inp[1]) ? node4205 : 16'b0000001111111111;
														assign node4205 = (inp[12]) ? node4207 : 16'b0000000111111111;
															assign node4207 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node4210 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node4213 = (inp[1]) ? node4219 : node4214;
													assign node4214 = (inp[9]) ? 16'b0000000011111111 : node4215;
														assign node4215 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node4219 = (inp[12]) ? node4221 : 16'b0000000011111111;
														assign node4221 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node4224 = (inp[12]) ? node4250 : node4225;
											assign node4225 = (inp[5]) ? node4237 : node4226;
												assign node4226 = (inp[1]) ? node4232 : node4227;
													assign node4227 = (inp[8]) ? 16'b0000000011111111 : node4228;
														assign node4228 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node4232 = (inp[14]) ? 16'b0000000011111111 : node4233;
														assign node4233 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node4237 = (inp[9]) ? node4245 : node4238;
													assign node4238 = (inp[1]) ? 16'b0000000001111111 : node4239;
														assign node4239 = (inp[0]) ? 16'b0000000011111111 : node4240;
															assign node4240 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node4245 = (inp[8]) ? 16'b0000000000111111 : node4246;
														assign node4246 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node4250 = (inp[1]) ? node4258 : node4251;
												assign node4251 = (inp[0]) ? 16'b0000000001111111 : node4252;
													assign node4252 = (inp[14]) ? 16'b0000000001111111 : node4253;
														assign node4253 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node4258 = (inp[9]) ? node4262 : node4259;
													assign node4259 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000001111111;
													assign node4262 = (inp[0]) ? 16'b0000000000111111 : node4263;
														assign node4263 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node4267 = (inp[8]) ? node4307 : node4268;
										assign node4268 = (inp[4]) ? node4288 : node4269;
											assign node4269 = (inp[12]) ? node4281 : node4270;
												assign node4270 = (inp[9]) ? node4274 : node4271;
													assign node4271 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node4274 = (inp[5]) ? node4278 : node4275;
														assign node4275 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node4278 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node4281 = (inp[14]) ? node4283 : 16'b0000000011111111;
													assign node4283 = (inp[1]) ? 16'b0000000001111111 : node4284;
														assign node4284 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node4288 = (inp[9]) ? node4302 : node4289;
												assign node4289 = (inp[1]) ? node4295 : node4290;
													assign node4290 = (inp[14]) ? 16'b0000000001111111 : node4291;
														assign node4291 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node4295 = (inp[0]) ? node4299 : node4296;
														assign node4296 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node4299 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node4302 = (inp[0]) ? node4304 : 16'b0000000001111111;
													assign node4304 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node4307 = (inp[14]) ? node4331 : node4308;
											assign node4308 = (inp[9]) ? node4316 : node4309;
												assign node4309 = (inp[12]) ? 16'b0000000001111111 : node4310;
													assign node4310 = (inp[4]) ? node4312 : 16'b0000000111111111;
														assign node4312 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node4316 = (inp[1]) ? node4320 : node4317;
													assign node4317 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node4320 = (inp[4]) ? node4328 : node4321;
														assign node4321 = (inp[12]) ? 16'b0000000000111111 : node4322;
															assign node4322 = (inp[0]) ? node4324 : 16'b0000000001111111;
																assign node4324 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node4328 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node4331 = (inp[9]) ? node4341 : node4332;
												assign node4332 = (inp[4]) ? node4338 : node4333;
													assign node4333 = (inp[0]) ? 16'b0000000000111111 : node4334;
														assign node4334 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node4338 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000000011111;
												assign node4341 = (inp[1]) ? node4343 : 16'b0000000000111111;
													assign node4343 = (inp[0]) ? node4347 : node4344;
														assign node4344 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node4347 = (inp[12]) ? 16'b0000000000001111 : node4348;
															assign node4348 = (inp[4]) ? 16'b0000000000011111 : 16'b0000000000111111;
					assign node4352 = (inp[2]) ? node5156 : node4353;
						assign node4353 = (inp[5]) ? node4733 : node4354;
							assign node4354 = (inp[9]) ? node4552 : node4355;
								assign node4355 = (inp[14]) ? node4453 : node4356;
									assign node4356 = (inp[12]) ? node4406 : node4357;
										assign node4357 = (inp[6]) ? node4379 : node4358;
											assign node4358 = (inp[1]) ? node4372 : node4359;
												assign node4359 = (inp[13]) ? node4365 : node4360;
													assign node4360 = (inp[8]) ? 16'b0000111111111111 : node4361;
														assign node4361 = (inp[0]) ? 16'b0000111111111111 : 16'b0011111111111111;
													assign node4365 = (inp[4]) ? 16'b0000011111111111 : node4366;
														assign node4366 = (inp[15]) ? 16'b0000011111111111 : node4367;
															assign node4367 = (inp[8]) ? 16'b0000111111111111 : 16'b0001111111111111;
												assign node4372 = (inp[15]) ? node4374 : 16'b0000011111111111;
													assign node4374 = (inp[4]) ? 16'b0000001111111111 : node4375;
														assign node4375 = (inp[0]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node4379 = (inp[13]) ? node4389 : node4380;
												assign node4380 = (inp[4]) ? node4384 : node4381;
													assign node4381 = (inp[1]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node4384 = (inp[0]) ? 16'b0000001111111111 : node4385;
														assign node4385 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node4389 = (inp[0]) ? node4397 : node4390;
													assign node4390 = (inp[4]) ? node4394 : node4391;
														assign node4391 = (inp[1]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node4394 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node4397 = (inp[1]) ? node4401 : node4398;
														assign node4398 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node4401 = (inp[4]) ? node4403 : 16'b0000000111111111;
															assign node4403 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node4406 = (inp[13]) ? node4442 : node4407;
											assign node4407 = (inp[8]) ? node4423 : node4408;
												assign node4408 = (inp[4]) ? node4416 : node4409;
													assign node4409 = (inp[15]) ? node4413 : node4410;
														assign node4410 = (inp[1]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node4413 = (inp[6]) ? 16'b0000011111111111 : 16'b0000001111111111;
													assign node4416 = (inp[0]) ? node4418 : 16'b0000011111111111;
														assign node4418 = (inp[15]) ? node4420 : 16'b0000001111111111;
															assign node4420 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node4423 = (inp[0]) ? node4429 : node4424;
													assign node4424 = (inp[4]) ? node4426 : 16'b0000001111111111;
														assign node4426 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node4429 = (inp[1]) ? node4433 : node4430;
														assign node4430 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node4433 = (inp[6]) ? node4437 : node4434;
															assign node4434 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
															assign node4437 = (inp[15]) ? 16'b0000000011111111 : node4438;
																assign node4438 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node4442 = (inp[1]) ? node4450 : node4443;
												assign node4443 = (inp[15]) ? 16'b0000000111111111 : node4444;
													assign node4444 = (inp[8]) ? 16'b0000000111111111 : node4445;
														assign node4445 = (inp[0]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node4450 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node4453 = (inp[12]) ? node4501 : node4454;
										assign node4454 = (inp[8]) ? node4482 : node4455;
											assign node4455 = (inp[4]) ? node4469 : node4456;
												assign node4456 = (inp[13]) ? node4460 : node4457;
													assign node4457 = (inp[6]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node4460 = (inp[0]) ? node4466 : node4461;
														assign node4461 = (inp[1]) ? 16'b0000001111111111 : node4462;
															assign node4462 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node4466 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node4469 = (inp[6]) ? node4477 : node4470;
													assign node4470 = (inp[13]) ? node4474 : node4471;
														assign node4471 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node4474 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node4477 = (inp[0]) ? 16'b0000000111111111 : node4478;
														assign node4478 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node4482 = (inp[15]) ? node4490 : node4483;
												assign node4483 = (inp[1]) ? node4485 : 16'b0000001111111111;
													assign node4485 = (inp[6]) ? 16'b0000000111111111 : node4486;
														assign node4486 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node4490 = (inp[13]) ? node4492 : 16'b0000000111111111;
													assign node4492 = (inp[0]) ? 16'b0000000011111111 : node4493;
														assign node4493 = (inp[4]) ? node4495 : 16'b0000000111111111;
															assign node4495 = (inp[1]) ? 16'b0000000011111111 : node4496;
																assign node4496 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node4501 = (inp[15]) ? node4529 : node4502;
											assign node4502 = (inp[13]) ? node4512 : node4503;
												assign node4503 = (inp[4]) ? node4507 : node4504;
													assign node4504 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node4507 = (inp[8]) ? 16'b0000000111111111 : node4508;
														assign node4508 = (inp[6]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node4512 = (inp[1]) ? node4522 : node4513;
													assign node4513 = (inp[4]) ? node4515 : 16'b0000000111111111;
														assign node4515 = (inp[8]) ? node4517 : 16'b0000000111111111;
															assign node4517 = (inp[6]) ? 16'b0000000011111111 : node4518;
																assign node4518 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node4522 = (inp[0]) ? 16'b0000000001111111 : node4523;
														assign node4523 = (inp[8]) ? 16'b0000000011111111 : node4524;
															assign node4524 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node4529 = (inp[4]) ? node4541 : node4530;
												assign node4530 = (inp[6]) ? node4532 : 16'b0000000111111111;
													assign node4532 = (inp[13]) ? 16'b0000000011111111 : node4533;
														assign node4533 = (inp[1]) ? node4535 : 16'b0000000111111111;
															assign node4535 = (inp[8]) ? 16'b0000000011111111 : node4536;
																assign node4536 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node4541 = (inp[6]) ? 16'b0000000001111111 : node4542;
													assign node4542 = (inp[8]) ? node4544 : 16'b0000000011111111;
														assign node4544 = (inp[1]) ? node4546 : 16'b0000000011111111;
															assign node4546 = (inp[13]) ? node4548 : 16'b0000000001111111;
																assign node4548 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
								assign node4552 = (inp[13]) ? node4644 : node4553;
									assign node4553 = (inp[0]) ? node4599 : node4554;
										assign node4554 = (inp[8]) ? node4584 : node4555;
											assign node4555 = (inp[6]) ? node4571 : node4556;
												assign node4556 = (inp[14]) ? node4566 : node4557;
													assign node4557 = (inp[12]) ? 16'b0000001111111111 : node4558;
														assign node4558 = (inp[15]) ? 16'b0000011111111111 : node4559;
															assign node4559 = (inp[4]) ? node4561 : 16'b0000111111111111;
																assign node4561 = (inp[1]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node4566 = (inp[4]) ? 16'b0000001111111111 : node4567;
														assign node4567 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node4571 = (inp[12]) ? node4579 : node4572;
													assign node4572 = (inp[4]) ? 16'b0000000111111111 : node4573;
														assign node4573 = (inp[15]) ? 16'b0000001111111111 : node4574;
															assign node4574 = (inp[1]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node4579 = (inp[14]) ? node4581 : 16'b0000000111111111;
														assign node4581 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node4584 = (inp[4]) ? node4592 : node4585;
												assign node4585 = (inp[1]) ? node4587 : 16'b0000001111111111;
													assign node4587 = (inp[15]) ? 16'b0000000011111111 : node4588;
														assign node4588 = (inp[6]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node4592 = (inp[6]) ? node4594 : 16'b0000000111111111;
													assign node4594 = (inp[12]) ? node4596 : 16'b0000000111111111;
														assign node4596 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node4599 = (inp[8]) ? node4625 : node4600;
											assign node4600 = (inp[4]) ? node4612 : node4601;
												assign node4601 = (inp[6]) ? node4603 : 16'b0000001111111111;
													assign node4603 = (inp[12]) ? 16'b0000000001111111 : node4604;
														assign node4604 = (inp[15]) ? 16'b0000000111111111 : node4605;
															assign node4605 = (inp[1]) ? 16'b0000000111111111 : node4606;
																assign node4606 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node4612 = (inp[15]) ? node4622 : node4613;
													assign node4613 = (inp[14]) ? node4617 : node4614;
														assign node4614 = (inp[6]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node4617 = (inp[12]) ? 16'b0000000011111111 : node4618;
															assign node4618 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node4622 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node4625 = (inp[14]) ? node4633 : node4626;
												assign node4626 = (inp[12]) ? node4628 : 16'b0000001111111111;
													assign node4628 = (inp[6]) ? node4630 : 16'b0000000011111111;
														assign node4630 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000001111111;
												assign node4633 = (inp[15]) ? node4637 : node4634;
													assign node4634 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node4637 = (inp[4]) ? node4639 : 16'b0000000001111111;
														assign node4639 = (inp[6]) ? node4641 : 16'b0000000001111111;
															assign node4641 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node4644 = (inp[4]) ? node4692 : node4645;
										assign node4645 = (inp[6]) ? node4677 : node4646;
											assign node4646 = (inp[14]) ? node4664 : node4647;
												assign node4647 = (inp[1]) ? node4649 : 16'b0000011111111111;
													assign node4649 = (inp[8]) ? 16'b0000000011111111 : node4650;
														assign node4650 = (inp[15]) ? node4656 : node4651;
															assign node4651 = (inp[12]) ? node4653 : 16'b0000001111111111;
																assign node4653 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
															assign node4656 = (inp[0]) ? node4660 : node4657;
																assign node4657 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
																assign node4660 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node4664 = (inp[0]) ? node4670 : node4665;
													assign node4665 = (inp[8]) ? node4667 : 16'b0000000111111111;
														assign node4667 = (inp[12]) ? 16'b0000000111111111 : 16'b0000000011111111;
													assign node4670 = (inp[1]) ? node4672 : 16'b0000000011111111;
														assign node4672 = (inp[15]) ? 16'b0000000011111111 : node4673;
															assign node4673 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node4677 = (inp[1]) ? node4685 : node4678;
												assign node4678 = (inp[12]) ? node4680 : 16'b0000000111111111;
													assign node4680 = (inp[0]) ? 16'b0000000011111111 : node4681;
														assign node4681 = (inp[15]) ? 16'b0000000111111111 : 16'b0000000011111111;
												assign node4685 = (inp[12]) ? node4687 : 16'b0000000011111111;
													assign node4687 = (inp[15]) ? 16'b0000000000111111 : node4688;
														assign node4688 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000111111111;
										assign node4692 = (inp[14]) ? node4714 : node4693;
											assign node4693 = (inp[15]) ? node4699 : node4694;
												assign node4694 = (inp[12]) ? 16'b0000000011111111 : node4695;
													assign node4695 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node4699 = (inp[0]) ? node4709 : node4700;
													assign node4700 = (inp[1]) ? node4706 : node4701;
														assign node4701 = (inp[12]) ? node4703 : 16'b0000001111111111;
															assign node4703 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node4706 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node4709 = (inp[8]) ? node4711 : 16'b0000000001111111;
														assign node4711 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node4714 = (inp[15]) ? node4724 : node4715;
												assign node4715 = (inp[1]) ? node4717 : 16'b0000000011111111;
													assign node4717 = (inp[0]) ? node4721 : node4718;
														assign node4718 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node4721 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node4724 = (inp[6]) ? node4728 : node4725;
													assign node4725 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node4728 = (inp[0]) ? 16'b0000000000111111 : node4729;
														assign node4729 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
							assign node4733 = (inp[14]) ? node4949 : node4734;
								assign node4734 = (inp[0]) ? node4844 : node4735;
									assign node4735 = (inp[13]) ? node4789 : node4736;
										assign node4736 = (inp[9]) ? node4748 : node4737;
											assign node4737 = (inp[1]) ? node4741 : node4738;
												assign node4738 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node4741 = (inp[12]) ? node4743 : 16'b0000001111111111;
													assign node4743 = (inp[4]) ? 16'b0000000111111111 : node4744;
														assign node4744 = (inp[6]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node4748 = (inp[15]) ? node4766 : node4749;
												assign node4749 = (inp[6]) ? node4757 : node4750;
													assign node4750 = (inp[4]) ? node4754 : node4751;
														assign node4751 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node4754 = (inp[1]) ? 16'b0000001111111111 : 16'b0000000111111111;
													assign node4757 = (inp[1]) ? node4763 : node4758;
														assign node4758 = (inp[12]) ? node4760 : 16'b0000001111111111;
															assign node4760 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node4763 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node4766 = (inp[4]) ? node4778 : node4767;
													assign node4767 = (inp[8]) ? node4775 : node4768;
														assign node4768 = (inp[6]) ? node4770 : 16'b0000001111111111;
															assign node4770 = (inp[1]) ? 16'b0000000111111111 : node4771;
																assign node4771 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node4775 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node4778 = (inp[8]) ? node4786 : node4779;
														assign node4779 = (inp[12]) ? 16'b0000000011111111 : node4780;
															assign node4780 = (inp[6]) ? node4782 : 16'b0000000111111111;
																assign node4782 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node4786 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node4789 = (inp[12]) ? node4823 : node4790;
											assign node4790 = (inp[15]) ? node4800 : node4791;
												assign node4791 = (inp[8]) ? 16'b0000001111111111 : node4792;
													assign node4792 = (inp[9]) ? 16'b0000000111111111 : node4793;
														assign node4793 = (inp[6]) ? node4795 : 16'b0000001111111111;
															assign node4795 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node4800 = (inp[6]) ? node4814 : node4801;
													assign node4801 = (inp[4]) ? node4809 : node4802;
														assign node4802 = (inp[8]) ? node4804 : 16'b0000001111111111;
															assign node4804 = (inp[9]) ? 16'b0000000111111111 : node4805;
																assign node4805 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node4809 = (inp[9]) ? node4811 : 16'b0000000111111111;
															assign node4811 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node4814 = (inp[1]) ? node4820 : node4815;
														assign node4815 = (inp[8]) ? 16'b0000000011111111 : node4816;
															assign node4816 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node4820 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node4823 = (inp[8]) ? node4837 : node4824;
												assign node4824 = (inp[4]) ? node4832 : node4825;
													assign node4825 = (inp[9]) ? node4827 : 16'b0000000111111111;
														assign node4827 = (inp[6]) ? 16'b0000000011111111 : node4828;
															assign node4828 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node4832 = (inp[1]) ? 16'b0000000011111111 : node4833;
														assign node4833 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node4837 = (inp[9]) ? 16'b0000000001111111 : node4838;
													assign node4838 = (inp[6]) ? 16'b0000000001111111 : node4839;
														assign node4839 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node4844 = (inp[15]) ? node4900 : node4845;
										assign node4845 = (inp[13]) ? node4873 : node4846;
											assign node4846 = (inp[9]) ? node4856 : node4847;
												assign node4847 = (inp[4]) ? node4851 : node4848;
													assign node4848 = (inp[6]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node4851 = (inp[6]) ? 16'b0000000011111111 : node4852;
														assign node4852 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node4856 = (inp[4]) ? node4868 : node4857;
													assign node4857 = (inp[1]) ? node4865 : node4858;
														assign node4858 = (inp[12]) ? node4860 : 16'b0000001111111111;
															assign node4860 = (inp[8]) ? 16'b0000000111111111 : node4861;
																assign node4861 = (inp[6]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node4865 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node4868 = (inp[12]) ? 16'b0000000011111111 : node4869;
														assign node4869 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node4873 = (inp[8]) ? node4885 : node4874;
												assign node4874 = (inp[9]) ? node4880 : node4875;
													assign node4875 = (inp[4]) ? 16'b0000000111111111 : node4876;
														assign node4876 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node4880 = (inp[12]) ? 16'b0000000011111111 : node4881;
														assign node4881 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node4885 = (inp[1]) ? node4895 : node4886;
													assign node4886 = (inp[12]) ? node4890 : node4887;
														assign node4887 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node4890 = (inp[9]) ? node4892 : 16'b0000000011111111;
															assign node4892 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node4895 = (inp[6]) ? node4897 : 16'b0000000001111111;
														assign node4897 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node4900 = (inp[12]) ? node4922 : node4901;
											assign node4901 = (inp[9]) ? node4913 : node4902;
												assign node4902 = (inp[6]) ? node4908 : node4903;
													assign node4903 = (inp[13]) ? node4905 : 16'b0000000111111111;
														assign node4905 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node4908 = (inp[8]) ? node4910 : 16'b0000000011111111;
														assign node4910 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node4913 = (inp[6]) ? node4917 : node4914;
													assign node4914 = (inp[8]) ? 16'b0000000111111111 : 16'b0000000011111111;
													assign node4917 = (inp[1]) ? 16'b0000000001111111 : node4918;
														assign node4918 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node4922 = (inp[4]) ? node4936 : node4923;
												assign node4923 = (inp[1]) ? node4927 : node4924;
													assign node4924 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node4927 = (inp[9]) ? node4931 : node4928;
														assign node4928 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node4931 = (inp[6]) ? node4933 : 16'b0000000001111111;
															assign node4933 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node4936 = (inp[9]) ? node4944 : node4937;
													assign node4937 = (inp[6]) ? node4939 : 16'b0000000001111111;
														assign node4939 = (inp[13]) ? 16'b0000000000111111 : node4940;
															assign node4940 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node4944 = (inp[6]) ? node4946 : 16'b0000000000111111;
														assign node4946 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
								assign node4949 = (inp[8]) ? node5041 : node4950;
									assign node4950 = (inp[6]) ? node5000 : node4951;
										assign node4951 = (inp[4]) ? node4983 : node4952;
											assign node4952 = (inp[12]) ? node4966 : node4953;
												assign node4953 = (inp[1]) ? 16'b0000000111111111 : node4954;
													assign node4954 = (inp[9]) ? node4958 : node4955;
														assign node4955 = (inp[0]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node4958 = (inp[13]) ? 16'b0000000111111111 : node4959;
															assign node4959 = (inp[0]) ? node4961 : 16'b0000001111111111;
																assign node4961 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node4966 = (inp[15]) ? node4978 : node4967;
													assign node4967 = (inp[1]) ? node4973 : node4968;
														assign node4968 = (inp[9]) ? 16'b0000000111111111 : node4969;
															assign node4969 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node4973 = (inp[0]) ? node4975 : 16'b0000000111111111;
															assign node4975 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node4978 = (inp[0]) ? 16'b0000000000111111 : node4979;
														assign node4979 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node4983 = (inp[15]) ? node4991 : node4984;
												assign node4984 = (inp[13]) ? 16'b0000000011111111 : node4985;
													assign node4985 = (inp[9]) ? 16'b0000000111111111 : node4986;
														assign node4986 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node4991 = (inp[0]) ? node4995 : node4992;
													assign node4992 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node4995 = (inp[13]) ? 16'b0000000001111111 : node4996;
														assign node4996 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node5000 = (inp[1]) ? node5016 : node5001;
											assign node5001 = (inp[12]) ? node5013 : node5002;
												assign node5002 = (inp[13]) ? node5008 : node5003;
													assign node5003 = (inp[0]) ? 16'b0000000111111111 : node5004;
														assign node5004 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node5008 = (inp[0]) ? 16'b0000000001111111 : node5009;
														assign node5009 = (inp[15]) ? 16'b0000000011111111 : 16'b0000001111111111;
												assign node5013 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node5016 = (inp[0]) ? node5026 : node5017;
												assign node5017 = (inp[15]) ? node5021 : node5018;
													assign node5018 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node5021 = (inp[9]) ? node5023 : 16'b0000000011111111;
														assign node5023 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node5026 = (inp[12]) ? node5032 : node5027;
													assign node5027 = (inp[15]) ? node5029 : 16'b0000000001111111;
														assign node5029 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node5032 = (inp[13]) ? node5038 : node5033;
														assign node5033 = (inp[9]) ? node5035 : 16'b0000000001111111;
															assign node5035 = (inp[4]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node5038 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node5041 = (inp[6]) ? node5093 : node5042;
										assign node5042 = (inp[12]) ? node5058 : node5043;
											assign node5043 = (inp[0]) ? node5049 : node5044;
												assign node5044 = (inp[13]) ? node5046 : 16'b0000000111111111;
													assign node5046 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node5049 = (inp[15]) ? node5051 : 16'b0000000011111111;
													assign node5051 = (inp[13]) ? node5055 : node5052;
														assign node5052 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node5055 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node5058 = (inp[15]) ? node5078 : node5059;
												assign node5059 = (inp[13]) ? node5065 : node5060;
													assign node5060 = (inp[4]) ? node5062 : 16'b0000000111111111;
														assign node5062 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node5065 = (inp[9]) ? node5071 : node5066;
														assign node5066 = (inp[1]) ? 16'b0000000001111111 : node5067;
															assign node5067 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node5071 = (inp[1]) ? 16'b0000000000111111 : node5072;
															assign node5072 = (inp[4]) ? node5074 : 16'b0000000001111111;
																assign node5074 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node5078 = (inp[0]) ? node5088 : node5079;
													assign node5079 = (inp[9]) ? node5081 : 16'b0000000001111111;
														assign node5081 = (inp[13]) ? node5083 : 16'b0000000001111111;
															assign node5083 = (inp[4]) ? 16'b0000000000111111 : node5084;
																assign node5084 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node5088 = (inp[9]) ? 16'b0000000000111111 : node5089;
														assign node5089 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node5093 = (inp[15]) ? node5125 : node5094;
											assign node5094 = (inp[9]) ? node5114 : node5095;
												assign node5095 = (inp[1]) ? node5103 : node5096;
													assign node5096 = (inp[13]) ? node5100 : node5097;
														assign node5097 = (inp[0]) ? 16'b0000000011111111 : 16'b0000001111111111;
														assign node5100 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node5103 = (inp[13]) ? node5109 : node5104;
														assign node5104 = (inp[4]) ? 16'b0000000001111111 : node5105;
															assign node5105 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node5109 = (inp[0]) ? node5111 : 16'b0000000001111111;
															assign node5111 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node5114 = (inp[0]) ? node5120 : node5115;
													assign node5115 = (inp[1]) ? node5117 : 16'b0000000001111111;
														assign node5117 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node5120 = (inp[13]) ? 16'b0000000000111111 : node5121;
														assign node5121 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node5125 = (inp[0]) ? node5149 : node5126;
												assign node5126 = (inp[1]) ? node5140 : node5127;
													assign node5127 = (inp[12]) ? node5135 : node5128;
														assign node5128 = (inp[13]) ? 16'b0000000001111111 : node5129;
															assign node5129 = (inp[9]) ? 16'b0000000011111111 : node5130;
																assign node5130 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node5135 = (inp[4]) ? node5137 : 16'b0000000001111111;
															assign node5137 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node5140 = (inp[13]) ? node5144 : node5141;
														assign node5141 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000000111111;
														assign node5144 = (inp[4]) ? node5146 : 16'b0000000000111111;
															assign node5146 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node5149 = (inp[4]) ? 16'b0000000000011111 : node5150;
													assign node5150 = (inp[9]) ? node5152 : 16'b0000000000111111;
														assign node5152 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000111111;
						assign node5156 = (inp[6]) ? node5508 : node5157;
							assign node5157 = (inp[9]) ? node5317 : node5158;
								assign node5158 = (inp[0]) ? node5244 : node5159;
									assign node5159 = (inp[13]) ? node5197 : node5160;
										assign node5160 = (inp[12]) ? node5178 : node5161;
											assign node5161 = (inp[8]) ? node5167 : node5162;
												assign node5162 = (inp[15]) ? node5164 : 16'b0000011111111111;
													assign node5164 = (inp[1]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node5167 = (inp[5]) ? node5171 : node5168;
													assign node5168 = (inp[15]) ? 16'b0000001111111111 : 16'b0000111111111111;
													assign node5171 = (inp[15]) ? 16'b0000000011111111 : node5172;
														assign node5172 = (inp[14]) ? 16'b0000000111111111 : node5173;
															assign node5173 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node5178 = (inp[5]) ? node5184 : node5179;
												assign node5179 = (inp[15]) ? node5181 : 16'b0000001111111111;
													assign node5181 = (inp[14]) ? 16'b0000001111111111 : 16'b0000000111111111;
												assign node5184 = (inp[4]) ? node5190 : node5185;
													assign node5185 = (inp[8]) ? 16'b0000000111111111 : node5186;
														assign node5186 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node5190 = (inp[14]) ? node5194 : node5191;
														assign node5191 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node5194 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node5197 = (inp[1]) ? node5227 : node5198;
											assign node5198 = (inp[4]) ? node5216 : node5199;
												assign node5199 = (inp[8]) ? node5209 : node5200;
													assign node5200 = (inp[5]) ? node5202 : 16'b0000001111111111;
														assign node5202 = (inp[12]) ? 16'b0000000111111111 : node5203;
															assign node5203 = (inp[15]) ? node5205 : 16'b0000001111111111;
																assign node5205 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node5209 = (inp[14]) ? 16'b0000000011111111 : node5210;
														assign node5210 = (inp[5]) ? 16'b0000000111111111 : node5211;
															assign node5211 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node5216 = (inp[15]) ? node5218 : 16'b0000000111111111;
													assign node5218 = (inp[8]) ? 16'b0000000001111111 : node5219;
														assign node5219 = (inp[5]) ? node5221 : 16'b0000000111111111;
															assign node5221 = (inp[14]) ? 16'b0000000011111111 : node5222;
																assign node5222 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node5227 = (inp[12]) ? node5235 : node5228;
												assign node5228 = (inp[15]) ? node5230 : 16'b0000001111111111;
													assign node5230 = (inp[14]) ? 16'b0000000011111111 : node5231;
														assign node5231 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node5235 = (inp[8]) ? 16'b0000000001111111 : node5236;
													assign node5236 = (inp[5]) ? 16'b0000000011111111 : node5237;
														assign node5237 = (inp[14]) ? node5239 : 16'b0000000111111111;
															assign node5239 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node5244 = (inp[4]) ? node5280 : node5245;
										assign node5245 = (inp[1]) ? node5263 : node5246;
											assign node5246 = (inp[8]) ? node5254 : node5247;
												assign node5247 = (inp[12]) ? node5251 : node5248;
													assign node5248 = (inp[15]) ? 16'b0000001111111111 : 16'b0000111111111111;
													assign node5251 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node5254 = (inp[13]) ? node5256 : 16'b0000000111111111;
													assign node5256 = (inp[15]) ? 16'b0000000011111111 : node5257;
														assign node5257 = (inp[5]) ? node5259 : 16'b0000000111111111;
															assign node5259 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node5263 = (inp[13]) ? node5275 : node5264;
												assign node5264 = (inp[12]) ? node5266 : 16'b0000000111111111;
													assign node5266 = (inp[8]) ? node5272 : node5267;
														assign node5267 = (inp[14]) ? node5269 : 16'b0000000111111111;
															assign node5269 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node5272 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node5275 = (inp[5]) ? node5277 : 16'b0000000111111111;
													assign node5277 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node5280 = (inp[15]) ? node5306 : node5281;
											assign node5281 = (inp[12]) ? node5295 : node5282;
												assign node5282 = (inp[8]) ? node5288 : node5283;
													assign node5283 = (inp[1]) ? 16'b0000000111111111 : node5284;
														assign node5284 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node5288 = (inp[1]) ? 16'b0000000011111111 : node5289;
														assign node5289 = (inp[5]) ? 16'b0000000011111111 : node5290;
															assign node5290 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node5295 = (inp[13]) ? node5301 : node5296;
													assign node5296 = (inp[8]) ? 16'b0000000001111111 : node5297;
														assign node5297 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node5301 = (inp[8]) ? node5303 : 16'b0000000001111111;
														assign node5303 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node5306 = (inp[1]) ? node5310 : node5307;
												assign node5307 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node5310 = (inp[5]) ? 16'b0000000000111111 : node5311;
													assign node5311 = (inp[12]) ? node5313 : 16'b0000000001111111;
														assign node5313 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
								assign node5317 = (inp[15]) ? node5425 : node5318;
									assign node5318 = (inp[4]) ? node5376 : node5319;
										assign node5319 = (inp[13]) ? node5353 : node5320;
											assign node5320 = (inp[0]) ? node5340 : node5321;
												assign node5321 = (inp[5]) ? node5331 : node5322;
													assign node5322 = (inp[14]) ? 16'b0000001111111111 : node5323;
														assign node5323 = (inp[8]) ? 16'b0000001111111111 : node5324;
															assign node5324 = (inp[1]) ? node5326 : 16'b0000011111111111;
																assign node5326 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node5331 = (inp[14]) ? node5337 : node5332;
														assign node5332 = (inp[1]) ? node5334 : 16'b0000001111111111;
															assign node5334 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node5337 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node5340 = (inp[8]) ? node5348 : node5341;
													assign node5341 = (inp[14]) ? node5343 : 16'b0000000111111111;
														assign node5343 = (inp[5]) ? 16'b0000000111111111 : node5344;
															assign node5344 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node5348 = (inp[14]) ? node5350 : 16'b0000000111111111;
														assign node5350 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node5353 = (inp[14]) ? node5363 : node5354;
												assign node5354 = (inp[1]) ? node5358 : node5355;
													assign node5355 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node5358 = (inp[5]) ? 16'b0000000011111111 : node5359;
														assign node5359 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node5363 = (inp[1]) ? node5369 : node5364;
													assign node5364 = (inp[8]) ? node5366 : 16'b0000000011111111;
														assign node5366 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node5369 = (inp[5]) ? node5373 : node5370;
														assign node5370 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node5373 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node5376 = (inp[5]) ? node5398 : node5377;
											assign node5377 = (inp[0]) ? node5385 : node5378;
												assign node5378 = (inp[13]) ? 16'b0000000011111111 : node5379;
													assign node5379 = (inp[14]) ? 16'b0000000111111111 : node5380;
														assign node5380 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node5385 = (inp[1]) ? node5391 : node5386;
													assign node5386 = (inp[13]) ? 16'b0000000011111111 : node5387;
														assign node5387 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node5391 = (inp[13]) ? 16'b0000000000111111 : node5392;
														assign node5392 = (inp[14]) ? 16'b0000000001111111 : node5393;
															assign node5393 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node5398 = (inp[14]) ? node5404 : node5399;
												assign node5399 = (inp[12]) ? 16'b0000000001111111 : node5400;
													assign node5400 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000111111111;
												assign node5404 = (inp[8]) ? node5416 : node5405;
													assign node5405 = (inp[1]) ? node5411 : node5406;
														assign node5406 = (inp[0]) ? 16'b0000000001111111 : node5407;
															assign node5407 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node5411 = (inp[0]) ? 16'b0000000000111111 : node5412;
															assign node5412 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node5416 = (inp[12]) ? node5418 : 16'b0000000000111111;
														assign node5418 = (inp[0]) ? node5420 : 16'b0000000000011111;
															assign node5420 = (inp[13]) ? node5422 : 16'b0000000000011111;
																assign node5422 = (inp[1]) ? 16'b0000000000001111 : 16'b0000000000011111;
									assign node5425 = (inp[12]) ? node5469 : node5426;
										assign node5426 = (inp[8]) ? node5456 : node5427;
											assign node5427 = (inp[4]) ? node5431 : node5428;
												assign node5428 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node5431 = (inp[5]) ? node5443 : node5432;
													assign node5432 = (inp[0]) ? node5440 : node5433;
														assign node5433 = (inp[14]) ? 16'b0000000011111111 : node5434;
															assign node5434 = (inp[1]) ? node5436 : 16'b0000000111111111;
																assign node5436 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node5440 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node5443 = (inp[1]) ? node5449 : node5444;
														assign node5444 = (inp[0]) ? 16'b0000000001111111 : node5445;
															assign node5445 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node5449 = (inp[14]) ? 16'b0000000000111111 : node5450;
															assign node5450 = (inp[0]) ? node5452 : 16'b0000000001111111;
																assign node5452 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node5456 = (inp[0]) ? node5462 : node5457;
												assign node5457 = (inp[14]) ? 16'b0000000001111111 : node5458;
													assign node5458 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node5462 = (inp[4]) ? node5466 : node5463;
													assign node5463 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node5466 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node5469 = (inp[1]) ? node5491 : node5470;
											assign node5470 = (inp[0]) ? node5480 : node5471;
												assign node5471 = (inp[13]) ? 16'b0000000001111111 : node5472;
													assign node5472 = (inp[14]) ? node5474 : 16'b0000000001111111;
														assign node5474 = (inp[8]) ? node5476 : 16'b0000000001111111;
															assign node5476 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node5480 = (inp[4]) ? node5488 : node5481;
													assign node5481 = (inp[13]) ? 16'b0000000000111111 : node5482;
														assign node5482 = (inp[8]) ? node5484 : 16'b0000000011111111;
															assign node5484 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node5488 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node5491 = (inp[8]) ? 16'b0000000000011111 : node5492;
												assign node5492 = (inp[0]) ? node5500 : node5493;
													assign node5493 = (inp[5]) ? node5495 : 16'b0000000011111111;
														assign node5495 = (inp[4]) ? 16'b0000000000111111 : node5496;
															assign node5496 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node5500 = (inp[14]) ? 16'b0000000000111111 : node5501;
														assign node5501 = (inp[13]) ? node5503 : 16'b0000000000111111;
															assign node5503 = (inp[4]) ? 16'b0000000000011111 : 16'b0000000000111111;
							assign node5508 = (inp[8]) ? node5690 : node5509;
								assign node5509 = (inp[1]) ? node5599 : node5510;
									assign node5510 = (inp[13]) ? node5566 : node5511;
										assign node5511 = (inp[4]) ? node5537 : node5512;
											assign node5512 = (inp[14]) ? node5526 : node5513;
												assign node5513 = (inp[9]) ? node5521 : node5514;
													assign node5514 = (inp[5]) ? node5516 : 16'b0000001111111111;
														assign node5516 = (inp[0]) ? node5518 : 16'b0000001111111111;
															assign node5518 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node5521 = (inp[15]) ? 16'b0000000111111111 : node5522;
														assign node5522 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node5526 = (inp[12]) ? 16'b0000000011111111 : node5527;
													assign node5527 = (inp[5]) ? node5529 : 16'b0000001111111111;
														assign node5529 = (inp[0]) ? 16'b0000000011111111 : node5530;
															assign node5530 = (inp[9]) ? node5532 : 16'b0000000111111111;
																assign node5532 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node5537 = (inp[5]) ? node5555 : node5538;
												assign node5538 = (inp[15]) ? node5550 : node5539;
													assign node5539 = (inp[12]) ? node5545 : node5540;
														assign node5540 = (inp[0]) ? 16'b0000000111111111 : node5541;
															assign node5541 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node5545 = (inp[9]) ? node5547 : 16'b0000000111111111;
															assign node5547 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node5550 = (inp[12]) ? node5552 : 16'b0000000011111111;
														assign node5552 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000011111111;
												assign node5555 = (inp[12]) ? node5559 : node5556;
													assign node5556 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node5559 = (inp[0]) ? node5561 : 16'b0000000001111111;
														assign node5561 = (inp[9]) ? node5563 : 16'b0000000000111111;
															assign node5563 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node5566 = (inp[14]) ? node5578 : node5567;
											assign node5567 = (inp[5]) ? node5573 : node5568;
												assign node5568 = (inp[12]) ? 16'b0000000011111111 : node5569;
													assign node5569 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node5573 = (inp[9]) ? 16'b0000000001111111 : node5574;
													assign node5574 = (inp[4]) ? 16'b0000000111111111 : 16'b0000000011111111;
											assign node5578 = (inp[15]) ? node5590 : node5579;
												assign node5579 = (inp[0]) ? node5587 : node5580;
													assign node5580 = (inp[5]) ? node5584 : node5581;
														assign node5581 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node5584 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000001111111;
													assign node5587 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node5590 = (inp[9]) ? node5592 : 16'b0000000000011111;
													assign node5592 = (inp[0]) ? 16'b0000000000111111 : node5593;
														assign node5593 = (inp[4]) ? node5595 : 16'b0000000001111111;
															assign node5595 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node5599 = (inp[9]) ? node5649 : node5600;
										assign node5600 = (inp[15]) ? node5626 : node5601;
											assign node5601 = (inp[0]) ? node5619 : node5602;
												assign node5602 = (inp[5]) ? node5610 : node5603;
													assign node5603 = (inp[4]) ? node5607 : node5604;
														assign node5604 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node5607 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node5610 = (inp[4]) ? 16'b0000000011111111 : node5611;
														assign node5611 = (inp[14]) ? node5613 : 16'b0000000111111111;
															assign node5613 = (inp[12]) ? 16'b0000000011111111 : node5614;
																assign node5614 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node5619 = (inp[4]) ? node5621 : 16'b0000000011111111;
													assign node5621 = (inp[13]) ? 16'b0000000001111111 : node5622;
														assign node5622 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node5626 = (inp[5]) ? node5642 : node5627;
												assign node5627 = (inp[4]) ? node5635 : node5628;
													assign node5628 = (inp[13]) ? node5632 : node5629;
														assign node5629 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node5632 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000011111111;
													assign node5635 = (inp[0]) ? node5639 : node5636;
														assign node5636 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node5639 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000001111111;
												assign node5642 = (inp[4]) ? 16'b0000000000111111 : node5643;
													assign node5643 = (inp[13]) ? node5645 : 16'b0000000011111111;
														assign node5645 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node5649 = (inp[5]) ? node5675 : node5650;
											assign node5650 = (inp[15]) ? node5664 : node5651;
												assign node5651 = (inp[13]) ? 16'b0000000001111111 : node5652;
													assign node5652 = (inp[0]) ? node5654 : 16'b0000000111111111;
														assign node5654 = (inp[12]) ? node5660 : node5655;
															assign node5655 = (inp[4]) ? node5657 : 16'b0000000011111111;
																assign node5657 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
															assign node5660 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node5664 = (inp[14]) ? node5666 : 16'b0000000001111111;
													assign node5666 = (inp[0]) ? 16'b0000000000001111 : node5667;
														assign node5667 = (inp[12]) ? node5669 : 16'b0000000001111111;
															assign node5669 = (inp[4]) ? node5671 : 16'b0000000000111111;
																assign node5671 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node5675 = (inp[4]) ? node5679 : node5676;
												assign node5676 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node5679 = (inp[12]) ? node5685 : node5680;
													assign node5680 = (inp[14]) ? node5682 : 16'b0000000000111111;
														assign node5682 = (inp[0]) ? 16'b0000000000001111 : 16'b0000000000111111;
													assign node5685 = (inp[15]) ? node5687 : 16'b0000000000011111;
														assign node5687 = (inp[0]) ? 16'b0000000000001111 : 16'b0000000000011111;
								assign node5690 = (inp[14]) ? node5776 : node5691;
									assign node5691 = (inp[4]) ? node5733 : node5692;
										assign node5692 = (inp[0]) ? node5714 : node5693;
											assign node5693 = (inp[12]) ? node5697 : node5694;
												assign node5694 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node5697 = (inp[1]) ? node5707 : node5698;
													assign node5698 = (inp[9]) ? node5700 : 16'b0000000011111111;
														assign node5700 = (inp[13]) ? node5702 : 16'b0000000011111111;
															assign node5702 = (inp[5]) ? 16'b0000000001111111 : node5703;
																assign node5703 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node5707 = (inp[5]) ? 16'b0000000001111111 : node5708;
														assign node5708 = (inp[9]) ? 16'b0000000001111111 : node5709;
															assign node5709 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node5714 = (inp[13]) ? node5730 : node5715;
												assign node5715 = (inp[12]) ? node5721 : node5716;
													assign node5716 = (inp[15]) ? node5718 : 16'b0000000011111111;
														assign node5718 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node5721 = (inp[5]) ? node5727 : node5722;
														assign node5722 = (inp[15]) ? 16'b0000000001111111 : node5723;
															assign node5723 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node5727 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node5730 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000000111111;
										assign node5733 = (inp[9]) ? node5749 : node5734;
											assign node5734 = (inp[5]) ? node5746 : node5735;
												assign node5735 = (inp[0]) ? node5739 : node5736;
													assign node5736 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node5739 = (inp[1]) ? node5743 : node5740;
														assign node5740 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node5743 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node5746 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node5749 = (inp[5]) ? node5767 : node5750;
												assign node5750 = (inp[12]) ? node5758 : node5751;
													assign node5751 = (inp[13]) ? 16'b0000000011111111 : node5752;
														assign node5752 = (inp[0]) ? node5754 : 16'b0000000001111111;
															assign node5754 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node5758 = (inp[0]) ? node5764 : node5759;
														assign node5759 = (inp[1]) ? 16'b0000000000111111 : node5760;
															assign node5760 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node5764 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000000011111;
												assign node5767 = (inp[12]) ? node5773 : node5768;
													assign node5768 = (inp[1]) ? node5770 : 16'b0000000001111111;
														assign node5770 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node5773 = (inp[13]) ? 16'b0000000000001111 : 16'b0000000000011111;
									assign node5776 = (inp[13]) ? node5818 : node5777;
										assign node5777 = (inp[0]) ? node5793 : node5778;
											assign node5778 = (inp[9]) ? node5788 : node5779;
												assign node5779 = (inp[1]) ? node5785 : node5780;
													assign node5780 = (inp[4]) ? 16'b0000000011111111 : node5781;
														assign node5781 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node5785 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000111111111;
												assign node5788 = (inp[4]) ? node5790 : 16'b0000000001111111;
													assign node5790 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node5793 = (inp[12]) ? node5807 : node5794;
												assign node5794 = (inp[15]) ? 16'b0000000000011111 : node5795;
													assign node5795 = (inp[9]) ? 16'b0000000000111111 : node5796;
														assign node5796 = (inp[5]) ? node5802 : node5797;
															assign node5797 = (inp[1]) ? node5799 : 16'b0000000011111111;
																assign node5799 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
															assign node5802 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node5807 = (inp[9]) ? node5809 : 16'b0000000000111111;
													assign node5809 = (inp[1]) ? node5815 : node5810;
														assign node5810 = (inp[5]) ? node5812 : 16'b0000000000111111;
															assign node5812 = (inp[4]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node5815 = (inp[4]) ? 16'b0000000000001111 : 16'b0000000000011111;
										assign node5818 = (inp[0]) ? node5846 : node5819;
											assign node5819 = (inp[12]) ? node5835 : node5820;
												assign node5820 = (inp[9]) ? node5824 : node5821;
													assign node5821 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node5824 = (inp[1]) ? node5832 : node5825;
														assign node5825 = (inp[4]) ? node5827 : 16'b0000000001111111;
															assign node5827 = (inp[15]) ? 16'b0000000000111111 : node5828;
																assign node5828 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node5832 = (inp[4]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node5835 = (inp[1]) ? node5841 : node5836;
													assign node5836 = (inp[4]) ? 16'b0000000000011111 : node5837;
														assign node5837 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node5841 = (inp[9]) ? 16'b0000000000000111 : node5842;
														assign node5842 = (inp[4]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node5846 = (inp[9]) ? node5858 : node5847;
												assign node5847 = (inp[4]) ? node5853 : node5848;
													assign node5848 = (inp[15]) ? node5850 : 16'b0000000001111111;
														assign node5850 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node5853 = (inp[1]) ? 16'b0000000000001111 : node5854;
														assign node5854 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node5858 = (inp[1]) ? node5864 : node5859;
													assign node5859 = (inp[4]) ? node5861 : 16'b0000000000011111;
														assign node5861 = (inp[15]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node5864 = (inp[15]) ? node5872 : node5865;
														assign node5865 = (inp[12]) ? 16'b0000000000001111 : node5866;
															assign node5866 = (inp[4]) ? node5868 : 16'b0000000000011111;
																assign node5868 = (inp[5]) ? 16'b0000000000001111 : 16'b0000000000011111;
														assign node5872 = (inp[5]) ? 16'b0000000000000111 : node5873;
															assign node5873 = (inp[4]) ? 16'b0000000000001111 : 16'b0000000000011111;
			assign node5877 = (inp[15]) ? node8951 : node5878;
				assign node5878 = (inp[12]) ? node7412 : node5879;
					assign node5879 = (inp[1]) ? node6607 : node5880;
						assign node5880 = (inp[4]) ? node6254 : node5881;
							assign node5881 = (inp[8]) ? node6075 : node5882;
								assign node5882 = (inp[5]) ? node5994 : node5883;
									assign node5883 = (inp[9]) ? node5939 : node5884;
										assign node5884 = (inp[14]) ? node5914 : node5885;
											assign node5885 = (inp[10]) ? node5897 : node5886;
												assign node5886 = (inp[0]) ? node5890 : node5887;
													assign node5887 = (inp[6]) ? 16'b0001111111111111 : 16'b0011111111111111;
													assign node5890 = (inp[13]) ? node5892 : 16'b0001111111111111;
														assign node5892 = (inp[3]) ? node5894 : 16'b0000111111111111;
															assign node5894 = (inp[2]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node5897 = (inp[6]) ? node5907 : node5898;
													assign node5898 = (inp[0]) ? node5902 : node5899;
														assign node5899 = (inp[13]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node5902 = (inp[3]) ? node5904 : 16'b0000111111111111;
															assign node5904 = (inp[13]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node5907 = (inp[3]) ? 16'b0000011111111111 : node5908;
														assign node5908 = (inp[2]) ? node5910 : 16'b0000111111111111;
															assign node5910 = (inp[13]) ? 16'b0000011111111111 : 16'b0000111111111111;
											assign node5914 = (inp[2]) ? node5928 : node5915;
												assign node5915 = (inp[0]) ? node5921 : node5916;
													assign node5916 = (inp[6]) ? 16'b0000111111111111 : node5917;
														assign node5917 = (inp[3]) ? 16'b0000111111111111 : 16'b0001111111111111;
													assign node5921 = (inp[3]) ? node5923 : 16'b0000111111111111;
														assign node5923 = (inp[13]) ? 16'b0000011111111111 : node5924;
															assign node5924 = (inp[6]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node5928 = (inp[13]) ? node5934 : node5929;
													assign node5929 = (inp[6]) ? 16'b0000011111111111 : node5930;
														assign node5930 = (inp[0]) ? 16'b0000111111111111 : 16'b0000011111111111;
													assign node5934 = (inp[0]) ? 16'b0000000011111111 : node5935;
														assign node5935 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
										assign node5939 = (inp[13]) ? node5963 : node5940;
											assign node5940 = (inp[10]) ? node5950 : node5941;
												assign node5941 = (inp[6]) ? 16'b0000011111111111 : node5942;
													assign node5942 = (inp[3]) ? 16'b0000111111111111 : node5943;
														assign node5943 = (inp[0]) ? 16'b0000111111111111 : node5944;
															assign node5944 = (inp[14]) ? 16'b0001111111111111 : 16'b0011111111111111;
												assign node5950 = (inp[0]) ? node5954 : node5951;
													assign node5951 = (inp[6]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node5954 = (inp[14]) ? 16'b0000001111111111 : node5955;
														assign node5955 = (inp[3]) ? node5957 : 16'b0000011111111111;
															assign node5957 = (inp[6]) ? 16'b0000001111111111 : node5958;
																assign node5958 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node5963 = (inp[0]) ? node5977 : node5964;
												assign node5964 = (inp[10]) ? node5972 : node5965;
													assign node5965 = (inp[14]) ? node5967 : 16'b0000011111111111;
														assign node5967 = (inp[6]) ? 16'b0000011111111111 : node5968;
															assign node5968 = (inp[3]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node5972 = (inp[3]) ? node5974 : 16'b0000011111111111;
														assign node5974 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node5977 = (inp[10]) ? node5985 : node5978;
													assign node5978 = (inp[3]) ? node5982 : node5979;
														assign node5979 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node5982 = (inp[6]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node5985 = (inp[6]) ? node5989 : node5986;
														assign node5986 = (inp[3]) ? 16'b0000000111111111 : 16'b0000011111111111;
														assign node5989 = (inp[14]) ? node5991 : 16'b0000000111111111;
															assign node5991 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node5994 = (inp[3]) ? node6042 : node5995;
										assign node5995 = (inp[6]) ? node6015 : node5996;
											assign node5996 = (inp[2]) ? node6010 : node5997;
												assign node5997 = (inp[10]) ? node6005 : node5998;
													assign node5998 = (inp[13]) ? node6002 : node5999;
														assign node5999 = (inp[14]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node6002 = (inp[14]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node6005 = (inp[14]) ? node6007 : 16'b0000011111111111;
														assign node6007 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node6010 = (inp[13]) ? node6012 : 16'b0000011111111111;
													assign node6012 = (inp[0]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node6015 = (inp[2]) ? node6027 : node6016;
												assign node6016 = (inp[9]) ? node6022 : node6017;
													assign node6017 = (inp[0]) ? node6019 : 16'b0000011111111111;
														assign node6019 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node6022 = (inp[13]) ? 16'b0000001111111111 : node6023;
														assign node6023 = (inp[14]) ? 16'b0000001111111111 : 16'b0000111111111111;
												assign node6027 = (inp[10]) ? node6035 : node6028;
													assign node6028 = (inp[14]) ? node6032 : node6029;
														assign node6029 = (inp[9]) ? 16'b0000001111111111 : 16'b0000111111111111;
														assign node6032 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node6035 = (inp[0]) ? node6039 : node6036;
														assign node6036 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node6039 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node6042 = (inp[9]) ? node6064 : node6043;
											assign node6043 = (inp[0]) ? node6053 : node6044;
												assign node6044 = (inp[14]) ? 16'b0000001111111111 : node6045;
													assign node6045 = (inp[2]) ? 16'b0000001111111111 : node6046;
														assign node6046 = (inp[10]) ? 16'b0000011111111111 : node6047;
															assign node6047 = (inp[6]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node6053 = (inp[14]) ? node6061 : node6054;
													assign node6054 = (inp[6]) ? node6058 : node6055;
														assign node6055 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node6058 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node6061 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node6064 = (inp[10]) ? node6072 : node6065;
												assign node6065 = (inp[13]) ? node6069 : node6066;
													assign node6066 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node6069 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node6072 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000001111111;
								assign node6075 = (inp[14]) ? node6169 : node6076;
									assign node6076 = (inp[2]) ? node6124 : node6077;
										assign node6077 = (inp[9]) ? node6105 : node6078;
											assign node6078 = (inp[0]) ? node6092 : node6079;
												assign node6079 = (inp[3]) ? node6083 : node6080;
													assign node6080 = (inp[13]) ? 16'b0000011111111111 : 16'b0001111111111111;
													assign node6083 = (inp[6]) ? 16'b0000001111111111 : node6084;
														assign node6084 = (inp[5]) ? node6086 : 16'b0000111111111111;
															assign node6086 = (inp[13]) ? 16'b0000011111111111 : node6087;
																assign node6087 = (inp[10]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node6092 = (inp[5]) ? node6098 : node6093;
													assign node6093 = (inp[3]) ? node6095 : 16'b0000111111111111;
														assign node6095 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node6098 = (inp[10]) ? node6100 : 16'b0000001111111111;
														assign node6100 = (inp[3]) ? 16'b0000001111111111 : node6101;
															assign node6101 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node6105 = (inp[6]) ? node6113 : node6106;
												assign node6106 = (inp[10]) ? node6108 : 16'b0000011111111111;
													assign node6108 = (inp[3]) ? 16'b0000001111111111 : node6109;
														assign node6109 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node6113 = (inp[13]) ? node6121 : node6114;
													assign node6114 = (inp[10]) ? node6118 : node6115;
														assign node6115 = (inp[0]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node6118 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node6121 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node6124 = (inp[10]) ? node6148 : node6125;
											assign node6125 = (inp[9]) ? node6135 : node6126;
												assign node6126 = (inp[3]) ? node6132 : node6127;
													assign node6127 = (inp[6]) ? 16'b0000011111111111 : node6128;
														assign node6128 = (inp[5]) ? 16'b0000011111111111 : 16'b0001111111111111;
													assign node6132 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node6135 = (inp[6]) ? node6143 : node6136;
													assign node6136 = (inp[5]) ? node6138 : 16'b0000001111111111;
														assign node6138 = (inp[13]) ? node6140 : 16'b0000001111111111;
															assign node6140 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node6143 = (inp[13]) ? 16'b0000000011111111 : node6144;
														assign node6144 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node6148 = (inp[3]) ? node6162 : node6149;
												assign node6149 = (inp[0]) ? node6157 : node6150;
													assign node6150 = (inp[9]) ? node6154 : node6151;
														assign node6151 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node6154 = (inp[5]) ? 16'b0000000011111111 : 16'b0000001111111111;
													assign node6157 = (inp[5]) ? node6159 : 16'b0000000111111111;
														assign node6159 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node6162 = (inp[13]) ? node6166 : node6163;
													assign node6163 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node6166 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node6169 = (inp[3]) ? node6217 : node6170;
										assign node6170 = (inp[0]) ? node6192 : node6171;
											assign node6171 = (inp[2]) ? node6189 : node6172;
												assign node6172 = (inp[9]) ? node6180 : node6173;
													assign node6173 = (inp[13]) ? node6177 : node6174;
														assign node6174 = (inp[6]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node6177 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node6180 = (inp[10]) ? node6186 : node6181;
														assign node6181 = (inp[6]) ? 16'b0000001111111111 : node6182;
															assign node6182 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node6186 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node6189 = (inp[6]) ? 16'b0000000011111111 : 16'b0000001111111111;
											assign node6192 = (inp[5]) ? node6208 : node6193;
												assign node6193 = (inp[9]) ? node6201 : node6194;
													assign node6194 = (inp[6]) ? node6198 : node6195;
														assign node6195 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node6198 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node6201 = (inp[6]) ? node6205 : node6202;
														assign node6202 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node6205 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node6208 = (inp[9]) ? node6214 : node6209;
													assign node6209 = (inp[2]) ? 16'b0000000011111111 : node6210;
														assign node6210 = (inp[6]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node6214 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000001111111;
										assign node6217 = (inp[10]) ? node6229 : node6218;
											assign node6218 = (inp[2]) ? node6222 : node6219;
												assign node6219 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node6222 = (inp[6]) ? node6224 : 16'b0000000111111111;
													assign node6224 = (inp[13]) ? 16'b0000000011111111 : node6225;
														assign node6225 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node6229 = (inp[9]) ? node6241 : node6230;
												assign node6230 = (inp[6]) ? node6236 : node6231;
													assign node6231 = (inp[5]) ? node6233 : 16'b0000000111111111;
														assign node6233 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node6236 = (inp[13]) ? 16'b0000000011111111 : node6237;
														assign node6237 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node6241 = (inp[0]) ? node6249 : node6242;
													assign node6242 = (inp[13]) ? node6246 : node6243;
														assign node6243 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node6246 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000001111111;
													assign node6249 = (inp[13]) ? 16'b0000000001111111 : node6250;
														assign node6250 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
							assign node6254 = (inp[13]) ? node6450 : node6255;
								assign node6255 = (inp[2]) ? node6373 : node6256;
									assign node6256 = (inp[8]) ? node6304 : node6257;
										assign node6257 = (inp[6]) ? node6283 : node6258;
											assign node6258 = (inp[14]) ? node6270 : node6259;
												assign node6259 = (inp[0]) ? node6263 : node6260;
													assign node6260 = (inp[3]) ? 16'b0000111111111111 : 16'b0011111111111111;
													assign node6263 = (inp[10]) ? node6267 : node6264;
														assign node6264 = (inp[3]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node6267 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node6270 = (inp[9]) ? node6278 : node6271;
													assign node6271 = (inp[0]) ? 16'b0000011111111111 : node6272;
														assign node6272 = (inp[3]) ? 16'b0000011111111111 : node6273;
															assign node6273 = (inp[5]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node6278 = (inp[0]) ? 16'b0000000111111111 : node6279;
														assign node6279 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node6283 = (inp[5]) ? node6291 : node6284;
												assign node6284 = (inp[0]) ? node6288 : node6285;
													assign node6285 = (inp[10]) ? 16'b0000001111111111 : 16'b0000111111111111;
													assign node6288 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node6291 = (inp[14]) ? node6301 : node6292;
													assign node6292 = (inp[9]) ? node6296 : node6293;
														assign node6293 = (inp[0]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node6296 = (inp[0]) ? 16'b0000000111111111 : node6297;
															assign node6297 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node6301 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node6304 = (inp[14]) ? node6344 : node6305;
											assign node6305 = (inp[10]) ? node6325 : node6306;
												assign node6306 = (inp[6]) ? node6318 : node6307;
													assign node6307 = (inp[0]) ? node6313 : node6308;
														assign node6308 = (inp[3]) ? node6310 : 16'b0001111111111111;
															assign node6310 = (inp[5]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node6313 = (inp[9]) ? node6315 : 16'b0000011111111111;
															assign node6315 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node6318 = (inp[0]) ? node6322 : node6319;
														assign node6319 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node6322 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node6325 = (inp[9]) ? node6341 : node6326;
													assign node6326 = (inp[6]) ? node6332 : node6327;
														assign node6327 = (inp[5]) ? 16'b0000001111111111 : node6328;
															assign node6328 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node6332 = (inp[0]) ? 16'b0000000111111111 : node6333;
															assign node6333 = (inp[5]) ? node6337 : node6334;
																assign node6334 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
																assign node6337 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node6341 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node6344 = (inp[3]) ? node6362 : node6345;
												assign node6345 = (inp[9]) ? node6353 : node6346;
													assign node6346 = (inp[5]) ? node6348 : 16'b0000011111111111;
														assign node6348 = (inp[6]) ? node6350 : 16'b0000001111111111;
															assign node6350 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node6353 = (inp[0]) ? node6357 : node6354;
														assign node6354 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node6357 = (inp[6]) ? node6359 : 16'b0000000111111111;
															assign node6359 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node6362 = (inp[10]) ? node6368 : node6363;
													assign node6363 = (inp[9]) ? 16'b0000000011111111 : node6364;
														assign node6364 = (inp[6]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node6368 = (inp[5]) ? 16'b0000000011111111 : node6369;
														assign node6369 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node6373 = (inp[10]) ? node6405 : node6374;
										assign node6374 = (inp[5]) ? node6396 : node6375;
											assign node6375 = (inp[8]) ? node6383 : node6376;
												assign node6376 = (inp[9]) ? node6380 : node6377;
													assign node6377 = (inp[14]) ? 16'b0000001111111111 : 16'b0000111111111111;
													assign node6380 = (inp[0]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node6383 = (inp[6]) ? node6391 : node6384;
													assign node6384 = (inp[0]) ? node6388 : node6385;
														assign node6385 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node6388 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node6391 = (inp[14]) ? node6393 : 16'b0000000111111111;
														assign node6393 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node6396 = (inp[6]) ? node6402 : node6397;
												assign node6397 = (inp[14]) ? 16'b0000000111111111 : node6398;
													assign node6398 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node6402 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000111111111;
										assign node6405 = (inp[9]) ? node6415 : node6406;
											assign node6406 = (inp[3]) ? node6408 : 16'b0000000111111111;
												assign node6408 = (inp[14]) ? node6410 : 16'b0000000111111111;
													assign node6410 = (inp[5]) ? 16'b0000000011111111 : node6411;
														assign node6411 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node6415 = (inp[6]) ? node6433 : node6416;
												assign node6416 = (inp[5]) ? node6426 : node6417;
													assign node6417 = (inp[14]) ? node6421 : node6418;
														assign node6418 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node6421 = (inp[8]) ? node6423 : 16'b0000000111111111;
															assign node6423 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node6426 = (inp[8]) ? 16'b0000000011111111 : node6427;
														assign node6427 = (inp[3]) ? 16'b0000000011111111 : node6428;
															assign node6428 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node6433 = (inp[0]) ? node6445 : node6434;
													assign node6434 = (inp[8]) ? node6440 : node6435;
														assign node6435 = (inp[14]) ? node6437 : 16'b0000000111111111;
															assign node6437 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node6440 = (inp[5]) ? node6442 : 16'b0000000011111111;
															assign node6442 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node6445 = (inp[14]) ? 16'b0000000001111111 : node6446;
														assign node6446 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
								assign node6450 = (inp[3]) ? node6516 : node6451;
									assign node6451 = (inp[5]) ? node6489 : node6452;
										assign node6452 = (inp[8]) ? node6482 : node6453;
											assign node6453 = (inp[9]) ? node6463 : node6454;
												assign node6454 = (inp[0]) ? node6456 : 16'b0000011111111111;
													assign node6456 = (inp[14]) ? node6458 : 16'b0000011111111111;
														assign node6458 = (inp[6]) ? 16'b0000001111111111 : node6459;
															assign node6459 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node6463 = (inp[6]) ? node6473 : node6464;
													assign node6464 = (inp[2]) ? node6466 : 16'b0000111111111111;
														assign node6466 = (inp[14]) ? 16'b0000000111111111 : node6467;
															assign node6467 = (inp[0]) ? 16'b0000001111111111 : node6468;
																assign node6468 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node6473 = (inp[10]) ? node6475 : 16'b0000001111111111;
														assign node6475 = (inp[0]) ? 16'b0000000111111111 : node6476;
															assign node6476 = (inp[14]) ? 16'b0000000111111111 : node6477;
																assign node6477 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node6482 = (inp[2]) ? node6484 : 16'b0000001111111111;
												assign node6484 = (inp[10]) ? 16'b0000000001111111 : node6485;
													assign node6485 = (inp[0]) ? 16'b0000000111111111 : 16'b0000000011111111;
										assign node6489 = (inp[6]) ? node6499 : node6490;
											assign node6490 = (inp[8]) ? 16'b0000000111111111 : node6491;
												assign node6491 = (inp[2]) ? node6493 : 16'b0000001111111111;
													assign node6493 = (inp[10]) ? 16'b0000000111111111 : node6494;
														assign node6494 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node6499 = (inp[8]) ? node6509 : node6500;
												assign node6500 = (inp[10]) ? node6504 : node6501;
													assign node6501 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node6504 = (inp[14]) ? 16'b0000000001111111 : node6505;
														assign node6505 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node6509 = (inp[14]) ? node6513 : node6510;
													assign node6510 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node6513 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node6516 = (inp[2]) ? node6564 : node6517;
										assign node6517 = (inp[6]) ? node6541 : node6518;
											assign node6518 = (inp[5]) ? node6526 : node6519;
												assign node6519 = (inp[9]) ? node6521 : 16'b0000001111111111;
													assign node6521 = (inp[8]) ? node6523 : 16'b0000001111111111;
														assign node6523 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node6526 = (inp[9]) ? node6536 : node6527;
													assign node6527 = (inp[8]) ? node6529 : 16'b0000000011111111;
														assign node6529 = (inp[10]) ? 16'b0000000111111111 : node6530;
															assign node6530 = (inp[14]) ? 16'b0000000111111111 : node6531;
																assign node6531 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node6536 = (inp[8]) ? 16'b0000000011111111 : node6537;
														assign node6537 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node6541 = (inp[8]) ? node6551 : node6542;
												assign node6542 = (inp[0]) ? node6548 : node6543;
													assign node6543 = (inp[14]) ? 16'b0000000111111111 : node6544;
														assign node6544 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node6548 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node6551 = (inp[9]) ? node6557 : node6552;
													assign node6552 = (inp[5]) ? node6554 : 16'b0000000111111111;
														assign node6554 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node6557 = (inp[0]) ? node6559 : 16'b0000000001111111;
														assign node6559 = (inp[14]) ? node6561 : 16'b0000000001111111;
															assign node6561 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node6564 = (inp[8]) ? node6588 : node6565;
											assign node6565 = (inp[0]) ? node6577 : node6566;
												assign node6566 = (inp[6]) ? node6570 : node6567;
													assign node6567 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node6570 = (inp[5]) ? node6572 : 16'b0000000011111111;
														assign node6572 = (inp[10]) ? node6574 : 16'b0000000011111111;
															assign node6574 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node6577 = (inp[9]) ? node6585 : node6578;
													assign node6578 = (inp[6]) ? node6580 : 16'b0000000111111111;
														assign node6580 = (inp[5]) ? node6582 : 16'b0000000011111111;
															assign node6582 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node6585 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node6588 = (inp[9]) ? node6598 : node6589;
												assign node6589 = (inp[10]) ? node6593 : node6590;
													assign node6590 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node6593 = (inp[0]) ? node6595 : 16'b0000000001111111;
														assign node6595 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node6598 = (inp[5]) ? node6600 : 16'b0000000001111111;
													assign node6600 = (inp[6]) ? node6604 : node6601;
														assign node6601 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node6604 = (inp[0]) ? 16'b0000000000001111 : 16'b0000000000011111;
						assign node6607 = (inp[6]) ? node7031 : node6608;
							assign node6608 = (inp[3]) ? node6812 : node6609;
								assign node6609 = (inp[8]) ? node6743 : node6610;
									assign node6610 = (inp[13]) ? node6678 : node6611;
										assign node6611 = (inp[10]) ? node6649 : node6612;
											assign node6612 = (inp[9]) ? node6630 : node6613;
												assign node6613 = (inp[4]) ? node6627 : node6614;
													assign node6614 = (inp[14]) ? 16'b0000111111111111 : node6615;
														assign node6615 = (inp[2]) ? node6621 : node6616;
															assign node6616 = (inp[0]) ? 16'b0001111111111111 : node6617;
																assign node6617 = (inp[5]) ? 16'b0001111111111111 : 16'b0011111111111111;
															assign node6621 = (inp[5]) ? node6623 : 16'b0001111111111111;
																assign node6623 = (inp[0]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node6627 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node6630 = (inp[5]) ? node6640 : node6631;
													assign node6631 = (inp[0]) ? node6635 : node6632;
														assign node6632 = (inp[14]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node6635 = (inp[2]) ? node6637 : 16'b0000011111111111;
															assign node6637 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node6640 = (inp[4]) ? node6646 : node6641;
														assign node6641 = (inp[2]) ? 16'b0000001111111111 : node6642;
															assign node6642 = (inp[0]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node6646 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node6649 = (inp[2]) ? node6663 : node6650;
												assign node6650 = (inp[5]) ? 16'b0000001111111111 : node6651;
													assign node6651 = (inp[0]) ? node6653 : 16'b0000111111111111;
														assign node6653 = (inp[9]) ? node6659 : node6654;
															assign node6654 = (inp[4]) ? node6656 : 16'b0000011111111111;
																assign node6656 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
															assign node6659 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node6663 = (inp[14]) ? node6675 : node6664;
													assign node6664 = (inp[0]) ? node6668 : node6665;
														assign node6665 = (inp[9]) ? 16'b0000011111111111 : 16'b0000001111111111;
														assign node6668 = (inp[5]) ? 16'b0000000111111111 : node6669;
															assign node6669 = (inp[4]) ? node6671 : 16'b0000001111111111;
																assign node6671 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node6675 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node6678 = (inp[2]) ? node6710 : node6679;
											assign node6679 = (inp[4]) ? node6695 : node6680;
												assign node6680 = (inp[10]) ? node6690 : node6681;
													assign node6681 = (inp[9]) ? node6687 : node6682;
														assign node6682 = (inp[5]) ? 16'b0000011111111111 : node6683;
															assign node6683 = (inp[0]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node6687 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node6690 = (inp[14]) ? 16'b0000000111111111 : node6691;
														assign node6691 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node6695 = (inp[14]) ? node6701 : node6696;
													assign node6696 = (inp[0]) ? 16'b0000001111111111 : node6697;
														assign node6697 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node6701 = (inp[0]) ? node6707 : node6702;
														assign node6702 = (inp[10]) ? node6704 : 16'b0000001111111111;
															assign node6704 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node6707 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node6710 = (inp[14]) ? node6728 : node6711;
												assign node6711 = (inp[5]) ? node6717 : node6712;
													assign node6712 = (inp[0]) ? 16'b0000001111111111 : node6713;
														assign node6713 = (inp[4]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node6717 = (inp[0]) ? node6725 : node6718;
														assign node6718 = (inp[10]) ? node6720 : 16'b0000001111111111;
															assign node6720 = (inp[9]) ? 16'b0000000111111111 : node6721;
																assign node6721 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node6725 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node6728 = (inp[4]) ? node6736 : node6729;
													assign node6729 = (inp[10]) ? 16'b0000000111111111 : node6730;
														assign node6730 = (inp[9]) ? 16'b0000000111111111 : node6731;
															assign node6731 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node6736 = (inp[10]) ? node6740 : node6737;
														assign node6737 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node6740 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node6743 = (inp[14]) ? node6777 : node6744;
										assign node6744 = (inp[4]) ? node6760 : node6745;
											assign node6745 = (inp[5]) ? node6753 : node6746;
												assign node6746 = (inp[9]) ? node6748 : 16'b0000111111111111;
													assign node6748 = (inp[2]) ? 16'b0000001111111111 : node6749;
														assign node6749 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node6753 = (inp[13]) ? node6755 : 16'b0000001111111111;
													assign node6755 = (inp[2]) ? 16'b0000000011111111 : node6756;
														assign node6756 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node6760 = (inp[5]) ? node6772 : node6761;
												assign node6761 = (inp[0]) ? node6765 : node6762;
													assign node6762 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node6765 = (inp[10]) ? node6767 : 16'b0000001111111111;
														assign node6767 = (inp[13]) ? node6769 : 16'b0000000111111111;
															assign node6769 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node6772 = (inp[0]) ? node6774 : 16'b0000000111111111;
													assign node6774 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node6777 = (inp[5]) ? node6799 : node6778;
											assign node6778 = (inp[10]) ? node6788 : node6779;
												assign node6779 = (inp[9]) ? node6785 : node6780;
													assign node6780 = (inp[4]) ? 16'b0000001111111111 : node6781;
														assign node6781 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node6785 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node6788 = (inp[2]) ? node6790 : 16'b0000000111111111;
													assign node6790 = (inp[4]) ? node6792 : 16'b0000000111111111;
														assign node6792 = (inp[13]) ? node6794 : 16'b0000000011111111;
															assign node6794 = (inp[0]) ? 16'b0000000001111111 : node6795;
																assign node6795 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node6799 = (inp[4]) ? node6809 : node6800;
												assign node6800 = (inp[9]) ? node6806 : node6801;
													assign node6801 = (inp[0]) ? node6803 : 16'b0000000111111111;
														assign node6803 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000111111111;
													assign node6806 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000001111111;
												assign node6809 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000000111111;
								assign node6812 = (inp[10]) ? node6916 : node6813;
									assign node6813 = (inp[5]) ? node6869 : node6814;
										assign node6814 = (inp[4]) ? node6834 : node6815;
											assign node6815 = (inp[9]) ? node6827 : node6816;
												assign node6816 = (inp[13]) ? node6822 : node6817;
													assign node6817 = (inp[14]) ? 16'b0000011111111111 : node6818;
														assign node6818 = (inp[8]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node6822 = (inp[2]) ? 16'b0000001111111111 : node6823;
														assign node6823 = (inp[0]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node6827 = (inp[8]) ? 16'b0000000111111111 : node6828;
													assign node6828 = (inp[13]) ? 16'b0000000111111111 : node6829;
														assign node6829 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node6834 = (inp[13]) ? node6854 : node6835;
												assign node6835 = (inp[9]) ? node6845 : node6836;
													assign node6836 = (inp[14]) ? node6842 : node6837;
														assign node6837 = (inp[0]) ? 16'b0000001111111111 : node6838;
															assign node6838 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node6842 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node6845 = (inp[8]) ? node6849 : node6846;
														assign node6846 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node6849 = (inp[14]) ? 16'b0000000011111111 : node6850;
															assign node6850 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node6854 = (inp[0]) ? node6864 : node6855;
													assign node6855 = (inp[2]) ? node6861 : node6856;
														assign node6856 = (inp[8]) ? 16'b0000000111111111 : node6857;
															assign node6857 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node6861 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node6864 = (inp[14]) ? 16'b0000000011111111 : node6865;
														assign node6865 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000111111111;
										assign node6869 = (inp[14]) ? node6895 : node6870;
											assign node6870 = (inp[0]) ? node6880 : node6871;
												assign node6871 = (inp[13]) ? node6875 : node6872;
													assign node6872 = (inp[9]) ? 16'b0000011111111111 : 16'b0000001111111111;
													assign node6875 = (inp[4]) ? 16'b0000000111111111 : node6876;
														assign node6876 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node6880 = (inp[9]) ? node6888 : node6881;
													assign node6881 = (inp[4]) ? node6885 : node6882;
														assign node6882 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node6885 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node6888 = (inp[4]) ? node6890 : 16'b0000000011111111;
														assign node6890 = (inp[8]) ? node6892 : 16'b0000000011111111;
															assign node6892 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node6895 = (inp[8]) ? node6909 : node6896;
												assign node6896 = (inp[13]) ? node6898 : 16'b0000000111111111;
													assign node6898 = (inp[0]) ? node6902 : node6899;
														assign node6899 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node6902 = (inp[2]) ? 16'b0000000001111111 : node6903;
															assign node6903 = (inp[9]) ? node6905 : 16'b0000000011111111;
																assign node6905 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node6909 = (inp[13]) ? node6913 : node6910;
													assign node6910 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node6913 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node6916 = (inp[0]) ? node6972 : node6917;
										assign node6917 = (inp[14]) ? node6941 : node6918;
											assign node6918 = (inp[13]) ? node6930 : node6919;
												assign node6919 = (inp[2]) ? node6925 : node6920;
													assign node6920 = (inp[9]) ? node6922 : 16'b0000011111111111;
														assign node6922 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node6925 = (inp[8]) ? 16'b0000000111111111 : node6926;
														assign node6926 = (inp[4]) ? 16'b0000001111111111 : 16'b0000000111111111;
												assign node6930 = (inp[5]) ? node6936 : node6931;
													assign node6931 = (inp[2]) ? 16'b0000000111111111 : node6932;
														assign node6932 = (inp[9]) ? 16'b0000000111111111 : 16'b0000011111111111;
													assign node6936 = (inp[9]) ? node6938 : 16'b0000000011111111;
														assign node6938 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node6941 = (inp[2]) ? node6953 : node6942;
												assign node6942 = (inp[9]) ? node6946 : node6943;
													assign node6943 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node6946 = (inp[4]) ? node6950 : node6947;
														assign node6947 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node6950 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node6953 = (inp[4]) ? node6961 : node6954;
													assign node6954 = (inp[13]) ? 16'b0000000001111111 : node6955;
														assign node6955 = (inp[8]) ? 16'b0000000011111111 : node6956;
															assign node6956 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node6961 = (inp[5]) ? node6965 : node6962;
														assign node6962 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node6965 = (inp[9]) ? 16'b0000000000111111 : node6966;
															assign node6966 = (inp[8]) ? node6968 : 16'b0000000001111111;
																assign node6968 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node6972 = (inp[9]) ? node7000 : node6973;
											assign node6973 = (inp[2]) ? node6985 : node6974;
												assign node6974 = (inp[4]) ? node6976 : 16'b0000000111111111;
													assign node6976 = (inp[5]) ? node6982 : node6977;
														assign node6977 = (inp[8]) ? 16'b0000000011111111 : node6978;
															assign node6978 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node6982 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node6985 = (inp[14]) ? node6991 : node6986;
													assign node6986 = (inp[8]) ? node6988 : 16'b0000000011111111;
														assign node6988 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000001111111;
													assign node6991 = (inp[5]) ? node6995 : node6992;
														assign node6992 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node6995 = (inp[4]) ? node6997 : 16'b0000000001111111;
															assign node6997 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node7000 = (inp[13]) ? node7018 : node7001;
												assign node7001 = (inp[2]) ? node7009 : node7002;
													assign node7002 = (inp[5]) ? node7004 : 16'b0000000011111111;
														assign node7004 = (inp[14]) ? node7006 : 16'b0000000011111111;
															assign node7006 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node7009 = (inp[14]) ? node7011 : 16'b0000000011111111;
														assign node7011 = (inp[5]) ? 16'b0000000000111111 : node7012;
															assign node7012 = (inp[8]) ? node7014 : 16'b0000000001111111;
																assign node7014 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node7018 = (inp[14]) ? node7024 : node7019;
													assign node7019 = (inp[5]) ? node7021 : 16'b0000000001111111;
														assign node7021 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node7024 = (inp[8]) ? node7028 : node7025;
														assign node7025 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node7028 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
							assign node7031 = (inp[9]) ? node7211 : node7032;
								assign node7032 = (inp[13]) ? node7116 : node7033;
									assign node7033 = (inp[14]) ? node7073 : node7034;
										assign node7034 = (inp[10]) ? node7056 : node7035;
											assign node7035 = (inp[0]) ? node7053 : node7036;
												assign node7036 = (inp[5]) ? node7044 : node7037;
													assign node7037 = (inp[3]) ? node7041 : node7038;
														assign node7038 = (inp[8]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node7041 = (inp[4]) ? 16'b0000011111111111 : 16'b0000001111111111;
													assign node7044 = (inp[8]) ? node7050 : node7045;
														assign node7045 = (inp[4]) ? 16'b0000001111111111 : node7046;
															assign node7046 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node7050 = (inp[3]) ? 16'b0000000011111111 : 16'b0000001111111111;
												assign node7053 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node7056 = (inp[4]) ? 16'b0000000111111111 : node7057;
												assign node7057 = (inp[5]) ? node7067 : node7058;
													assign node7058 = (inp[0]) ? node7064 : node7059;
														assign node7059 = (inp[8]) ? 16'b0000001111111111 : node7060;
															assign node7060 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node7064 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node7067 = (inp[3]) ? node7069 : 16'b0000001111111111;
														assign node7069 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node7073 = (inp[0]) ? node7097 : node7074;
											assign node7074 = (inp[5]) ? node7088 : node7075;
												assign node7075 = (inp[2]) ? node7081 : node7076;
													assign node7076 = (inp[3]) ? node7078 : 16'b0000001111111111;
														assign node7078 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node7081 = (inp[8]) ? 16'b0000000111111111 : node7082;
														assign node7082 = (inp[3]) ? 16'b0000000111111111 : node7083;
															assign node7083 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node7088 = (inp[4]) ? node7090 : 16'b0000000111111111;
													assign node7090 = (inp[8]) ? 16'b0000000011111111 : node7091;
														assign node7091 = (inp[3]) ? 16'b0000000011111111 : node7092;
															assign node7092 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node7097 = (inp[8]) ? node7105 : node7098;
												assign node7098 = (inp[10]) ? node7100 : 16'b0000001111111111;
													assign node7100 = (inp[3]) ? 16'b0000000011111111 : node7101;
														assign node7101 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node7105 = (inp[4]) ? node7107 : 16'b0000000011111111;
													assign node7107 = (inp[10]) ? 16'b0000000001111111 : node7108;
														assign node7108 = (inp[5]) ? 16'b0000000001111111 : node7109;
															assign node7109 = (inp[3]) ? node7111 : 16'b0000000011111111;
																assign node7111 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node7116 = (inp[2]) ? node7168 : node7117;
										assign node7117 = (inp[3]) ? node7137 : node7118;
											assign node7118 = (inp[4]) ? node7126 : node7119;
												assign node7119 = (inp[5]) ? node7121 : 16'b0000001111111111;
													assign node7121 = (inp[0]) ? 16'b0000001111111111 : node7122;
														assign node7122 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node7126 = (inp[8]) ? node7132 : node7127;
													assign node7127 = (inp[10]) ? 16'b0000000111111111 : node7128;
														assign node7128 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node7132 = (inp[0]) ? 16'b0000000011111111 : node7133;
														assign node7133 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node7137 = (inp[14]) ? node7155 : node7138;
												assign node7138 = (inp[5]) ? node7144 : node7139;
													assign node7139 = (inp[4]) ? 16'b0000000111111111 : node7140;
														assign node7140 = (inp[8]) ? 16'b0000000111111111 : 16'b0000011111111111;
													assign node7144 = (inp[4]) ? node7152 : node7145;
														assign node7145 = (inp[8]) ? 16'b0000000011111111 : node7146;
															assign node7146 = (inp[10]) ? node7148 : 16'b0000000111111111;
																assign node7148 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node7152 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node7155 = (inp[10]) ? node7163 : node7156;
													assign node7156 = (inp[0]) ? node7158 : 16'b0000000011111111;
														assign node7158 = (inp[5]) ? node7160 : 16'b0000000011111111;
															assign node7160 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node7163 = (inp[5]) ? 16'b0000000001111111 : node7164;
														assign node7164 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node7168 = (inp[10]) ? node7186 : node7169;
											assign node7169 = (inp[8]) ? node7175 : node7170;
												assign node7170 = (inp[3]) ? 16'b0000000111111111 : node7171;
													assign node7171 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node7175 = (inp[5]) ? node7181 : node7176;
													assign node7176 = (inp[14]) ? 16'b0000000001111111 : node7177;
														assign node7177 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node7181 = (inp[0]) ? 16'b0000000001111111 : node7182;
														assign node7182 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node7186 = (inp[5]) ? node7196 : node7187;
												assign node7187 = (inp[3]) ? node7189 : 16'b0000000011111111;
													assign node7189 = (inp[0]) ? 16'b0000000001111111 : node7190;
														assign node7190 = (inp[14]) ? 16'b0000000001111111 : node7191;
															assign node7191 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node7196 = (inp[0]) ? node7202 : node7197;
													assign node7197 = (inp[8]) ? node7199 : 16'b0000000001111111;
														assign node7199 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000011111111;
													assign node7202 = (inp[3]) ? node7208 : node7203;
														assign node7203 = (inp[8]) ? 16'b0000000000111111 : node7204;
															assign node7204 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node7208 = (inp[4]) ? 16'b0000000000011111 : 16'b0000000000111111;
								assign node7211 = (inp[3]) ? node7317 : node7212;
									assign node7212 = (inp[5]) ? node7264 : node7213;
										assign node7213 = (inp[10]) ? node7235 : node7214;
											assign node7214 = (inp[4]) ? node7230 : node7215;
												assign node7215 = (inp[2]) ? 16'b0000000111111111 : node7216;
													assign node7216 = (inp[14]) ? node7220 : node7217;
														assign node7217 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node7220 = (inp[0]) ? node7226 : node7221;
															assign node7221 = (inp[8]) ? node7223 : 16'b0000001111111111;
																assign node7223 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
															assign node7226 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node7230 = (inp[13]) ? node7232 : 16'b0000001111111111;
													assign node7232 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node7235 = (inp[13]) ? node7249 : node7236;
												assign node7236 = (inp[4]) ? node7242 : node7237;
													assign node7237 = (inp[14]) ? 16'b0000000011111111 : node7238;
														assign node7238 = (inp[8]) ? 16'b0000001111111111 : 16'b0000000111111111;
													assign node7242 = (inp[0]) ? 16'b0000000011111111 : node7243;
														assign node7243 = (inp[8]) ? 16'b0000000011111111 : node7244;
															assign node7244 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node7249 = (inp[14]) ? node7261 : node7250;
													assign node7250 = (inp[8]) ? node7258 : node7251;
														assign node7251 = (inp[2]) ? 16'b0000000011111111 : node7252;
															assign node7252 = (inp[4]) ? node7254 : 16'b0000000111111111;
																assign node7254 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node7258 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node7261 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node7264 = (inp[14]) ? node7294 : node7265;
											assign node7265 = (inp[13]) ? node7285 : node7266;
												assign node7266 = (inp[4]) ? node7276 : node7267;
													assign node7267 = (inp[8]) ? node7273 : node7268;
														assign node7268 = (inp[10]) ? 16'b0000000111111111 : node7269;
															assign node7269 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node7273 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node7276 = (inp[2]) ? node7280 : node7277;
														assign node7277 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node7280 = (inp[0]) ? node7282 : 16'b0000000011111111;
															assign node7282 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node7285 = (inp[4]) ? node7291 : node7286;
													assign node7286 = (inp[2]) ? node7288 : 16'b0000001111111111;
														assign node7288 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node7291 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node7294 = (inp[13]) ? node7304 : node7295;
												assign node7295 = (inp[2]) ? node7299 : node7296;
													assign node7296 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node7299 = (inp[4]) ? node7301 : 16'b0000000001111111;
														assign node7301 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node7304 = (inp[0]) ? node7310 : node7305;
													assign node7305 = (inp[2]) ? 16'b0000000000111111 : node7306;
														assign node7306 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node7310 = (inp[8]) ? 16'b0000000000011111 : node7311;
														assign node7311 = (inp[2]) ? 16'b0000000000111111 : node7312;
															assign node7312 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node7317 = (inp[10]) ? node7369 : node7318;
										assign node7318 = (inp[14]) ? node7342 : node7319;
											assign node7319 = (inp[8]) ? node7335 : node7320;
												assign node7320 = (inp[5]) ? node7330 : node7321;
													assign node7321 = (inp[0]) ? node7327 : node7322;
														assign node7322 = (inp[13]) ? 16'b0000000111111111 : node7323;
															assign node7323 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node7327 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node7330 = (inp[4]) ? node7332 : 16'b0000000011111111;
														assign node7332 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000011111111;
												assign node7335 = (inp[0]) ? node7337 : 16'b0000000011111111;
													assign node7337 = (inp[5]) ? 16'b0000000001111111 : node7338;
														assign node7338 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node7342 = (inp[4]) ? node7354 : node7343;
												assign node7343 = (inp[0]) ? node7349 : node7344;
													assign node7344 = (inp[2]) ? 16'b0000000011111111 : node7345;
														assign node7345 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node7349 = (inp[2]) ? node7351 : 16'b0000000011111111;
														assign node7351 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node7354 = (inp[2]) ? node7360 : node7355;
													assign node7355 = (inp[8]) ? 16'b0000000000111111 : node7356;
														assign node7356 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node7360 = (inp[13]) ? node7362 : 16'b0000000000111111;
														assign node7362 = (inp[8]) ? node7364 : 16'b0000000000111111;
															assign node7364 = (inp[5]) ? node7366 : 16'b0000000000011111;
																assign node7366 = (inp[0]) ? 16'b0000000000001111 : 16'b0000000000011111;
										assign node7369 = (inp[0]) ? node7393 : node7370;
											assign node7370 = (inp[2]) ? node7382 : node7371;
												assign node7371 = (inp[8]) ? node7377 : node7372;
													assign node7372 = (inp[13]) ? node7374 : 16'b0000000011111111;
														assign node7374 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node7377 = (inp[5]) ? node7379 : 16'b0000000001111111;
														assign node7379 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node7382 = (inp[14]) ? node7390 : node7383;
													assign node7383 = (inp[5]) ? node7387 : node7384;
														assign node7384 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node7387 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node7390 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000000011111;
											assign node7393 = (inp[4]) ? node7399 : node7394;
												assign node7394 = (inp[14]) ? 16'b0000000000111111 : node7395;
													assign node7395 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node7399 = (inp[13]) ? node7403 : node7400;
													assign node7400 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node7403 = (inp[14]) ? node7407 : node7404;
														assign node7404 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node7407 = (inp[2]) ? node7409 : 16'b0000000000011111;
															assign node7409 = (inp[5]) ? 16'b0000000000000111 : 16'b0000000000001111;
					assign node7412 = (inp[13]) ? node8142 : node7413;
						assign node7413 = (inp[1]) ? node7759 : node7414;
							assign node7414 = (inp[0]) ? node7576 : node7415;
								assign node7415 = (inp[9]) ? node7493 : node7416;
									assign node7416 = (inp[14]) ? node7452 : node7417;
										assign node7417 = (inp[6]) ? node7441 : node7418;
											assign node7418 = (inp[10]) ? node7432 : node7419;
												assign node7419 = (inp[5]) ? node7427 : node7420;
													assign node7420 = (inp[4]) ? node7422 : 16'b0001111111111111;
														assign node7422 = (inp[3]) ? node7424 : 16'b0000111111111111;
															assign node7424 = (inp[8]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node7427 = (inp[4]) ? 16'b0000011111111111 : node7428;
														assign node7428 = (inp[3]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node7432 = (inp[4]) ? 16'b0000000111111111 : node7433;
													assign node7433 = (inp[2]) ? 16'b0000001111111111 : node7434;
														assign node7434 = (inp[5]) ? 16'b0000011111111111 : node7435;
															assign node7435 = (inp[3]) ? 16'b0000011111111111 : 16'b0000111111111111;
											assign node7441 = (inp[3]) ? node7445 : node7442;
												assign node7442 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node7445 = (inp[4]) ? node7447 : 16'b0000001111111111;
													assign node7447 = (inp[10]) ? 16'b0000000111111111 : node7448;
														assign node7448 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node7452 = (inp[10]) ? node7468 : node7453;
											assign node7453 = (inp[2]) ? node7461 : node7454;
												assign node7454 = (inp[4]) ? 16'b0000001111111111 : node7455;
													assign node7455 = (inp[8]) ? 16'b0000001111111111 : node7456;
														assign node7456 = (inp[5]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node7461 = (inp[8]) ? node7463 : 16'b0000001111111111;
													assign node7463 = (inp[3]) ? 16'b0000000111111111 : node7464;
														assign node7464 = (inp[6]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node7468 = (inp[6]) ? node7482 : node7469;
												assign node7469 = (inp[4]) ? node7475 : node7470;
													assign node7470 = (inp[3]) ? 16'b0000001111111111 : node7471;
														assign node7471 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node7475 = (inp[5]) ? node7477 : 16'b0000001111111111;
														assign node7477 = (inp[2]) ? node7479 : 16'b0000000111111111;
															assign node7479 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node7482 = (inp[2]) ? node7488 : node7483;
													assign node7483 = (inp[3]) ? node7485 : 16'b0000000111111111;
														assign node7485 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node7488 = (inp[8]) ? node7490 : 16'b0000000011111111;
														assign node7490 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node7493 = (inp[5]) ? node7535 : node7494;
										assign node7494 = (inp[6]) ? node7518 : node7495;
											assign node7495 = (inp[14]) ? node7511 : node7496;
												assign node7496 = (inp[3]) ? node7502 : node7497;
													assign node7497 = (inp[10]) ? node7499 : 16'b0000111111111111;
														assign node7499 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node7502 = (inp[8]) ? node7504 : 16'b0000001111111111;
														assign node7504 = (inp[4]) ? node7506 : 16'b0000001111111111;
															assign node7506 = (inp[10]) ? 16'b0000000111111111 : node7507;
																assign node7507 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node7511 = (inp[4]) ? 16'b0000000111111111 : node7512;
													assign node7512 = (inp[10]) ? node7514 : 16'b0000001111111111;
														assign node7514 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node7518 = (inp[8]) ? node7526 : node7519;
												assign node7519 = (inp[3]) ? node7523 : node7520;
													assign node7520 = (inp[4]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node7523 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node7526 = (inp[2]) ? 16'b0000000011111111 : node7527;
													assign node7527 = (inp[10]) ? node7531 : node7528;
														assign node7528 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node7531 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node7535 = (inp[2]) ? node7561 : node7536;
											assign node7536 = (inp[10]) ? node7548 : node7537;
												assign node7537 = (inp[3]) ? 16'b0000000111111111 : node7538;
													assign node7538 = (inp[4]) ? node7540 : 16'b0000000111111111;
														assign node7540 = (inp[6]) ? node7542 : 16'b0000000111111111;
															assign node7542 = (inp[14]) ? node7544 : 16'b0000000111111111;
																assign node7544 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node7548 = (inp[4]) ? node7558 : node7549;
													assign node7549 = (inp[6]) ? 16'b0000000011111111 : node7550;
														assign node7550 = (inp[14]) ? 16'b0000000111111111 : node7551;
															assign node7551 = (inp[3]) ? node7553 : 16'b0000001111111111;
																assign node7553 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node7558 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node7561 = (inp[4]) ? node7565 : node7562;
												assign node7562 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node7565 = (inp[10]) ? node7569 : node7566;
													assign node7566 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node7569 = (inp[6]) ? node7573 : node7570;
														assign node7570 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000001111111;
														assign node7573 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
								assign node7576 = (inp[10]) ? node7666 : node7577;
									assign node7577 = (inp[3]) ? node7629 : node7578;
										assign node7578 = (inp[2]) ? node7602 : node7579;
											assign node7579 = (inp[6]) ? node7589 : node7580;
												assign node7580 = (inp[5]) ? node7586 : node7581;
													assign node7581 = (inp[8]) ? 16'b0000011111111111 : node7582;
														assign node7582 = (inp[4]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node7586 = (inp[9]) ? 16'b0000011111111111 : 16'b0000001111111111;
												assign node7589 = (inp[5]) ? node7599 : node7590;
													assign node7590 = (inp[14]) ? node7596 : node7591;
														assign node7591 = (inp[9]) ? node7593 : 16'b0000111111111111;
															assign node7593 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node7596 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node7599 = (inp[4]) ? 16'b0000000111111111 : 16'b0000000011111111;
											assign node7602 = (inp[9]) ? node7614 : node7603;
												assign node7603 = (inp[8]) ? node7609 : node7604;
													assign node7604 = (inp[4]) ? node7606 : 16'b0000111111111111;
														assign node7606 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node7609 = (inp[14]) ? 16'b0000000111111111 : node7610;
														assign node7610 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node7614 = (inp[5]) ? node7624 : node7615;
													assign node7615 = (inp[14]) ? node7617 : 16'b0000000111111111;
														assign node7617 = (inp[6]) ? node7619 : 16'b0000000111111111;
															assign node7619 = (inp[8]) ? 16'b0000000011111111 : node7620;
																assign node7620 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node7624 = (inp[4]) ? node7626 : 16'b0000000011111111;
														assign node7626 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node7629 = (inp[4]) ? node7643 : node7630;
											assign node7630 = (inp[6]) ? node7636 : node7631;
												assign node7631 = (inp[5]) ? node7633 : 16'b0000011111111111;
													assign node7633 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node7636 = (inp[5]) ? node7638 : 16'b0000000111111111;
													assign node7638 = (inp[2]) ? node7640 : 16'b0000000111111111;
														assign node7640 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node7643 = (inp[9]) ? node7659 : node7644;
												assign node7644 = (inp[14]) ? node7650 : node7645;
													assign node7645 = (inp[5]) ? 16'b0000000111111111 : node7646;
														assign node7646 = (inp[2]) ? 16'b0000001111111111 : 16'b0000000111111111;
													assign node7650 = (inp[8]) ? node7654 : node7651;
														assign node7651 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node7654 = (inp[6]) ? node7656 : 16'b0000000011111111;
															assign node7656 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node7659 = (inp[8]) ? node7663 : node7660;
													assign node7660 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node7663 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node7666 = (inp[2]) ? node7708 : node7667;
										assign node7667 = (inp[14]) ? node7693 : node7668;
											assign node7668 = (inp[5]) ? node7684 : node7669;
												assign node7669 = (inp[8]) ? node7675 : node7670;
													assign node7670 = (inp[3]) ? 16'b0000001111111111 : node7671;
														assign node7671 = (inp[4]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node7675 = (inp[6]) ? 16'b0000000011111111 : node7676;
														assign node7676 = (inp[9]) ? 16'b0000000111111111 : node7677;
															assign node7677 = (inp[4]) ? node7679 : 16'b0000001111111111;
																assign node7679 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node7684 = (inp[9]) ? 16'b0000000011111111 : node7685;
													assign node7685 = (inp[8]) ? 16'b0000000011111111 : node7686;
														assign node7686 = (inp[3]) ? 16'b0000000111111111 : node7687;
															assign node7687 = (inp[6]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node7693 = (inp[9]) ? node7699 : node7694;
												assign node7694 = (inp[5]) ? node7696 : 16'b0000000111111111;
													assign node7696 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node7699 = (inp[3]) ? node7701 : 16'b0000000111111111;
													assign node7701 = (inp[5]) ? node7703 : 16'b0000000001111111;
														assign node7703 = (inp[8]) ? 16'b0000000000011111 : node7704;
															assign node7704 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node7708 = (inp[6]) ? node7736 : node7709;
											assign node7709 = (inp[8]) ? node7721 : node7710;
												assign node7710 = (inp[9]) ? node7712 : 16'b0000000111111111;
													assign node7712 = (inp[5]) ? node7716 : node7713;
														assign node7713 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node7716 = (inp[4]) ? 16'b0000000001111111 : node7717;
															assign node7717 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node7721 = (inp[4]) ? node7729 : node7722;
													assign node7722 = (inp[9]) ? 16'b0000000001111111 : node7723;
														assign node7723 = (inp[3]) ? 16'b0000000011111111 : node7724;
															assign node7724 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node7729 = (inp[5]) ? 16'b0000000001111111 : node7730;
														assign node7730 = (inp[14]) ? node7732 : 16'b0000000011111111;
															assign node7732 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node7736 = (inp[4]) ? node7740 : node7737;
												assign node7737 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node7740 = (inp[5]) ? node7750 : node7741;
													assign node7741 = (inp[3]) ? 16'b0000000000111111 : node7742;
														assign node7742 = (inp[14]) ? 16'b0000000001111111 : node7743;
															assign node7743 = (inp[8]) ? node7745 : 16'b0000000011111111;
																assign node7745 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node7750 = (inp[9]) ? node7756 : node7751;
														assign node7751 = (inp[8]) ? node7753 : 16'b0000000001111111;
															assign node7753 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node7756 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
							assign node7759 = (inp[9]) ? node7939 : node7760;
								assign node7760 = (inp[5]) ? node7864 : node7761;
									assign node7761 = (inp[3]) ? node7805 : node7762;
										assign node7762 = (inp[2]) ? node7780 : node7763;
											assign node7763 = (inp[10]) ? node7777 : node7764;
												assign node7764 = (inp[14]) ? node7768 : node7765;
													assign node7765 = (inp[8]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node7768 = (inp[0]) ? 16'b0000001111111111 : node7769;
														assign node7769 = (inp[6]) ? 16'b0000001111111111 : node7770;
															assign node7770 = (inp[4]) ? node7772 : 16'b0000011111111111;
																assign node7772 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node7777 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node7780 = (inp[14]) ? node7794 : node7781;
												assign node7781 = (inp[10]) ? node7787 : node7782;
													assign node7782 = (inp[8]) ? 16'b0000001111111111 : node7783;
														assign node7783 = (inp[0]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node7787 = (inp[8]) ? 16'b0000000111111111 : node7788;
														assign node7788 = (inp[4]) ? 16'b0000000111111111 : node7789;
															assign node7789 = (inp[6]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node7794 = (inp[4]) ? node7800 : node7795;
													assign node7795 = (inp[8]) ? 16'b0000000111111111 : node7796;
														assign node7796 = (inp[6]) ? 16'b0000000111111111 : 16'b0000011111111111;
													assign node7800 = (inp[8]) ? 16'b0000000011111111 : node7801;
														assign node7801 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node7805 = (inp[0]) ? node7837 : node7806;
											assign node7806 = (inp[2]) ? node7826 : node7807;
												assign node7807 = (inp[14]) ? node7821 : node7808;
													assign node7808 = (inp[6]) ? node7810 : 16'b0000011111111111;
														assign node7810 = (inp[8]) ? node7816 : node7811;
															assign node7811 = (inp[4]) ? node7813 : 16'b0000001111111111;
																assign node7813 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
															assign node7816 = (inp[4]) ? 16'b0000000111111111 : node7817;
																assign node7817 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node7821 = (inp[10]) ? 16'b0000000111111111 : node7822;
														assign node7822 = (inp[6]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node7826 = (inp[10]) ? node7828 : 16'b0000000111111111;
													assign node7828 = (inp[6]) ? node7832 : node7829;
														assign node7829 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node7832 = (inp[14]) ? node7834 : 16'b0000000011111111;
															assign node7834 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node7837 = (inp[2]) ? node7849 : node7838;
												assign node7838 = (inp[8]) ? node7840 : 16'b0000000111111111;
													assign node7840 = (inp[10]) ? node7844 : node7841;
														assign node7841 = (inp[6]) ? 16'b0000000011111111 : 16'b0000001111111111;
														assign node7844 = (inp[14]) ? node7846 : 16'b0000000011111111;
															assign node7846 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node7849 = (inp[6]) ? node7855 : node7850;
													assign node7850 = (inp[8]) ? node7852 : 16'b0000000011111111;
														assign node7852 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node7855 = (inp[4]) ? node7861 : node7856;
														assign node7856 = (inp[14]) ? 16'b0000000001111111 : node7857;
															assign node7857 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node7861 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node7864 = (inp[2]) ? node7908 : node7865;
										assign node7865 = (inp[10]) ? node7885 : node7866;
											assign node7866 = (inp[14]) ? node7874 : node7867;
												assign node7867 = (inp[4]) ? node7871 : node7868;
													assign node7868 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node7871 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node7874 = (inp[0]) ? node7880 : node7875;
													assign node7875 = (inp[3]) ? 16'b0000000111111111 : node7876;
														assign node7876 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node7880 = (inp[6]) ? node7882 : 16'b0000000111111111;
														assign node7882 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node7885 = (inp[8]) ? node7895 : node7886;
												assign node7886 = (inp[3]) ? 16'b0000000011111111 : node7887;
													assign node7887 = (inp[4]) ? 16'b0000000011111111 : node7888;
														assign node7888 = (inp[6]) ? node7890 : 16'b0000000111111111;
															assign node7890 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node7895 = (inp[4]) ? node7905 : node7896;
													assign node7896 = (inp[3]) ? node7902 : node7897;
														assign node7897 = (inp[14]) ? node7899 : 16'b0000001111111111;
															assign node7899 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node7902 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node7905 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node7908 = (inp[3]) ? node7924 : node7909;
											assign node7909 = (inp[6]) ? node7915 : node7910;
												assign node7910 = (inp[10]) ? 16'b0000000011111111 : node7911;
													assign node7911 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node7915 = (inp[14]) ? node7917 : 16'b0000000111111111;
													assign node7917 = (inp[0]) ? node7919 : 16'b0000000001111111;
														assign node7919 = (inp[10]) ? node7921 : 16'b0000000001111111;
															assign node7921 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node7924 = (inp[0]) ? node7930 : node7925;
												assign node7925 = (inp[10]) ? 16'b0000000001111111 : node7926;
													assign node7926 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000111111111;
												assign node7930 = (inp[4]) ? node7934 : node7931;
													assign node7931 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node7934 = (inp[14]) ? node7936 : 16'b0000000000111111;
														assign node7936 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000111111;
								assign node7939 = (inp[8]) ? node8063 : node7940;
									assign node7940 = (inp[3]) ? node8002 : node7941;
										assign node7941 = (inp[6]) ? node7971 : node7942;
											assign node7942 = (inp[10]) ? node7958 : node7943;
												assign node7943 = (inp[2]) ? node7951 : node7944;
													assign node7944 = (inp[0]) ? node7946 : 16'b0000001111111111;
														assign node7946 = (inp[4]) ? 16'b0000000111111111 : node7947;
															assign node7947 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node7951 = (inp[0]) ? 16'b0000000011111111 : node7952;
														assign node7952 = (inp[14]) ? 16'b0000000111111111 : node7953;
															assign node7953 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node7958 = (inp[5]) ? node7964 : node7959;
													assign node7959 = (inp[14]) ? 16'b0000000111111111 : node7960;
														assign node7960 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node7964 = (inp[14]) ? node7968 : node7965;
														assign node7965 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node7968 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node7971 = (inp[14]) ? node7987 : node7972;
												assign node7972 = (inp[0]) ? node7978 : node7973;
													assign node7973 = (inp[10]) ? node7975 : 16'b0000001111111111;
														assign node7975 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node7978 = (inp[10]) ? 16'b0000000011111111 : node7979;
														assign node7979 = (inp[4]) ? 16'b0000000011111111 : node7980;
															assign node7980 = (inp[5]) ? node7982 : 16'b0000000111111111;
																assign node7982 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node7987 = (inp[5]) ? node7993 : node7988;
													assign node7988 = (inp[0]) ? node7990 : 16'b0000000011111111;
														assign node7990 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node7993 = (inp[0]) ? node7995 : 16'b0000000001111111;
														assign node7995 = (inp[4]) ? node7997 : 16'b0000000001111111;
															assign node7997 = (inp[10]) ? 16'b0000000000111111 : node7998;
																assign node7998 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node8002 = (inp[0]) ? node8034 : node8003;
											assign node8003 = (inp[2]) ? node8019 : node8004;
												assign node8004 = (inp[10]) ? node8014 : node8005;
													assign node8005 = (inp[6]) ? node8009 : node8006;
														assign node8006 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node8009 = (inp[14]) ? node8011 : 16'b0000000111111111;
															assign node8011 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node8014 = (inp[6]) ? node8016 : 16'b0000000111111111;
														assign node8016 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node8019 = (inp[6]) ? node8029 : node8020;
													assign node8020 = (inp[4]) ? 16'b0000000011111111 : node8021;
														assign node8021 = (inp[14]) ? node8023 : 16'b0000000011111111;
															assign node8023 = (inp[10]) ? node8025 : 16'b0000000011111111;
																assign node8025 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node8029 = (inp[5]) ? node8031 : 16'b0000000011111111;
														assign node8031 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node8034 = (inp[6]) ? node8048 : node8035;
												assign node8035 = (inp[5]) ? node8041 : node8036;
													assign node8036 = (inp[14]) ? node8038 : 16'b0000000111111111;
														assign node8038 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node8041 = (inp[14]) ? node8045 : node8042;
														assign node8042 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node8045 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node8048 = (inp[14]) ? node8056 : node8049;
													assign node8049 = (inp[10]) ? node8053 : node8050;
														assign node8050 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node8053 = (inp[4]) ? 16'b0000000000011111 : 16'b0000000001111111;
													assign node8056 = (inp[5]) ? 16'b0000000000011111 : node8057;
														assign node8057 = (inp[2]) ? node8059 : 16'b0000000000111111;
															assign node8059 = (inp[4]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node8063 = (inp[10]) ? node8103 : node8064;
										assign node8064 = (inp[4]) ? node8076 : node8065;
											assign node8065 = (inp[14]) ? node8071 : node8066;
												assign node8066 = (inp[0]) ? 16'b0000000011111111 : node8067;
													assign node8067 = (inp[3]) ? 16'b0000001111111111 : 16'b0000000111111111;
												assign node8071 = (inp[6]) ? 16'b0000000001111111 : node8072;
													assign node8072 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node8076 = (inp[6]) ? node8092 : node8077;
												assign node8077 = (inp[2]) ? node8083 : node8078;
													assign node8078 = (inp[0]) ? node8080 : 16'b0000000011111111;
														assign node8080 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node8083 = (inp[5]) ? node8087 : node8084;
														assign node8084 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node8087 = (inp[0]) ? node8089 : 16'b0000000001111111;
															assign node8089 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node8092 = (inp[3]) ? 16'b0000000000111111 : node8093;
													assign node8093 = (inp[5]) ? node8095 : 16'b0000000001111111;
														assign node8095 = (inp[0]) ? 16'b0000000000111111 : node8096;
															assign node8096 = (inp[14]) ? node8098 : 16'b0000000001111111;
																assign node8098 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node8103 = (inp[0]) ? node8123 : node8104;
											assign node8104 = (inp[4]) ? node8114 : node8105;
												assign node8105 = (inp[5]) ? node8109 : node8106;
													assign node8106 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000111111111;
													assign node8109 = (inp[3]) ? 16'b0000000001111111 : node8110;
														assign node8110 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node8114 = (inp[14]) ? node8120 : node8115;
													assign node8115 = (inp[6]) ? node8117 : 16'b0000000001111111;
														assign node8117 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node8120 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node8123 = (inp[5]) ? node8133 : node8124;
												assign node8124 = (inp[6]) ? 16'b0000000000111111 : node8125;
													assign node8125 = (inp[4]) ? node8127 : 16'b0000000000111111;
														assign node8127 = (inp[14]) ? node8129 : 16'b0000000000111111;
															assign node8129 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node8133 = (inp[6]) ? node8135 : 16'b0000000000111111;
													assign node8135 = (inp[3]) ? node8137 : 16'b0000000000011111;
														assign node8137 = (inp[4]) ? node8139 : 16'b0000000000001111;
															assign node8139 = (inp[14]) ? 16'b0000000000000111 : 16'b0000000000001111;
						assign node8142 = (inp[6]) ? node8552 : node8143;
							assign node8143 = (inp[0]) ? node8357 : node8144;
								assign node8144 = (inp[5]) ? node8238 : node8145;
									assign node8145 = (inp[9]) ? node8185 : node8146;
										assign node8146 = (inp[3]) ? node8168 : node8147;
											assign node8147 = (inp[14]) ? node8157 : node8148;
												assign node8148 = (inp[2]) ? node8154 : node8149;
													assign node8149 = (inp[10]) ? 16'b0000011111111111 : node8150;
														assign node8150 = (inp[4]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node8154 = (inp[1]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node8157 = (inp[1]) ? node8165 : node8158;
													assign node8158 = (inp[4]) ? 16'b0000001111111111 : node8159;
														assign node8159 = (inp[2]) ? node8161 : 16'b0000011111111111;
															assign node8161 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node8165 = (inp[8]) ? 16'b0000000011111111 : 16'b0000001111111111;
											assign node8168 = (inp[14]) ? node8178 : node8169;
												assign node8169 = (inp[2]) ? 16'b0000000111111111 : node8170;
													assign node8170 = (inp[8]) ? node8174 : node8171;
														assign node8171 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node8174 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node8178 = (inp[10]) ? 16'b0000000000111111 : node8179;
													assign node8179 = (inp[1]) ? node8181 : 16'b0000000111111111;
														assign node8181 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node8185 = (inp[1]) ? node8207 : node8186;
											assign node8186 = (inp[8]) ? node8196 : node8187;
												assign node8187 = (inp[10]) ? node8193 : node8188;
													assign node8188 = (inp[4]) ? 16'b0000001111111111 : node8189;
														assign node8189 = (inp[14]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node8193 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node8196 = (inp[4]) ? node8200 : node8197;
													assign node8197 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node8200 = (inp[10]) ? node8204 : node8201;
														assign node8201 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node8204 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node8207 = (inp[2]) ? node8221 : node8208;
												assign node8208 = (inp[14]) ? 16'b0000000011111111 : node8209;
													assign node8209 = (inp[4]) ? node8215 : node8210;
														assign node8210 = (inp[10]) ? 16'b0000000111111111 : node8211;
															assign node8211 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node8215 = (inp[8]) ? node8217 : 16'b0000000111111111;
															assign node8217 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node8221 = (inp[8]) ? node8233 : node8222;
													assign node8222 = (inp[4]) ? node8228 : node8223;
														assign node8223 = (inp[10]) ? node8225 : 16'b0000000111111111;
															assign node8225 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node8228 = (inp[14]) ? node8230 : 16'b0000000011111111;
															assign node8230 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node8233 = (inp[10]) ? node8235 : 16'b0000000011111111;
														assign node8235 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node8238 = (inp[9]) ? node8302 : node8239;
										assign node8239 = (inp[3]) ? node8275 : node8240;
											assign node8240 = (inp[8]) ? node8256 : node8241;
												assign node8241 = (inp[2]) ? 16'b0000000111111111 : node8242;
													assign node8242 = (inp[1]) ? node8252 : node8243;
														assign node8243 = (inp[14]) ? node8247 : node8244;
															assign node8244 = (inp[10]) ? 16'b0000011111111111 : 16'b0000111111111111;
															assign node8247 = (inp[4]) ? 16'b0000001111111111 : node8248;
																assign node8248 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node8252 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node8256 = (inp[1]) ? node8270 : node8257;
													assign node8257 = (inp[10]) ? node8263 : node8258;
														assign node8258 = (inp[4]) ? 16'b0000000111111111 : node8259;
															assign node8259 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node8263 = (inp[14]) ? node8265 : 16'b0000000111111111;
															assign node8265 = (inp[2]) ? 16'b0000000011111111 : node8266;
																assign node8266 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node8270 = (inp[4]) ? node8272 : 16'b0000000011111111;
														assign node8272 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node8275 = (inp[2]) ? node8297 : node8276;
												assign node8276 = (inp[14]) ? node8290 : node8277;
													assign node8277 = (inp[4]) ? node8285 : node8278;
														assign node8278 = (inp[8]) ? node8280 : 16'b0000001111111111;
															assign node8280 = (inp[10]) ? node8282 : 16'b0000000111111111;
																assign node8282 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node8285 = (inp[10]) ? 16'b0000000011111111 : node8286;
															assign node8286 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node8290 = (inp[8]) ? node8294 : node8291;
														assign node8291 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node8294 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node8297 = (inp[8]) ? 16'b0000000001111111 : node8298;
													assign node8298 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000001111111;
										assign node8302 = (inp[4]) ? node8326 : node8303;
											assign node8303 = (inp[3]) ? node8315 : node8304;
												assign node8304 = (inp[1]) ? node8306 : 16'b0000000111111111;
													assign node8306 = (inp[2]) ? node8312 : node8307;
														assign node8307 = (inp[10]) ? node8309 : 16'b0000000111111111;
															assign node8309 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node8312 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node8315 = (inp[2]) ? node8321 : node8316;
													assign node8316 = (inp[10]) ? node8318 : 16'b0000000011111111;
														assign node8318 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node8321 = (inp[10]) ? 16'b0000000000011111 : node8322;
														assign node8322 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node8326 = (inp[14]) ? node8346 : node8327;
												assign node8327 = (inp[1]) ? node8339 : node8328;
													assign node8328 = (inp[10]) ? node8332 : node8329;
														assign node8329 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node8332 = (inp[8]) ? 16'b0000000001111111 : node8333;
															assign node8333 = (inp[2]) ? node8335 : 16'b0000000011111111;
																assign node8335 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node8339 = (inp[3]) ? 16'b0000000000111111 : node8340;
														assign node8340 = (inp[8]) ? 16'b0000000001111111 : node8341;
															assign node8341 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node8346 = (inp[3]) ? node8352 : node8347;
													assign node8347 = (inp[10]) ? node8349 : 16'b0000000001111111;
														assign node8349 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000001111111;
													assign node8352 = (inp[8]) ? 16'b0000000000111111 : node8353;
														assign node8353 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
								assign node8357 = (inp[10]) ? node8461 : node8358;
									assign node8358 = (inp[1]) ? node8398 : node8359;
										assign node8359 = (inp[8]) ? node8383 : node8360;
											assign node8360 = (inp[4]) ? node8370 : node8361;
												assign node8361 = (inp[9]) ? 16'b0000000111111111 : node8362;
													assign node8362 = (inp[2]) ? node8364 : 16'b0000011111111111;
														assign node8364 = (inp[3]) ? node8366 : 16'b0000001111111111;
															assign node8366 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node8370 = (inp[14]) ? node8380 : node8371;
													assign node8371 = (inp[2]) ? node8377 : node8372;
														assign node8372 = (inp[5]) ? 16'b0000000111111111 : node8373;
															assign node8373 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node8377 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node8380 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node8383 = (inp[9]) ? node8395 : node8384;
												assign node8384 = (inp[14]) ? 16'b0000000011111111 : node8385;
													assign node8385 = (inp[5]) ? node8389 : node8386;
														assign node8386 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node8389 = (inp[3]) ? 16'b0000000011111111 : node8390;
															assign node8390 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node8395 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node8398 = (inp[4]) ? node8426 : node8399;
											assign node8399 = (inp[8]) ? node8417 : node8400;
												assign node8400 = (inp[2]) ? node8408 : node8401;
													assign node8401 = (inp[3]) ? 16'b0000000011111111 : node8402;
														assign node8402 = (inp[14]) ? node8404 : 16'b0000001111111111;
															assign node8404 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node8408 = (inp[5]) ? node8414 : node8409;
														assign node8409 = (inp[14]) ? node8411 : 16'b0000000111111111;
															assign node8411 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node8414 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node8417 = (inp[9]) ? node8419 : 16'b0000000011111111;
													assign node8419 = (inp[3]) ? node8423 : node8420;
														assign node8420 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node8423 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node8426 = (inp[3]) ? node8446 : node8427;
												assign node8427 = (inp[5]) ? node8435 : node8428;
													assign node8428 = (inp[14]) ? node8432 : node8429;
														assign node8429 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node8432 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node8435 = (inp[14]) ? node8443 : node8436;
														assign node8436 = (inp[9]) ? 16'b0000000001111111 : node8437;
															assign node8437 = (inp[2]) ? node8439 : 16'b0000000011111111;
																assign node8439 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node8443 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node8446 = (inp[2]) ? node8456 : node8447;
													assign node8447 = (inp[5]) ? 16'b0000000001111111 : node8448;
														assign node8448 = (inp[8]) ? node8450 : 16'b0000000011111111;
															assign node8450 = (inp[9]) ? 16'b0000000000111111 : node8451;
																assign node8451 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node8456 = (inp[9]) ? node8458 : 16'b0000000000111111;
														assign node8458 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node8461 = (inp[5]) ? node8501 : node8462;
										assign node8462 = (inp[1]) ? node8484 : node8463;
											assign node8463 = (inp[9]) ? node8475 : node8464;
												assign node8464 = (inp[2]) ? node8466 : 16'b0000001111111111;
													assign node8466 = (inp[8]) ? node8470 : node8467;
														assign node8467 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node8470 = (inp[14]) ? node8472 : 16'b0000000011111111;
															assign node8472 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node8475 = (inp[3]) ? node8477 : 16'b0000000011111111;
													assign node8477 = (inp[4]) ? 16'b0000000001111111 : node8478;
														assign node8478 = (inp[14]) ? node8480 : 16'b0000000011111111;
															assign node8480 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node8484 = (inp[14]) ? node8494 : node8485;
												assign node8485 = (inp[3]) ? node8487 : 16'b0000000111111111;
													assign node8487 = (inp[4]) ? 16'b0000000000111111 : node8488;
														assign node8488 = (inp[8]) ? node8490 : 16'b0000000011111111;
															assign node8490 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node8494 = (inp[8]) ? 16'b0000000001111111 : node8495;
													assign node8495 = (inp[9]) ? node8497 : 16'b0000000001111111;
														assign node8497 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node8501 = (inp[2]) ? node8525 : node8502;
											assign node8502 = (inp[8]) ? node8514 : node8503;
												assign node8503 = (inp[3]) ? node8509 : node8504;
													assign node8504 = (inp[9]) ? 16'b0000000011111111 : node8505;
														assign node8505 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node8509 = (inp[4]) ? 16'b0000000001111111 : node8510;
														assign node8510 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node8514 = (inp[9]) ? node8522 : node8515;
													assign node8515 = (inp[14]) ? 16'b0000000000111111 : node8516;
														assign node8516 = (inp[1]) ? 16'b0000000001111111 : node8517;
															assign node8517 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node8522 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node8525 = (inp[3]) ? node8543 : node8526;
												assign node8526 = (inp[8]) ? node8534 : node8527;
													assign node8527 = (inp[1]) ? node8529 : 16'b0000000011111111;
														assign node8529 = (inp[9]) ? node8531 : 16'b0000000001111111;
															assign node8531 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node8534 = (inp[1]) ? 16'b0000000000011111 : node8535;
														assign node8535 = (inp[14]) ? 16'b0000000000111111 : node8536;
															assign node8536 = (inp[9]) ? node8538 : 16'b0000000001111111;
																assign node8538 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node8543 = (inp[8]) ? 16'b0000000000011111 : node8544;
													assign node8544 = (inp[4]) ? node8546 : 16'b0000000000111111;
														assign node8546 = (inp[9]) ? node8548 : 16'b0000000000111111;
															assign node8548 = (inp[1]) ? 16'b0000000000001111 : 16'b0000000000011111;
							assign node8552 = (inp[4]) ? node8778 : node8553;
								assign node8553 = (inp[1]) ? node8667 : node8554;
									assign node8554 = (inp[9]) ? node8618 : node8555;
										assign node8555 = (inp[8]) ? node8585 : node8556;
											assign node8556 = (inp[5]) ? node8574 : node8557;
												assign node8557 = (inp[14]) ? node8565 : node8558;
													assign node8558 = (inp[3]) ? node8562 : node8559;
														assign node8559 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node8562 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node8565 = (inp[2]) ? node8571 : node8566;
														assign node8566 = (inp[3]) ? 16'b0000000111111111 : node8567;
															assign node8567 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node8571 = (inp[10]) ? 16'b0000000111111111 : 16'b0000000011111111;
												assign node8574 = (inp[10]) ? node8580 : node8575;
													assign node8575 = (inp[14]) ? node8577 : 16'b0000000111111111;
														assign node8577 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node8580 = (inp[0]) ? 16'b0000000011111111 : node8581;
														assign node8581 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node8585 = (inp[10]) ? node8603 : node8586;
												assign node8586 = (inp[14]) ? node8598 : node8587;
													assign node8587 = (inp[2]) ? node8595 : node8588;
														assign node8588 = (inp[3]) ? 16'b0000000111111111 : node8589;
															assign node8589 = (inp[5]) ? node8591 : 16'b0000001111111111;
																assign node8591 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node8595 = (inp[3]) ? 16'b0000000111111111 : 16'b0000000011111111;
													assign node8598 = (inp[0]) ? 16'b0000000001111111 : node8599;
														assign node8599 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node8603 = (inp[0]) ? node8609 : node8604;
													assign node8604 = (inp[14]) ? node8606 : 16'b0000001111111111;
														assign node8606 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node8609 = (inp[2]) ? node8611 : 16'b0000000001111111;
														assign node8611 = (inp[5]) ? node8613 : 16'b0000000000111111;
															assign node8613 = (inp[3]) ? node8615 : 16'b0000000000111111;
																assign node8615 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node8618 = (inp[14]) ? node8644 : node8619;
											assign node8619 = (inp[2]) ? node8635 : node8620;
												assign node8620 = (inp[10]) ? node8630 : node8621;
													assign node8621 = (inp[3]) ? node8623 : 16'b0000000111111111;
														assign node8623 = (inp[5]) ? node8625 : 16'b0000000111111111;
															assign node8625 = (inp[8]) ? 16'b0000000011111111 : node8626;
																assign node8626 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node8630 = (inp[3]) ? 16'b0000000001111111 : node8631;
														assign node8631 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node8635 = (inp[8]) ? node8637 : 16'b0000000011111111;
													assign node8637 = (inp[3]) ? node8639 : 16'b0000000011111111;
														assign node8639 = (inp[5]) ? node8641 : 16'b0000000001111111;
															assign node8641 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node8644 = (inp[3]) ? node8652 : node8645;
												assign node8645 = (inp[2]) ? node8647 : 16'b0000000011111111;
													assign node8647 = (inp[8]) ? 16'b0000000001111111 : node8648;
														assign node8648 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node8652 = (inp[5]) ? node8658 : node8653;
													assign node8653 = (inp[10]) ? 16'b0000000001111111 : node8654;
														assign node8654 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node8658 = (inp[2]) ? node8664 : node8659;
														assign node8659 = (inp[0]) ? node8661 : 16'b0000000000111111;
															assign node8661 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node8664 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node8667 = (inp[8]) ? node8709 : node8668;
										assign node8668 = (inp[3]) ? node8692 : node8669;
											assign node8669 = (inp[14]) ? node8677 : node8670;
												assign node8670 = (inp[10]) ? node8674 : node8671;
													assign node8671 = (inp[5]) ? 16'b0000001111111111 : 16'b0000000111111111;
													assign node8674 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node8677 = (inp[9]) ? node8689 : node8678;
													assign node8678 = (inp[5]) ? node8684 : node8679;
														assign node8679 = (inp[2]) ? node8681 : 16'b0000000111111111;
															assign node8681 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node8684 = (inp[0]) ? node8686 : 16'b0000000011111111;
															assign node8686 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node8689 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node8692 = (inp[5]) ? node8702 : node8693;
												assign node8693 = (inp[9]) ? 16'b0000000001111111 : node8694;
													assign node8694 = (inp[0]) ? node8696 : 16'b0000000111111111;
														assign node8696 = (inp[2]) ? 16'b0000000001111111 : node8697;
															assign node8697 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node8702 = (inp[10]) ? 16'b0000000000111111 : node8703;
													assign node8703 = (inp[2]) ? 16'b0000000000111111 : node8704;
														assign node8704 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node8709 = (inp[14]) ? node8737 : node8710;
											assign node8710 = (inp[3]) ? node8728 : node8711;
												assign node8711 = (inp[10]) ? node8721 : node8712;
													assign node8712 = (inp[2]) ? node8716 : node8713;
														assign node8713 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node8716 = (inp[0]) ? node8718 : 16'b0000000011111111;
															assign node8718 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node8721 = (inp[9]) ? node8725 : node8722;
														assign node8722 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node8725 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000000111111;
												assign node8728 = (inp[5]) ? node8732 : node8729;
													assign node8729 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node8732 = (inp[10]) ? 16'b0000000000111111 : node8733;
														assign node8733 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000011111111;
											assign node8737 = (inp[2]) ? node8759 : node8738;
												assign node8738 = (inp[10]) ? node8748 : node8739;
													assign node8739 = (inp[9]) ? node8745 : node8740;
														assign node8740 = (inp[5]) ? node8742 : 16'b0000000011111111;
															assign node8742 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000011111111;
														assign node8745 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node8748 = (inp[9]) ? node8752 : node8749;
														assign node8749 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node8752 = (inp[5]) ? 16'b0000000000011111 : node8753;
															assign node8753 = (inp[0]) ? node8755 : 16'b0000000000111111;
																assign node8755 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node8759 = (inp[9]) ? node8771 : node8760;
													assign node8760 = (inp[10]) ? node8764 : node8761;
														assign node8761 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node8764 = (inp[5]) ? node8766 : 16'b0000000000111111;
															assign node8766 = (inp[3]) ? node8768 : 16'b0000000000011111;
																assign node8768 = (inp[0]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node8771 = (inp[10]) ? node8773 : 16'b0000000000011111;
														assign node8773 = (inp[5]) ? node8775 : 16'b0000000000011111;
															assign node8775 = (inp[3]) ? 16'b0000000000000111 : 16'b0000000000001111;
								assign node8778 = (inp[10]) ? node8874 : node8779;
									assign node8779 = (inp[2]) ? node8819 : node8780;
										assign node8780 = (inp[1]) ? node8800 : node8781;
											assign node8781 = (inp[8]) ? node8789 : node8782;
												assign node8782 = (inp[0]) ? node8784 : 16'b0000000111111111;
													assign node8784 = (inp[3]) ? 16'b0000000001111111 : node8785;
														assign node8785 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node8789 = (inp[3]) ? node8795 : node8790;
													assign node8790 = (inp[14]) ? 16'b0000000011111111 : node8791;
														assign node8791 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node8795 = (inp[0]) ? 16'b0000000000111111 : node8796;
														assign node8796 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node8800 = (inp[8]) ? node8810 : node8801;
												assign node8801 = (inp[0]) ? node8803 : 16'b0000000011111111;
													assign node8803 = (inp[5]) ? node8805 : 16'b0000000011111111;
														assign node8805 = (inp[9]) ? node8807 : 16'b0000000001111111;
															assign node8807 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node8810 = (inp[5]) ? node8814 : node8811;
													assign node8811 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000011111111;
													assign node8814 = (inp[14]) ? 16'b0000000000111111 : node8815;
														assign node8815 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node8819 = (inp[14]) ? node8841 : node8820;
											assign node8820 = (inp[0]) ? node8832 : node8821;
												assign node8821 = (inp[3]) ? node8827 : node8822;
													assign node8822 = (inp[5]) ? 16'b0000000011111111 : node8823;
														assign node8823 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node8827 = (inp[5]) ? node8829 : 16'b0000000001111111;
														assign node8829 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000011111111;
												assign node8832 = (inp[9]) ? node8834 : 16'b0000000001111111;
													assign node8834 = (inp[5]) ? 16'b0000000000111111 : node8835;
														assign node8835 = (inp[8]) ? node8837 : 16'b0000000011111111;
															assign node8837 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node8841 = (inp[8]) ? node8849 : node8842;
												assign node8842 = (inp[1]) ? 16'b0000000000111111 : node8843;
													assign node8843 = (inp[3]) ? 16'b0000000000111111 : node8844;
														assign node8844 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000011111111;
												assign node8849 = (inp[5]) ? node8859 : node8850;
													assign node8850 = (inp[1]) ? node8852 : 16'b0000000001111111;
														assign node8852 = (inp[3]) ? node8856 : node8853;
															assign node8853 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000000111111;
															assign node8856 = (inp[0]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node8859 = (inp[0]) ? node8861 : 16'b0000000000011111;
														assign node8861 = (inp[9]) ? node8869 : node8862;
															assign node8862 = (inp[3]) ? node8866 : node8863;
																assign node8863 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000111111;
																assign node8866 = (inp[1]) ? 16'b0000000000001111 : 16'b0000000000011111;
															assign node8869 = (inp[3]) ? node8871 : 16'b0000000000001111;
																assign node8871 = (inp[1]) ? 16'b0000000000000111 : 16'b0000000000001111;
									assign node8874 = (inp[5]) ? node8908 : node8875;
										assign node8875 = (inp[0]) ? node8895 : node8876;
											assign node8876 = (inp[9]) ? node8880 : node8877;
												assign node8877 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node8880 = (inp[3]) ? node8890 : node8881;
													assign node8881 = (inp[8]) ? node8883 : 16'b0000000001111111;
														assign node8883 = (inp[2]) ? node8885 : 16'b0000000001111111;
															assign node8885 = (inp[1]) ? node8887 : 16'b0000000000111111;
																assign node8887 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node8890 = (inp[14]) ? 16'b0000000000111111 : node8891;
														assign node8891 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node8895 = (inp[1]) ? node8901 : node8896;
												assign node8896 = (inp[14]) ? 16'b0000000000111111 : node8897;
													assign node8897 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node8901 = (inp[3]) ? node8903 : 16'b0000000001111111;
													assign node8903 = (inp[9]) ? node8905 : 16'b0000000000011111;
														assign node8905 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000001111;
										assign node8908 = (inp[9]) ? node8924 : node8909;
											assign node8909 = (inp[14]) ? node8921 : node8910;
												assign node8910 = (inp[3]) ? node8918 : node8911;
													assign node8911 = (inp[2]) ? node8915 : node8912;
														assign node8912 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000111111111;
														assign node8915 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node8918 = (inp[1]) ? 16'b0000000000001111 : 16'b0000000000111111;
												assign node8921 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node8924 = (inp[8]) ? node8934 : node8925;
												assign node8925 = (inp[14]) ? node8931 : node8926;
													assign node8926 = (inp[2]) ? node8928 : 16'b0000000000111111;
														assign node8928 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node8931 = (inp[3]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node8934 = (inp[3]) ? node8940 : node8935;
													assign node8935 = (inp[2]) ? node8937 : 16'b0000000001111111;
														assign node8937 = (inp[0]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node8940 = (inp[2]) ? node8948 : node8941;
														assign node8941 = (inp[14]) ? node8943 : 16'b0000000000011111;
															assign node8943 = (inp[0]) ? 16'b0000000000001111 : node8944;
																assign node8944 = (inp[1]) ? 16'b0000000000001111 : 16'b0000000000011111;
														assign node8948 = (inp[0]) ? 16'b0000000000000111 : 16'b0000000000001111;
				assign node8951 = (inp[3]) ? node10389 : node8952;
					assign node8952 = (inp[4]) ? node9694 : node8953;
						assign node8953 = (inp[6]) ? node9339 : node8954;
							assign node8954 = (inp[12]) ? node9150 : node8955;
								assign node8955 = (inp[5]) ? node9047 : node8956;
									assign node8956 = (inp[10]) ? node9004 : node8957;
										assign node8957 = (inp[8]) ? node8987 : node8958;
											assign node8958 = (inp[0]) ? node8974 : node8959;
												assign node8959 = (inp[2]) ? node8965 : node8960;
													assign node8960 = (inp[9]) ? 16'b0000111111111111 : node8961;
														assign node8961 = (inp[13]) ? 16'b0000111111111111 : 16'b0001111111111111;
													assign node8965 = (inp[14]) ? node8971 : node8966;
														assign node8966 = (inp[13]) ? node8968 : 16'b0000111111111111;
															assign node8968 = (inp[9]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node8971 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node8974 = (inp[1]) ? node8984 : node8975;
													assign node8975 = (inp[13]) ? node8979 : node8976;
														assign node8976 = (inp[9]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node8979 = (inp[9]) ? node8981 : 16'b0000011111111111;
															assign node8981 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node8984 = (inp[14]) ? 16'b0000011111111111 : 16'b0000001111111111;
											assign node8987 = (inp[2]) ? node8997 : node8988;
												assign node8988 = (inp[14]) ? node8990 : 16'b0000011111111111;
													assign node8990 = (inp[1]) ? 16'b0000001111111111 : node8991;
														assign node8991 = (inp[9]) ? node8993 : 16'b0000011111111111;
															assign node8993 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node8997 = (inp[14]) ? node8999 : 16'b0000001111111111;
													assign node8999 = (inp[0]) ? node9001 : 16'b0000000111111111;
														assign node9001 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node9004 = (inp[0]) ? node9026 : node9005;
											assign node9005 = (inp[13]) ? node9015 : node9006;
												assign node9006 = (inp[14]) ? node9010 : node9007;
													assign node9007 = (inp[9]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node9010 = (inp[9]) ? node9012 : 16'b0000011111111111;
														assign node9012 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node9015 = (inp[2]) ? node9019 : node9016;
													assign node9016 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node9019 = (inp[1]) ? node9021 : 16'b0000001111111111;
														assign node9021 = (inp[9]) ? node9023 : 16'b0000000111111111;
															assign node9023 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node9026 = (inp[1]) ? node9038 : node9027;
												assign node9027 = (inp[13]) ? node9033 : node9028;
													assign node9028 = (inp[2]) ? node9030 : 16'b0000001111111111;
														assign node9030 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node9033 = (inp[2]) ? 16'b0000000011111111 : node9034;
														assign node9034 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node9038 = (inp[8]) ? node9040 : 16'b0000000111111111;
													assign node9040 = (inp[2]) ? 16'b0000000011111111 : node9041;
														assign node9041 = (inp[14]) ? node9043 : 16'b0000000111111111;
															assign node9043 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node9047 = (inp[8]) ? node9103 : node9048;
										assign node9048 = (inp[13]) ? node9080 : node9049;
											assign node9049 = (inp[2]) ? node9065 : node9050;
												assign node9050 = (inp[1]) ? node9056 : node9051;
													assign node9051 = (inp[10]) ? node9053 : 16'b0000111111111111;
														assign node9053 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node9056 = (inp[14]) ? 16'b0000000111111111 : node9057;
														assign node9057 = (inp[0]) ? 16'b0000001111111111 : node9058;
															assign node9058 = (inp[9]) ? node9060 : 16'b0000011111111111;
																assign node9060 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node9065 = (inp[1]) ? node9071 : node9066;
													assign node9066 = (inp[10]) ? 16'b0000000111111111 : node9067;
														assign node9067 = (inp[0]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node9071 = (inp[0]) ? 16'b0000000111111111 : node9072;
														assign node9072 = (inp[14]) ? node9074 : 16'b0000001111111111;
															assign node9074 = (inp[10]) ? 16'b0000000111111111 : node9075;
																assign node9075 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node9080 = (inp[0]) ? node9090 : node9081;
												assign node9081 = (inp[1]) ? node9083 : 16'b0000011111111111;
													assign node9083 = (inp[10]) ? 16'b0000000111111111 : node9084;
														assign node9084 = (inp[14]) ? node9086 : 16'b0000001111111111;
															assign node9086 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node9090 = (inp[14]) ? node9098 : node9091;
													assign node9091 = (inp[2]) ? node9095 : node9092;
														assign node9092 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node9095 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node9098 = (inp[9]) ? node9100 : 16'b0000000011111111;
														assign node9100 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node9103 = (inp[13]) ? node9125 : node9104;
											assign node9104 = (inp[10]) ? node9112 : node9105;
												assign node9105 = (inp[9]) ? 16'b0000000111111111 : node9106;
													assign node9106 = (inp[1]) ? 16'b0000000111111111 : node9107;
														assign node9107 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node9112 = (inp[2]) ? node9114 : 16'b0000000111111111;
													assign node9114 = (inp[0]) ? node9122 : node9115;
														assign node9115 = (inp[1]) ? 16'b0000000011111111 : node9116;
															assign node9116 = (inp[14]) ? node9118 : 16'b0000000111111111;
																assign node9118 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node9122 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node9125 = (inp[2]) ? node9143 : node9126;
												assign node9126 = (inp[0]) ? node9134 : node9127;
													assign node9127 = (inp[10]) ? node9131 : node9128;
														assign node9128 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node9131 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node9134 = (inp[14]) ? 16'b0000000011111111 : node9135;
														assign node9135 = (inp[1]) ? 16'b0000000011111111 : node9136;
															assign node9136 = (inp[10]) ? node9138 : 16'b0000000111111111;
																assign node9138 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node9143 = (inp[1]) ? 16'b0000000001111111 : node9144;
													assign node9144 = (inp[9]) ? 16'b0000000011111111 : node9145;
														assign node9145 = (inp[0]) ? 16'b0000000011111111 : 16'b0000001111111111;
								assign node9150 = (inp[5]) ? node9246 : node9151;
									assign node9151 = (inp[10]) ? node9193 : node9152;
										assign node9152 = (inp[9]) ? node9174 : node9153;
											assign node9153 = (inp[8]) ? node9167 : node9154;
												assign node9154 = (inp[0]) ? 16'b0000001111111111 : node9155;
													assign node9155 = (inp[13]) ? node9163 : node9156;
														assign node9156 = (inp[14]) ? node9158 : 16'b0000111111111111;
															assign node9158 = (inp[2]) ? 16'b0000011111111111 : node9159;
																assign node9159 = (inp[1]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node9163 = (inp[14]) ? 16'b0000000111111111 : 16'b0000011111111111;
												assign node9167 = (inp[1]) ? node9171 : node9168;
													assign node9168 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node9171 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node9174 = (inp[13]) ? node9184 : node9175;
												assign node9175 = (inp[1]) ? node9181 : node9176;
													assign node9176 = (inp[2]) ? node9178 : 16'b0000001111111111;
														assign node9178 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node9181 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node9184 = (inp[14]) ? node9190 : node9185;
													assign node9185 = (inp[0]) ? node9187 : 16'b0000000111111111;
														assign node9187 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node9190 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node9193 = (inp[8]) ? node9229 : node9194;
											assign node9194 = (inp[0]) ? node9212 : node9195;
												assign node9195 = (inp[14]) ? node9201 : node9196;
													assign node9196 = (inp[2]) ? 16'b0000001111111111 : node9197;
														assign node9197 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node9201 = (inp[9]) ? node9207 : node9202;
														assign node9202 = (inp[2]) ? 16'b0000000111111111 : node9203;
															assign node9203 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node9207 = (inp[2]) ? 16'b0000000001111111 : node9208;
															assign node9208 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node9212 = (inp[13]) ? node9220 : node9213;
													assign node9213 = (inp[14]) ? node9217 : node9214;
														assign node9214 = (inp[1]) ? 16'b0000001111111111 : 16'b0000000111111111;
														assign node9217 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node9220 = (inp[14]) ? 16'b0000000011111111 : node9221;
														assign node9221 = (inp[2]) ? node9223 : 16'b0000000111111111;
															assign node9223 = (inp[1]) ? 16'b0000000011111111 : node9224;
																assign node9224 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node9229 = (inp[0]) ? node9239 : node9230;
												assign node9230 = (inp[13]) ? node9234 : node9231;
													assign node9231 = (inp[1]) ? 16'b0000000011111111 : 16'b0000001111111111;
													assign node9234 = (inp[9]) ? node9236 : 16'b0000000011111111;
														assign node9236 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node9239 = (inp[13]) ? 16'b0000000001111111 : node9240;
													assign node9240 = (inp[9]) ? 16'b0000000011111111 : node9241;
														assign node9241 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node9246 = (inp[0]) ? node9298 : node9247;
										assign node9247 = (inp[9]) ? node9279 : node9248;
											assign node9248 = (inp[8]) ? node9262 : node9249;
												assign node9249 = (inp[2]) ? node9255 : node9250;
													assign node9250 = (inp[14]) ? node9252 : 16'b0000001111111111;
														assign node9252 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node9255 = (inp[14]) ? node9259 : node9256;
														assign node9256 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node9259 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node9262 = (inp[13]) ? node9272 : node9263;
													assign node9263 = (inp[14]) ? node9265 : 16'b0000000111111111;
														assign node9265 = (inp[1]) ? 16'b0000000011111111 : node9266;
															assign node9266 = (inp[10]) ? node9268 : 16'b0000000111111111;
																assign node9268 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node9272 = (inp[1]) ? node9276 : node9273;
														assign node9273 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node9276 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node9279 = (inp[2]) ? node9285 : node9280;
												assign node9280 = (inp[13]) ? 16'b0000000011111111 : node9281;
													assign node9281 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node9285 = (inp[8]) ? node9295 : node9286;
													assign node9286 = (inp[13]) ? node9292 : node9287;
														assign node9287 = (inp[14]) ? 16'b0000000011111111 : node9288;
															assign node9288 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node9292 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node9295 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node9298 = (inp[14]) ? node9324 : node9299;
											assign node9299 = (inp[9]) ? node9309 : node9300;
												assign node9300 = (inp[10]) ? node9304 : node9301;
													assign node9301 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node9304 = (inp[13]) ? 16'b0000000011111111 : node9305;
														assign node9305 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node9309 = (inp[2]) ? node9317 : node9310;
													assign node9310 = (inp[13]) ? node9314 : node9311;
														assign node9311 = (inp[8]) ? 16'b0000000111111111 : 16'b0000000011111111;
														assign node9314 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node9317 = (inp[10]) ? node9321 : node9318;
														assign node9318 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node9321 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node9324 = (inp[10]) ? node9332 : node9325;
												assign node9325 = (inp[9]) ? 16'b0000000001111111 : node9326;
													assign node9326 = (inp[8]) ? 16'b0000000011111111 : node9327;
														assign node9327 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node9332 = (inp[1]) ? 16'b0000000000111111 : node9333;
													assign node9333 = (inp[13]) ? node9335 : 16'b0000000001111111;
														assign node9335 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
							assign node9339 = (inp[8]) ? node9511 : node9340;
								assign node9340 = (inp[13]) ? node9426 : node9341;
									assign node9341 = (inp[12]) ? node9381 : node9342;
										assign node9342 = (inp[14]) ? node9362 : node9343;
											assign node9343 = (inp[5]) ? node9353 : node9344;
												assign node9344 = (inp[1]) ? node9348 : node9345;
													assign node9345 = (inp[10]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node9348 = (inp[9]) ? node9350 : 16'b0000001111111111;
														assign node9350 = (inp[0]) ? 16'b0000001111111111 : 16'b0000000111111111;
												assign node9353 = (inp[10]) ? node9355 : 16'b0000001111111111;
													assign node9355 = (inp[9]) ? node9359 : node9356;
														assign node9356 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node9359 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node9362 = (inp[2]) ? node9372 : node9363;
												assign node9363 = (inp[1]) ? node9369 : node9364;
													assign node9364 = (inp[9]) ? node9366 : 16'b0000111111111111;
														assign node9366 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node9369 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node9372 = (inp[10]) ? 16'b0000000011111111 : node9373;
													assign node9373 = (inp[9]) ? 16'b0000000011111111 : node9374;
														assign node9374 = (inp[1]) ? node9376 : 16'b0000000111111111;
															assign node9376 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node9381 = (inp[9]) ? node9405 : node9382;
											assign node9382 = (inp[1]) ? node9398 : node9383;
												assign node9383 = (inp[10]) ? node9387 : node9384;
													assign node9384 = (inp[0]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node9387 = (inp[5]) ? node9395 : node9388;
														assign node9388 = (inp[0]) ? node9390 : 16'b0000001111111111;
															assign node9390 = (inp[14]) ? 16'b0000000111111111 : node9391;
																assign node9391 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node9395 = (inp[14]) ? 16'b0000000111111111 : 16'b0000000011111111;
												assign node9398 = (inp[10]) ? node9400 : 16'b0000000111111111;
													assign node9400 = (inp[0]) ? node9402 : 16'b0000000111111111;
														assign node9402 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node9405 = (inp[5]) ? node9417 : node9406;
												assign node9406 = (inp[2]) ? node9412 : node9407;
													assign node9407 = (inp[1]) ? node9409 : 16'b0000000111111111;
														assign node9409 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node9412 = (inp[10]) ? 16'b0000000011111111 : node9413;
														assign node9413 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node9417 = (inp[1]) ? node9423 : node9418;
													assign node9418 = (inp[2]) ? 16'b0000000011111111 : node9419;
														assign node9419 = (inp[0]) ? 16'b0000000011111111 : 16'b0000001111111111;
													assign node9423 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node9426 = (inp[2]) ? node9482 : node9427;
										assign node9427 = (inp[9]) ? node9459 : node9428;
											assign node9428 = (inp[14]) ? node9448 : node9429;
												assign node9429 = (inp[5]) ? node9437 : node9430;
													assign node9430 = (inp[1]) ? node9432 : 16'b0000000111111111;
														assign node9432 = (inp[0]) ? 16'b0000001111111111 : node9433;
															assign node9433 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node9437 = (inp[1]) ? node9443 : node9438;
														assign node9438 = (inp[12]) ? node9440 : 16'b0000001111111111;
															assign node9440 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node9443 = (inp[10]) ? node9445 : 16'b0000000111111111;
															assign node9445 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node9448 = (inp[1]) ? node9456 : node9449;
													assign node9449 = (inp[12]) ? node9453 : node9450;
														assign node9450 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node9453 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node9456 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node9459 = (inp[12]) ? node9473 : node9460;
												assign node9460 = (inp[1]) ? node9466 : node9461;
													assign node9461 = (inp[0]) ? 16'b0000000001111111 : node9462;
														assign node9462 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node9466 = (inp[14]) ? node9468 : 16'b0000000011111111;
														assign node9468 = (inp[10]) ? node9470 : 16'b0000000011111111;
															assign node9470 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node9473 = (inp[10]) ? node9477 : node9474;
													assign node9474 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node9477 = (inp[14]) ? node9479 : 16'b0000000001111111;
														assign node9479 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node9482 = (inp[14]) ? node9498 : node9483;
											assign node9483 = (inp[5]) ? node9489 : node9484;
												assign node9484 = (inp[12]) ? 16'b0000000011111111 : node9485;
													assign node9485 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node9489 = (inp[0]) ? node9493 : node9490;
													assign node9490 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node9493 = (inp[1]) ? 16'b0000000000111111 : node9494;
														assign node9494 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node9498 = (inp[12]) ? node9504 : node9499;
												assign node9499 = (inp[1]) ? node9501 : 16'b0000000011111111;
													assign node9501 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node9504 = (inp[0]) ? node9506 : 16'b0000000001111111;
													assign node9506 = (inp[10]) ? node9508 : 16'b0000000001111111;
														assign node9508 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
								assign node9511 = (inp[1]) ? node9599 : node9512;
									assign node9512 = (inp[9]) ? node9554 : node9513;
										assign node9513 = (inp[12]) ? node9537 : node9514;
											assign node9514 = (inp[5]) ? node9522 : node9515;
												assign node9515 = (inp[14]) ? 16'b0000001111111111 : node9516;
													assign node9516 = (inp[13]) ? 16'b0000001111111111 : node9517;
														assign node9517 = (inp[10]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node9522 = (inp[2]) ? node9532 : node9523;
													assign node9523 = (inp[14]) ? 16'b0000000111111111 : node9524;
														assign node9524 = (inp[13]) ? 16'b0000000111111111 : node9525;
															assign node9525 = (inp[10]) ? node9527 : 16'b0000001111111111;
																assign node9527 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node9532 = (inp[0]) ? node9534 : 16'b0000000111111111;
														assign node9534 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node9537 = (inp[10]) ? node9549 : node9538;
												assign node9538 = (inp[0]) ? node9540 : 16'b0000000111111111;
													assign node9540 = (inp[5]) ? node9544 : node9541;
														assign node9541 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node9544 = (inp[13]) ? node9546 : 16'b0000000011111111;
															assign node9546 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node9549 = (inp[5]) ? 16'b0000000001111111 : node9550;
													assign node9550 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000111111111;
										assign node9554 = (inp[2]) ? node9578 : node9555;
											assign node9555 = (inp[0]) ? node9565 : node9556;
												assign node9556 = (inp[10]) ? node9560 : node9557;
													assign node9557 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node9560 = (inp[5]) ? 16'b0000000001111111 : node9561;
														assign node9561 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node9565 = (inp[13]) ? node9573 : node9566;
													assign node9566 = (inp[14]) ? node9570 : node9567;
														assign node9567 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node9570 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node9573 = (inp[10]) ? node9575 : 16'b0000000001111111;
														assign node9575 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node9578 = (inp[12]) ? node9590 : node9579;
												assign node9579 = (inp[5]) ? node9585 : node9580;
													assign node9580 = (inp[10]) ? 16'b0000000011111111 : node9581;
														assign node9581 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node9585 = (inp[10]) ? node9587 : 16'b0000000001111111;
														assign node9587 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000001111111;
												assign node9590 = (inp[0]) ? node9594 : node9591;
													assign node9591 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000011111111;
													assign node9594 = (inp[5]) ? node9596 : 16'b0000000000111111;
														assign node9596 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node9599 = (inp[0]) ? node9645 : node9600;
										assign node9600 = (inp[5]) ? node9626 : node9601;
											assign node9601 = (inp[12]) ? node9613 : node9602;
												assign node9602 = (inp[9]) ? node9608 : node9603;
													assign node9603 = (inp[13]) ? 16'b0000000011111111 : node9604;
														assign node9604 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node9608 = (inp[10]) ? node9610 : 16'b0000000011111111;
														assign node9610 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node9613 = (inp[13]) ? node9623 : node9614;
													assign node9614 = (inp[10]) ? node9616 : 16'b0000000011111111;
														assign node9616 = (inp[2]) ? 16'b0000000001111111 : node9617;
															assign node9617 = (inp[9]) ? node9619 : 16'b0000000011111111;
																assign node9619 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node9623 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node9626 = (inp[2]) ? node9634 : node9627;
												assign node9627 = (inp[9]) ? node9629 : 16'b0000000011111111;
													assign node9629 = (inp[10]) ? 16'b0000000000111111 : node9630;
														assign node9630 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000111111111;
												assign node9634 = (inp[9]) ? node9640 : node9635;
													assign node9635 = (inp[10]) ? node9637 : 16'b0000000001111111;
														assign node9637 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node9640 = (inp[14]) ? 16'b0000000000011111 : node9641;
														assign node9641 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node9645 = (inp[9]) ? node9671 : node9646;
											assign node9646 = (inp[14]) ? node9656 : node9647;
												assign node9647 = (inp[12]) ? node9651 : node9648;
													assign node9648 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000001111111;
													assign node9651 = (inp[13]) ? 16'b0000000001111111 : node9652;
														assign node9652 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000111111111;
												assign node9656 = (inp[10]) ? node9664 : node9657;
													assign node9657 = (inp[12]) ? node9661 : node9658;
														assign node9658 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node9661 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node9664 = (inp[5]) ? node9666 : 16'b0000000000111111;
														assign node9666 = (inp[12]) ? 16'b0000000000011111 : node9667;
															assign node9667 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node9671 = (inp[5]) ? node9681 : node9672;
												assign node9672 = (inp[12]) ? node9674 : 16'b0000000001111111;
													assign node9674 = (inp[13]) ? node9678 : node9675;
														assign node9675 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node9678 = (inp[2]) ? 16'b0000000000001111 : 16'b0000000000111111;
												assign node9681 = (inp[12]) ? node9689 : node9682;
													assign node9682 = (inp[10]) ? node9686 : node9683;
														assign node9683 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000011111111;
														assign node9686 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node9689 = (inp[2]) ? node9691 : 16'b0000000000011111;
														assign node9691 = (inp[13]) ? 16'b0000000000001111 : 16'b0000000000011111;
						assign node9694 = (inp[10]) ? node10012 : node9695;
							assign node9695 = (inp[0]) ? node9853 : node9696;
								assign node9696 = (inp[6]) ? node9784 : node9697;
									assign node9697 = (inp[14]) ? node9749 : node9698;
										assign node9698 = (inp[8]) ? node9716 : node9699;
											assign node9699 = (inp[9]) ? node9705 : node9700;
												assign node9700 = (inp[2]) ? 16'b0000011111111111 : node9701;
													assign node9701 = (inp[12]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node9705 = (inp[13]) ? node9711 : node9706;
													assign node9706 = (inp[12]) ? 16'b0000001111111111 : node9707;
														assign node9707 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node9711 = (inp[12]) ? node9713 : 16'b0000001111111111;
														assign node9713 = (inp[5]) ? 16'b0000000011111111 : 16'b0000001111111111;
											assign node9716 = (inp[2]) ? node9734 : node9717;
												assign node9717 = (inp[1]) ? node9729 : node9718;
													assign node9718 = (inp[12]) ? node9726 : node9719;
														assign node9719 = (inp[13]) ? 16'b0000001111111111 : node9720;
															assign node9720 = (inp[9]) ? node9722 : 16'b0000011111111111;
																assign node9722 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node9726 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node9729 = (inp[5]) ? node9731 : 16'b0000000111111111;
														assign node9731 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node9734 = (inp[12]) ? node9736 : 16'b0000000011111111;
													assign node9736 = (inp[5]) ? 16'b0000000011111111 : node9737;
														assign node9737 = (inp[9]) ? node9743 : node9738;
															assign node9738 = (inp[1]) ? 16'b0000000111111111 : node9739;
																assign node9739 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
															assign node9743 = (inp[13]) ? 16'b0000000011111111 : node9744;
																assign node9744 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node9749 = (inp[12]) ? node9759 : node9750;
											assign node9750 = (inp[2]) ? 16'b0000000111111111 : node9751;
												assign node9751 = (inp[8]) ? 16'b0000000111111111 : node9752;
													assign node9752 = (inp[5]) ? node9754 : 16'b0000001111111111;
														assign node9754 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node9759 = (inp[9]) ? node9771 : node9760;
												assign node9760 = (inp[13]) ? node9762 : 16'b0000000111111111;
													assign node9762 = (inp[2]) ? node9768 : node9763;
														assign node9763 = (inp[1]) ? node9765 : 16'b0000000111111111;
															assign node9765 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node9768 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node9771 = (inp[8]) ? node9779 : node9772;
													assign node9772 = (inp[2]) ? node9774 : 16'b0000000111111111;
														assign node9774 = (inp[5]) ? node9776 : 16'b0000000011111111;
															assign node9776 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node9779 = (inp[13]) ? 16'b0000000000111111 : node9780;
														assign node9780 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node9784 = (inp[9]) ? node9822 : node9785;
										assign node9785 = (inp[8]) ? node9803 : node9786;
											assign node9786 = (inp[12]) ? node9792 : node9787;
												assign node9787 = (inp[2]) ? 16'b0000001111111111 : node9788;
													assign node9788 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node9792 = (inp[2]) ? node9800 : node9793;
													assign node9793 = (inp[14]) ? 16'b0000000111111111 : node9794;
														assign node9794 = (inp[13]) ? 16'b0000000111111111 : node9795;
															assign node9795 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node9800 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000001111111;
											assign node9803 = (inp[12]) ? node9819 : node9804;
												assign node9804 = (inp[2]) ? node9812 : node9805;
													assign node9805 = (inp[14]) ? node9807 : 16'b0000000111111111;
														assign node9807 = (inp[13]) ? 16'b0000000011111111 : node9808;
															assign node9808 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node9812 = (inp[1]) ? node9816 : node9813;
														assign node9813 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node9816 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node9819 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000011111111;
										assign node9822 = (inp[12]) ? node9838 : node9823;
											assign node9823 = (inp[1]) ? node9829 : node9824;
												assign node9824 = (inp[5]) ? 16'b0000000011111111 : node9825;
													assign node9825 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node9829 = (inp[13]) ? node9833 : node9830;
													assign node9830 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000111111111;
													assign node9833 = (inp[8]) ? 16'b0000000000011111 : node9834;
														assign node9834 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node9838 = (inp[2]) ? node9846 : node9839;
												assign node9839 = (inp[14]) ? node9843 : node9840;
													assign node9840 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node9843 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000000111111;
												assign node9846 = (inp[13]) ? node9850 : node9847;
													assign node9847 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000000111111;
													assign node9850 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
								assign node9853 = (inp[14]) ? node9929 : node9854;
									assign node9854 = (inp[12]) ? node9892 : node9855;
										assign node9855 = (inp[13]) ? node9877 : node9856;
											assign node9856 = (inp[8]) ? node9864 : node9857;
												assign node9857 = (inp[9]) ? node9859 : 16'b0000001111111111;
													assign node9859 = (inp[1]) ? 16'b0000000111111111 : node9860;
														assign node9860 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node9864 = (inp[6]) ? node9872 : node9865;
													assign node9865 = (inp[5]) ? node9869 : node9866;
														assign node9866 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node9869 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node9872 = (inp[9]) ? 16'b0000000001111111 : node9873;
														assign node9873 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node9877 = (inp[1]) ? node9885 : node9878;
												assign node9878 = (inp[5]) ? 16'b0000000011111111 : node9879;
													assign node9879 = (inp[9]) ? node9881 : 16'b0000000111111111;
														assign node9881 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node9885 = (inp[6]) ? node9887 : 16'b0000000011111111;
													assign node9887 = (inp[9]) ? 16'b0000000001111111 : node9888;
														assign node9888 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node9892 = (inp[13]) ? node9912 : node9893;
											assign node9893 = (inp[8]) ? node9905 : node9894;
												assign node9894 = (inp[9]) ? node9902 : node9895;
													assign node9895 = (inp[1]) ? node9899 : node9896;
														assign node9896 = (inp[6]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node9899 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node9902 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000001111111;
												assign node9905 = (inp[5]) ? node9907 : 16'b0000000011111111;
													assign node9907 = (inp[1]) ? 16'b0000000000111111 : node9908;
														assign node9908 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node9912 = (inp[9]) ? node9924 : node9913;
												assign node9913 = (inp[8]) ? node9919 : node9914;
													assign node9914 = (inp[2]) ? 16'b0000000001111111 : node9915;
														assign node9915 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node9919 = (inp[2]) ? node9921 : 16'b0000000001111111;
														assign node9921 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node9924 = (inp[8]) ? 16'b0000000000011111 : node9925;
													assign node9925 = (inp[6]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node9929 = (inp[6]) ? node9977 : node9930;
										assign node9930 = (inp[13]) ? node9950 : node9931;
											assign node9931 = (inp[8]) ? node9937 : node9932;
												assign node9932 = (inp[12]) ? node9934 : 16'b0000000111111111;
													assign node9934 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node9937 = (inp[1]) ? node9945 : node9938;
													assign node9938 = (inp[12]) ? node9942 : node9939;
														assign node9939 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node9942 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000001111111;
													assign node9945 = (inp[9]) ? 16'b0000000001111111 : node9946;
														assign node9946 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node9950 = (inp[5]) ? node9966 : node9951;
												assign node9951 = (inp[1]) ? node9959 : node9952;
													assign node9952 = (inp[12]) ? node9956 : node9953;
														assign node9953 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node9956 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node9959 = (inp[2]) ? node9963 : node9960;
														assign node9960 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node9963 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node9966 = (inp[9]) ? node9968 : 16'b0000000001111111;
													assign node9968 = (inp[8]) ? node9972 : node9969;
														assign node9969 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node9972 = (inp[12]) ? 16'b0000000000111111 : node9973;
															assign node9973 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node9977 = (inp[2]) ? node9991 : node9978;
											assign node9978 = (inp[1]) ? node9984 : node9979;
												assign node9979 = (inp[9]) ? 16'b0000000001111111 : node9980;
													assign node9980 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000111111111;
												assign node9984 = (inp[12]) ? node9988 : node9985;
													assign node9985 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node9988 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000000011111;
											assign node9991 = (inp[5]) ? node10001 : node9992;
												assign node9992 = (inp[13]) ? node9996 : node9993;
													assign node9993 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node9996 = (inp[12]) ? node9998 : 16'b0000000001111111;
														assign node9998 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node10001 = (inp[9]) ? node10007 : node10002;
													assign node10002 = (inp[13]) ? node10004 : 16'b0000000000111111;
														assign node10004 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node10007 = (inp[8]) ? 16'b0000000000011111 : node10008;
														assign node10008 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
							assign node10012 = (inp[14]) ? node10180 : node10013;
								assign node10013 = (inp[5]) ? node10091 : node10014;
									assign node10014 = (inp[12]) ? node10062 : node10015;
										assign node10015 = (inp[0]) ? node10043 : node10016;
											assign node10016 = (inp[13]) ? node10030 : node10017;
												assign node10017 = (inp[8]) ? node10023 : node10018;
													assign node10018 = (inp[1]) ? node10020 : 16'b0000001111111111;
														assign node10020 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node10023 = (inp[9]) ? node10027 : node10024;
														assign node10024 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node10027 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node10030 = (inp[8]) ? node10032 : 16'b0000000111111111;
													assign node10032 = (inp[2]) ? node10040 : node10033;
														assign node10033 = (inp[6]) ? 16'b0000000011111111 : node10034;
															assign node10034 = (inp[1]) ? node10036 : 16'b0000000111111111;
																assign node10036 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node10040 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node10043 = (inp[9]) ? node10055 : node10044;
												assign node10044 = (inp[1]) ? node10046 : 16'b0000000111111111;
													assign node10046 = (inp[13]) ? node10050 : node10047;
														assign node10047 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node10050 = (inp[8]) ? node10052 : 16'b0000000011111111;
															assign node10052 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node10055 = (inp[8]) ? node10059 : node10056;
													assign node10056 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node10059 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node10062 = (inp[6]) ? node10076 : node10063;
											assign node10063 = (inp[2]) ? node10069 : node10064;
												assign node10064 = (inp[13]) ? 16'b0000000111111111 : node10065;
													assign node10065 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node10069 = (inp[1]) ? 16'b0000000001111111 : node10070;
													assign node10070 = (inp[8]) ? node10072 : 16'b0000000011111111;
														assign node10072 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node10076 = (inp[8]) ? node10084 : node10077;
												assign node10077 = (inp[9]) ? 16'b0000000001111111 : node10078;
													assign node10078 = (inp[0]) ? 16'b0000000001111111 : node10079;
														assign node10079 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node10084 = (inp[2]) ? 16'b0000000000111111 : node10085;
													assign node10085 = (inp[13]) ? node10087 : 16'b0000000011111111;
														assign node10087 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node10091 = (inp[1]) ? node10139 : node10092;
										assign node10092 = (inp[0]) ? node10118 : node10093;
											assign node10093 = (inp[13]) ? node10101 : node10094;
												assign node10094 = (inp[9]) ? 16'b0000000011111111 : node10095;
													assign node10095 = (inp[2]) ? 16'b0000000111111111 : node10096;
														assign node10096 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node10101 = (inp[12]) ? node10109 : node10102;
													assign node10102 = (inp[2]) ? node10104 : 16'b0000000111111111;
														assign node10104 = (inp[8]) ? node10106 : 16'b0000000011111111;
															assign node10106 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node10109 = (inp[2]) ? node10113 : node10110;
														assign node10110 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node10113 = (inp[9]) ? 16'b0000000000111111 : node10114;
															assign node10114 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node10118 = (inp[2]) ? node10136 : node10119;
												assign node10119 = (inp[8]) ? node10125 : node10120;
													assign node10120 = (inp[13]) ? node10122 : 16'b0000000011111111;
														assign node10122 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000011111111;
													assign node10125 = (inp[12]) ? 16'b0000000000011111 : node10126;
														assign node10126 = (inp[6]) ? node10130 : node10127;
															assign node10127 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
															assign node10130 = (inp[13]) ? node10132 : 16'b0000000001111111;
																assign node10132 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node10136 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node10139 = (inp[9]) ? node10163 : node10140;
											assign node10140 = (inp[8]) ? node10150 : node10141;
												assign node10141 = (inp[0]) ? node10145 : node10142;
													assign node10142 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node10145 = (inp[12]) ? 16'b0000000001111111 : node10146;
														assign node10146 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node10150 = (inp[13]) ? node10156 : node10151;
													assign node10151 = (inp[2]) ? 16'b0000000000111111 : node10152;
														assign node10152 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node10156 = (inp[2]) ? node10158 : 16'b0000000000111111;
														assign node10158 = (inp[6]) ? node10160 : 16'b0000000000111111;
															assign node10160 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node10163 = (inp[0]) ? node10171 : node10164;
												assign node10164 = (inp[12]) ? node10166 : 16'b0000000001111111;
													assign node10166 = (inp[13]) ? 16'b0000000000011111 : node10167;
														assign node10167 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node10171 = (inp[12]) ? node10175 : node10172;
													assign node10172 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000000011111;
													assign node10175 = (inp[13]) ? node10177 : 16'b0000000000011111;
														assign node10177 = (inp[8]) ? 16'b0000000000001111 : 16'b0000000000011111;
								assign node10180 = (inp[6]) ? node10280 : node10181;
									assign node10181 = (inp[2]) ? node10227 : node10182;
										assign node10182 = (inp[8]) ? node10204 : node10183;
											assign node10183 = (inp[9]) ? node10195 : node10184;
												assign node10184 = (inp[0]) ? node10186 : 16'b0000000111111111;
													assign node10186 = (inp[5]) ? node10190 : node10187;
														assign node10187 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node10190 = (inp[13]) ? node10192 : 16'b0000000011111111;
															assign node10192 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node10195 = (inp[0]) ? node10199 : node10196;
													assign node10196 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node10199 = (inp[13]) ? 16'b0000000001111111 : node10200;
														assign node10200 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node10204 = (inp[1]) ? node10212 : node10205;
												assign node10205 = (inp[0]) ? node10207 : 16'b0000000011111111;
													assign node10207 = (inp[12]) ? 16'b0000000000111111 : node10208;
														assign node10208 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node10212 = (inp[9]) ? node10220 : node10213;
													assign node10213 = (inp[13]) ? node10217 : node10214;
														assign node10214 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node10217 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000000111111;
													assign node10220 = (inp[0]) ? node10224 : node10221;
														assign node10221 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node10224 = (inp[13]) ? 16'b0000000000001111 : 16'b0000000000011111;
										assign node10227 = (inp[5]) ? node10257 : node10228;
											assign node10228 = (inp[0]) ? node10238 : node10229;
												assign node10229 = (inp[9]) ? node10231 : 16'b0000000011111111;
													assign node10231 = (inp[12]) ? node10233 : 16'b0000000000111111;
														assign node10233 = (inp[13]) ? 16'b0000000001111111 : node10234;
															assign node10234 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node10238 = (inp[1]) ? node10248 : node10239;
													assign node10239 = (inp[12]) ? node10241 : 16'b0000000001111111;
														assign node10241 = (inp[8]) ? 16'b0000000000111111 : node10242;
															assign node10242 = (inp[9]) ? node10244 : 16'b0000000001111111;
																assign node10244 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node10248 = (inp[8]) ? node10252 : node10249;
														assign node10249 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node10252 = (inp[9]) ? node10254 : 16'b0000000000111111;
															assign node10254 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node10257 = (inp[13]) ? node10267 : node10258;
												assign node10258 = (inp[12]) ? node10260 : 16'b0000000011111111;
													assign node10260 = (inp[1]) ? node10264 : node10261;
														assign node10261 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node10264 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node10267 = (inp[9]) ? node10273 : node10268;
													assign node10268 = (inp[8]) ? node10270 : 16'b0000000000111111;
														assign node10270 = (inp[1]) ? 16'b0000000000001111 : 16'b0000000000111111;
													assign node10273 = (inp[12]) ? node10275 : 16'b0000000000011111;
														assign node10275 = (inp[8]) ? 16'b0000000000001111 : node10276;
															assign node10276 = (inp[0]) ? 16'b0000000000001111 : 16'b0000000000011111;
									assign node10280 = (inp[13]) ? node10330 : node10281;
										assign node10281 = (inp[12]) ? node10307 : node10282;
											assign node10282 = (inp[1]) ? node10298 : node10283;
												assign node10283 = (inp[2]) ? node10293 : node10284;
													assign node10284 = (inp[0]) ? node10288 : node10285;
														assign node10285 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node10288 = (inp[8]) ? 16'b0000000001111111 : node10289;
															assign node10289 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node10293 = (inp[0]) ? node10295 : 16'b0000000001111111;
														assign node10295 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node10298 = (inp[9]) ? 16'b0000000000111111 : node10299;
													assign node10299 = (inp[5]) ? node10303 : node10300;
														assign node10300 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node10303 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node10307 = (inp[5]) ? node10313 : node10308;
												assign node10308 = (inp[1]) ? node10310 : 16'b0000000001111111;
													assign node10310 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node10313 = (inp[0]) ? node10323 : node10314;
													assign node10314 = (inp[9]) ? node10318 : node10315;
														assign node10315 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node10318 = (inp[2]) ? node10320 : 16'b0000000000111111;
															assign node10320 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node10323 = (inp[2]) ? node10327 : node10324;
														assign node10324 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node10327 = (inp[8]) ? 16'b0000000000000111 : 16'b0000000000011111;
										assign node10330 = (inp[8]) ? node10356 : node10331;
											assign node10331 = (inp[0]) ? node10347 : node10332;
												assign node10332 = (inp[1]) ? node10342 : node10333;
													assign node10333 = (inp[9]) ? node10337 : node10334;
														assign node10334 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node10337 = (inp[5]) ? node10339 : 16'b0000000001111111;
															assign node10339 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node10342 = (inp[12]) ? node10344 : 16'b0000000000111111;
														assign node10344 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node10347 = (inp[2]) ? node10353 : node10348;
													assign node10348 = (inp[5]) ? node10350 : 16'b0000000000111111;
														assign node10350 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000001111111;
													assign node10353 = (inp[12]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node10356 = (inp[5]) ? node10372 : node10357;
												assign node10357 = (inp[1]) ? node10363 : node10358;
													assign node10358 = (inp[9]) ? node10360 : 16'b0000000000111111;
														assign node10360 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node10363 = (inp[0]) ? 16'b0000000000011111 : node10364;
														assign node10364 = (inp[2]) ? node10366 : 16'b0000000000111111;
															assign node10366 = (inp[12]) ? 16'b0000000000011111 : node10367;
																assign node10367 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node10372 = (inp[9]) ? node10380 : node10373;
													assign node10373 = (inp[12]) ? 16'b0000000000011111 : node10374;
														assign node10374 = (inp[1]) ? 16'b0000000000011111 : node10375;
															assign node10375 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node10380 = (inp[1]) ? node10386 : node10381;
														assign node10381 = (inp[12]) ? 16'b0000000000001111 : node10382;
															assign node10382 = (inp[0]) ? 16'b0000000000001111 : 16'b0000000000011111;
														assign node10386 = (inp[0]) ? 16'b0000000000001111 : 16'b0000000000000111;
					assign node10389 = (inp[2]) ? node11117 : node10390;
						assign node10390 = (inp[9]) ? node10744 : node10391;
							assign node10391 = (inp[13]) ? node10575 : node10392;
								assign node10392 = (inp[6]) ? node10498 : node10393;
									assign node10393 = (inp[5]) ? node10439 : node10394;
										assign node10394 = (inp[4]) ? node10416 : node10395;
											assign node10395 = (inp[1]) ? node10403 : node10396;
												assign node10396 = (inp[8]) ? node10398 : 16'b0000011111111111;
													assign node10398 = (inp[14]) ? 16'b0000001111111111 : node10399;
														assign node10399 = (inp[0]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node10403 = (inp[0]) ? node10411 : node10404;
													assign node10404 = (inp[14]) ? node10408 : node10405;
														assign node10405 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node10408 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node10411 = (inp[8]) ? 16'b0000000111111111 : node10412;
														assign node10412 = (inp[12]) ? 16'b0000000011111111 : 16'b0000001111111111;
											assign node10416 = (inp[1]) ? node10430 : node10417;
												assign node10417 = (inp[14]) ? 16'b0000000111111111 : node10418;
													assign node10418 = (inp[10]) ? node10422 : node10419;
														assign node10419 = (inp[12]) ? 16'b0000001111111111 : 16'b0000111111111111;
														assign node10422 = (inp[12]) ? 16'b0000000111111111 : node10423;
															assign node10423 = (inp[0]) ? node10425 : 16'b0000001111111111;
																assign node10425 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node10430 = (inp[12]) ? 16'b0000000011111111 : node10431;
													assign node10431 = (inp[0]) ? node10435 : node10432;
														assign node10432 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node10435 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node10439 = (inp[10]) ? node10465 : node10440;
											assign node10440 = (inp[12]) ? node10452 : node10441;
												assign node10441 = (inp[1]) ? node10447 : node10442;
													assign node10442 = (inp[4]) ? node10444 : 16'b0000011111111111;
														assign node10444 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node10447 = (inp[14]) ? 16'b0000000111111111 : node10448;
														assign node10448 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node10452 = (inp[4]) ? node10458 : node10453;
													assign node10453 = (inp[8]) ? node10455 : 16'b0000000111111111;
														assign node10455 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node10458 = (inp[14]) ? node10462 : node10459;
														assign node10459 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node10462 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node10465 = (inp[12]) ? node10483 : node10466;
												assign node10466 = (inp[8]) ? node10470 : node10467;
													assign node10467 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node10470 = (inp[14]) ? node10478 : node10471;
														assign node10471 = (inp[4]) ? node10473 : 16'b0000000111111111;
															assign node10473 = (inp[0]) ? 16'b0000000011111111 : node10474;
																assign node10474 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node10478 = (inp[1]) ? node10480 : 16'b0000000011111111;
															assign node10480 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node10483 = (inp[1]) ? node10489 : node10484;
													assign node10484 = (inp[0]) ? node10486 : 16'b0000000011111111;
														assign node10486 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node10489 = (inp[14]) ? node10493 : node10490;
														assign node10490 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node10493 = (inp[0]) ? node10495 : 16'b0000000001111111;
															assign node10495 = (inp[4]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node10498 = (inp[0]) ? node10540 : node10499;
										assign node10499 = (inp[5]) ? node10523 : node10500;
											assign node10500 = (inp[4]) ? node10506 : node10501;
												assign node10501 = (inp[8]) ? node10503 : 16'b0000001111111111;
													assign node10503 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node10506 = (inp[8]) ? node10512 : node10507;
													assign node10507 = (inp[10]) ? node10509 : 16'b0000011111111111;
														assign node10509 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node10512 = (inp[1]) ? node10516 : node10513;
														assign node10513 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node10516 = (inp[10]) ? node10518 : 16'b0000000011111111;
															assign node10518 = (inp[14]) ? node10520 : 16'b0000000001111111;
																assign node10520 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node10523 = (inp[1]) ? node10531 : node10524;
												assign node10524 = (inp[10]) ? 16'b0000000011111111 : node10525;
													assign node10525 = (inp[8]) ? node10527 : 16'b0000000111111111;
														assign node10527 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node10531 = (inp[12]) ? node10533 : 16'b0000000011111111;
													assign node10533 = (inp[4]) ? 16'b0000000001111111 : node10534;
														assign node10534 = (inp[8]) ? node10536 : 16'b0000000011111111;
															assign node10536 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node10540 = (inp[14]) ? node10562 : node10541;
											assign node10541 = (inp[8]) ? node10553 : node10542;
												assign node10542 = (inp[12]) ? node10546 : node10543;
													assign node10543 = (inp[10]) ? 16'b0000001111111111 : 16'b0000000111111111;
													assign node10546 = (inp[1]) ? node10550 : node10547;
														assign node10547 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node10550 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node10553 = (inp[12]) ? node10559 : node10554;
													assign node10554 = (inp[1]) ? node10556 : 16'b0000000011111111;
														assign node10556 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node10559 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000001111111;
											assign node10562 = (inp[8]) ? node10568 : node10563;
												assign node10563 = (inp[1]) ? node10565 : 16'b0000000001111111;
													assign node10565 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node10568 = (inp[4]) ? node10570 : 16'b0000000001111111;
													assign node10570 = (inp[10]) ? 16'b0000000000111111 : node10571;
														assign node10571 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
								assign node10575 = (inp[4]) ? node10653 : node10576;
									assign node10576 = (inp[10]) ? node10604 : node10577;
										assign node10577 = (inp[5]) ? node10589 : node10578;
											assign node10578 = (inp[8]) ? node10582 : node10579;
												assign node10579 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node10582 = (inp[0]) ? node10584 : 16'b0000000111111111;
													assign node10584 = (inp[1]) ? 16'b0000000011111111 : node10585;
														assign node10585 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node10589 = (inp[8]) ? node10599 : node10590;
												assign node10590 = (inp[6]) ? node10594 : node10591;
													assign node10591 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node10594 = (inp[0]) ? 16'b0000000001111111 : node10595;
														assign node10595 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node10599 = (inp[1]) ? node10601 : 16'b0000000011111111;
													assign node10601 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node10604 = (inp[1]) ? node10638 : node10605;
											assign node10605 = (inp[0]) ? node10623 : node10606;
												assign node10606 = (inp[5]) ? node10618 : node10607;
													assign node10607 = (inp[6]) ? node10613 : node10608;
														assign node10608 = (inp[8]) ? node10610 : 16'b0000001111111111;
															assign node10610 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node10613 = (inp[12]) ? node10615 : 16'b0000000111111111;
															assign node10615 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node10618 = (inp[12]) ? 16'b0000000011111111 : node10619;
														assign node10619 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node10623 = (inp[14]) ? node10631 : node10624;
													assign node10624 = (inp[5]) ? node10628 : node10625;
														assign node10625 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node10628 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node10631 = (inp[12]) ? node10635 : node10632;
														assign node10632 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node10635 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node10638 = (inp[8]) ? node10644 : node10639;
												assign node10639 = (inp[6]) ? node10641 : 16'b0000000111111111;
													assign node10641 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node10644 = (inp[5]) ? node10646 : 16'b0000000001111111;
													assign node10646 = (inp[6]) ? node10648 : 16'b0000000001111111;
														assign node10648 = (inp[14]) ? 16'b0000000000111111 : node10649;
															assign node10649 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node10653 = (inp[12]) ? node10689 : node10654;
										assign node10654 = (inp[10]) ? node10676 : node10655;
											assign node10655 = (inp[14]) ? node10663 : node10656;
												assign node10656 = (inp[1]) ? 16'b0000000011111111 : node10657;
													assign node10657 = (inp[0]) ? node10659 : 16'b0000001111111111;
														assign node10659 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node10663 = (inp[8]) ? 16'b0000000001111111 : node10664;
													assign node10664 = (inp[1]) ? node10670 : node10665;
														assign node10665 = (inp[5]) ? node10667 : 16'b0000000011111111;
															assign node10667 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node10670 = (inp[0]) ? 16'b0000000001111111 : node10671;
															assign node10671 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node10676 = (inp[6]) ? node10682 : node10677;
												assign node10677 = (inp[0]) ? node10679 : 16'b0000000011111111;
													assign node10679 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node10682 = (inp[1]) ? node10684 : 16'b0000000001111111;
													assign node10684 = (inp[0]) ? node10686 : 16'b0000000000111111;
														assign node10686 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node10689 = (inp[14]) ? node10717 : node10690;
											assign node10690 = (inp[1]) ? node10704 : node10691;
												assign node10691 = (inp[0]) ? node10697 : node10692;
													assign node10692 = (inp[10]) ? node10694 : 16'b0000000111111111;
														assign node10694 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node10697 = (inp[5]) ? node10701 : node10698;
														assign node10698 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node10701 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node10704 = (inp[0]) ? node10712 : node10705;
													assign node10705 = (inp[5]) ? 16'b0000000001111111 : node10706;
														assign node10706 = (inp[6]) ? node10708 : 16'b0000000001111111;
															assign node10708 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node10712 = (inp[10]) ? 16'b0000000000111111 : node10713;
														assign node10713 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node10717 = (inp[6]) ? node10727 : node10718;
												assign node10718 = (inp[1]) ? node10720 : 16'b0000000001111111;
													assign node10720 = (inp[10]) ? node10724 : node10721;
														assign node10721 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node10724 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node10727 = (inp[0]) ? node10737 : node10728;
													assign node10728 = (inp[5]) ? node10734 : node10729;
														assign node10729 = (inp[8]) ? 16'b0000000000111111 : node10730;
															assign node10730 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node10734 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node10737 = (inp[8]) ? node10739 : 16'b0000000000011111;
														assign node10739 = (inp[5]) ? node10741 : 16'b0000000000001111;
															assign node10741 = (inp[10]) ? 16'b0000000000000111 : 16'b0000000000001111;
							assign node10744 = (inp[5]) ? node10938 : node10745;
								assign node10745 = (inp[0]) ? node10835 : node10746;
									assign node10746 = (inp[12]) ? node10786 : node10747;
										assign node10747 = (inp[13]) ? node10767 : node10748;
											assign node10748 = (inp[4]) ? node10760 : node10749;
												assign node10749 = (inp[10]) ? node10757 : node10750;
													assign node10750 = (inp[8]) ? node10754 : node10751;
														assign node10751 = (inp[1]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node10754 = (inp[6]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node10757 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node10760 = (inp[1]) ? node10764 : node10761;
													assign node10761 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node10764 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node10767 = (inp[10]) ? node10779 : node10768;
												assign node10768 = (inp[8]) ? node10774 : node10769;
													assign node10769 = (inp[14]) ? node10771 : 16'b0000000111111111;
														assign node10771 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node10774 = (inp[4]) ? 16'b0000000011111111 : node10775;
														assign node10775 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node10779 = (inp[8]) ? node10781 : 16'b0000000011111111;
													assign node10781 = (inp[14]) ? node10783 : 16'b0000000001111111;
														assign node10783 = (inp[6]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node10786 = (inp[8]) ? node10818 : node10787;
											assign node10787 = (inp[1]) ? node10803 : node10788;
												assign node10788 = (inp[6]) ? node10794 : node10789;
													assign node10789 = (inp[4]) ? node10791 : 16'b0000000111111111;
														assign node10791 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node10794 = (inp[14]) ? node10800 : node10795;
														assign node10795 = (inp[4]) ? 16'b0000000011111111 : node10796;
															assign node10796 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node10800 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node10803 = (inp[4]) ? node10813 : node10804;
													assign node10804 = (inp[14]) ? node10810 : node10805;
														assign node10805 = (inp[6]) ? 16'b0000000011111111 : node10806;
															assign node10806 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node10810 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node10813 = (inp[13]) ? node10815 : 16'b0000000011111111;
														assign node10815 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node10818 = (inp[6]) ? node10826 : node10819;
												assign node10819 = (inp[13]) ? node10821 : 16'b0000000011111111;
													assign node10821 = (inp[10]) ? node10823 : 16'b0000000011111111;
														assign node10823 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node10826 = (inp[4]) ? node10832 : node10827;
													assign node10827 = (inp[10]) ? node10829 : 16'b0000000011111111;
														assign node10829 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node10832 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node10835 = (inp[14]) ? node10879 : node10836;
										assign node10836 = (inp[6]) ? node10858 : node10837;
											assign node10837 = (inp[8]) ? node10853 : node10838;
												assign node10838 = (inp[12]) ? node10842 : node10839;
													assign node10839 = (inp[10]) ? 16'b0000000111111111 : 16'b0000011111111111;
													assign node10842 = (inp[10]) ? node10848 : node10843;
														assign node10843 = (inp[13]) ? 16'b0000000011111111 : node10844;
															assign node10844 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node10848 = (inp[1]) ? node10850 : 16'b0000000011111111;
															assign node10850 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node10853 = (inp[12]) ? node10855 : 16'b0000000011111111;
													assign node10855 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000011111111;
											assign node10858 = (inp[10]) ? node10866 : node10859;
												assign node10859 = (inp[1]) ? node10863 : node10860;
													assign node10860 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node10863 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node10866 = (inp[13]) ? node10874 : node10867;
													assign node10867 = (inp[1]) ? node10871 : node10868;
														assign node10868 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000001111111;
														assign node10871 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node10874 = (inp[1]) ? node10876 : 16'b0000000000011111;
														assign node10876 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node10879 = (inp[12]) ? node10911 : node10880;
											assign node10880 = (inp[1]) ? node10896 : node10881;
												assign node10881 = (inp[4]) ? node10887 : node10882;
													assign node10882 = (inp[10]) ? node10884 : 16'b0000000111111111;
														assign node10884 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node10887 = (inp[8]) ? node10891 : node10888;
														assign node10888 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node10891 = (inp[10]) ? node10893 : 16'b0000000001111111;
															assign node10893 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node10896 = (inp[10]) ? node10902 : node10897;
													assign node10897 = (inp[13]) ? node10899 : 16'b0000000001111111;
														assign node10899 = (inp[4]) ? 16'b0000000000011111 : 16'b0000000001111111;
													assign node10902 = (inp[6]) ? node10904 : 16'b0000000000111111;
														assign node10904 = (inp[8]) ? 16'b0000000000011111 : node10905;
															assign node10905 = (inp[13]) ? node10907 : 16'b0000000000111111;
																assign node10907 = (inp[4]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node10911 = (inp[13]) ? node10925 : node10912;
												assign node10912 = (inp[6]) ? node10920 : node10913;
													assign node10913 = (inp[4]) ? 16'b0000000000111111 : node10914;
														assign node10914 = (inp[8]) ? node10916 : 16'b0000000001111111;
															assign node10916 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node10920 = (inp[4]) ? node10922 : 16'b0000000000111111;
														assign node10922 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node10925 = (inp[6]) ? node10933 : node10926;
													assign node10926 = (inp[8]) ? node10928 : 16'b0000000000111111;
														assign node10928 = (inp[4]) ? 16'b0000000000011111 : node10929;
															assign node10929 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node10933 = (inp[1]) ? node10935 : 16'b0000000000001111;
														assign node10935 = (inp[10]) ? 16'b0000000000000111 : 16'b0000000000001111;
								assign node10938 = (inp[12]) ? node11034 : node10939;
									assign node10939 = (inp[13]) ? node10983 : node10940;
										assign node10940 = (inp[10]) ? node10962 : node10941;
											assign node10941 = (inp[8]) ? node10953 : node10942;
												assign node10942 = (inp[1]) ? node10948 : node10943;
													assign node10943 = (inp[14]) ? 16'b0000000111111111 : node10944;
														assign node10944 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node10948 = (inp[0]) ? node10950 : 16'b0000001111111111;
														assign node10950 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node10953 = (inp[6]) ? 16'b0000000001111111 : node10954;
													assign node10954 = (inp[14]) ? node10958 : node10955;
														assign node10955 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node10958 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node10962 = (inp[1]) ? node10978 : node10963;
												assign node10963 = (inp[0]) ? node10973 : node10964;
													assign node10964 = (inp[4]) ? node10966 : 16'b0000000111111111;
														assign node10966 = (inp[6]) ? 16'b0000000001111111 : node10967;
															assign node10967 = (inp[8]) ? node10969 : 16'b0000000011111111;
																assign node10969 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node10973 = (inp[6]) ? 16'b0000000001111111 : node10974;
														assign node10974 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000011111111;
												assign node10978 = (inp[14]) ? node10980 : 16'b0000000000111111;
													assign node10980 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node10983 = (inp[4]) ? node11007 : node10984;
											assign node10984 = (inp[14]) ? node10998 : node10985;
												assign node10985 = (inp[8]) ? 16'b0000000001111111 : node10986;
													assign node10986 = (inp[1]) ? node10990 : node10987;
														assign node10987 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node10990 = (inp[0]) ? node10994 : node10991;
															assign node10991 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
															assign node10994 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node10998 = (inp[6]) ? 16'b0000000000111111 : node10999;
													assign node10999 = (inp[1]) ? node11001 : 16'b0000000001111111;
														assign node11001 = (inp[8]) ? node11003 : 16'b0000000001111111;
															assign node11003 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node11007 = (inp[10]) ? node11021 : node11008;
												assign node11008 = (inp[0]) ? node11014 : node11009;
													assign node11009 = (inp[6]) ? node11011 : 16'b0000000011111111;
														assign node11011 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node11014 = (inp[14]) ? node11016 : 16'b0000000001111111;
														assign node11016 = (inp[6]) ? node11018 : 16'b0000000000111111;
															assign node11018 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node11021 = (inp[6]) ? node11027 : node11022;
													assign node11022 = (inp[8]) ? node11024 : 16'b0000000001111111;
														assign node11024 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node11027 = (inp[0]) ? node11029 : 16'b0000000000011111;
														assign node11029 = (inp[8]) ? 16'b0000000000001111 : node11030;
															assign node11030 = (inp[14]) ? 16'b0000000000001111 : 16'b0000000000011111;
									assign node11034 = (inp[0]) ? node11074 : node11035;
										assign node11035 = (inp[8]) ? node11061 : node11036;
											assign node11036 = (inp[14]) ? node11046 : node11037;
												assign node11037 = (inp[4]) ? node11043 : node11038;
													assign node11038 = (inp[13]) ? node11040 : 16'b0000000011111111;
														assign node11040 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node11043 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node11046 = (inp[6]) ? node11052 : node11047;
													assign node11047 = (inp[13]) ? node11049 : 16'b0000000001111111;
														assign node11049 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node11052 = (inp[4]) ? node11058 : node11053;
														assign node11053 = (inp[1]) ? 16'b0000000000111111 : node11054;
															assign node11054 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node11058 = (inp[13]) ? 16'b0000000000001111 : 16'b0000000000111111;
											assign node11061 = (inp[14]) ? node11071 : node11062;
												assign node11062 = (inp[4]) ? node11066 : node11063;
													assign node11063 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000011111111;
													assign node11066 = (inp[13]) ? node11068 : 16'b0000000000111111;
														assign node11068 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node11071 = (inp[4]) ? 16'b0000000000000111 : 16'b0000000000011111;
										assign node11074 = (inp[1]) ? node11096 : node11075;
											assign node11075 = (inp[10]) ? node11089 : node11076;
												assign node11076 = (inp[4]) ? node11082 : node11077;
													assign node11077 = (inp[6]) ? node11079 : 16'b0000000011111111;
														assign node11079 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node11082 = (inp[13]) ? 16'b0000000000011111 : node11083;
														assign node11083 = (inp[14]) ? 16'b0000000000111111 : node11084;
															assign node11084 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node11089 = (inp[4]) ? node11093 : node11090;
													assign node11090 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node11093 = (inp[6]) ? 16'b0000000000011111 : 16'b0000000000001111;
											assign node11096 = (inp[13]) ? node11106 : node11097;
												assign node11097 = (inp[6]) ? node11101 : node11098;
													assign node11098 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node11101 = (inp[10]) ? node11103 : 16'b0000000000011111;
														assign node11103 = (inp[14]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node11106 = (inp[10]) ? node11112 : node11107;
													assign node11107 = (inp[14]) ? 16'b0000000000001111 : node11108;
														assign node11108 = (inp[6]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node11112 = (inp[14]) ? node11114 : 16'b0000000000001111;
														assign node11114 = (inp[6]) ? 16'b0000000000000111 : 16'b0000000000011111;
						assign node11117 = (inp[14]) ? node11503 : node11118;
							assign node11118 = (inp[13]) ? node11316 : node11119;
								assign node11119 = (inp[0]) ? node11215 : node11120;
									assign node11120 = (inp[12]) ? node11168 : node11121;
										assign node11121 = (inp[4]) ? node11141 : node11122;
											assign node11122 = (inp[5]) ? node11134 : node11123;
												assign node11123 = (inp[9]) ? node11129 : node11124;
													assign node11124 = (inp[10]) ? node11126 : 16'b0000001111111111;
														assign node11126 = (inp[6]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node11129 = (inp[1]) ? node11131 : 16'b0000000111111111;
														assign node11131 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node11134 = (inp[10]) ? node11136 : 16'b0000000111111111;
													assign node11136 = (inp[6]) ? 16'b0000000011111111 : node11137;
														assign node11137 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node11141 = (inp[9]) ? node11153 : node11142;
												assign node11142 = (inp[1]) ? 16'b0000000011111111 : node11143;
													assign node11143 = (inp[10]) ? node11145 : 16'b0000000111111111;
														assign node11145 = (inp[8]) ? node11147 : 16'b0000000111111111;
															assign node11147 = (inp[5]) ? 16'b0000000011111111 : node11148;
																assign node11148 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node11153 = (inp[8]) ? node11163 : node11154;
													assign node11154 = (inp[1]) ? node11158 : node11155;
														assign node11155 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node11158 = (inp[10]) ? node11160 : 16'b0000000011111111;
															assign node11160 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node11163 = (inp[1]) ? node11165 : 16'b0000000001111111;
														assign node11165 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node11168 = (inp[10]) ? node11196 : node11169;
											assign node11169 = (inp[6]) ? node11187 : node11170;
												assign node11170 = (inp[8]) ? node11180 : node11171;
													assign node11171 = (inp[5]) ? node11173 : 16'b0000011111111111;
														assign node11173 = (inp[1]) ? 16'b0000000111111111 : node11174;
															assign node11174 = (inp[9]) ? 16'b0000000111111111 : node11175;
																assign node11175 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node11180 = (inp[5]) ? node11182 : 16'b0000000111111111;
														assign node11182 = (inp[1]) ? node11184 : 16'b0000000011111111;
															assign node11184 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node11187 = (inp[4]) ? node11193 : node11188;
													assign node11188 = (inp[5]) ? node11190 : 16'b0000000011111111;
														assign node11190 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node11193 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node11196 = (inp[8]) ? node11206 : node11197;
												assign node11197 = (inp[5]) ? node11199 : 16'b0000000011111111;
													assign node11199 = (inp[6]) ? 16'b0000000000111111 : node11200;
														assign node11200 = (inp[9]) ? 16'b0000000001111111 : node11201;
															assign node11201 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node11206 = (inp[5]) ? node11208 : 16'b0000000001111111;
													assign node11208 = (inp[1]) ? 16'b0000000000011111 : node11209;
														assign node11209 = (inp[9]) ? node11211 : 16'b0000000001111111;
															assign node11211 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node11215 = (inp[4]) ? node11265 : node11216;
										assign node11216 = (inp[9]) ? node11240 : node11217;
											assign node11217 = (inp[8]) ? node11233 : node11218;
												assign node11218 = (inp[12]) ? node11224 : node11219;
													assign node11219 = (inp[1]) ? node11221 : 16'b0000000111111111;
														assign node11221 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node11224 = (inp[10]) ? node11226 : 16'b0000000111111111;
														assign node11226 = (inp[6]) ? 16'b0000000011111111 : node11227;
															assign node11227 = (inp[5]) ? 16'b0000000011111111 : node11228;
																assign node11228 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node11233 = (inp[10]) ? 16'b0000000001111111 : node11234;
													assign node11234 = (inp[5]) ? 16'b0000000011111111 : node11235;
														assign node11235 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node11240 = (inp[10]) ? node11256 : node11241;
												assign node11241 = (inp[8]) ? node11247 : node11242;
													assign node11242 = (inp[5]) ? node11244 : 16'b0000000011111111;
														assign node11244 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node11247 = (inp[5]) ? node11253 : node11248;
														assign node11248 = (inp[6]) ? 16'b0000000001111111 : node11249;
															assign node11249 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node11253 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node11256 = (inp[5]) ? 16'b0000000000111111 : node11257;
													assign node11257 = (inp[8]) ? node11259 : 16'b0000000001111111;
														assign node11259 = (inp[6]) ? 16'b0000000000011111 : node11260;
															assign node11260 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node11265 = (inp[5]) ? node11283 : node11266;
											assign node11266 = (inp[1]) ? node11268 : 16'b0000000001111111;
												assign node11268 = (inp[12]) ? node11276 : node11269;
													assign node11269 = (inp[10]) ? node11273 : node11270;
														assign node11270 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node11273 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node11276 = (inp[8]) ? node11280 : node11277;
														assign node11277 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node11280 = (inp[6]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node11283 = (inp[10]) ? node11305 : node11284;
												assign node11284 = (inp[8]) ? node11294 : node11285;
													assign node11285 = (inp[6]) ? node11289 : node11286;
														assign node11286 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000111111111;
														assign node11289 = (inp[12]) ? node11291 : 16'b0000000001111111;
															assign node11291 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node11294 = (inp[9]) ? node11302 : node11295;
														assign node11295 = (inp[12]) ? 16'b0000000000111111 : node11296;
															assign node11296 = (inp[1]) ? node11298 : 16'b0000000001111111;
																assign node11298 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node11302 = (inp[6]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node11305 = (inp[6]) ? 16'b0000000000011111 : node11306;
													assign node11306 = (inp[1]) ? node11310 : node11307;
														assign node11307 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node11310 = (inp[12]) ? node11312 : 16'b0000000000111111;
															assign node11312 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
								assign node11316 = (inp[9]) ? node11396 : node11317;
									assign node11317 = (inp[6]) ? node11349 : node11318;
										assign node11318 = (inp[8]) ? node11334 : node11319;
											assign node11319 = (inp[10]) ? node11325 : node11320;
												assign node11320 = (inp[1]) ? 16'b0000000011111111 : node11321;
													assign node11321 = (inp[5]) ? 16'b0000000111111111 : 16'b0000011111111111;
												assign node11325 = (inp[4]) ? 16'b0000000001111111 : node11326;
													assign node11326 = (inp[0]) ? node11330 : node11327;
														assign node11327 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node11330 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node11334 = (inp[5]) ? node11344 : node11335;
												assign node11335 = (inp[10]) ? node11339 : node11336;
													assign node11336 = (inp[4]) ? 16'b0000000111111111 : 16'b0000000011111111;
													assign node11339 = (inp[1]) ? 16'b0000000001111111 : node11340;
														assign node11340 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000111111111;
												assign node11344 = (inp[10]) ? node11346 : 16'b0000000001111111;
													assign node11346 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node11349 = (inp[10]) ? node11379 : node11350;
											assign node11350 = (inp[5]) ? node11368 : node11351;
												assign node11351 = (inp[12]) ? node11359 : node11352;
													assign node11352 = (inp[0]) ? node11356 : node11353;
														assign node11353 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node11356 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node11359 = (inp[1]) ? node11363 : node11360;
														assign node11360 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000111111111;
														assign node11363 = (inp[4]) ? node11365 : 16'b0000000001111111;
															assign node11365 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node11368 = (inp[12]) ? node11374 : node11369;
													assign node11369 = (inp[8]) ? node11371 : 16'b0000000001111111;
														assign node11371 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node11374 = (inp[0]) ? 16'b0000000000011111 : node11375;
														assign node11375 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node11379 = (inp[5]) ? node11389 : node11380;
												assign node11380 = (inp[8]) ? 16'b0000000000111111 : node11381;
													assign node11381 = (inp[4]) ? 16'b0000000000111111 : node11382;
														assign node11382 = (inp[12]) ? node11384 : 16'b0000000001111111;
															assign node11384 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node11389 = (inp[1]) ? node11391 : 16'b0000000000111111;
													assign node11391 = (inp[12]) ? 16'b0000000000011111 : node11392;
														assign node11392 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000000011111;
									assign node11396 = (inp[10]) ? node11436 : node11397;
										assign node11397 = (inp[12]) ? node11409 : node11398;
											assign node11398 = (inp[0]) ? 16'b0000000001111111 : node11399;
												assign node11399 = (inp[1]) ? node11405 : node11400;
													assign node11400 = (inp[5]) ? node11402 : 16'b0000000011111111;
														assign node11402 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node11405 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node11409 = (inp[1]) ? node11427 : node11410;
												assign node11410 = (inp[4]) ? node11418 : node11411;
													assign node11411 = (inp[6]) ? 16'b0000000001111111 : node11412;
														assign node11412 = (inp[5]) ? node11414 : 16'b0000000011111111;
															assign node11414 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node11418 = (inp[8]) ? node11424 : node11419;
														assign node11419 = (inp[6]) ? 16'b0000000000111111 : node11420;
															assign node11420 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node11424 = (inp[6]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node11427 = (inp[4]) ? node11431 : node11428;
													assign node11428 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node11431 = (inp[5]) ? node11433 : 16'b0000000000011111;
														assign node11433 = (inp[0]) ? 16'b0000000000001111 : 16'b0000000000011111;
										assign node11436 = (inp[6]) ? node11462 : node11437;
											assign node11437 = (inp[4]) ? node11451 : node11438;
												assign node11438 = (inp[8]) ? node11446 : node11439;
													assign node11439 = (inp[1]) ? node11441 : 16'b0000000011111111;
														assign node11441 = (inp[5]) ? node11443 : 16'b0000000001111111;
															assign node11443 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node11446 = (inp[12]) ? node11448 : 16'b0000000000111111;
														assign node11448 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node11451 = (inp[8]) ? node11455 : node11452;
													assign node11452 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node11455 = (inp[0]) ? node11457 : 16'b0000000000011111;
														assign node11457 = (inp[5]) ? node11459 : 16'b0000000000011111;
															assign node11459 = (inp[1]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node11462 = (inp[12]) ? node11480 : node11463;
												assign node11463 = (inp[0]) ? node11473 : node11464;
													assign node11464 = (inp[5]) ? node11468 : node11465;
														assign node11465 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node11468 = (inp[1]) ? node11470 : 16'b0000000000111111;
															assign node11470 = (inp[4]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node11473 = (inp[8]) ? 16'b0000000000001111 : node11474;
														assign node11474 = (inp[1]) ? 16'b0000000000011111 : node11475;
															assign node11475 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node11480 = (inp[5]) ? node11490 : node11481;
													assign node11481 = (inp[4]) ? node11483 : 16'b0000000000011111;
														assign node11483 = (inp[0]) ? node11485 : 16'b0000000000011111;
															assign node11485 = (inp[8]) ? 16'b0000000000001111 : node11486;
																assign node11486 = (inp[1]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node11490 = (inp[8]) ? node11496 : node11491;
														assign node11491 = (inp[0]) ? 16'b0000000000001111 : node11492;
															assign node11492 = (inp[4]) ? 16'b0000000000001111 : 16'b0000000000111111;
														assign node11496 = (inp[1]) ? node11498 : 16'b0000000000001111;
															assign node11498 = (inp[4]) ? 16'b0000000000000011 : node11499;
																assign node11499 = (inp[0]) ? 16'b0000000000000111 : 16'b0000000000001111;
							assign node11503 = (inp[6]) ? node11713 : node11504;
								assign node11504 = (inp[0]) ? node11610 : node11505;
									assign node11505 = (inp[10]) ? node11551 : node11506;
										assign node11506 = (inp[5]) ? node11528 : node11507;
											assign node11507 = (inp[9]) ? node11519 : node11508;
												assign node11508 = (inp[12]) ? node11512 : node11509;
													assign node11509 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node11512 = (inp[13]) ? 16'b0000000011111111 : node11513;
														assign node11513 = (inp[8]) ? 16'b0000000011111111 : node11514;
															assign node11514 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node11519 = (inp[1]) ? node11521 : 16'b0000000011111111;
													assign node11521 = (inp[13]) ? 16'b0000000001111111 : node11522;
														assign node11522 = (inp[8]) ? 16'b0000000011111111 : node11523;
															assign node11523 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node11528 = (inp[9]) ? node11534 : node11529;
												assign node11529 = (inp[8]) ? 16'b0000000011111111 : node11530;
													assign node11530 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node11534 = (inp[1]) ? node11544 : node11535;
													assign node11535 = (inp[4]) ? node11539 : node11536;
														assign node11536 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000011111111;
														assign node11539 = (inp[12]) ? node11541 : 16'b0000000001111111;
															assign node11541 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node11544 = (inp[12]) ? node11548 : node11545;
														assign node11545 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node11548 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node11551 = (inp[9]) ? node11583 : node11552;
											assign node11552 = (inp[12]) ? node11566 : node11553;
												assign node11553 = (inp[13]) ? node11555 : 16'b0000000011111111;
													assign node11555 = (inp[5]) ? node11559 : node11556;
														assign node11556 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000111111111;
														assign node11559 = (inp[1]) ? 16'b0000000001111111 : node11560;
															assign node11560 = (inp[4]) ? 16'b0000000001111111 : node11561;
																assign node11561 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node11566 = (inp[1]) ? node11574 : node11567;
													assign node11567 = (inp[8]) ? node11571 : node11568;
														assign node11568 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node11571 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node11574 = (inp[8]) ? node11578 : node11575;
														assign node11575 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node11578 = (inp[4]) ? node11580 : 16'b0000000000111111;
															assign node11580 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node11583 = (inp[13]) ? node11595 : node11584;
												assign node11584 = (inp[1]) ? node11590 : node11585;
													assign node11585 = (inp[12]) ? 16'b0000000001111111 : node11586;
														assign node11586 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node11590 = (inp[12]) ? node11592 : 16'b0000000001111111;
														assign node11592 = (inp[4]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node11595 = (inp[12]) ? node11605 : node11596;
													assign node11596 = (inp[5]) ? node11598 : 16'b0000000000111111;
														assign node11598 = (inp[8]) ? 16'b0000000000011111 : node11599;
															assign node11599 = (inp[4]) ? node11601 : 16'b0000000000111111;
																assign node11601 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node11605 = (inp[1]) ? 16'b0000000000011111 : node11606;
														assign node11606 = (inp[5]) ? 16'b0000000000001111 : 16'b0000000000011111;
									assign node11610 = (inp[9]) ? node11654 : node11611;
										assign node11611 = (inp[10]) ? node11635 : node11612;
											assign node11612 = (inp[1]) ? node11624 : node11613;
												assign node11613 = (inp[12]) ? node11617 : node11614;
													assign node11614 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node11617 = (inp[5]) ? node11621 : node11618;
														assign node11618 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node11621 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node11624 = (inp[8]) ? node11632 : node11625;
													assign node11625 = (inp[4]) ? node11629 : node11626;
														assign node11626 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node11629 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node11632 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000000011111;
											assign node11635 = (inp[13]) ? node11643 : node11636;
												assign node11636 = (inp[12]) ? 16'b0000000000111111 : node11637;
													assign node11637 = (inp[4]) ? node11639 : 16'b0000000011111111;
														assign node11639 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node11643 = (inp[4]) ? node11649 : node11644;
													assign node11644 = (inp[1]) ? node11646 : 16'b0000000000111111;
														assign node11646 = (inp[8]) ? 16'b0000000000001111 : 16'b0000000000111111;
													assign node11649 = (inp[12]) ? 16'b0000000000011111 : node11650;
														assign node11650 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node11654 = (inp[4]) ? node11690 : node11655;
											assign node11655 = (inp[12]) ? node11677 : node11656;
												assign node11656 = (inp[1]) ? node11666 : node11657;
													assign node11657 = (inp[8]) ? node11663 : node11658;
														assign node11658 = (inp[10]) ? node11660 : 16'b0000000001111111;
															assign node11660 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node11663 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node11666 = (inp[8]) ? node11672 : node11667;
														assign node11667 = (inp[5]) ? 16'b0000000000111111 : node11668;
															assign node11668 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000011111111;
														assign node11672 = (inp[13]) ? node11674 : 16'b0000000000111111;
															assign node11674 = (inp[5]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node11677 = (inp[1]) ? node11683 : node11678;
													assign node11678 = (inp[10]) ? 16'b0000000000011111 : node11679;
														assign node11679 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node11683 = (inp[10]) ? 16'b0000000000000111 : node11684;
														assign node11684 = (inp[8]) ? node11686 : 16'b0000000000011111;
															assign node11686 = (inp[13]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node11690 = (inp[5]) ? node11700 : node11691;
												assign node11691 = (inp[8]) ? node11695 : node11692;
													assign node11692 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node11695 = (inp[12]) ? node11697 : 16'b0000000000011111;
														assign node11697 = (inp[1]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node11700 = (inp[13]) ? node11708 : node11701;
													assign node11701 = (inp[1]) ? node11703 : 16'b0000000000011111;
														assign node11703 = (inp[12]) ? node11705 : 16'b0000000000001111;
															assign node11705 = (inp[10]) ? 16'b0000000000000111 : 16'b0000000000001111;
													assign node11708 = (inp[8]) ? node11710 : 16'b0000000000001111;
														assign node11710 = (inp[1]) ? 16'b0000000000000011 : 16'b0000000000000111;
								assign node11713 = (inp[12]) ? node11813 : node11714;
									assign node11714 = (inp[9]) ? node11768 : node11715;
										assign node11715 = (inp[10]) ? node11741 : node11716;
											assign node11716 = (inp[0]) ? node11730 : node11717;
												assign node11717 = (inp[4]) ? node11721 : node11718;
													assign node11718 = (inp[5]) ? 16'b0000000011111111 : 16'b0000001111111111;
													assign node11721 = (inp[1]) ? 16'b0000000001111111 : node11722;
														assign node11722 = (inp[13]) ? node11724 : 16'b0000000011111111;
															assign node11724 = (inp[5]) ? 16'b0000000001111111 : node11725;
																assign node11725 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node11730 = (inp[5]) ? node11736 : node11731;
													assign node11731 = (inp[4]) ? node11733 : 16'b0000000001111111;
														assign node11733 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000000111111;
													assign node11736 = (inp[13]) ? node11738 : 16'b0000000000111111;
														assign node11738 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000000011111;
											assign node11741 = (inp[8]) ? node11755 : node11742;
												assign node11742 = (inp[0]) ? node11746 : node11743;
													assign node11743 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000111111111;
													assign node11746 = (inp[1]) ? node11748 : 16'b0000000001111111;
														assign node11748 = (inp[4]) ? 16'b0000000000111111 : node11749;
															assign node11749 = (inp[13]) ? 16'b0000000000111111 : node11750;
																assign node11750 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node11755 = (inp[1]) ? node11763 : node11756;
													assign node11756 = (inp[0]) ? 16'b0000000000011111 : node11757;
														assign node11757 = (inp[13]) ? 16'b0000000000111111 : node11758;
															assign node11758 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node11763 = (inp[4]) ? node11765 : 16'b0000000000011111;
														assign node11765 = (inp[0]) ? 16'b0000000000000111 : 16'b0000000000001111;
										assign node11768 = (inp[13]) ? node11790 : node11769;
											assign node11769 = (inp[5]) ? node11777 : node11770;
												assign node11770 = (inp[8]) ? node11772 : 16'b0000000001111111;
													assign node11772 = (inp[4]) ? 16'b0000000000111111 : node11773;
														assign node11773 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node11777 = (inp[4]) ? node11787 : node11778;
													assign node11778 = (inp[10]) ? node11780 : 16'b0000000001111111;
														assign node11780 = (inp[8]) ? node11782 : 16'b0000000000111111;
															assign node11782 = (inp[1]) ? 16'b0000000000011111 : node11783;
																assign node11783 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node11787 = (inp[1]) ? 16'b0000000000000111 : 16'b0000000000011111;
											assign node11790 = (inp[5]) ? node11806 : node11791;
												assign node11791 = (inp[8]) ? node11799 : node11792;
													assign node11792 = (inp[10]) ? node11794 : 16'b0000000001111111;
														assign node11794 = (inp[0]) ? 16'b0000000000011111 : node11795;
															assign node11795 = (inp[4]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node11799 = (inp[4]) ? node11803 : node11800;
														assign node11800 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node11803 = (inp[1]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node11806 = (inp[10]) ? node11808 : 16'b0000000000011111;
													assign node11808 = (inp[8]) ? 16'b0000000000001111 : node11809;
														assign node11809 = (inp[1]) ? 16'b0000000000001111 : 16'b0000000000011111;
									assign node11813 = (inp[0]) ? node11855 : node11814;
										assign node11814 = (inp[1]) ? node11832 : node11815;
											assign node11815 = (inp[8]) ? node11821 : node11816;
												assign node11816 = (inp[9]) ? node11818 : 16'b0000000001111111;
													assign node11818 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node11821 = (inp[10]) ? 16'b0000000000011111 : node11822;
													assign node11822 = (inp[4]) ? node11828 : node11823;
														assign node11823 = (inp[13]) ? node11825 : 16'b0000000001111111;
															assign node11825 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000001111111;
														assign node11828 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node11832 = (inp[4]) ? node11840 : node11833;
												assign node11833 = (inp[10]) ? node11835 : 16'b0000000000111111;
													assign node11835 = (inp[9]) ? 16'b0000000000011111 : node11836;
														assign node11836 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node11840 = (inp[13]) ? node11846 : node11841;
													assign node11841 = (inp[5]) ? 16'b0000000000011111 : node11842;
														assign node11842 = (inp[9]) ? 16'b0000000000001111 : 16'b0000000000111111;
													assign node11846 = (inp[10]) ? node11848 : 16'b0000000000001111;
														assign node11848 = (inp[9]) ? 16'b0000000000000111 : node11849;
															assign node11849 = (inp[5]) ? node11851 : 16'b0000000000001111;
																assign node11851 = (inp[8]) ? 16'b0000000000000111 : 16'b0000000000001111;
										assign node11855 = (inp[1]) ? node11885 : node11856;
											assign node11856 = (inp[9]) ? node11872 : node11857;
												assign node11857 = (inp[13]) ? node11865 : node11858;
													assign node11858 = (inp[10]) ? node11862 : node11859;
														assign node11859 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node11862 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node11865 = (inp[8]) ? node11867 : 16'b0000000000111111;
														assign node11867 = (inp[5]) ? node11869 : 16'b0000000000011111;
															assign node11869 = (inp[4]) ? 16'b0000000000000111 : 16'b0000000000001111;
												assign node11872 = (inp[13]) ? node11878 : node11873;
													assign node11873 = (inp[10]) ? 16'b0000000000001111 : node11874;
														assign node11874 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node11878 = (inp[5]) ? node11880 : 16'b0000000000001111;
														assign node11880 = (inp[8]) ? node11882 : 16'b0000000000001111;
															assign node11882 = (inp[4]) ? 16'b0000000000000111 : 16'b0000000000001111;
											assign node11885 = (inp[8]) ? node11897 : node11886;
												assign node11886 = (inp[13]) ? node11892 : node11887;
													assign node11887 = (inp[5]) ? node11889 : 16'b0000000000011111;
														assign node11889 = (inp[10]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node11892 = (inp[5]) ? node11894 : 16'b0000000000001111;
														assign node11894 = (inp[10]) ? 16'b0000000000000111 : 16'b0000000000001111;
												assign node11897 = (inp[4]) ? node11911 : node11898;
													assign node11898 = (inp[10]) ? node11902 : node11899;
														assign node11899 = (inp[9]) ? 16'b0000000000001111 : 16'b0000000000011111;
														assign node11902 = (inp[9]) ? node11908 : node11903;
															assign node11903 = (inp[5]) ? node11905 : 16'b0000000000001111;
																assign node11905 = (inp[13]) ? 16'b0000000000000111 : 16'b0000000000001111;
															assign node11908 = (inp[13]) ? 16'b0000000000000011 : 16'b0000000000000111;
													assign node11911 = (inp[9]) ? node11913 : 16'b0000000000000111;
														assign node11913 = (inp[5]) ? 16'b0000000000000011 : 16'b0000000000000111;
		assign node11916 = (inp[0]) ? node18124 : node11917;
			assign node11917 = (inp[12]) ? node15031 : node11918;
				assign node11918 = (inp[9]) ? node13464 : node11919;
					assign node11919 = (inp[2]) ? node12709 : node11920;
						assign node11920 = (inp[14]) ? node12298 : node11921;
							assign node11921 = (inp[5]) ? node12115 : node11922;
								assign node11922 = (inp[10]) ? node12016 : node11923;
									assign node11923 = (inp[8]) ? node11969 : node11924;
										assign node11924 = (inp[6]) ? node11952 : node11925;
											assign node11925 = (inp[4]) ? node11937 : node11926;
												assign node11926 = (inp[11]) ? node11932 : node11927;
													assign node11927 = (inp[15]) ? 16'b0001111111111111 : node11928;
														assign node11928 = (inp[1]) ? 16'b0001111111111111 : 16'b0011111111111111;
													assign node11932 = (inp[13]) ? 16'b0000111111111111 : node11933;
														assign node11933 = (inp[15]) ? 16'b0000111111111111 : 16'b0001111111111111;
												assign node11937 = (inp[13]) ? node11943 : node11938;
													assign node11938 = (inp[11]) ? 16'b0000111111111111 : node11939;
														assign node11939 = (inp[1]) ? 16'b0000111111111111 : 16'b0001111111111111;
													assign node11943 = (inp[11]) ? 16'b0000011111111111 : node11944;
														assign node11944 = (inp[15]) ? node11948 : node11945;
															assign node11945 = (inp[3]) ? 16'b0000111111111111 : 16'b0001111111111111;
															assign node11948 = (inp[3]) ? 16'b0000011111111111 : 16'b0000111111111111;
											assign node11952 = (inp[11]) ? node11966 : node11953;
												assign node11953 = (inp[13]) ? node11955 : 16'b0000111111111111;
													assign node11955 = (inp[4]) ? 16'b0000011111111111 : node11956;
														assign node11956 = (inp[1]) ? node11960 : node11957;
															assign node11957 = (inp[3]) ? 16'b0000111111111111 : 16'b0001111111111111;
															assign node11960 = (inp[15]) ? 16'b0000011111111111 : node11961;
																assign node11961 = (inp[3]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node11966 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
										assign node11969 = (inp[3]) ? node11991 : node11970;
											assign node11970 = (inp[1]) ? node11984 : node11971;
												assign node11971 = (inp[4]) ? node11973 : 16'b0000111111111111;
													assign node11973 = (inp[11]) ? node11981 : node11974;
														assign node11974 = (inp[6]) ? 16'b0000011111111111 : node11975;
															assign node11975 = (inp[15]) ? 16'b0000111111111111 : node11976;
																assign node11976 = (inp[13]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node11981 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node11984 = (inp[4]) ? 16'b0000001111111111 : node11985;
													assign node11985 = (inp[11]) ? node11987 : 16'b0000011111111111;
														assign node11987 = (inp[15]) ? 16'b0000001111111111 : 16'b0000111111111111;
											assign node11991 = (inp[4]) ? node12005 : node11992;
												assign node11992 = (inp[15]) ? node11996 : node11993;
													assign node11993 = (inp[11]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node11996 = (inp[1]) ? node11998 : 16'b0000011111111111;
														assign node11998 = (inp[6]) ? 16'b0000000111111111 : node11999;
															assign node11999 = (inp[11]) ? node12001 : 16'b0000001111111111;
																assign node12001 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node12005 = (inp[11]) ? node12011 : node12006;
													assign node12006 = (inp[13]) ? 16'b0000001111111111 : node12007;
														assign node12007 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node12011 = (inp[6]) ? 16'b0000000111111111 : node12012;
														assign node12012 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
									assign node12016 = (inp[4]) ? node12074 : node12017;
										assign node12017 = (inp[13]) ? node12043 : node12018;
											assign node12018 = (inp[6]) ? node12030 : node12019;
												assign node12019 = (inp[3]) ? node12025 : node12020;
													assign node12020 = (inp[11]) ? 16'b0000111111111111 : node12021;
														assign node12021 = (inp[8]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node12025 = (inp[11]) ? 16'b0000011111111111 : node12026;
														assign node12026 = (inp[15]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node12030 = (inp[15]) ? node12032 : 16'b0000111111111111;
													assign node12032 = (inp[1]) ? 16'b0000001111111111 : node12033;
														assign node12033 = (inp[3]) ? node12039 : node12034;
															assign node12034 = (inp[8]) ? 16'b0000011111111111 : node12035;
																assign node12035 = (inp[11]) ? 16'b0000011111111111 : 16'b0000111111111111;
															assign node12039 = (inp[11]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node12043 = (inp[15]) ? node12061 : node12044;
												assign node12044 = (inp[11]) ? node12054 : node12045;
													assign node12045 = (inp[1]) ? 16'b0000001111111111 : node12046;
														assign node12046 = (inp[3]) ? 16'b0000011111111111 : node12047;
															assign node12047 = (inp[8]) ? node12049 : 16'b0000111111111111;
																assign node12049 = (inp[6]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node12054 = (inp[6]) ? node12058 : node12055;
														assign node12055 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node12058 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node12061 = (inp[8]) ? node12067 : node12062;
													assign node12062 = (inp[1]) ? node12064 : 16'b0000011111111111;
														assign node12064 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node12067 = (inp[11]) ? 16'b0000000001111111 : node12068;
														assign node12068 = (inp[1]) ? node12070 : 16'b0000000111111111;
															assign node12070 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node12074 = (inp[6]) ? node12090 : node12075;
											assign node12075 = (inp[15]) ? node12083 : node12076;
												assign node12076 = (inp[8]) ? 16'b0000001111111111 : node12077;
													assign node12077 = (inp[13]) ? 16'b0000001111111111 : node12078;
														assign node12078 = (inp[1]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node12083 = (inp[3]) ? 16'b0000000111111111 : node12084;
													assign node12084 = (inp[13]) ? 16'b0000001111111111 : node12085;
														assign node12085 = (inp[1]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node12090 = (inp[11]) ? node12104 : node12091;
												assign node12091 = (inp[3]) ? node12099 : node12092;
													assign node12092 = (inp[15]) ? 16'b0000001111111111 : node12093;
														assign node12093 = (inp[8]) ? node12095 : 16'b0000011111111111;
															assign node12095 = (inp[1]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node12099 = (inp[8]) ? node12101 : 16'b0000001111111111;
														assign node12101 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node12104 = (inp[15]) ? node12108 : node12105;
													assign node12105 = (inp[3]) ? 16'b0000000111111111 : 16'b0000000011111111;
													assign node12108 = (inp[3]) ? node12112 : node12109;
														assign node12109 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node12112 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
								assign node12115 = (inp[4]) ? node12217 : node12116;
									assign node12116 = (inp[8]) ? node12176 : node12117;
										assign node12117 = (inp[6]) ? node12143 : node12118;
											assign node12118 = (inp[3]) ? node12130 : node12119;
												assign node12119 = (inp[10]) ? 16'b0000011111111111 : node12120;
													assign node12120 = (inp[11]) ? node12124 : node12121;
														assign node12121 = (inp[15]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node12124 = (inp[15]) ? node12126 : 16'b0000111111111111;
															assign node12126 = (inp[13]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node12130 = (inp[1]) ? node12138 : node12131;
													assign node12131 = (inp[11]) ? 16'b0000011111111111 : node12132;
														assign node12132 = (inp[15]) ? 16'b0000011111111111 : node12133;
															assign node12133 = (inp[13]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node12138 = (inp[10]) ? 16'b0000001111111111 : node12139;
														assign node12139 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node12143 = (inp[11]) ? node12157 : node12144;
												assign node12144 = (inp[3]) ? node12150 : node12145;
													assign node12145 = (inp[13]) ? 16'b0000011111111111 : node12146;
														assign node12146 = (inp[1]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node12150 = (inp[13]) ? node12154 : node12151;
														assign node12151 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node12154 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node12157 = (inp[1]) ? node12167 : node12158;
													assign node12158 = (inp[15]) ? node12164 : node12159;
														assign node12159 = (inp[13]) ? 16'b0000001111111111 : node12160;
															assign node12160 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node12164 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node12167 = (inp[15]) ? 16'b0000000011111111 : node12168;
														assign node12168 = (inp[3]) ? 16'b0000000111111111 : node12169;
															assign node12169 = (inp[13]) ? node12171 : 16'b0000001111111111;
																assign node12171 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node12176 = (inp[15]) ? node12194 : node12177;
											assign node12177 = (inp[11]) ? node12187 : node12178;
												assign node12178 = (inp[13]) ? node12182 : node12179;
													assign node12179 = (inp[3]) ? 16'b0000111111111111 : 16'b0000011111111111;
													assign node12182 = (inp[1]) ? 16'b0000001111111111 : node12183;
														assign node12183 = (inp[6]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node12187 = (inp[3]) ? 16'b0000000111111111 : node12188;
													assign node12188 = (inp[6]) ? node12190 : 16'b0000001111111111;
														assign node12190 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node12194 = (inp[1]) ? node12210 : node12195;
												assign node12195 = (inp[10]) ? node12203 : node12196;
													assign node12196 = (inp[11]) ? node12198 : 16'b0000001111111111;
														assign node12198 = (inp[6]) ? 16'b0000000111111111 : node12199;
															assign node12199 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node12203 = (inp[11]) ? node12207 : node12204;
														assign node12204 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node12207 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000111111111;
												assign node12210 = (inp[6]) ? 16'b0000000011111111 : node12211;
													assign node12211 = (inp[13]) ? node12213 : 16'b0000000111111111;
														assign node12213 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000111111111;
									assign node12217 = (inp[15]) ? node12259 : node12218;
										assign node12218 = (inp[3]) ? node12242 : node12219;
											assign node12219 = (inp[10]) ? node12231 : node12220;
												assign node12220 = (inp[8]) ? node12224 : node12221;
													assign node12221 = (inp[1]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node12224 = (inp[6]) ? 16'b0000001111111111 : node12225;
														assign node12225 = (inp[11]) ? node12227 : 16'b0000011111111111;
															assign node12227 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node12231 = (inp[11]) ? node12239 : node12232;
													assign node12232 = (inp[1]) ? node12236 : node12233;
														assign node12233 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node12236 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node12239 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node12242 = (inp[8]) ? node12254 : node12243;
												assign node12243 = (inp[1]) ? node12245 : 16'b0000001111111111;
													assign node12245 = (inp[6]) ? node12249 : node12246;
														assign node12246 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node12249 = (inp[13]) ? 16'b0000000011111111 : node12250;
															assign node12250 = (inp[10]) ? 16'b0000000011111111 : 16'b0000001111111111;
												assign node12254 = (inp[10]) ? 16'b0000000011111111 : node12255;
													assign node12255 = (inp[13]) ? 16'b0000000111111111 : 16'b0000000011111111;
										assign node12259 = (inp[3]) ? node12271 : node12260;
											assign node12260 = (inp[8]) ? node12266 : node12261;
												assign node12261 = (inp[13]) ? 16'b0000000111111111 : node12262;
													assign node12262 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node12266 = (inp[11]) ? 16'b0000000011111111 : node12267;
													assign node12267 = (inp[6]) ? 16'b0000001111111111 : 16'b0000000111111111;
											assign node12271 = (inp[13]) ? node12281 : node12272;
												assign node12272 = (inp[8]) ? node12274 : 16'b0000000111111111;
													assign node12274 = (inp[1]) ? 16'b0000000001111111 : node12275;
														assign node12275 = (inp[10]) ? node12277 : 16'b0000000111111111;
															assign node12277 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node12281 = (inp[1]) ? node12293 : node12282;
													assign node12282 = (inp[8]) ? node12286 : node12283;
														assign node12283 = (inp[6]) ? 16'b0000000111111111 : 16'b0000000011111111;
														assign node12286 = (inp[10]) ? 16'b0000000001111111 : node12287;
															assign node12287 = (inp[6]) ? node12289 : 16'b0000000011111111;
																assign node12289 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node12293 = (inp[6]) ? node12295 : 16'b0000000011111111;
														assign node12295 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
							assign node12298 = (inp[13]) ? node12468 : node12299;
								assign node12299 = (inp[4]) ? node12375 : node12300;
									assign node12300 = (inp[11]) ? node12338 : node12301;
										assign node12301 = (inp[8]) ? node12315 : node12302;
											assign node12302 = (inp[15]) ? 16'b0000001111111111 : node12303;
												assign node12303 = (inp[3]) ? 16'b0000011111111111 : node12304;
													assign node12304 = (inp[5]) ? node12306 : 16'b0000111111111111;
														assign node12306 = (inp[10]) ? node12308 : 16'b0000111111111111;
															assign node12308 = (inp[6]) ? 16'b0000011111111111 : node12309;
																assign node12309 = (inp[1]) ? 16'b0000011111111111 : 16'b0000111111111111;
											assign node12315 = (inp[10]) ? node12331 : node12316;
												assign node12316 = (inp[1]) ? node12326 : node12317;
													assign node12317 = (inp[15]) ? node12321 : node12318;
														assign node12318 = (inp[6]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node12321 = (inp[5]) ? node12323 : 16'b0000011111111111;
															assign node12323 = (inp[6]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node12326 = (inp[3]) ? 16'b0000001111111111 : node12327;
														assign node12327 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node12331 = (inp[6]) ? node12333 : 16'b0000001111111111;
													assign node12333 = (inp[3]) ? node12335 : 16'b0000001111111111;
														assign node12335 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node12338 = (inp[3]) ? node12356 : node12339;
											assign node12339 = (inp[15]) ? node12347 : node12340;
												assign node12340 = (inp[1]) ? 16'b0000001111111111 : node12341;
													assign node12341 = (inp[5]) ? 16'b0000001111111111 : node12342;
														assign node12342 = (inp[10]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node12347 = (inp[10]) ? node12349 : 16'b0000001111111111;
													assign node12349 = (inp[1]) ? 16'b0000000111111111 : node12350;
														assign node12350 = (inp[6]) ? node12352 : 16'b0000001111111111;
															assign node12352 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node12356 = (inp[8]) ? node12362 : node12357;
												assign node12357 = (inp[5]) ? node12359 : 16'b0000001111111111;
													assign node12359 = (inp[6]) ? 16'b0000000011111111 : 16'b0000001111111111;
												assign node12362 = (inp[6]) ? node12368 : node12363;
													assign node12363 = (inp[15]) ? node12365 : 16'b0000001111111111;
														assign node12365 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node12368 = (inp[15]) ? node12372 : node12369;
														assign node12369 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node12372 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node12375 = (inp[8]) ? node12415 : node12376;
										assign node12376 = (inp[3]) ? node12398 : node12377;
											assign node12377 = (inp[15]) ? node12385 : node12378;
												assign node12378 = (inp[6]) ? node12380 : 16'b0000011111111111;
													assign node12380 = (inp[10]) ? node12382 : 16'b0000001111111111;
														assign node12382 = (inp[11]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node12385 = (inp[10]) ? node12391 : node12386;
													assign node12386 = (inp[11]) ? 16'b0000001111111111 : node12387;
														assign node12387 = (inp[1]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node12391 = (inp[1]) ? node12395 : node12392;
														assign node12392 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node12395 = (inp[6]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node12398 = (inp[11]) ? node12408 : node12399;
												assign node12399 = (inp[5]) ? node12401 : 16'b0000011111111111;
													assign node12401 = (inp[10]) ? node12403 : 16'b0000001111111111;
														assign node12403 = (inp[6]) ? 16'b0000000111111111 : node12404;
															assign node12404 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node12408 = (inp[5]) ? node12410 : 16'b0000000111111111;
													assign node12410 = (inp[1]) ? node12412 : 16'b0000000111111111;
														assign node12412 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node12415 = (inp[1]) ? node12449 : node12416;
											assign node12416 = (inp[3]) ? node12442 : node12417;
												assign node12417 = (inp[5]) ? node12429 : node12418;
													assign node12418 = (inp[15]) ? node12424 : node12419;
														assign node12419 = (inp[6]) ? node12421 : 16'b0000111111111111;
															assign node12421 = (inp[11]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node12424 = (inp[6]) ? node12426 : 16'b0000001111111111;
															assign node12426 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node12429 = (inp[6]) ? node12435 : node12430;
														assign node12430 = (inp[11]) ? node12432 : 16'b0000011111111111;
															assign node12432 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node12435 = (inp[15]) ? node12437 : 16'b0000000111111111;
															assign node12437 = (inp[10]) ? 16'b0000000011111111 : node12438;
																assign node12438 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node12442 = (inp[15]) ? node12444 : 16'b0000000111111111;
													assign node12444 = (inp[6]) ? node12446 : 16'b0000000111111111;
														assign node12446 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node12449 = (inp[5]) ? node12461 : node12450;
												assign node12450 = (inp[10]) ? node12452 : 16'b0000000111111111;
													assign node12452 = (inp[11]) ? node12458 : node12453;
														assign node12453 = (inp[6]) ? node12455 : 16'b0000000111111111;
															assign node12455 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000111111111;
														assign node12458 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node12461 = (inp[3]) ? 16'b0000000001111111 : node12462;
													assign node12462 = (inp[6]) ? node12464 : 16'b0000000011111111;
														assign node12464 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
								assign node12468 = (inp[5]) ? node12590 : node12469;
									assign node12469 = (inp[10]) ? node12523 : node12470;
										assign node12470 = (inp[1]) ? node12492 : node12471;
											assign node12471 = (inp[15]) ? node12477 : node12472;
												assign node12472 = (inp[6]) ? node12474 : 16'b0000011111111111;
													assign node12474 = (inp[4]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node12477 = (inp[8]) ? node12485 : node12478;
													assign node12478 = (inp[11]) ? 16'b0000001111111111 : node12479;
														assign node12479 = (inp[4]) ? 16'b0000001111111111 : node12480;
															assign node12480 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node12485 = (inp[11]) ? node12489 : node12486;
														assign node12486 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node12489 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node12492 = (inp[6]) ? node12510 : node12493;
												assign node12493 = (inp[8]) ? node12501 : node12494;
													assign node12494 = (inp[3]) ? node12496 : 16'b0000011111111111;
														assign node12496 = (inp[11]) ? node12498 : 16'b0000001111111111;
															assign node12498 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node12501 = (inp[4]) ? 16'b0000000011111111 : node12502;
														assign node12502 = (inp[11]) ? node12504 : 16'b0000001111111111;
															assign node12504 = (inp[15]) ? 16'b0000000111111111 : node12505;
																assign node12505 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node12510 = (inp[15]) ? node12516 : node12511;
													assign node12511 = (inp[3]) ? 16'b0000000111111111 : node12512;
														assign node12512 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node12516 = (inp[8]) ? 16'b0000000011111111 : node12517;
														assign node12517 = (inp[3]) ? node12519 : 16'b0000000111111111;
															assign node12519 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node12523 = (inp[6]) ? node12561 : node12524;
											assign node12524 = (inp[1]) ? node12540 : node12525;
												assign node12525 = (inp[15]) ? node12535 : node12526;
													assign node12526 = (inp[11]) ? node12532 : node12527;
														assign node12527 = (inp[4]) ? node12529 : 16'b0000011111111111;
															assign node12529 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node12532 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node12535 = (inp[4]) ? 16'b0000000111111111 : node12536;
														assign node12536 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node12540 = (inp[11]) ? node12550 : node12541;
													assign node12541 = (inp[3]) ? node12543 : 16'b0000001111111111;
														assign node12543 = (inp[15]) ? node12545 : 16'b0000000111111111;
															assign node12545 = (inp[4]) ? 16'b0000000011111111 : node12546;
																assign node12546 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node12550 = (inp[3]) ? node12558 : node12551;
														assign node12551 = (inp[4]) ? 16'b0000000011111111 : node12552;
															assign node12552 = (inp[15]) ? node12554 : 16'b0000000111111111;
																assign node12554 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node12558 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000001111111;
											assign node12561 = (inp[11]) ? node12575 : node12562;
												assign node12562 = (inp[3]) ? node12568 : node12563;
													assign node12563 = (inp[15]) ? 16'b0000000111111111 : node12564;
														assign node12564 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node12568 = (inp[8]) ? node12570 : 16'b0000000111111111;
														assign node12570 = (inp[15]) ? node12572 : 16'b0000000011111111;
															assign node12572 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node12575 = (inp[15]) ? node12583 : node12576;
													assign node12576 = (inp[3]) ? node12578 : 16'b0000000011111111;
														assign node12578 = (inp[8]) ? 16'b0000000001111111 : node12579;
															assign node12579 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node12583 = (inp[8]) ? node12585 : 16'b0000000001111111;
														assign node12585 = (inp[4]) ? 16'b0000000000111111 : node12586;
															assign node12586 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node12590 = (inp[15]) ? node12650 : node12591;
										assign node12591 = (inp[8]) ? node12625 : node12592;
											assign node12592 = (inp[10]) ? node12610 : node12593;
												assign node12593 = (inp[1]) ? node12601 : node12594;
													assign node12594 = (inp[3]) ? 16'b0000001111111111 : node12595;
														assign node12595 = (inp[4]) ? node12597 : 16'b0000011111111111;
															assign node12597 = (inp[11]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node12601 = (inp[6]) ? node12607 : node12602;
														assign node12602 = (inp[3]) ? node12604 : 16'b0000001111111111;
															assign node12604 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node12607 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node12610 = (inp[11]) ? node12618 : node12611;
													assign node12611 = (inp[6]) ? node12615 : node12612;
														assign node12612 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node12615 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node12618 = (inp[4]) ? 16'b0000000001111111 : node12619;
														assign node12619 = (inp[1]) ? 16'b0000000011111111 : node12620;
															assign node12620 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node12625 = (inp[6]) ? node12641 : node12626;
												assign node12626 = (inp[4]) ? node12634 : node12627;
													assign node12627 = (inp[11]) ? node12629 : 16'b0000000111111111;
														assign node12629 = (inp[1]) ? 16'b0000000011111111 : node12630;
															assign node12630 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node12634 = (inp[1]) ? node12638 : node12635;
														assign node12635 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node12638 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node12641 = (inp[1]) ? node12647 : node12642;
													assign node12642 = (inp[4]) ? node12644 : 16'b0000000111111111;
														assign node12644 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node12647 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node12650 = (inp[10]) ? node12682 : node12651;
											assign node12651 = (inp[6]) ? node12667 : node12652;
												assign node12652 = (inp[3]) ? node12660 : node12653;
													assign node12653 = (inp[1]) ? node12657 : node12654;
														assign node12654 = (inp[11]) ? 16'b0000000111111111 : 16'b0000011111111111;
														assign node12657 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node12660 = (inp[1]) ? node12664 : node12661;
														assign node12661 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node12664 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node12667 = (inp[8]) ? node12677 : node12668;
													assign node12668 = (inp[4]) ? node12670 : 16'b0000000011111111;
														assign node12670 = (inp[1]) ? node12672 : 16'b0000000011111111;
															assign node12672 = (inp[3]) ? 16'b0000000001111111 : node12673;
																assign node12673 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node12677 = (inp[3]) ? 16'b0000000000111111 : node12678;
														assign node12678 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node12682 = (inp[3]) ? node12702 : node12683;
												assign node12683 = (inp[8]) ? node12693 : node12684;
													assign node12684 = (inp[1]) ? node12686 : 16'b0000000111111111;
														assign node12686 = (inp[4]) ? 16'b0000000001111111 : node12687;
															assign node12687 = (inp[11]) ? node12689 : 16'b0000000011111111;
																assign node12689 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node12693 = (inp[11]) ? node12695 : 16'b0000000001111111;
														assign node12695 = (inp[1]) ? 16'b0000000000111111 : node12696;
															assign node12696 = (inp[6]) ? node12698 : 16'b0000000001111111;
																assign node12698 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node12702 = (inp[8]) ? node12706 : node12703;
													assign node12703 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000011111111;
													assign node12706 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000111111;
						assign node12709 = (inp[10]) ? node13071 : node12710;
							assign node12710 = (inp[15]) ? node12898 : node12711;
								assign node12711 = (inp[4]) ? node12813 : node12712;
									assign node12712 = (inp[1]) ? node12770 : node12713;
										assign node12713 = (inp[13]) ? node12753 : node12714;
											assign node12714 = (inp[11]) ? node12730 : node12715;
												assign node12715 = (inp[14]) ? node12721 : node12716;
													assign node12716 = (inp[8]) ? 16'b0000111111111111 : node12717;
														assign node12717 = (inp[6]) ? 16'b0000111111111111 : 16'b0001111111111111;
													assign node12721 = (inp[8]) ? 16'b0000011111111111 : node12722;
														assign node12722 = (inp[5]) ? 16'b0000011111111111 : node12723;
															assign node12723 = (inp[3]) ? 16'b0000111111111111 : node12724;
																assign node12724 = (inp[6]) ? 16'b0000111111111111 : 16'b0001111111111111;
												assign node12730 = (inp[8]) ? node12748 : node12731;
													assign node12731 = (inp[6]) ? node12739 : node12732;
														assign node12732 = (inp[5]) ? node12734 : 16'b0000111111111111;
															assign node12734 = (inp[14]) ? 16'b0000011111111111 : node12735;
																assign node12735 = (inp[3]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node12739 = (inp[14]) ? node12745 : node12740;
															assign node12740 = (inp[5]) ? node12742 : 16'b0000011111111111;
																assign node12742 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
															assign node12745 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node12748 = (inp[3]) ? node12750 : 16'b0000001111111111;
														assign node12750 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node12753 = (inp[8]) ? node12763 : node12754;
												assign node12754 = (inp[14]) ? node12756 : 16'b0000011111111111;
													assign node12756 = (inp[5]) ? node12760 : node12757;
														assign node12757 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node12760 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node12763 = (inp[6]) ? node12765 : 16'b0000001111111111;
													assign node12765 = (inp[3]) ? 16'b0000000011111111 : node12766;
														assign node12766 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node12770 = (inp[3]) ? node12798 : node12771;
											assign node12771 = (inp[5]) ? node12789 : node12772;
												assign node12772 = (inp[11]) ? node12782 : node12773;
													assign node12773 = (inp[14]) ? node12779 : node12774;
														assign node12774 = (inp[6]) ? 16'b0000011111111111 : node12775;
															assign node12775 = (inp[13]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node12779 = (inp[8]) ? 16'b0000000111111111 : 16'b0000011111111111;
													assign node12782 = (inp[13]) ? 16'b0000001111111111 : node12783;
														assign node12783 = (inp[6]) ? 16'b0000001111111111 : node12784;
															assign node12784 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node12789 = (inp[13]) ? node12791 : 16'b0000001111111111;
													assign node12791 = (inp[14]) ? node12795 : node12792;
														assign node12792 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node12795 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node12798 = (inp[11]) ? node12802 : node12799;
												assign node12799 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node12802 = (inp[8]) ? node12804 : 16'b0000000111111111;
													assign node12804 = (inp[5]) ? node12808 : node12805;
														assign node12805 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node12808 = (inp[6]) ? node12810 : 16'b0000000011111111;
															assign node12810 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node12813 = (inp[3]) ? node12857 : node12814;
										assign node12814 = (inp[13]) ? node12830 : node12815;
											assign node12815 = (inp[8]) ? node12823 : node12816;
												assign node12816 = (inp[11]) ? node12820 : node12817;
													assign node12817 = (inp[1]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node12820 = (inp[1]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node12823 = (inp[5]) ? node12825 : 16'b0000001111111111;
													assign node12825 = (inp[6]) ? node12827 : 16'b0000001111111111;
														assign node12827 = (inp[11]) ? 16'b0000000111111111 : 16'b0000000011111111;
											assign node12830 = (inp[11]) ? node12840 : node12831;
												assign node12831 = (inp[14]) ? 16'b0000001111111111 : node12832;
													assign node12832 = (inp[8]) ? node12834 : 16'b0000001111111111;
														assign node12834 = (inp[6]) ? 16'b0000000111111111 : node12835;
															assign node12835 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node12840 = (inp[8]) ? node12850 : node12841;
													assign node12841 = (inp[6]) ? node12847 : node12842;
														assign node12842 = (inp[5]) ? 16'b0000000111111111 : node12843;
															assign node12843 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node12847 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node12850 = (inp[5]) ? node12854 : node12851;
														assign node12851 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node12854 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node12857 = (inp[13]) ? node12879 : node12858;
											assign node12858 = (inp[5]) ? node12870 : node12859;
												assign node12859 = (inp[11]) ? node12865 : node12860;
													assign node12860 = (inp[14]) ? node12862 : 16'b0000011111111111;
														assign node12862 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node12865 = (inp[14]) ? 16'b0000000111111111 : node12866;
														assign node12866 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node12870 = (inp[6]) ? node12872 : 16'b0000000111111111;
													assign node12872 = (inp[11]) ? node12876 : node12873;
														assign node12873 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node12876 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node12879 = (inp[5]) ? node12891 : node12880;
												assign node12880 = (inp[8]) ? 16'b0000000011111111 : node12881;
													assign node12881 = (inp[14]) ? node12883 : 16'b0000001111111111;
														assign node12883 = (inp[1]) ? node12885 : 16'b0000000111111111;
															assign node12885 = (inp[11]) ? 16'b0000000011111111 : node12886;
																assign node12886 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node12891 = (inp[1]) ? node12893 : 16'b0000000011111111;
													assign node12893 = (inp[14]) ? 16'b0000000001111111 : node12894;
														assign node12894 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000001111111;
								assign node12898 = (inp[13]) ? node12992 : node12899;
									assign node12899 = (inp[14]) ? node12941 : node12900;
										assign node12900 = (inp[5]) ? node12922 : node12901;
											assign node12901 = (inp[1]) ? node12909 : node12902;
												assign node12902 = (inp[6]) ? node12906 : node12903;
													assign node12903 = (inp[3]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node12906 = (inp[4]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node12909 = (inp[4]) ? node12917 : node12910;
													assign node12910 = (inp[11]) ? 16'b0000001111111111 : node12911;
														assign node12911 = (inp[3]) ? node12913 : 16'b0000011111111111;
															assign node12913 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node12917 = (inp[3]) ? node12919 : 16'b0000001111111111;
														assign node12919 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node12922 = (inp[1]) ? node12934 : node12923;
												assign node12923 = (inp[8]) ? node12929 : node12924;
													assign node12924 = (inp[3]) ? node12926 : 16'b0000001111111111;
														assign node12926 = (inp[4]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node12929 = (inp[3]) ? 16'b0000000111111111 : node12930;
														assign node12930 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node12934 = (inp[8]) ? node12936 : 16'b0000000111111111;
													assign node12936 = (inp[11]) ? 16'b0000000001111111 : node12937;
														assign node12937 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node12941 = (inp[6]) ? node12969 : node12942;
											assign node12942 = (inp[8]) ? node12960 : node12943;
												assign node12943 = (inp[4]) ? node12951 : node12944;
													assign node12944 = (inp[1]) ? node12948 : node12945;
														assign node12945 = (inp[11]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node12948 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node12951 = (inp[3]) ? node12955 : node12952;
														assign node12952 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node12955 = (inp[11]) ? 16'b0000000011111111 : node12956;
															assign node12956 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node12960 = (inp[11]) ? node12964 : node12961;
													assign node12961 = (inp[3]) ? 16'b0000000011111111 : 16'b0000001111111111;
													assign node12964 = (inp[4]) ? 16'b0000000011111111 : node12965;
														assign node12965 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node12969 = (inp[11]) ? node12977 : node12970;
												assign node12970 = (inp[1]) ? 16'b0000000011111111 : node12971;
													assign node12971 = (inp[8]) ? node12973 : 16'b0000000111111111;
														assign node12973 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node12977 = (inp[8]) ? node12985 : node12978;
													assign node12978 = (inp[3]) ? node12982 : node12979;
														assign node12979 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node12982 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node12985 = (inp[3]) ? 16'b0000000001111111 : node12986;
														assign node12986 = (inp[4]) ? 16'b0000000001111111 : node12987;
															assign node12987 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node12992 = (inp[14]) ? node13052 : node12993;
										assign node12993 = (inp[8]) ? node13017 : node12994;
											assign node12994 = (inp[5]) ? node13004 : node12995;
												assign node12995 = (inp[4]) ? node12999 : node12996;
													assign node12996 = (inp[1]) ? 16'b0000000111111111 : 16'b0000011111111111;
													assign node12999 = (inp[3]) ? 16'b0000000111111111 : node13000;
														assign node13000 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node13004 = (inp[4]) ? node13012 : node13005;
													assign node13005 = (inp[6]) ? node13009 : node13006;
														assign node13006 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node13009 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node13012 = (inp[3]) ? 16'b0000000000111111 : node13013;
														assign node13013 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node13017 = (inp[6]) ? node13029 : node13018;
												assign node13018 = (inp[1]) ? node13026 : node13019;
													assign node13019 = (inp[3]) ? node13023 : node13020;
														assign node13020 = (inp[5]) ? 16'b0000001111111111 : 16'b0000000111111111;
														assign node13023 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node13026 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node13029 = (inp[4]) ? node13039 : node13030;
													assign node13030 = (inp[11]) ? node13032 : 16'b0000000111111111;
														assign node13032 = (inp[1]) ? 16'b0000000001111111 : node13033;
															assign node13033 = (inp[3]) ? node13035 : 16'b0000000011111111;
																assign node13035 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node13039 = (inp[5]) ? node13045 : node13040;
														assign node13040 = (inp[1]) ? 16'b0000000001111111 : node13041;
															assign node13041 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node13045 = (inp[1]) ? 16'b0000000000111111 : node13046;
															assign node13046 = (inp[11]) ? node13048 : 16'b0000000001111111;
																assign node13048 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node13052 = (inp[4]) ? node13060 : node13053;
											assign node13053 = (inp[5]) ? 16'b0000000001111111 : node13054;
												assign node13054 = (inp[3]) ? node13056 : 16'b0000000111111111;
													assign node13056 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node13060 = (inp[3]) ? node13062 : 16'b0000000001111111;
												assign node13062 = (inp[5]) ? node13066 : node13063;
													assign node13063 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node13066 = (inp[1]) ? node13068 : 16'b0000000000111111;
														assign node13068 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
							assign node13071 = (inp[11]) ? node13261 : node13072;
								assign node13072 = (inp[1]) ? node13162 : node13073;
									assign node13073 = (inp[5]) ? node13125 : node13074;
										assign node13074 = (inp[13]) ? node13100 : node13075;
											assign node13075 = (inp[8]) ? node13089 : node13076;
												assign node13076 = (inp[3]) ? 16'b0000001111111111 : node13077;
													assign node13077 = (inp[4]) ? node13085 : node13078;
														assign node13078 = (inp[6]) ? 16'b0000011111111111 : node13079;
															assign node13079 = (inp[14]) ? node13081 : 16'b0000111111111111;
																assign node13081 = (inp[15]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node13085 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node13089 = (inp[15]) ? node13095 : node13090;
													assign node13090 = (inp[3]) ? 16'b0000001111111111 : node13091;
														assign node13091 = (inp[6]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node13095 = (inp[6]) ? 16'b0000000111111111 : node13096;
														assign node13096 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node13100 = (inp[15]) ? node13108 : node13101;
												assign node13101 = (inp[3]) ? 16'b0000000111111111 : node13102;
													assign node13102 = (inp[4]) ? 16'b0000001111111111 : node13103;
														assign node13103 = (inp[6]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node13108 = (inp[8]) ? node13116 : node13109;
													assign node13109 = (inp[14]) ? node13111 : 16'b0000001111111111;
														assign node13111 = (inp[3]) ? node13113 : 16'b0000000111111111;
															assign node13113 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node13116 = (inp[14]) ? node13122 : node13117;
														assign node13117 = (inp[6]) ? 16'b0000000011111111 : node13118;
															assign node13118 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node13122 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node13125 = (inp[4]) ? node13143 : node13126;
											assign node13126 = (inp[14]) ? node13134 : node13127;
												assign node13127 = (inp[8]) ? node13129 : 16'b0000001111111111;
													assign node13129 = (inp[15]) ? node13131 : 16'b0000001111111111;
														assign node13131 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node13134 = (inp[8]) ? node13136 : 16'b0000000111111111;
													assign node13136 = (inp[13]) ? 16'b0000000001111111 : node13137;
														assign node13137 = (inp[3]) ? 16'b0000000011111111 : node13138;
															assign node13138 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node13143 = (inp[6]) ? node13149 : node13144;
												assign node13144 = (inp[13]) ? node13146 : 16'b0000000111111111;
													assign node13146 = (inp[15]) ? 16'b0000000111111111 : 16'b0000000011111111;
												assign node13149 = (inp[14]) ? node13157 : node13150;
													assign node13150 = (inp[8]) ? 16'b0000000011111111 : node13151;
														assign node13151 = (inp[3]) ? 16'b0000000011111111 : node13152;
															assign node13152 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node13157 = (inp[8]) ? 16'b0000000001111111 : node13158;
														assign node13158 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node13162 = (inp[6]) ? node13216 : node13163;
										assign node13163 = (inp[15]) ? node13185 : node13164;
											assign node13164 = (inp[14]) ? node13174 : node13165;
												assign node13165 = (inp[8]) ? 16'b0000000111111111 : node13166;
													assign node13166 = (inp[3]) ? node13168 : 16'b0000001111111111;
														assign node13168 = (inp[4]) ? 16'b0000000111111111 : node13169;
															assign node13169 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node13174 = (inp[13]) ? node13180 : node13175;
													assign node13175 = (inp[5]) ? 16'b0000000111111111 : node13176;
														assign node13176 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node13180 = (inp[5]) ? node13182 : 16'b0000000111111111;
														assign node13182 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node13185 = (inp[3]) ? node13203 : node13186;
												assign node13186 = (inp[14]) ? node13194 : node13187;
													assign node13187 = (inp[4]) ? node13189 : 16'b0000000111111111;
														assign node13189 = (inp[5]) ? node13191 : 16'b0000000111111111;
															assign node13191 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node13194 = (inp[13]) ? node13198 : node13195;
														assign node13195 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node13198 = (inp[4]) ? node13200 : 16'b0000000011111111;
															assign node13200 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node13203 = (inp[5]) ? node13209 : node13204;
													assign node13204 = (inp[4]) ? 16'b0000000011111111 : node13205;
														assign node13205 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node13209 = (inp[4]) ? node13211 : 16'b0000000011111111;
														assign node13211 = (inp[8]) ? node13213 : 16'b0000000001111111;
															assign node13213 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node13216 = (inp[5]) ? node13238 : node13217;
											assign node13217 = (inp[13]) ? node13227 : node13218;
												assign node13218 = (inp[14]) ? node13222 : node13219;
													assign node13219 = (inp[4]) ? 16'b0000000111111111 : 16'b0000011111111111;
													assign node13222 = (inp[8]) ? node13224 : 16'b0000000011111111;
														assign node13224 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node13227 = (inp[4]) ? node13233 : node13228;
													assign node13228 = (inp[8]) ? node13230 : 16'b0000000111111111;
														assign node13230 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node13233 = (inp[15]) ? node13235 : 16'b0000000001111111;
														assign node13235 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node13238 = (inp[14]) ? node13246 : node13239;
												assign node13239 = (inp[8]) ? 16'b0000000001111111 : node13240;
													assign node13240 = (inp[4]) ? 16'b0000000001111111 : node13241;
														assign node13241 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node13246 = (inp[13]) ? node13256 : node13247;
													assign node13247 = (inp[15]) ? node13253 : node13248;
														assign node13248 = (inp[3]) ? 16'b0000000001111111 : node13249;
															assign node13249 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node13253 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node13256 = (inp[8]) ? node13258 : 16'b0000000000111111;
														assign node13258 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
								assign node13261 = (inp[15]) ? node13357 : node13262;
									assign node13262 = (inp[14]) ? node13298 : node13263;
										assign node13263 = (inp[4]) ? node13279 : node13264;
											assign node13264 = (inp[1]) ? node13268 : node13265;
												assign node13265 = (inp[6]) ? 16'b0000000111111111 : 16'b0000011111111111;
												assign node13268 = (inp[3]) ? node13270 : 16'b0000000111111111;
													assign node13270 = (inp[8]) ? 16'b0000000011111111 : node13271;
														assign node13271 = (inp[13]) ? 16'b0000000011111111 : node13272;
															assign node13272 = (inp[5]) ? 16'b0000000111111111 : node13273;
																assign node13273 = (inp[6]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node13279 = (inp[13]) ? node13287 : node13280;
												assign node13280 = (inp[1]) ? node13282 : 16'b0000000111111111;
													assign node13282 = (inp[6]) ? node13284 : 16'b0000000111111111;
														assign node13284 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node13287 = (inp[3]) ? node13295 : node13288;
													assign node13288 = (inp[8]) ? 16'b0000000011111111 : node13289;
														assign node13289 = (inp[6]) ? 16'b0000000011111111 : node13290;
															assign node13290 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node13295 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node13298 = (inp[8]) ? node13328 : node13299;
											assign node13299 = (inp[4]) ? node13319 : node13300;
												assign node13300 = (inp[13]) ? node13310 : node13301;
													assign node13301 = (inp[3]) ? node13305 : node13302;
														assign node13302 = (inp[6]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node13305 = (inp[6]) ? 16'b0000000011111111 : node13306;
															assign node13306 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node13310 = (inp[6]) ? node13316 : node13311;
														assign node13311 = (inp[1]) ? 16'b0000000011111111 : node13312;
															assign node13312 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node13316 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node13319 = (inp[1]) ? node13321 : 16'b0000000011111111;
													assign node13321 = (inp[3]) ? node13325 : node13322;
														assign node13322 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node13325 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node13328 = (inp[13]) ? node13342 : node13329;
												assign node13329 = (inp[6]) ? 16'b0000000000111111 : node13330;
													assign node13330 = (inp[3]) ? node13334 : node13331;
														assign node13331 = (inp[4]) ? 16'b0000000011111111 : 16'b0000001111111111;
														assign node13334 = (inp[5]) ? node13336 : 16'b0000000011111111;
															assign node13336 = (inp[1]) ? 16'b0000000001111111 : node13337;
																assign node13337 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node13342 = (inp[1]) ? node13348 : node13343;
													assign node13343 = (inp[6]) ? 16'b0000000001111111 : node13344;
														assign node13344 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node13348 = (inp[5]) ? node13352 : node13349;
														assign node13349 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node13352 = (inp[4]) ? node13354 : 16'b0000000000111111;
															assign node13354 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node13357 = (inp[14]) ? node13407 : node13358;
										assign node13358 = (inp[4]) ? node13382 : node13359;
											assign node13359 = (inp[8]) ? node13371 : node13360;
												assign node13360 = (inp[1]) ? 16'b0000000011111111 : node13361;
													assign node13361 = (inp[3]) ? 16'b0000000011111111 : node13362;
														assign node13362 = (inp[6]) ? node13364 : 16'b0000001111111111;
															assign node13364 = (inp[13]) ? 16'b0000000111111111 : node13365;
																assign node13365 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node13371 = (inp[5]) ? node13377 : node13372;
													assign node13372 = (inp[3]) ? 16'b0000000011111111 : node13373;
														assign node13373 = (inp[13]) ? 16'b0000000011111111 : 16'b0000001111111111;
													assign node13377 = (inp[1]) ? node13379 : 16'b0000000001111111;
														assign node13379 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000011111111;
											assign node13382 = (inp[6]) ? node13394 : node13383;
												assign node13383 = (inp[1]) ? node13389 : node13384;
													assign node13384 = (inp[8]) ? node13386 : 16'b0000000111111111;
														assign node13386 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node13389 = (inp[13]) ? 16'b0000000001111111 : node13390;
														assign node13390 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node13394 = (inp[8]) ? node13402 : node13395;
													assign node13395 = (inp[3]) ? node13397 : 16'b0000000001111111;
														assign node13397 = (inp[13]) ? node13399 : 16'b0000000001111111;
															assign node13399 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node13402 = (inp[5]) ? 16'b0000000000011111 : node13403;
														assign node13403 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node13407 = (inp[8]) ? node13439 : node13408;
											assign node13408 = (inp[4]) ? node13422 : node13409;
												assign node13409 = (inp[5]) ? node13413 : node13410;
													assign node13410 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000111111111;
													assign node13413 = (inp[13]) ? node13415 : 16'b0000000011111111;
														assign node13415 = (inp[6]) ? 16'b0000000001111111 : node13416;
															assign node13416 = (inp[1]) ? 16'b0000000001111111 : node13417;
																assign node13417 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node13422 = (inp[1]) ? node13432 : node13423;
													assign node13423 = (inp[5]) ? node13425 : 16'b0000000001111111;
														assign node13425 = (inp[6]) ? 16'b0000000000111111 : node13426;
															assign node13426 = (inp[13]) ? node13428 : 16'b0000000001111111;
																assign node13428 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node13432 = (inp[13]) ? node13436 : node13433;
														assign node13433 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node13436 = (inp[6]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node13439 = (inp[1]) ? node13447 : node13440;
												assign node13440 = (inp[4]) ? 16'b0000000000111111 : node13441;
													assign node13441 = (inp[6]) ? node13443 : 16'b0000000001111111;
														assign node13443 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node13447 = (inp[6]) ? node13461 : node13448;
													assign node13448 = (inp[3]) ? node13450 : 16'b0000000000111111;
														assign node13450 = (inp[5]) ? node13456 : node13451;
															assign node13451 = (inp[4]) ? node13453 : 16'b0000000000111111;
																assign node13453 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
															assign node13456 = (inp[13]) ? node13458 : 16'b0000000000011111;
																assign node13458 = (inp[4]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node13461 = (inp[4]) ? 16'b0000000000001111 : 16'b0000000000011111;
					assign node13464 = (inp[2]) ? node14262 : node13465;
						assign node13465 = (inp[6]) ? node13867 : node13466;
							assign node13466 = (inp[11]) ? node13660 : node13467;
								assign node13467 = (inp[5]) ? node13583 : node13468;
									assign node13468 = (inp[13]) ? node13530 : node13469;
										assign node13469 = (inp[15]) ? node13509 : node13470;
											assign node13470 = (inp[1]) ? node13490 : node13471;
												assign node13471 = (inp[14]) ? node13483 : node13472;
													assign node13472 = (inp[3]) ? node13478 : node13473;
														assign node13473 = (inp[10]) ? 16'b0000111111111111 : node13474;
															assign node13474 = (inp[4]) ? 16'b0001111111111111 : 16'b0011111111111111;
														assign node13478 = (inp[10]) ? 16'b0000011111111111 : node13479;
															assign node13479 = (inp[4]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node13483 = (inp[10]) ? 16'b0000001111111111 : node13484;
														assign node13484 = (inp[3]) ? 16'b0000001111111111 : node13485;
															assign node13485 = (inp[4]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node13490 = (inp[4]) ? node13500 : node13491;
													assign node13491 = (inp[8]) ? node13495 : node13492;
														assign node13492 = (inp[14]) ? 16'b0000111111111111 : 16'b0000011111111111;
														assign node13495 = (inp[3]) ? node13497 : 16'b0000011111111111;
															assign node13497 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node13500 = (inp[3]) ? node13506 : node13501;
														assign node13501 = (inp[10]) ? 16'b0000001111111111 : node13502;
															assign node13502 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node13506 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node13509 = (inp[3]) ? node13521 : node13510;
												assign node13510 = (inp[14]) ? node13518 : node13511;
													assign node13511 = (inp[4]) ? node13515 : node13512;
														assign node13512 = (inp[1]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node13515 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node13518 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node13521 = (inp[4]) ? 16'b0000000111111111 : node13522;
													assign node13522 = (inp[10]) ? node13524 : 16'b0000001111111111;
														assign node13524 = (inp[14]) ? 16'b0000000111111111 : node13525;
															assign node13525 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node13530 = (inp[14]) ? node13558 : node13531;
											assign node13531 = (inp[10]) ? node13545 : node13532;
												assign node13532 = (inp[1]) ? node13540 : node13533;
													assign node13533 = (inp[4]) ? node13535 : 16'b0000111111111111;
														assign node13535 = (inp[3]) ? node13537 : 16'b0000011111111111;
															assign node13537 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node13540 = (inp[4]) ? 16'b0000000111111111 : node13541;
														assign node13541 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node13545 = (inp[8]) ? 16'b0000000111111111 : node13546;
													assign node13546 = (inp[15]) ? node13550 : node13547;
														assign node13547 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node13550 = (inp[1]) ? node13552 : 16'b0000001111111111;
															assign node13552 = (inp[4]) ? node13554 : 16'b0000000111111111;
																assign node13554 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node13558 = (inp[3]) ? node13566 : node13559;
												assign node13559 = (inp[1]) ? 16'b0000000111111111 : node13560;
													assign node13560 = (inp[10]) ? 16'b0000000111111111 : node13561;
														assign node13561 = (inp[4]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node13566 = (inp[10]) ? node13576 : node13567;
													assign node13567 = (inp[1]) ? node13571 : node13568;
														assign node13568 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node13571 = (inp[8]) ? node13573 : 16'b0000000111111111;
															assign node13573 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node13576 = (inp[15]) ? node13580 : node13577;
														assign node13577 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node13580 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000011111111;
									assign node13583 = (inp[10]) ? node13615 : node13584;
										assign node13584 = (inp[15]) ? node13600 : node13585;
											assign node13585 = (inp[4]) ? node13597 : node13586;
												assign node13586 = (inp[8]) ? node13594 : node13587;
													assign node13587 = (inp[13]) ? 16'b0000011111111111 : node13588;
														assign node13588 = (inp[1]) ? 16'b0000011111111111 : node13589;
															assign node13589 = (inp[14]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node13594 = (inp[3]) ? 16'b0000000111111111 : 16'b0000011111111111;
												assign node13597 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node13600 = (inp[8]) ? node13608 : node13601;
												assign node13601 = (inp[1]) ? node13603 : 16'b0000001111111111;
													assign node13603 = (inp[14]) ? 16'b0000000111111111 : node13604;
														assign node13604 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node13608 = (inp[4]) ? node13612 : node13609;
													assign node13609 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node13612 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node13615 = (inp[14]) ? node13643 : node13616;
											assign node13616 = (inp[1]) ? node13628 : node13617;
												assign node13617 = (inp[13]) ? 16'b0000000111111111 : node13618;
													assign node13618 = (inp[8]) ? node13620 : 16'b0000001111111111;
														assign node13620 = (inp[4]) ? node13622 : 16'b0000001111111111;
															assign node13622 = (inp[3]) ? node13624 : 16'b0000000111111111;
																assign node13624 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node13628 = (inp[13]) ? node13638 : node13629;
													assign node13629 = (inp[3]) ? node13635 : node13630;
														assign node13630 = (inp[15]) ? 16'b0000000111111111 : node13631;
															assign node13631 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node13635 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node13638 = (inp[8]) ? 16'b0000000011111111 : node13639;
														assign node13639 = (inp[4]) ? 16'b0000000011111111 : 16'b0000001111111111;
											assign node13643 = (inp[15]) ? node13649 : node13644;
												assign node13644 = (inp[4]) ? 16'b0000000011111111 : node13645;
													assign node13645 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node13649 = (inp[8]) ? node13655 : node13650;
													assign node13650 = (inp[13]) ? node13652 : 16'b0000000011111111;
														assign node13652 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000001111111;
													assign node13655 = (inp[3]) ? node13657 : 16'b0000000001111111;
														assign node13657 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
								assign node13660 = (inp[4]) ? node13762 : node13661;
									assign node13661 = (inp[1]) ? node13709 : node13662;
										assign node13662 = (inp[8]) ? node13686 : node13663;
											assign node13663 = (inp[13]) ? node13679 : node13664;
												assign node13664 = (inp[5]) ? node13674 : node13665;
													assign node13665 = (inp[3]) ? node13669 : node13666;
														assign node13666 = (inp[15]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node13669 = (inp[14]) ? node13671 : 16'b0000011111111111;
															assign node13671 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node13674 = (inp[3]) ? 16'b0000001111111111 : node13675;
														assign node13675 = (inp[15]) ? 16'b0000000111111111 : 16'b0000011111111111;
												assign node13679 = (inp[10]) ? node13683 : node13680;
													assign node13680 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node13683 = (inp[15]) ? 16'b0000000111111111 : 16'b0000000011111111;
											assign node13686 = (inp[10]) ? node13702 : node13687;
												assign node13687 = (inp[15]) ? node13695 : node13688;
													assign node13688 = (inp[3]) ? node13692 : node13689;
														assign node13689 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node13692 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node13695 = (inp[3]) ? node13699 : node13696;
														assign node13696 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node13699 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node13702 = (inp[3]) ? node13704 : 16'b0000000111111111;
													assign node13704 = (inp[14]) ? 16'b0000000001111111 : node13705;
														assign node13705 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node13709 = (inp[10]) ? node13741 : node13710;
											assign node13710 = (inp[8]) ? node13728 : node13711;
												assign node13711 = (inp[3]) ? node13717 : node13712;
													assign node13712 = (inp[13]) ? 16'b0000000111111111 : node13713;
														assign node13713 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node13717 = (inp[5]) ? node13725 : node13718;
														assign node13718 = (inp[14]) ? node13720 : 16'b0000001111111111;
															assign node13720 = (inp[15]) ? 16'b0000000111111111 : node13721;
																assign node13721 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node13725 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node13728 = (inp[15]) ? node13736 : node13729;
													assign node13729 = (inp[14]) ? node13731 : 16'b0000001111111111;
														assign node13731 = (inp[3]) ? node13733 : 16'b0000000111111111;
															assign node13733 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node13736 = (inp[13]) ? node13738 : 16'b0000000011111111;
														assign node13738 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node13741 = (inp[15]) ? node13751 : node13742;
												assign node13742 = (inp[13]) ? 16'b0000000001111111 : node13743;
													assign node13743 = (inp[14]) ? node13747 : node13744;
														assign node13744 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node13747 = (inp[8]) ? 16'b0000000111111111 : 16'b0000000011111111;
												assign node13751 = (inp[14]) ? node13753 : 16'b0000000011111111;
													assign node13753 = (inp[3]) ? node13757 : node13754;
														assign node13754 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node13757 = (inp[8]) ? node13759 : 16'b0000000001111111;
															assign node13759 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node13762 = (inp[8]) ? node13808 : node13763;
										assign node13763 = (inp[15]) ? node13787 : node13764;
											assign node13764 = (inp[1]) ? node13776 : node13765;
												assign node13765 = (inp[3]) ? 16'b0000000111111111 : node13766;
													assign node13766 = (inp[5]) ? node13768 : 16'b0000001111111111;
														assign node13768 = (inp[10]) ? node13772 : node13769;
															assign node13769 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
															assign node13772 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node13776 = (inp[14]) ? node13782 : node13777;
													assign node13777 = (inp[13]) ? node13779 : 16'b0000000111111111;
														assign node13779 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node13782 = (inp[13]) ? 16'b0000000011111111 : node13783;
														assign node13783 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node13787 = (inp[10]) ? node13801 : node13788;
												assign node13788 = (inp[3]) ? node13794 : node13789;
													assign node13789 = (inp[5]) ? 16'b0000000011111111 : node13790;
														assign node13790 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node13794 = (inp[14]) ? node13798 : node13795;
														assign node13795 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node13798 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node13801 = (inp[3]) ? node13803 : 16'b0000000011111111;
													assign node13803 = (inp[13]) ? node13805 : 16'b0000000001111111;
														assign node13805 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node13808 = (inp[10]) ? node13838 : node13809;
											assign node13809 = (inp[15]) ? node13821 : node13810;
												assign node13810 = (inp[5]) ? node13816 : node13811;
													assign node13811 = (inp[13]) ? node13813 : 16'b0000000111111111;
														assign node13813 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node13816 = (inp[13]) ? 16'b0000000011111111 : node13817;
														assign node13817 = (inp[1]) ? 16'b0000000011111111 : 16'b0000001111111111;
												assign node13821 = (inp[1]) ? node13833 : node13822;
													assign node13822 = (inp[3]) ? node13826 : node13823;
														assign node13823 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node13826 = (inp[14]) ? node13828 : 16'b0000000011111111;
															assign node13828 = (inp[13]) ? 16'b0000000001111111 : node13829;
																assign node13829 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node13833 = (inp[3]) ? 16'b0000000001111111 : node13834;
														assign node13834 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node13838 = (inp[13]) ? node13852 : node13839;
												assign node13839 = (inp[5]) ? node13845 : node13840;
													assign node13840 = (inp[15]) ? node13842 : 16'b0000000011111111;
														assign node13842 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node13845 = (inp[3]) ? node13849 : node13846;
														assign node13846 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000111111111;
														assign node13849 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node13852 = (inp[15]) ? node13860 : node13853;
													assign node13853 = (inp[3]) ? 16'b0000000000111111 : node13854;
														assign node13854 = (inp[5]) ? node13856 : 16'b0000000001111111;
															assign node13856 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node13860 = (inp[1]) ? node13862 : 16'b0000000000111111;
														assign node13862 = (inp[5]) ? node13864 : 16'b0000000000011111;
															assign node13864 = (inp[14]) ? 16'b0000000000001111 : 16'b0000000000011111;
							assign node13867 = (inp[14]) ? node14067 : node13868;
								assign node13868 = (inp[13]) ? node13980 : node13869;
									assign node13869 = (inp[15]) ? node13929 : node13870;
										assign node13870 = (inp[11]) ? node13906 : node13871;
											assign node13871 = (inp[1]) ? node13893 : node13872;
												assign node13872 = (inp[5]) ? node13882 : node13873;
													assign node13873 = (inp[3]) ? 16'b0000011111111111 : node13874;
														assign node13874 = (inp[10]) ? node13878 : node13875;
															assign node13875 = (inp[4]) ? 16'b0000111111111111 : 16'b0001111111111111;
															assign node13878 = (inp[4]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node13882 = (inp[4]) ? node13890 : node13883;
														assign node13883 = (inp[8]) ? node13885 : 16'b0000011111111111;
															assign node13885 = (inp[3]) ? 16'b0000001111111111 : node13886;
																assign node13886 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node13890 = (inp[10]) ? 16'b0000001111111111 : 16'b0000000111111111;
												assign node13893 = (inp[3]) ? node13899 : node13894;
													assign node13894 = (inp[8]) ? 16'b0000001111111111 : node13895;
														assign node13895 = (inp[4]) ? 16'b0000011111111111 : 16'b0000001111111111;
													assign node13899 = (inp[4]) ? node13903 : node13900;
														assign node13900 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node13903 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node13906 = (inp[5]) ? node13918 : node13907;
												assign node13907 = (inp[8]) ? node13915 : node13908;
													assign node13908 = (inp[4]) ? node13912 : node13909;
														assign node13909 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node13912 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node13915 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node13918 = (inp[1]) ? node13922 : node13919;
													assign node13919 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node13922 = (inp[4]) ? 16'b0000000011111111 : node13923;
														assign node13923 = (inp[8]) ? node13925 : 16'b0000000011111111;
															assign node13925 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node13929 = (inp[8]) ? node13947 : node13930;
											assign node13930 = (inp[1]) ? node13940 : node13931;
												assign node13931 = (inp[11]) ? node13933 : 16'b0000001111111111;
													assign node13933 = (inp[4]) ? node13937 : node13934;
														assign node13934 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node13937 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node13940 = (inp[11]) ? node13942 : 16'b0000000111111111;
													assign node13942 = (inp[4]) ? 16'b0000000011111111 : node13943;
														assign node13943 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node13947 = (inp[1]) ? node13967 : node13948;
												assign node13948 = (inp[4]) ? node13958 : node13949;
													assign node13949 = (inp[10]) ? node13951 : 16'b0000001111111111;
														assign node13951 = (inp[5]) ? 16'b0000000111111111 : node13952;
															assign node13952 = (inp[11]) ? 16'b0000000111111111 : node13953;
																assign node13953 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node13958 = (inp[10]) ? 16'b0000000001111111 : node13959;
														assign node13959 = (inp[3]) ? node13961 : 16'b0000000011111111;
															assign node13961 = (inp[5]) ? node13963 : 16'b0000000011111111;
																assign node13963 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node13967 = (inp[5]) ? node13975 : node13968;
													assign node13968 = (inp[11]) ? 16'b0000000001111111 : node13969;
														assign node13969 = (inp[4]) ? node13971 : 16'b0000000011111111;
															assign node13971 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node13975 = (inp[11]) ? node13977 : 16'b0000000001111111;
														assign node13977 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000001111111;
									assign node13980 = (inp[3]) ? node14028 : node13981;
										assign node13981 = (inp[5]) ? node14005 : node13982;
											assign node13982 = (inp[10]) ? node13996 : node13983;
												assign node13983 = (inp[11]) ? node13991 : node13984;
													assign node13984 = (inp[15]) ? 16'b0000001111111111 : node13985;
														assign node13985 = (inp[8]) ? 16'b0000001111111111 : node13986;
															assign node13986 = (inp[4]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node13991 = (inp[1]) ? node13993 : 16'b0000001111111111;
														assign node13993 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node13996 = (inp[11]) ? node14000 : node13997;
													assign node13997 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node14000 = (inp[1]) ? 16'b0000000011111111 : node14001;
														assign node14001 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node14005 = (inp[1]) ? node14009 : node14006;
												assign node14006 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node14009 = (inp[15]) ? node14021 : node14010;
													assign node14010 = (inp[11]) ? node14014 : node14011;
														assign node14011 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node14014 = (inp[8]) ? 16'b0000000001111111 : node14015;
															assign node14015 = (inp[10]) ? node14017 : 16'b0000000011111111;
																assign node14017 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node14021 = (inp[10]) ? node14025 : node14022;
														assign node14022 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node14025 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node14028 = (inp[4]) ? node14046 : node14029;
											assign node14029 = (inp[10]) ? node14039 : node14030;
												assign node14030 = (inp[5]) ? 16'b0000000011111111 : node14031;
													assign node14031 = (inp[15]) ? node14033 : 16'b0000000111111111;
														assign node14033 = (inp[8]) ? 16'b0000000011111111 : node14034;
															assign node14034 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node14039 = (inp[11]) ? node14041 : 16'b0000000011111111;
													assign node14041 = (inp[8]) ? node14043 : 16'b0000000001111111;
														assign node14043 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node14046 = (inp[1]) ? node14054 : node14047;
												assign node14047 = (inp[11]) ? 16'b0000000001111111 : node14048;
													assign node14048 = (inp[8]) ? 16'b0000000001111111 : node14049;
														assign node14049 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node14054 = (inp[10]) ? node14062 : node14055;
													assign node14055 = (inp[15]) ? node14059 : node14056;
														assign node14056 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node14059 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node14062 = (inp[15]) ? 16'b0000000000111111 : node14063;
														assign node14063 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
								assign node14067 = (inp[10]) ? node14155 : node14068;
									assign node14068 = (inp[3]) ? node14116 : node14069;
										assign node14069 = (inp[4]) ? node14081 : node14070;
											assign node14070 = (inp[13]) ? node14076 : node14071;
												assign node14071 = (inp[1]) ? node14073 : 16'b0000001111111111;
													assign node14073 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node14076 = (inp[8]) ? 16'b0000000011111111 : node14077;
													assign node14077 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node14081 = (inp[13]) ? node14103 : node14082;
												assign node14082 = (inp[15]) ? node14094 : node14083;
													assign node14083 = (inp[11]) ? node14091 : node14084;
														assign node14084 = (inp[8]) ? 16'b0000000011111111 : node14085;
															assign node14085 = (inp[5]) ? node14087 : 16'b0000001111111111;
																assign node14087 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node14091 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node14094 = (inp[5]) ? node14096 : 16'b0000000111111111;
														assign node14096 = (inp[11]) ? node14098 : 16'b0000000011111111;
															assign node14098 = (inp[1]) ? node14100 : 16'b0000000011111111;
																assign node14100 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node14103 = (inp[15]) ? node14107 : node14104;
													assign node14104 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node14107 = (inp[8]) ? node14111 : node14108;
														assign node14108 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node14111 = (inp[1]) ? node14113 : 16'b0000000001111111;
															assign node14113 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node14116 = (inp[11]) ? node14132 : node14117;
											assign node14117 = (inp[1]) ? node14121 : node14118;
												assign node14118 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node14121 = (inp[8]) ? 16'b0000000001111111 : node14122;
													assign node14122 = (inp[5]) ? node14126 : node14123;
														assign node14123 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node14126 = (inp[15]) ? node14128 : 16'b0000000011111111;
															assign node14128 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node14132 = (inp[8]) ? node14148 : node14133;
												assign node14133 = (inp[13]) ? node14141 : node14134;
													assign node14134 = (inp[15]) ? 16'b0000000001111111 : node14135;
														assign node14135 = (inp[5]) ? 16'b0000000001111111 : node14136;
															assign node14136 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node14141 = (inp[4]) ? node14143 : 16'b0000000001111111;
														assign node14143 = (inp[5]) ? 16'b0000000000111111 : node14144;
															assign node14144 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node14148 = (inp[5]) ? 16'b0000000000111111 : node14149;
													assign node14149 = (inp[1]) ? node14151 : 16'b0000000000111111;
														assign node14151 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node14155 = (inp[4]) ? node14213 : node14156;
										assign node14156 = (inp[1]) ? node14182 : node14157;
											assign node14157 = (inp[11]) ? node14169 : node14158;
												assign node14158 = (inp[13]) ? node14162 : node14159;
													assign node14159 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node14162 = (inp[5]) ? 16'b0000000001111111 : node14163;
														assign node14163 = (inp[8]) ? 16'b0000000011111111 : node14164;
															assign node14164 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node14169 = (inp[8]) ? node14175 : node14170;
													assign node14170 = (inp[13]) ? node14172 : 16'b0000000011111111;
														assign node14172 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000011111111;
													assign node14175 = (inp[5]) ? node14177 : 16'b0000000001111111;
														assign node14177 = (inp[13]) ? 16'b0000000001111111 : node14178;
															assign node14178 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node14182 = (inp[5]) ? node14200 : node14183;
												assign node14183 = (inp[3]) ? node14189 : node14184;
													assign node14184 = (inp[13]) ? node14186 : 16'b0000000011111111;
														assign node14186 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node14189 = (inp[8]) ? node14195 : node14190;
														assign node14190 = (inp[13]) ? 16'b0000000001111111 : node14191;
															assign node14191 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node14195 = (inp[13]) ? 16'b0000000000011111 : node14196;
															assign node14196 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node14200 = (inp[11]) ? node14208 : node14201;
													assign node14201 = (inp[15]) ? node14203 : 16'b0000000001111111;
														assign node14203 = (inp[3]) ? 16'b0000000000111111 : node14204;
															assign node14204 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node14208 = (inp[8]) ? node14210 : 16'b0000000000111111;
														assign node14210 = (inp[15]) ? 16'b0000000000001111 : 16'b0000000000011111;
										assign node14213 = (inp[15]) ? node14233 : node14214;
											assign node14214 = (inp[3]) ? node14220 : node14215;
												assign node14215 = (inp[5]) ? 16'b0000000001111111 : node14216;
													assign node14216 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node14220 = (inp[1]) ? node14222 : 16'b0000000001111111;
													assign node14222 = (inp[11]) ? node14228 : node14223;
														assign node14223 = (inp[5]) ? 16'b0000000000111111 : node14224;
															assign node14224 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node14228 = (inp[13]) ? node14230 : 16'b0000000000111111;
															assign node14230 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node14233 = (inp[13]) ? node14249 : node14234;
												assign node14234 = (inp[5]) ? node14242 : node14235;
													assign node14235 = (inp[1]) ? node14239 : node14236;
														assign node14236 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node14239 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node14242 = (inp[3]) ? node14246 : node14243;
														assign node14243 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node14246 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node14249 = (inp[5]) ? node14255 : node14250;
													assign node14250 = (inp[3]) ? node14252 : 16'b0000000000111111;
														assign node14252 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node14255 = (inp[1]) ? node14259 : node14256;
														assign node14256 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node14259 = (inp[3]) ? 16'b0000000000001111 : 16'b0000000000011111;
						assign node14262 = (inp[1]) ? node14648 : node14263;
							assign node14263 = (inp[5]) ? node14465 : node14264;
								assign node14264 = (inp[4]) ? node14372 : node14265;
									assign node14265 = (inp[6]) ? node14325 : node14266;
										assign node14266 = (inp[13]) ? node14292 : node14267;
											assign node14267 = (inp[14]) ? node14281 : node14268;
												assign node14268 = (inp[3]) ? 16'b0000001111111111 : node14269;
													assign node14269 = (inp[15]) ? node14277 : node14270;
														assign node14270 = (inp[10]) ? 16'b0000011111111111 : node14271;
															assign node14271 = (inp[8]) ? 16'b0000111111111111 : node14272;
																assign node14272 = (inp[11]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node14277 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node14281 = (inp[15]) ? node14287 : node14282;
													assign node14282 = (inp[10]) ? 16'b0000001111111111 : node14283;
														assign node14283 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node14287 = (inp[3]) ? 16'b0000000001111111 : node14288;
														assign node14288 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node14292 = (inp[14]) ? node14310 : node14293;
												assign node14293 = (inp[3]) ? node14307 : node14294;
													assign node14294 = (inp[10]) ? node14300 : node14295;
														assign node14295 = (inp[8]) ? 16'b0000001111111111 : node14296;
															assign node14296 = (inp[11]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node14300 = (inp[11]) ? node14302 : 16'b0000001111111111;
															assign node14302 = (inp[15]) ? 16'b0000000111111111 : node14303;
																assign node14303 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node14307 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node14310 = (inp[11]) ? node14318 : node14311;
													assign node14311 = (inp[8]) ? node14315 : node14312;
														assign node14312 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node14315 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node14318 = (inp[10]) ? 16'b0000000001111111 : node14319;
														assign node14319 = (inp[3]) ? 16'b0000000011111111 : node14320;
															assign node14320 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node14325 = (inp[15]) ? node14343 : node14326;
											assign node14326 = (inp[13]) ? node14334 : node14327;
												assign node14327 = (inp[10]) ? 16'b0000000111111111 : node14328;
													assign node14328 = (inp[14]) ? 16'b0000001111111111 : node14329;
														assign node14329 = (inp[3]) ? 16'b0000011111111111 : 16'b0000001111111111;
												assign node14334 = (inp[11]) ? node14338 : node14335;
													assign node14335 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node14338 = (inp[8]) ? node14340 : 16'b0000000001111111;
														assign node14340 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node14343 = (inp[11]) ? node14359 : node14344;
												assign node14344 = (inp[8]) ? node14356 : node14345;
													assign node14345 = (inp[14]) ? node14349 : node14346;
														assign node14346 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node14349 = (inp[3]) ? 16'b0000000011111111 : node14350;
															assign node14350 = (inp[13]) ? node14352 : 16'b0000000111111111;
																assign node14352 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node14356 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node14359 = (inp[14]) ? node14367 : node14360;
													assign node14360 = (inp[3]) ? node14364 : node14361;
														assign node14361 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node14364 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node14367 = (inp[13]) ? 16'b0000000000111111 : node14368;
														assign node14368 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node14372 = (inp[15]) ? node14412 : node14373;
										assign node14373 = (inp[14]) ? node14393 : node14374;
											assign node14374 = (inp[6]) ? node14384 : node14375;
												assign node14375 = (inp[13]) ? node14381 : node14376;
													assign node14376 = (inp[3]) ? 16'b0000001111111111 : node14377;
														assign node14377 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node14381 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node14384 = (inp[11]) ? node14386 : 16'b0000000111111111;
													assign node14386 = (inp[13]) ? 16'b0000000011111111 : node14387;
														assign node14387 = (inp[3]) ? 16'b0000000011111111 : node14388;
															assign node14388 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node14393 = (inp[6]) ? node14403 : node14394;
												assign node14394 = (inp[10]) ? 16'b0000000011111111 : node14395;
													assign node14395 = (inp[11]) ? 16'b0000000011111111 : node14396;
														assign node14396 = (inp[8]) ? 16'b0000000111111111 : node14397;
															assign node14397 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node14403 = (inp[8]) ? node14405 : 16'b0000000011111111;
													assign node14405 = (inp[3]) ? node14407 : 16'b0000000011111111;
														assign node14407 = (inp[13]) ? node14409 : 16'b0000000001111111;
															assign node14409 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node14412 = (inp[11]) ? node14436 : node14413;
											assign node14413 = (inp[8]) ? node14419 : node14414;
												assign node14414 = (inp[13]) ? 16'b0000000001111111 : node14415;
													assign node14415 = (inp[6]) ? 16'b0000001111111111 : 16'b0000000111111111;
												assign node14419 = (inp[3]) ? node14431 : node14420;
													assign node14420 = (inp[14]) ? node14428 : node14421;
														assign node14421 = (inp[6]) ? 16'b0000000011111111 : node14422;
															assign node14422 = (inp[10]) ? node14424 : 16'b0000000111111111;
																assign node14424 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node14428 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node14431 = (inp[6]) ? 16'b0000000001111111 : node14432;
														assign node14432 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node14436 = (inp[13]) ? node14446 : node14437;
												assign node14437 = (inp[14]) ? node14443 : node14438;
													assign node14438 = (inp[6]) ? node14440 : 16'b0000000011111111;
														assign node14440 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node14443 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node14446 = (inp[3]) ? node14456 : node14447;
													assign node14447 = (inp[14]) ? node14451 : node14448;
														assign node14448 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node14451 = (inp[6]) ? 16'b0000000000111111 : node14452;
															assign node14452 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node14456 = (inp[10]) ? node14460 : node14457;
														assign node14457 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000000111111;
														assign node14460 = (inp[8]) ? node14462 : 16'b0000000000111111;
															assign node14462 = (inp[6]) ? 16'b0000000000011111 : 16'b0000000000111111;
								assign node14465 = (inp[8]) ? node14555 : node14466;
									assign node14466 = (inp[6]) ? node14514 : node14467;
										assign node14467 = (inp[3]) ? node14487 : node14468;
											assign node14468 = (inp[14]) ? node14476 : node14469;
												assign node14469 = (inp[4]) ? node14473 : node14470;
													assign node14470 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node14473 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node14476 = (inp[15]) ? node14482 : node14477;
													assign node14477 = (inp[13]) ? node14479 : 16'b0000001111111111;
														assign node14479 = (inp[4]) ? 16'b0000000111111111 : 16'b0000000011111111;
													assign node14482 = (inp[4]) ? 16'b0000000011111111 : node14483;
														assign node14483 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node14487 = (inp[4]) ? node14503 : node14488;
												assign node14488 = (inp[10]) ? node14498 : node14489;
													assign node14489 = (inp[13]) ? 16'b0000000011111111 : node14490;
														assign node14490 = (inp[11]) ? 16'b0000000111111111 : node14491;
															assign node14491 = (inp[15]) ? node14493 : 16'b0000001111111111;
																assign node14493 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node14498 = (inp[11]) ? 16'b0000000001111111 : node14499;
														assign node14499 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node14503 = (inp[15]) ? node14505 : 16'b0000000011111111;
													assign node14505 = (inp[10]) ? node14509 : node14506;
														assign node14506 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node14509 = (inp[14]) ? 16'b0000000000111111 : node14510;
															assign node14510 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node14514 = (inp[3]) ? node14536 : node14515;
											assign node14515 = (inp[14]) ? node14527 : node14516;
												assign node14516 = (inp[15]) ? node14522 : node14517;
													assign node14517 = (inp[13]) ? 16'b0000000011111111 : node14518;
														assign node14518 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node14522 = (inp[10]) ? 16'b0000000001111111 : node14523;
														assign node14523 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node14527 = (inp[10]) ? node14533 : node14528;
													assign node14528 = (inp[15]) ? node14530 : 16'b0000000011111111;
														assign node14530 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node14533 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node14536 = (inp[13]) ? node14550 : node14537;
												assign node14537 = (inp[15]) ? node14545 : node14538;
													assign node14538 = (inp[4]) ? 16'b0000000001111111 : node14539;
														assign node14539 = (inp[11]) ? 16'b0000000011111111 : node14540;
															assign node14540 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node14545 = (inp[10]) ? node14547 : 16'b0000000001111111;
														assign node14547 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node14550 = (inp[11]) ? 16'b0000000000111111 : node14551;
													assign node14551 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000000111111;
									assign node14555 = (inp[14]) ? node14609 : node14556;
										assign node14556 = (inp[11]) ? node14588 : node14557;
											assign node14557 = (inp[15]) ? node14577 : node14558;
												assign node14558 = (inp[13]) ? node14570 : node14559;
													assign node14559 = (inp[10]) ? node14563 : node14560;
														assign node14560 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node14563 = (inp[4]) ? node14565 : 16'b0000000111111111;
															assign node14565 = (inp[6]) ? 16'b0000000011111111 : node14566;
																assign node14566 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node14570 = (inp[6]) ? node14572 : 16'b0000000001111111;
														assign node14572 = (inp[4]) ? 16'b0000000011111111 : node14573;
															assign node14573 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node14577 = (inp[10]) ? node14579 : 16'b0000000011111111;
													assign node14579 = (inp[3]) ? 16'b0000000000111111 : node14580;
														assign node14580 = (inp[6]) ? 16'b0000000001111111 : node14581;
															assign node14581 = (inp[13]) ? node14583 : 16'b0000000011111111;
																assign node14583 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node14588 = (inp[15]) ? node14596 : node14589;
												assign node14589 = (inp[3]) ? node14593 : node14590;
													assign node14590 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node14593 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node14596 = (inp[6]) ? node14598 : 16'b0000000001111111;
													assign node14598 = (inp[13]) ? node14606 : node14599;
														assign node14599 = (inp[4]) ? node14601 : 16'b0000000001111111;
															assign node14601 = (inp[10]) ? 16'b0000000000111111 : node14602;
																assign node14602 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node14606 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node14609 = (inp[10]) ? node14631 : node14610;
											assign node14610 = (inp[13]) ? node14614 : node14611;
												assign node14611 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000001111111;
												assign node14614 = (inp[3]) ? node14626 : node14615;
													assign node14615 = (inp[15]) ? node14621 : node14616;
														assign node14616 = (inp[4]) ? node14618 : 16'b0000000011111111;
															assign node14618 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node14621 = (inp[11]) ? 16'b0000000000111111 : node14622;
															assign node14622 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node14626 = (inp[6]) ? 16'b0000000000011111 : node14627;
														assign node14627 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node14631 = (inp[6]) ? node14641 : node14632;
												assign node14632 = (inp[13]) ? node14638 : node14633;
													assign node14633 = (inp[4]) ? node14635 : 16'b0000000001111111;
														assign node14635 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node14638 = (inp[4]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node14641 = (inp[3]) ? node14645 : node14642;
													assign node14642 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node14645 = (inp[4]) ? 16'b0000000000001111 : 16'b0000000000011111;
							assign node14648 = (inp[13]) ? node14818 : node14649;
								assign node14649 = (inp[3]) ? node14729 : node14650;
									assign node14650 = (inp[11]) ? node14682 : node14651;
										assign node14651 = (inp[6]) ? node14663 : node14652;
											assign node14652 = (inp[14]) ? node14660 : node14653;
												assign node14653 = (inp[10]) ? 16'b0000001111111111 : node14654;
													assign node14654 = (inp[8]) ? 16'b0000000111111111 : node14655;
														assign node14655 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node14660 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node14663 = (inp[4]) ? node14673 : node14664;
												assign node14664 = (inp[8]) ? node14666 : 16'b0000000111111111;
													assign node14666 = (inp[5]) ? 16'b0000000011111111 : node14667;
														assign node14667 = (inp[10]) ? node14669 : 16'b0000000111111111;
															assign node14669 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node14673 = (inp[5]) ? node14675 : 16'b0000000111111111;
													assign node14675 = (inp[15]) ? 16'b0000000001111111 : node14676;
														assign node14676 = (inp[14]) ? node14678 : 16'b0000000011111111;
															assign node14678 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node14682 = (inp[14]) ? node14706 : node14683;
											assign node14683 = (inp[4]) ? node14699 : node14684;
												assign node14684 = (inp[15]) ? node14690 : node14685;
													assign node14685 = (inp[5]) ? 16'b0000000111111111 : node14686;
														assign node14686 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node14690 = (inp[10]) ? 16'b0000000011111111 : node14691;
														assign node14691 = (inp[8]) ? 16'b0000000011111111 : node14692;
															assign node14692 = (inp[6]) ? node14694 : 16'b0000000111111111;
																assign node14694 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node14699 = (inp[15]) ? node14703 : node14700;
													assign node14700 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node14703 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node14706 = (inp[10]) ? node14720 : node14707;
												assign node14707 = (inp[5]) ? node14711 : node14708;
													assign node14708 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node14711 = (inp[15]) ? 16'b0000000000111111 : node14712;
														assign node14712 = (inp[8]) ? 16'b0000000001111111 : node14713;
															assign node14713 = (inp[4]) ? node14715 : 16'b0000000011111111;
																assign node14715 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node14720 = (inp[5]) ? 16'b0000000000011111 : node14721;
													assign node14721 = (inp[15]) ? 16'b0000000000111111 : node14722;
														assign node14722 = (inp[6]) ? node14724 : 16'b0000000011111111;
															assign node14724 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node14729 = (inp[15]) ? node14779 : node14730;
										assign node14730 = (inp[6]) ? node14756 : node14731;
											assign node14731 = (inp[5]) ? node14737 : node14732;
												assign node14732 = (inp[4]) ? node14734 : 16'b0000000111111111;
													assign node14734 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node14737 = (inp[10]) ? node14747 : node14738;
													assign node14738 = (inp[4]) ? 16'b0000000011111111 : node14739;
														assign node14739 = (inp[11]) ? node14741 : 16'b0000000111111111;
															assign node14741 = (inp[8]) ? 16'b0000000011111111 : node14742;
																assign node14742 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node14747 = (inp[14]) ? node14753 : node14748;
														assign node14748 = (inp[11]) ? node14750 : 16'b0000000011111111;
															assign node14750 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node14753 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node14756 = (inp[5]) ? node14766 : node14757;
												assign node14757 = (inp[10]) ? node14759 : 16'b0000000011111111;
													assign node14759 = (inp[4]) ? 16'b0000000001111111 : node14760;
														assign node14760 = (inp[14]) ? 16'b0000000001111111 : node14761;
															assign node14761 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node14766 = (inp[4]) ? node14774 : node14767;
													assign node14767 = (inp[11]) ? node14769 : 16'b0000000011111111;
														assign node14769 = (inp[14]) ? node14771 : 16'b0000000001111111;
															assign node14771 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node14774 = (inp[11]) ? 16'b0000000000001111 : node14775;
														assign node14775 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node14779 = (inp[4]) ? node14795 : node14780;
											assign node14780 = (inp[14]) ? node14790 : node14781;
												assign node14781 = (inp[8]) ? node14785 : node14782;
													assign node14782 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node14785 = (inp[10]) ? 16'b0000000000111111 : node14786;
														assign node14786 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node14790 = (inp[6]) ? node14792 : 16'b0000000001111111;
													assign node14792 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000001111111;
											assign node14795 = (inp[6]) ? node14807 : node14796;
												assign node14796 = (inp[8]) ? 16'b0000000000011111 : node14797;
													assign node14797 = (inp[11]) ? node14799 : 16'b0000000011111111;
														assign node14799 = (inp[10]) ? 16'b0000000000111111 : node14800;
															assign node14800 = (inp[5]) ? node14802 : 16'b0000000001111111;
																assign node14802 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node14807 = (inp[10]) ? node14811 : node14808;
													assign node14808 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node14811 = (inp[14]) ? 16'b0000000000001111 : node14812;
														assign node14812 = (inp[8]) ? node14814 : 16'b0000000000011111;
															assign node14814 = (inp[5]) ? 16'b0000000000001111 : 16'b0000000000011111;
								assign node14818 = (inp[11]) ? node14920 : node14819;
									assign node14819 = (inp[3]) ? node14869 : node14820;
										assign node14820 = (inp[8]) ? node14840 : node14821;
											assign node14821 = (inp[14]) ? node14833 : node14822;
												assign node14822 = (inp[4]) ? node14824 : 16'b0000000111111111;
													assign node14824 = (inp[15]) ? node14830 : node14825;
														assign node14825 = (inp[5]) ? node14827 : 16'b0000000111111111;
															assign node14827 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node14830 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node14833 = (inp[5]) ? 16'b0000000001111111 : node14834;
													assign node14834 = (inp[6]) ? node14836 : 16'b0000000011111111;
														assign node14836 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node14840 = (inp[10]) ? node14858 : node14841;
												assign node14841 = (inp[6]) ? node14849 : node14842;
													assign node14842 = (inp[5]) ? node14846 : node14843;
														assign node14843 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node14846 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node14849 = (inp[14]) ? node14855 : node14850;
														assign node14850 = (inp[5]) ? 16'b0000000001111111 : node14851;
															assign node14851 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node14855 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node14858 = (inp[5]) ? node14862 : node14859;
													assign node14859 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node14862 = (inp[4]) ? node14864 : 16'b0000000000011111;
														assign node14864 = (inp[14]) ? node14866 : 16'b0000000000111111;
															assign node14866 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node14869 = (inp[4]) ? node14903 : node14870;
											assign node14870 = (inp[6]) ? node14892 : node14871;
												assign node14871 = (inp[8]) ? node14879 : node14872;
													assign node14872 = (inp[14]) ? node14874 : 16'b0000001111111111;
														assign node14874 = (inp[5]) ? node14876 : 16'b0000000011111111;
															assign node14876 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node14879 = (inp[5]) ? node14885 : node14880;
														assign node14880 = (inp[10]) ? 16'b0000000001111111 : node14881;
															assign node14881 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node14885 = (inp[14]) ? node14887 : 16'b0000000001111111;
															assign node14887 = (inp[10]) ? 16'b0000000000111111 : node14888;
																assign node14888 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node14892 = (inp[14]) ? node14896 : node14893;
													assign node14893 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node14896 = (inp[8]) ? 16'b0000000000011111 : node14897;
														assign node14897 = (inp[15]) ? node14899 : 16'b0000000000111111;
															assign node14899 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node14903 = (inp[15]) ? node14909 : node14904;
												assign node14904 = (inp[6]) ? node14906 : 16'b0000000000111111;
													assign node14906 = (inp[10]) ? 16'b0000000000001111 : 16'b0000000000111111;
												assign node14909 = (inp[14]) ? node14915 : node14910;
													assign node14910 = (inp[6]) ? node14912 : 16'b0000000001111111;
														assign node14912 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node14915 = (inp[6]) ? node14917 : 16'b0000000000011111;
														assign node14917 = (inp[8]) ? 16'b0000000000001111 : 16'b0000000000011111;
									assign node14920 = (inp[4]) ? node14978 : node14921;
										assign node14921 = (inp[14]) ? node14947 : node14922;
											assign node14922 = (inp[15]) ? 16'b0000000000111111 : node14923;
												assign node14923 = (inp[8]) ? node14935 : node14924;
													assign node14924 = (inp[6]) ? node14928 : node14925;
														assign node14925 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node14928 = (inp[5]) ? node14930 : 16'b0000000011111111;
															assign node14930 = (inp[3]) ? 16'b0000000001111111 : node14931;
																assign node14931 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node14935 = (inp[6]) ? node14941 : node14936;
														assign node14936 = (inp[10]) ? 16'b0000000001111111 : node14937;
															assign node14937 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node14941 = (inp[10]) ? 16'b0000000000111111 : node14942;
															assign node14942 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000011111111;
											assign node14947 = (inp[8]) ? node14959 : node14948;
												assign node14948 = (inp[5]) ? 16'b0000000000111111 : node14949;
													assign node14949 = (inp[6]) ? 16'b0000000000111111 : node14950;
														assign node14950 = (inp[15]) ? node14952 : 16'b0000000001111111;
															assign node14952 = (inp[3]) ? node14954 : 16'b0000000001111111;
																assign node14954 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node14959 = (inp[10]) ? node14963 : node14960;
													assign node14960 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node14963 = (inp[3]) ? node14971 : node14964;
														assign node14964 = (inp[15]) ? node14966 : 16'b0000000000011111;
															assign node14966 = (inp[5]) ? node14968 : 16'b0000000000011111;
																assign node14968 = (inp[6]) ? 16'b0000000000001111 : 16'b0000000000011111;
														assign node14971 = (inp[15]) ? node14975 : node14972;
															assign node14972 = (inp[6]) ? 16'b0000000000001111 : 16'b0000000000011111;
															assign node14975 = (inp[6]) ? 16'b0000000000000111 : 16'b0000000000001111;
										assign node14978 = (inp[6]) ? node15000 : node14979;
											assign node14979 = (inp[8]) ? node14985 : node14980;
												assign node14980 = (inp[15]) ? 16'b0000000000111111 : node14981;
													assign node14981 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node14985 = (inp[5]) ? node14993 : node14986;
													assign node14986 = (inp[3]) ? node14990 : node14987;
														assign node14987 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node14990 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000000011111;
													assign node14993 = (inp[15]) ? node14997 : node14994;
														assign node14994 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node14997 = (inp[14]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node15000 = (inp[3]) ? node15012 : node15001;
												assign node15001 = (inp[10]) ? 16'b0000000000011111 : node15002;
													assign node15002 = (inp[8]) ? node15004 : 16'b0000000000111111;
														assign node15004 = (inp[15]) ? 16'b0000000000011111 : node15005;
															assign node15005 = (inp[14]) ? node15007 : 16'b0000000000111111;
																assign node15007 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node15012 = (inp[8]) ? node15022 : node15013;
													assign node15013 = (inp[14]) ? node15019 : node15014;
														assign node15014 = (inp[10]) ? 16'b0000000000011111 : node15015;
															assign node15015 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node15019 = (inp[5]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node15022 = (inp[5]) ? node15024 : 16'b0000000000011111;
														assign node15024 = (inp[15]) ? 16'b0000000000000111 : node15025;
															assign node15025 = (inp[10]) ? node15027 : 16'b0000000000001111;
																assign node15027 = (inp[14]) ? 16'b0000000000000111 : 16'b0000000000001111;
				assign node15031 = (inp[13]) ? node16559 : node15032;
					assign node15032 = (inp[14]) ? node15746 : node15033;
						assign node15033 = (inp[1]) ? node15383 : node15034;
							assign node15034 = (inp[8]) ? node15206 : node15035;
								assign node15035 = (inp[5]) ? node15127 : node15036;
									assign node15036 = (inp[10]) ? node15076 : node15037;
										assign node15037 = (inp[4]) ? node15049 : node15038;
											assign node15038 = (inp[2]) ? node15044 : node15039;
												assign node15039 = (inp[3]) ? 16'b0000111111111111 : node15040;
													assign node15040 = (inp[11]) ? 16'b0000111111111111 : 16'b0001111111111111;
												assign node15044 = (inp[6]) ? 16'b0000001111111111 : node15045;
													assign node15045 = (inp[3]) ? 16'b0000011111111111 : 16'b0001111111111111;
											assign node15049 = (inp[9]) ? node15061 : node15050;
												assign node15050 = (inp[3]) ? node15056 : node15051;
													assign node15051 = (inp[11]) ? node15053 : 16'b0000111111111111;
														assign node15053 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node15056 = (inp[15]) ? node15058 : 16'b0000001111111111;
														assign node15058 = (inp[6]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node15061 = (inp[15]) ? node15067 : node15062;
													assign node15062 = (inp[6]) ? node15064 : 16'b0000001111111111;
														assign node15064 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node15067 = (inp[6]) ? 16'b0000000111111111 : node15068;
														assign node15068 = (inp[3]) ? 16'b0000000111111111 : node15069;
															assign node15069 = (inp[11]) ? node15071 : 16'b0000001111111111;
																assign node15071 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node15076 = (inp[11]) ? node15104 : node15077;
											assign node15077 = (inp[6]) ? node15087 : node15078;
												assign node15078 = (inp[15]) ? node15082 : node15079;
													assign node15079 = (inp[3]) ? 16'b0000001111111111 : 16'b0000111111111111;
													assign node15082 = (inp[4]) ? 16'b0000001111111111 : node15083;
														assign node15083 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node15087 = (inp[2]) ? node15097 : node15088;
													assign node15088 = (inp[3]) ? node15094 : node15089;
														assign node15089 = (inp[9]) ? 16'b0000001111111111 : node15090;
															assign node15090 = (inp[4]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node15094 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node15097 = (inp[4]) ? node15101 : node15098;
														assign node15098 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node15101 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node15104 = (inp[4]) ? node15122 : node15105;
												assign node15105 = (inp[3]) ? node15113 : node15106;
													assign node15106 = (inp[9]) ? node15110 : node15107;
														assign node15107 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node15110 = (inp[6]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node15113 = (inp[2]) ? node15117 : node15114;
														assign node15114 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node15117 = (inp[6]) ? node15119 : 16'b0000000111111111;
															assign node15119 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node15122 = (inp[3]) ? node15124 : 16'b0000000011111111;
													assign node15124 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node15127 = (inp[10]) ? node15169 : node15128;
										assign node15128 = (inp[15]) ? node15146 : node15129;
											assign node15129 = (inp[3]) ? node15137 : node15130;
												assign node15130 = (inp[11]) ? node15132 : 16'b0000011111111111;
													assign node15132 = (inp[4]) ? 16'b0000000111111111 : node15133;
														assign node15133 = (inp[2]) ? 16'b0000001111111111 : 16'b0000111111111111;
												assign node15137 = (inp[6]) ? node15139 : 16'b0000001111111111;
													assign node15139 = (inp[4]) ? 16'b0000000011111111 : node15140;
														assign node15140 = (inp[9]) ? node15142 : 16'b0000001111111111;
															assign node15142 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node15146 = (inp[11]) ? node15158 : node15147;
												assign node15147 = (inp[4]) ? node15155 : node15148;
													assign node15148 = (inp[6]) ? node15152 : node15149;
														assign node15149 = (inp[3]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node15152 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node15155 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node15158 = (inp[9]) ? node15164 : node15159;
													assign node15159 = (inp[2]) ? node15161 : 16'b0000001111111111;
														assign node15161 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node15164 = (inp[3]) ? 16'b0000000011111111 : node15165;
														assign node15165 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node15169 = (inp[6]) ? node15187 : node15170;
											assign node15170 = (inp[9]) ? node15178 : node15171;
												assign node15171 = (inp[4]) ? node15175 : node15172;
													assign node15172 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node15175 = (inp[11]) ? 16'b0000000011111111 : 16'b0000001111111111;
												assign node15178 = (inp[11]) ? node15180 : 16'b0000000111111111;
													assign node15180 = (inp[2]) ? node15184 : node15181;
														assign node15181 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node15184 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node15187 = (inp[4]) ? node15197 : node15188;
												assign node15188 = (inp[9]) ? node15192 : node15189;
													assign node15189 = (inp[3]) ? 16'b0000000011111111 : 16'b0000001111111111;
													assign node15192 = (inp[11]) ? node15194 : 16'b0000000011111111;
														assign node15194 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node15197 = (inp[3]) ? 16'b0000000000011111 : node15198;
													assign node15198 = (inp[2]) ? node15200 : 16'b0000000011111111;
														assign node15200 = (inp[11]) ? node15202 : 16'b0000000001111111;
															assign node15202 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
								assign node15206 = (inp[11]) ? node15292 : node15207;
									assign node15207 = (inp[3]) ? node15253 : node15208;
										assign node15208 = (inp[2]) ? node15232 : node15209;
											assign node15209 = (inp[5]) ? node15223 : node15210;
												assign node15210 = (inp[9]) ? node15218 : node15211;
													assign node15211 = (inp[10]) ? node15215 : node15212;
														assign node15212 = (inp[4]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node15215 = (inp[6]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node15218 = (inp[6]) ? node15220 : 16'b0000001111111111;
														assign node15220 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node15223 = (inp[9]) ? node15225 : 16'b0000001111111111;
													assign node15225 = (inp[15]) ? 16'b0000000011111111 : node15226;
														assign node15226 = (inp[10]) ? 16'b0000000111111111 : node15227;
															assign node15227 = (inp[6]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node15232 = (inp[6]) ? node15246 : node15233;
												assign node15233 = (inp[10]) ? node15237 : node15234;
													assign node15234 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node15237 = (inp[9]) ? 16'b0000000111111111 : node15238;
														assign node15238 = (inp[4]) ? 16'b0000000111111111 : node15239;
															assign node15239 = (inp[15]) ? node15241 : 16'b0000001111111111;
																assign node15241 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node15246 = (inp[15]) ? 16'b0000000011111111 : node15247;
													assign node15247 = (inp[10]) ? node15249 : 16'b0000000111111111;
														assign node15249 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node15253 = (inp[6]) ? node15275 : node15254;
											assign node15254 = (inp[10]) ? node15260 : node15255;
												assign node15255 = (inp[4]) ? 16'b0000000111111111 : node15256;
													assign node15256 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node15260 = (inp[9]) ? node15270 : node15261;
													assign node15261 = (inp[4]) ? node15267 : node15262;
														assign node15262 = (inp[2]) ? 16'b0000000111111111 : node15263;
															assign node15263 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node15267 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node15270 = (inp[2]) ? node15272 : 16'b0000000111111111;
														assign node15272 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000001111111;
											assign node15275 = (inp[4]) ? node15283 : node15276;
												assign node15276 = (inp[5]) ? node15280 : node15277;
													assign node15277 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node15280 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000111111111;
												assign node15283 = (inp[10]) ? node15285 : 16'b0000000011111111;
													assign node15285 = (inp[15]) ? node15287 : 16'b0000000011111111;
														assign node15287 = (inp[2]) ? node15289 : 16'b0000000000111111;
															assign node15289 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node15292 = (inp[3]) ? node15340 : node15293;
										assign node15293 = (inp[2]) ? node15317 : node15294;
											assign node15294 = (inp[15]) ? node15304 : node15295;
												assign node15295 = (inp[4]) ? node15299 : node15296;
													assign node15296 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node15299 = (inp[10]) ? node15301 : 16'b0000001111111111;
														assign node15301 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node15304 = (inp[6]) ? node15314 : node15305;
													assign node15305 = (inp[10]) ? node15307 : 16'b0000000111111111;
														assign node15307 = (inp[5]) ? node15309 : 16'b0000000111111111;
															assign node15309 = (inp[4]) ? 16'b0000000011111111 : node15310;
																assign node15310 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node15314 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000011111111;
											assign node15317 = (inp[9]) ? node15331 : node15318;
												assign node15318 = (inp[10]) ? node15322 : node15319;
													assign node15319 = (inp[15]) ? 16'b0000001111111111 : 16'b0000000111111111;
													assign node15322 = (inp[6]) ? node15326 : node15323;
														assign node15323 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node15326 = (inp[5]) ? node15328 : 16'b0000000011111111;
															assign node15328 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node15331 = (inp[4]) ? node15335 : node15332;
													assign node15332 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node15335 = (inp[6]) ? 16'b0000000001111111 : node15336;
														assign node15336 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node15340 = (inp[10]) ? node15364 : node15341;
											assign node15341 = (inp[15]) ? node15357 : node15342;
												assign node15342 = (inp[4]) ? node15348 : node15343;
													assign node15343 = (inp[9]) ? node15345 : 16'b0000000111111111;
														assign node15345 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node15348 = (inp[2]) ? node15352 : node15349;
														assign node15349 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node15352 = (inp[5]) ? node15354 : 16'b0000000011111111;
															assign node15354 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node15357 = (inp[2]) ? node15359 : 16'b0000000011111111;
													assign node15359 = (inp[9]) ? 16'b0000000001111111 : node15360;
														assign node15360 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node15364 = (inp[4]) ? node15376 : node15365;
												assign node15365 = (inp[5]) ? node15367 : 16'b0000000011111111;
													assign node15367 = (inp[9]) ? node15373 : node15368;
														assign node15368 = (inp[6]) ? 16'b0000000001111111 : node15369;
															assign node15369 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node15373 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node15376 = (inp[2]) ? node15378 : 16'b0000000001111111;
													assign node15378 = (inp[9]) ? node15380 : 16'b0000000000111111;
														assign node15380 = (inp[6]) ? 16'b0000000000001111 : 16'b0000000000011111;
							assign node15383 = (inp[8]) ? node15567 : node15384;
								assign node15384 = (inp[15]) ? node15480 : node15385;
									assign node15385 = (inp[11]) ? node15437 : node15386;
										assign node15386 = (inp[2]) ? node15410 : node15387;
											assign node15387 = (inp[9]) ? node15397 : node15388;
												assign node15388 = (inp[3]) ? node15392 : node15389;
													assign node15389 = (inp[5]) ? 16'b0000011111111111 : 16'b0001111111111111;
													assign node15392 = (inp[6]) ? 16'b0000001111111111 : node15393;
														assign node15393 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node15397 = (inp[10]) ? node15403 : node15398;
													assign node15398 = (inp[4]) ? 16'b0000001111111111 : node15399;
														assign node15399 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node15403 = (inp[6]) ? 16'b0000000111111111 : node15404;
														assign node15404 = (inp[5]) ? node15406 : 16'b0000001111111111;
															assign node15406 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node15410 = (inp[5]) ? node15420 : node15411;
												assign node15411 = (inp[9]) ? 16'b0000000111111111 : node15412;
													assign node15412 = (inp[4]) ? node15416 : node15413;
														assign node15413 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node15416 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node15420 = (inp[3]) ? node15428 : node15421;
													assign node15421 = (inp[6]) ? 16'b0000000011111111 : node15422;
														assign node15422 = (inp[4]) ? node15424 : 16'b0000001111111111;
															assign node15424 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node15428 = (inp[10]) ? node15432 : node15429;
														assign node15429 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node15432 = (inp[9]) ? node15434 : 16'b0000000011111111;
															assign node15434 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node15437 = (inp[10]) ? node15455 : node15438;
											assign node15438 = (inp[9]) ? node15448 : node15439;
												assign node15439 = (inp[6]) ? node15445 : node15440;
													assign node15440 = (inp[4]) ? node15442 : 16'b0000011111111111;
														assign node15442 = (inp[2]) ? 16'b0000001111111111 : 16'b0000000111111111;
													assign node15445 = (inp[3]) ? 16'b0000001111111111 : 16'b0000000111111111;
												assign node15448 = (inp[5]) ? 16'b0000000011111111 : node15449;
													assign node15449 = (inp[6]) ? 16'b0000000001111111 : node15450;
														assign node15450 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node15455 = (inp[2]) ? node15473 : node15456;
												assign node15456 = (inp[4]) ? node15468 : node15457;
													assign node15457 = (inp[9]) ? node15461 : node15458;
														assign node15458 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node15461 = (inp[3]) ? node15463 : 16'b0000001111111111;
															assign node15463 = (inp[5]) ? 16'b0000000011111111 : node15464;
																assign node15464 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node15468 = (inp[3]) ? node15470 : 16'b0000000011111111;
														assign node15470 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node15473 = (inp[5]) ? 16'b0000000001111111 : node15474;
													assign node15474 = (inp[6]) ? 16'b0000000000111111 : node15475;
														assign node15475 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node15480 = (inp[5]) ? node15532 : node15481;
										assign node15481 = (inp[11]) ? node15503 : node15482;
											assign node15482 = (inp[10]) ? node15492 : node15483;
												assign node15483 = (inp[6]) ? node15487 : node15484;
													assign node15484 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node15487 = (inp[2]) ? 16'b0000000111111111 : node15488;
														assign node15488 = (inp[4]) ? 16'b0000000111111111 : 16'b0000011111111111;
												assign node15492 = (inp[9]) ? node15494 : 16'b0000000111111111;
													assign node15494 = (inp[6]) ? 16'b0000000001111111 : node15495;
														assign node15495 = (inp[4]) ? 16'b0000000011111111 : node15496;
															assign node15496 = (inp[3]) ? node15498 : 16'b0000000111111111;
																assign node15498 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node15503 = (inp[2]) ? node15511 : node15504;
												assign node15504 = (inp[4]) ? node15506 : 16'b0000000111111111;
													assign node15506 = (inp[3]) ? 16'b0000000011111111 : node15507;
														assign node15507 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node15511 = (inp[4]) ? node15521 : node15512;
													assign node15512 = (inp[3]) ? 16'b0000000011111111 : node15513;
														assign node15513 = (inp[10]) ? node15515 : 16'b0000000111111111;
															assign node15515 = (inp[9]) ? 16'b0000000011111111 : node15516;
																assign node15516 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node15521 = (inp[3]) ? node15529 : node15522;
														assign node15522 = (inp[10]) ? 16'b0000000001111111 : node15523;
															assign node15523 = (inp[9]) ? node15525 : 16'b0000000011111111;
																assign node15525 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node15529 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node15532 = (inp[6]) ? node15556 : node15533;
											assign node15533 = (inp[3]) ? node15543 : node15534;
												assign node15534 = (inp[11]) ? node15536 : 16'b0000000111111111;
													assign node15536 = (inp[9]) ? node15538 : 16'b0000000111111111;
														assign node15538 = (inp[2]) ? node15540 : 16'b0000000011111111;
															assign node15540 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000011111111;
												assign node15543 = (inp[9]) ? node15551 : node15544;
													assign node15544 = (inp[2]) ? node15546 : 16'b0000000111111111;
														assign node15546 = (inp[4]) ? node15548 : 16'b0000000011111111;
															assign node15548 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000011111111;
													assign node15551 = (inp[11]) ? node15553 : 16'b0000000001111111;
														assign node15553 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node15556 = (inp[11]) ? 16'b0000000000111111 : node15557;
												assign node15557 = (inp[9]) ? node15559 : 16'b0000000001111111;
													assign node15559 = (inp[3]) ? node15561 : 16'b0000000001111111;
														assign node15561 = (inp[4]) ? node15563 : 16'b0000000000111111;
															assign node15563 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
								assign node15567 = (inp[3]) ? node15649 : node15568;
									assign node15568 = (inp[11]) ? node15610 : node15569;
										assign node15569 = (inp[4]) ? node15591 : node15570;
											assign node15570 = (inp[10]) ? node15580 : node15571;
												assign node15571 = (inp[5]) ? node15575 : node15572;
													assign node15572 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node15575 = (inp[9]) ? 16'b0000000111111111 : node15576;
														assign node15576 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node15580 = (inp[15]) ? node15586 : node15581;
													assign node15581 = (inp[5]) ? 16'b0000000111111111 : node15582;
														assign node15582 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node15586 = (inp[6]) ? 16'b0000000011111111 : node15587;
														assign node15587 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node15591 = (inp[9]) ? node15603 : node15592;
												assign node15592 = (inp[2]) ? node15598 : node15593;
													assign node15593 = (inp[15]) ? 16'b0000000111111111 : node15594;
														assign node15594 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node15598 = (inp[15]) ? 16'b0000000011111111 : node15599;
														assign node15599 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node15603 = (inp[10]) ? node15605 : 16'b0000000011111111;
													assign node15605 = (inp[15]) ? 16'b0000000001111111 : node15606;
														assign node15606 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000011111111;
										assign node15610 = (inp[5]) ? node15628 : node15611;
											assign node15611 = (inp[6]) ? node15621 : node15612;
												assign node15612 = (inp[10]) ? 16'b0000000011111111 : node15613;
													assign node15613 = (inp[4]) ? node15615 : 16'b0000000111111111;
														assign node15615 = (inp[9]) ? 16'b0000000011111111 : node15616;
															assign node15616 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node15621 = (inp[9]) ? node15625 : node15622;
													assign node15622 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node15625 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node15628 = (inp[15]) ? node15638 : node15629;
												assign node15629 = (inp[9]) ? node15635 : node15630;
													assign node15630 = (inp[10]) ? node15632 : 16'b0000000111111111;
														assign node15632 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node15635 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node15638 = (inp[4]) ? node15644 : node15639;
													assign node15639 = (inp[6]) ? node15641 : 16'b0000000001111111;
														assign node15641 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node15644 = (inp[6]) ? node15646 : 16'b0000000000111111;
														assign node15646 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node15649 = (inp[4]) ? node15709 : node15650;
										assign node15650 = (inp[5]) ? node15684 : node15651;
											assign node15651 = (inp[9]) ? node15669 : node15652;
												assign node15652 = (inp[15]) ? node15660 : node15653;
													assign node15653 = (inp[11]) ? node15657 : node15654;
														assign node15654 = (inp[6]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node15657 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node15660 = (inp[11]) ? node15664 : node15661;
														assign node15661 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node15664 = (inp[2]) ? 16'b0000000011111111 : node15665;
															assign node15665 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node15669 = (inp[2]) ? node15679 : node15670;
													assign node15670 = (inp[11]) ? node15674 : node15671;
														assign node15671 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node15674 = (inp[10]) ? node15676 : 16'b0000000011111111;
															assign node15676 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node15679 = (inp[15]) ? node15681 : 16'b0000000001111111;
														assign node15681 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node15684 = (inp[2]) ? node15698 : node15685;
												assign node15685 = (inp[10]) ? node15693 : node15686;
													assign node15686 = (inp[11]) ? 16'b0000000001111111 : node15687;
														assign node15687 = (inp[9]) ? node15689 : 16'b0000000011111111;
															assign node15689 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node15693 = (inp[11]) ? node15695 : 16'b0000000001111111;
														assign node15695 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node15698 = (inp[9]) ? node15704 : node15699;
													assign node15699 = (inp[15]) ? 16'b0000000001111111 : node15700;
														assign node15700 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node15704 = (inp[15]) ? 16'b0000000000011111 : node15705;
														assign node15705 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node15709 = (inp[2]) ? node15719 : node15710;
											assign node15710 = (inp[5]) ? node15714 : node15711;
												assign node15711 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node15714 = (inp[11]) ? 16'b0000000000111111 : node15715;
													assign node15715 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000011111111;
											assign node15719 = (inp[11]) ? node15737 : node15720;
												assign node15720 = (inp[15]) ? node15724 : node15721;
													assign node15721 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node15724 = (inp[9]) ? node15730 : node15725;
														assign node15725 = (inp[6]) ? node15727 : 16'b0000000001111111;
															assign node15727 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node15730 = (inp[5]) ? 16'b0000000000011111 : node15731;
															assign node15731 = (inp[10]) ? node15733 : 16'b0000000000111111;
																assign node15733 = (inp[6]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node15737 = (inp[9]) ? node15743 : node15738;
													assign node15738 = (inp[6]) ? node15740 : 16'b0000000000111111;
														assign node15740 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node15743 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000111111;
						assign node15746 = (inp[5]) ? node16144 : node15747;
							assign node15747 = (inp[11]) ? node15927 : node15748;
								assign node15748 = (inp[8]) ? node15848 : node15749;
									assign node15749 = (inp[9]) ? node15791 : node15750;
										assign node15750 = (inp[3]) ? node15766 : node15751;
											assign node15751 = (inp[4]) ? node15759 : node15752;
												assign node15752 = (inp[1]) ? node15754 : 16'b0000011111111111;
													assign node15754 = (inp[2]) ? 16'b0000001111111111 : node15755;
														assign node15755 = (inp[6]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node15759 = (inp[1]) ? 16'b0000001111111111 : node15760;
													assign node15760 = (inp[6]) ? node15762 : 16'b0000111111111111;
														assign node15762 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node15766 = (inp[15]) ? node15784 : node15767;
												assign node15767 = (inp[10]) ? node15771 : node15768;
													assign node15768 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node15771 = (inp[2]) ? node15777 : node15772;
														assign node15772 = (inp[6]) ? node15774 : 16'b0000001111111111;
															assign node15774 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node15777 = (inp[6]) ? node15779 : 16'b0000000111111111;
															assign node15779 = (inp[4]) ? 16'b0000000011111111 : node15780;
																assign node15780 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node15784 = (inp[10]) ? node15788 : node15785;
													assign node15785 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node15788 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node15791 = (inp[2]) ? node15823 : node15792;
											assign node15792 = (inp[15]) ? node15812 : node15793;
												assign node15793 = (inp[10]) ? node15805 : node15794;
													assign node15794 = (inp[1]) ? node15798 : node15795;
														assign node15795 = (inp[3]) ? 16'b0000001111111111 : 16'b0000111111111111;
														assign node15798 = (inp[6]) ? 16'b0000000111111111 : node15799;
															assign node15799 = (inp[4]) ? node15801 : 16'b0000001111111111;
																assign node15801 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node15805 = (inp[1]) ? node15809 : node15806;
														assign node15806 = (inp[6]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node15809 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node15812 = (inp[3]) ? node15814 : 16'b0000000111111111;
													assign node15814 = (inp[4]) ? node15820 : node15815;
														assign node15815 = (inp[10]) ? node15817 : 16'b0000000111111111;
															assign node15817 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node15820 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node15823 = (inp[3]) ? node15837 : node15824;
												assign node15824 = (inp[10]) ? node15832 : node15825;
													assign node15825 = (inp[6]) ? node15827 : 16'b0000001111111111;
														assign node15827 = (inp[15]) ? 16'b0000000011111111 : node15828;
															assign node15828 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node15832 = (inp[4]) ? node15834 : 16'b0000000011111111;
														assign node15834 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000001111111;
												assign node15837 = (inp[1]) ? node15843 : node15838;
													assign node15838 = (inp[6]) ? node15840 : 16'b0000000111111111;
														assign node15840 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node15843 = (inp[10]) ? node15845 : 16'b0000000001111111;
														assign node15845 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node15848 = (inp[1]) ? node15882 : node15849;
										assign node15849 = (inp[6]) ? node15865 : node15850;
											assign node15850 = (inp[3]) ? node15856 : node15851;
												assign node15851 = (inp[2]) ? node15853 : 16'b0000001111111111;
													assign node15853 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node15856 = (inp[2]) ? 16'b0000000011111111 : node15857;
													assign node15857 = (inp[15]) ? node15861 : node15858;
														assign node15858 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node15861 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node15865 = (inp[4]) ? node15875 : node15866;
												assign node15866 = (inp[2]) ? 16'b0000000011111111 : node15867;
													assign node15867 = (inp[15]) ? node15871 : node15868;
														assign node15868 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node15871 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node15875 = (inp[9]) ? 16'b0000000001111111 : node15876;
													assign node15876 = (inp[15]) ? 16'b0000000001111111 : node15877;
														assign node15877 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node15882 = (inp[4]) ? node15910 : node15883;
											assign node15883 = (inp[2]) ? node15895 : node15884;
												assign node15884 = (inp[9]) ? node15890 : node15885;
													assign node15885 = (inp[15]) ? node15887 : 16'b0000001111111111;
														assign node15887 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node15890 = (inp[10]) ? node15892 : 16'b0000000011111111;
														assign node15892 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000111111111;
												assign node15895 = (inp[3]) ? node15905 : node15896;
													assign node15896 = (inp[9]) ? node15902 : node15897;
														assign node15897 = (inp[10]) ? 16'b0000000011111111 : node15898;
															assign node15898 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node15902 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node15905 = (inp[6]) ? node15907 : 16'b0000000001111111;
														assign node15907 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node15910 = (inp[15]) ? node15920 : node15911;
												assign node15911 = (inp[3]) ? node15917 : node15912;
													assign node15912 = (inp[9]) ? 16'b0000000001111111 : node15913;
														assign node15913 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node15917 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000000111111;
												assign node15920 = (inp[3]) ? node15924 : node15921;
													assign node15921 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node15924 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
								assign node15927 = (inp[1]) ? node16021 : node15928;
									assign node15928 = (inp[2]) ? node15978 : node15929;
										assign node15929 = (inp[10]) ? node15951 : node15930;
											assign node15930 = (inp[15]) ? node15948 : node15931;
												assign node15931 = (inp[4]) ? node15939 : node15932;
													assign node15932 = (inp[6]) ? node15934 : 16'b0000111111111111;
														assign node15934 = (inp[8]) ? node15936 : 16'b0000001111111111;
															assign node15936 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node15939 = (inp[9]) ? 16'b0000000111111111 : node15940;
														assign node15940 = (inp[3]) ? 16'b0000000111111111 : node15941;
															assign node15941 = (inp[8]) ? node15943 : 16'b0000001111111111;
																assign node15943 = (inp[6]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node15948 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000111111111;
											assign node15951 = (inp[6]) ? node15969 : node15952;
												assign node15952 = (inp[3]) ? node15958 : node15953;
													assign node15953 = (inp[9]) ? 16'b0000000111111111 : node15954;
														assign node15954 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node15958 = (inp[15]) ? node15966 : node15959;
														assign node15959 = (inp[4]) ? node15961 : 16'b0000000111111111;
															assign node15961 = (inp[9]) ? 16'b0000000011111111 : node15962;
																assign node15962 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node15966 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node15969 = (inp[8]) ? node15973 : node15970;
													assign node15970 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000111111111;
													assign node15973 = (inp[15]) ? node15975 : 16'b0000000001111111;
														assign node15975 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node15978 = (inp[3]) ? node15996 : node15979;
											assign node15979 = (inp[9]) ? node15987 : node15980;
												assign node15980 = (inp[15]) ? node15982 : 16'b0000000111111111;
													assign node15982 = (inp[4]) ? 16'b0000000011111111 : node15983;
														assign node15983 = (inp[10]) ? 16'b0000000011111111 : 16'b0000001111111111;
												assign node15987 = (inp[8]) ? node15989 : 16'b0000000011111111;
													assign node15989 = (inp[10]) ? 16'b0000000001111111 : node15990;
														assign node15990 = (inp[15]) ? node15992 : 16'b0000000011111111;
															assign node15992 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node15996 = (inp[15]) ? node16014 : node15997;
												assign node15997 = (inp[8]) ? node16009 : node15998;
													assign node15998 = (inp[6]) ? node16000 : 16'b0000000111111111;
														assign node16000 = (inp[4]) ? node16004 : node16001;
															assign node16001 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
															assign node16004 = (inp[10]) ? 16'b0000000001111111 : node16005;
																assign node16005 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node16009 = (inp[10]) ? node16011 : 16'b0000000001111111;
														assign node16011 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node16014 = (inp[9]) ? 16'b0000000000111111 : node16015;
													assign node16015 = (inp[8]) ? node16017 : 16'b0000000001111111;
														assign node16017 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node16021 = (inp[10]) ? node16077 : node16022;
										assign node16022 = (inp[8]) ? node16046 : node16023;
											assign node16023 = (inp[4]) ? node16037 : node16024;
												assign node16024 = (inp[9]) ? node16030 : node16025;
													assign node16025 = (inp[6]) ? node16027 : 16'b0000000111111111;
														assign node16027 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node16030 = (inp[2]) ? node16034 : node16031;
														assign node16031 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node16034 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node16037 = (inp[6]) ? node16039 : 16'b0000000011111111;
													assign node16039 = (inp[3]) ? node16043 : node16040;
														assign node16040 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node16043 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node16046 = (inp[9]) ? node16062 : node16047;
												assign node16047 = (inp[3]) ? node16053 : node16048;
													assign node16048 = (inp[6]) ? node16050 : 16'b0000000011111111;
														assign node16050 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node16053 = (inp[2]) ? node16057 : node16054;
														assign node16054 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node16057 = (inp[6]) ? 16'b0000000000111111 : node16058;
															assign node16058 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node16062 = (inp[4]) ? node16070 : node16063;
													assign node16063 = (inp[6]) ? node16065 : 16'b0000000111111111;
														assign node16065 = (inp[15]) ? node16067 : 16'b0000000001111111;
															assign node16067 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node16070 = (inp[6]) ? node16074 : node16071;
														assign node16071 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node16074 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node16077 = (inp[2]) ? node16115 : node16078;
											assign node16078 = (inp[8]) ? node16098 : node16079;
												assign node16079 = (inp[3]) ? node16091 : node16080;
													assign node16080 = (inp[15]) ? node16084 : node16081;
														assign node16081 = (inp[6]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node16084 = (inp[6]) ? 16'b0000000011111111 : node16085;
															assign node16085 = (inp[4]) ? 16'b0000000011111111 : node16086;
																assign node16086 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node16091 = (inp[9]) ? node16095 : node16092;
														assign node16092 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node16095 = (inp[6]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node16098 = (inp[3]) ? node16104 : node16099;
													assign node16099 = (inp[15]) ? node16101 : 16'b0000000001111111;
														assign node16101 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000000111111;
													assign node16104 = (inp[4]) ? node16108 : node16105;
														assign node16105 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node16108 = (inp[6]) ? node16110 : 16'b0000000000111111;
															assign node16110 = (inp[15]) ? node16112 : 16'b0000000000011111;
																assign node16112 = (inp[9]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node16115 = (inp[8]) ? node16133 : node16116;
												assign node16116 = (inp[15]) ? node16122 : node16117;
													assign node16117 = (inp[3]) ? node16119 : 16'b0000000000111111;
														assign node16119 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node16122 = (inp[9]) ? node16124 : 16'b0000000000111111;
														assign node16124 = (inp[6]) ? node16130 : node16125;
															assign node16125 = (inp[4]) ? node16127 : 16'b0000000000111111;
																assign node16127 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000000111111;
															assign node16130 = (inp[4]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node16133 = (inp[3]) ? node16137 : node16134;
													assign node16134 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node16137 = (inp[9]) ? 16'b0000000000001111 : node16138;
														assign node16138 = (inp[6]) ? node16140 : 16'b0000000000011111;
															assign node16140 = (inp[4]) ? 16'b0000000000001111 : 16'b0000000000011111;
							assign node16144 = (inp[9]) ? node16366 : node16145;
								assign node16145 = (inp[4]) ? node16255 : node16146;
									assign node16146 = (inp[15]) ? node16198 : node16147;
										assign node16147 = (inp[2]) ? node16179 : node16148;
											assign node16148 = (inp[10]) ? node16162 : node16149;
												assign node16149 = (inp[8]) ? node16155 : node16150;
													assign node16150 = (inp[6]) ? 16'b0000001111111111 : node16151;
														assign node16151 = (inp[11]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node16155 = (inp[6]) ? 16'b0000000111111111 : node16156;
														assign node16156 = (inp[1]) ? node16158 : 16'b0000001111111111;
															assign node16158 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node16162 = (inp[3]) ? node16166 : node16163;
													assign node16163 = (inp[6]) ? 16'b0000000011111111 : 16'b0000001111111111;
													assign node16166 = (inp[8]) ? node16172 : node16167;
														assign node16167 = (inp[11]) ? 16'b0000000011111111 : node16168;
															assign node16168 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node16172 = (inp[1]) ? 16'b0000000001111111 : node16173;
															assign node16173 = (inp[11]) ? node16175 : 16'b0000000011111111;
																assign node16175 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node16179 = (inp[11]) ? node16187 : node16180;
												assign node16180 = (inp[1]) ? node16184 : node16181;
													assign node16181 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node16184 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node16187 = (inp[3]) ? node16193 : node16188;
													assign node16188 = (inp[6]) ? node16190 : 16'b0000000011111111;
														assign node16190 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node16193 = (inp[1]) ? 16'b0000000001111111 : node16194;
														assign node16194 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node16198 = (inp[3]) ? node16226 : node16199;
											assign node16199 = (inp[10]) ? node16215 : node16200;
												assign node16200 = (inp[11]) ? node16210 : node16201;
													assign node16201 = (inp[8]) ? node16207 : node16202;
														assign node16202 = (inp[1]) ? 16'b0000000111111111 : node16203;
															assign node16203 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node16207 = (inp[1]) ? 16'b0000000111111111 : 16'b0000000011111111;
													assign node16210 = (inp[1]) ? 16'b0000000011111111 : node16211;
														assign node16211 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node16215 = (inp[2]) ? 16'b0000000001111111 : node16216;
													assign node16216 = (inp[6]) ? node16218 : 16'b0000000011111111;
														assign node16218 = (inp[1]) ? node16222 : node16219;
															assign node16219 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
															assign node16222 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node16226 = (inp[6]) ? node16240 : node16227;
												assign node16227 = (inp[8]) ? node16237 : node16228;
													assign node16228 = (inp[2]) ? node16234 : node16229;
														assign node16229 = (inp[10]) ? 16'b0000000011111111 : node16230;
															assign node16230 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node16234 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000011111111;
													assign node16237 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node16240 = (inp[1]) ? node16246 : node16241;
													assign node16241 = (inp[10]) ? node16243 : 16'b0000000001111111;
														assign node16243 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node16246 = (inp[8]) ? node16252 : node16247;
														assign node16247 = (inp[10]) ? 16'b0000000000111111 : node16248;
															assign node16248 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node16252 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node16255 = (inp[8]) ? node16313 : node16256;
										assign node16256 = (inp[11]) ? node16280 : node16257;
											assign node16257 = (inp[6]) ? node16269 : node16258;
												assign node16258 = (inp[3]) ? node16264 : node16259;
													assign node16259 = (inp[10]) ? 16'b0000000011111111 : node16260;
														assign node16260 = (inp[1]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node16264 = (inp[10]) ? 16'b0000000011111111 : node16265;
														assign node16265 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node16269 = (inp[10]) ? node16271 : 16'b0000000011111111;
													assign node16271 = (inp[15]) ? 16'b0000000000111111 : node16272;
														assign node16272 = (inp[1]) ? 16'b0000000001111111 : node16273;
															assign node16273 = (inp[3]) ? node16275 : 16'b0000000011111111;
																assign node16275 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node16280 = (inp[3]) ? node16300 : node16281;
												assign node16281 = (inp[2]) ? node16289 : node16282;
													assign node16282 = (inp[1]) ? node16286 : node16283;
														assign node16283 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node16286 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node16289 = (inp[15]) ? node16293 : node16290;
														assign node16290 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000111111111;
														assign node16293 = (inp[10]) ? 16'b0000000000111111 : node16294;
															assign node16294 = (inp[6]) ? node16296 : 16'b0000000001111111;
																assign node16296 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node16300 = (inp[6]) ? node16306 : node16301;
													assign node16301 = (inp[10]) ? node16303 : 16'b0000000001111111;
														assign node16303 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000000111111;
													assign node16306 = (inp[1]) ? node16310 : node16307;
														assign node16307 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node16310 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node16313 = (inp[11]) ? node16341 : node16314;
											assign node16314 = (inp[6]) ? node16328 : node16315;
												assign node16315 = (inp[15]) ? node16319 : node16316;
													assign node16316 = (inp[1]) ? 16'b0000000111111111 : 16'b0000000011111111;
													assign node16319 = (inp[2]) ? node16323 : node16320;
														assign node16320 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000001111111;
														assign node16323 = (inp[1]) ? 16'b0000000000111111 : node16324;
															assign node16324 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node16328 = (inp[15]) ? node16336 : node16329;
													assign node16329 = (inp[1]) ? node16331 : 16'b0000000001111111;
														assign node16331 = (inp[10]) ? node16333 : 16'b0000000001111111;
															assign node16333 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node16336 = (inp[1]) ? node16338 : 16'b0000000000111111;
														assign node16338 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node16341 = (inp[6]) ? node16355 : node16342;
												assign node16342 = (inp[1]) ? node16346 : node16343;
													assign node16343 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node16346 = (inp[10]) ? node16352 : node16347;
														assign node16347 = (inp[15]) ? 16'b0000000000111111 : node16348;
															assign node16348 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node16352 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node16355 = (inp[3]) ? node16361 : node16356;
													assign node16356 = (inp[10]) ? 16'b0000000000011111 : node16357;
														assign node16357 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node16361 = (inp[1]) ? node16363 : 16'b0000000000011111;
														assign node16363 = (inp[10]) ? 16'b0000000000001111 : 16'b0000000000011111;
								assign node16366 = (inp[8]) ? node16478 : node16367;
									assign node16367 = (inp[6]) ? node16427 : node16368;
										assign node16368 = (inp[1]) ? node16394 : node16369;
											assign node16369 = (inp[15]) ? node16383 : node16370;
												assign node16370 = (inp[2]) ? node16374 : node16371;
													assign node16371 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node16374 = (inp[10]) ? 16'b0000000011111111 : node16375;
														assign node16375 = (inp[4]) ? 16'b0000000011111111 : node16376;
															assign node16376 = (inp[3]) ? node16378 : 16'b0000000111111111;
																assign node16378 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node16383 = (inp[10]) ? 16'b0000000001111111 : node16384;
													assign node16384 = (inp[2]) ? node16388 : node16385;
														assign node16385 = (inp[11]) ? 16'b0000000111111111 : 16'b0000000011111111;
														assign node16388 = (inp[11]) ? node16390 : 16'b0000000011111111;
															assign node16390 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node16394 = (inp[11]) ? node16408 : node16395;
												assign node16395 = (inp[3]) ? node16401 : node16396;
													assign node16396 = (inp[4]) ? node16398 : 16'b0000000011111111;
														assign node16398 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node16401 = (inp[10]) ? node16405 : node16402;
														assign node16402 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node16405 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node16408 = (inp[15]) ? node16420 : node16409;
													assign node16409 = (inp[2]) ? node16415 : node16410;
														assign node16410 = (inp[10]) ? 16'b0000000001111111 : node16411;
															assign node16411 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node16415 = (inp[10]) ? 16'b0000000000111111 : node16416;
															assign node16416 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node16420 = (inp[10]) ? node16424 : node16421;
														assign node16421 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node16424 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node16427 = (inp[2]) ? node16449 : node16428;
											assign node16428 = (inp[4]) ? node16442 : node16429;
												assign node16429 = (inp[10]) ? node16437 : node16430;
													assign node16430 = (inp[11]) ? node16432 : 16'b0000000111111111;
														assign node16432 = (inp[1]) ? node16434 : 16'b0000000011111111;
															assign node16434 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node16437 = (inp[11]) ? node16439 : 16'b0000000001111111;
														assign node16439 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node16442 = (inp[3]) ? node16444 : 16'b0000000001111111;
													assign node16444 = (inp[11]) ? 16'b0000000000111111 : node16445;
														assign node16445 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node16449 = (inp[4]) ? node16461 : node16450;
												assign node16450 = (inp[10]) ? node16452 : 16'b0000000001111111;
													assign node16452 = (inp[15]) ? node16454 : 16'b0000000001111111;
														assign node16454 = (inp[1]) ? 16'b0000000000011111 : node16455;
															assign node16455 = (inp[3]) ? 16'b0000000000111111 : node16456;
																assign node16456 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node16461 = (inp[1]) ? node16469 : node16462;
													assign node16462 = (inp[10]) ? node16464 : 16'b0000000000111111;
														assign node16464 = (inp[15]) ? 16'b0000000000011111 : node16465;
															assign node16465 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node16469 = (inp[10]) ? node16473 : node16470;
														assign node16470 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node16473 = (inp[11]) ? node16475 : 16'b0000000000011111;
															assign node16475 = (inp[3]) ? 16'b0000000000001111 : 16'b0000000000011111;
									assign node16478 = (inp[4]) ? node16526 : node16479;
										assign node16479 = (inp[10]) ? node16505 : node16480;
											assign node16480 = (inp[15]) ? node16490 : node16481;
												assign node16481 = (inp[11]) ? node16485 : node16482;
													assign node16482 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000111111111;
													assign node16485 = (inp[2]) ? node16487 : 16'b0000000001111111;
														assign node16487 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node16490 = (inp[2]) ? node16498 : node16491;
													assign node16491 = (inp[3]) ? node16493 : 16'b0000000011111111;
														assign node16493 = (inp[6]) ? 16'b0000000000111111 : node16494;
															assign node16494 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node16498 = (inp[3]) ? node16500 : 16'b0000000000111111;
														assign node16500 = (inp[1]) ? node16502 : 16'b0000000000111111;
															assign node16502 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node16505 = (inp[11]) ? node16517 : node16506;
												assign node16506 = (inp[1]) ? node16514 : node16507;
													assign node16507 = (inp[6]) ? node16509 : 16'b0000000001111111;
														assign node16509 = (inp[2]) ? 16'b0000000000111111 : node16510;
															assign node16510 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node16514 = (inp[6]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node16517 = (inp[2]) ? node16519 : 16'b0000000000111111;
													assign node16519 = (inp[1]) ? node16523 : node16520;
														assign node16520 = (inp[6]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node16523 = (inp[3]) ? 16'b0000000000001111 : 16'b0000000000011111;
										assign node16526 = (inp[2]) ? node16540 : node16527;
											assign node16527 = (inp[6]) ? node16537 : node16528;
												assign node16528 = (inp[15]) ? node16534 : node16529;
													assign node16529 = (inp[1]) ? 16'b0000000001111111 : node16530;
														assign node16530 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node16534 = (inp[1]) ? 16'b0000000000001111 : 16'b0000000000111111;
												assign node16537 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node16540 = (inp[3]) ? node16556 : node16541;
												assign node16541 = (inp[15]) ? node16549 : node16542;
													assign node16542 = (inp[6]) ? 16'b0000000000011111 : node16543;
														assign node16543 = (inp[11]) ? node16545 : 16'b0000000000111111;
															assign node16545 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node16549 = (inp[11]) ? node16551 : 16'b0000000000011111;
														assign node16551 = (inp[6]) ? 16'b0000000000001111 : node16552;
															assign node16552 = (inp[10]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node16556 = (inp[1]) ? 16'b0000000000001111 : 16'b0000000000011111;
					assign node16559 = (inp[10]) ? node17331 : node16560;
						assign node16560 = (inp[3]) ? node16938 : node16561;
							assign node16561 = (inp[11]) ? node16739 : node16562;
								assign node16562 = (inp[5]) ? node16666 : node16563;
									assign node16563 = (inp[14]) ? node16617 : node16564;
										assign node16564 = (inp[2]) ? node16592 : node16565;
											assign node16565 = (inp[1]) ? node16579 : node16566;
												assign node16566 = (inp[4]) ? node16576 : node16567;
													assign node16567 = (inp[9]) ? 16'b0000011111111111 : node16568;
														assign node16568 = (inp[15]) ? node16570 : 16'b0000111111111111;
															assign node16570 = (inp[6]) ? 16'b0000011111111111 : node16571;
																assign node16571 = (inp[8]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node16576 = (inp[6]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node16579 = (inp[6]) ? node16585 : node16580;
													assign node16580 = (inp[4]) ? 16'b0000001111111111 : node16581;
														assign node16581 = (inp[8]) ? 16'b0000001111111111 : 16'b0000111111111111;
													assign node16585 = (inp[4]) ? node16587 : 16'b0000001111111111;
														assign node16587 = (inp[15]) ? node16589 : 16'b0000000111111111;
															assign node16589 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node16592 = (inp[15]) ? node16602 : node16593;
												assign node16593 = (inp[8]) ? 16'b0000000111111111 : node16594;
													assign node16594 = (inp[9]) ? node16596 : 16'b0000011111111111;
														assign node16596 = (inp[6]) ? 16'b0000001111111111 : node16597;
															assign node16597 = (inp[4]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node16602 = (inp[8]) ? node16612 : node16603;
													assign node16603 = (inp[4]) ? node16609 : node16604;
														assign node16604 = (inp[1]) ? 16'b0000000111111111 : node16605;
															assign node16605 = (inp[6]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node16609 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node16612 = (inp[6]) ? 16'b0000000011111111 : node16613;
														assign node16613 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node16617 = (inp[2]) ? node16649 : node16618;
											assign node16618 = (inp[1]) ? node16636 : node16619;
												assign node16619 = (inp[4]) ? node16631 : node16620;
													assign node16620 = (inp[15]) ? node16624 : node16621;
														assign node16621 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node16624 = (inp[8]) ? node16626 : 16'b0000001111111111;
															assign node16626 = (inp[6]) ? 16'b0000000111111111 : node16627;
																assign node16627 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node16631 = (inp[9]) ? 16'b0000000111111111 : node16632;
														assign node16632 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node16636 = (inp[6]) ? node16646 : node16637;
													assign node16637 = (inp[8]) ? node16639 : 16'b0000000111111111;
														assign node16639 = (inp[4]) ? 16'b0000000011111111 : node16640;
															assign node16640 = (inp[9]) ? node16642 : 16'b0000000111111111;
																assign node16642 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node16646 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node16649 = (inp[15]) ? node16655 : node16650;
												assign node16650 = (inp[4]) ? 16'b0000000011111111 : node16651;
													assign node16651 = (inp[6]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node16655 = (inp[1]) ? 16'b0000000001111111 : node16656;
													assign node16656 = (inp[4]) ? node16658 : 16'b0000000011111111;
														assign node16658 = (inp[8]) ? 16'b0000000001111111 : node16659;
															assign node16659 = (inp[6]) ? node16661 : 16'b0000000111111111;
																assign node16661 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node16666 = (inp[6]) ? node16700 : node16667;
										assign node16667 = (inp[1]) ? node16679 : node16668;
											assign node16668 = (inp[14]) ? 16'b0000000111111111 : node16669;
												assign node16669 = (inp[15]) ? node16673 : node16670;
													assign node16670 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node16673 = (inp[4]) ? 16'b0000000111111111 : node16674;
														assign node16674 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node16679 = (inp[15]) ? node16683 : node16680;
												assign node16680 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node16683 = (inp[14]) ? node16697 : node16684;
													assign node16684 = (inp[4]) ? node16692 : node16685;
														assign node16685 = (inp[9]) ? 16'b0000000011111111 : node16686;
															assign node16686 = (inp[8]) ? node16688 : 16'b0000000111111111;
																assign node16688 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node16692 = (inp[9]) ? 16'b0000000001111111 : node16693;
															assign node16693 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node16697 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node16700 = (inp[9]) ? node16724 : node16701;
											assign node16701 = (inp[1]) ? node16711 : node16702;
												assign node16702 = (inp[2]) ? 16'b0000000011111111 : node16703;
													assign node16703 = (inp[15]) ? node16707 : node16704;
														assign node16704 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node16707 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node16711 = (inp[4]) ? node16719 : node16712;
													assign node16712 = (inp[8]) ? node16716 : node16713;
														assign node16713 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node16716 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000011111111;
													assign node16719 = (inp[8]) ? 16'b0000000001111111 : node16720;
														assign node16720 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000001111111;
											assign node16724 = (inp[15]) ? node16732 : node16725;
												assign node16725 = (inp[8]) ? 16'b0000000001111111 : node16726;
													assign node16726 = (inp[4]) ? node16728 : 16'b0000000011111111;
														assign node16728 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000001111111;
												assign node16732 = (inp[4]) ? node16736 : node16733;
													assign node16733 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node16736 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
								assign node16739 = (inp[2]) ? node16835 : node16740;
									assign node16740 = (inp[8]) ? node16790 : node16741;
										assign node16741 = (inp[4]) ? node16767 : node16742;
											assign node16742 = (inp[14]) ? node16756 : node16743;
												assign node16743 = (inp[5]) ? 16'b0000000111111111 : node16744;
													assign node16744 = (inp[15]) ? node16750 : node16745;
														assign node16745 = (inp[9]) ? node16747 : 16'b0000011111111111;
															assign node16747 = (inp[1]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node16750 = (inp[1]) ? node16752 : 16'b0000001111111111;
															assign node16752 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node16756 = (inp[5]) ? node16762 : node16757;
													assign node16757 = (inp[15]) ? node16759 : 16'b0000001111111111;
														assign node16759 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node16762 = (inp[6]) ? node16764 : 16'b0000000011111111;
														assign node16764 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000111111111;
											assign node16767 = (inp[15]) ? node16783 : node16768;
												assign node16768 = (inp[1]) ? node16776 : node16769;
													assign node16769 = (inp[6]) ? node16773 : node16770;
														assign node16770 = (inp[9]) ? 16'b0000000011111111 : 16'b0000001111111111;
														assign node16773 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node16776 = (inp[5]) ? node16780 : node16777;
														assign node16777 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node16780 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node16783 = (inp[14]) ? 16'b0000000001111111 : node16784;
													assign node16784 = (inp[1]) ? 16'b0000000011111111 : node16785;
														assign node16785 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node16790 = (inp[1]) ? node16814 : node16791;
											assign node16791 = (inp[14]) ? node16801 : node16792;
												assign node16792 = (inp[9]) ? node16798 : node16793;
													assign node16793 = (inp[4]) ? 16'b0000000111111111 : node16794;
														assign node16794 = (inp[6]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node16798 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000111111111;
												assign node16801 = (inp[5]) ? node16807 : node16802;
													assign node16802 = (inp[4]) ? node16804 : 16'b0000000111111111;
														assign node16804 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node16807 = (inp[9]) ? node16811 : node16808;
														assign node16808 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node16811 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node16814 = (inp[5]) ? node16828 : node16815;
												assign node16815 = (inp[9]) ? node16825 : node16816;
													assign node16816 = (inp[15]) ? node16818 : 16'b0000000011111111;
														assign node16818 = (inp[14]) ? node16820 : 16'b0000000011111111;
															assign node16820 = (inp[4]) ? 16'b0000000001111111 : node16821;
																assign node16821 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node16825 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000001111111;
												assign node16828 = (inp[14]) ? node16830 : 16'b0000000001111111;
													assign node16830 = (inp[6]) ? 16'b0000000000111111 : node16831;
														assign node16831 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node16835 = (inp[1]) ? node16881 : node16836;
										assign node16836 = (inp[15]) ? node16864 : node16837;
											assign node16837 = (inp[8]) ? node16849 : node16838;
												assign node16838 = (inp[4]) ? node16844 : node16839;
													assign node16839 = (inp[14]) ? node16841 : 16'b0000001111111111;
														assign node16841 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node16844 = (inp[9]) ? 16'b0000000011111111 : node16845;
														assign node16845 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node16849 = (inp[14]) ? node16859 : node16850;
													assign node16850 = (inp[4]) ? node16854 : node16851;
														assign node16851 = (inp[6]) ? 16'b0000000111111111 : 16'b0000000011111111;
														assign node16854 = (inp[6]) ? node16856 : 16'b0000000011111111;
															assign node16856 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node16859 = (inp[5]) ? 16'b0000000001111111 : node16860;
														assign node16860 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000111111111;
											assign node16864 = (inp[14]) ? node16868 : node16865;
												assign node16865 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node16868 = (inp[8]) ? node16876 : node16869;
													assign node16869 = (inp[4]) ? node16871 : 16'b0000000001111111;
														assign node16871 = (inp[6]) ? node16873 : 16'b0000000001111111;
															assign node16873 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node16876 = (inp[6]) ? 16'b0000000000111111 : node16877;
														assign node16877 = (inp[4]) ? 16'b0000000000011111 : 16'b0000000001111111;
										assign node16881 = (inp[6]) ? node16909 : node16882;
											assign node16882 = (inp[14]) ? node16890 : node16883;
												assign node16883 = (inp[9]) ? 16'b0000000000111111 : node16884;
													assign node16884 = (inp[15]) ? 16'b0000000011111111 : node16885;
														assign node16885 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node16890 = (inp[4]) ? node16902 : node16891;
													assign node16891 = (inp[15]) ? node16895 : node16892;
														assign node16892 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node16895 = (inp[5]) ? node16897 : 16'b0000000001111111;
															assign node16897 = (inp[9]) ? 16'b0000000000111111 : node16898;
																assign node16898 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node16902 = (inp[15]) ? node16904 : 16'b0000000000111111;
														assign node16904 = (inp[9]) ? 16'b0000000000011111 : node16905;
															assign node16905 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node16909 = (inp[15]) ? node16923 : node16910;
												assign node16910 = (inp[4]) ? node16916 : node16911;
													assign node16911 = (inp[8]) ? 16'b0000000000111111 : node16912;
														assign node16912 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node16916 = (inp[9]) ? 16'b0000000000011111 : node16917;
														assign node16917 = (inp[14]) ? 16'b0000000000111111 : node16918;
															assign node16918 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node16923 = (inp[8]) ? node16929 : node16924;
													assign node16924 = (inp[4]) ? node16926 : 16'b0000000000111111;
														assign node16926 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node16929 = (inp[5]) ? node16931 : 16'b0000000000011111;
														assign node16931 = (inp[9]) ? 16'b0000000000001111 : node16932;
															assign node16932 = (inp[14]) ? node16934 : 16'b0000000000011111;
																assign node16934 = (inp[4]) ? 16'b0000000000001111 : 16'b0000000000011111;
							assign node16938 = (inp[14]) ? node17150 : node16939;
								assign node16939 = (inp[11]) ? node17047 : node16940;
									assign node16940 = (inp[15]) ? node16984 : node16941;
										assign node16941 = (inp[4]) ? node16961 : node16942;
											assign node16942 = (inp[1]) ? node16950 : node16943;
												assign node16943 = (inp[8]) ? 16'b0000000111111111 : node16944;
													assign node16944 = (inp[5]) ? 16'b0000001111111111 : node16945;
														assign node16945 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node16950 = (inp[6]) ? node16956 : node16951;
													assign node16951 = (inp[5]) ? 16'b0000000111111111 : node16952;
														assign node16952 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node16956 = (inp[5]) ? 16'b0000000011111111 : node16957;
														assign node16957 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node16961 = (inp[2]) ? node16973 : node16962;
												assign node16962 = (inp[9]) ? node16968 : node16963;
													assign node16963 = (inp[6]) ? node16965 : 16'b0000001111111111;
														assign node16965 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node16968 = (inp[1]) ? 16'b0000000011111111 : node16969;
														assign node16969 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node16973 = (inp[1]) ? node16981 : node16974;
													assign node16974 = (inp[9]) ? node16978 : node16975;
														assign node16975 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node16978 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node16981 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000000111111;
										assign node16984 = (inp[8]) ? node17010 : node16985;
											assign node16985 = (inp[5]) ? node17001 : node16986;
												assign node16986 = (inp[4]) ? node16990 : node16987;
													assign node16987 = (inp[6]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node16990 = (inp[2]) ? node16998 : node16991;
														assign node16991 = (inp[1]) ? 16'b0000000011111111 : node16992;
															assign node16992 = (inp[9]) ? node16994 : 16'b0000000111111111;
																assign node16994 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node16998 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node17001 = (inp[1]) ? node17005 : node17002;
													assign node17002 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node17005 = (inp[6]) ? 16'b0000000001111111 : node17006;
														assign node17006 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node17010 = (inp[1]) ? node17034 : node17011;
												assign node17011 = (inp[9]) ? node17025 : node17012;
													assign node17012 = (inp[5]) ? node17018 : node17013;
														assign node17013 = (inp[2]) ? 16'b0000000011111111 : node17014;
															assign node17014 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node17018 = (inp[2]) ? node17020 : 16'b0000000011111111;
															assign node17020 = (inp[6]) ? 16'b0000000001111111 : node17021;
																assign node17021 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node17025 = (inp[5]) ? node17029 : node17026;
														assign node17026 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node17029 = (inp[4]) ? node17031 : 16'b0000000001111111;
															assign node17031 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node17034 = (inp[4]) ? node17044 : node17035;
													assign node17035 = (inp[5]) ? node17039 : node17036;
														assign node17036 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node17039 = (inp[2]) ? 16'b0000000000111111 : node17040;
															assign node17040 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node17044 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node17047 = (inp[9]) ? node17097 : node17048;
										assign node17048 = (inp[2]) ? node17072 : node17049;
											assign node17049 = (inp[15]) ? node17065 : node17050;
												assign node17050 = (inp[1]) ? node17056 : node17051;
													assign node17051 = (inp[5]) ? 16'b0000000111111111 : node17052;
														assign node17052 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node17056 = (inp[4]) ? node17058 : 16'b0000000111111111;
														assign node17058 = (inp[5]) ? 16'b0000000001111111 : node17059;
															assign node17059 = (inp[8]) ? node17061 : 16'b0000000011111111;
																assign node17061 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node17065 = (inp[1]) ? 16'b0000000001111111 : node17066;
													assign node17066 = (inp[4]) ? node17068 : 16'b0000000011111111;
														assign node17068 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000011111111;
											assign node17072 = (inp[4]) ? node17090 : node17073;
												assign node17073 = (inp[1]) ? node17081 : node17074;
													assign node17074 = (inp[8]) ? node17078 : node17075;
														assign node17075 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node17078 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node17081 = (inp[5]) ? node17087 : node17082;
														assign node17082 = (inp[15]) ? 16'b0000000001111111 : node17083;
															assign node17083 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node17087 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000000111111;
												assign node17090 = (inp[5]) ? 16'b0000000000111111 : node17091;
													assign node17091 = (inp[8]) ? node17093 : 16'b0000000001111111;
														assign node17093 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node17097 = (inp[15]) ? node17123 : node17098;
											assign node17098 = (inp[4]) ? node17114 : node17099;
												assign node17099 = (inp[2]) ? node17107 : node17100;
													assign node17100 = (inp[1]) ? node17104 : node17101;
														assign node17101 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node17104 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node17107 = (inp[5]) ? 16'b0000000001111111 : node17108;
														assign node17108 = (inp[6]) ? node17110 : 16'b0000000011111111;
															assign node17110 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node17114 = (inp[5]) ? node17118 : node17115;
													assign node17115 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node17118 = (inp[1]) ? node17120 : 16'b0000000000111111;
														assign node17120 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node17123 = (inp[6]) ? node17135 : node17124;
												assign node17124 = (inp[2]) ? node17130 : node17125;
													assign node17125 = (inp[8]) ? node17127 : 16'b0000000011111111;
														assign node17127 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node17130 = (inp[8]) ? 16'b0000000000111111 : node17131;
														assign node17131 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node17135 = (inp[8]) ? node17139 : node17136;
													assign node17136 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node17139 = (inp[4]) ? node17145 : node17140;
														assign node17140 = (inp[5]) ? 16'b0000000000011111 : node17141;
															assign node17141 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node17145 = (inp[1]) ? node17147 : 16'b0000000000011111;
															assign node17147 = (inp[2]) ? 16'b0000000000000111 : 16'b0000000000001111;
								assign node17150 = (inp[8]) ? node17226 : node17151;
									assign node17151 = (inp[9]) ? node17183 : node17152;
										assign node17152 = (inp[5]) ? node17172 : node17153;
											assign node17153 = (inp[4]) ? node17165 : node17154;
												assign node17154 = (inp[6]) ? node17160 : node17155;
													assign node17155 = (inp[2]) ? node17157 : 16'b0000000111111111;
														assign node17157 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node17160 = (inp[2]) ? 16'b0000000001111111 : node17161;
														assign node17161 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node17165 = (inp[11]) ? 16'b0000000001111111 : node17166;
													assign node17166 = (inp[2]) ? node17168 : 16'b0000000011111111;
														assign node17168 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node17172 = (inp[1]) ? node17178 : node17173;
												assign node17173 = (inp[4]) ? node17175 : 16'b0000000001111111;
													assign node17175 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node17178 = (inp[11]) ? 16'b0000000000111111 : node17179;
													assign node17179 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node17183 = (inp[4]) ? node17203 : node17184;
											assign node17184 = (inp[2]) ? node17192 : node17185;
												assign node17185 = (inp[15]) ? 16'b0000000001111111 : node17186;
													assign node17186 = (inp[11]) ? 16'b0000000011111111 : node17187;
														assign node17187 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node17192 = (inp[6]) ? node17198 : node17193;
													assign node17193 = (inp[5]) ? node17195 : 16'b0000000011111111;
														assign node17195 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node17198 = (inp[11]) ? 16'b0000000000111111 : node17199;
														assign node17199 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node17203 = (inp[15]) ? node17215 : node17204;
												assign node17204 = (inp[1]) ? node17208 : node17205;
													assign node17205 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000001111111;
													assign node17208 = (inp[2]) ? node17212 : node17209;
														assign node17209 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node17212 = (inp[5]) ? 16'b0000000000001111 : 16'b0000000000111111;
												assign node17215 = (inp[1]) ? node17221 : node17216;
													assign node17216 = (inp[2]) ? node17218 : 16'b0000000000111111;
														assign node17218 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node17221 = (inp[5]) ? 16'b0000000000000111 : node17222;
														assign node17222 = (inp[6]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node17226 = (inp[5]) ? node17280 : node17227;
										assign node17227 = (inp[15]) ? node17255 : node17228;
											assign node17228 = (inp[6]) ? node17242 : node17229;
												assign node17229 = (inp[2]) ? node17239 : node17230;
													assign node17230 = (inp[4]) ? node17234 : node17231;
														assign node17231 = (inp[11]) ? 16'b0000000011111111 : 16'b0000001111111111;
														assign node17234 = (inp[9]) ? node17236 : 16'b0000000011111111;
															assign node17236 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node17239 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node17242 = (inp[9]) ? node17248 : node17243;
													assign node17243 = (inp[2]) ? node17245 : 16'b0000000001111111;
														assign node17245 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000000111111;
													assign node17248 = (inp[2]) ? node17250 : 16'b0000000000111111;
														assign node17250 = (inp[4]) ? node17252 : 16'b0000000000111111;
															assign node17252 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node17255 = (inp[11]) ? node17265 : node17256;
												assign node17256 = (inp[2]) ? node17258 : 16'b0000000001111111;
													assign node17258 = (inp[1]) ? node17262 : node17259;
														assign node17259 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node17262 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node17265 = (inp[1]) ? node17271 : node17266;
													assign node17266 = (inp[9]) ? node17268 : 16'b0000000000111111;
														assign node17268 = (inp[6]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node17271 = (inp[6]) ? node17277 : node17272;
														assign node17272 = (inp[9]) ? node17274 : 16'b0000000000011111;
															assign node17274 = (inp[4]) ? 16'b0000000000001111 : 16'b0000000000011111;
														assign node17277 = (inp[2]) ? 16'b0000000000000111 : 16'b0000000000001111;
										assign node17280 = (inp[11]) ? node17310 : node17281;
											assign node17281 = (inp[1]) ? node17295 : node17282;
												assign node17282 = (inp[2]) ? node17290 : node17283;
													assign node17283 = (inp[6]) ? node17285 : 16'b0000000001111111;
														assign node17285 = (inp[4]) ? 16'b0000000000111111 : node17286;
															assign node17286 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node17290 = (inp[4]) ? node17292 : 16'b0000000000111111;
														assign node17292 = (inp[6]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node17295 = (inp[9]) ? node17305 : node17296;
													assign node17296 = (inp[6]) ? 16'b0000000000011111 : node17297;
														assign node17297 = (inp[4]) ? node17299 : 16'b0000000000111111;
															assign node17299 = (inp[2]) ? node17301 : 16'b0000000000111111;
																assign node17301 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node17305 = (inp[15]) ? 16'b0000000000001111 : node17306;
														assign node17306 = (inp[4]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node17310 = (inp[6]) ? node17316 : node17311;
												assign node17311 = (inp[1]) ? 16'b0000000000011111 : node17312;
													assign node17312 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node17316 = (inp[4]) ? node17318 : 16'b0000000000111111;
													assign node17318 = (inp[15]) ? node17324 : node17319;
														assign node17319 = (inp[2]) ? 16'b0000000000001111 : node17320;
															assign node17320 = (inp[1]) ? 16'b0000000000001111 : 16'b0000000000011111;
														assign node17324 = (inp[9]) ? node17326 : 16'b0000000000001111;
															assign node17326 = (inp[2]) ? 16'b0000000000000111 : node17327;
																assign node17327 = (inp[1]) ? 16'b0000000000000111 : 16'b0000000000001111;
						assign node17331 = (inp[9]) ? node17709 : node17332;
							assign node17332 = (inp[2]) ? node17504 : node17333;
								assign node17333 = (inp[8]) ? node17417 : node17334;
									assign node17334 = (inp[15]) ? node17374 : node17335;
										assign node17335 = (inp[11]) ? node17353 : node17336;
											assign node17336 = (inp[5]) ? node17350 : node17337;
												assign node17337 = (inp[1]) ? node17343 : node17338;
													assign node17338 = (inp[14]) ? 16'b0000000111111111 : node17339;
														assign node17339 = (inp[6]) ? 16'b0000011111111111 : 16'b0000001111111111;
													assign node17343 = (inp[14]) ? node17345 : 16'b0000000111111111;
														assign node17345 = (inp[3]) ? 16'b0000000111111111 : node17346;
															assign node17346 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node17350 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node17353 = (inp[5]) ? node17367 : node17354;
												assign node17354 = (inp[6]) ? node17362 : node17355;
													assign node17355 = (inp[4]) ? node17359 : node17356;
														assign node17356 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node17359 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node17362 = (inp[3]) ? 16'b0000000011111111 : node17363;
														assign node17363 = (inp[1]) ? 16'b0000000111111111 : 16'b0000000011111111;
												assign node17367 = (inp[14]) ? 16'b0000000000011111 : node17368;
													assign node17368 = (inp[3]) ? node17370 : 16'b0000000011111111;
														assign node17370 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node17374 = (inp[11]) ? node17404 : node17375;
											assign node17375 = (inp[6]) ? node17393 : node17376;
												assign node17376 = (inp[3]) ? node17384 : node17377;
													assign node17377 = (inp[1]) ? node17381 : node17378;
														assign node17378 = (inp[4]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node17381 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node17384 = (inp[1]) ? node17388 : node17385;
														assign node17385 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node17388 = (inp[14]) ? node17390 : 16'b0000000011111111;
															assign node17390 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node17393 = (inp[3]) ? node17399 : node17394;
													assign node17394 = (inp[14]) ? node17396 : 16'b0000000011111111;
														assign node17396 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node17399 = (inp[4]) ? node17401 : 16'b0000000001111111;
														assign node17401 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node17404 = (inp[4]) ? node17408 : node17405;
												assign node17405 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000001111111;
												assign node17408 = (inp[14]) ? node17410 : 16'b0000000001111111;
													assign node17410 = (inp[6]) ? node17412 : 16'b0000000000011111;
														assign node17412 = (inp[1]) ? node17414 : 16'b0000000000111111;
															assign node17414 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node17417 = (inp[1]) ? node17455 : node17418;
										assign node17418 = (inp[11]) ? node17438 : node17419;
											assign node17419 = (inp[3]) ? node17427 : node17420;
												assign node17420 = (inp[5]) ? node17424 : node17421;
													assign node17421 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node17424 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node17427 = (inp[14]) ? node17431 : node17428;
													assign node17428 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node17431 = (inp[4]) ? node17433 : 16'b0000000011111111;
														assign node17433 = (inp[6]) ? 16'b0000000001111111 : node17434;
															assign node17434 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node17438 = (inp[14]) ? node17448 : node17439;
												assign node17439 = (inp[5]) ? node17441 : 16'b0000000011111111;
													assign node17441 = (inp[3]) ? node17445 : node17442;
														assign node17442 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node17445 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node17448 = (inp[15]) ? node17452 : node17449;
													assign node17449 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000011111111;
													assign node17452 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node17455 = (inp[3]) ? node17481 : node17456;
											assign node17456 = (inp[6]) ? node17470 : node17457;
												assign node17457 = (inp[4]) ? node17463 : node17458;
													assign node17458 = (inp[14]) ? node17460 : 16'b0000000011111111;
														assign node17460 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000001111111;
													assign node17463 = (inp[15]) ? 16'b0000000001111111 : node17464;
														assign node17464 = (inp[14]) ? 16'b0000000001111111 : node17465;
															assign node17465 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node17470 = (inp[14]) ? 16'b0000000000111111 : node17471;
													assign node17471 = (inp[15]) ? 16'b0000000000111111 : node17472;
														assign node17472 = (inp[4]) ? 16'b0000000001111111 : node17473;
															assign node17473 = (inp[5]) ? node17475 : 16'b0000000011111111;
																assign node17475 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node17481 = (inp[4]) ? node17493 : node17482;
												assign node17482 = (inp[14]) ? node17488 : node17483;
													assign node17483 = (inp[15]) ? 16'b0000000001111111 : node17484;
														assign node17484 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000001111111;
													assign node17488 = (inp[6]) ? node17490 : 16'b0000000000111111;
														assign node17490 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node17493 = (inp[5]) ? node17495 : 16'b0000000000111111;
													assign node17495 = (inp[11]) ? node17499 : node17496;
														assign node17496 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000000011111;
														assign node17499 = (inp[6]) ? node17501 : 16'b0000000000011111;
															assign node17501 = (inp[14]) ? 16'b0000000000001111 : 16'b0000000000011111;
								assign node17504 = (inp[15]) ? node17604 : node17505;
									assign node17505 = (inp[6]) ? node17561 : node17506;
										assign node17506 = (inp[3]) ? node17530 : node17507;
											assign node17507 = (inp[8]) ? node17519 : node17508;
												assign node17508 = (inp[1]) ? node17514 : node17509;
													assign node17509 = (inp[5]) ? node17511 : 16'b0000000111111111;
														assign node17511 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node17514 = (inp[5]) ? 16'b0000000001111111 : node17515;
														assign node17515 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000111111111;
												assign node17519 = (inp[14]) ? node17525 : node17520;
													assign node17520 = (inp[11]) ? 16'b0000000001111111 : node17521;
														assign node17521 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node17525 = (inp[4]) ? node17527 : 16'b0000000001111111;
														assign node17527 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node17530 = (inp[4]) ? node17548 : node17531;
												assign node17531 = (inp[14]) ? node17539 : node17532;
													assign node17532 = (inp[8]) ? node17536 : node17533;
														assign node17533 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node17536 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node17539 = (inp[1]) ? 16'b0000000001111111 : node17540;
														assign node17540 = (inp[11]) ? 16'b0000000001111111 : node17541;
															assign node17541 = (inp[8]) ? node17543 : 16'b0000000011111111;
																assign node17543 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node17548 = (inp[11]) ? node17558 : node17549;
													assign node17549 = (inp[1]) ? node17551 : 16'b0000000011111111;
														assign node17551 = (inp[8]) ? 16'b0000000000011111 : node17552;
															assign node17552 = (inp[5]) ? node17554 : 16'b0000000001111111;
																assign node17554 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node17558 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node17561 = (inp[8]) ? node17583 : node17562;
											assign node17562 = (inp[14]) ? node17572 : node17563;
												assign node17563 = (inp[4]) ? 16'b0000000001111111 : node17564;
													assign node17564 = (inp[1]) ? node17566 : 16'b0000000011111111;
														assign node17566 = (inp[5]) ? 16'b0000000001111111 : node17567;
															assign node17567 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node17572 = (inp[1]) ? node17580 : node17573;
													assign node17573 = (inp[3]) ? node17577 : node17574;
														assign node17574 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node17577 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node17580 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node17583 = (inp[5]) ? node17593 : node17584;
												assign node17584 = (inp[14]) ? node17590 : node17585;
													assign node17585 = (inp[4]) ? node17587 : 16'b0000000001111111;
														assign node17587 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node17590 = (inp[4]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node17593 = (inp[4]) ? node17597 : node17594;
													assign node17594 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node17597 = (inp[3]) ? node17599 : 16'b0000000000111111;
														assign node17599 = (inp[14]) ? node17601 : 16'b0000000000011111;
															assign node17601 = (inp[1]) ? 16'b0000000000001111 : 16'b0000000000011111;
									assign node17604 = (inp[4]) ? node17654 : node17605;
										assign node17605 = (inp[6]) ? node17629 : node17606;
											assign node17606 = (inp[3]) ? node17620 : node17607;
												assign node17607 = (inp[1]) ? node17613 : node17608;
													assign node17608 = (inp[14]) ? 16'b0000000011111111 : node17609;
														assign node17609 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node17613 = (inp[14]) ? node17617 : node17614;
														assign node17614 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000001111111;
														assign node17617 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node17620 = (inp[14]) ? 16'b0000000000111111 : node17621;
													assign node17621 = (inp[5]) ? node17623 : 16'b0000000011111111;
														assign node17623 = (inp[8]) ? node17625 : 16'b0000000001111111;
															assign node17625 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node17629 = (inp[1]) ? node17643 : node17630;
												assign node17630 = (inp[8]) ? node17638 : node17631;
													assign node17631 = (inp[14]) ? 16'b0000000000011111 : node17632;
														assign node17632 = (inp[5]) ? 16'b0000000001111111 : node17633;
															assign node17633 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node17638 = (inp[11]) ? 16'b0000000000111111 : node17639;
														assign node17639 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node17643 = (inp[3]) ? node17649 : node17644;
													assign node17644 = (inp[8]) ? node17646 : 16'b0000000000111111;
														assign node17646 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node17649 = (inp[14]) ? node17651 : 16'b0000000000011111;
														assign node17651 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node17654 = (inp[11]) ? node17678 : node17655;
											assign node17655 = (inp[1]) ? node17663 : node17656;
												assign node17656 = (inp[5]) ? 16'b0000000000111111 : node17657;
													assign node17657 = (inp[8]) ? 16'b0000000001111111 : node17658;
														assign node17658 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000111111111;
												assign node17663 = (inp[6]) ? node17671 : node17664;
													assign node17664 = (inp[3]) ? node17668 : node17665;
														assign node17665 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node17668 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node17671 = (inp[14]) ? node17675 : node17672;
														assign node17672 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000000011111;
														assign node17675 = (inp[8]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node17678 = (inp[6]) ? node17698 : node17679;
												assign node17679 = (inp[3]) ? node17687 : node17680;
													assign node17680 = (inp[1]) ? node17684 : node17681;
														assign node17681 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node17684 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node17687 = (inp[1]) ? node17691 : node17688;
														assign node17688 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node17691 = (inp[14]) ? 16'b0000000000001111 : node17692;
															assign node17692 = (inp[8]) ? node17694 : 16'b0000000000011111;
																assign node17694 = (inp[5]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node17698 = (inp[8]) ? node17704 : node17699;
													assign node17699 = (inp[1]) ? node17701 : 16'b0000000000011111;
														assign node17701 = (inp[3]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node17704 = (inp[3]) ? node17706 : 16'b0000000000001111;
														assign node17706 = (inp[1]) ? 16'b0000000000000011 : 16'b0000000000000111;
							assign node17709 = (inp[8]) ? node17903 : node17710;
								assign node17710 = (inp[15]) ? node17794 : node17711;
									assign node17711 = (inp[1]) ? node17759 : node17712;
										assign node17712 = (inp[14]) ? node17740 : node17713;
											assign node17713 = (inp[11]) ? node17729 : node17714;
												assign node17714 = (inp[6]) ? node17720 : node17715;
													assign node17715 = (inp[2]) ? node17717 : 16'b0000000111111111;
														assign node17717 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node17720 = (inp[4]) ? node17724 : node17721;
														assign node17721 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node17724 = (inp[3]) ? node17726 : 16'b0000000011111111;
															assign node17726 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node17729 = (inp[3]) ? node17735 : node17730;
													assign node17730 = (inp[6]) ? 16'b0000000001111111 : node17731;
														assign node17731 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node17735 = (inp[2]) ? node17737 : 16'b0000000001111111;
														assign node17737 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node17740 = (inp[4]) ? node17746 : node17741;
												assign node17741 = (inp[11]) ? 16'b0000000001111111 : node17742;
													assign node17742 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node17746 = (inp[5]) ? 16'b0000000000111111 : node17747;
													assign node17747 = (inp[11]) ? node17751 : node17748;
														assign node17748 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node17751 = (inp[3]) ? node17753 : 16'b0000000001111111;
															assign node17753 = (inp[6]) ? 16'b0000000000111111 : node17754;
																assign node17754 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node17759 = (inp[11]) ? node17785 : node17760;
											assign node17760 = (inp[14]) ? node17770 : node17761;
												assign node17761 = (inp[5]) ? node17765 : node17762;
													assign node17762 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node17765 = (inp[3]) ? node17767 : 16'b0000000001111111;
														assign node17767 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node17770 = (inp[2]) ? node17776 : node17771;
													assign node17771 = (inp[5]) ? node17773 : 16'b0000000011111111;
														assign node17773 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node17776 = (inp[4]) ? node17780 : node17777;
														assign node17777 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node17780 = (inp[5]) ? 16'b0000000000111111 : node17781;
															assign node17781 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node17785 = (inp[14]) ? node17787 : 16'b0000000000111111;
												assign node17787 = (inp[5]) ? node17791 : node17788;
													assign node17788 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node17791 = (inp[4]) ? 16'b0000000000001111 : 16'b0000000000011111;
									assign node17794 = (inp[2]) ? node17844 : node17795;
										assign node17795 = (inp[4]) ? node17817 : node17796;
											assign node17796 = (inp[6]) ? node17806 : node17797;
												assign node17797 = (inp[3]) ? node17801 : node17798;
													assign node17798 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node17801 = (inp[1]) ? 16'b0000000000111111 : node17802;
														assign node17802 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node17806 = (inp[11]) ? node17810 : node17807;
													assign node17807 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000001111111;
													assign node17810 = (inp[14]) ? 16'b0000000000011111 : node17811;
														assign node17811 = (inp[5]) ? node17813 : 16'b0000000001111111;
															assign node17813 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node17817 = (inp[3]) ? node17833 : node17818;
												assign node17818 = (inp[6]) ? node17828 : node17819;
													assign node17819 = (inp[14]) ? node17823 : node17820;
														assign node17820 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node17823 = (inp[1]) ? node17825 : 16'b0000000001111111;
															assign node17825 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node17828 = (inp[5]) ? node17830 : 16'b0000000000111111;
														assign node17830 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node17833 = (inp[5]) ? 16'b0000000000011111 : node17834;
													assign node17834 = (inp[14]) ? node17840 : node17835;
														assign node17835 = (inp[1]) ? 16'b0000000000111111 : node17836;
															assign node17836 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node17840 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node17844 = (inp[6]) ? node17868 : node17845;
											assign node17845 = (inp[3]) ? node17859 : node17846;
												assign node17846 = (inp[5]) ? node17848 : 16'b0000000001111111;
													assign node17848 = (inp[11]) ? node17856 : node17849;
														assign node17849 = (inp[1]) ? 16'b0000000000011111 : node17850;
															assign node17850 = (inp[4]) ? 16'b0000000001111111 : node17851;
																assign node17851 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node17856 = (inp[4]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node17859 = (inp[14]) ? node17861 : 16'b0000000000111111;
													assign node17861 = (inp[5]) ? node17863 : 16'b0000000000111111;
														assign node17863 = (inp[1]) ? 16'b0000000000001111 : node17864;
															assign node17864 = (inp[11]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node17868 = (inp[1]) ? node17886 : node17869;
												assign node17869 = (inp[4]) ? node17875 : node17870;
													assign node17870 = (inp[14]) ? node17872 : 16'b0000000000111111;
														assign node17872 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node17875 = (inp[3]) ? node17879 : node17876;
														assign node17876 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000001111111;
														assign node17879 = (inp[14]) ? node17881 : 16'b0000000000011111;
															assign node17881 = (inp[5]) ? 16'b0000000000001111 : node17882;
																assign node17882 = (inp[11]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node17886 = (inp[3]) ? node17900 : node17887;
													assign node17887 = (inp[4]) ? node17897 : node17888;
														assign node17888 = (inp[5]) ? node17892 : node17889;
															assign node17889 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
															assign node17892 = (inp[14]) ? node17894 : 16'b0000000000011111;
																assign node17894 = (inp[11]) ? 16'b0000000000001111 : 16'b0000000000011111;
														assign node17897 = (inp[14]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node17900 = (inp[4]) ? 16'b0000000000001111 : 16'b0000000000000111;
								assign node17903 = (inp[6]) ? node17999 : node17904;
									assign node17904 = (inp[3]) ? node17952 : node17905;
										assign node17905 = (inp[1]) ? node17929 : node17906;
											assign node17906 = (inp[2]) ? node17924 : node17907;
												assign node17907 = (inp[11]) ? node17915 : node17908;
													assign node17908 = (inp[5]) ? 16'b0000000011111111 : node17909;
														assign node17909 = (inp[15]) ? 16'b0000000111111111 : node17910;
															assign node17910 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node17915 = (inp[4]) ? node17919 : node17916;
														assign node17916 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node17919 = (inp[5]) ? 16'b0000000001111111 : node17920;
															assign node17920 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node17924 = (inp[11]) ? node17926 : 16'b0000000001111111;
													assign node17926 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node17929 = (inp[2]) ? node17943 : node17930;
												assign node17930 = (inp[11]) ? node17936 : node17931;
													assign node17931 = (inp[14]) ? 16'b0000000000111111 : node17932;
														assign node17932 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node17936 = (inp[15]) ? node17940 : node17937;
														assign node17937 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000000111111;
														assign node17940 = (inp[4]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node17943 = (inp[15]) ? node17949 : node17944;
													assign node17944 = (inp[5]) ? node17946 : 16'b0000000000111111;
														assign node17946 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node17949 = (inp[5]) ? 16'b0000000000000111 : 16'b0000000000011111;
										assign node17952 = (inp[1]) ? node17978 : node17953;
											assign node17953 = (inp[15]) ? node17963 : node17954;
												assign node17954 = (inp[4]) ? node17960 : node17955;
													assign node17955 = (inp[11]) ? node17957 : 16'b0000000001111111;
														assign node17957 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node17960 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node17963 = (inp[5]) ? node17971 : node17964;
													assign node17964 = (inp[14]) ? node17968 : node17965;
														assign node17965 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node17968 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node17971 = (inp[14]) ? node17975 : node17972;
														assign node17972 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000000011111;
														assign node17975 = (inp[11]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node17978 = (inp[15]) ? node17992 : node17979;
												assign node17979 = (inp[4]) ? node17985 : node17980;
													assign node17980 = (inp[5]) ? node17982 : 16'b0000000001111111;
														assign node17982 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node17985 = (inp[14]) ? node17987 : 16'b0000000000011111;
														assign node17987 = (inp[11]) ? node17989 : 16'b0000000000011111;
															assign node17989 = (inp[2]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node17992 = (inp[5]) ? 16'b0000000000001111 : node17993;
													assign node17993 = (inp[4]) ? node17995 : 16'b0000000000011111;
														assign node17995 = (inp[14]) ? 16'b0000000000001111 : 16'b0000000000011111;
									assign node17999 = (inp[4]) ? node18049 : node18000;
										assign node18000 = (inp[11]) ? node18022 : node18001;
											assign node18001 = (inp[1]) ? node18009 : node18002;
												assign node18002 = (inp[5]) ? node18004 : 16'b0000000001111111;
													assign node18004 = (inp[15]) ? 16'b0000000000111111 : node18005;
														assign node18005 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node18009 = (inp[15]) ? node18017 : node18010;
													assign node18010 = (inp[3]) ? 16'b0000000000111111 : node18011;
														assign node18011 = (inp[14]) ? 16'b0000000000111111 : node18012;
															assign node18012 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node18017 = (inp[5]) ? 16'b0000000000001111 : node18018;
														assign node18018 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node18022 = (inp[5]) ? node18036 : node18023;
												assign node18023 = (inp[15]) ? node18033 : node18024;
													assign node18024 = (inp[14]) ? node18030 : node18025;
														assign node18025 = (inp[3]) ? 16'b0000000000111111 : node18026;
															assign node18026 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node18030 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node18033 = (inp[14]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node18036 = (inp[2]) ? node18042 : node18037;
													assign node18037 = (inp[1]) ? node18039 : 16'b0000000000011111;
														assign node18039 = (inp[3]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node18042 = (inp[15]) ? node18044 : 16'b0000000000001111;
														assign node18044 = (inp[1]) ? 16'b0000000000000111 : node18045;
															assign node18045 = (inp[3]) ? 16'b0000000000000111 : 16'b0000000000001111;
										assign node18049 = (inp[14]) ? node18089 : node18050;
											assign node18050 = (inp[11]) ? node18064 : node18051;
												assign node18051 = (inp[5]) ? node18057 : node18052;
													assign node18052 = (inp[15]) ? 16'b0000000000111111 : node18053;
														assign node18053 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node18057 = (inp[2]) ? node18061 : node18058;
														assign node18058 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node18061 = (inp[3]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node18064 = (inp[15]) ? node18080 : node18065;
													assign node18065 = (inp[2]) ? node18069 : node18066;
														assign node18066 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node18069 = (inp[3]) ? node18075 : node18070;
															assign node18070 = (inp[5]) ? node18072 : 16'b0000000000011111;
																assign node18072 = (inp[1]) ? 16'b0000000000001111 : 16'b0000000000011111;
															assign node18075 = (inp[1]) ? 16'b0000000000001111 : node18076;
																assign node18076 = (inp[5]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node18080 = (inp[3]) ? node18084 : node18081;
														assign node18081 = (inp[1]) ? 16'b0000000000001111 : 16'b0000000000011111;
														assign node18084 = (inp[2]) ? node18086 : 16'b0000000000001111;
															assign node18086 = (inp[5]) ? 16'b0000000000000111 : 16'b0000000000001111;
											assign node18089 = (inp[5]) ? node18105 : node18090;
												assign node18090 = (inp[1]) ? node18098 : node18091;
													assign node18091 = (inp[2]) ? node18095 : node18092;
														assign node18092 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000001111111;
														assign node18095 = (inp[3]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node18098 = (inp[11]) ? node18102 : node18099;
														assign node18099 = (inp[15]) ? 16'b0000000000001111 : 16'b0000000000011111;
														assign node18102 = (inp[3]) ? 16'b0000000000000111 : 16'b0000000000001111;
												assign node18105 = (inp[3]) ? node18111 : node18106;
													assign node18106 = (inp[1]) ? node18108 : 16'b0000000000011111;
														assign node18108 = (inp[11]) ? 16'b0000000000000111 : 16'b0000000000001111;
													assign node18111 = (inp[15]) ? node18117 : node18112;
														assign node18112 = (inp[11]) ? 16'b0000000000000111 : node18113;
															assign node18113 = (inp[1]) ? 16'b0000000000000111 : 16'b0000000000001111;
														assign node18117 = (inp[11]) ? node18121 : node18118;
															assign node18118 = (inp[1]) ? 16'b0000000000000011 : 16'b0000000000000111;
															assign node18121 = (inp[1]) ? 16'b0000000000000001 : 16'b0000000000000011;
			assign node18124 = (inp[8]) ? node21132 : node18125;
				assign node18125 = (inp[5]) ? node19643 : node18126;
					assign node18126 = (inp[13]) ? node18866 : node18127;
						assign node18127 = (inp[15]) ? node18527 : node18128;
							assign node18128 = (inp[6]) ? node18312 : node18129;
								assign node18129 = (inp[14]) ? node18219 : node18130;
									assign node18130 = (inp[11]) ? node18176 : node18131;
										assign node18131 = (inp[10]) ? node18159 : node18132;
											assign node18132 = (inp[12]) ? node18142 : node18133;
												assign node18133 = (inp[3]) ? node18139 : node18134;
													assign node18134 = (inp[4]) ? 16'b0000111111111111 : node18135;
														assign node18135 = (inp[2]) ? 16'b0000111111111111 : 16'b0001111111111111;
													assign node18139 = (inp[1]) ? 16'b0000111111111111 : 16'b0000011111111111;
												assign node18142 = (inp[4]) ? node18152 : node18143;
													assign node18143 = (inp[2]) ? 16'b0000011111111111 : node18144;
														assign node18144 = (inp[1]) ? 16'b0000011111111111 : node18145;
															assign node18145 = (inp[3]) ? 16'b0000111111111111 : node18146;
																assign node18146 = (inp[9]) ? 16'b0000111111111111 : 16'b0001111111111111;
													assign node18152 = (inp[9]) ? 16'b0000001111111111 : node18153;
														assign node18153 = (inp[1]) ? node18155 : 16'b0000011111111111;
															assign node18155 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node18159 = (inp[12]) ? node18169 : node18160;
												assign node18160 = (inp[4]) ? node18166 : node18161;
													assign node18161 = (inp[9]) ? node18163 : 16'b0000111111111111;
														assign node18163 = (inp[1]) ? 16'b0000000111111111 : 16'b0000011111111111;
													assign node18166 = (inp[9]) ? 16'b0000011111111111 : 16'b0000001111111111;
												assign node18169 = (inp[3]) ? node18171 : 16'b0000001111111111;
													assign node18171 = (inp[1]) ? 16'b0000000011111111 : node18172;
														assign node18172 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node18176 = (inp[3]) ? node18200 : node18177;
											assign node18177 = (inp[9]) ? node18195 : node18178;
												assign node18178 = (inp[1]) ? node18188 : node18179;
													assign node18179 = (inp[12]) ? 16'b0000001111111111 : node18180;
														assign node18180 = (inp[4]) ? 16'b0000011111111111 : node18181;
															assign node18181 = (inp[2]) ? 16'b0000111111111111 : node18182;
																assign node18182 = (inp[10]) ? 16'b0000111111111111 : 16'b0001111111111111;
													assign node18188 = (inp[4]) ? node18192 : node18189;
														assign node18189 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node18192 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node18195 = (inp[12]) ? node18197 : 16'b0000001111111111;
													assign node18197 = (inp[10]) ? 16'b0000000011111111 : 16'b0000001111111111;
											assign node18200 = (inp[2]) ? node18212 : node18201;
												assign node18201 = (inp[10]) ? node18205 : node18202;
													assign node18202 = (inp[12]) ? 16'b0000011111111111 : 16'b0000001111111111;
													assign node18205 = (inp[9]) ? node18209 : node18206;
														assign node18206 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node18209 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node18212 = (inp[1]) ? node18214 : 16'b0000000111111111;
													assign node18214 = (inp[12]) ? 16'b0000000011111111 : node18215;
														assign node18215 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node18219 = (inp[10]) ? node18271 : node18220;
										assign node18220 = (inp[12]) ? node18246 : node18221;
											assign node18221 = (inp[11]) ? node18235 : node18222;
												assign node18222 = (inp[9]) ? node18230 : node18223;
													assign node18223 = (inp[3]) ? node18227 : node18224;
														assign node18224 = (inp[2]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node18227 = (inp[1]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node18230 = (inp[3]) ? node18232 : 16'b0000000111111111;
														assign node18232 = (inp[4]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node18235 = (inp[4]) ? node18241 : node18236;
													assign node18236 = (inp[2]) ? 16'b0000001111111111 : node18237;
														assign node18237 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node18241 = (inp[1]) ? 16'b0000000111111111 : node18242;
														assign node18242 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node18246 = (inp[9]) ? node18262 : node18247;
												assign node18247 = (inp[4]) ? node18255 : node18248;
													assign node18248 = (inp[3]) ? node18252 : node18249;
														assign node18249 = (inp[1]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node18252 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node18255 = (inp[3]) ? node18259 : node18256;
														assign node18256 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node18259 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node18262 = (inp[1]) ? node18266 : node18263;
													assign node18263 = (inp[3]) ? 16'b0000000111111111 : 16'b0000000011111111;
													assign node18266 = (inp[3]) ? node18268 : 16'b0000000011111111;
														assign node18268 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node18271 = (inp[2]) ? node18291 : node18272;
											assign node18272 = (inp[3]) ? node18284 : node18273;
												assign node18273 = (inp[9]) ? 16'b0000000111111111 : node18274;
													assign node18274 = (inp[12]) ? node18276 : 16'b0000111111111111;
														assign node18276 = (inp[1]) ? node18280 : node18277;
															assign node18277 = (inp[11]) ? 16'b0000001111111111 : 16'b0000011111111111;
															assign node18280 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node18284 = (inp[4]) ? node18286 : 16'b0000000111111111;
													assign node18286 = (inp[1]) ? node18288 : 16'b0000000111111111;
														assign node18288 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node18291 = (inp[3]) ? node18307 : node18292;
												assign node18292 = (inp[4]) ? node18300 : node18293;
													assign node18293 = (inp[1]) ? node18297 : node18294;
														assign node18294 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node18297 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node18300 = (inp[11]) ? 16'b0000000001111111 : node18301;
														assign node18301 = (inp[9]) ? 16'b0000000001111111 : node18302;
															assign node18302 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node18307 = (inp[9]) ? 16'b0000000001111111 : node18308;
													assign node18308 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000001111111;
								assign node18312 = (inp[12]) ? node18436 : node18313;
									assign node18313 = (inp[1]) ? node18385 : node18314;
										assign node18314 = (inp[2]) ? node18356 : node18315;
											assign node18315 = (inp[11]) ? node18339 : node18316;
												assign node18316 = (inp[9]) ? node18324 : node18317;
													assign node18317 = (inp[14]) ? node18319 : 16'b0000111111111111;
														assign node18319 = (inp[3]) ? node18321 : 16'b0000011111111111;
															assign node18321 = (inp[4]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node18324 = (inp[10]) ? node18330 : node18325;
														assign node18325 = (inp[4]) ? node18327 : 16'b0000011111111111;
															assign node18327 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node18330 = (inp[4]) ? node18336 : node18331;
															assign node18331 = (inp[3]) ? 16'b0000001111111111 : node18332;
																assign node18332 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
															assign node18336 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node18339 = (inp[4]) ? node18349 : node18340;
													assign node18340 = (inp[9]) ? node18344 : node18341;
														assign node18341 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node18344 = (inp[3]) ? node18346 : 16'b0000001111111111;
															assign node18346 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node18349 = (inp[9]) ? node18353 : node18350;
														assign node18350 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node18353 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node18356 = (inp[10]) ? node18374 : node18357;
												assign node18357 = (inp[11]) ? node18367 : node18358;
													assign node18358 = (inp[4]) ? node18360 : 16'b0000011111111111;
														assign node18360 = (inp[9]) ? 16'b0000000111111111 : node18361;
															assign node18361 = (inp[14]) ? node18363 : 16'b0000001111111111;
																assign node18363 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node18367 = (inp[14]) ? node18371 : node18368;
														assign node18368 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node18371 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node18374 = (inp[14]) ? 16'b0000000000111111 : node18375;
													assign node18375 = (inp[3]) ? 16'b0000000011111111 : node18376;
														assign node18376 = (inp[9]) ? node18378 : 16'b0000000111111111;
															assign node18378 = (inp[4]) ? node18380 : 16'b0000000111111111;
																assign node18380 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node18385 = (inp[3]) ? node18409 : node18386;
											assign node18386 = (inp[10]) ? node18394 : node18387;
												assign node18387 = (inp[14]) ? 16'b0000000111111111 : node18388;
													assign node18388 = (inp[9]) ? 16'b0000001111111111 : node18389;
														assign node18389 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node18394 = (inp[11]) ? node18404 : node18395;
													assign node18395 = (inp[9]) ? node18399 : node18396;
														assign node18396 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node18399 = (inp[2]) ? node18401 : 16'b0000000111111111;
															assign node18401 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node18404 = (inp[9]) ? 16'b0000000001111111 : node18405;
														assign node18405 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node18409 = (inp[10]) ? node18425 : node18410;
												assign node18410 = (inp[9]) ? node18414 : node18411;
													assign node18411 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node18414 = (inp[11]) ? node18420 : node18415;
														assign node18415 = (inp[14]) ? node18417 : 16'b0000000111111111;
															assign node18417 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node18420 = (inp[2]) ? node18422 : 16'b0000000011111111;
															assign node18422 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node18425 = (inp[4]) ? node18427 : 16'b0000000011111111;
													assign node18427 = (inp[9]) ? node18433 : node18428;
														assign node18428 = (inp[2]) ? 16'b0000000001111111 : node18429;
															assign node18429 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node18433 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000001111111;
									assign node18436 = (inp[10]) ? node18478 : node18437;
										assign node18437 = (inp[4]) ? node18459 : node18438;
											assign node18438 = (inp[11]) ? node18448 : node18439;
												assign node18439 = (inp[1]) ? 16'b0000000111111111 : node18440;
													assign node18440 = (inp[3]) ? 16'b0000001111111111 : node18441;
														assign node18441 = (inp[14]) ? node18443 : 16'b0000011111111111;
															assign node18443 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node18448 = (inp[2]) ? node18454 : node18449;
													assign node18449 = (inp[9]) ? 16'b0000000111111111 : node18450;
														assign node18450 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node18454 = (inp[14]) ? 16'b0000000001111111 : node18455;
														assign node18455 = (inp[1]) ? 16'b0000000111111111 : 16'b0000000011111111;
											assign node18459 = (inp[1]) ? node18471 : node18460;
												assign node18460 = (inp[14]) ? node18466 : node18461;
													assign node18461 = (inp[2]) ? 16'b0000000011111111 : node18462;
														assign node18462 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node18466 = (inp[9]) ? node18468 : 16'b0000000011111111;
														assign node18468 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node18471 = (inp[9]) ? 16'b0000000001111111 : node18472;
													assign node18472 = (inp[11]) ? 16'b0000000001111111 : node18473;
														assign node18473 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node18478 = (inp[9]) ? node18504 : node18479;
											assign node18479 = (inp[4]) ? node18489 : node18480;
												assign node18480 = (inp[1]) ? node18482 : 16'b0000000111111111;
													assign node18482 = (inp[2]) ? node18486 : node18483;
														assign node18483 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node18486 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node18489 = (inp[1]) ? node18497 : node18490;
													assign node18490 = (inp[14]) ? 16'b0000000001111111 : node18491;
														assign node18491 = (inp[2]) ? 16'b0000000011111111 : node18492;
															assign node18492 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node18497 = (inp[11]) ? 16'b0000000000111111 : node18498;
														assign node18498 = (inp[14]) ? 16'b0000000001111111 : node18499;
															assign node18499 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node18504 = (inp[14]) ? node18514 : node18505;
												assign node18505 = (inp[4]) ? 16'b0000000001111111 : node18506;
													assign node18506 = (inp[3]) ? 16'b0000000001111111 : node18507;
														assign node18507 = (inp[11]) ? node18509 : 16'b0000000011111111;
															assign node18509 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node18514 = (inp[3]) ? node18518 : node18515;
													assign node18515 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node18518 = (inp[11]) ? node18524 : node18519;
														assign node18519 = (inp[2]) ? node18521 : 16'b0000000000111111;
															assign node18521 = (inp[4]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node18524 = (inp[4]) ? 16'b0000000000001111 : 16'b0000000000011111;
							assign node18527 = (inp[11]) ? node18691 : node18528;
								assign node18528 = (inp[1]) ? node18596 : node18529;
									assign node18529 = (inp[4]) ? node18569 : node18530;
										assign node18530 = (inp[12]) ? node18548 : node18531;
											assign node18531 = (inp[6]) ? node18533 : 16'b0000001111111111;
												assign node18533 = (inp[14]) ? node18537 : node18534;
													assign node18534 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node18537 = (inp[9]) ? node18545 : node18538;
														assign node18538 = (inp[10]) ? 16'b0000000111111111 : node18539;
															assign node18539 = (inp[2]) ? 16'b0000001111111111 : node18540;
																assign node18540 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node18545 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node18548 = (inp[6]) ? node18562 : node18549;
												assign node18549 = (inp[2]) ? node18551 : 16'b0000001111111111;
													assign node18551 = (inp[14]) ? node18557 : node18552;
														assign node18552 = (inp[10]) ? node18554 : 16'b0000001111111111;
															assign node18554 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node18557 = (inp[10]) ? node18559 : 16'b0000000011111111;
															assign node18559 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node18562 = (inp[3]) ? 16'b0000000011111111 : node18563;
													assign node18563 = (inp[9]) ? node18565 : 16'b0000000111111111;
														assign node18565 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node18569 = (inp[10]) ? node18583 : node18570;
											assign node18570 = (inp[3]) ? node18576 : node18571;
												assign node18571 = (inp[2]) ? node18573 : 16'b0000011111111111;
													assign node18573 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node18576 = (inp[9]) ? node18578 : 16'b0000000111111111;
													assign node18578 = (inp[2]) ? 16'b0000000000111111 : node18579;
														assign node18579 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node18583 = (inp[6]) ? node18591 : node18584;
												assign node18584 = (inp[3]) ? 16'b0000000011111111 : node18585;
													assign node18585 = (inp[9]) ? node18587 : 16'b0000001111111111;
														assign node18587 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node18591 = (inp[2]) ? node18593 : 16'b0000000011111111;
													assign node18593 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node18596 = (inp[14]) ? node18646 : node18597;
										assign node18597 = (inp[2]) ? node18619 : node18598;
											assign node18598 = (inp[9]) ? node18608 : node18599;
												assign node18599 = (inp[12]) ? node18603 : node18600;
													assign node18600 = (inp[10]) ? 16'b0000001111111111 : 16'b0000111111111111;
													assign node18603 = (inp[4]) ? node18605 : 16'b0000001111111111;
														assign node18605 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node18608 = (inp[12]) ? node18614 : node18609;
													assign node18609 = (inp[4]) ? 16'b0000000111111111 : node18610;
														assign node18610 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node18614 = (inp[3]) ? 16'b0000000011111111 : node18615;
														assign node18615 = (inp[10]) ? 16'b0000000011111111 : 16'b0000001111111111;
											assign node18619 = (inp[12]) ? node18635 : node18620;
												assign node18620 = (inp[3]) ? node18626 : node18621;
													assign node18621 = (inp[6]) ? 16'b0000000011111111 : node18622;
														assign node18622 = (inp[10]) ? 16'b0000000111111111 : 16'b0000011111111111;
													assign node18626 = (inp[10]) ? node18628 : 16'b0000000111111111;
														assign node18628 = (inp[9]) ? node18630 : 16'b0000000011111111;
															assign node18630 = (inp[4]) ? node18632 : 16'b0000000001111111;
																assign node18632 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node18635 = (inp[6]) ? node18641 : node18636;
													assign node18636 = (inp[10]) ? node18638 : 16'b0000000011111111;
														assign node18638 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node18641 = (inp[3]) ? 16'b0000000001111111 : node18642;
														assign node18642 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node18646 = (inp[2]) ? node18668 : node18647;
											assign node18647 = (inp[6]) ? node18655 : node18648;
												assign node18648 = (inp[3]) ? 16'b0000000011111111 : node18649;
													assign node18649 = (inp[12]) ? node18651 : 16'b0000000111111111;
														assign node18651 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node18655 = (inp[9]) ? node18663 : node18656;
													assign node18656 = (inp[10]) ? node18660 : node18657;
														assign node18657 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node18660 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node18663 = (inp[10]) ? node18665 : 16'b0000000001111111;
														assign node18665 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node18668 = (inp[9]) ? node18682 : node18669;
												assign node18669 = (inp[3]) ? node18673 : node18670;
													assign node18670 = (inp[6]) ? 16'b0000000111111111 : 16'b0000000011111111;
													assign node18673 = (inp[12]) ? node18677 : node18674;
														assign node18674 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node18677 = (inp[6]) ? node18679 : 16'b0000000001111111;
															assign node18679 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node18682 = (inp[4]) ? node18688 : node18683;
													assign node18683 = (inp[12]) ? node18685 : 16'b0000000001111111;
														assign node18685 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node18688 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
								assign node18691 = (inp[6]) ? node18779 : node18692;
									assign node18692 = (inp[4]) ? node18748 : node18693;
										assign node18693 = (inp[14]) ? node18725 : node18694;
											assign node18694 = (inp[10]) ? node18710 : node18695;
												assign node18695 = (inp[12]) ? node18701 : node18696;
													assign node18696 = (inp[9]) ? 16'b0000001111111111 : node18697;
														assign node18697 = (inp[2]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node18701 = (inp[3]) ? node18705 : node18702;
														assign node18702 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node18705 = (inp[2]) ? node18707 : 16'b0000000111111111;
															assign node18707 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node18710 = (inp[9]) ? node18718 : node18711;
													assign node18711 = (inp[12]) ? 16'b0000000011111111 : node18712;
														assign node18712 = (inp[2]) ? node18714 : 16'b0000001111111111;
															assign node18714 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node18718 = (inp[3]) ? node18720 : 16'b0000000011111111;
														assign node18720 = (inp[12]) ? 16'b0000000001111111 : node18721;
															assign node18721 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node18725 = (inp[12]) ? node18733 : node18726;
												assign node18726 = (inp[9]) ? 16'b0000000011111111 : node18727;
													assign node18727 = (inp[2]) ? node18729 : 16'b0000000111111111;
														assign node18729 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node18733 = (inp[3]) ? node18739 : node18734;
													assign node18734 = (inp[2]) ? 16'b0000000011111111 : node18735;
														assign node18735 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node18739 = (inp[10]) ? node18745 : node18740;
														assign node18740 = (inp[2]) ? node18742 : 16'b0000000011111111;
															assign node18742 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node18745 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node18748 = (inp[14]) ? node18770 : node18749;
											assign node18749 = (inp[12]) ? node18757 : node18750;
												assign node18750 = (inp[9]) ? node18752 : 16'b0000000111111111;
													assign node18752 = (inp[10]) ? node18754 : 16'b0000000111111111;
														assign node18754 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node18757 = (inp[1]) ? node18765 : node18758;
													assign node18758 = (inp[3]) ? node18760 : 16'b0000000111111111;
														assign node18760 = (inp[9]) ? 16'b0000000001111111 : node18761;
															assign node18761 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node18765 = (inp[9]) ? node18767 : 16'b0000000001111111;
														assign node18767 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000001111111;
											assign node18770 = (inp[1]) ? 16'b0000000000111111 : node18771;
												assign node18771 = (inp[3]) ? 16'b0000000001111111 : node18772;
													assign node18772 = (inp[12]) ? node18774 : 16'b0000000011111111;
														assign node18774 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node18779 = (inp[14]) ? node18825 : node18780;
										assign node18780 = (inp[3]) ? node18802 : node18781;
											assign node18781 = (inp[9]) ? node18787 : node18782;
												assign node18782 = (inp[12]) ? node18784 : 16'b0000000111111111;
													assign node18784 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node18787 = (inp[1]) ? node18797 : node18788;
													assign node18788 = (inp[10]) ? node18794 : node18789;
														assign node18789 = (inp[4]) ? node18791 : 16'b0000000111111111;
															assign node18791 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node18794 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node18797 = (inp[4]) ? 16'b0000000000111111 : node18798;
														assign node18798 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node18802 = (inp[1]) ? node18816 : node18803;
												assign node18803 = (inp[9]) ? node18809 : node18804;
													assign node18804 = (inp[4]) ? node18806 : 16'b0000000011111111;
														assign node18806 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node18809 = (inp[10]) ? node18813 : node18810;
														assign node18810 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node18813 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000001111111;
												assign node18816 = (inp[9]) ? 16'b0000000000111111 : node18817;
													assign node18817 = (inp[4]) ? node18819 : 16'b0000000001111111;
														assign node18819 = (inp[2]) ? 16'b0000000000111111 : node18820;
															assign node18820 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node18825 = (inp[1]) ? node18849 : node18826;
											assign node18826 = (inp[2]) ? node18836 : node18827;
												assign node18827 = (inp[10]) ? node18831 : node18828;
													assign node18828 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node18831 = (inp[4]) ? 16'b0000000001111111 : node18832;
														assign node18832 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node18836 = (inp[3]) ? node18842 : node18837;
													assign node18837 = (inp[10]) ? node18839 : 16'b0000000001111111;
														assign node18839 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000001111111;
													assign node18842 = (inp[12]) ? node18844 : 16'b0000000000111111;
														assign node18844 = (inp[4]) ? node18846 : 16'b0000000000111111;
															assign node18846 = (inp[9]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node18849 = (inp[10]) ? node18859 : node18850;
												assign node18850 = (inp[3]) ? node18852 : 16'b0000000001111111;
													assign node18852 = (inp[12]) ? node18856 : node18853;
														assign node18853 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node18856 = (inp[4]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node18859 = (inp[4]) ? 16'b0000000000011111 : node18860;
													assign node18860 = (inp[3]) ? node18862 : 16'b0000000000111111;
														assign node18862 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
						assign node18866 = (inp[4]) ? node19248 : node18867;
							assign node18867 = (inp[3]) ? node19057 : node18868;
								assign node18868 = (inp[9]) ? node18970 : node18869;
									assign node18869 = (inp[14]) ? node18931 : node18870;
										assign node18870 = (inp[15]) ? node18902 : node18871;
											assign node18871 = (inp[11]) ? node18889 : node18872;
												assign node18872 = (inp[1]) ? node18884 : node18873;
													assign node18873 = (inp[12]) ? node18881 : node18874;
														assign node18874 = (inp[10]) ? 16'b0000011111111111 : node18875;
															assign node18875 = (inp[2]) ? node18877 : 16'b0000111111111111;
																assign node18877 = (inp[6]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node18881 = (inp[6]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node18884 = (inp[6]) ? node18886 : 16'b0000001111111111;
														assign node18886 = (inp[2]) ? 16'b0000000111111111 : 16'b0000011111111111;
												assign node18889 = (inp[10]) ? node18893 : node18890;
													assign node18890 = (inp[1]) ? 16'b0000011111111111 : 16'b0000001111111111;
													assign node18893 = (inp[1]) ? node18899 : node18894;
														assign node18894 = (inp[2]) ? 16'b0000000111111111 : node18895;
															assign node18895 = (inp[6]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node18899 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node18902 = (inp[6]) ? node18918 : node18903;
												assign node18903 = (inp[2]) ? node18913 : node18904;
													assign node18904 = (inp[1]) ? node18908 : node18905;
														assign node18905 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node18908 = (inp[12]) ? 16'b0000000111111111 : node18909;
															assign node18909 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node18913 = (inp[1]) ? node18915 : 16'b0000000111111111;
														assign node18915 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node18918 = (inp[11]) ? 16'b0000000011111111 : node18919;
													assign node18919 = (inp[1]) ? node18923 : node18920;
														assign node18920 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node18923 = (inp[12]) ? node18925 : 16'b0000000111111111;
															assign node18925 = (inp[2]) ? 16'b0000000011111111 : node18926;
																assign node18926 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node18931 = (inp[2]) ? node18947 : node18932;
											assign node18932 = (inp[6]) ? node18940 : node18933;
												assign node18933 = (inp[1]) ? node18935 : 16'b0000001111111111;
													assign node18935 = (inp[12]) ? 16'b0000000011111111 : node18936;
														assign node18936 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node18940 = (inp[15]) ? node18942 : 16'b0000000111111111;
													assign node18942 = (inp[11]) ? 16'b0000000011111111 : node18943;
														assign node18943 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node18947 = (inp[11]) ? node18961 : node18948;
												assign node18948 = (inp[6]) ? node18954 : node18949;
													assign node18949 = (inp[12]) ? 16'b0000000111111111 : node18950;
														assign node18950 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node18954 = (inp[10]) ? 16'b0000000001111111 : node18955;
														assign node18955 = (inp[12]) ? 16'b0000000011111111 : node18956;
															assign node18956 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node18961 = (inp[1]) ? node18967 : node18962;
													assign node18962 = (inp[6]) ? node18964 : 16'b0000000011111111;
														assign node18964 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node18967 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node18970 = (inp[2]) ? node19016 : node18971;
										assign node18971 = (inp[1]) ? node18993 : node18972;
											assign node18972 = (inp[10]) ? node18982 : node18973;
												assign node18973 = (inp[14]) ? node18975 : 16'b0000001111111111;
													assign node18975 = (inp[12]) ? node18979 : node18976;
														assign node18976 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node18979 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node18982 = (inp[15]) ? node18988 : node18983;
													assign node18983 = (inp[11]) ? 16'b0000000111111111 : node18984;
														assign node18984 = (inp[12]) ? 16'b0000001111111111 : 16'b0000000111111111;
													assign node18988 = (inp[11]) ? node18990 : 16'b0000000111111111;
														assign node18990 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node18993 = (inp[12]) ? node19001 : node18994;
												assign node18994 = (inp[6]) ? node18996 : 16'b0000001111111111;
													assign node18996 = (inp[15]) ? 16'b0000000011111111 : node18997;
														assign node18997 = (inp[14]) ? 16'b0000000111111111 : 16'b0000000011111111;
												assign node19001 = (inp[10]) ? node19011 : node19002;
													assign node19002 = (inp[6]) ? 16'b0000000011111111 : node19003;
														assign node19003 = (inp[11]) ? 16'b0000000011111111 : node19004;
															assign node19004 = (inp[14]) ? node19006 : 16'b0000000111111111;
																assign node19006 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node19011 = (inp[14]) ? node19013 : 16'b0000000011111111;
														assign node19013 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node19016 = (inp[6]) ? node19028 : node19017;
											assign node19017 = (inp[15]) ? node19021 : node19018;
												assign node19018 = (inp[10]) ? 16'b0000000011111111 : 16'b0000001111111111;
												assign node19021 = (inp[14]) ? 16'b0000000001111111 : node19022;
													assign node19022 = (inp[1]) ? 16'b0000000001111111 : node19023;
														assign node19023 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node19028 = (inp[11]) ? node19044 : node19029;
												assign node19029 = (inp[15]) ? node19035 : node19030;
													assign node19030 = (inp[12]) ? 16'b0000000011111111 : node19031;
														assign node19031 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node19035 = (inp[14]) ? node19039 : node19036;
														assign node19036 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node19039 = (inp[10]) ? 16'b0000000000111111 : node19040;
															assign node19040 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node19044 = (inp[15]) ? node19050 : node19045;
													assign node19045 = (inp[14]) ? node19047 : 16'b0000000001111111;
														assign node19047 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node19050 = (inp[14]) ? 16'b0000000000001111 : node19051;
														assign node19051 = (inp[1]) ? node19053 : 16'b0000000000111111;
															assign node19053 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000111111;
								assign node19057 = (inp[1]) ? node19163 : node19058;
									assign node19058 = (inp[11]) ? node19110 : node19059;
										assign node19059 = (inp[12]) ? node19079 : node19060;
											assign node19060 = (inp[14]) ? node19070 : node19061;
												assign node19061 = (inp[9]) ? 16'b0000000111111111 : node19062;
													assign node19062 = (inp[6]) ? node19066 : node19063;
														assign node19063 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node19066 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node19070 = (inp[2]) ? 16'b0000000011111111 : node19071;
													assign node19071 = (inp[10]) ? node19075 : node19072;
														assign node19072 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node19075 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node19079 = (inp[10]) ? node19099 : node19080;
												assign node19080 = (inp[14]) ? node19096 : node19081;
													assign node19081 = (inp[9]) ? node19087 : node19082;
														assign node19082 = (inp[2]) ? node19084 : 16'b0000001111111111;
															assign node19084 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node19087 = (inp[2]) ? node19091 : node19088;
															assign node19088 = (inp[6]) ? 16'b0000000111111111 : 16'b0000001111111111;
															assign node19091 = (inp[6]) ? 16'b0000000011111111 : node19092;
																assign node19092 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node19096 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node19099 = (inp[2]) ? node19101 : 16'b0000000011111111;
													assign node19101 = (inp[6]) ? node19105 : node19102;
														assign node19102 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node19105 = (inp[14]) ? node19107 : 16'b0000000001111111;
															assign node19107 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node19110 = (inp[15]) ? node19140 : node19111;
											assign node19111 = (inp[9]) ? node19121 : node19112;
												assign node19112 = (inp[10]) ? 16'b0000000011111111 : node19113;
													assign node19113 = (inp[2]) ? node19115 : 16'b0000001111111111;
														assign node19115 = (inp[12]) ? 16'b0000000011111111 : node19116;
															assign node19116 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node19121 = (inp[10]) ? node19135 : node19122;
													assign node19122 = (inp[14]) ? node19130 : node19123;
														assign node19123 = (inp[12]) ? 16'b0000000011111111 : node19124;
															assign node19124 = (inp[2]) ? node19126 : 16'b0000000111111111;
																assign node19126 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node19130 = (inp[2]) ? 16'b0000000001111111 : node19131;
															assign node19131 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node19135 = (inp[2]) ? 16'b0000000001111111 : node19136;
														assign node19136 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node19140 = (inp[6]) ? node19148 : node19141;
												assign node19141 = (inp[9]) ? node19145 : node19142;
													assign node19142 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node19145 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000001111111;
												assign node19148 = (inp[10]) ? node19156 : node19149;
													assign node19149 = (inp[14]) ? node19153 : node19150;
														assign node19150 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node19153 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node19156 = (inp[9]) ? node19160 : node19157;
														assign node19157 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node19160 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node19163 = (inp[6]) ? node19203 : node19164;
										assign node19164 = (inp[15]) ? node19188 : node19165;
											assign node19165 = (inp[2]) ? node19175 : node19166;
												assign node19166 = (inp[9]) ? node19168 : 16'b0000000111111111;
													assign node19168 = (inp[11]) ? node19172 : node19169;
														assign node19169 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node19172 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node19175 = (inp[12]) ? node19183 : node19176;
													assign node19176 = (inp[9]) ? node19178 : 16'b0000000011111111;
														assign node19178 = (inp[14]) ? 16'b0000000001111111 : node19179;
															assign node19179 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node19183 = (inp[9]) ? 16'b0000000001111111 : node19184;
														assign node19184 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node19188 = (inp[14]) ? node19194 : node19189;
												assign node19189 = (inp[10]) ? 16'b0000000001111111 : node19190;
													assign node19190 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node19194 = (inp[11]) ? node19200 : node19195;
													assign node19195 = (inp[2]) ? node19197 : 16'b0000000001111111;
														assign node19197 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node19200 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node19203 = (inp[2]) ? node19233 : node19204;
											assign node19204 = (inp[14]) ? node19220 : node19205;
												assign node19205 = (inp[9]) ? node19217 : node19206;
													assign node19206 = (inp[10]) ? node19212 : node19207;
														assign node19207 = (inp[12]) ? node19209 : 16'b0000000011111111;
															assign node19209 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node19212 = (inp[15]) ? 16'b0000000001111111 : node19213;
															assign node19213 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node19217 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node19220 = (inp[11]) ? node19228 : node19221;
													assign node19221 = (inp[12]) ? node19225 : node19222;
														assign node19222 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node19225 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node19228 = (inp[10]) ? node19230 : 16'b0000000000111111;
														assign node19230 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node19233 = (inp[11]) ? node19243 : node19234;
												assign node19234 = (inp[15]) ? 16'b0000000000111111 : node19235;
													assign node19235 = (inp[10]) ? node19237 : 16'b0000000000111111;
														assign node19237 = (inp[14]) ? node19239 : 16'b0000000000111111;
															assign node19239 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node19243 = (inp[12]) ? 16'b0000000000011111 : node19244;
													assign node19244 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
							assign node19248 = (inp[2]) ? node19454 : node19249;
								assign node19249 = (inp[9]) ? node19341 : node19250;
									assign node19250 = (inp[14]) ? node19280 : node19251;
										assign node19251 = (inp[3]) ? node19267 : node19252;
											assign node19252 = (inp[10]) ? node19260 : node19253;
												assign node19253 = (inp[1]) ? 16'b0000000111111111 : node19254;
													assign node19254 = (inp[11]) ? 16'b0000001111111111 : node19255;
														assign node19255 = (inp[6]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node19260 = (inp[15]) ? 16'b0000000011111111 : node19261;
													assign node19261 = (inp[1]) ? node19263 : 16'b0000000111111111;
														assign node19263 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node19267 = (inp[15]) ? node19273 : node19268;
												assign node19268 = (inp[6]) ? node19270 : 16'b0000000111111111;
													assign node19270 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node19273 = (inp[12]) ? node19275 : 16'b0000000011111111;
													assign node19275 = (inp[11]) ? 16'b0000000001111111 : node19276;
														assign node19276 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node19280 = (inp[6]) ? node19312 : node19281;
											assign node19281 = (inp[1]) ? node19299 : node19282;
												assign node19282 = (inp[12]) ? node19292 : node19283;
													assign node19283 = (inp[15]) ? node19289 : node19284;
														assign node19284 = (inp[11]) ? 16'b0000000111111111 : node19285;
															assign node19285 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node19289 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node19292 = (inp[15]) ? node19296 : node19293;
														assign node19293 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node19296 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node19299 = (inp[3]) ? node19307 : node19300;
													assign node19300 = (inp[12]) ? node19304 : node19301;
														assign node19301 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node19304 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node19307 = (inp[15]) ? node19309 : 16'b0000000001111111;
														assign node19309 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node19312 = (inp[11]) ? node19324 : node19313;
												assign node19313 = (inp[10]) ? node19319 : node19314;
													assign node19314 = (inp[3]) ? 16'b0000000001111111 : node19315;
														assign node19315 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node19319 = (inp[1]) ? 16'b0000000001111111 : node19320;
														assign node19320 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node19324 = (inp[12]) ? node19334 : node19325;
													assign node19325 = (inp[3]) ? node19331 : node19326;
														assign node19326 = (inp[15]) ? node19328 : 16'b0000000011111111;
															assign node19328 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node19331 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node19334 = (inp[10]) ? node19336 : 16'b0000000001111111;
														assign node19336 = (inp[3]) ? 16'b0000000000011111 : node19337;
															assign node19337 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node19341 = (inp[15]) ? node19395 : node19342;
										assign node19342 = (inp[3]) ? node19370 : node19343;
											assign node19343 = (inp[12]) ? node19359 : node19344;
												assign node19344 = (inp[10]) ? node19354 : node19345;
													assign node19345 = (inp[1]) ? node19349 : node19346;
														assign node19346 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node19349 = (inp[14]) ? node19351 : 16'b0000000111111111;
															assign node19351 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node19354 = (inp[11]) ? 16'b0000000011111111 : node19355;
														assign node19355 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node19359 = (inp[10]) ? node19365 : node19360;
													assign node19360 = (inp[14]) ? 16'b0000000011111111 : node19361;
														assign node19361 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node19365 = (inp[1]) ? node19367 : 16'b0000000011111111;
														assign node19367 = (inp[6]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node19370 = (inp[11]) ? node19386 : node19371;
												assign node19371 = (inp[1]) ? node19377 : node19372;
													assign node19372 = (inp[14]) ? 16'b0000000011111111 : node19373;
														assign node19373 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node19377 = (inp[12]) ? node19383 : node19378;
														assign node19378 = (inp[14]) ? 16'b0000000001111111 : node19379;
															assign node19379 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node19383 = (inp[6]) ? 16'b0000000000011111 : 16'b0000000001111111;
												assign node19386 = (inp[6]) ? node19392 : node19387;
													assign node19387 = (inp[10]) ? node19389 : 16'b0000000001111111;
														assign node19389 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node19392 = (inp[14]) ? 16'b0000000000001111 : 16'b0000000000111111;
										assign node19395 = (inp[14]) ? node19427 : node19396;
											assign node19396 = (inp[11]) ? node19408 : node19397;
												assign node19397 = (inp[10]) ? node19401 : node19398;
													assign node19398 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node19401 = (inp[1]) ? node19403 : 16'b0000000001111111;
														assign node19403 = (inp[6]) ? 16'b0000000000111111 : node19404;
															assign node19404 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node19408 = (inp[3]) ? node19412 : node19409;
													assign node19409 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000001111111;
													assign node19412 = (inp[1]) ? node19420 : node19413;
														assign node19413 = (inp[12]) ? node19415 : 16'b0000000001111111;
															assign node19415 = (inp[6]) ? 16'b0000000000111111 : node19416;
																assign node19416 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node19420 = (inp[10]) ? 16'b0000000000011111 : node19421;
															assign node19421 = (inp[6]) ? 16'b0000000000111111 : node19422;
																assign node19422 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node19427 = (inp[6]) ? node19435 : node19428;
												assign node19428 = (inp[11]) ? 16'b0000000000111111 : node19429;
													assign node19429 = (inp[1]) ? node19431 : 16'b0000000000111111;
														assign node19431 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node19435 = (inp[11]) ? node19443 : node19436;
													assign node19436 = (inp[1]) ? node19438 : 16'b0000000001111111;
														assign node19438 = (inp[12]) ? node19440 : 16'b0000000000111111;
															assign node19440 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node19443 = (inp[1]) ? node19447 : node19444;
														assign node19444 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000001111111;
														assign node19447 = (inp[3]) ? 16'b0000000000001111 : node19448;
															assign node19448 = (inp[10]) ? node19450 : 16'b0000000000011111;
																assign node19450 = (inp[12]) ? 16'b0000000000001111 : 16'b0000000000011111;
								assign node19454 = (inp[10]) ? node19546 : node19455;
									assign node19455 = (inp[14]) ? node19505 : node19456;
										assign node19456 = (inp[11]) ? node19486 : node19457;
											assign node19457 = (inp[6]) ? node19473 : node19458;
												assign node19458 = (inp[15]) ? node19468 : node19459;
													assign node19459 = (inp[3]) ? 16'b0000000011111111 : node19460;
														assign node19460 = (inp[9]) ? node19462 : 16'b0000001111111111;
															assign node19462 = (inp[1]) ? 16'b0000000111111111 : node19463;
																assign node19463 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node19468 = (inp[12]) ? 16'b0000000001111111 : node19469;
														assign node19469 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node19473 = (inp[9]) ? node19479 : node19474;
													assign node19474 = (inp[1]) ? 16'b0000000011111111 : node19475;
														assign node19475 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node19479 = (inp[12]) ? node19483 : node19480;
														assign node19480 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node19483 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node19486 = (inp[9]) ? node19490 : node19487;
												assign node19487 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node19490 = (inp[12]) ? 16'b0000000000111111 : node19491;
													assign node19491 = (inp[6]) ? node19499 : node19492;
														assign node19492 = (inp[1]) ? node19494 : 16'b0000000011111111;
															assign node19494 = (inp[3]) ? 16'b0000000001111111 : node19495;
																assign node19495 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node19499 = (inp[1]) ? node19501 : 16'b0000000001111111;
															assign node19501 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node19505 = (inp[6]) ? node19523 : node19506;
											assign node19506 = (inp[9]) ? node19514 : node19507;
												assign node19507 = (inp[11]) ? node19509 : 16'b0000000011111111;
													assign node19509 = (inp[15]) ? 16'b0000000001111111 : node19510;
														assign node19510 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node19514 = (inp[1]) ? node19520 : node19515;
													assign node19515 = (inp[11]) ? node19517 : 16'b0000000001111111;
														assign node19517 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node19520 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000001111111;
											assign node19523 = (inp[9]) ? node19529 : node19524;
												assign node19524 = (inp[3]) ? 16'b0000000000111111 : node19525;
													assign node19525 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node19529 = (inp[12]) ? node19539 : node19530;
													assign node19530 = (inp[3]) ? node19536 : node19531;
														assign node19531 = (inp[11]) ? 16'b0000000000111111 : node19532;
															assign node19532 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node19536 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node19539 = (inp[1]) ? node19541 : 16'b0000000000111111;
														assign node19541 = (inp[3]) ? node19543 : 16'b0000000000011111;
															assign node19543 = (inp[11]) ? 16'b0000000000000111 : 16'b0000000000001111;
									assign node19546 = (inp[6]) ? node19596 : node19547;
										assign node19547 = (inp[11]) ? node19569 : node19548;
											assign node19548 = (inp[3]) ? node19562 : node19549;
												assign node19549 = (inp[14]) ? node19555 : node19550;
													assign node19550 = (inp[15]) ? node19552 : 16'b0000000011111111;
														assign node19552 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node19555 = (inp[9]) ? node19559 : node19556;
														assign node19556 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node19559 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node19562 = (inp[15]) ? node19564 : 16'b0000000001111111;
													assign node19564 = (inp[14]) ? 16'b0000000000011111 : node19565;
														assign node19565 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000000111111;
											assign node19569 = (inp[12]) ? node19581 : node19570;
												assign node19570 = (inp[15]) ? node19576 : node19571;
													assign node19571 = (inp[14]) ? 16'b0000000001111111 : node19572;
														assign node19572 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node19576 = (inp[14]) ? 16'b0000000000111111 : node19577;
														assign node19577 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node19581 = (inp[15]) ? node19593 : node19582;
													assign node19582 = (inp[1]) ? node19590 : node19583;
														assign node19583 = (inp[9]) ? node19585 : 16'b0000000001111111;
															assign node19585 = (inp[3]) ? 16'b0000000000111111 : node19586;
																assign node19586 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node19590 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node19593 = (inp[3]) ? 16'b0000000000001111 : 16'b0000000000011111;
										assign node19596 = (inp[11]) ? node19612 : node19597;
											assign node19597 = (inp[12]) ? node19605 : node19598;
												assign node19598 = (inp[9]) ? 16'b0000000000111111 : node19599;
													assign node19599 = (inp[15]) ? 16'b0000000001111111 : node19600;
														assign node19600 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node19605 = (inp[14]) ? 16'b0000000000011111 : node19606;
													assign node19606 = (inp[9]) ? 16'b0000000000111111 : node19607;
														assign node19607 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node19612 = (inp[9]) ? node19626 : node19613;
												assign node19613 = (inp[14]) ? node19619 : node19614;
													assign node19614 = (inp[15]) ? 16'b0000000000011111 : node19615;
														assign node19615 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000001111111;
													assign node19619 = (inp[12]) ? node19621 : 16'b0000000000011111;
														assign node19621 = (inp[1]) ? node19623 : 16'b0000000000011111;
															assign node19623 = (inp[15]) ? 16'b0000000000000111 : 16'b0000000000001111;
												assign node19626 = (inp[3]) ? node19628 : 16'b0000000000111111;
													assign node19628 = (inp[1]) ? node19636 : node19629;
														assign node19629 = (inp[15]) ? 16'b0000000000001111 : node19630;
															assign node19630 = (inp[12]) ? node19632 : 16'b0000000000011111;
																assign node19632 = (inp[14]) ? 16'b0000000000001111 : 16'b0000000000011111;
														assign node19636 = (inp[12]) ? node19638 : 16'b0000000000001111;
															assign node19638 = (inp[15]) ? 16'b0000000000000011 : node19639;
																assign node19639 = (inp[14]) ? 16'b0000000000000111 : 16'b0000000000001111;
					assign node19643 = (inp[1]) ? node20373 : node19644;
						assign node19644 = (inp[3]) ? node20016 : node19645;
							assign node19645 = (inp[10]) ? node19831 : node19646;
								assign node19646 = (inp[12]) ? node19738 : node19647;
									assign node19647 = (inp[15]) ? node19703 : node19648;
										assign node19648 = (inp[4]) ? node19678 : node19649;
											assign node19649 = (inp[11]) ? node19667 : node19650;
												assign node19650 = (inp[9]) ? node19658 : node19651;
													assign node19651 = (inp[6]) ? node19655 : node19652;
														assign node19652 = (inp[13]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node19655 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node19658 = (inp[2]) ? 16'b0000001111111111 : node19659;
														assign node19659 = (inp[6]) ? 16'b0000001111111111 : node19660;
															assign node19660 = (inp[13]) ? node19662 : 16'b0000011111111111;
																assign node19662 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node19667 = (inp[9]) ? node19675 : node19668;
													assign node19668 = (inp[14]) ? node19670 : 16'b0000001111111111;
														assign node19670 = (inp[6]) ? node19672 : 16'b0000001111111111;
															assign node19672 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node19675 = (inp[6]) ? 16'b0000000011111111 : 16'b0000001111111111;
											assign node19678 = (inp[14]) ? node19694 : node19679;
												assign node19679 = (inp[9]) ? node19685 : node19680;
													assign node19680 = (inp[13]) ? 16'b0000001111111111 : node19681;
														assign node19681 = (inp[6]) ? 16'b0000001111111111 : 16'b0000111111111111;
													assign node19685 = (inp[6]) ? 16'b0000000011111111 : node19686;
														assign node19686 = (inp[11]) ? node19688 : 16'b0000001111111111;
															assign node19688 = (inp[13]) ? 16'b0000000111111111 : node19689;
																assign node19689 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node19694 = (inp[2]) ? 16'b0000000011111111 : node19695;
													assign node19695 = (inp[9]) ? node19699 : node19696;
														assign node19696 = (inp[6]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node19699 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node19703 = (inp[9]) ? node19719 : node19704;
											assign node19704 = (inp[2]) ? node19714 : node19705;
												assign node19705 = (inp[6]) ? node19711 : node19706;
													assign node19706 = (inp[4]) ? 16'b0000001111111111 : node19707;
														assign node19707 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node19711 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node19714 = (inp[13]) ? node19716 : 16'b0000000111111111;
													assign node19716 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node19719 = (inp[4]) ? node19731 : node19720;
												assign node19720 = (inp[13]) ? node19728 : node19721;
													assign node19721 = (inp[6]) ? node19723 : 16'b0000001111111111;
														assign node19723 = (inp[2]) ? node19725 : 16'b0000000111111111;
															assign node19725 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000111111111;
													assign node19728 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node19731 = (inp[6]) ? node19733 : 16'b0000000011111111;
													assign node19733 = (inp[2]) ? 16'b0000000001111111 : node19734;
														assign node19734 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node19738 = (inp[4]) ? node19790 : node19739;
										assign node19739 = (inp[14]) ? node19771 : node19740;
											assign node19740 = (inp[9]) ? node19754 : node19741;
												assign node19741 = (inp[2]) ? node19749 : node19742;
													assign node19742 = (inp[13]) ? 16'b0000000111111111 : node19743;
														assign node19743 = (inp[15]) ? 16'b0000001111111111 : node19744;
															assign node19744 = (inp[6]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node19749 = (inp[15]) ? 16'b0000000111111111 : node19750;
														assign node19750 = (inp[6]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node19754 = (inp[13]) ? node19762 : node19755;
													assign node19755 = (inp[15]) ? node19759 : node19756;
														assign node19756 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node19759 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node19762 = (inp[6]) ? node19764 : 16'b0000000111111111;
														assign node19764 = (inp[11]) ? 16'b0000000001111111 : node19765;
															assign node19765 = (inp[2]) ? node19767 : 16'b0000000011111111;
																assign node19767 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node19771 = (inp[9]) ? node19775 : node19772;
												assign node19772 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node19775 = (inp[13]) ? node19783 : node19776;
													assign node19776 = (inp[2]) ? node19780 : node19777;
														assign node19777 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node19780 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node19783 = (inp[6]) ? 16'b0000000000111111 : node19784;
														assign node19784 = (inp[11]) ? 16'b0000000001111111 : node19785;
															assign node19785 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node19790 = (inp[13]) ? node19812 : node19791;
											assign node19791 = (inp[6]) ? node19797 : node19792;
												assign node19792 = (inp[14]) ? 16'b0000000011111111 : node19793;
													assign node19793 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node19797 = (inp[11]) ? node19803 : node19798;
													assign node19798 = (inp[15]) ? node19800 : 16'b0000000011111111;
														assign node19800 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node19803 = (inp[15]) ? node19809 : node19804;
														assign node19804 = (inp[2]) ? 16'b0000000001111111 : node19805;
															assign node19805 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node19809 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node19812 = (inp[15]) ? node19822 : node19813;
												assign node19813 = (inp[9]) ? node19817 : node19814;
													assign node19814 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node19817 = (inp[14]) ? 16'b0000000000111111 : node19818;
														assign node19818 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node19822 = (inp[9]) ? node19826 : node19823;
													assign node19823 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000011111111;
													assign node19826 = (inp[11]) ? node19828 : 16'b0000000000111111;
														assign node19828 = (inp[6]) ? 16'b0000000000011111 : 16'b0000000000111111;
								assign node19831 = (inp[14]) ? node19923 : node19832;
									assign node19832 = (inp[4]) ? node19882 : node19833;
										assign node19833 = (inp[9]) ? node19861 : node19834;
											assign node19834 = (inp[6]) ? node19852 : node19835;
												assign node19835 = (inp[2]) ? node19845 : node19836;
													assign node19836 = (inp[15]) ? 16'b0000001111111111 : node19837;
														assign node19837 = (inp[11]) ? 16'b0000001111111111 : node19838;
															assign node19838 = (inp[12]) ? 16'b0000011111111111 : node19839;
																assign node19839 = (inp[13]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node19845 = (inp[12]) ? node19849 : node19846;
														assign node19846 = (inp[13]) ? 16'b0000000111111111 : 16'b0000011111111111;
														assign node19849 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node19852 = (inp[12]) ? 16'b0000000011111111 : node19853;
													assign node19853 = (inp[2]) ? node19857 : node19854;
														assign node19854 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node19857 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node19861 = (inp[6]) ? node19875 : node19862;
												assign node19862 = (inp[12]) ? node19870 : node19863;
													assign node19863 = (inp[15]) ? node19867 : node19864;
														assign node19864 = (inp[2]) ? 16'b0000000111111111 : 16'b0000011111111111;
														assign node19867 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node19870 = (inp[2]) ? 16'b0000000011111111 : node19871;
														assign node19871 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node19875 = (inp[12]) ? node19879 : node19876;
													assign node19876 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node19879 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node19882 = (inp[6]) ? node19904 : node19883;
											assign node19883 = (inp[9]) ? node19899 : node19884;
												assign node19884 = (inp[15]) ? node19890 : node19885;
													assign node19885 = (inp[13]) ? 16'b0000000111111111 : node19886;
														assign node19886 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node19890 = (inp[11]) ? node19894 : node19891;
														assign node19891 = (inp[12]) ? 16'b0000000111111111 : 16'b0000000011111111;
														assign node19894 = (inp[12]) ? node19896 : 16'b0000000011111111;
															assign node19896 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node19899 = (inp[12]) ? 16'b0000000001111111 : node19900;
													assign node19900 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node19904 = (inp[12]) ? node19912 : node19905;
												assign node19905 = (inp[15]) ? node19907 : 16'b0000000011111111;
													assign node19907 = (inp[9]) ? 16'b0000000001111111 : node19908;
														assign node19908 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node19912 = (inp[15]) ? 16'b0000000000111111 : node19913;
													assign node19913 = (inp[11]) ? node19915 : 16'b0000000011111111;
														assign node19915 = (inp[2]) ? node19917 : 16'b0000000001111111;
															assign node19917 = (inp[9]) ? 16'b0000000000111111 : node19918;
																assign node19918 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node19923 = (inp[6]) ? node19969 : node19924;
										assign node19924 = (inp[11]) ? node19954 : node19925;
											assign node19925 = (inp[12]) ? node19933 : node19926;
												assign node19926 = (inp[9]) ? 16'b0000000011111111 : node19927;
													assign node19927 = (inp[13]) ? 16'b0000000011111111 : node19928;
														assign node19928 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node19933 = (inp[15]) ? node19941 : node19934;
													assign node19934 = (inp[4]) ? node19938 : node19935;
														assign node19935 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node19938 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node19941 = (inp[4]) ? node19947 : node19942;
														assign node19942 = (inp[9]) ? node19944 : 16'b0000000001111111;
															assign node19944 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node19947 = (inp[13]) ? 16'b0000000001111111 : node19948;
															assign node19948 = (inp[9]) ? 16'b0000000001111111 : node19949;
																assign node19949 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node19954 = (inp[13]) ? node19962 : node19955;
												assign node19955 = (inp[9]) ? 16'b0000000001111111 : node19956;
													assign node19956 = (inp[4]) ? node19958 : 16'b0000000011111111;
														assign node19958 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node19962 = (inp[15]) ? node19964 : 16'b0000000001111111;
													assign node19964 = (inp[4]) ? node19966 : 16'b0000000001111111;
														assign node19966 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node19969 = (inp[4]) ? node19989 : node19970;
											assign node19970 = (inp[9]) ? node19978 : node19971;
												assign node19971 = (inp[11]) ? 16'b0000000001111111 : node19972;
													assign node19972 = (inp[15]) ? 16'b0000000011111111 : node19973;
														assign node19973 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node19978 = (inp[11]) ? node19984 : node19979;
													assign node19979 = (inp[12]) ? 16'b0000000001111111 : node19980;
														assign node19980 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node19984 = (inp[12]) ? 16'b0000000000111111 : node19985;
														assign node19985 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node19989 = (inp[12]) ? node19999 : node19990;
												assign node19990 = (inp[15]) ? node19996 : node19991;
													assign node19991 = (inp[9]) ? 16'b0000000000111111 : node19992;
														assign node19992 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node19996 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node19999 = (inp[2]) ? node20009 : node20000;
													assign node20000 = (inp[13]) ? node20002 : 16'b0000000000111111;
														assign node20002 = (inp[15]) ? 16'b0000000000011111 : node20003;
															assign node20003 = (inp[9]) ? node20005 : 16'b0000000000111111;
																assign node20005 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node20009 = (inp[11]) ? node20013 : node20010;
														assign node20010 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node20013 = (inp[9]) ? 16'b0000000000001111 : 16'b0000000000011111;
							assign node20016 = (inp[9]) ? node20176 : node20017;
								assign node20017 = (inp[10]) ? node20095 : node20018;
									assign node20018 = (inp[2]) ? node20058 : node20019;
										assign node20019 = (inp[15]) ? node20049 : node20020;
											assign node20020 = (inp[4]) ? node20038 : node20021;
												assign node20021 = (inp[12]) ? node20031 : node20022;
													assign node20022 = (inp[14]) ? node20024 : 16'b0000001111111111;
														assign node20024 = (inp[11]) ? node20026 : 16'b0000001111111111;
															assign node20026 = (inp[13]) ? node20028 : 16'b0000000111111111;
																assign node20028 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node20031 = (inp[6]) ? node20033 : 16'b0000001111111111;
														assign node20033 = (inp[14]) ? 16'b0000000011111111 : node20034;
															assign node20034 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node20038 = (inp[11]) ? node20044 : node20039;
													assign node20039 = (inp[13]) ? node20041 : 16'b0000000111111111;
														assign node20041 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node20044 = (inp[12]) ? node20046 : 16'b0000000011111111;
														assign node20046 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000011111111;
											assign node20049 = (inp[13]) ? node20055 : node20050;
												assign node20050 = (inp[4]) ? 16'b0000000011111111 : node20051;
													assign node20051 = (inp[12]) ? 16'b0000000111111111 : 16'b0000000011111111;
												assign node20055 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node20058 = (inp[11]) ? node20076 : node20059;
											assign node20059 = (inp[12]) ? node20067 : node20060;
												assign node20060 = (inp[4]) ? node20062 : 16'b0000000111111111;
													assign node20062 = (inp[6]) ? 16'b0000000011111111 : node20063;
														assign node20063 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node20067 = (inp[4]) ? 16'b0000000001111111 : node20068;
													assign node20068 = (inp[13]) ? 16'b0000000011111111 : node20069;
														assign node20069 = (inp[14]) ? node20071 : 16'b0000000111111111;
															assign node20071 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node20076 = (inp[4]) ? node20082 : node20077;
												assign node20077 = (inp[14]) ? 16'b0000000001111111 : node20078;
													assign node20078 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000111111111;
												assign node20082 = (inp[15]) ? node20088 : node20083;
													assign node20083 = (inp[6]) ? 16'b0000000000111111 : node20084;
														assign node20084 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000011111111;
													assign node20088 = (inp[6]) ? node20090 : 16'b0000000000111111;
														assign node20090 = (inp[14]) ? node20092 : 16'b0000000000111111;
															assign node20092 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node20095 = (inp[13]) ? node20137 : node20096;
										assign node20096 = (inp[6]) ? node20114 : node20097;
											assign node20097 = (inp[11]) ? node20107 : node20098;
												assign node20098 = (inp[12]) ? node20104 : node20099;
													assign node20099 = (inp[15]) ? 16'b0000000111111111 : node20100;
														assign node20100 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node20104 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node20107 = (inp[12]) ? node20109 : 16'b0000000011111111;
													assign node20109 = (inp[2]) ? node20111 : 16'b0000000001111111;
														assign node20111 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node20114 = (inp[14]) ? node20126 : node20115;
												assign node20115 = (inp[2]) ? 16'b0000000001111111 : node20116;
													assign node20116 = (inp[12]) ? node20122 : node20117;
														assign node20117 = (inp[11]) ? 16'b0000000011111111 : node20118;
															assign node20118 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node20122 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node20126 = (inp[15]) ? node20132 : node20127;
													assign node20127 = (inp[12]) ? node20129 : 16'b0000000001111111;
														assign node20129 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node20132 = (inp[11]) ? 16'b0000000000111111 : node20133;
														assign node20133 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node20137 = (inp[15]) ? node20163 : node20138;
											assign node20138 = (inp[6]) ? node20152 : node20139;
												assign node20139 = (inp[11]) ? node20147 : node20140;
													assign node20140 = (inp[4]) ? node20144 : node20141;
														assign node20141 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node20144 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node20147 = (inp[4]) ? node20149 : 16'b0000000001111111;
														assign node20149 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000001111111;
												assign node20152 = (inp[12]) ? node20158 : node20153;
													assign node20153 = (inp[4]) ? node20155 : 16'b0000000001111111;
														assign node20155 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node20158 = (inp[4]) ? 16'b0000000000111111 : node20159;
														assign node20159 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node20163 = (inp[2]) ? node20167 : node20164;
												assign node20164 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node20167 = (inp[6]) ? 16'b0000000000000111 : node20168;
													assign node20168 = (inp[14]) ? 16'b0000000000011111 : node20169;
														assign node20169 = (inp[4]) ? node20171 : 16'b0000000000111111;
															assign node20171 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
								assign node20176 = (inp[10]) ? node20274 : node20177;
									assign node20177 = (inp[6]) ? node20231 : node20178;
										assign node20178 = (inp[4]) ? node20202 : node20179;
											assign node20179 = (inp[11]) ? node20191 : node20180;
												assign node20180 = (inp[15]) ? node20186 : node20181;
													assign node20181 = (inp[14]) ? node20183 : 16'b0000000111111111;
														assign node20183 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node20186 = (inp[14]) ? 16'b0000000011111111 : node20187;
														assign node20187 = (inp[12]) ? 16'b0000000011111111 : 16'b0000001111111111;
												assign node20191 = (inp[15]) ? node20193 : 16'b0000000011111111;
													assign node20193 = (inp[14]) ? 16'b0000000000111111 : node20194;
														assign node20194 = (inp[13]) ? 16'b0000000001111111 : node20195;
															assign node20195 = (inp[2]) ? node20197 : 16'b0000000011111111;
																assign node20197 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node20202 = (inp[13]) ? node20216 : node20203;
												assign node20203 = (inp[2]) ? node20209 : node20204;
													assign node20204 = (inp[12]) ? 16'b0000000011111111 : node20205;
														assign node20205 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node20209 = (inp[11]) ? node20213 : node20210;
														assign node20210 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node20213 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node20216 = (inp[11]) ? node20226 : node20217;
													assign node20217 = (inp[14]) ? node20219 : 16'b0000000000111111;
														assign node20219 = (inp[12]) ? 16'b0000000001111111 : node20220;
															assign node20220 = (inp[15]) ? 16'b0000000001111111 : node20221;
																assign node20221 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node20226 = (inp[14]) ? node20228 : 16'b0000000001111111;
														assign node20228 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node20231 = (inp[11]) ? node20251 : node20232;
											assign node20232 = (inp[15]) ? node20240 : node20233;
												assign node20233 = (inp[2]) ? node20235 : 16'b0000000011111111;
													assign node20235 = (inp[14]) ? node20237 : 16'b0000000001111111;
														assign node20237 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node20240 = (inp[4]) ? node20246 : node20241;
													assign node20241 = (inp[13]) ? 16'b0000000001111111 : node20242;
														assign node20242 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node20246 = (inp[14]) ? 16'b0000000000011111 : node20247;
														assign node20247 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node20251 = (inp[15]) ? node20259 : node20252;
												assign node20252 = (inp[4]) ? 16'b0000000000111111 : node20253;
													assign node20253 = (inp[12]) ? node20255 : 16'b0000000001111111;
														assign node20255 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node20259 = (inp[12]) ? node20269 : node20260;
													assign node20260 = (inp[2]) ? node20266 : node20261;
														assign node20261 = (inp[14]) ? 16'b0000000000111111 : node20262;
															assign node20262 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node20266 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node20269 = (inp[2]) ? node20271 : 16'b0000000000011111;
														assign node20271 = (inp[13]) ? 16'b0000000000001111 : 16'b0000000000011111;
									assign node20274 = (inp[11]) ? node20312 : node20275;
										assign node20275 = (inp[15]) ? node20293 : node20276;
											assign node20276 = (inp[6]) ? node20288 : node20277;
												assign node20277 = (inp[2]) ? node20283 : node20278;
													assign node20278 = (inp[4]) ? 16'b0000000011111111 : node20279;
														assign node20279 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node20283 = (inp[4]) ? 16'b0000000001111111 : node20284;
														assign node20284 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node20288 = (inp[4]) ? node20290 : 16'b0000000001111111;
													assign node20290 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000000111111;
											assign node20293 = (inp[2]) ? node20303 : node20294;
												assign node20294 = (inp[4]) ? 16'b0000000000111111 : node20295;
													assign node20295 = (inp[12]) ? node20297 : 16'b0000000001111111;
														assign node20297 = (inp[6]) ? 16'b0000000000111111 : node20298;
															assign node20298 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node20303 = (inp[6]) ? node20309 : node20304;
													assign node20304 = (inp[4]) ? node20306 : 16'b0000000000111111;
														assign node20306 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node20309 = (inp[4]) ? 16'b0000000000000111 : 16'b0000000000011111;
										assign node20312 = (inp[14]) ? node20340 : node20313;
											assign node20313 = (inp[4]) ? node20323 : node20314;
												assign node20314 = (inp[2]) ? 16'b0000000000111111 : node20315;
													assign node20315 = (inp[12]) ? node20319 : node20316;
														assign node20316 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000111111111;
														assign node20319 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node20323 = (inp[15]) ? node20331 : node20324;
													assign node20324 = (inp[2]) ? node20328 : node20325;
														assign node20325 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node20328 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node20331 = (inp[6]) ? node20335 : node20332;
														assign node20332 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000001111111;
														assign node20335 = (inp[12]) ? node20337 : 16'b0000000000011111;
															assign node20337 = (inp[13]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node20340 = (inp[6]) ? node20356 : node20341;
												assign node20341 = (inp[15]) ? node20347 : node20342;
													assign node20342 = (inp[4]) ? 16'b0000000000111111 : node20343;
														assign node20343 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node20347 = (inp[13]) ? node20351 : node20348;
														assign node20348 = (inp[4]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node20351 = (inp[4]) ? 16'b0000000000001111 : node20352;
															assign node20352 = (inp[12]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node20356 = (inp[15]) ? node20364 : node20357;
													assign node20357 = (inp[12]) ? node20359 : 16'b0000000000111111;
														assign node20359 = (inp[13]) ? 16'b0000000000001111 : node20360;
															assign node20360 = (inp[4]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node20364 = (inp[13]) ? node20366 : 16'b0000000000001111;
														assign node20366 = (inp[2]) ? node20368 : 16'b0000000000001111;
															assign node20368 = (inp[12]) ? node20370 : 16'b0000000000000111;
																assign node20370 = (inp[4]) ? 16'b0000000000000011 : 16'b0000000000000111;
						assign node20373 = (inp[14]) ? node20767 : node20374;
							assign node20374 = (inp[13]) ? node20568 : node20375;
								assign node20375 = (inp[11]) ? node20467 : node20376;
									assign node20376 = (inp[2]) ? node20422 : node20377;
										assign node20377 = (inp[4]) ? node20399 : node20378;
											assign node20378 = (inp[10]) ? node20388 : node20379;
												assign node20379 = (inp[6]) ? 16'b0000000111111111 : node20380;
													assign node20380 = (inp[9]) ? node20382 : 16'b0000011111111111;
														assign node20382 = (inp[12]) ? 16'b0000000111111111 : node20383;
															assign node20383 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node20388 = (inp[12]) ? 16'b0000000011111111 : node20389;
													assign node20389 = (inp[6]) ? node20395 : node20390;
														assign node20390 = (inp[3]) ? 16'b0000000111111111 : node20391;
															assign node20391 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node20395 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node20399 = (inp[3]) ? node20411 : node20400;
												assign node20400 = (inp[12]) ? 16'b0000000011111111 : node20401;
													assign node20401 = (inp[15]) ? node20403 : 16'b0000001111111111;
														assign node20403 = (inp[9]) ? node20405 : 16'b0000000111111111;
															assign node20405 = (inp[6]) ? 16'b0000000011111111 : node20406;
																assign node20406 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node20411 = (inp[6]) ? node20413 : 16'b0000000011111111;
													assign node20413 = (inp[9]) ? node20419 : node20414;
														assign node20414 = (inp[10]) ? node20416 : 16'b0000000011111111;
															assign node20416 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node20419 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node20422 = (inp[15]) ? node20442 : node20423;
											assign node20423 = (inp[10]) ? node20431 : node20424;
												assign node20424 = (inp[3]) ? node20426 : 16'b0000000111111111;
													assign node20426 = (inp[4]) ? 16'b0000000011111111 : node20427;
														assign node20427 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000111111111;
												assign node20431 = (inp[9]) ? 16'b0000000000011111 : node20432;
													assign node20432 = (inp[4]) ? node20434 : 16'b0000000011111111;
														assign node20434 = (inp[3]) ? node20436 : 16'b0000000011111111;
															assign node20436 = (inp[12]) ? 16'b0000000001111111 : node20437;
																assign node20437 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node20442 = (inp[12]) ? node20452 : node20443;
												assign node20443 = (inp[6]) ? node20447 : node20444;
													assign node20444 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000111111111;
													assign node20447 = (inp[4]) ? 16'b0000000001111111 : node20448;
														assign node20448 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node20452 = (inp[3]) ? node20456 : node20453;
													assign node20453 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node20456 = (inp[9]) ? node20458 : 16'b0000000000111111;
														assign node20458 = (inp[4]) ? node20464 : node20459;
															assign node20459 = (inp[10]) ? node20461 : 16'b0000000000111111;
																assign node20461 = (inp[6]) ? 16'b0000000000011111 : 16'b0000000000111111;
															assign node20464 = (inp[10]) ? 16'b0000000000001111 : 16'b0000000000011111;
									assign node20467 = (inp[10]) ? node20517 : node20468;
										assign node20468 = (inp[3]) ? node20488 : node20469;
											assign node20469 = (inp[12]) ? node20477 : node20470;
												assign node20470 = (inp[15]) ? node20472 : 16'b0000000111111111;
													assign node20472 = (inp[9]) ? 16'b0000000011111111 : node20473;
														assign node20473 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node20477 = (inp[6]) ? node20485 : node20478;
													assign node20478 = (inp[2]) ? node20482 : node20479;
														assign node20479 = (inp[4]) ? 16'b0000000111111111 : 16'b0000000011111111;
														assign node20482 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node20485 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node20488 = (inp[9]) ? node20510 : node20489;
												assign node20489 = (inp[6]) ? node20499 : node20490;
													assign node20490 = (inp[2]) ? node20494 : node20491;
														assign node20491 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node20494 = (inp[12]) ? 16'b0000000000111111 : node20495;
															assign node20495 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node20499 = (inp[15]) ? node20505 : node20500;
														assign node20500 = (inp[4]) ? 16'b0000000001111111 : node20501;
															assign node20501 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node20505 = (inp[4]) ? node20507 : 16'b0000000001111111;
															assign node20507 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node20510 = (inp[6]) ? node20514 : node20511;
													assign node20511 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000000111111;
													assign node20514 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node20517 = (inp[12]) ? node20539 : node20518;
											assign node20518 = (inp[9]) ? node20530 : node20519;
												assign node20519 = (inp[3]) ? node20525 : node20520;
													assign node20520 = (inp[15]) ? node20522 : 16'b0000000111111111;
														assign node20522 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node20525 = (inp[6]) ? node20527 : 16'b0000000001111111;
														assign node20527 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node20530 = (inp[15]) ? 16'b0000000000111111 : node20531;
													assign node20531 = (inp[4]) ? node20535 : node20532;
														assign node20532 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node20535 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node20539 = (inp[15]) ? node20553 : node20540;
												assign node20540 = (inp[6]) ? node20546 : node20541;
													assign node20541 = (inp[4]) ? node20543 : 16'b0000000011111111;
														assign node20543 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node20546 = (inp[4]) ? 16'b0000000000011111 : node20547;
														assign node20547 = (inp[3]) ? 16'b0000000000111111 : node20548;
															assign node20548 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node20553 = (inp[3]) ? node20559 : node20554;
													assign node20554 = (inp[4]) ? node20556 : 16'b0000000001111111;
														assign node20556 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node20559 = (inp[9]) ? node20565 : node20560;
														assign node20560 = (inp[6]) ? 16'b0000000000011111 : node20561;
															assign node20561 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node20565 = (inp[4]) ? 16'b0000000000001111 : 16'b0000000000011111;
								assign node20568 = (inp[11]) ? node20674 : node20569;
									assign node20569 = (inp[6]) ? node20627 : node20570;
										assign node20570 = (inp[4]) ? node20592 : node20571;
											assign node20571 = (inp[10]) ? node20579 : node20572;
												assign node20572 = (inp[12]) ? 16'b0000000011111111 : node20573;
													assign node20573 = (inp[9]) ? node20575 : 16'b0000011111111111;
														assign node20575 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node20579 = (inp[3]) ? node20585 : node20580;
													assign node20580 = (inp[9]) ? node20582 : 16'b0000000011111111;
														assign node20582 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node20585 = (inp[2]) ? 16'b0000000001111111 : node20586;
														assign node20586 = (inp[15]) ? 16'b0000000001111111 : node20587;
															assign node20587 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node20592 = (inp[15]) ? node20612 : node20593;
												assign node20593 = (inp[2]) ? node20605 : node20594;
													assign node20594 = (inp[9]) ? node20598 : node20595;
														assign node20595 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node20598 = (inp[10]) ? node20600 : 16'b0000000011111111;
															assign node20600 = (inp[3]) ? 16'b0000000001111111 : node20601;
																assign node20601 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node20605 = (inp[3]) ? 16'b0000000000111111 : node20606;
														assign node20606 = (inp[10]) ? 16'b0000000001111111 : node20607;
															assign node20607 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node20612 = (inp[12]) ? node20622 : node20613;
													assign node20613 = (inp[9]) ? node20615 : 16'b0000000011111111;
														assign node20615 = (inp[3]) ? 16'b0000000000111111 : node20616;
															assign node20616 = (inp[10]) ? node20618 : 16'b0000000001111111;
																assign node20618 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node20622 = (inp[10]) ? 16'b0000000000011111 : node20623;
														assign node20623 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node20627 = (inp[9]) ? node20647 : node20628;
											assign node20628 = (inp[12]) ? node20638 : node20629;
												assign node20629 = (inp[3]) ? 16'b0000000001111111 : node20630;
													assign node20630 = (inp[15]) ? 16'b0000000011111111 : node20631;
														assign node20631 = (inp[10]) ? node20633 : 16'b0000000111111111;
															assign node20633 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node20638 = (inp[3]) ? node20644 : node20639;
													assign node20639 = (inp[10]) ? node20641 : 16'b0000000001111111;
														assign node20641 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000000111111;
													assign node20644 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node20647 = (inp[4]) ? node20663 : node20648;
												assign node20648 = (inp[10]) ? node20658 : node20649;
													assign node20649 = (inp[12]) ? node20651 : 16'b0000000001111111;
														assign node20651 = (inp[15]) ? node20653 : 16'b0000000001111111;
															assign node20653 = (inp[2]) ? 16'b0000000000111111 : node20654;
																assign node20654 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node20658 = (inp[3]) ? 16'b0000000000011111 : node20659;
														assign node20659 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node20663 = (inp[12]) ? node20671 : node20664;
													assign node20664 = (inp[2]) ? 16'b0000000000011111 : node20665;
														assign node20665 = (inp[15]) ? 16'b0000000000111111 : node20666;
															assign node20666 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node20671 = (inp[10]) ? 16'b0000000000001111 : 16'b0000000000011111;
									assign node20674 = (inp[3]) ? node20730 : node20675;
										assign node20675 = (inp[2]) ? node20703 : node20676;
											assign node20676 = (inp[6]) ? node20690 : node20677;
												assign node20677 = (inp[15]) ? node20683 : node20678;
													assign node20678 = (inp[12]) ? node20680 : 16'b0000000011111111;
														assign node20680 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node20683 = (inp[12]) ? 16'b0000000001111111 : node20684;
														assign node20684 = (inp[10]) ? 16'b0000000001111111 : node20685;
															assign node20685 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node20690 = (inp[15]) ? node20696 : node20691;
													assign node20691 = (inp[9]) ? 16'b0000000000111111 : node20692;
														assign node20692 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node20696 = (inp[10]) ? 16'b0000000000011111 : node20697;
														assign node20697 = (inp[4]) ? 16'b0000000000111111 : node20698;
															assign node20698 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node20703 = (inp[4]) ? node20713 : node20704;
												assign node20704 = (inp[9]) ? node20710 : node20705;
													assign node20705 = (inp[6]) ? node20707 : 16'b0000000001111111;
														assign node20707 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node20710 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000000011111;
												assign node20713 = (inp[6]) ? node20723 : node20714;
													assign node20714 = (inp[15]) ? node20720 : node20715;
														assign node20715 = (inp[10]) ? 16'b0000000000111111 : node20716;
															assign node20716 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node20720 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node20723 = (inp[10]) ? node20727 : node20724;
														assign node20724 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000000011111;
														assign node20727 = (inp[12]) ? 16'b0000000000001111 : 16'b0000000000011111;
										assign node20730 = (inp[12]) ? node20750 : node20731;
											assign node20731 = (inp[15]) ? node20739 : node20732;
												assign node20732 = (inp[10]) ? 16'b0000000000111111 : node20733;
													assign node20733 = (inp[4]) ? node20735 : 16'b0000000011111111;
														assign node20735 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node20739 = (inp[4]) ? node20745 : node20740;
													assign node20740 = (inp[2]) ? 16'b0000000000011111 : node20741;
														assign node20741 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node20745 = (inp[6]) ? node20747 : 16'b0000000000011111;
														assign node20747 = (inp[9]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node20750 = (inp[4]) ? node20760 : node20751;
												assign node20751 = (inp[6]) ? 16'b0000000000001111 : node20752;
													assign node20752 = (inp[2]) ? node20754 : 16'b0000000000111111;
														assign node20754 = (inp[9]) ? 16'b0000000000011111 : node20755;
															assign node20755 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node20760 = (inp[2]) ? node20764 : node20761;
													assign node20761 = (inp[6]) ? 16'b0000000000011111 : 16'b0000000000001111;
													assign node20764 = (inp[15]) ? 16'b0000000000000111 : 16'b0000000000001111;
							assign node20767 = (inp[9]) ? node20949 : node20768;
								assign node20768 = (inp[2]) ? node20862 : node20769;
									assign node20769 = (inp[12]) ? node20815 : node20770;
										assign node20770 = (inp[15]) ? node20794 : node20771;
											assign node20771 = (inp[10]) ? node20777 : node20772;
												assign node20772 = (inp[6]) ? 16'b0000000011111111 : node20773;
													assign node20773 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node20777 = (inp[13]) ? node20785 : node20778;
													assign node20778 = (inp[3]) ? node20780 : 16'b0000000111111111;
														assign node20780 = (inp[6]) ? node20782 : 16'b0000000011111111;
															assign node20782 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node20785 = (inp[6]) ? 16'b0000000001111111 : node20786;
														assign node20786 = (inp[4]) ? node20788 : 16'b0000000011111111;
															assign node20788 = (inp[3]) ? 16'b0000000001111111 : node20789;
																assign node20789 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node20794 = (inp[10]) ? node20802 : node20795;
												assign node20795 = (inp[13]) ? node20797 : 16'b0000000011111111;
													assign node20797 = (inp[3]) ? 16'b0000000001111111 : node20798;
														assign node20798 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node20802 = (inp[13]) ? node20808 : node20803;
													assign node20803 = (inp[11]) ? node20805 : 16'b0000000011111111;
														assign node20805 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node20808 = (inp[4]) ? node20810 : 16'b0000000001111111;
														assign node20810 = (inp[11]) ? 16'b0000000000011111 : node20811;
															assign node20811 = (inp[6]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node20815 = (inp[3]) ? node20835 : node20816;
											assign node20816 = (inp[4]) ? node20824 : node20817;
												assign node20817 = (inp[13]) ? node20819 : 16'b0000000011111111;
													assign node20819 = (inp[6]) ? 16'b0000000001111111 : node20820;
														assign node20820 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node20824 = (inp[10]) ? 16'b0000000000111111 : node20825;
													assign node20825 = (inp[15]) ? node20827 : 16'b0000000001111111;
														assign node20827 = (inp[13]) ? 16'b0000000000111111 : node20828;
															assign node20828 = (inp[11]) ? 16'b0000000000111111 : node20829;
																assign node20829 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node20835 = (inp[13]) ? node20847 : node20836;
												assign node20836 = (inp[4]) ? node20840 : node20837;
													assign node20837 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node20840 = (inp[15]) ? node20844 : node20841;
														assign node20841 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node20844 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node20847 = (inp[6]) ? node20849 : 16'b0000000000111111;
													assign node20849 = (inp[4]) ? node20853 : node20850;
														assign node20850 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node20853 = (inp[15]) ? node20857 : node20854;
															assign node20854 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000111111;
															assign node20857 = (inp[10]) ? 16'b0000000000001111 : node20858;
																assign node20858 = (inp[11]) ? 16'b0000000000001111 : 16'b0000000000011111;
									assign node20862 = (inp[11]) ? node20900 : node20863;
										assign node20863 = (inp[13]) ? node20881 : node20864;
											assign node20864 = (inp[10]) ? node20872 : node20865;
												assign node20865 = (inp[4]) ? node20869 : node20866;
													assign node20866 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node20869 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000001111111;
												assign node20872 = (inp[6]) ? 16'b0000000000111111 : node20873;
													assign node20873 = (inp[3]) ? node20877 : node20874;
														assign node20874 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000011111111;
														assign node20877 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node20881 = (inp[6]) ? node20891 : node20882;
												assign node20882 = (inp[12]) ? node20884 : 16'b0000000000111111;
													assign node20884 = (inp[15]) ? 16'b0000000000111111 : node20885;
														assign node20885 = (inp[3]) ? node20887 : 16'b0000000001111111;
															assign node20887 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node20891 = (inp[10]) ? 16'b0000000000011111 : node20892;
													assign node20892 = (inp[3]) ? 16'b0000000000111111 : node20893;
														assign node20893 = (inp[12]) ? node20895 : 16'b0000000000111111;
															assign node20895 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node20900 = (inp[10]) ? node20922 : node20901;
											assign node20901 = (inp[3]) ? node20913 : node20902;
												assign node20902 = (inp[13]) ? node20906 : node20903;
													assign node20903 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node20906 = (inp[12]) ? 16'b0000000000111111 : node20907;
														assign node20907 = (inp[4]) ? node20909 : 16'b0000000001111111;
															assign node20909 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node20913 = (inp[13]) ? 16'b0000000000011111 : node20914;
													assign node20914 = (inp[6]) ? 16'b0000000000011111 : node20915;
														assign node20915 = (inp[15]) ? node20917 : 16'b0000000001111111;
															assign node20917 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node20922 = (inp[3]) ? node20934 : node20923;
												assign node20923 = (inp[6]) ? 16'b0000000000011111 : node20924;
													assign node20924 = (inp[13]) ? node20926 : 16'b0000000000111111;
														assign node20926 = (inp[12]) ? node20928 : 16'b0000000000111111;
															assign node20928 = (inp[15]) ? 16'b0000000000011111 : node20929;
																assign node20929 = (inp[4]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node20934 = (inp[6]) ? node20944 : node20935;
													assign node20935 = (inp[4]) ? node20939 : node20936;
														assign node20936 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node20939 = (inp[13]) ? node20941 : 16'b0000000000011111;
															assign node20941 = (inp[12]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node20944 = (inp[12]) ? 16'b0000000000001111 : node20945;
														assign node20945 = (inp[4]) ? 16'b0000000000000111 : 16'b0000000000001111;
								assign node20949 = (inp[11]) ? node21033 : node20950;
									assign node20950 = (inp[2]) ? node20986 : node20951;
										assign node20951 = (inp[3]) ? node20967 : node20952;
											assign node20952 = (inp[15]) ? node20958 : node20953;
												assign node20953 = (inp[10]) ? node20955 : 16'b0000000011111111;
													assign node20955 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node20958 = (inp[10]) ? node20962 : node20959;
													assign node20959 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node20962 = (inp[12]) ? 16'b0000000000111111 : node20963;
														assign node20963 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node20967 = (inp[13]) ? node20977 : node20968;
												assign node20968 = (inp[12]) ? 16'b0000000000111111 : node20969;
													assign node20969 = (inp[10]) ? node20971 : 16'b0000000111111111;
														assign node20971 = (inp[4]) ? node20973 : 16'b0000000001111111;
															assign node20973 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node20977 = (inp[12]) ? 16'b0000000000011111 : node20978;
													assign node20978 = (inp[6]) ? node20980 : 16'b0000000000111111;
														assign node20980 = (inp[10]) ? 16'b0000000000011111 : node20981;
															assign node20981 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node20986 = (inp[4]) ? node21014 : node20987;
											assign node20987 = (inp[6]) ? node21005 : node20988;
												assign node20988 = (inp[15]) ? node20996 : node20989;
													assign node20989 = (inp[3]) ? node20991 : 16'b0000000011111111;
														assign node20991 = (inp[13]) ? node20993 : 16'b0000000001111111;
															assign node20993 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node20996 = (inp[3]) ? node21002 : node20997;
														assign node20997 = (inp[12]) ? node20999 : 16'b0000000001111111;
															assign node20999 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node21002 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node21005 = (inp[12]) ? node21007 : 16'b0000000000111111;
													assign node21007 = (inp[3]) ? node21009 : 16'b0000000000111111;
														assign node21009 = (inp[10]) ? 16'b0000000000001111 : node21010;
															assign node21010 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node21014 = (inp[15]) ? node21024 : node21015;
												assign node21015 = (inp[10]) ? node21017 : 16'b0000000000111111;
													assign node21017 = (inp[12]) ? 16'b0000000000001111 : node21018;
														assign node21018 = (inp[6]) ? 16'b0000000000011111 : node21019;
															assign node21019 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node21024 = (inp[12]) ? node21030 : node21025;
													assign node21025 = (inp[10]) ? node21027 : 16'b0000000000011111;
														assign node21027 = (inp[6]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node21030 = (inp[13]) ? 16'b0000000000000111 : 16'b0000000000001111;
									assign node21033 = (inp[13]) ? node21077 : node21034;
										assign node21034 = (inp[6]) ? node21048 : node21035;
											assign node21035 = (inp[10]) ? node21043 : node21036;
												assign node21036 = (inp[15]) ? node21038 : 16'b0000000001111111;
													assign node21038 = (inp[3]) ? 16'b0000000001111111 : node21039;
														assign node21039 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node21043 = (inp[15]) ? node21045 : 16'b0000000000111111;
													assign node21045 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node21048 = (inp[12]) ? node21062 : node21049;
												assign node21049 = (inp[2]) ? node21057 : node21050;
													assign node21050 = (inp[15]) ? node21054 : node21051;
														assign node21051 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node21054 = (inp[4]) ? 16'b0000000000001111 : 16'b0000000000111111;
													assign node21057 = (inp[3]) ? node21059 : 16'b0000000000011111;
														assign node21059 = (inp[10]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node21062 = (inp[15]) ? node21074 : node21063;
													assign node21063 = (inp[4]) ? node21067 : node21064;
														assign node21064 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node21067 = (inp[2]) ? 16'b0000000000001111 : node21068;
															assign node21068 = (inp[3]) ? node21070 : 16'b0000000000011111;
																assign node21070 = (inp[10]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node21074 = (inp[3]) ? 16'b0000000000000111 : 16'b0000000000001111;
										assign node21077 = (inp[3]) ? node21107 : node21078;
											assign node21078 = (inp[4]) ? node21094 : node21079;
												assign node21079 = (inp[15]) ? node21085 : node21080;
													assign node21080 = (inp[10]) ? node21082 : 16'b0000000000111111;
														assign node21082 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node21085 = (inp[2]) ? node21087 : 16'b0000000000111111;
														assign node21087 = (inp[6]) ? 16'b0000000000001111 : node21088;
															assign node21088 = (inp[10]) ? node21090 : 16'b0000000000011111;
																assign node21090 = (inp[12]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node21094 = (inp[12]) ? node21100 : node21095;
													assign node21095 = (inp[6]) ? node21097 : 16'b0000000000011111;
														assign node21097 = (inp[2]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node21100 = (inp[10]) ? 16'b0000000000000111 : node21101;
														assign node21101 = (inp[2]) ? 16'b0000000000001111 : node21102;
															assign node21102 = (inp[6]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node21107 = (inp[15]) ? node21123 : node21108;
												assign node21108 = (inp[12]) ? node21116 : node21109;
													assign node21109 = (inp[6]) ? node21113 : node21110;
														assign node21110 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node21113 = (inp[2]) ? 16'b0000000000000111 : 16'b0000000000001111;
													assign node21116 = (inp[10]) ? 16'b0000000000001111 : node21117;
														assign node21117 = (inp[2]) ? 16'b0000000000001111 : node21118;
															assign node21118 = (inp[4]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node21123 = (inp[10]) ? node21127 : node21124;
													assign node21124 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000001111;
													assign node21127 = (inp[12]) ? node21129 : 16'b0000000000000111;
														assign node21129 = (inp[6]) ? 16'b0000000000000011 : 16'b0000000000000111;
				assign node21132 = (inp[4]) ? node22738 : node21133;
					assign node21133 = (inp[14]) ? node21913 : node21134;
						assign node21134 = (inp[12]) ? node21506 : node21135;
							assign node21135 = (inp[3]) ? node21313 : node21136;
								assign node21136 = (inp[2]) ? node21222 : node21137;
									assign node21137 = (inp[9]) ? node21183 : node21138;
										assign node21138 = (inp[5]) ? node21164 : node21139;
											assign node21139 = (inp[15]) ? node21151 : node21140;
												assign node21140 = (inp[6]) ? node21142 : 16'b0000011111111111;
													assign node21142 = (inp[13]) ? node21144 : 16'b0000011111111111;
														assign node21144 = (inp[11]) ? 16'b0000001111111111 : node21145;
															assign node21145 = (inp[10]) ? 16'b0000001111111111 : node21146;
																assign node21146 = (inp[1]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node21151 = (inp[11]) ? node21159 : node21152;
													assign node21152 = (inp[6]) ? node21156 : node21153;
														assign node21153 = (inp[10]) ? 16'b0000001111111111 : 16'b0000111111111111;
														assign node21156 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node21159 = (inp[1]) ? 16'b0000000111111111 : node21160;
														assign node21160 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node21164 = (inp[1]) ? node21172 : node21165;
												assign node21165 = (inp[15]) ? 16'b0000000111111111 : node21166;
													assign node21166 = (inp[13]) ? node21168 : 16'b0000001111111111;
														assign node21168 = (inp[11]) ? 16'b0000001111111111 : 16'b0000000111111111;
												assign node21172 = (inp[13]) ? 16'b0000000011111111 : node21173;
													assign node21173 = (inp[11]) ? node21177 : node21174;
														assign node21174 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node21177 = (inp[6]) ? node21179 : 16'b0000000111111111;
															assign node21179 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node21183 = (inp[1]) ? node21205 : node21184;
											assign node21184 = (inp[11]) ? node21186 : 16'b0000001111111111;
												assign node21186 = (inp[6]) ? node21196 : node21187;
													assign node21187 = (inp[13]) ? node21193 : node21188;
														assign node21188 = (inp[15]) ? 16'b0000001111111111 : node21189;
															assign node21189 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node21193 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node21196 = (inp[10]) ? node21202 : node21197;
														assign node21197 = (inp[13]) ? node21199 : 16'b0000000111111111;
															assign node21199 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node21202 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000001111111;
											assign node21205 = (inp[10]) ? node21213 : node21206;
												assign node21206 = (inp[13]) ? 16'b0000000011111111 : node21207;
													assign node21207 = (inp[15]) ? 16'b0000000011111111 : node21208;
														assign node21208 = (inp[5]) ? 16'b0000001111111111 : 16'b0000000111111111;
												assign node21213 = (inp[13]) ? node21215 : 16'b0000000011111111;
													assign node21215 = (inp[15]) ? node21219 : node21216;
														assign node21216 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000001111111;
														assign node21219 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node21222 = (inp[13]) ? node21266 : node21223;
										assign node21223 = (inp[1]) ? node21247 : node21224;
											assign node21224 = (inp[6]) ? node21232 : node21225;
												assign node21225 = (inp[5]) ? 16'b0000000111111111 : node21226;
													assign node21226 = (inp[9]) ? 16'b0000001111111111 : node21227;
														assign node21227 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node21232 = (inp[11]) ? node21236 : node21233;
													assign node21233 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node21236 = (inp[15]) ? node21242 : node21237;
														assign node21237 = (inp[5]) ? node21239 : 16'b0000000111111111;
															assign node21239 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node21242 = (inp[9]) ? node21244 : 16'b0000000011111111;
															assign node21244 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node21247 = (inp[11]) ? node21255 : node21248;
												assign node21248 = (inp[15]) ? 16'b0000000011111111 : node21249;
													assign node21249 = (inp[10]) ? node21251 : 16'b0000000111111111;
														assign node21251 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node21255 = (inp[5]) ? node21259 : node21256;
													assign node21256 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node21259 = (inp[9]) ? node21261 : 16'b0000000011111111;
														assign node21261 = (inp[10]) ? node21263 : 16'b0000000001111111;
															assign node21263 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node21266 = (inp[1]) ? node21292 : node21267;
											assign node21267 = (inp[15]) ? node21283 : node21268;
												assign node21268 = (inp[11]) ? node21276 : node21269;
													assign node21269 = (inp[5]) ? node21271 : 16'b0000000111111111;
														assign node21271 = (inp[9]) ? 16'b0000000011111111 : node21272;
															assign node21272 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node21276 = (inp[10]) ? node21278 : 16'b0000001111111111;
														assign node21278 = (inp[6]) ? node21280 : 16'b0000000011111111;
															assign node21280 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node21283 = (inp[6]) ? node21285 : 16'b0000000011111111;
													assign node21285 = (inp[9]) ? node21287 : 16'b0000000011111111;
														assign node21287 = (inp[5]) ? 16'b0000000001111111 : node21288;
															assign node21288 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node21292 = (inp[9]) ? node21304 : node21293;
												assign node21293 = (inp[5]) ? node21299 : node21294;
													assign node21294 = (inp[11]) ? node21296 : 16'b0000000111111111;
														assign node21296 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node21299 = (inp[10]) ? 16'b0000000001111111 : node21300;
														assign node21300 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node21304 = (inp[5]) ? 16'b0000000000001111 : node21305;
													assign node21305 = (inp[11]) ? node21309 : node21306;
														assign node21306 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node21309 = (inp[6]) ? 16'b0000000000011111 : 16'b0000000001111111;
								assign node21313 = (inp[9]) ? node21429 : node21314;
									assign node21314 = (inp[15]) ? node21366 : node21315;
										assign node21315 = (inp[1]) ? node21341 : node21316;
											assign node21316 = (inp[13]) ? node21330 : node21317;
												assign node21317 = (inp[10]) ? node21323 : node21318;
													assign node21318 = (inp[5]) ? 16'b0000001111111111 : node21319;
														assign node21319 = (inp[11]) ? 16'b0000001111111111 : 16'b0000111111111111;
													assign node21323 = (inp[2]) ? 16'b0000000111111111 : node21324;
														assign node21324 = (inp[11]) ? 16'b0000000111111111 : node21325;
															assign node21325 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node21330 = (inp[5]) ? 16'b0000000011111111 : node21331;
													assign node21331 = (inp[6]) ? node21333 : 16'b0000001111111111;
														assign node21333 = (inp[10]) ? 16'b0000000011111111 : node21334;
															assign node21334 = (inp[11]) ? node21336 : 16'b0000000111111111;
																assign node21336 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node21341 = (inp[10]) ? node21349 : node21342;
												assign node21342 = (inp[11]) ? 16'b0000000011111111 : node21343;
													assign node21343 = (inp[6]) ? node21345 : 16'b0000000111111111;
														assign node21345 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node21349 = (inp[5]) ? node21361 : node21350;
													assign node21350 = (inp[13]) ? node21356 : node21351;
														assign node21351 = (inp[6]) ? 16'b0000000011111111 : node21352;
															assign node21352 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node21356 = (inp[6]) ? node21358 : 16'b0000000011111111;
															assign node21358 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node21361 = (inp[6]) ? node21363 : 16'b0000000001111111;
														assign node21363 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node21366 = (inp[5]) ? node21398 : node21367;
											assign node21367 = (inp[10]) ? node21381 : node21368;
												assign node21368 = (inp[13]) ? node21374 : node21369;
													assign node21369 = (inp[1]) ? 16'b0000000001111111 : node21370;
														assign node21370 = (inp[11]) ? 16'b0000001111111111 : 16'b0000000111111111;
													assign node21374 = (inp[1]) ? node21376 : 16'b0000000011111111;
														assign node21376 = (inp[2]) ? 16'b0000000011111111 : node21377;
															assign node21377 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node21381 = (inp[13]) ? node21393 : node21382;
													assign node21382 = (inp[2]) ? node21384 : 16'b0000000111111111;
														assign node21384 = (inp[6]) ? node21388 : node21385;
															assign node21385 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
															assign node21388 = (inp[1]) ? 16'b0000000001111111 : node21389;
																assign node21389 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node21393 = (inp[1]) ? 16'b0000000001111111 : node21394;
														assign node21394 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node21398 = (inp[2]) ? node21416 : node21399;
												assign node21399 = (inp[1]) ? node21407 : node21400;
													assign node21400 = (inp[6]) ? node21404 : node21401;
														assign node21401 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node21404 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node21407 = (inp[6]) ? node21413 : node21408;
														assign node21408 = (inp[11]) ? node21410 : 16'b0000000001111111;
															assign node21410 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node21413 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node21416 = (inp[1]) ? node21426 : node21417;
													assign node21417 = (inp[6]) ? node21421 : node21418;
														assign node21418 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node21421 = (inp[13]) ? node21423 : 16'b0000000001111111;
															assign node21423 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node21426 = (inp[6]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node21429 = (inp[6]) ? node21465 : node21430;
										assign node21430 = (inp[1]) ? node21448 : node21431;
											assign node21431 = (inp[15]) ? node21435 : node21432;
												assign node21432 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node21435 = (inp[2]) ? node21441 : node21436;
													assign node21436 = (inp[13]) ? 16'b0000000011111111 : node21437;
														assign node21437 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node21441 = (inp[13]) ? node21443 : 16'b0000000011111111;
														assign node21443 = (inp[5]) ? 16'b0000000001111111 : node21444;
															assign node21444 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node21448 = (inp[5]) ? node21456 : node21449;
												assign node21449 = (inp[11]) ? 16'b0000000001111111 : node21450;
													assign node21450 = (inp[15]) ? 16'b0000000011111111 : node21451;
														assign node21451 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node21456 = (inp[11]) ? node21462 : node21457;
													assign node21457 = (inp[13]) ? node21459 : 16'b0000000000111111;
														assign node21459 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node21462 = (inp[2]) ? 16'b0000000000001111 : 16'b0000000000011111;
										assign node21465 = (inp[11]) ? node21487 : node21466;
											assign node21466 = (inp[2]) ? node21478 : node21467;
												assign node21467 = (inp[1]) ? node21475 : node21468;
													assign node21468 = (inp[13]) ? node21472 : node21469;
														assign node21469 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node21472 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node21475 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node21478 = (inp[5]) ? node21484 : node21479;
													assign node21479 = (inp[13]) ? 16'b0000000000111111 : node21480;
														assign node21480 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node21484 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node21487 = (inp[1]) ? node21499 : node21488;
												assign node21488 = (inp[13]) ? 16'b0000000000111111 : node21489;
													assign node21489 = (inp[15]) ? node21491 : 16'b0000000001111111;
														assign node21491 = (inp[10]) ? node21495 : node21492;
															assign node21492 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
															assign node21495 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node21499 = (inp[5]) ? node21501 : 16'b0000000000111111;
													assign node21501 = (inp[13]) ? node21503 : 16'b0000000000011111;
														assign node21503 = (inp[10]) ? 16'b0000000000001111 : 16'b0000000000011111;
							assign node21506 = (inp[6]) ? node21710 : node21507;
								assign node21507 = (inp[3]) ? node21597 : node21508;
									assign node21508 = (inp[15]) ? node21554 : node21509;
										assign node21509 = (inp[2]) ? node21525 : node21510;
											assign node21510 = (inp[9]) ? node21518 : node21511;
												assign node21511 = (inp[11]) ? node21513 : 16'b0000001111111111;
													assign node21513 = (inp[5]) ? 16'b0000000111111111 : node21514;
														assign node21514 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node21518 = (inp[1]) ? node21520 : 16'b0000000111111111;
													assign node21520 = (inp[10]) ? node21522 : 16'b0000000111111111;
														assign node21522 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node21525 = (inp[10]) ? node21547 : node21526;
												assign node21526 = (inp[13]) ? node21536 : node21527;
													assign node21527 = (inp[11]) ? node21533 : node21528;
														assign node21528 = (inp[5]) ? 16'b0000000111111111 : node21529;
															assign node21529 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node21533 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node21536 = (inp[11]) ? node21544 : node21537;
														assign node21537 = (inp[9]) ? node21539 : 16'b0000000111111111;
															assign node21539 = (inp[1]) ? 16'b0000000011111111 : node21540;
																assign node21540 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node21544 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node21547 = (inp[5]) ? node21549 : 16'b0000000011111111;
													assign node21549 = (inp[11]) ? 16'b0000000000111111 : node21550;
														assign node21550 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000111111111;
										assign node21554 = (inp[2]) ? node21576 : node21555;
											assign node21555 = (inp[9]) ? node21569 : node21556;
												assign node21556 = (inp[5]) ? node21558 : 16'b0000000111111111;
													assign node21558 = (inp[13]) ? node21566 : node21559;
														assign node21559 = (inp[11]) ? node21561 : 16'b0000000111111111;
															assign node21561 = (inp[1]) ? 16'b0000000011111111 : node21562;
																assign node21562 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node21566 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node21569 = (inp[11]) ? 16'b0000000001111111 : node21570;
													assign node21570 = (inp[1]) ? node21572 : 16'b0000000111111111;
														assign node21572 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node21576 = (inp[1]) ? node21590 : node21577;
												assign node21577 = (inp[10]) ? node21583 : node21578;
													assign node21578 = (inp[9]) ? node21580 : 16'b0000000011111111;
														assign node21580 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node21583 = (inp[9]) ? node21587 : node21584;
														assign node21584 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node21587 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node21590 = (inp[5]) ? node21592 : 16'b0000000001111111;
													assign node21592 = (inp[11]) ? 16'b0000000000111111 : node21593;
														assign node21593 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node21597 = (inp[5]) ? node21649 : node21598;
										assign node21598 = (inp[10]) ? node21620 : node21599;
											assign node21599 = (inp[9]) ? node21607 : node21600;
												assign node21600 = (inp[15]) ? node21604 : node21601;
													assign node21601 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node21604 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node21607 = (inp[15]) ? node21615 : node21608;
													assign node21608 = (inp[1]) ? 16'b0000000011111111 : node21609;
														assign node21609 = (inp[13]) ? 16'b0000000011111111 : node21610;
															assign node21610 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node21615 = (inp[1]) ? 16'b0000000001111111 : node21616;
														assign node21616 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node21620 = (inp[9]) ? node21634 : node21621;
												assign node21621 = (inp[15]) ? node21631 : node21622;
													assign node21622 = (inp[2]) ? 16'b0000000011111111 : node21623;
														assign node21623 = (inp[1]) ? node21625 : 16'b0000000111111111;
															assign node21625 = (inp[13]) ? 16'b0000000011111111 : node21626;
																assign node21626 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node21631 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000011111111;
												assign node21634 = (inp[2]) ? node21642 : node21635;
													assign node21635 = (inp[1]) ? node21639 : node21636;
														assign node21636 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node21639 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node21642 = (inp[1]) ? node21644 : 16'b0000000000111111;
														assign node21644 = (inp[13]) ? 16'b0000000000001111 : node21645;
															assign node21645 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node21649 = (inp[10]) ? node21679 : node21650;
											assign node21650 = (inp[15]) ? node21662 : node21651;
												assign node21651 = (inp[9]) ? node21657 : node21652;
													assign node21652 = (inp[2]) ? 16'b0000000011111111 : node21653;
														assign node21653 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node21657 = (inp[1]) ? 16'b0000000001111111 : node21658;
														assign node21658 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node21662 = (inp[13]) ? node21670 : node21663;
													assign node21663 = (inp[2]) ? node21665 : 16'b0000000001111111;
														assign node21665 = (inp[1]) ? node21667 : 16'b0000000001111111;
															assign node21667 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node21670 = (inp[9]) ? node21676 : node21671;
														assign node21671 = (inp[1]) ? node21673 : 16'b0000000000111111;
															assign node21673 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node21676 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node21679 = (inp[11]) ? node21697 : node21680;
												assign node21680 = (inp[9]) ? node21688 : node21681;
													assign node21681 = (inp[15]) ? node21685 : node21682;
														assign node21682 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node21685 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node21688 = (inp[1]) ? node21692 : node21689;
														assign node21689 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node21692 = (inp[2]) ? 16'b0000000000011111 : node21693;
															assign node21693 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node21697 = (inp[13]) ? node21699 : 16'b0000000000111111;
													assign node21699 = (inp[2]) ? node21703 : node21700;
														assign node21700 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node21703 = (inp[15]) ? 16'b0000000000001111 : node21704;
															assign node21704 = (inp[9]) ? node21706 : 16'b0000000000011111;
																assign node21706 = (inp[1]) ? 16'b0000000000001111 : 16'b0000000000011111;
								assign node21710 = (inp[1]) ? node21822 : node21711;
									assign node21711 = (inp[5]) ? node21753 : node21712;
										assign node21712 = (inp[11]) ? node21736 : node21713;
											assign node21713 = (inp[2]) ? node21725 : node21714;
												assign node21714 = (inp[15]) ? node21716 : 16'b0000000111111111;
													assign node21716 = (inp[3]) ? 16'b0000000011111111 : node21717;
														assign node21717 = (inp[13]) ? node21719 : 16'b0000000111111111;
															assign node21719 = (inp[10]) ? 16'b0000000011111111 : node21720;
																assign node21720 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node21725 = (inp[10]) ? node21729 : node21726;
													assign node21726 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node21729 = (inp[3]) ? node21733 : node21730;
														assign node21730 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node21733 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node21736 = (inp[9]) ? node21738 : 16'b0000000011111111;
												assign node21738 = (inp[2]) ? node21746 : node21739;
													assign node21739 = (inp[3]) ? node21743 : node21740;
														assign node21740 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node21743 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node21746 = (inp[13]) ? node21750 : node21747;
														assign node21747 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node21750 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node21753 = (inp[13]) ? node21793 : node21754;
											assign node21754 = (inp[10]) ? node21776 : node21755;
												assign node21755 = (inp[11]) ? node21767 : node21756;
													assign node21756 = (inp[3]) ? node21764 : node21757;
														assign node21757 = (inp[2]) ? 16'b0000000001111111 : node21758;
															assign node21758 = (inp[15]) ? node21760 : 16'b0000000111111111;
																assign node21760 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node21764 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node21767 = (inp[3]) ? node21771 : node21768;
														assign node21768 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node21771 = (inp[2]) ? node21773 : 16'b0000000001111111;
															assign node21773 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node21776 = (inp[9]) ? node21778 : 16'b0000000001111111;
													assign node21778 = (inp[11]) ? node21788 : node21779;
														assign node21779 = (inp[3]) ? node21783 : node21780;
															assign node21780 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
															assign node21783 = (inp[15]) ? 16'b0000000000111111 : node21784;
																assign node21784 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node21788 = (inp[2]) ? node21790 : 16'b0000000000111111;
															assign node21790 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node21793 = (inp[3]) ? node21803 : node21794;
												assign node21794 = (inp[10]) ? 16'b0000000000111111 : node21795;
													assign node21795 = (inp[2]) ? node21799 : node21796;
														assign node21796 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node21799 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node21803 = (inp[15]) ? node21811 : node21804;
													assign node21804 = (inp[10]) ? node21808 : node21805;
														assign node21805 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node21808 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node21811 = (inp[10]) ? node21817 : node21812;
														assign node21812 = (inp[11]) ? node21814 : 16'b0000000000011111;
															assign node21814 = (inp[2]) ? 16'b0000000000001111 : 16'b0000000000011111;
														assign node21817 = (inp[11]) ? 16'b0000000000001111 : node21818;
															assign node21818 = (inp[2]) ? 16'b0000000000001111 : 16'b0000000000011111;
									assign node21822 = (inp[3]) ? node21872 : node21823;
										assign node21823 = (inp[9]) ? node21855 : node21824;
											assign node21824 = (inp[11]) ? node21840 : node21825;
												assign node21825 = (inp[5]) ? node21835 : node21826;
													assign node21826 = (inp[2]) ? node21828 : 16'b0000000111111111;
														assign node21828 = (inp[13]) ? 16'b0000000001111111 : node21829;
															assign node21829 = (inp[10]) ? 16'b0000000011111111 : node21830;
																assign node21830 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node21835 = (inp[13]) ? node21837 : 16'b0000000001111111;
														assign node21837 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node21840 = (inp[13]) ? node21846 : node21841;
													assign node21841 = (inp[2]) ? node21843 : 16'b0000000011111111;
														assign node21843 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node21846 = (inp[15]) ? node21850 : node21847;
														assign node21847 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node21850 = (inp[2]) ? 16'b0000000000011111 : node21851;
															assign node21851 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node21855 = (inp[2]) ? 16'b0000000000111111 : node21856;
												assign node21856 = (inp[11]) ? node21866 : node21857;
													assign node21857 = (inp[13]) ? node21859 : 16'b0000000001111111;
														assign node21859 = (inp[10]) ? node21863 : node21860;
															assign node21860 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
															assign node21863 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node21866 = (inp[10]) ? 16'b0000000000011111 : node21867;
														assign node21867 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node21872 = (inp[11]) ? node21888 : node21873;
											assign node21873 = (inp[9]) ? node21881 : node21874;
												assign node21874 = (inp[10]) ? 16'b0000000000111111 : node21875;
													assign node21875 = (inp[2]) ? node21877 : 16'b0000000001111111;
														assign node21877 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node21881 = (inp[10]) ? node21883 : 16'b0000000000111111;
													assign node21883 = (inp[15]) ? node21885 : 16'b0000000000011111;
														assign node21885 = (inp[2]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node21888 = (inp[2]) ? node21904 : node21889;
												assign node21889 = (inp[9]) ? node21895 : node21890;
													assign node21890 = (inp[15]) ? 16'b0000000000111111 : node21891;
														assign node21891 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node21895 = (inp[5]) ? node21901 : node21896;
														assign node21896 = (inp[10]) ? 16'b0000000000011111 : node21897;
															assign node21897 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node21901 = (inp[13]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node21904 = (inp[9]) ? node21910 : node21905;
													assign node21905 = (inp[13]) ? node21907 : 16'b0000000000011111;
														assign node21907 = (inp[5]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node21910 = (inp[15]) ? 16'b0000000000001111 : 16'b0000000000111111;
						assign node21913 = (inp[15]) ? node22347 : node21914;
							assign node21914 = (inp[13]) ? node22130 : node21915;
								assign node21915 = (inp[5]) ? node22019 : node21916;
									assign node21916 = (inp[11]) ? node21974 : node21917;
										assign node21917 = (inp[2]) ? node21943 : node21918;
											assign node21918 = (inp[3]) ? node21934 : node21919;
												assign node21919 = (inp[12]) ? node21927 : node21920;
													assign node21920 = (inp[6]) ? 16'b0000001111111111 : node21921;
														assign node21921 = (inp[1]) ? node21923 : 16'b0000111111111111;
															assign node21923 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node21927 = (inp[6]) ? node21929 : 16'b0000001111111111;
														assign node21929 = (inp[1]) ? node21931 : 16'b0000000111111111;
															assign node21931 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node21934 = (inp[1]) ? node21938 : node21935;
													assign node21935 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node21938 = (inp[10]) ? 16'b0000000011111111 : node21939;
														assign node21939 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node21943 = (inp[12]) ? node21967 : node21944;
												assign node21944 = (inp[1]) ? node21960 : node21945;
													assign node21945 = (inp[9]) ? node21949 : node21946;
														assign node21946 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node21949 = (inp[6]) ? node21955 : node21950;
															assign node21950 = (inp[3]) ? node21952 : 16'b0000000111111111;
																assign node21952 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
															assign node21955 = (inp[3]) ? 16'b0000000011111111 : node21956;
																assign node21956 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node21960 = (inp[3]) ? node21964 : node21961;
														assign node21961 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node21964 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node21967 = (inp[9]) ? 16'b0000000001111111 : node21968;
													assign node21968 = (inp[10]) ? node21970 : 16'b0000000111111111;
														assign node21970 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node21974 = (inp[1]) ? node22000 : node21975;
											assign node21975 = (inp[9]) ? node21993 : node21976;
												assign node21976 = (inp[6]) ? node21984 : node21977;
													assign node21977 = (inp[10]) ? node21981 : node21978;
														assign node21978 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node21981 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node21984 = (inp[12]) ? node21988 : node21985;
														assign node21985 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node21988 = (inp[2]) ? node21990 : 16'b0000000011111111;
															assign node21990 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node21993 = (inp[2]) ? 16'b0000000001111111 : node21994;
													assign node21994 = (inp[10]) ? node21996 : 16'b0000000011111111;
														assign node21996 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000001111111;
											assign node22000 = (inp[3]) ? node22014 : node22001;
												assign node22001 = (inp[2]) ? node22003 : 16'b0000000111111111;
													assign node22003 = (inp[9]) ? node22011 : node22004;
														assign node22004 = (inp[12]) ? 16'b0000000001111111 : node22005;
															assign node22005 = (inp[10]) ? node22007 : 16'b0000000011111111;
																assign node22007 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node22011 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node22014 = (inp[9]) ? node22016 : 16'b0000000001111111;
													assign node22016 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000001111111;
									assign node22019 = (inp[10]) ? node22075 : node22020;
										assign node22020 = (inp[2]) ? node22050 : node22021;
											assign node22021 = (inp[9]) ? node22039 : node22022;
												assign node22022 = (inp[3]) ? node22030 : node22023;
													assign node22023 = (inp[6]) ? 16'b0000000111111111 : node22024;
														assign node22024 = (inp[1]) ? node22026 : 16'b0000001111111111;
															assign node22026 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node22030 = (inp[12]) ? node22036 : node22031;
														assign node22031 = (inp[6]) ? node22033 : 16'b0000001111111111;
															assign node22033 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node22036 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node22039 = (inp[3]) ? node22047 : node22040;
													assign node22040 = (inp[6]) ? node22044 : node22041;
														assign node22041 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node22044 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node22047 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node22050 = (inp[3]) ? node22064 : node22051;
												assign node22051 = (inp[9]) ? node22057 : node22052;
													assign node22052 = (inp[6]) ? node22054 : 16'b0000000011111111;
														assign node22054 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000001111111;
													assign node22057 = (inp[12]) ? node22061 : node22058;
														assign node22058 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node22061 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000001111111;
												assign node22064 = (inp[6]) ? node22072 : node22065;
													assign node22065 = (inp[9]) ? node22069 : node22066;
														assign node22066 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node22069 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node22072 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node22075 = (inp[6]) ? node22107 : node22076;
											assign node22076 = (inp[12]) ? node22090 : node22077;
												assign node22077 = (inp[3]) ? node22085 : node22078;
													assign node22078 = (inp[1]) ? node22082 : node22079;
														assign node22079 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node22082 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node22085 = (inp[11]) ? node22087 : 16'b0000000011111111;
														assign node22087 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node22090 = (inp[1]) ? node22094 : node22091;
													assign node22091 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node22094 = (inp[9]) ? node22100 : node22095;
														assign node22095 = (inp[3]) ? 16'b0000000000111111 : node22096;
															assign node22096 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node22100 = (inp[11]) ? node22102 : 16'b0000000000111111;
															assign node22102 = (inp[2]) ? 16'b0000000000011111 : node22103;
																assign node22103 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node22107 = (inp[9]) ? node22111 : node22108;
												assign node22108 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node22111 = (inp[1]) ? node22125 : node22112;
													assign node22112 = (inp[12]) ? node22118 : node22113;
														assign node22113 = (inp[11]) ? 16'b0000000000111111 : node22114;
															assign node22114 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node22118 = (inp[2]) ? 16'b0000000000011111 : node22119;
															assign node22119 = (inp[11]) ? node22121 : 16'b0000000000111111;
																assign node22121 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node22125 = (inp[3]) ? node22127 : 16'b0000000000011111;
														assign node22127 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
								assign node22130 = (inp[1]) ? node22238 : node22131;
									assign node22131 = (inp[2]) ? node22197 : node22132;
										assign node22132 = (inp[11]) ? node22160 : node22133;
											assign node22133 = (inp[9]) ? node22147 : node22134;
												assign node22134 = (inp[3]) ? node22142 : node22135;
													assign node22135 = (inp[12]) ? node22137 : 16'b0000000111111111;
														assign node22137 = (inp[6]) ? 16'b0000000111111111 : node22138;
															assign node22138 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node22142 = (inp[10]) ? 16'b0000000001111111 : node22143;
														assign node22143 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node22147 = (inp[12]) ? node22153 : node22148;
													assign node22148 = (inp[10]) ? node22150 : 16'b0000000011111111;
														assign node22150 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node22153 = (inp[10]) ? node22157 : node22154;
														assign node22154 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node22157 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node22160 = (inp[6]) ? node22182 : node22161;
												assign node22161 = (inp[12]) ? node22171 : node22162;
													assign node22162 = (inp[5]) ? node22164 : 16'b0000000111111111;
														assign node22164 = (inp[10]) ? 16'b0000000001111111 : node22165;
															assign node22165 = (inp[9]) ? node22167 : 16'b0000000011111111;
																assign node22167 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node22171 = (inp[5]) ? node22177 : node22172;
														assign node22172 = (inp[3]) ? 16'b0000000001111111 : node22173;
															assign node22173 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node22177 = (inp[10]) ? node22179 : 16'b0000000001111111;
															assign node22179 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node22182 = (inp[3]) ? node22186 : node22183;
													assign node22183 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node22186 = (inp[5]) ? node22194 : node22187;
														assign node22187 = (inp[10]) ? 16'b0000000000011111 : node22188;
															assign node22188 = (inp[12]) ? node22190 : 16'b0000000001111111;
																assign node22190 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node22194 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node22197 = (inp[3]) ? node22225 : node22198;
											assign node22198 = (inp[12]) ? node22204 : node22199;
												assign node22199 = (inp[5]) ? node22201 : 16'b0000000011111111;
													assign node22201 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node22204 = (inp[10]) ? node22214 : node22205;
													assign node22205 = (inp[5]) ? node22209 : node22206;
														assign node22206 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node22209 = (inp[9]) ? 16'b0000000000111111 : node22210;
															assign node22210 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node22214 = (inp[5]) ? node22222 : node22215;
														assign node22215 = (inp[11]) ? 16'b0000000000111111 : node22216;
															assign node22216 = (inp[9]) ? node22218 : 16'b0000000001111111;
																assign node22218 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node22222 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node22225 = (inp[11]) ? node22229 : node22226;
												assign node22226 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node22229 = (inp[12]) ? 16'b0000000000001111 : node22230;
													assign node22230 = (inp[5]) ? node22232 : 16'b0000000001111111;
														assign node22232 = (inp[9]) ? 16'b0000000000011111 : node22233;
															assign node22233 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node22238 = (inp[10]) ? node22294 : node22239;
										assign node22239 = (inp[2]) ? node22271 : node22240;
											assign node22240 = (inp[9]) ? node22258 : node22241;
												assign node22241 = (inp[6]) ? node22251 : node22242;
													assign node22242 = (inp[5]) ? node22244 : 16'b0000000011111111;
														assign node22244 = (inp[12]) ? node22246 : 16'b0000000011111111;
															assign node22246 = (inp[11]) ? node22248 : 16'b0000000011111111;
																assign node22248 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node22251 = (inp[3]) ? node22255 : node22252;
														assign node22252 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node22255 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node22258 = (inp[3]) ? node22264 : node22259;
													assign node22259 = (inp[5]) ? node22261 : 16'b0000000001111111;
														assign node22261 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node22264 = (inp[12]) ? node22268 : node22265;
														assign node22265 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000011111111;
														assign node22268 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node22271 = (inp[12]) ? node22277 : node22272;
												assign node22272 = (inp[5]) ? 16'b0000000000111111 : node22273;
													assign node22273 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node22277 = (inp[9]) ? node22285 : node22278;
													assign node22278 = (inp[3]) ? node22280 : 16'b0000000001111111;
														assign node22280 = (inp[6]) ? node22282 : 16'b0000000000111111;
															assign node22282 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node22285 = (inp[6]) ? node22289 : node22286;
														assign node22286 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node22289 = (inp[11]) ? node22291 : 16'b0000000000011111;
															assign node22291 = (inp[3]) ? 16'b0000000000001111 : 16'b0000000000011111;
										assign node22294 = (inp[12]) ? node22316 : node22295;
											assign node22295 = (inp[6]) ? node22305 : node22296;
												assign node22296 = (inp[5]) ? node22300 : node22297;
													assign node22297 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000001111111;
													assign node22300 = (inp[11]) ? 16'b0000000000011111 : node22301;
														assign node22301 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000011111111;
												assign node22305 = (inp[2]) ? node22313 : node22306;
													assign node22306 = (inp[3]) ? node22308 : 16'b0000000000111111;
														assign node22308 = (inp[9]) ? 16'b0000000000011111 : node22309;
															assign node22309 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node22313 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000000001111;
											assign node22316 = (inp[9]) ? node22334 : node22317;
												assign node22317 = (inp[11]) ? node22327 : node22318;
													assign node22318 = (inp[3]) ? node22320 : 16'b0000000000111111;
														assign node22320 = (inp[5]) ? node22324 : node22321;
															assign node22321 = (inp[6]) ? 16'b0000000000011111 : 16'b0000000000111111;
															assign node22324 = (inp[6]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node22327 = (inp[6]) ? node22329 : 16'b0000000000011111;
														assign node22329 = (inp[3]) ? node22331 : 16'b0000000000011111;
															assign node22331 = (inp[5]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node22334 = (inp[3]) ? node22336 : 16'b0000000000011111;
													assign node22336 = (inp[11]) ? node22340 : node22337;
														assign node22337 = (inp[6]) ? 16'b0000000000011111 : 16'b0000000000001111;
														assign node22340 = (inp[6]) ? 16'b0000000000000111 : node22341;
															assign node22341 = (inp[5]) ? node22343 : 16'b0000000000001111;
																assign node22343 = (inp[2]) ? 16'b0000000000000111 : 16'b0000000000001111;
							assign node22347 = (inp[10]) ? node22535 : node22348;
								assign node22348 = (inp[11]) ? node22452 : node22349;
									assign node22349 = (inp[3]) ? node22411 : node22350;
										assign node22350 = (inp[1]) ? node22382 : node22351;
											assign node22351 = (inp[5]) ? node22371 : node22352;
												assign node22352 = (inp[9]) ? node22358 : node22353;
													assign node22353 = (inp[13]) ? 16'b0000000111111111 : node22354;
														assign node22354 = (inp[2]) ? 16'b0000001111111111 : 16'b0000000111111111;
													assign node22358 = (inp[13]) ? node22364 : node22359;
														assign node22359 = (inp[6]) ? node22361 : 16'b0000000111111111;
															assign node22361 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node22364 = (inp[2]) ? 16'b0000000001111111 : node22365;
															assign node22365 = (inp[6]) ? 16'b0000000011111111 : node22366;
																assign node22366 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node22371 = (inp[13]) ? node22377 : node22372;
													assign node22372 = (inp[12]) ? node22374 : 16'b0000000011111111;
														assign node22374 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node22377 = (inp[9]) ? 16'b0000000000111111 : node22378;
														assign node22378 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node22382 = (inp[9]) ? node22398 : node22383;
												assign node22383 = (inp[12]) ? node22389 : node22384;
													assign node22384 = (inp[13]) ? 16'b0000000011111111 : node22385;
														assign node22385 = (inp[2]) ? 16'b0000000111111111 : 16'b0000000011111111;
													assign node22389 = (inp[5]) ? node22393 : node22390;
														assign node22390 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node22393 = (inp[2]) ? 16'b0000000000111111 : node22394;
															assign node22394 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node22398 = (inp[13]) ? node22402 : node22399;
													assign node22399 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node22402 = (inp[5]) ? node22408 : node22403;
														assign node22403 = (inp[2]) ? 16'b0000000000111111 : node22404;
															assign node22404 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node22408 = (inp[6]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node22411 = (inp[9]) ? node22431 : node22412;
											assign node22412 = (inp[5]) ? node22426 : node22413;
												assign node22413 = (inp[13]) ? node22419 : node22414;
													assign node22414 = (inp[12]) ? node22416 : 16'b0000000011111111;
														assign node22416 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000001111111;
													assign node22419 = (inp[2]) ? 16'b0000000000111111 : node22420;
														assign node22420 = (inp[1]) ? 16'b0000000001111111 : node22421;
															assign node22421 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node22426 = (inp[1]) ? 16'b0000000000111111 : node22427;
													assign node22427 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node22431 = (inp[6]) ? node22445 : node22432;
												assign node22432 = (inp[2]) ? node22438 : node22433;
													assign node22433 = (inp[5]) ? 16'b0000000001111111 : node22434;
														assign node22434 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node22438 = (inp[5]) ? node22442 : node22439;
														assign node22439 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node22442 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node22445 = (inp[5]) ? node22447 : 16'b0000000000111111;
													assign node22447 = (inp[13]) ? 16'b0000000000001111 : node22448;
														assign node22448 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node22452 = (inp[13]) ? node22486 : node22453;
										assign node22453 = (inp[1]) ? node22467 : node22454;
											assign node22454 = (inp[12]) ? node22462 : node22455;
												assign node22455 = (inp[3]) ? node22457 : 16'b0000000011111111;
													assign node22457 = (inp[5]) ? 16'b0000000001111111 : node22458;
														assign node22458 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node22462 = (inp[5]) ? 16'b0000000000111111 : node22463;
													assign node22463 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node22467 = (inp[2]) ? node22483 : node22468;
												assign node22468 = (inp[9]) ? node22476 : node22469;
													assign node22469 = (inp[6]) ? node22471 : 16'b0000000001111111;
														assign node22471 = (inp[3]) ? 16'b0000000000111111 : node22472;
															assign node22472 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node22476 = (inp[3]) ? node22478 : 16'b0000000000111111;
														assign node22478 = (inp[5]) ? node22480 : 16'b0000000000111111;
															assign node22480 = (inp[6]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node22483 = (inp[3]) ? 16'b0000000000001111 : 16'b0000000000011111;
										assign node22486 = (inp[9]) ? node22508 : node22487;
											assign node22487 = (inp[12]) ? node22501 : node22488;
												assign node22488 = (inp[2]) ? node22490 : 16'b0000000011111111;
													assign node22490 = (inp[1]) ? node22496 : node22491;
														assign node22491 = (inp[6]) ? node22493 : 16'b0000000001111111;
															assign node22493 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node22496 = (inp[3]) ? 16'b0000000000011111 : node22497;
															assign node22497 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node22501 = (inp[6]) ? node22503 : 16'b0000000000001111;
													assign node22503 = (inp[3]) ? 16'b0000000000011111 : node22504;
														assign node22504 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node22508 = (inp[2]) ? node22520 : node22509;
												assign node22509 = (inp[6]) ? node22511 : 16'b0000000000111111;
													assign node22511 = (inp[12]) ? 16'b0000000000011111 : node22512;
														assign node22512 = (inp[1]) ? node22514 : 16'b0000000000111111;
															assign node22514 = (inp[3]) ? 16'b0000000000011111 : node22515;
																assign node22515 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node22520 = (inp[5]) ? node22526 : node22521;
													assign node22521 = (inp[12]) ? node22523 : 16'b0000000000011111;
														assign node22523 = (inp[6]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node22526 = (inp[12]) ? node22532 : node22527;
														assign node22527 = (inp[6]) ? 16'b0000000000001111 : node22528;
															assign node22528 = (inp[3]) ? 16'b0000000000001111 : 16'b0000000000011111;
														assign node22532 = (inp[1]) ? 16'b0000000000000011 : 16'b0000000000001111;
								assign node22535 = (inp[6]) ? node22633 : node22536;
									assign node22536 = (inp[2]) ? node22584 : node22537;
										assign node22537 = (inp[13]) ? node22567 : node22538;
											assign node22538 = (inp[1]) ? node22550 : node22539;
												assign node22539 = (inp[5]) ? node22543 : node22540;
													assign node22540 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node22543 = (inp[12]) ? 16'b0000000000111111 : node22544;
														assign node22544 = (inp[9]) ? 16'b0000000001111111 : node22545;
															assign node22545 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node22550 = (inp[12]) ? node22558 : node22551;
													assign node22551 = (inp[11]) ? node22553 : 16'b0000000011111111;
														assign node22553 = (inp[9]) ? node22555 : 16'b0000000001111111;
															assign node22555 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node22558 = (inp[11]) ? 16'b0000000000011111 : node22559;
														assign node22559 = (inp[9]) ? 16'b0000000000111111 : node22560;
															assign node22560 = (inp[5]) ? node22562 : 16'b0000000001111111;
																assign node22562 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node22567 = (inp[5]) ? node22575 : node22568;
												assign node22568 = (inp[1]) ? node22570 : 16'b0000000001111111;
													assign node22570 = (inp[12]) ? 16'b0000000000001111 : node22571;
														assign node22571 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node22575 = (inp[9]) ? node22579 : node22576;
													assign node22576 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000001111111;
													assign node22579 = (inp[3]) ? node22581 : 16'b0000000000011111;
														assign node22581 = (inp[12]) ? 16'b0000000000001111 : 16'b0000000000011111;
										assign node22584 = (inp[3]) ? node22610 : node22585;
											assign node22585 = (inp[11]) ? node22603 : node22586;
												assign node22586 = (inp[12]) ? node22594 : node22587;
													assign node22587 = (inp[5]) ? node22589 : 16'b0000000011111111;
														assign node22589 = (inp[13]) ? node22591 : 16'b0000000001111111;
															assign node22591 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node22594 = (inp[9]) ? node22600 : node22595;
														assign node22595 = (inp[1]) ? 16'b0000000000111111 : node22596;
															assign node22596 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node22600 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node22603 = (inp[1]) ? node22605 : 16'b0000000000111111;
													assign node22605 = (inp[12]) ? 16'b0000000000011111 : node22606;
														assign node22606 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node22610 = (inp[5]) ? node22618 : node22611;
												assign node22611 = (inp[12]) ? node22613 : 16'b0000000000111111;
													assign node22613 = (inp[1]) ? 16'b0000000000001111 : node22614;
														assign node22614 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node22618 = (inp[9]) ? node22624 : node22619;
													assign node22619 = (inp[1]) ? node22621 : 16'b0000000000111111;
														assign node22621 = (inp[13]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node22624 = (inp[13]) ? node22630 : node22625;
														assign node22625 = (inp[12]) ? 16'b0000000000001111 : node22626;
															assign node22626 = (inp[1]) ? 16'b0000000000001111 : 16'b0000000000011111;
														assign node22630 = (inp[12]) ? 16'b0000000000000111 : 16'b0000000000001111;
									assign node22633 = (inp[12]) ? node22685 : node22634;
										assign node22634 = (inp[2]) ? node22656 : node22635;
											assign node22635 = (inp[3]) ? node22647 : node22636;
												assign node22636 = (inp[5]) ? node22644 : node22637;
													assign node22637 = (inp[1]) ? node22641 : node22638;
														assign node22638 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node22641 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node22644 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node22647 = (inp[11]) ? node22649 : 16'b0000000000111111;
													assign node22649 = (inp[5]) ? 16'b0000000000011111 : node22650;
														assign node22650 = (inp[9]) ? node22652 : 16'b0000000000111111;
															assign node22652 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node22656 = (inp[5]) ? node22672 : node22657;
												assign node22657 = (inp[13]) ? node22665 : node22658;
													assign node22658 = (inp[11]) ? node22660 : 16'b0000000000011111;
														assign node22660 = (inp[3]) ? 16'b0000000000111111 : node22661;
															assign node22661 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node22665 = (inp[3]) ? 16'b0000000000011111 : node22666;
														assign node22666 = (inp[11]) ? node22668 : 16'b0000000000011111;
															assign node22668 = (inp[1]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node22672 = (inp[13]) ? node22676 : node22673;
													assign node22673 = (inp[1]) ? 16'b0000000000000111 : 16'b0000000000011111;
													assign node22676 = (inp[11]) ? 16'b0000000000001111 : node22677;
														assign node22677 = (inp[9]) ? 16'b0000000000001111 : node22678;
															assign node22678 = (inp[1]) ? node22680 : 16'b0000000000011111;
																assign node22680 = (inp[3]) ? 16'b0000000000001111 : 16'b0000000000011111;
										assign node22685 = (inp[2]) ? node22711 : node22686;
											assign node22686 = (inp[13]) ? node22704 : node22687;
												assign node22687 = (inp[3]) ? node22695 : node22688;
													assign node22688 = (inp[11]) ? 16'b0000000000011111 : node22689;
														assign node22689 = (inp[1]) ? node22691 : 16'b0000000000111111;
															assign node22691 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node22695 = (inp[11]) ? node22697 : 16'b0000000000011111;
														assign node22697 = (inp[5]) ? 16'b0000000000001111 : node22698;
															assign node22698 = (inp[1]) ? node22700 : 16'b0000000000011111;
																assign node22700 = (inp[9]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node22704 = (inp[5]) ? node22706 : 16'b0000000000011111;
													assign node22706 = (inp[11]) ? 16'b0000000000001111 : node22707;
														assign node22707 = (inp[9]) ? 16'b0000000000000111 : 16'b0000000000001111;
											assign node22711 = (inp[11]) ? node22729 : node22712;
												assign node22712 = (inp[9]) ? node22720 : node22713;
													assign node22713 = (inp[1]) ? node22717 : node22714;
														assign node22714 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node22717 = (inp[5]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node22720 = (inp[5]) ? node22722 : 16'b0000000000001111;
														assign node22722 = (inp[1]) ? node22724 : 16'b0000000000001111;
															assign node22724 = (inp[3]) ? 16'b0000000000000111 : node22725;
																assign node22725 = (inp[13]) ? 16'b0000000000000111 : 16'b0000000000001111;
												assign node22729 = (inp[5]) ? node22731 : 16'b0000000000001111;
													assign node22731 = (inp[9]) ? 16'b0000000000000011 : node22732;
														assign node22732 = (inp[1]) ? node22734 : 16'b0000000000000111;
															assign node22734 = (inp[13]) ? 16'b0000000000000011 : 16'b0000000000000111;
					assign node22738 = (inp[1]) ? node23494 : node22739;
						assign node22739 = (inp[10]) ? node23081 : node22740;
							assign node22740 = (inp[14]) ? node22918 : node22741;
								assign node22741 = (inp[5]) ? node22837 : node22742;
									assign node22742 = (inp[9]) ? node22798 : node22743;
										assign node22743 = (inp[12]) ? node22777 : node22744;
											assign node22744 = (inp[15]) ? node22760 : node22745;
												assign node22745 = (inp[11]) ? node22753 : node22746;
													assign node22746 = (inp[13]) ? node22750 : node22747;
														assign node22747 = (inp[6]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node22750 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node22753 = (inp[3]) ? node22757 : node22754;
														assign node22754 = (inp[6]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node22757 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node22760 = (inp[2]) ? node22772 : node22761;
													assign node22761 = (inp[3]) ? node22767 : node22762;
														assign node22762 = (inp[13]) ? 16'b0000000111111111 : node22763;
															assign node22763 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node22767 = (inp[13]) ? node22769 : 16'b0000000111111111;
															assign node22769 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node22772 = (inp[6]) ? node22774 : 16'b0000000111111111;
														assign node22774 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node22777 = (inp[3]) ? node22789 : node22778;
												assign node22778 = (inp[6]) ? node22784 : node22779;
													assign node22779 = (inp[11]) ? 16'b0000000111111111 : node22780;
														assign node22780 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node22784 = (inp[15]) ? 16'b0000000001111111 : node22785;
														assign node22785 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node22789 = (inp[11]) ? node22793 : node22790;
													assign node22790 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node22793 = (inp[6]) ? node22795 : 16'b0000000001111111;
														assign node22795 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node22798 = (inp[6]) ? node22812 : node22799;
											assign node22799 = (inp[13]) ? node22807 : node22800;
												assign node22800 = (inp[12]) ? node22804 : node22801;
													assign node22801 = (inp[15]) ? 16'b0000000011111111 : 16'b0000001111111111;
													assign node22804 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node22807 = (inp[2]) ? node22809 : 16'b0000000011111111;
													assign node22809 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node22812 = (inp[3]) ? node22824 : node22813;
												assign node22813 = (inp[11]) ? node22819 : node22814;
													assign node22814 = (inp[2]) ? node22816 : 16'b0000000011111111;
														assign node22816 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node22819 = (inp[2]) ? 16'b0000000000011111 : node22820;
														assign node22820 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node22824 = (inp[15]) ? node22832 : node22825;
													assign node22825 = (inp[2]) ? node22827 : 16'b0000000001111111;
														assign node22827 = (inp[12]) ? node22829 : 16'b0000000001111111;
															assign node22829 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node22832 = (inp[2]) ? 16'b0000000000011111 : node22833;
														assign node22833 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node22837 = (inp[3]) ? node22875 : node22838;
										assign node22838 = (inp[12]) ? node22856 : node22839;
											assign node22839 = (inp[6]) ? node22853 : node22840;
												assign node22840 = (inp[15]) ? node22850 : node22841;
													assign node22841 = (inp[13]) ? node22843 : 16'b0000001111111111;
														assign node22843 = (inp[2]) ? 16'b0000000011111111 : node22844;
															assign node22844 = (inp[11]) ? node22846 : 16'b0000000111111111;
																assign node22846 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node22850 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node22853 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node22856 = (inp[6]) ? node22868 : node22857;
												assign node22857 = (inp[15]) ? node22863 : node22858;
													assign node22858 = (inp[9]) ? 16'b0000000001111111 : node22859;
														assign node22859 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node22863 = (inp[9]) ? node22865 : 16'b0000000001111111;
														assign node22865 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node22868 = (inp[15]) ? 16'b0000000000111111 : node22869;
													assign node22869 = (inp[13]) ? node22871 : 16'b0000000001111111;
														assign node22871 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node22875 = (inp[2]) ? node22893 : node22876;
											assign node22876 = (inp[13]) ? node22884 : node22877;
												assign node22877 = (inp[9]) ? 16'b0000000001111111 : node22878;
													assign node22878 = (inp[12]) ? node22880 : 16'b0000000011111111;
														assign node22880 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node22884 = (inp[6]) ? 16'b0000000000111111 : node22885;
													assign node22885 = (inp[11]) ? node22889 : node22886;
														assign node22886 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node22889 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node22893 = (inp[13]) ? node22905 : node22894;
												assign node22894 = (inp[9]) ? node22900 : node22895;
													assign node22895 = (inp[15]) ? node22897 : 16'b0000000001111111;
														assign node22897 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node22900 = (inp[6]) ? 16'b0000000000111111 : node22901;
														assign node22901 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node22905 = (inp[12]) ? node22911 : node22906;
													assign node22906 = (inp[11]) ? 16'b0000000000111111 : node22907;
														assign node22907 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node22911 = (inp[9]) ? node22913 : 16'b0000000000001111;
														assign node22913 = (inp[15]) ? 16'b0000000000011111 : node22914;
															assign node22914 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
								assign node22918 = (inp[6]) ? node23004 : node22919;
									assign node22919 = (inp[5]) ? node22961 : node22920;
										assign node22920 = (inp[9]) ? node22944 : node22921;
											assign node22921 = (inp[3]) ? node22935 : node22922;
												assign node22922 = (inp[2]) ? node22926 : node22923;
													assign node22923 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node22926 = (inp[13]) ? node22930 : node22927;
														assign node22927 = (inp[15]) ? 16'b0000000011111111 : 16'b0000001111111111;
														assign node22930 = (inp[11]) ? node22932 : 16'b0000000011111111;
															assign node22932 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node22935 = (inp[12]) ? node22941 : node22936;
													assign node22936 = (inp[2]) ? 16'b0000000011111111 : node22937;
														assign node22937 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node22941 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node22944 = (inp[11]) ? node22952 : node22945;
												assign node22945 = (inp[13]) ? 16'b0000000001111111 : node22946;
													assign node22946 = (inp[15]) ? node22948 : 16'b0000000011111111;
														assign node22948 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node22952 = (inp[2]) ? 16'b0000000000111111 : node22953;
													assign node22953 = (inp[13]) ? node22955 : 16'b0000000011111111;
														assign node22955 = (inp[15]) ? node22957 : 16'b0000000001111111;
															assign node22957 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000001111111;
										assign node22961 = (inp[2]) ? node22981 : node22962;
											assign node22962 = (inp[13]) ? node22966 : node22963;
												assign node22963 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node22966 = (inp[11]) ? node22976 : node22967;
													assign node22967 = (inp[9]) ? node22969 : 16'b0000000011111111;
														assign node22969 = (inp[15]) ? node22971 : 16'b0000000001111111;
															assign node22971 = (inp[3]) ? 16'b0000000000111111 : node22972;
																assign node22972 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node22976 = (inp[12]) ? node22978 : 16'b0000000000111111;
														assign node22978 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node22981 = (inp[15]) ? node22995 : node22982;
												assign node22982 = (inp[12]) ? node22988 : node22983;
													assign node22983 = (inp[9]) ? node22985 : 16'b0000000001111111;
														assign node22985 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node22988 = (inp[9]) ? 16'b0000000001111111 : node22989;
														assign node22989 = (inp[13]) ? node22991 : 16'b0000000000111111;
															assign node22991 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node22995 = (inp[11]) ? 16'b0000000000011111 : node22996;
													assign node22996 = (inp[3]) ? node22998 : 16'b0000000000111111;
														assign node22998 = (inp[13]) ? 16'b0000000000011111 : node22999;
															assign node22999 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node23004 = (inp[11]) ? node23050 : node23005;
										assign node23005 = (inp[15]) ? node23027 : node23006;
											assign node23006 = (inp[3]) ? node23020 : node23007;
												assign node23007 = (inp[9]) ? node23011 : node23008;
													assign node23008 = (inp[12]) ? 16'b0000000111111111 : 16'b0000000011111111;
													assign node23011 = (inp[12]) ? 16'b0000000001111111 : node23012;
														assign node23012 = (inp[13]) ? node23014 : 16'b0000000011111111;
															assign node23014 = (inp[2]) ? 16'b0000000001111111 : node23015;
																assign node23015 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node23020 = (inp[12]) ? node23024 : node23021;
													assign node23021 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node23024 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node23027 = (inp[13]) ? node23041 : node23028;
												assign node23028 = (inp[3]) ? node23034 : node23029;
													assign node23029 = (inp[2]) ? node23031 : 16'b0000000011111111;
														assign node23031 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node23034 = (inp[9]) ? node23038 : node23035;
														assign node23035 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node23038 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node23041 = (inp[3]) ? 16'b0000000000011111 : node23042;
													assign node23042 = (inp[2]) ? node23044 : 16'b0000000000111111;
														assign node23044 = (inp[9]) ? 16'b0000000000011111 : node23045;
															assign node23045 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node23050 = (inp[3]) ? node23056 : node23051;
											assign node23051 = (inp[5]) ? node23053 : 16'b0000000000111111;
												assign node23053 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000001111111;
											assign node23056 = (inp[9]) ? node23068 : node23057;
												assign node23057 = (inp[2]) ? node23065 : node23058;
													assign node23058 = (inp[13]) ? node23060 : 16'b0000000000111111;
														assign node23060 = (inp[12]) ? node23062 : 16'b0000000000111111;
															assign node23062 = (inp[15]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node23065 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000001111;
												assign node23068 = (inp[12]) ? node23074 : node23069;
													assign node23069 = (inp[13]) ? 16'b0000000000011111 : node23070;
														assign node23070 = (inp[2]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node23074 = (inp[15]) ? 16'b0000000000000111 : node23075;
														assign node23075 = (inp[5]) ? node23077 : 16'b0000000000011111;
															assign node23077 = (inp[2]) ? 16'b0000000000000111 : 16'b0000000000001111;
							assign node23081 = (inp[13]) ? node23277 : node23082;
								assign node23082 = (inp[3]) ? node23168 : node23083;
									assign node23083 = (inp[5]) ? node23125 : node23084;
										assign node23084 = (inp[15]) ? node23106 : node23085;
											assign node23085 = (inp[2]) ? node23099 : node23086;
												assign node23086 = (inp[9]) ? node23092 : node23087;
													assign node23087 = (inp[11]) ? 16'b0000000111111111 : node23088;
														assign node23088 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node23092 = (inp[14]) ? 16'b0000000001111111 : node23093;
														assign node23093 = (inp[11]) ? node23095 : 16'b0000000111111111;
															assign node23095 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node23099 = (inp[14]) ? 16'b0000000001111111 : node23100;
													assign node23100 = (inp[11]) ? 16'b0000000011111111 : node23101;
														assign node23101 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node23106 = (inp[6]) ? node23116 : node23107;
												assign node23107 = (inp[12]) ? node23113 : node23108;
													assign node23108 = (inp[2]) ? 16'b0000000011111111 : node23109;
														assign node23109 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node23113 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000011111111;
												assign node23116 = (inp[11]) ? node23118 : 16'b0000000001111111;
													assign node23118 = (inp[12]) ? node23122 : node23119;
														assign node23119 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node23122 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node23125 = (inp[9]) ? node23141 : node23126;
											assign node23126 = (inp[12]) ? node23138 : node23127;
												assign node23127 = (inp[15]) ? 16'b0000000001111111 : node23128;
													assign node23128 = (inp[2]) ? node23132 : node23129;
														assign node23129 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node23132 = (inp[14]) ? node23134 : 16'b0000000011111111;
															assign node23134 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node23138 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node23141 = (inp[12]) ? node23155 : node23142;
												assign node23142 = (inp[2]) ? node23150 : node23143;
													assign node23143 = (inp[15]) ? node23147 : node23144;
														assign node23144 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node23147 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node23150 = (inp[6]) ? 16'b0000000000111111 : node23151;
														assign node23151 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node23155 = (inp[11]) ? node23163 : node23156;
													assign node23156 = (inp[15]) ? 16'b0000000000111111 : node23157;
														assign node23157 = (inp[14]) ? node23159 : 16'b0000000000111111;
															assign node23159 = (inp[6]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node23163 = (inp[15]) ? 16'b0000000000011111 : node23164;
														assign node23164 = (inp[2]) ? 16'b0000000000001111 : 16'b0000000000011111;
									assign node23168 = (inp[14]) ? node23222 : node23169;
										assign node23169 = (inp[12]) ? node23193 : node23170;
											assign node23170 = (inp[2]) ? node23184 : node23171;
												assign node23171 = (inp[5]) ? node23177 : node23172;
													assign node23172 = (inp[6]) ? node23174 : 16'b0000000011111111;
														assign node23174 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node23177 = (inp[15]) ? 16'b0000000001111111 : node23178;
														assign node23178 = (inp[11]) ? node23180 : 16'b0000000111111111;
															assign node23180 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node23184 = (inp[6]) ? node23190 : node23185;
													assign node23185 = (inp[9]) ? node23187 : 16'b0000000001111111;
														assign node23187 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node23190 = (inp[5]) ? 16'b0000000000001111 : 16'b0000000000111111;
											assign node23193 = (inp[11]) ? node23209 : node23194;
												assign node23194 = (inp[5]) ? node23202 : node23195;
													assign node23195 = (inp[2]) ? node23199 : node23196;
														assign node23196 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node23199 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node23202 = (inp[6]) ? 16'b0000000000111111 : node23203;
														assign node23203 = (inp[9]) ? 16'b0000000000111111 : node23204;
															assign node23204 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node23209 = (inp[15]) ? node23217 : node23210;
													assign node23210 = (inp[2]) ? node23212 : 16'b0000000000111111;
														assign node23212 = (inp[5]) ? node23214 : 16'b0000000000111111;
															assign node23214 = (inp[6]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node23217 = (inp[6]) ? 16'b0000000000011111 : node23218;
														assign node23218 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000001111111;
										assign node23222 = (inp[15]) ? node23252 : node23223;
											assign node23223 = (inp[5]) ? node23239 : node23224;
												assign node23224 = (inp[9]) ? node23230 : node23225;
													assign node23225 = (inp[11]) ? node23227 : 16'b0000000001111111;
														assign node23227 = (inp[6]) ? 16'b0000000000011111 : 16'b0000000001111111;
													assign node23230 = (inp[2]) ? node23236 : node23231;
														assign node23231 = (inp[12]) ? node23233 : 16'b0000000001111111;
															assign node23233 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node23236 = (inp[6]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node23239 = (inp[6]) ? node23245 : node23240;
													assign node23240 = (inp[2]) ? 16'b0000000000011111 : node23241;
														assign node23241 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node23245 = (inp[2]) ? 16'b0000000000001111 : node23246;
														assign node23246 = (inp[12]) ? node23248 : 16'b0000000000111111;
															assign node23248 = (inp[11]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node23252 = (inp[12]) ? node23266 : node23253;
												assign node23253 = (inp[11]) ? node23261 : node23254;
													assign node23254 = (inp[9]) ? 16'b0000000000011111 : node23255;
														assign node23255 = (inp[6]) ? 16'b0000000000111111 : node23256;
															assign node23256 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node23261 = (inp[5]) ? 16'b0000000000011111 : node23262;
														assign node23262 = (inp[6]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node23266 = (inp[9]) ? node23272 : node23267;
													assign node23267 = (inp[6]) ? 16'b0000000000011111 : node23268;
														assign node23268 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node23272 = (inp[11]) ? node23274 : 16'b0000000000001111;
														assign node23274 = (inp[5]) ? 16'b0000000000000111 : 16'b0000000000001111;
								assign node23277 = (inp[11]) ? node23397 : node23278;
									assign node23278 = (inp[6]) ? node23332 : node23279;
										assign node23279 = (inp[5]) ? node23297 : node23280;
											assign node23280 = (inp[9]) ? node23288 : node23281;
												assign node23281 = (inp[15]) ? 16'b0000000001111111 : node23282;
													assign node23282 = (inp[3]) ? node23284 : 16'b0000000011111111;
														assign node23284 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node23288 = (inp[12]) ? node23294 : node23289;
													assign node23289 = (inp[3]) ? node23291 : 16'b0000000001111111;
														assign node23291 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node23294 = (inp[2]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node23297 = (inp[14]) ? node23319 : node23298;
												assign node23298 = (inp[12]) ? node23312 : node23299;
													assign node23299 = (inp[3]) ? node23305 : node23300;
														assign node23300 = (inp[9]) ? node23302 : 16'b0000000011111111;
															assign node23302 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node23305 = (inp[15]) ? 16'b0000000000111111 : node23306;
															assign node23306 = (inp[2]) ? 16'b0000000001111111 : node23307;
																assign node23307 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node23312 = (inp[15]) ? node23314 : 16'b0000000000111111;
														assign node23314 = (inp[3]) ? node23316 : 16'b0000000000111111;
															assign node23316 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node23319 = (inp[9]) ? node23321 : 16'b0000000000111111;
													assign node23321 = (inp[15]) ? node23327 : node23322;
														assign node23322 = (inp[3]) ? node23324 : 16'b0000000000111111;
															assign node23324 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node23327 = (inp[2]) ? node23329 : 16'b0000000000011111;
															assign node23329 = (inp[3]) ? 16'b0000000000001111 : 16'b0000000000011111;
										assign node23332 = (inp[3]) ? node23368 : node23333;
											assign node23333 = (inp[15]) ? node23353 : node23334;
												assign node23334 = (inp[2]) ? node23346 : node23335;
													assign node23335 = (inp[12]) ? node23339 : node23336;
														assign node23336 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node23339 = (inp[9]) ? 16'b0000000000111111 : node23340;
															assign node23340 = (inp[5]) ? node23342 : 16'b0000000001111111;
																assign node23342 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node23346 = (inp[5]) ? node23350 : node23347;
														assign node23347 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node23350 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node23353 = (inp[2]) ? node23363 : node23354;
													assign node23354 = (inp[14]) ? node23356 : 16'b0000000000111111;
														assign node23356 = (inp[12]) ? 16'b0000000000011111 : node23357;
															assign node23357 = (inp[5]) ? node23359 : 16'b0000000001111111;
																assign node23359 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node23363 = (inp[9]) ? 16'b0000000000011111 : node23364;
														assign node23364 = (inp[12]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node23368 = (inp[9]) ? node23376 : node23369;
												assign node23369 = (inp[12]) ? 16'b0000000000011111 : node23370;
													assign node23370 = (inp[14]) ? node23372 : 16'b0000000000111111;
														assign node23372 = (inp[2]) ? 16'b0000000000001111 : 16'b0000000000111111;
												assign node23376 = (inp[5]) ? node23384 : node23377;
													assign node23377 = (inp[2]) ? 16'b0000000000001111 : node23378;
														assign node23378 = (inp[12]) ? 16'b0000000000011111 : node23379;
															assign node23379 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node23384 = (inp[12]) ? node23388 : node23385;
														assign node23385 = (inp[14]) ? 16'b0000000000001111 : 16'b0000000000011111;
														assign node23388 = (inp[2]) ? node23392 : node23389;
															assign node23389 = (inp[14]) ? 16'b0000000000000111 : 16'b0000000000001111;
															assign node23392 = (inp[15]) ? node23394 : 16'b0000000000000111;
																assign node23394 = (inp[14]) ? 16'b0000000000000011 : 16'b0000000000000111;
									assign node23397 = (inp[9]) ? node23455 : node23398;
										assign node23398 = (inp[12]) ? node23424 : node23399;
											assign node23399 = (inp[5]) ? node23411 : node23400;
												assign node23400 = (inp[3]) ? node23404 : node23401;
													assign node23401 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node23404 = (inp[2]) ? node23406 : 16'b0000000000111111;
														assign node23406 = (inp[14]) ? node23408 : 16'b0000000000111111;
															assign node23408 = (inp[6]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node23411 = (inp[3]) ? node23419 : node23412;
													assign node23412 = (inp[14]) ? node23414 : 16'b0000000000111111;
														assign node23414 = (inp[6]) ? 16'b0000000000011111 : node23415;
															assign node23415 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node23419 = (inp[6]) ? node23421 : 16'b0000000000011111;
														assign node23421 = (inp[14]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node23424 = (inp[2]) ? node23436 : node23425;
												assign node23425 = (inp[15]) ? node23431 : node23426;
													assign node23426 = (inp[6]) ? node23428 : 16'b0000000001111111;
														assign node23428 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node23431 = (inp[5]) ? 16'b0000000000001111 : node23432;
														assign node23432 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node23436 = (inp[6]) ? node23448 : node23437;
													assign node23437 = (inp[15]) ? node23441 : node23438;
														assign node23438 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node23441 = (inp[3]) ? 16'b0000000000001111 : node23442;
															assign node23442 = (inp[14]) ? node23444 : 16'b0000000000011111;
																assign node23444 = (inp[5]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node23448 = (inp[15]) ? node23450 : 16'b0000000000001111;
														assign node23450 = (inp[5]) ? node23452 : 16'b0000000000001111;
															assign node23452 = (inp[14]) ? 16'b0000000000000111 : 16'b0000000000001111;
										assign node23455 = (inp[3]) ? node23473 : node23456;
											assign node23456 = (inp[14]) ? node23466 : node23457;
												assign node23457 = (inp[12]) ? node23461 : node23458;
													assign node23458 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node23461 = (inp[15]) ? 16'b0000000000001111 : node23462;
														assign node23462 = (inp[6]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node23466 = (inp[5]) ? node23468 : 16'b0000000000011111;
													assign node23468 = (inp[12]) ? 16'b0000000000001111 : node23469;
														assign node23469 = (inp[15]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node23473 = (inp[12]) ? node23481 : node23474;
												assign node23474 = (inp[14]) ? node23478 : node23475;
													assign node23475 = (inp[5]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node23478 = (inp[6]) ? 16'b0000000000000111 : 16'b0000000000001111;
												assign node23481 = (inp[15]) ? node23485 : node23482;
													assign node23482 = (inp[6]) ? 16'b0000000000001111 : 16'b0000000000000111;
													assign node23485 = (inp[2]) ? node23487 : 16'b0000000000000111;
														assign node23487 = (inp[6]) ? node23489 : 16'b0000000000000111;
															assign node23489 = (inp[5]) ? 16'b0000000000000011 : node23490;
																assign node23490 = (inp[14]) ? 16'b0000000000000011 : 16'b0000000000000111;
						assign node23494 = (inp[2]) ? node23876 : node23495;
							assign node23495 = (inp[15]) ? node23669 : node23496;
								assign node23496 = (inp[14]) ? node23572 : node23497;
									assign node23497 = (inp[11]) ? node23541 : node23498;
										assign node23498 = (inp[10]) ? node23514 : node23499;
											assign node23499 = (inp[3]) ? node23509 : node23500;
												assign node23500 = (inp[5]) ? node23504 : node23501;
													assign node23501 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node23504 = (inp[6]) ? 16'b0000000011111111 : node23505;
														assign node23505 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000111111111;
												assign node23509 = (inp[9]) ? node23511 : 16'b0000000011111111;
													assign node23511 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node23514 = (inp[13]) ? node23528 : node23515;
												assign node23515 = (inp[5]) ? node23523 : node23516;
													assign node23516 = (inp[12]) ? node23518 : 16'b0000000011111111;
														assign node23518 = (inp[6]) ? 16'b0000000001111111 : node23519;
															assign node23519 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node23523 = (inp[3]) ? 16'b0000000001111111 : node23524;
														assign node23524 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node23528 = (inp[12]) ? node23538 : node23529;
													assign node23529 = (inp[6]) ? node23533 : node23530;
														assign node23530 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node23533 = (inp[9]) ? node23535 : 16'b0000000001111111;
															assign node23535 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node23538 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node23541 = (inp[10]) ? node23555 : node23542;
											assign node23542 = (inp[6]) ? node23548 : node23543;
												assign node23543 = (inp[3]) ? node23545 : 16'b0000000111111111;
													assign node23545 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node23548 = (inp[9]) ? node23550 : 16'b0000000001111111;
													assign node23550 = (inp[3]) ? 16'b0000000000011111 : node23551;
														assign node23551 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node23555 = (inp[5]) ? node23565 : node23556;
												assign node23556 = (inp[12]) ? 16'b0000000000111111 : node23557;
													assign node23557 = (inp[13]) ? 16'b0000000000111111 : node23558;
														assign node23558 = (inp[9]) ? node23560 : 16'b0000000001111111;
															assign node23560 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node23565 = (inp[6]) ? node23567 : 16'b0000000001111111;
													assign node23567 = (inp[9]) ? 16'b0000000000001111 : node23568;
														assign node23568 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node23572 = (inp[12]) ? node23636 : node23573;
										assign node23573 = (inp[5]) ? node23607 : node23574;
											assign node23574 = (inp[11]) ? node23594 : node23575;
												assign node23575 = (inp[13]) ? node23581 : node23576;
													assign node23576 = (inp[10]) ? 16'b0000000011111111 : node23577;
														assign node23577 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node23581 = (inp[9]) ? node23591 : node23582;
														assign node23582 = (inp[6]) ? node23586 : node23583;
															assign node23583 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
															assign node23586 = (inp[10]) ? 16'b0000000001111111 : node23587;
																assign node23587 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node23591 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node23594 = (inp[13]) ? node23598 : node23595;
													assign node23595 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node23598 = (inp[6]) ? 16'b0000000000111111 : node23599;
														assign node23599 = (inp[10]) ? 16'b0000000000111111 : node23600;
															assign node23600 = (inp[3]) ? node23602 : 16'b0000000001111111;
																assign node23602 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node23607 = (inp[3]) ? node23623 : node23608;
												assign node23608 = (inp[13]) ? node23612 : node23609;
													assign node23609 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000111111111;
													assign node23612 = (inp[9]) ? node23620 : node23613;
														assign node23613 = (inp[11]) ? node23615 : 16'b0000000001111111;
															assign node23615 = (inp[10]) ? 16'b0000000000111111 : node23616;
																assign node23616 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node23620 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node23623 = (inp[6]) ? node23629 : node23624;
													assign node23624 = (inp[10]) ? node23626 : 16'b0000000001111111;
														assign node23626 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node23629 = (inp[13]) ? node23631 : 16'b0000000000011111;
														assign node23631 = (inp[11]) ? 16'b0000000000000111 : node23632;
															assign node23632 = (inp[9]) ? 16'b0000000000001111 : 16'b0000000000011111;
										assign node23636 = (inp[3]) ? node23652 : node23637;
											assign node23637 = (inp[13]) ? node23643 : node23638;
												assign node23638 = (inp[10]) ? 16'b0000000000111111 : node23639;
													assign node23639 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node23643 = (inp[6]) ? node23647 : node23644;
													assign node23644 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000000011111;
													assign node23647 = (inp[11]) ? node23649 : 16'b0000000000011111;
														assign node23649 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node23652 = (inp[6]) ? node23660 : node23653;
												assign node23653 = (inp[9]) ? 16'b0000000000011111 : node23654;
													assign node23654 = (inp[5]) ? 16'b0000000000011111 : node23655;
														assign node23655 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node23660 = (inp[11]) ? node23662 : 16'b0000000000011111;
													assign node23662 = (inp[9]) ? node23666 : node23663;
														assign node23663 = (inp[5]) ? 16'b0000000000001111 : 16'b0000000000011111;
														assign node23666 = (inp[5]) ? 16'b0000000000000111 : 16'b0000000000001111;
								assign node23669 = (inp[11]) ? node23767 : node23670;
									assign node23670 = (inp[6]) ? node23708 : node23671;
										assign node23671 = (inp[12]) ? node23693 : node23672;
											assign node23672 = (inp[3]) ? node23686 : node23673;
												assign node23673 = (inp[14]) ? node23681 : node23674;
													assign node23674 = (inp[9]) ? node23676 : 16'b0000000011111111;
														assign node23676 = (inp[13]) ? node23678 : 16'b0000000011111111;
															assign node23678 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node23681 = (inp[5]) ? node23683 : 16'b0000000001111111;
														assign node23683 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node23686 = (inp[14]) ? 16'b0000000000011111 : node23687;
													assign node23687 = (inp[10]) ? node23689 : 16'b0000000001111111;
														assign node23689 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node23693 = (inp[13]) ? node23701 : node23694;
												assign node23694 = (inp[5]) ? 16'b0000000000111111 : node23695;
													assign node23695 = (inp[10]) ? node23697 : 16'b0000000001111111;
														assign node23697 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node23701 = (inp[3]) ? 16'b0000000000011111 : node23702;
													assign node23702 = (inp[14]) ? node23704 : 16'b0000000001111111;
														assign node23704 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node23708 = (inp[9]) ? node23736 : node23709;
											assign node23709 = (inp[13]) ? node23725 : node23710;
												assign node23710 = (inp[3]) ? node23716 : node23711;
													assign node23711 = (inp[12]) ? 16'b0000000001111111 : node23712;
														assign node23712 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node23716 = (inp[5]) ? 16'b0000000000111111 : node23717;
														assign node23717 = (inp[12]) ? node23719 : 16'b0000000001111111;
															assign node23719 = (inp[10]) ? 16'b0000000000111111 : node23720;
																assign node23720 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node23725 = (inp[3]) ? node23731 : node23726;
													assign node23726 = (inp[5]) ? 16'b0000000000111111 : node23727;
														assign node23727 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node23731 = (inp[10]) ? node23733 : 16'b0000000000111111;
														assign node23733 = (inp[14]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node23736 = (inp[5]) ? node23756 : node23737;
												assign node23737 = (inp[10]) ? node23747 : node23738;
													assign node23738 = (inp[14]) ? node23744 : node23739;
														assign node23739 = (inp[3]) ? 16'b0000000000111111 : node23740;
															assign node23740 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node23744 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node23747 = (inp[3]) ? node23751 : node23748;
														assign node23748 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node23751 = (inp[14]) ? node23753 : 16'b0000000000011111;
															assign node23753 = (inp[12]) ? 16'b0000000000000111 : 16'b0000000000001111;
												assign node23756 = (inp[3]) ? 16'b0000000000001111 : node23757;
													assign node23757 = (inp[13]) ? node23761 : node23758;
														assign node23758 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node23761 = (inp[10]) ? 16'b0000000000001111 : node23762;
															assign node23762 = (inp[14]) ? 16'b0000000000001111 : 16'b0000000000011111;
									assign node23767 = (inp[3]) ? node23835 : node23768;
										assign node23768 = (inp[13]) ? node23792 : node23769;
											assign node23769 = (inp[6]) ? node23779 : node23770;
												assign node23770 = (inp[10]) ? 16'b0000000011111111 : node23771;
													assign node23771 = (inp[14]) ? node23773 : 16'b0000000001111111;
														assign node23773 = (inp[9]) ? 16'b0000000000111111 : node23774;
															assign node23774 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node23779 = (inp[12]) ? node23787 : node23780;
													assign node23780 = (inp[14]) ? node23784 : node23781;
														assign node23781 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node23784 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node23787 = (inp[14]) ? node23789 : 16'b0000000000011111;
														assign node23789 = (inp[5]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node23792 = (inp[5]) ? node23814 : node23793;
												assign node23793 = (inp[9]) ? node23803 : node23794;
													assign node23794 = (inp[6]) ? node23798 : node23795;
														assign node23795 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000011111111;
														assign node23798 = (inp[12]) ? 16'b0000000000011111 : node23799;
															assign node23799 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node23803 = (inp[10]) ? node23807 : node23804;
														assign node23804 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node23807 = (inp[12]) ? node23809 : 16'b0000000000011111;
															assign node23809 = (inp[14]) ? 16'b0000000000001111 : node23810;
																assign node23810 = (inp[6]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node23814 = (inp[14]) ? node23824 : node23815;
													assign node23815 = (inp[12]) ? node23817 : 16'b0000000000111111;
														assign node23817 = (inp[10]) ? node23819 : 16'b0000000000011111;
															assign node23819 = (inp[6]) ? 16'b0000000000001111 : node23820;
																assign node23820 = (inp[9]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node23824 = (inp[9]) ? node23828 : node23825;
														assign node23825 = (inp[10]) ? 16'b0000000000000111 : 16'b0000000000001111;
														assign node23828 = (inp[12]) ? 16'b0000000000001111 : node23829;
															assign node23829 = (inp[10]) ? 16'b0000000000001111 : node23830;
																assign node23830 = (inp[6]) ? 16'b0000000000001111 : 16'b0000000000011111;
										assign node23835 = (inp[6]) ? node23847 : node23836;
											assign node23836 = (inp[12]) ? node23842 : node23837;
												assign node23837 = (inp[13]) ? 16'b0000000000011111 : node23838;
													assign node23838 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000011111111;
												assign node23842 = (inp[13]) ? 16'b0000000000001111 : node23843;
													assign node23843 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000000001111;
											assign node23847 = (inp[13]) ? node23857 : node23848;
												assign node23848 = (inp[10]) ? node23854 : node23849;
													assign node23849 = (inp[5]) ? node23851 : 16'b0000000000011111;
														assign node23851 = (inp[9]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node23854 = (inp[12]) ? 16'b0000000000000111 : 16'b0000000000001111;
												assign node23857 = (inp[5]) ? node23861 : node23858;
													assign node23858 = (inp[14]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node23861 = (inp[12]) ? node23865 : node23862;
														assign node23862 = (inp[14]) ? 16'b0000000000000111 : 16'b0000000000001111;
														assign node23865 = (inp[10]) ? node23871 : node23866;
															assign node23866 = (inp[9]) ? node23868 : 16'b0000000000000111;
																assign node23868 = (inp[14]) ? 16'b0000000000000011 : 16'b0000000000000111;
															assign node23871 = (inp[14]) ? node23873 : 16'b0000000000000011;
																assign node23873 = (inp[9]) ? 16'b0000000000000001 : 16'b0000000000000011;
							assign node23876 = (inp[11]) ? node24058 : node23877;
								assign node23877 = (inp[9]) ? node23955 : node23878;
									assign node23878 = (inp[12]) ? node23916 : node23879;
										assign node23879 = (inp[14]) ? node23893 : node23880;
											assign node23880 = (inp[15]) ? node23890 : node23881;
												assign node23881 = (inp[3]) ? 16'b0000000011111111 : node23882;
													assign node23882 = (inp[13]) ? node23884 : 16'b0000000111111111;
														assign node23884 = (inp[5]) ? 16'b0000000001111111 : node23885;
															assign node23885 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node23890 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node23893 = (inp[15]) ? node23911 : node23894;
												assign node23894 = (inp[10]) ? node23900 : node23895;
													assign node23895 = (inp[3]) ? node23897 : 16'b0000000011111111;
														assign node23897 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node23900 = (inp[3]) ? node23904 : node23901;
														assign node23901 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node23904 = (inp[6]) ? node23906 : 16'b0000000000111111;
															assign node23906 = (inp[5]) ? 16'b0000000000011111 : node23907;
																assign node23907 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node23911 = (inp[6]) ? node23913 : 16'b0000000000111111;
													assign node23913 = (inp[13]) ? 16'b0000000000001111 : 16'b0000000000111111;
										assign node23916 = (inp[15]) ? node23938 : node23917;
											assign node23917 = (inp[6]) ? node23927 : node23918;
												assign node23918 = (inp[3]) ? 16'b0000000000111111 : node23919;
													assign node23919 = (inp[10]) ? node23921 : 16'b0000000001111111;
														assign node23921 = (inp[14]) ? 16'b0000000000111111 : node23922;
															assign node23922 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node23927 = (inp[14]) ? node23933 : node23928;
													assign node23928 = (inp[5]) ? 16'b0000000000111111 : node23929;
														assign node23929 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node23933 = (inp[3]) ? 16'b0000000000001111 : node23934;
														assign node23934 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node23938 = (inp[10]) ? node23946 : node23939;
												assign node23939 = (inp[14]) ? node23943 : node23940;
													assign node23940 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000000011111;
													assign node23943 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000000001111;
												assign node23946 = (inp[6]) ? 16'b0000000000000111 : node23947;
													assign node23947 = (inp[3]) ? node23949 : 16'b0000000000011111;
														assign node23949 = (inp[5]) ? node23951 : 16'b0000000000011111;
															assign node23951 = (inp[14]) ? 16'b0000000000000111 : 16'b0000000000001111;
									assign node23955 = (inp[14]) ? node23997 : node23956;
										assign node23956 = (inp[15]) ? node23974 : node23957;
											assign node23957 = (inp[12]) ? node23967 : node23958;
												assign node23958 = (inp[3]) ? node23960 : 16'b0000000001111111;
													assign node23960 = (inp[5]) ? 16'b0000000000011111 : node23961;
														assign node23961 = (inp[13]) ? 16'b0000000000111111 : node23962;
															assign node23962 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000011111111;
												assign node23967 = (inp[13]) ? 16'b0000000000011111 : node23968;
													assign node23968 = (inp[3]) ? node23970 : 16'b0000000000111111;
														assign node23970 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node23974 = (inp[10]) ? node23982 : node23975;
												assign node23975 = (inp[13]) ? 16'b0000000000011111 : node23976;
													assign node23976 = (inp[6]) ? node23978 : 16'b0000000001111111;
														assign node23978 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node23982 = (inp[6]) ? node23994 : node23983;
													assign node23983 = (inp[12]) ? node23991 : node23984;
														assign node23984 = (inp[5]) ? 16'b0000000000011111 : node23985;
															assign node23985 = (inp[13]) ? node23987 : 16'b0000000000111111;
																assign node23987 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node23991 = (inp[3]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node23994 = (inp[3]) ? 16'b0000000000000111 : 16'b0000000000001111;
										assign node23997 = (inp[6]) ? node24031 : node23998;
											assign node23998 = (inp[3]) ? node24014 : node23999;
												assign node23999 = (inp[5]) ? node24005 : node24000;
													assign node24000 = (inp[13]) ? 16'b0000000000111111 : node24001;
														assign node24001 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node24005 = (inp[10]) ? node24011 : node24006;
														assign node24006 = (inp[15]) ? node24008 : 16'b0000000000111111;
															assign node24008 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node24011 = (inp[15]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node24014 = (inp[10]) ? node24022 : node24015;
													assign node24015 = (inp[15]) ? node24019 : node24016;
														assign node24016 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node24019 = (inp[12]) ? 16'b0000000000000111 : 16'b0000000000011111;
													assign node24022 = (inp[12]) ? 16'b0000000000001111 : node24023;
														assign node24023 = (inp[13]) ? node24025 : 16'b0000000000011111;
															assign node24025 = (inp[5]) ? 16'b0000000000001111 : node24026;
																assign node24026 = (inp[15]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node24031 = (inp[13]) ? node24045 : node24032;
												assign node24032 = (inp[15]) ? node24038 : node24033;
													assign node24033 = (inp[10]) ? node24035 : 16'b0000000000011111;
														assign node24035 = (inp[3]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node24038 = (inp[5]) ? 16'b0000000000001111 : node24039;
														assign node24039 = (inp[12]) ? node24041 : 16'b0000000000001111;
															assign node24041 = (inp[10]) ? 16'b0000000000000111 : 16'b0000000000001111;
												assign node24045 = (inp[5]) ? 16'b0000000000000111 : node24046;
													assign node24046 = (inp[10]) ? node24050 : node24047;
														assign node24047 = (inp[15]) ? 16'b0000000000001111 : 16'b0000000000011111;
														assign node24050 = (inp[3]) ? node24052 : 16'b0000000000001111;
															assign node24052 = (inp[12]) ? 16'b0000000000000111 : node24053;
																assign node24053 = (inp[15]) ? 16'b0000000000000111 : 16'b0000000000001111;
								assign node24058 = (inp[6]) ? node24166 : node24059;
									assign node24059 = (inp[12]) ? node24115 : node24060;
										assign node24060 = (inp[10]) ? node24082 : node24061;
											assign node24061 = (inp[3]) ? node24073 : node24062;
												assign node24062 = (inp[9]) ? node24070 : node24063;
													assign node24063 = (inp[5]) ? 16'b0000000001111111 : node24064;
														assign node24064 = (inp[15]) ? 16'b0000000001111111 : node24065;
															assign node24065 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node24070 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000001111111;
												assign node24073 = (inp[9]) ? node24077 : node24074;
													assign node24074 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000001111111;
													assign node24077 = (inp[13]) ? 16'b0000000000011111 : node24078;
														assign node24078 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node24082 = (inp[13]) ? node24100 : node24083;
												assign node24083 = (inp[9]) ? node24095 : node24084;
													assign node24084 = (inp[14]) ? node24090 : node24085;
														assign node24085 = (inp[3]) ? 16'b0000000000111111 : node24086;
															assign node24086 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node24090 = (inp[5]) ? node24092 : 16'b0000000000111111;
															assign node24092 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node24095 = (inp[3]) ? node24097 : 16'b0000000000011111;
														assign node24097 = (inp[14]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node24100 = (inp[14]) ? node24104 : node24101;
													assign node24101 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000000011111;
													assign node24104 = (inp[5]) ? node24110 : node24105;
														assign node24105 = (inp[3]) ? 16'b0000000000001111 : node24106;
															assign node24106 = (inp[15]) ? 16'b0000000000001111 : 16'b0000000000011111;
														assign node24110 = (inp[9]) ? node24112 : 16'b0000000000001111;
															assign node24112 = (inp[3]) ? 16'b0000000000000011 : 16'b0000000000000111;
										assign node24115 = (inp[14]) ? node24143 : node24116;
											assign node24116 = (inp[10]) ? node24130 : node24117;
												assign node24117 = (inp[9]) ? node24125 : node24118;
													assign node24118 = (inp[13]) ? node24120 : 16'b0000000001111111;
														assign node24120 = (inp[3]) ? node24122 : 16'b0000000000111111;
															assign node24122 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node24125 = (inp[13]) ? 16'b0000000000011111 : node24126;
														assign node24126 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000001111111;
												assign node24130 = (inp[3]) ? node24136 : node24131;
													assign node24131 = (inp[9]) ? node24133 : 16'b0000000000011111;
														assign node24133 = (inp[13]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node24136 = (inp[15]) ? node24138 : 16'b0000000000001111;
														assign node24138 = (inp[5]) ? node24140 : 16'b0000000000001111;
															assign node24140 = (inp[13]) ? 16'b0000000000000011 : 16'b0000000000000111;
											assign node24143 = (inp[13]) ? node24155 : node24144;
												assign node24144 = (inp[3]) ? node24150 : node24145;
													assign node24145 = (inp[15]) ? node24147 : 16'b0000000000111111;
														assign node24147 = (inp[5]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node24150 = (inp[15]) ? node24152 : 16'b0000000000001111;
														assign node24152 = (inp[10]) ? 16'b0000000000000111 : 16'b0000000000001111;
												assign node24155 = (inp[3]) ? node24161 : node24156;
													assign node24156 = (inp[10]) ? 16'b0000000000000111 : node24157;
														assign node24157 = (inp[15]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node24161 = (inp[10]) ? 16'b0000000000000111 : node24162;
														assign node24162 = (inp[9]) ? 16'b0000000000000011 : 16'b0000000000000111;
									assign node24166 = (inp[10]) ? node24218 : node24167;
										assign node24167 = (inp[14]) ? node24189 : node24168;
											assign node24168 = (inp[13]) ? node24184 : node24169;
												assign node24169 = (inp[9]) ? node24177 : node24170;
													assign node24170 = (inp[5]) ? node24174 : node24171;
														assign node24171 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node24174 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node24177 = (inp[12]) ? 16'b0000000000001111 : node24178;
														assign node24178 = (inp[15]) ? 16'b0000000000011111 : node24179;
															assign node24179 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node24184 = (inp[15]) ? node24186 : 16'b0000000000011111;
													assign node24186 = (inp[9]) ? 16'b0000000000000111 : 16'b0000000000001111;
											assign node24189 = (inp[3]) ? node24203 : node24190;
												assign node24190 = (inp[5]) ? node24198 : node24191;
													assign node24191 = (inp[12]) ? node24193 : 16'b0000000000011111;
														assign node24193 = (inp[13]) ? node24195 : 16'b0000000000011111;
															assign node24195 = (inp[9]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node24198 = (inp[12]) ? 16'b0000000000000111 : node24199;
														assign node24199 = (inp[15]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node24203 = (inp[12]) ? node24213 : node24204;
													assign node24204 = (inp[5]) ? node24210 : node24205;
														assign node24205 = (inp[13]) ? 16'b0000000000001111 : node24206;
															assign node24206 = (inp[9]) ? 16'b0000000000001111 : 16'b0000000000011111;
														assign node24210 = (inp[13]) ? 16'b0000000000000111 : 16'b0000000000001111;
													assign node24213 = (inp[13]) ? 16'b0000000000000011 : node24214;
														assign node24214 = (inp[9]) ? 16'b0000000000000111 : 16'b0000000000001111;
										assign node24218 = (inp[5]) ? node24248 : node24219;
											assign node24219 = (inp[3]) ? node24233 : node24220;
												assign node24220 = (inp[9]) ? node24228 : node24221;
													assign node24221 = (inp[14]) ? 16'b0000000000111111 : node24222;
														assign node24222 = (inp[12]) ? 16'b0000000000011111 : node24223;
															assign node24223 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node24228 = (inp[15]) ? 16'b0000000000011111 : node24229;
														assign node24229 = (inp[12]) ? 16'b0000000000000111 : 16'b0000000000001111;
												assign node24233 = (inp[9]) ? node24241 : node24234;
													assign node24234 = (inp[14]) ? node24238 : node24235;
														assign node24235 = (inp[13]) ? 16'b0000000000001111 : 16'b0000000000011111;
														assign node24238 = (inp[13]) ? 16'b0000000000000111 : 16'b0000000000001111;
													assign node24241 = (inp[15]) ? node24245 : node24242;
														assign node24242 = (inp[14]) ? 16'b0000000000000111 : 16'b0000000000001111;
														assign node24245 = (inp[14]) ? 16'b0000000000000011 : 16'b0000000000000111;
											assign node24248 = (inp[13]) ? node24258 : node24249;
												assign node24249 = (inp[9]) ? 16'b0000000000000111 : node24250;
													assign node24250 = (inp[3]) ? node24254 : node24251;
														assign node24251 = (inp[12]) ? 16'b0000000000001111 : 16'b0000000000011111;
														assign node24254 = (inp[12]) ? 16'b0000000000000111 : 16'b0000000000001111;
												assign node24258 = (inp[14]) ? node24268 : node24259;
													assign node24259 = (inp[9]) ? node24263 : node24260;
														assign node24260 = (inp[15]) ? 16'b0000000000000111 : 16'b0000000000001111;
														assign node24263 = (inp[15]) ? node24265 : 16'b0000000000000111;
															assign node24265 = (inp[12]) ? 16'b0000000000000011 : 16'b0000000000000111;
													assign node24268 = (inp[9]) ? node24276 : node24269;
														assign node24269 = (inp[3]) ? node24271 : 16'b0000000000000111;
															assign node24271 = (inp[15]) ? node24273 : 16'b0000000000000011;
																assign node24273 = (inp[12]) ? 16'b0000000000000001 : 16'b0000000000000011;
														assign node24276 = (inp[12]) ? node24278 : 16'b0000000000000001;
															assign node24278 = (inp[3]) ? 16'b0000000000000000 : 16'b0000000000000001;

endmodule