module dtc_split75_bm75 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node7;
	wire [3-1:0] node8;
	wire [3-1:0] node9;
	wire [3-1:0] node12;
	wire [3-1:0] node15;
	wire [3-1:0] node16;
	wire [3-1:0] node20;
	wire [3-1:0] node21;
	wire [3-1:0] node22;
	wire [3-1:0] node25;
	wire [3-1:0] node28;
	wire [3-1:0] node29;
	wire [3-1:0] node32;
	wire [3-1:0] node35;
	wire [3-1:0] node36;
	wire [3-1:0] node37;
	wire [3-1:0] node38;
	wire [3-1:0] node41;
	wire [3-1:0] node44;
	wire [3-1:0] node45;
	wire [3-1:0] node48;
	wire [3-1:0] node51;
	wire [3-1:0] node52;
	wire [3-1:0] node53;
	wire [3-1:0] node56;
	wire [3-1:0] node59;
	wire [3-1:0] node60;
	wire [3-1:0] node63;
	wire [3-1:0] node66;
	wire [3-1:0] node67;
	wire [3-1:0] node68;
	wire [3-1:0] node70;
	wire [3-1:0] node72;
	wire [3-1:0] node76;
	wire [3-1:0] node77;
	wire [3-1:0] node78;
	wire [3-1:0] node80;
	wire [3-1:0] node84;
	wire [3-1:0] node85;
	wire [3-1:0] node86;
	wire [3-1:0] node89;
	wire [3-1:0] node92;
	wire [3-1:0] node93;
	wire [3-1:0] node96;
	wire [3-1:0] node99;
	wire [3-1:0] node100;
	wire [3-1:0] node101;
	wire [3-1:0] node102;
	wire [3-1:0] node103;
	wire [3-1:0] node105;
	wire [3-1:0] node110;
	wire [3-1:0] node111;
	wire [3-1:0] node112;
	wire [3-1:0] node113;
	wire [3-1:0] node117;
	wire [3-1:0] node118;
	wire [3-1:0] node122;
	wire [3-1:0] node123;
	wire [3-1:0] node125;
	wire [3-1:0] node129;
	wire [3-1:0] node131;
	wire [3-1:0] node132;
	wire [3-1:0] node133;
	wire [3-1:0] node134;
	wire [3-1:0] node140;
	wire [3-1:0] node141;
	wire [3-1:0] node142;
	wire [3-1:0] node143;
	wire [3-1:0] node144;
	wire [3-1:0] node145;
	wire [3-1:0] node146;
	wire [3-1:0] node149;
	wire [3-1:0] node152;
	wire [3-1:0] node153;
	wire [3-1:0] node156;
	wire [3-1:0] node159;
	wire [3-1:0] node160;
	wire [3-1:0] node161;
	wire [3-1:0] node164;
	wire [3-1:0] node167;
	wire [3-1:0] node168;
	wire [3-1:0] node171;
	wire [3-1:0] node174;
	wire [3-1:0] node175;
	wire [3-1:0] node176;
	wire [3-1:0] node177;
	wire [3-1:0] node180;
	wire [3-1:0] node183;
	wire [3-1:0] node184;
	wire [3-1:0] node187;
	wire [3-1:0] node190;
	wire [3-1:0] node191;
	wire [3-1:0] node192;
	wire [3-1:0] node195;
	wire [3-1:0] node198;
	wire [3-1:0] node199;
	wire [3-1:0] node202;
	wire [3-1:0] node205;
	wire [3-1:0] node206;
	wire [3-1:0] node207;
	wire [3-1:0] node208;
	wire [3-1:0] node210;
	wire [3-1:0] node213;
	wire [3-1:0] node214;
	wire [3-1:0] node217;
	wire [3-1:0] node220;
	wire [3-1:0] node221;
	wire [3-1:0] node222;
	wire [3-1:0] node225;
	wire [3-1:0] node228;
	wire [3-1:0] node229;
	wire [3-1:0] node232;
	wire [3-1:0] node235;
	wire [3-1:0] node236;
	wire [3-1:0] node237;
	wire [3-1:0] node238;
	wire [3-1:0] node241;
	wire [3-1:0] node244;
	wire [3-1:0] node245;
	wire [3-1:0] node248;
	wire [3-1:0] node251;
	wire [3-1:0] node252;
	wire [3-1:0] node253;
	wire [3-1:0] node256;
	wire [3-1:0] node259;
	wire [3-1:0] node260;
	wire [3-1:0] node263;
	wire [3-1:0] node266;
	wire [3-1:0] node267;
	wire [3-1:0] node268;
	wire [3-1:0] node269;
	wire [3-1:0] node270;
	wire [3-1:0] node271;
	wire [3-1:0] node274;
	wire [3-1:0] node277;
	wire [3-1:0] node279;
	wire [3-1:0] node282;
	wire [3-1:0] node283;
	wire [3-1:0] node284;
	wire [3-1:0] node287;
	wire [3-1:0] node290;
	wire [3-1:0] node291;
	wire [3-1:0] node294;
	wire [3-1:0] node297;
	wire [3-1:0] node298;
	wire [3-1:0] node299;
	wire [3-1:0] node300;
	wire [3-1:0] node303;
	wire [3-1:0] node306;
	wire [3-1:0] node308;
	wire [3-1:0] node311;
	wire [3-1:0] node312;
	wire [3-1:0] node313;
	wire [3-1:0] node316;
	wire [3-1:0] node319;
	wire [3-1:0] node320;
	wire [3-1:0] node323;
	wire [3-1:0] node326;
	wire [3-1:0] node327;
	wire [3-1:0] node328;
	wire [3-1:0] node329;
	wire [3-1:0] node330;
	wire [3-1:0] node335;
	wire [3-1:0] node336;
	wire [3-1:0] node337;
	wire [3-1:0] node340;
	wire [3-1:0] node343;
	wire [3-1:0] node345;
	wire [3-1:0] node348;
	wire [3-1:0] node349;
	wire [3-1:0] node350;
	wire [3-1:0] node351;
	wire [3-1:0] node354;
	wire [3-1:0] node357;
	wire [3-1:0] node358;
	wire [3-1:0] node362;
	wire [3-1:0] node363;
	wire [3-1:0] node364;
	wire [3-1:0] node367;
	wire [3-1:0] node370;
	wire [3-1:0] node371;
	wire [3-1:0] node374;
	wire [3-1:0] node377;
	wire [3-1:0] node378;
	wire [3-1:0] node379;
	wire [3-1:0] node380;
	wire [3-1:0] node381;
	wire [3-1:0] node382;
	wire [3-1:0] node383;
	wire [3-1:0] node384;
	wire [3-1:0] node388;
	wire [3-1:0] node389;
	wire [3-1:0] node392;
	wire [3-1:0] node395;
	wire [3-1:0] node396;
	wire [3-1:0] node397;
	wire [3-1:0] node400;
	wire [3-1:0] node403;
	wire [3-1:0] node404;
	wire [3-1:0] node407;
	wire [3-1:0] node410;
	wire [3-1:0] node411;
	wire [3-1:0] node412;
	wire [3-1:0] node413;
	wire [3-1:0] node416;
	wire [3-1:0] node419;
	wire [3-1:0] node420;
	wire [3-1:0] node423;
	wire [3-1:0] node426;
	wire [3-1:0] node427;
	wire [3-1:0] node428;
	wire [3-1:0] node432;
	wire [3-1:0] node433;
	wire [3-1:0] node436;
	wire [3-1:0] node439;
	wire [3-1:0] node440;
	wire [3-1:0] node441;
	wire [3-1:0] node442;
	wire [3-1:0] node443;
	wire [3-1:0] node446;
	wire [3-1:0] node449;
	wire [3-1:0] node450;
	wire [3-1:0] node453;
	wire [3-1:0] node456;
	wire [3-1:0] node457;
	wire [3-1:0] node458;
	wire [3-1:0] node461;
	wire [3-1:0] node464;
	wire [3-1:0] node465;
	wire [3-1:0] node468;
	wire [3-1:0] node471;
	wire [3-1:0] node472;
	wire [3-1:0] node473;
	wire [3-1:0] node474;
	wire [3-1:0] node477;
	wire [3-1:0] node480;
	wire [3-1:0] node481;
	wire [3-1:0] node484;
	wire [3-1:0] node487;
	wire [3-1:0] node488;
	wire [3-1:0] node489;
	wire [3-1:0] node492;
	wire [3-1:0] node495;
	wire [3-1:0] node496;
	wire [3-1:0] node499;
	wire [3-1:0] node502;
	wire [3-1:0] node503;
	wire [3-1:0] node504;
	wire [3-1:0] node505;
	wire [3-1:0] node506;
	wire [3-1:0] node507;
	wire [3-1:0] node510;
	wire [3-1:0] node513;
	wire [3-1:0] node514;
	wire [3-1:0] node517;
	wire [3-1:0] node520;
	wire [3-1:0] node521;
	wire [3-1:0] node522;
	wire [3-1:0] node525;
	wire [3-1:0] node528;
	wire [3-1:0] node529;
	wire [3-1:0] node532;
	wire [3-1:0] node535;
	wire [3-1:0] node536;
	wire [3-1:0] node537;
	wire [3-1:0] node539;
	wire [3-1:0] node542;
	wire [3-1:0] node543;
	wire [3-1:0] node546;
	wire [3-1:0] node549;
	wire [3-1:0] node550;
	wire [3-1:0] node551;
	wire [3-1:0] node555;
	wire [3-1:0] node556;
	wire [3-1:0] node559;
	wire [3-1:0] node562;
	wire [3-1:0] node563;
	wire [3-1:0] node564;
	wire [3-1:0] node566;
	wire [3-1:0] node567;
	wire [3-1:0] node571;
	wire [3-1:0] node572;
	wire [3-1:0] node573;
	wire [3-1:0] node576;
	wire [3-1:0] node579;
	wire [3-1:0] node580;
	wire [3-1:0] node584;
	wire [3-1:0] node585;
	wire [3-1:0] node586;
	wire [3-1:0] node587;
	wire [3-1:0] node590;
	wire [3-1:0] node593;
	wire [3-1:0] node594;
	wire [3-1:0] node598;
	wire [3-1:0] node599;
	wire [3-1:0] node600;
	wire [3-1:0] node603;
	wire [3-1:0] node606;
	wire [3-1:0] node607;
	wire [3-1:0] node610;
	wire [3-1:0] node613;
	wire [3-1:0] node614;
	wire [3-1:0] node615;
	wire [3-1:0] node616;
	wire [3-1:0] node617;
	wire [3-1:0] node618;
	wire [3-1:0] node619;
	wire [3-1:0] node622;
	wire [3-1:0] node625;
	wire [3-1:0] node626;
	wire [3-1:0] node629;
	wire [3-1:0] node632;
	wire [3-1:0] node633;
	wire [3-1:0] node634;
	wire [3-1:0] node637;
	wire [3-1:0] node640;
	wire [3-1:0] node641;
	wire [3-1:0] node644;
	wire [3-1:0] node647;
	wire [3-1:0] node648;
	wire [3-1:0] node649;
	wire [3-1:0] node650;
	wire [3-1:0] node654;
	wire [3-1:0] node655;
	wire [3-1:0] node658;
	wire [3-1:0] node661;
	wire [3-1:0] node662;
	wire [3-1:0] node663;
	wire [3-1:0] node667;
	wire [3-1:0] node668;
	wire [3-1:0] node671;
	wire [3-1:0] node674;
	wire [3-1:0] node675;
	wire [3-1:0] node676;
	wire [3-1:0] node677;
	wire [3-1:0] node678;
	wire [3-1:0] node681;
	wire [3-1:0] node684;
	wire [3-1:0] node685;
	wire [3-1:0] node688;
	wire [3-1:0] node691;
	wire [3-1:0] node692;
	wire [3-1:0] node693;
	wire [3-1:0] node696;
	wire [3-1:0] node699;
	wire [3-1:0] node700;
	wire [3-1:0] node703;
	wire [3-1:0] node706;
	wire [3-1:0] node707;
	wire [3-1:0] node708;
	wire [3-1:0] node709;
	wire [3-1:0] node712;
	wire [3-1:0] node715;
	wire [3-1:0] node716;
	wire [3-1:0] node719;
	wire [3-1:0] node722;
	wire [3-1:0] node723;
	wire [3-1:0] node724;
	wire [3-1:0] node727;
	wire [3-1:0] node730;
	wire [3-1:0] node731;
	wire [3-1:0] node734;
	wire [3-1:0] node737;
	wire [3-1:0] node738;
	wire [3-1:0] node739;
	wire [3-1:0] node740;
	wire [3-1:0] node741;
	wire [3-1:0] node742;
	wire [3-1:0] node745;
	wire [3-1:0] node748;
	wire [3-1:0] node749;
	wire [3-1:0] node752;
	wire [3-1:0] node755;
	wire [3-1:0] node756;
	wire [3-1:0] node757;
	wire [3-1:0] node760;
	wire [3-1:0] node763;
	wire [3-1:0] node764;
	wire [3-1:0] node767;
	wire [3-1:0] node770;
	wire [3-1:0] node771;
	wire [3-1:0] node772;
	wire [3-1:0] node773;
	wire [3-1:0] node777;
	wire [3-1:0] node779;
	wire [3-1:0] node782;
	wire [3-1:0] node783;
	wire [3-1:0] node784;
	wire [3-1:0] node787;
	wire [3-1:0] node790;
	wire [3-1:0] node791;
	wire [3-1:0] node794;
	wire [3-1:0] node797;
	wire [3-1:0] node798;
	wire [3-1:0] node799;
	wire [3-1:0] node800;
	wire [3-1:0] node802;
	wire [3-1:0] node805;
	wire [3-1:0] node806;
	wire [3-1:0] node809;
	wire [3-1:0] node812;
	wire [3-1:0] node813;
	wire [3-1:0] node814;
	wire [3-1:0] node817;
	wire [3-1:0] node820;
	wire [3-1:0] node821;
	wire [3-1:0] node824;
	wire [3-1:0] node827;
	wire [3-1:0] node828;
	wire [3-1:0] node829;
	wire [3-1:0] node830;
	wire [3-1:0] node833;
	wire [3-1:0] node836;
	wire [3-1:0] node837;
	wire [3-1:0] node840;
	wire [3-1:0] node843;
	wire [3-1:0] node844;
	wire [3-1:0] node845;
	wire [3-1:0] node848;
	wire [3-1:0] node851;
	wire [3-1:0] node852;
	wire [3-1:0] node855;
	wire [3-1:0] node858;
	wire [3-1:0] node859;
	wire [3-1:0] node860;
	wire [3-1:0] node861;
	wire [3-1:0] node862;
	wire [3-1:0] node863;
	wire [3-1:0] node864;
	wire [3-1:0] node865;
	wire [3-1:0] node866;
	wire [3-1:0] node869;
	wire [3-1:0] node872;
	wire [3-1:0] node873;
	wire [3-1:0] node876;
	wire [3-1:0] node879;
	wire [3-1:0] node880;
	wire [3-1:0] node881;
	wire [3-1:0] node884;
	wire [3-1:0] node887;
	wire [3-1:0] node888;
	wire [3-1:0] node891;
	wire [3-1:0] node894;
	wire [3-1:0] node895;
	wire [3-1:0] node896;
	wire [3-1:0] node897;
	wire [3-1:0] node900;
	wire [3-1:0] node903;
	wire [3-1:0] node904;
	wire [3-1:0] node908;
	wire [3-1:0] node910;
	wire [3-1:0] node911;
	wire [3-1:0] node914;
	wire [3-1:0] node917;
	wire [3-1:0] node918;
	wire [3-1:0] node919;
	wire [3-1:0] node920;
	wire [3-1:0] node921;
	wire [3-1:0] node924;
	wire [3-1:0] node927;
	wire [3-1:0] node928;
	wire [3-1:0] node932;
	wire [3-1:0] node933;
	wire [3-1:0] node934;
	wire [3-1:0] node937;
	wire [3-1:0] node940;
	wire [3-1:0] node941;
	wire [3-1:0] node944;
	wire [3-1:0] node947;
	wire [3-1:0] node948;
	wire [3-1:0] node949;
	wire [3-1:0] node950;
	wire [3-1:0] node953;
	wire [3-1:0] node956;
	wire [3-1:0] node957;
	wire [3-1:0] node960;
	wire [3-1:0] node963;
	wire [3-1:0] node964;
	wire [3-1:0] node965;
	wire [3-1:0] node968;
	wire [3-1:0] node971;
	wire [3-1:0] node972;
	wire [3-1:0] node975;
	wire [3-1:0] node978;
	wire [3-1:0] node979;
	wire [3-1:0] node980;
	wire [3-1:0] node981;
	wire [3-1:0] node982;
	wire [3-1:0] node984;
	wire [3-1:0] node987;
	wire [3-1:0] node988;
	wire [3-1:0] node991;
	wire [3-1:0] node994;
	wire [3-1:0] node995;
	wire [3-1:0] node996;
	wire [3-1:0] node999;
	wire [3-1:0] node1002;
	wire [3-1:0] node1003;
	wire [3-1:0] node1006;
	wire [3-1:0] node1009;
	wire [3-1:0] node1010;
	wire [3-1:0] node1011;
	wire [3-1:0] node1012;
	wire [3-1:0] node1015;
	wire [3-1:0] node1018;
	wire [3-1:0] node1019;
	wire [3-1:0] node1022;
	wire [3-1:0] node1025;
	wire [3-1:0] node1026;
	wire [3-1:0] node1027;
	wire [3-1:0] node1030;
	wire [3-1:0] node1033;
	wire [3-1:0] node1034;
	wire [3-1:0] node1037;
	wire [3-1:0] node1040;
	wire [3-1:0] node1041;
	wire [3-1:0] node1042;
	wire [3-1:0] node1043;
	wire [3-1:0] node1044;
	wire [3-1:0] node1047;
	wire [3-1:0] node1050;
	wire [3-1:0] node1051;
	wire [3-1:0] node1054;
	wire [3-1:0] node1057;
	wire [3-1:0] node1058;
	wire [3-1:0] node1059;
	wire [3-1:0] node1062;
	wire [3-1:0] node1065;
	wire [3-1:0] node1066;
	wire [3-1:0] node1069;
	wire [3-1:0] node1072;
	wire [3-1:0] node1073;
	wire [3-1:0] node1074;
	wire [3-1:0] node1075;
	wire [3-1:0] node1078;
	wire [3-1:0] node1081;
	wire [3-1:0] node1082;
	wire [3-1:0] node1085;
	wire [3-1:0] node1088;
	wire [3-1:0] node1089;
	wire [3-1:0] node1090;
	wire [3-1:0] node1093;
	wire [3-1:0] node1096;
	wire [3-1:0] node1097;
	wire [3-1:0] node1101;
	wire [3-1:0] node1102;
	wire [3-1:0] node1103;
	wire [3-1:0] node1104;
	wire [3-1:0] node1105;
	wire [3-1:0] node1106;
	wire [3-1:0] node1108;
	wire [3-1:0] node1111;
	wire [3-1:0] node1112;
	wire [3-1:0] node1115;
	wire [3-1:0] node1118;
	wire [3-1:0] node1119;
	wire [3-1:0] node1121;
	wire [3-1:0] node1125;
	wire [3-1:0] node1127;
	wire [3-1:0] node1129;
	wire [3-1:0] node1130;
	wire [3-1:0] node1134;
	wire [3-1:0] node1135;
	wire [3-1:0] node1136;
	wire [3-1:0] node1137;
	wire [3-1:0] node1138;
	wire [3-1:0] node1141;
	wire [3-1:0] node1144;
	wire [3-1:0] node1145;
	wire [3-1:0] node1148;
	wire [3-1:0] node1151;
	wire [3-1:0] node1152;
	wire [3-1:0] node1153;
	wire [3-1:0] node1156;
	wire [3-1:0] node1159;
	wire [3-1:0] node1160;
	wire [3-1:0] node1163;
	wire [3-1:0] node1166;
	wire [3-1:0] node1167;
	wire [3-1:0] node1168;
	wire [3-1:0] node1170;
	wire [3-1:0] node1173;
	wire [3-1:0] node1174;
	wire [3-1:0] node1177;
	wire [3-1:0] node1180;
	wire [3-1:0] node1182;
	wire [3-1:0] node1184;
	wire [3-1:0] node1187;
	wire [3-1:0] node1188;
	wire [3-1:0] node1189;
	wire [3-1:0] node1190;
	wire [3-1:0] node1191;
	wire [3-1:0] node1192;
	wire [3-1:0] node1195;
	wire [3-1:0] node1198;
	wire [3-1:0] node1199;
	wire [3-1:0] node1202;
	wire [3-1:0] node1205;
	wire [3-1:0] node1206;
	wire [3-1:0] node1207;
	wire [3-1:0] node1210;
	wire [3-1:0] node1213;
	wire [3-1:0] node1214;
	wire [3-1:0] node1217;
	wire [3-1:0] node1220;
	wire [3-1:0] node1221;
	wire [3-1:0] node1222;
	wire [3-1:0] node1223;
	wire [3-1:0] node1226;
	wire [3-1:0] node1229;
	wire [3-1:0] node1230;
	wire [3-1:0] node1233;
	wire [3-1:0] node1236;
	wire [3-1:0] node1238;
	wire [3-1:0] node1240;
	wire [3-1:0] node1243;
	wire [3-1:0] node1244;
	wire [3-1:0] node1245;
	wire [3-1:0] node1246;
	wire [3-1:0] node1247;
	wire [3-1:0] node1250;
	wire [3-1:0] node1253;
	wire [3-1:0] node1254;
	wire [3-1:0] node1257;
	wire [3-1:0] node1260;
	wire [3-1:0] node1261;
	wire [3-1:0] node1262;
	wire [3-1:0] node1265;
	wire [3-1:0] node1268;
	wire [3-1:0] node1269;
	wire [3-1:0] node1272;
	wire [3-1:0] node1275;
	wire [3-1:0] node1276;
	wire [3-1:0] node1277;
	wire [3-1:0] node1278;
	wire [3-1:0] node1281;
	wire [3-1:0] node1284;
	wire [3-1:0] node1285;
	wire [3-1:0] node1288;
	wire [3-1:0] node1291;
	wire [3-1:0] node1292;
	wire [3-1:0] node1293;
	wire [3-1:0] node1297;
	wire [3-1:0] node1298;
	wire [3-1:0] node1301;
	wire [3-1:0] node1304;
	wire [3-1:0] node1305;
	wire [3-1:0] node1306;
	wire [3-1:0] node1307;
	wire [3-1:0] node1308;
	wire [3-1:0] node1309;
	wire [3-1:0] node1310;
	wire [3-1:0] node1312;
	wire [3-1:0] node1315;
	wire [3-1:0] node1316;
	wire [3-1:0] node1319;
	wire [3-1:0] node1322;
	wire [3-1:0] node1323;
	wire [3-1:0] node1325;
	wire [3-1:0] node1330;
	wire [3-1:0] node1331;
	wire [3-1:0] node1332;
	wire [3-1:0] node1333;
	wire [3-1:0] node1334;
	wire [3-1:0] node1337;
	wire [3-1:0] node1340;
	wire [3-1:0] node1341;
	wire [3-1:0] node1344;
	wire [3-1:0] node1347;
	wire [3-1:0] node1348;
	wire [3-1:0] node1350;
	wire [3-1:0] node1353;
	wire [3-1:0] node1354;
	wire [3-1:0] node1357;
	wire [3-1:0] node1360;
	wire [3-1:0] node1361;
	wire [3-1:0] node1362;
	wire [3-1:0] node1364;
	wire [3-1:0] node1368;
	wire [3-1:0] node1369;
	wire [3-1:0] node1370;
	wire [3-1:0] node1374;
	wire [3-1:0] node1375;
	wire [3-1:0] node1379;
	wire [3-1:0] node1380;
	wire [3-1:0] node1381;
	wire [3-1:0] node1382;
	wire [3-1:0] node1383;
	wire [3-1:0] node1384;
	wire [3-1:0] node1387;
	wire [3-1:0] node1390;
	wire [3-1:0] node1391;
	wire [3-1:0] node1394;
	wire [3-1:0] node1397;
	wire [3-1:0] node1398;
	wire [3-1:0] node1399;
	wire [3-1:0] node1402;
	wire [3-1:0] node1405;
	wire [3-1:0] node1406;
	wire [3-1:0] node1409;
	wire [3-1:0] node1412;
	wire [3-1:0] node1413;
	wire [3-1:0] node1414;
	wire [3-1:0] node1416;
	wire [3-1:0] node1419;
	wire [3-1:0] node1420;
	wire [3-1:0] node1423;
	wire [3-1:0] node1426;
	wire [3-1:0] node1428;
	wire [3-1:0] node1430;
	wire [3-1:0] node1433;
	wire [3-1:0] node1434;
	wire [3-1:0] node1435;
	wire [3-1:0] node1436;
	wire [3-1:0] node1437;
	wire [3-1:0] node1441;
	wire [3-1:0] node1442;
	wire [3-1:0] node1445;
	wire [3-1:0] node1448;
	wire [3-1:0] node1449;
	wire [3-1:0] node1450;
	wire [3-1:0] node1453;
	wire [3-1:0] node1456;
	wire [3-1:0] node1457;
	wire [3-1:0] node1460;
	wire [3-1:0] node1463;
	wire [3-1:0] node1464;
	wire [3-1:0] node1465;
	wire [3-1:0] node1466;
	wire [3-1:0] node1469;
	wire [3-1:0] node1472;
	wire [3-1:0] node1473;
	wire [3-1:0] node1476;
	wire [3-1:0] node1479;
	wire [3-1:0] node1480;
	wire [3-1:0] node1481;
	wire [3-1:0] node1484;
	wire [3-1:0] node1487;
	wire [3-1:0] node1488;
	wire [3-1:0] node1491;
	wire [3-1:0] node1494;
	wire [3-1:0] node1495;
	wire [3-1:0] node1496;
	wire [3-1:0] node1497;
	wire [3-1:0] node1498;
	wire [3-1:0] node1500;
	wire [3-1:0] node1502;
	wire [3-1:0] node1508;
	wire [3-1:0] node1509;
	wire [3-1:0] node1510;
	wire [3-1:0] node1512;
	wire [3-1:0] node1514;
	wire [3-1:0] node1515;
	wire [3-1:0] node1520;
	wire [3-1:0] node1521;
	wire [3-1:0] node1522;
	wire [3-1:0] node1523;
	wire [3-1:0] node1524;
	wire [3-1:0] node1527;
	wire [3-1:0] node1530;
	wire [3-1:0] node1531;
	wire [3-1:0] node1534;
	wire [3-1:0] node1537;
	wire [3-1:0] node1538;
	wire [3-1:0] node1540;
	wire [3-1:0] node1543;
	wire [3-1:0] node1544;
	wire [3-1:0] node1547;
	wire [3-1:0] node1550;
	wire [3-1:0] node1552;
	wire [3-1:0] node1554;
	wire [3-1:0] node1555;
	wire [3-1:0] node1558;

	assign outp = (inp[3]) ? node858 : node1;
		assign node1 = (inp[9]) ? node377 : node2;
			assign node2 = (inp[4]) ? node140 : node3;
				assign node3 = (inp[6]) ? node99 : node4;
					assign node4 = (inp[0]) ? node66 : node5;
						assign node5 = (inp[5]) ? node35 : node6;
							assign node6 = (inp[10]) ? node20 : node7;
								assign node7 = (inp[1]) ? node15 : node8;
									assign node8 = (inp[7]) ? node12 : node9;
										assign node9 = (inp[11]) ? 3'b101 : 3'b011;
										assign node12 = (inp[11]) ? 3'b011 : 3'b111;
									assign node15 = (inp[7]) ? 3'b111 : node16;
										assign node16 = (inp[2]) ? 3'b111 : 3'b011;
								assign node20 = (inp[7]) ? node28 : node21;
									assign node21 = (inp[2]) ? node25 : node22;
										assign node22 = (inp[8]) ? 3'b101 : 3'b101;
										assign node25 = (inp[11]) ? 3'b001 : 3'b011;
									assign node28 = (inp[1]) ? node32 : node29;
										assign node29 = (inp[11]) ? 3'b101 : 3'b011;
										assign node32 = (inp[11]) ? 3'b011 : 3'b111;
							assign node35 = (inp[1]) ? node51 : node36;
								assign node36 = (inp[11]) ? node44 : node37;
									assign node37 = (inp[10]) ? node41 : node38;
										assign node38 = (inp[7]) ? 3'b011 : 3'b101;
										assign node41 = (inp[7]) ? 3'b101 : 3'b001;
									assign node44 = (inp[7]) ? node48 : node45;
										assign node45 = (inp[10]) ? 3'b110 : 3'b001;
										assign node48 = (inp[10]) ? 3'b001 : 3'b101;
								assign node51 = (inp[10]) ? node59 : node52;
									assign node52 = (inp[7]) ? node56 : node53;
										assign node53 = (inp[2]) ? 3'b011 : 3'b101;
										assign node56 = (inp[11]) ? 3'b011 : 3'b111;
									assign node59 = (inp[7]) ? node63 : node60;
										assign node60 = (inp[8]) ? 3'b101 : 3'b001;
										assign node63 = (inp[11]) ? 3'b101 : 3'b001;
						assign node66 = (inp[10]) ? node76 : node67;
							assign node67 = (inp[7]) ? 3'b111 : node68;
								assign node68 = (inp[11]) ? node70 : 3'b111;
									assign node70 = (inp[5]) ? node72 : 3'b111;
										assign node72 = (inp[1]) ? 3'b111 : 3'b011;
							assign node76 = (inp[5]) ? node84 : node77;
								assign node77 = (inp[1]) ? 3'b111 : node78;
									assign node78 = (inp[7]) ? node80 : 3'b011;
										assign node80 = (inp[2]) ? 3'b111 : 3'b111;
								assign node84 = (inp[7]) ? node92 : node85;
									assign node85 = (inp[1]) ? node89 : node86;
										assign node86 = (inp[11]) ? 3'b101 : 3'b101;
										assign node89 = (inp[8]) ? 3'b011 : 3'b101;
									assign node92 = (inp[11]) ? node96 : node93;
										assign node93 = (inp[1]) ? 3'b111 : 3'b011;
										assign node96 = (inp[2]) ? 3'b011 : 3'b011;
					assign node99 = (inp[0]) ? node129 : node100;
						assign node100 = (inp[5]) ? node110 : node101;
							assign node101 = (inp[2]) ? 3'b111 : node102;
								assign node102 = (inp[7]) ? 3'b111 : node103;
									assign node103 = (inp[10]) ? node105 : 3'b111;
										assign node105 = (inp[8]) ? 3'b111 : 3'b011;
							assign node110 = (inp[1]) ? node122 : node111;
								assign node111 = (inp[10]) ? node117 : node112;
									assign node112 = (inp[7]) ? 3'b111 : node113;
										assign node113 = (inp[8]) ? 3'b111 : 3'b011;
									assign node117 = (inp[11]) ? 3'b101 : node118;
										assign node118 = (inp[8]) ? 3'b011 : 3'b011;
								assign node122 = (inp[7]) ? 3'b111 : node123;
									assign node123 = (inp[10]) ? node125 : 3'b111;
										assign node125 = (inp[2]) ? 3'b011 : 3'b011;
						assign node129 = (inp[5]) ? node131 : 3'b111;
							assign node131 = (inp[1]) ? 3'b111 : node132;
								assign node132 = (inp[8]) ? 3'b111 : node133;
									assign node133 = (inp[7]) ? 3'b111 : node134;
										assign node134 = (inp[10]) ? 3'b011 : 3'b111;
				assign node140 = (inp[6]) ? node266 : node141;
					assign node141 = (inp[0]) ? node205 : node142;
						assign node142 = (inp[10]) ? node174 : node143;
							assign node143 = (inp[5]) ? node159 : node144;
								assign node144 = (inp[7]) ? node152 : node145;
									assign node145 = (inp[1]) ? node149 : node146;
										assign node146 = (inp[11]) ? 3'b110 : 3'b001;
										assign node149 = (inp[8]) ? 3'b101 : 3'b001;
									assign node152 = (inp[1]) ? node156 : node153;
										assign node153 = (inp[8]) ? 3'b101 : 3'b001;
										assign node156 = (inp[2]) ? 3'b001 : 3'b101;
								assign node159 = (inp[7]) ? node167 : node160;
									assign node160 = (inp[1]) ? node164 : node161;
										assign node161 = (inp[11]) ? 3'b010 : 3'b110;
										assign node164 = (inp[11]) ? 3'b110 : 3'b001;
									assign node167 = (inp[1]) ? node171 : node168;
										assign node168 = (inp[8]) ? 3'b001 : 3'b110;
										assign node171 = (inp[8]) ? 3'b001 : 3'b001;
							assign node174 = (inp[5]) ? node190 : node175;
								assign node175 = (inp[7]) ? node183 : node176;
									assign node176 = (inp[8]) ? node180 : node177;
										assign node177 = (inp[1]) ? 3'b110 : 3'b010;
										assign node180 = (inp[11]) ? 3'b110 : 3'b000;
									assign node183 = (inp[1]) ? node187 : node184;
										assign node184 = (inp[8]) ? 3'b001 : 3'b110;
										assign node187 = (inp[2]) ? 3'b001 : 3'b001;
								assign node190 = (inp[11]) ? node198 : node191;
									assign node191 = (inp[7]) ? node195 : node192;
										assign node192 = (inp[1]) ? 3'b010 : 3'b010;
										assign node195 = (inp[1]) ? 3'b110 : 3'b010;
									assign node198 = (inp[2]) ? node202 : node199;
										assign node199 = (inp[1]) ? 3'b010 : 3'b010;
										assign node202 = (inp[1]) ? 3'b010 : 3'b010;
						assign node205 = (inp[5]) ? node235 : node206;
							assign node206 = (inp[1]) ? node220 : node207;
								assign node207 = (inp[7]) ? node213 : node208;
									assign node208 = (inp[10]) ? node210 : 3'b101;
										assign node210 = (inp[8]) ? 3'b001 : 3'b000;
									assign node213 = (inp[10]) ? node217 : node214;
										assign node214 = (inp[2]) ? 3'b011 : 3'b011;
										assign node217 = (inp[8]) ? 3'b001 : 3'b101;
								assign node220 = (inp[10]) ? node228 : node221;
									assign node221 = (inp[7]) ? node225 : node222;
										assign node222 = (inp[8]) ? 3'b011 : 3'b011;
										assign node225 = (inp[11]) ? 3'b011 : 3'b111;
									assign node228 = (inp[7]) ? node232 : node229;
										assign node229 = (inp[11]) ? 3'b001 : 3'b101;
										assign node232 = (inp[11]) ? 3'b101 : 3'b011;
							assign node235 = (inp[7]) ? node251 : node236;
								assign node236 = (inp[10]) ? node244 : node237;
									assign node237 = (inp[1]) ? node241 : node238;
										assign node238 = (inp[8]) ? 3'b001 : 3'b000;
										assign node241 = (inp[2]) ? 3'b101 : 3'b101;
									assign node244 = (inp[1]) ? node248 : node245;
										assign node245 = (inp[11]) ? 3'b110 : 3'b110;
										assign node248 = (inp[2]) ? 3'b000 : 3'b001;
								assign node251 = (inp[10]) ? node259 : node252;
									assign node252 = (inp[1]) ? node256 : node253;
										assign node253 = (inp[8]) ? 3'b101 : 3'b101;
										assign node256 = (inp[8]) ? 3'b011 : 3'b101;
									assign node259 = (inp[1]) ? node263 : node260;
										assign node260 = (inp[2]) ? 3'b001 : 3'b001;
										assign node263 = (inp[11]) ? 3'b001 : 3'b101;
					assign node266 = (inp[0]) ? node326 : node267;
						assign node267 = (inp[1]) ? node297 : node268;
							assign node268 = (inp[2]) ? node282 : node269;
								assign node269 = (inp[5]) ? node277 : node270;
									assign node270 = (inp[10]) ? node274 : node271;
										assign node271 = (inp[8]) ? 3'b111 : 3'b101;
										assign node274 = (inp[7]) ? 3'b101 : 3'b001;
									assign node277 = (inp[8]) ? node279 : 3'b001;
										assign node279 = (inp[10]) ? 3'b001 : 3'b101;
								assign node282 = (inp[10]) ? node290 : node283;
									assign node283 = (inp[7]) ? node287 : node284;
										assign node284 = (inp[8]) ? 3'b001 : 3'b101;
										assign node287 = (inp[5]) ? 3'b101 : 3'b011;
									assign node290 = (inp[7]) ? node294 : node291;
										assign node291 = (inp[5]) ? 3'b110 : 3'b001;
										assign node294 = (inp[5]) ? 3'b001 : 3'b101;
							assign node297 = (inp[5]) ? node311 : node298;
								assign node298 = (inp[2]) ? node306 : node299;
									assign node299 = (inp[7]) ? node303 : node300;
										assign node300 = (inp[10]) ? 3'b101 : 3'b011;
										assign node303 = (inp[10]) ? 3'b011 : 3'b111;
									assign node306 = (inp[8]) ? node308 : 3'b011;
										assign node308 = (inp[11]) ? 3'b011 : 3'b111;
								assign node311 = (inp[10]) ? node319 : node312;
									assign node312 = (inp[7]) ? node316 : node313;
										assign node313 = (inp[11]) ? 3'b101 : 3'b101;
										assign node316 = (inp[11]) ? 3'b011 : 3'b011;
									assign node319 = (inp[7]) ? node323 : node320;
										assign node320 = (inp[11]) ? 3'b000 : 3'b001;
										assign node323 = (inp[8]) ? 3'b101 : 3'b001;
						assign node326 = (inp[10]) ? node348 : node327;
							assign node327 = (inp[5]) ? node335 : node328;
								assign node328 = (inp[7]) ? 3'b111 : node329;
									assign node329 = (inp[8]) ? 3'b111 : node330;
										assign node330 = (inp[1]) ? 3'b111 : 3'b011;
								assign node335 = (inp[7]) ? node343 : node336;
									assign node336 = (inp[1]) ? node340 : node337;
										assign node337 = (inp[8]) ? 3'b011 : 3'b011;
										assign node340 = (inp[8]) ? 3'b111 : 3'b011;
									assign node343 = (inp[11]) ? node345 : 3'b111;
										assign node345 = (inp[1]) ? 3'b111 : 3'b011;
							assign node348 = (inp[5]) ? node362 : node349;
								assign node349 = (inp[7]) ? node357 : node350;
									assign node350 = (inp[1]) ? node354 : node351;
										assign node351 = (inp[11]) ? 3'b101 : 3'b011;
										assign node354 = (inp[11]) ? 3'b011 : 3'b111;
									assign node357 = (inp[1]) ? 3'b111 : node358;
										assign node358 = (inp[2]) ? 3'b111 : 3'b011;
								assign node362 = (inp[7]) ? node370 : node363;
									assign node363 = (inp[1]) ? node367 : node364;
										assign node364 = (inp[11]) ? 3'b001 : 3'b101;
										assign node367 = (inp[8]) ? 3'b011 : 3'b101;
									assign node370 = (inp[1]) ? node374 : node371;
										assign node371 = (inp[8]) ? 3'b011 : 3'b101;
										assign node374 = (inp[11]) ? 3'b011 : 3'b111;
			assign node377 = (inp[4]) ? node613 : node378;
				assign node378 = (inp[6]) ? node502 : node379;
					assign node379 = (inp[0]) ? node439 : node380;
						assign node380 = (inp[10]) ? node410 : node381;
							assign node381 = (inp[5]) ? node395 : node382;
								assign node382 = (inp[7]) ? node388 : node383;
									assign node383 = (inp[11]) ? 3'b001 : node384;
										assign node384 = (inp[2]) ? 3'b001 : 3'b000;
									assign node388 = (inp[1]) ? node392 : node389;
										assign node389 = (inp[8]) ? 3'b101 : 3'b001;
										assign node392 = (inp[2]) ? 3'b101 : 3'b101;
								assign node395 = (inp[11]) ? node403 : node396;
									assign node396 = (inp[7]) ? node400 : node397;
										assign node397 = (inp[1]) ? 3'b001 : 3'b110;
										assign node400 = (inp[8]) ? 3'b001 : 3'b001;
									assign node403 = (inp[7]) ? node407 : node404;
										assign node404 = (inp[2]) ? 3'b110 : 3'b010;
										assign node407 = (inp[8]) ? 3'b001 : 3'b110;
							assign node410 = (inp[5]) ? node426 : node411;
								assign node411 = (inp[1]) ? node419 : node412;
									assign node412 = (inp[11]) ? node416 : node413;
										assign node413 = (inp[7]) ? 3'b001 : 3'b110;
										assign node416 = (inp[7]) ? 3'b110 : 3'b010;
									assign node419 = (inp[11]) ? node423 : node420;
										assign node420 = (inp[8]) ? 3'b001 : 3'b001;
										assign node423 = (inp[7]) ? 3'b001 : 3'b110;
								assign node426 = (inp[7]) ? node432 : node427;
									assign node427 = (inp[1]) ? 3'b010 : node428;
										assign node428 = (inp[2]) ? 3'b010 : 3'b100;
									assign node432 = (inp[11]) ? node436 : node433;
										assign node433 = (inp[2]) ? 3'b110 : 3'b110;
										assign node436 = (inp[1]) ? 3'b110 : 3'b010;
						assign node439 = (inp[10]) ? node471 : node440;
							assign node440 = (inp[5]) ? node456 : node441;
								assign node441 = (inp[7]) ? node449 : node442;
									assign node442 = (inp[1]) ? node446 : node443;
										assign node443 = (inp[2]) ? 3'b001 : 3'b101;
										assign node446 = (inp[8]) ? 3'b011 : 3'b011;
									assign node449 = (inp[8]) ? node453 : node450;
										assign node450 = (inp[1]) ? 3'b011 : 3'b011;
										assign node453 = (inp[1]) ? 3'b111 : 3'b011;
								assign node456 = (inp[11]) ? node464 : node457;
									assign node457 = (inp[7]) ? node461 : node458;
										assign node458 = (inp[1]) ? 3'b101 : 3'b001;
										assign node461 = (inp[2]) ? 3'b011 : 3'b101;
									assign node464 = (inp[7]) ? node468 : node465;
										assign node465 = (inp[1]) ? 3'b101 : 3'b001;
										assign node468 = (inp[2]) ? 3'b101 : 3'b101;
							assign node471 = (inp[5]) ? node487 : node472;
								assign node472 = (inp[1]) ? node480 : node473;
									assign node473 = (inp[8]) ? node477 : node474;
										assign node474 = (inp[7]) ? 3'b101 : 3'b001;
										assign node477 = (inp[7]) ? 3'b011 : 3'b001;
									assign node480 = (inp[2]) ? node484 : node481;
										assign node481 = (inp[8]) ? 3'b101 : 3'b101;
										assign node484 = (inp[7]) ? 3'b011 : 3'b101;
								assign node487 = (inp[7]) ? node495 : node488;
									assign node488 = (inp[11]) ? node492 : node489;
										assign node489 = (inp[1]) ? 3'b001 : 3'b110;
										assign node492 = (inp[8]) ? 3'b110 : 3'b110;
									assign node495 = (inp[1]) ? node499 : node496;
										assign node496 = (inp[8]) ? 3'b001 : 3'b000;
										assign node499 = (inp[2]) ? 3'b101 : 3'b001;
					assign node502 = (inp[0]) ? node562 : node503;
						assign node503 = (inp[10]) ? node535 : node504;
							assign node504 = (inp[5]) ? node520 : node505;
								assign node505 = (inp[11]) ? node513 : node506;
									assign node506 = (inp[7]) ? node510 : node507;
										assign node507 = (inp[2]) ? 3'b011 : 3'b011;
										assign node510 = (inp[1]) ? 3'b111 : 3'b011;
									assign node513 = (inp[1]) ? node517 : node514;
										assign node514 = (inp[7]) ? 3'b011 : 3'b101;
										assign node517 = (inp[7]) ? 3'b111 : 3'b011;
								assign node520 = (inp[2]) ? node528 : node521;
									assign node521 = (inp[11]) ? node525 : node522;
										assign node522 = (inp[8]) ? 3'b101 : 3'b001;
										assign node525 = (inp[1]) ? 3'b001 : 3'b001;
									assign node528 = (inp[7]) ? node532 : node529;
										assign node529 = (inp[1]) ? 3'b101 : 3'b001;
										assign node532 = (inp[1]) ? 3'b011 : 3'b001;
							assign node535 = (inp[1]) ? node549 : node536;
								assign node536 = (inp[5]) ? node542 : node537;
									assign node537 = (inp[7]) ? node539 : 3'b001;
										assign node539 = (inp[2]) ? 3'b101 : 3'b101;
									assign node542 = (inp[7]) ? node546 : node543;
										assign node543 = (inp[8]) ? 3'b110 : 3'b110;
										assign node546 = (inp[8]) ? 3'b001 : 3'b001;
								assign node549 = (inp[5]) ? node555 : node550;
									assign node550 = (inp[7]) ? 3'b011 : node551;
										assign node551 = (inp[2]) ? 3'b101 : 3'b101;
									assign node555 = (inp[11]) ? node559 : node556;
										assign node556 = (inp[7]) ? 3'b101 : 3'b001;
										assign node559 = (inp[7]) ? 3'b001 : 3'b001;
						assign node562 = (inp[10]) ? node584 : node563;
							assign node563 = (inp[5]) ? node571 : node564;
								assign node564 = (inp[11]) ? node566 : 3'b111;
									assign node566 = (inp[7]) ? 3'b111 : node567;
										assign node567 = (inp[8]) ? 3'b111 : 3'b111;
								assign node571 = (inp[1]) ? node579 : node572;
									assign node572 = (inp[11]) ? node576 : node573;
										assign node573 = (inp[7]) ? 3'b111 : 3'b011;
										assign node576 = (inp[7]) ? 3'b011 : 3'b101;
									assign node579 = (inp[7]) ? 3'b111 : node580;
										assign node580 = (inp[2]) ? 3'b111 : 3'b011;
							assign node584 = (inp[5]) ? node598 : node585;
								assign node585 = (inp[7]) ? node593 : node586;
									assign node586 = (inp[11]) ? node590 : node587;
										assign node587 = (inp[1]) ? 3'b111 : 3'b011;
										assign node590 = (inp[1]) ? 3'b011 : 3'b101;
									assign node593 = (inp[8]) ? 3'b111 : node594;
										assign node594 = (inp[11]) ? 3'b011 : 3'b111;
								assign node598 = (inp[1]) ? node606 : node599;
									assign node599 = (inp[11]) ? node603 : node600;
										assign node600 = (inp[7]) ? 3'b001 : 3'b101;
										assign node603 = (inp[2]) ? 3'b001 : 3'b101;
									assign node606 = (inp[2]) ? node610 : node607;
										assign node607 = (inp[7]) ? 3'b011 : 3'b101;
										assign node610 = (inp[11]) ? 3'b011 : 3'b011;
				assign node613 = (inp[6]) ? node737 : node614;
					assign node614 = (inp[0]) ? node674 : node615;
						assign node615 = (inp[5]) ? node647 : node616;
							assign node616 = (inp[10]) ? node632 : node617;
								assign node617 = (inp[7]) ? node625 : node618;
									assign node618 = (inp[1]) ? node622 : node619;
										assign node619 = (inp[2]) ? 3'b010 : 3'b100;
										assign node622 = (inp[8]) ? 3'b010 : 3'b010;
									assign node625 = (inp[1]) ? node629 : node626;
										assign node626 = (inp[11]) ? 3'b010 : 3'b110;
										assign node629 = (inp[11]) ? 3'b110 : 3'b110;
								assign node632 = (inp[7]) ? node640 : node633;
									assign node633 = (inp[11]) ? node637 : node634;
										assign node634 = (inp[8]) ? 3'b000 : 3'b100;
										assign node637 = (inp[2]) ? 3'b100 : 3'b000;
									assign node640 = (inp[1]) ? node644 : node641;
										assign node641 = (inp[11]) ? 3'b100 : 3'b010;
										assign node644 = (inp[2]) ? 3'b010 : 3'b010;
							assign node647 = (inp[10]) ? node661 : node648;
								assign node648 = (inp[7]) ? node654 : node649;
									assign node649 = (inp[1]) ? 3'b100 : node650;
										assign node650 = (inp[2]) ? 3'b100 : 3'b000;
									assign node654 = (inp[11]) ? node658 : node655;
										assign node655 = (inp[8]) ? 3'b010 : 3'b010;
										assign node658 = (inp[1]) ? 3'b010 : 3'b100;
								assign node661 = (inp[1]) ? node667 : node662;
									assign node662 = (inp[11]) ? 3'b000 : node663;
										assign node663 = (inp[8]) ? 3'b100 : 3'b000;
									assign node667 = (inp[7]) ? node671 : node668;
										assign node668 = (inp[11]) ? 3'b000 : 3'b000;
										assign node671 = (inp[11]) ? 3'b100 : 3'b100;
						assign node674 = (inp[10]) ? node706 : node675;
							assign node675 = (inp[5]) ? node691 : node676;
								assign node676 = (inp[7]) ? node684 : node677;
									assign node677 = (inp[11]) ? node681 : node678;
										assign node678 = (inp[1]) ? 3'b001 : 3'b110;
										assign node681 = (inp[8]) ? 3'b110 : 3'b110;
									assign node684 = (inp[1]) ? node688 : node685;
										assign node685 = (inp[11]) ? 3'b001 : 3'b001;
										assign node688 = (inp[8]) ? 3'b101 : 3'b001;
								assign node691 = (inp[7]) ? node699 : node692;
									assign node692 = (inp[2]) ? node696 : node693;
										assign node693 = (inp[8]) ? 3'b010 : 3'b010;
										assign node696 = (inp[11]) ? 3'b010 : 3'b110;
									assign node699 = (inp[1]) ? node703 : node700;
										assign node700 = (inp[8]) ? 3'b110 : 3'b010;
										assign node703 = (inp[8]) ? 3'b001 : 3'b110;
							assign node706 = (inp[5]) ? node722 : node707;
								assign node707 = (inp[7]) ? node715 : node708;
									assign node708 = (inp[1]) ? node712 : node709;
										assign node709 = (inp[11]) ? 3'b000 : 3'b010;
										assign node712 = (inp[11]) ? 3'b010 : 3'b110;
									assign node715 = (inp[1]) ? node719 : node716;
										assign node716 = (inp[11]) ? 3'b010 : 3'b110;
										assign node719 = (inp[11]) ? 3'b110 : 3'b001;
								assign node722 = (inp[7]) ? node730 : node723;
									assign node723 = (inp[1]) ? node727 : node724;
										assign node724 = (inp[8]) ? 3'b100 : 3'b100;
										assign node727 = (inp[11]) ? 3'b100 : 3'b010;
									assign node730 = (inp[1]) ? node734 : node731;
										assign node731 = (inp[11]) ? 3'b100 : 3'b010;
										assign node734 = (inp[2]) ? 3'b110 : 3'b010;
					assign node737 = (inp[0]) ? node797 : node738;
						assign node738 = (inp[10]) ? node770 : node739;
							assign node739 = (inp[5]) ? node755 : node740;
								assign node740 = (inp[7]) ? node748 : node741;
									assign node741 = (inp[1]) ? node745 : node742;
										assign node742 = (inp[2]) ? 3'b110 : 3'b110;
										assign node745 = (inp[8]) ? 3'b001 : 3'b001;
									assign node748 = (inp[11]) ? node752 : node749;
										assign node749 = (inp[1]) ? 3'b101 : 3'b001;
										assign node752 = (inp[2]) ? 3'b001 : 3'b001;
								assign node755 = (inp[1]) ? node763 : node756;
									assign node756 = (inp[7]) ? node760 : node757;
										assign node757 = (inp[8]) ? 3'b010 : 3'b000;
										assign node760 = (inp[8]) ? 3'b110 : 3'b010;
									assign node763 = (inp[7]) ? node767 : node764;
										assign node764 = (inp[8]) ? 3'b110 : 3'b110;
										assign node767 = (inp[11]) ? 3'b110 : 3'b001;
							assign node770 = (inp[7]) ? node782 : node771;
								assign node771 = (inp[5]) ? node777 : node772;
									assign node772 = (inp[8]) ? 3'b110 : node773;
										assign node773 = (inp[2]) ? 3'b010 : 3'b110;
									assign node777 = (inp[1]) ? node779 : 3'b100;
										assign node779 = (inp[11]) ? 3'b100 : 3'b010;
								assign node782 = (inp[5]) ? node790 : node783;
									assign node783 = (inp[11]) ? node787 : node784;
										assign node784 = (inp[1]) ? 3'b001 : 3'b110;
										assign node787 = (inp[2]) ? 3'b110 : 3'b110;
									assign node790 = (inp[1]) ? node794 : node791;
										assign node791 = (inp[2]) ? 3'b010 : 3'b010;
										assign node794 = (inp[2]) ? 3'b110 : 3'b010;
						assign node797 = (inp[11]) ? node827 : node798;
							assign node798 = (inp[5]) ? node812 : node799;
								assign node799 = (inp[1]) ? node805 : node800;
									assign node800 = (inp[10]) ? node802 : 3'b101;
										assign node802 = (inp[7]) ? 3'b101 : 3'b001;
									assign node805 = (inp[10]) ? node809 : node806;
										assign node806 = (inp[7]) ? 3'b111 : 3'b011;
										assign node809 = (inp[2]) ? 3'b101 : 3'b101;
								assign node812 = (inp[10]) ? node820 : node813;
									assign node813 = (inp[8]) ? node817 : node814;
										assign node814 = (inp[7]) ? 3'b101 : 3'b001;
										assign node817 = (inp[7]) ? 3'b011 : 3'b001;
									assign node820 = (inp[2]) ? node824 : node821;
										assign node821 = (inp[8]) ? 3'b001 : 3'b010;
										assign node824 = (inp[8]) ? 3'b001 : 3'b001;
							assign node827 = (inp[5]) ? node843 : node828;
								assign node828 = (inp[10]) ? node836 : node829;
									assign node829 = (inp[1]) ? node833 : node830;
										assign node830 = (inp[7]) ? 3'b101 : 3'b001;
										assign node833 = (inp[7]) ? 3'b011 : 3'b101;
									assign node836 = (inp[7]) ? node840 : node837;
										assign node837 = (inp[1]) ? 3'b001 : 3'b110;
										assign node840 = (inp[2]) ? 3'b101 : 3'b001;
								assign node843 = (inp[7]) ? node851 : node844;
									assign node844 = (inp[10]) ? node848 : node845;
										assign node845 = (inp[1]) ? 3'b001 : 3'b110;
										assign node848 = (inp[1]) ? 3'b110 : 3'b010;
									assign node851 = (inp[10]) ? node855 : node852;
										assign node852 = (inp[1]) ? 3'b101 : 3'b001;
										assign node855 = (inp[1]) ? 3'b001 : 3'b110;
		assign node858 = (inp[9]) ? node1304 : node859;
			assign node859 = (inp[4]) ? node1101 : node860;
				assign node860 = (inp[6]) ? node978 : node861;
					assign node861 = (inp[0]) ? node917 : node862;
						assign node862 = (inp[10]) ? node894 : node863;
							assign node863 = (inp[5]) ? node879 : node864;
								assign node864 = (inp[7]) ? node872 : node865;
									assign node865 = (inp[1]) ? node869 : node866;
										assign node866 = (inp[2]) ? 3'b010 : 3'b100;
										assign node869 = (inp[11]) ? 3'b010 : 3'b110;
									assign node872 = (inp[2]) ? node876 : node873;
										assign node873 = (inp[1]) ? 3'b110 : 3'b010;
										assign node876 = (inp[1]) ? 3'b110 : 3'b110;
								assign node879 = (inp[11]) ? node887 : node880;
									assign node880 = (inp[1]) ? node884 : node881;
										assign node881 = (inp[7]) ? 3'b010 : 3'b100;
										assign node884 = (inp[7]) ? 3'b010 : 3'b010;
									assign node887 = (inp[1]) ? node891 : node888;
										assign node888 = (inp[7]) ? 3'b100 : 3'b000;
										assign node891 = (inp[7]) ? 3'b000 : 3'b100;
							assign node894 = (inp[5]) ? node908 : node895;
								assign node895 = (inp[11]) ? node903 : node896;
									assign node896 = (inp[1]) ? node900 : node897;
										assign node897 = (inp[2]) ? 3'b100 : 3'b000;
										assign node900 = (inp[2]) ? 3'b010 : 3'b010;
									assign node903 = (inp[7]) ? 3'b100 : node904;
										assign node904 = (inp[1]) ? 3'b100 : 3'b000;
								assign node908 = (inp[7]) ? node910 : 3'b000;
									assign node910 = (inp[1]) ? node914 : node911;
										assign node911 = (inp[11]) ? 3'b000 : 3'b100;
										assign node914 = (inp[11]) ? 3'b100 : 3'b100;
						assign node917 = (inp[10]) ? node947 : node918;
							assign node918 = (inp[5]) ? node932 : node919;
								assign node919 = (inp[1]) ? node927 : node920;
									assign node920 = (inp[7]) ? node924 : node921;
										assign node921 = (inp[8]) ? 3'b110 : 3'b110;
										assign node924 = (inp[2]) ? 3'b001 : 3'b001;
									assign node927 = (inp[11]) ? 3'b001 : node928;
										assign node928 = (inp[7]) ? 3'b101 : 3'b001;
								assign node932 = (inp[7]) ? node940 : node933;
									assign node933 = (inp[1]) ? node937 : node934;
										assign node934 = (inp[2]) ? 3'b010 : 3'b000;
										assign node937 = (inp[2]) ? 3'b110 : 3'b010;
									assign node940 = (inp[2]) ? node944 : node941;
										assign node941 = (inp[1]) ? 3'b110 : 3'b110;
										assign node944 = (inp[1]) ? 3'b001 : 3'b110;
							assign node947 = (inp[5]) ? node963 : node948;
								assign node948 = (inp[7]) ? node956 : node949;
									assign node949 = (inp[1]) ? node953 : node950;
										assign node950 = (inp[11]) ? 3'b010 : 3'b010;
										assign node953 = (inp[11]) ? 3'b010 : 3'b110;
									assign node956 = (inp[1]) ? node960 : node957;
										assign node957 = (inp[8]) ? 3'b110 : 3'b110;
										assign node960 = (inp[8]) ? 3'b001 : 3'b110;
								assign node963 = (inp[11]) ? node971 : node964;
									assign node964 = (inp[8]) ? node968 : node965;
										assign node965 = (inp[7]) ? 3'b010 : 3'b000;
										assign node968 = (inp[1]) ? 3'b010 : 3'b010;
									assign node971 = (inp[1]) ? node975 : node972;
										assign node972 = (inp[8]) ? 3'b100 : 3'b100;
										assign node975 = (inp[7]) ? 3'b010 : 3'b100;
					assign node978 = (inp[0]) ? node1040 : node979;
						assign node979 = (inp[10]) ? node1009 : node980;
							assign node980 = (inp[1]) ? node994 : node981;
								assign node981 = (inp[5]) ? node987 : node982;
									assign node982 = (inp[11]) ? node984 : 3'b001;
										assign node984 = (inp[7]) ? 3'b000 : 3'b110;
									assign node987 = (inp[7]) ? node991 : node988;
										assign node988 = (inp[8]) ? 3'b010 : 3'b010;
										assign node991 = (inp[2]) ? 3'b110 : 3'b110;
								assign node994 = (inp[11]) ? node1002 : node995;
									assign node995 = (inp[8]) ? node999 : node996;
										assign node996 = (inp[5]) ? 3'b001 : 3'b001;
										assign node999 = (inp[7]) ? 3'b001 : 3'b101;
									assign node1002 = (inp[8]) ? node1006 : node1003;
										assign node1003 = (inp[5]) ? 3'b110 : 3'b100;
										assign node1006 = (inp[5]) ? 3'b000 : 3'b001;
							assign node1009 = (inp[5]) ? node1025 : node1010;
								assign node1010 = (inp[7]) ? node1018 : node1011;
									assign node1011 = (inp[1]) ? node1015 : node1012;
										assign node1012 = (inp[8]) ? 3'b010 : 3'b000;
										assign node1015 = (inp[2]) ? 3'b110 : 3'b110;
									assign node1018 = (inp[11]) ? node1022 : node1019;
										assign node1019 = (inp[1]) ? 3'b001 : 3'b000;
										assign node1022 = (inp[8]) ? 3'b110 : 3'b110;
								assign node1025 = (inp[7]) ? node1033 : node1026;
									assign node1026 = (inp[1]) ? node1030 : node1027;
										assign node1027 = (inp[2]) ? 3'b100 : 3'b100;
										assign node1030 = (inp[11]) ? 3'b010 : 3'b010;
									assign node1033 = (inp[11]) ? node1037 : node1034;
										assign node1034 = (inp[1]) ? 3'b110 : 3'b010;
										assign node1037 = (inp[2]) ? 3'b010 : 3'b010;
						assign node1040 = (inp[7]) ? node1072 : node1041;
							assign node1041 = (inp[5]) ? node1057 : node1042;
								assign node1042 = (inp[10]) ? node1050 : node1043;
									assign node1043 = (inp[1]) ? node1047 : node1044;
										assign node1044 = (inp[11]) ? 3'b101 : 3'b101;
										assign node1047 = (inp[11]) ? 3'b101 : 3'b001;
									assign node1050 = (inp[11]) ? node1054 : node1051;
										assign node1051 = (inp[1]) ? 3'b101 : 3'b001;
										assign node1054 = (inp[1]) ? 3'b001 : 3'b110;
								assign node1057 = (inp[10]) ? node1065 : node1058;
									assign node1058 = (inp[11]) ? node1062 : node1059;
										assign node1059 = (inp[1]) ? 3'b001 : 3'b001;
										assign node1062 = (inp[8]) ? 3'b001 : 3'b110;
									assign node1065 = (inp[11]) ? node1069 : node1066;
										assign node1066 = (inp[1]) ? 3'b001 : 3'b110;
										assign node1069 = (inp[1]) ? 3'b110 : 3'b010;
							assign node1072 = (inp[1]) ? node1088 : node1073;
								assign node1073 = (inp[5]) ? node1081 : node1074;
									assign node1074 = (inp[2]) ? node1078 : node1075;
										assign node1075 = (inp[10]) ? 3'b001 : 3'b101;
										assign node1078 = (inp[10]) ? 3'b101 : 3'b011;
									assign node1081 = (inp[8]) ? node1085 : node1082;
										assign node1082 = (inp[10]) ? 3'b110 : 3'b001;
										assign node1085 = (inp[10]) ? 3'b001 : 3'b101;
								assign node1088 = (inp[5]) ? node1096 : node1089;
									assign node1089 = (inp[10]) ? node1093 : node1090;
										assign node1090 = (inp[11]) ? 3'b011 : 3'b111;
										assign node1093 = (inp[11]) ? 3'b101 : 3'b011;
									assign node1096 = (inp[10]) ? 3'b001 : node1097;
										assign node1097 = (inp[11]) ? 3'b101 : 3'b011;
				assign node1101 = (inp[6]) ? node1187 : node1102;
					assign node1102 = (inp[0]) ? node1134 : node1103;
						assign node1103 = (inp[10]) ? node1125 : node1104;
							assign node1104 = (inp[5]) ? node1118 : node1105;
								assign node1105 = (inp[7]) ? node1111 : node1106;
									assign node1106 = (inp[8]) ? node1108 : 3'b000;
										assign node1108 = (inp[2]) ? 3'b000 : 3'b000;
									assign node1111 = (inp[11]) ? node1115 : node1112;
										assign node1112 = (inp[1]) ? 3'b100 : 3'b100;
										assign node1115 = (inp[1]) ? 3'b100 : 3'b000;
								assign node1118 = (inp[11]) ? 3'b000 : node1119;
									assign node1119 = (inp[7]) ? node1121 : 3'b000;
										assign node1121 = (inp[1]) ? 3'b000 : 3'b000;
							assign node1125 = (inp[1]) ? node1127 : 3'b000;
								assign node1127 = (inp[8]) ? node1129 : 3'b000;
									assign node1129 = (inp[11]) ? 3'b000 : node1130;
										assign node1130 = (inp[7]) ? 3'b000 : 3'b000;
						assign node1134 = (inp[10]) ? node1166 : node1135;
							assign node1135 = (inp[5]) ? node1151 : node1136;
								assign node1136 = (inp[7]) ? node1144 : node1137;
									assign node1137 = (inp[11]) ? node1141 : node1138;
										assign node1138 = (inp[1]) ? 3'b010 : 3'b100;
										assign node1141 = (inp[8]) ? 3'b000 : 3'b100;
									assign node1144 = (inp[1]) ? node1148 : node1145;
										assign node1145 = (inp[8]) ? 3'b010 : 3'b000;
										assign node1148 = (inp[11]) ? 3'b010 : 3'b110;
								assign node1151 = (inp[7]) ? node1159 : node1152;
									assign node1152 = (inp[1]) ? node1156 : node1153;
										assign node1153 = (inp[8]) ? 3'b000 : 3'b000;
										assign node1156 = (inp[11]) ? 3'b000 : 3'b100;
									assign node1159 = (inp[1]) ? node1163 : node1160;
										assign node1160 = (inp[11]) ? 3'b000 : 3'b100;
										assign node1163 = (inp[8]) ? 3'b010 : 3'b000;
							assign node1166 = (inp[5]) ? node1180 : node1167;
								assign node1167 = (inp[7]) ? node1173 : node1168;
									assign node1168 = (inp[8]) ? node1170 : 3'b000;
										assign node1170 = (inp[2]) ? 3'b100 : 3'b000;
									assign node1173 = (inp[2]) ? node1177 : node1174;
										assign node1174 = (inp[1]) ? 3'b100 : 3'b000;
										assign node1177 = (inp[1]) ? 3'b010 : 3'b100;
								assign node1180 = (inp[1]) ? node1182 : 3'b000;
									assign node1182 = (inp[7]) ? node1184 : 3'b000;
										assign node1184 = (inp[8]) ? 3'b100 : 3'b000;
					assign node1187 = (inp[0]) ? node1243 : node1188;
						assign node1188 = (inp[5]) ? node1220 : node1189;
							assign node1189 = (inp[10]) ? node1205 : node1190;
								assign node1190 = (inp[1]) ? node1198 : node1191;
									assign node1191 = (inp[7]) ? node1195 : node1192;
										assign node1192 = (inp[2]) ? 3'b100 : 3'b000;
										assign node1195 = (inp[8]) ? 3'b010 : 3'b010;
									assign node1198 = (inp[7]) ? node1202 : node1199;
										assign node1199 = (inp[2]) ? 3'b010 : 3'b010;
										assign node1202 = (inp[11]) ? 3'b010 : 3'b110;
								assign node1205 = (inp[2]) ? node1213 : node1206;
									assign node1206 = (inp[11]) ? node1210 : node1207;
										assign node1207 = (inp[1]) ? 3'b100 : 3'b100;
										assign node1210 = (inp[7]) ? 3'b100 : 3'b000;
									assign node1213 = (inp[7]) ? node1217 : node1214;
										assign node1214 = (inp[8]) ? 3'b100 : 3'b000;
										assign node1217 = (inp[1]) ? 3'b010 : 3'b100;
							assign node1220 = (inp[10]) ? node1236 : node1221;
								assign node1221 = (inp[11]) ? node1229 : node1222;
									assign node1222 = (inp[7]) ? node1226 : node1223;
										assign node1223 = (inp[1]) ? 3'b100 : 3'b000;
										assign node1226 = (inp[1]) ? 3'b010 : 3'b100;
									assign node1229 = (inp[1]) ? node1233 : node1230;
										assign node1230 = (inp[7]) ? 3'b100 : 3'b000;
										assign node1233 = (inp[8]) ? 3'b100 : 3'b100;
								assign node1236 = (inp[7]) ? node1238 : 3'b000;
									assign node1238 = (inp[1]) ? node1240 : 3'b000;
										assign node1240 = (inp[11]) ? 3'b000 : 3'b100;
						assign node1243 = (inp[5]) ? node1275 : node1244;
							assign node1244 = (inp[10]) ? node1260 : node1245;
								assign node1245 = (inp[7]) ? node1253 : node1246;
									assign node1246 = (inp[1]) ? node1250 : node1247;
										assign node1247 = (inp[11]) ? 3'b010 : 3'b110;
										assign node1250 = (inp[8]) ? 3'b001 : 3'b110;
									assign node1253 = (inp[1]) ? node1257 : node1254;
										assign node1254 = (inp[2]) ? 3'b001 : 3'b110;
										assign node1257 = (inp[11]) ? 3'b001 : 3'b001;
								assign node1260 = (inp[11]) ? node1268 : node1261;
									assign node1261 = (inp[1]) ? node1265 : node1262;
										assign node1262 = (inp[7]) ? 3'b110 : 3'b000;
										assign node1265 = (inp[7]) ? 3'b110 : 3'b110;
									assign node1268 = (inp[8]) ? node1272 : node1269;
										assign node1269 = (inp[2]) ? 3'b100 : 3'b010;
										assign node1272 = (inp[7]) ? 3'b010 : 3'b010;
							assign node1275 = (inp[7]) ? node1291 : node1276;
								assign node1276 = (inp[10]) ? node1284 : node1277;
									assign node1277 = (inp[1]) ? node1281 : node1278;
										assign node1278 = (inp[8]) ? 3'b010 : 3'b100;
										assign node1281 = (inp[11]) ? 3'b010 : 3'b110;
									assign node1284 = (inp[8]) ? node1288 : node1285;
										assign node1285 = (inp[1]) ? 3'b100 : 3'b000;
										assign node1288 = (inp[11]) ? 3'b100 : 3'b100;
								assign node1291 = (inp[10]) ? node1297 : node1292;
									assign node1292 = (inp[2]) ? 3'b110 : node1293;
										assign node1293 = (inp[8]) ? 3'b110 : 3'b010;
									assign node1297 = (inp[11]) ? node1301 : node1298;
										assign node1298 = (inp[1]) ? 3'b010 : 3'b010;
										assign node1301 = (inp[1]) ? 3'b010 : 3'b100;
			assign node1304 = (inp[4]) ? node1494 : node1305;
				assign node1305 = (inp[6]) ? node1379 : node1306;
					assign node1306 = (inp[0]) ? node1330 : node1307;
						assign node1307 = (inp[10]) ? 3'b000 : node1308;
							assign node1308 = (inp[5]) ? node1322 : node1309;
								assign node1309 = (inp[7]) ? node1315 : node1310;
									assign node1310 = (inp[1]) ? node1312 : 3'b000;
										assign node1312 = (inp[8]) ? 3'b000 : 3'b000;
									assign node1315 = (inp[1]) ? node1319 : node1316;
										assign node1316 = (inp[2]) ? 3'b000 : 3'b000;
										assign node1319 = (inp[8]) ? 3'b100 : 3'b100;
								assign node1322 = (inp[11]) ? 3'b000 : node1323;
									assign node1323 = (inp[7]) ? node1325 : 3'b000;
										assign node1325 = (inp[1]) ? 3'b000 : 3'b000;
						assign node1330 = (inp[5]) ? node1360 : node1331;
							assign node1331 = (inp[10]) ? node1347 : node1332;
								assign node1332 = (inp[11]) ? node1340 : node1333;
									assign node1333 = (inp[7]) ? node1337 : node1334;
										assign node1334 = (inp[1]) ? 3'b010 : 3'b100;
										assign node1337 = (inp[1]) ? 3'b110 : 3'b010;
									assign node1340 = (inp[1]) ? node1344 : node1341;
										assign node1341 = (inp[8]) ? 3'b100 : 3'b100;
										assign node1344 = (inp[8]) ? 3'b010 : 3'b100;
								assign node1347 = (inp[7]) ? node1353 : node1348;
									assign node1348 = (inp[1]) ? node1350 : 3'b000;
										assign node1350 = (inp[2]) ? 3'b100 : 3'b000;
									assign node1353 = (inp[11]) ? node1357 : node1354;
										assign node1354 = (inp[1]) ? 3'b010 : 3'b100;
										assign node1357 = (inp[1]) ? 3'b100 : 3'b000;
							assign node1360 = (inp[7]) ? node1368 : node1361;
								assign node1361 = (inp[10]) ? 3'b000 : node1362;
									assign node1362 = (inp[8]) ? node1364 : 3'b000;
										assign node1364 = (inp[1]) ? 3'b000 : 3'b000;
								assign node1368 = (inp[10]) ? node1374 : node1369;
									assign node1369 = (inp[2]) ? 3'b010 : node1370;
										assign node1370 = (inp[8]) ? 3'b100 : 3'b100;
									assign node1374 = (inp[11]) ? 3'b000 : node1375;
										assign node1375 = (inp[1]) ? 3'b100 : 3'b000;
					assign node1379 = (inp[0]) ? node1433 : node1380;
						assign node1380 = (inp[5]) ? node1412 : node1381;
							assign node1381 = (inp[10]) ? node1397 : node1382;
								assign node1382 = (inp[7]) ? node1390 : node1383;
									assign node1383 = (inp[11]) ? node1387 : node1384;
										assign node1384 = (inp[2]) ? 3'b010 : 3'b100;
										assign node1387 = (inp[2]) ? 3'b100 : 3'b100;
									assign node1390 = (inp[2]) ? node1394 : node1391;
										assign node1391 = (inp[8]) ? 3'b010 : 3'b000;
										assign node1394 = (inp[1]) ? 3'b110 : 3'b010;
								assign node1397 = (inp[7]) ? node1405 : node1398;
									assign node1398 = (inp[8]) ? node1402 : node1399;
										assign node1399 = (inp[1]) ? 3'b000 : 3'b000;
										assign node1402 = (inp[2]) ? 3'b100 : 3'b000;
									assign node1405 = (inp[1]) ? node1409 : node1406;
										assign node1406 = (inp[8]) ? 3'b100 : 3'b100;
										assign node1409 = (inp[11]) ? 3'b100 : 3'b010;
							assign node1412 = (inp[10]) ? node1426 : node1413;
								assign node1413 = (inp[7]) ? node1419 : node1414;
									assign node1414 = (inp[1]) ? node1416 : 3'b000;
										assign node1416 = (inp[11]) ? 3'b000 : 3'b100;
									assign node1419 = (inp[1]) ? node1423 : node1420;
										assign node1420 = (inp[11]) ? 3'b000 : 3'b100;
										assign node1423 = (inp[11]) ? 3'b100 : 3'b010;
								assign node1426 = (inp[7]) ? node1428 : 3'b000;
									assign node1428 = (inp[1]) ? node1430 : 3'b000;
										assign node1430 = (inp[2]) ? 3'b100 : 3'b000;
						assign node1433 = (inp[5]) ? node1463 : node1434;
							assign node1434 = (inp[10]) ? node1448 : node1435;
								assign node1435 = (inp[7]) ? node1441 : node1436;
									assign node1436 = (inp[11]) ? 3'b110 : node1437;
										assign node1437 = (inp[1]) ? 3'b000 : 3'b110;
									assign node1441 = (inp[8]) ? node1445 : node1442;
										assign node1442 = (inp[1]) ? 3'b001 : 3'b110;
										assign node1445 = (inp[1]) ? 3'b101 : 3'b001;
								assign node1448 = (inp[7]) ? node1456 : node1449;
									assign node1449 = (inp[1]) ? node1453 : node1450;
										assign node1450 = (inp[8]) ? 3'b010 : 3'b100;
										assign node1453 = (inp[2]) ? 3'b010 : 3'b010;
									assign node1456 = (inp[1]) ? node1460 : node1457;
										assign node1457 = (inp[11]) ? 3'b010 : 3'b110;
										assign node1460 = (inp[11]) ? 3'b110 : 3'b110;
							assign node1463 = (inp[1]) ? node1479 : node1464;
								assign node1464 = (inp[10]) ? node1472 : node1465;
									assign node1465 = (inp[8]) ? node1469 : node1466;
										assign node1466 = (inp[7]) ? 3'b110 : 3'b100;
										assign node1469 = (inp[11]) ? 3'b010 : 3'b110;
									assign node1472 = (inp[7]) ? node1476 : node1473;
										assign node1473 = (inp[11]) ? 3'b000 : 3'b100;
										assign node1476 = (inp[8]) ? 3'b000 : 3'b100;
								assign node1479 = (inp[10]) ? node1487 : node1480;
									assign node1480 = (inp[7]) ? node1484 : node1481;
										assign node1481 = (inp[11]) ? 3'b010 : 3'b010;
										assign node1484 = (inp[2]) ? 3'b110 : 3'b110;
									assign node1487 = (inp[7]) ? node1491 : node1488;
										assign node1488 = (inp[8]) ? 3'b010 : 3'b100;
										assign node1491 = (inp[11]) ? 3'b010 : 3'b010;
				assign node1494 = (inp[6]) ? node1508 : node1495;
					assign node1495 = (inp[10]) ? 3'b000 : node1496;
						assign node1496 = (inp[5]) ? 3'b000 : node1497;
							assign node1497 = (inp[11]) ? 3'b000 : node1498;
								assign node1498 = (inp[7]) ? node1500 : 3'b000;
									assign node1500 = (inp[0]) ? node1502 : 3'b000;
										assign node1502 = (inp[1]) ? 3'b100 : 3'b000;
					assign node1508 = (inp[0]) ? node1520 : node1509;
						assign node1509 = (inp[10]) ? 3'b000 : node1510;
							assign node1510 = (inp[1]) ? node1512 : 3'b000;
								assign node1512 = (inp[7]) ? node1514 : 3'b000;
									assign node1514 = (inp[5]) ? 3'b000 : node1515;
										assign node1515 = (inp[2]) ? 3'b100 : 3'b000;
						assign node1520 = (inp[10]) ? node1550 : node1521;
							assign node1521 = (inp[5]) ? node1537 : node1522;
								assign node1522 = (inp[7]) ? node1530 : node1523;
									assign node1523 = (inp[1]) ? node1527 : node1524;
										assign node1524 = (inp[11]) ? 3'b000 : 3'b100;
										assign node1527 = (inp[11]) ? 3'b100 : 3'b100;
									assign node1530 = (inp[11]) ? node1534 : node1531;
										assign node1531 = (inp[8]) ? 3'b010 : 3'b010;
										assign node1534 = (inp[1]) ? 3'b010 : 3'b100;
								assign node1537 = (inp[7]) ? node1543 : node1538;
									assign node1538 = (inp[8]) ? node1540 : 3'b000;
										assign node1540 = (inp[2]) ? 3'b000 : 3'b000;
									assign node1543 = (inp[8]) ? node1547 : node1544;
										assign node1544 = (inp[1]) ? 3'b100 : 3'b000;
										assign node1547 = (inp[2]) ? 3'b100 : 3'b100;
							assign node1550 = (inp[1]) ? node1552 : 3'b000;
								assign node1552 = (inp[7]) ? node1554 : 3'b000;
									assign node1554 = (inp[5]) ? node1558 : node1555;
										assign node1555 = (inp[2]) ? 3'b010 : 3'b100;
										assign node1558 = (inp[2]) ? 3'b000 : 3'b000;

endmodule