module dtc_split25_bm71 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node7;
	wire [3-1:0] node8;
	wire [3-1:0] node9;
	wire [3-1:0] node13;
	wire [3-1:0] node14;
	wire [3-1:0] node17;
	wire [3-1:0] node20;
	wire [3-1:0] node23;
	wire [3-1:0] node25;
	wire [3-1:0] node27;
	wire [3-1:0] node29;
	wire [3-1:0] node32;
	wire [3-1:0] node33;
	wire [3-1:0] node34;
	wire [3-1:0] node35;
	wire [3-1:0] node36;
	wire [3-1:0] node39;
	wire [3-1:0] node43;
	wire [3-1:0] node45;
	wire [3-1:0] node48;
	wire [3-1:0] node49;
	wire [3-1:0] node51;
	wire [3-1:0] node53;
	wire [3-1:0] node56;
	wire [3-1:0] node58;
	wire [3-1:0] node59;
	wire [3-1:0] node62;
	wire [3-1:0] node63;
	wire [3-1:0] node67;
	wire [3-1:0] node68;
	wire [3-1:0] node69;
	wire [3-1:0] node70;
	wire [3-1:0] node71;
	wire [3-1:0] node72;
	wire [3-1:0] node79;
	wire [3-1:0] node80;
	wire [3-1:0] node81;
	wire [3-1:0] node82;
	wire [3-1:0] node83;
	wire [3-1:0] node88;
	wire [3-1:0] node89;
	wire [3-1:0] node91;
	wire [3-1:0] node94;
	wire [3-1:0] node96;
	wire [3-1:0] node99;
	wire [3-1:0] node100;
	wire [3-1:0] node101;
	wire [3-1:0] node103;
	wire [3-1:0] node108;
	wire [3-1:0] node109;
	wire [3-1:0] node110;
	wire [3-1:0] node111;
	wire [3-1:0] node112;
	wire [3-1:0] node113;
	wire [3-1:0] node120;
	wire [3-1:0] node121;
	wire [3-1:0] node122;
	wire [3-1:0] node123;
	wire [3-1:0] node124;
	wire [3-1:0] node125;
	wire [3-1:0] node129;
	wire [3-1:0] node132;
	wire [3-1:0] node134;
	wire [3-1:0] node136;
	wire [3-1:0] node139;
	wire [3-1:0] node140;
	wire [3-1:0] node141;
	wire [3-1:0] node142;
	wire [3-1:0] node146;
	wire [3-1:0] node149;
	wire [3-1:0] node150;
	wire [3-1:0] node152;
	wire [3-1:0] node155;
	wire [3-1:0] node158;
	wire [3-1:0] node159;
	wire [3-1:0] node161;
	wire [3-1:0] node165;
	wire [3-1:0] node167;
	wire [3-1:0] node168;
	wire [3-1:0] node169;
	wire [3-1:0] node170;
	wire [3-1:0] node171;
	wire [3-1:0] node172;
	wire [3-1:0] node173;
	wire [3-1:0] node177;
	wire [3-1:0] node180;
	wire [3-1:0] node181;
	wire [3-1:0] node188;
	wire [3-1:0] node189;
	wire [3-1:0] node190;
	wire [3-1:0] node191;
	wire [3-1:0] node192;
	wire [3-1:0] node193;
	wire [3-1:0] node194;
	wire [3-1:0] node195;
	wire [3-1:0] node199;
	wire [3-1:0] node200;
	wire [3-1:0] node203;
	wire [3-1:0] node206;
	wire [3-1:0] node207;
	wire [3-1:0] node208;
	wire [3-1:0] node209;
	wire [3-1:0] node210;
	wire [3-1:0] node215;
	wire [3-1:0] node218;
	wire [3-1:0] node219;
	wire [3-1:0] node220;
	wire [3-1:0] node222;
	wire [3-1:0] node226;
	wire [3-1:0] node229;
	wire [3-1:0] node230;
	wire [3-1:0] node231;
	wire [3-1:0] node234;
	wire [3-1:0] node236;
	wire [3-1:0] node239;
	wire [3-1:0] node240;
	wire [3-1:0] node241;
	wire [3-1:0] node245;
	wire [3-1:0] node246;
	wire [3-1:0] node247;
	wire [3-1:0] node250;
	wire [3-1:0] node254;
	wire [3-1:0] node255;
	wire [3-1:0] node256;
	wire [3-1:0] node258;
	wire [3-1:0] node260;
	wire [3-1:0] node263;
	wire [3-1:0] node264;
	wire [3-1:0] node265;
	wire [3-1:0] node266;
	wire [3-1:0] node270;
	wire [3-1:0] node273;
	wire [3-1:0] node274;
	wire [3-1:0] node275;
	wire [3-1:0] node278;
	wire [3-1:0] node282;
	wire [3-1:0] node284;
	wire [3-1:0] node285;
	wire [3-1:0] node287;
	wire [3-1:0] node290;
	wire [3-1:0] node293;
	wire [3-1:0] node294;
	wire [3-1:0] node295;
	wire [3-1:0] node296;
	wire [3-1:0] node297;
	wire [3-1:0] node298;
	wire [3-1:0] node299;
	wire [3-1:0] node303;
	wire [3-1:0] node304;
	wire [3-1:0] node308;
	wire [3-1:0] node309;
	wire [3-1:0] node312;
	wire [3-1:0] node314;
	wire [3-1:0] node317;
	wire [3-1:0] node318;
	wire [3-1:0] node319;
	wire [3-1:0] node321;
	wire [3-1:0] node322;
	wire [3-1:0] node326;
	wire [3-1:0] node329;
	wire [3-1:0] node330;
	wire [3-1:0] node333;
	wire [3-1:0] node334;
	wire [3-1:0] node338;
	wire [3-1:0] node339;
	wire [3-1:0] node340;
	wire [3-1:0] node342;
	wire [3-1:0] node345;
	wire [3-1:0] node346;
	wire [3-1:0] node349;
	wire [3-1:0] node352;
	wire [3-1:0] node353;
	wire [3-1:0] node354;
	wire [3-1:0] node356;
	wire [3-1:0] node360;
	wire [3-1:0] node361;
	wire [3-1:0] node364;
	wire [3-1:0] node367;
	wire [3-1:0] node368;
	wire [3-1:0] node369;
	wire [3-1:0] node370;
	wire [3-1:0] node371;
	wire [3-1:0] node372;
	wire [3-1:0] node377;
	wire [3-1:0] node378;
	wire [3-1:0] node380;
	wire [3-1:0] node384;
	wire [3-1:0] node385;
	wire [3-1:0] node386;
	wire [3-1:0] node388;
	wire [3-1:0] node390;
	wire [3-1:0] node393;
	wire [3-1:0] node396;
	wire [3-1:0] node397;
	wire [3-1:0] node400;
	wire [3-1:0] node402;
	wire [3-1:0] node403;
	wire [3-1:0] node407;
	wire [3-1:0] node408;
	wire [3-1:0] node409;
	wire [3-1:0] node410;
	wire [3-1:0] node411;
	wire [3-1:0] node412;
	wire [3-1:0] node417;
	wire [3-1:0] node418;
	wire [3-1:0] node419;
	wire [3-1:0] node423;
	wire [3-1:0] node426;
	wire [3-1:0] node428;
	wire [3-1:0] node431;
	wire [3-1:0] node432;
	wire [3-1:0] node434;
	wire [3-1:0] node435;
	wire [3-1:0] node436;
	wire [3-1:0] node437;
	wire [3-1:0] node441;
	wire [3-1:0] node444;
	wire [3-1:0] node447;
	wire [3-1:0] node448;
	wire [3-1:0] node451;
	wire [3-1:0] node453;
	wire [3-1:0] node456;
	wire [3-1:0] node457;
	wire [3-1:0] node458;
	wire [3-1:0] node459;
	wire [3-1:0] node460;
	wire [3-1:0] node461;
	wire [3-1:0] node462;
	wire [3-1:0] node465;
	wire [3-1:0] node468;
	wire [3-1:0] node469;
	wire [3-1:0] node470;
	wire [3-1:0] node472;
	wire [3-1:0] node476;
	wire [3-1:0] node479;
	wire [3-1:0] node480;
	wire [3-1:0] node481;
	wire [3-1:0] node482;
	wire [3-1:0] node486;
	wire [3-1:0] node487;
	wire [3-1:0] node491;
	wire [3-1:0] node492;
	wire [3-1:0] node493;
	wire [3-1:0] node498;
	wire [3-1:0] node500;
	wire [3-1:0] node501;
	wire [3-1:0] node502;
	wire [3-1:0] node506;
	wire [3-1:0] node508;
	wire [3-1:0] node509;
	wire [3-1:0] node513;
	wire [3-1:0] node514;
	wire [3-1:0] node515;
	wire [3-1:0] node517;
	wire [3-1:0] node518;
	wire [3-1:0] node519;
	wire [3-1:0] node523;
	wire [3-1:0] node524;
	wire [3-1:0] node528;
	wire [3-1:0] node529;
	wire [3-1:0] node531;
	wire [3-1:0] node533;
	wire [3-1:0] node536;
	wire [3-1:0] node537;
	wire [3-1:0] node539;
	wire [3-1:0] node541;
	wire [3-1:0] node544;
	wire [3-1:0] node547;
	wire [3-1:0] node548;
	wire [3-1:0] node549;
	wire [3-1:0] node550;
	wire [3-1:0] node552;
	wire [3-1:0] node555;
	wire [3-1:0] node556;
	wire [3-1:0] node560;
	wire [3-1:0] node561;
	wire [3-1:0] node563;
	wire [3-1:0] node566;
	wire [3-1:0] node569;
	wire [3-1:0] node570;
	wire [3-1:0] node571;
	wire [3-1:0] node573;
	wire [3-1:0] node576;
	wire [3-1:0] node579;
	wire [3-1:0] node581;
	wire [3-1:0] node584;
	wire [3-1:0] node585;
	wire [3-1:0] node586;
	wire [3-1:0] node588;
	wire [3-1:0] node589;
	wire [3-1:0] node594;
	wire [3-1:0] node595;
	wire [3-1:0] node596;
	wire [3-1:0] node597;
	wire [3-1:0] node598;
	wire [3-1:0] node600;
	wire [3-1:0] node602;
	wire [3-1:0] node605;
	wire [3-1:0] node606;
	wire [3-1:0] node610;
	wire [3-1:0] node611;
	wire [3-1:0] node614;
	wire [3-1:0] node616;
	wire [3-1:0] node619;
	wire [3-1:0] node620;
	wire [3-1:0] node621;
	wire [3-1:0] node625;
	wire [3-1:0] node626;
	wire [3-1:0] node629;
	wire [3-1:0] node630;
	wire [3-1:0] node634;
	wire [3-1:0] node635;
	wire [3-1:0] node636;
	wire [3-1:0] node637;
	wire [3-1:0] node638;

	assign outp = (inp[6]) ? node188 : node1;
		assign node1 = (inp[9]) ? node165 : node2;
			assign node2 = (inp[0]) ? node108 : node3;
				assign node3 = (inp[10]) ? node67 : node4;
					assign node4 = (inp[7]) ? node32 : node5;
						assign node5 = (inp[1]) ? node23 : node6;
							assign node6 = (inp[2]) ? node20 : node7;
								assign node7 = (inp[4]) ? node13 : node8;
									assign node8 = (inp[5]) ? 3'b110 : node9;
										assign node9 = (inp[8]) ? 3'b001 : 3'b110;
									assign node13 = (inp[11]) ? node17 : node14;
										assign node14 = (inp[8]) ? 3'b110 : 3'b010;
										assign node17 = (inp[8]) ? 3'b010 : 3'b100;
								assign node20 = (inp[11]) ? 3'b100 : 3'b110;
							assign node23 = (inp[4]) ? node25 : 3'b000;
								assign node25 = (inp[5]) ? node27 : 3'b100;
									assign node27 = (inp[8]) ? node29 : 3'b100;
										assign node29 = (inp[11]) ? 3'b100 : 3'b010;
						assign node32 = (inp[11]) ? node48 : node33;
							assign node33 = (inp[4]) ? node43 : node34;
								assign node34 = (inp[1]) ? 3'b001 : node35;
									assign node35 = (inp[8]) ? node39 : node36;
										assign node36 = (inp[3]) ? 3'b001 : 3'b101;
										assign node39 = (inp[2]) ? 3'b101 : 3'b011;
								assign node43 = (inp[1]) ? node45 : 3'b001;
									assign node45 = (inp[3]) ? 3'b010 : 3'b110;
							assign node48 = (inp[4]) ? node56 : node49;
								assign node49 = (inp[8]) ? node51 : 3'b110;
									assign node51 = (inp[2]) ? node53 : 3'b110;
										assign node53 = (inp[3]) ? 3'b010 : 3'b110;
								assign node56 = (inp[3]) ? node58 : 3'b110;
									assign node58 = (inp[2]) ? node62 : node59;
										assign node59 = (inp[8]) ? 3'b001 : 3'b010;
										assign node62 = (inp[1]) ? 3'b100 : node63;
											assign node63 = (inp[8]) ? 3'b110 : 3'b010;
					assign node67 = (inp[7]) ? node79 : node68;
						assign node68 = (inp[11]) ? 3'b000 : node69;
							assign node69 = (inp[1]) ? 3'b000 : node70;
								assign node70 = (inp[2]) ? 3'b000 : node71;
									assign node71 = (inp[8]) ? 3'b100 : node72;
										assign node72 = (inp[3]) ? 3'b000 : 3'b100;
						assign node79 = (inp[8]) ? node99 : node80;
							assign node80 = (inp[1]) ? node88 : node81;
								assign node81 = (inp[11]) ? 3'b100 : node82;
									assign node82 = (inp[2]) ? 3'b100 : node83;
										assign node83 = (inp[3]) ? 3'b010 : 3'b110;
								assign node88 = (inp[2]) ? node94 : node89;
									assign node89 = (inp[3]) ? node91 : 3'b100;
										assign node91 = (inp[11]) ? 3'b000 : 3'b100;
									assign node94 = (inp[5]) ? node96 : 3'b000;
										assign node96 = (inp[11]) ? 3'b000 : 3'b100;
							assign node99 = (inp[3]) ? 3'b010 : node100;
								assign node100 = (inp[1]) ? 3'b100 : node101;
									assign node101 = (inp[2]) ? node103 : 3'b110;
										assign node103 = (inp[4]) ? 3'b010 : 3'b110;
				assign node108 = (inp[7]) ? node120 : node109;
					assign node109 = (inp[3]) ? 3'b000 : node110;
						assign node110 = (inp[11]) ? 3'b000 : node111;
							assign node111 = (inp[1]) ? 3'b000 : node112;
								assign node112 = (inp[10]) ? 3'b000 : node113;
									assign node113 = (inp[2]) ? 3'b000 : 3'b100;
					assign node120 = (inp[10]) ? node158 : node121;
						assign node121 = (inp[11]) ? node139 : node122;
							assign node122 = (inp[1]) ? node132 : node123;
								assign node123 = (inp[4]) ? node129 : node124;
									assign node124 = (inp[8]) ? 3'b010 : node125;
										assign node125 = (inp[5]) ? 3'b100 : 3'b010;
									assign node129 = (inp[8]) ? 3'b110 : 3'b100;
								assign node132 = (inp[4]) ? node134 : 3'b100;
									assign node134 = (inp[3]) ? node136 : 3'b010;
										assign node136 = (inp[8]) ? 3'b100 : 3'b000;
							assign node139 = (inp[3]) ? node149 : node140;
								assign node140 = (inp[4]) ? node146 : node141;
									assign node141 = (inp[1]) ? 3'b000 : node142;
										assign node142 = (inp[2]) ? 3'b000 : 3'b010;
									assign node146 = (inp[2]) ? 3'b000 : 3'b100;
								assign node149 = (inp[1]) ? node155 : node150;
									assign node150 = (inp[2]) ? node152 : 3'b100;
										assign node152 = (inp[8]) ? 3'b100 : 3'b000;
									assign node155 = (inp[4]) ? 3'b000 : 3'b100;
						assign node158 = (inp[1]) ? 3'b000 : node159;
							assign node159 = (inp[8]) ? node161 : 3'b000;
								assign node161 = (inp[2]) ? 3'b000 : 3'b100;
			assign node165 = (inp[7]) ? node167 : 3'b000;
				assign node167 = (inp[10]) ? 3'b000 : node168;
					assign node168 = (inp[0]) ? 3'b000 : node169;
						assign node169 = (inp[1]) ? 3'b000 : node170;
							assign node170 = (inp[11]) ? node180 : node171;
								assign node171 = (inp[8]) ? node177 : node172;
									assign node172 = (inp[3]) ? 3'b000 : node173;
										assign node173 = (inp[2]) ? 3'b000 : 3'b100;
									assign node177 = (inp[2]) ? 3'b100 : 3'b010;
								assign node180 = (inp[2]) ? 3'b000 : node181;
									assign node181 = (inp[3]) ? 3'b000 : 3'b100;
		assign node188 = (inp[9]) ? node456 : node189;
			assign node189 = (inp[0]) ? node293 : node190;
				assign node190 = (inp[7]) ? node254 : node191;
					assign node191 = (inp[10]) ? node229 : node192;
						assign node192 = (inp[1]) ? node206 : node193;
							assign node193 = (inp[11]) ? node199 : node194;
								assign node194 = (inp[8]) ? 3'b111 : node195;
									assign node195 = (inp[2]) ? 3'b011 : 3'b111;
								assign node199 = (inp[2]) ? node203 : node200;
									assign node200 = (inp[8]) ? 3'b111 : 3'b011;
									assign node203 = (inp[8]) ? 3'b011 : 3'b101;
							assign node206 = (inp[3]) ? node218 : node207;
								assign node207 = (inp[2]) ? node215 : node208;
									assign node208 = (inp[4]) ? 3'b101 : node209;
										assign node209 = (inp[11]) ? 3'b011 : node210;
											assign node210 = (inp[8]) ? 3'b111 : 3'b011;
									assign node215 = (inp[11]) ? 3'b001 : 3'b101;
								assign node218 = (inp[11]) ? node226 : node219;
									assign node219 = (inp[8]) ? 3'b011 : node220;
										assign node220 = (inp[2]) ? node222 : 3'b101;
											assign node222 = (inp[4]) ? 3'b001 : 3'b101;
									assign node226 = (inp[8]) ? 3'b101 : 3'b110;
						assign node229 = (inp[1]) ? node239 : node230;
							assign node230 = (inp[8]) ? node234 : node231;
								assign node231 = (inp[11]) ? 3'b110 : 3'b001;
								assign node234 = (inp[4]) ? node236 : 3'b101;
									assign node236 = (inp[11]) ? 3'b001 : 3'b101;
							assign node239 = (inp[3]) ? node245 : node240;
								assign node240 = (inp[11]) ? 3'b110 : node241;
									assign node241 = (inp[8]) ? 3'b001 : 3'b110;
								assign node245 = (inp[8]) ? 3'b010 : node246;
									assign node246 = (inp[11]) ? node250 : node247;
										assign node247 = (inp[2]) ? 3'b010 : 3'b110;
										assign node250 = (inp[2]) ? 3'b100 : 3'b010;
					assign node254 = (inp[8]) ? node282 : node255;
						assign node255 = (inp[10]) ? node263 : node256;
							assign node256 = (inp[11]) ? node258 : 3'b111;
								assign node258 = (inp[1]) ? node260 : 3'b111;
									assign node260 = (inp[4]) ? 3'b101 : 3'b011;
							assign node263 = (inp[1]) ? node273 : node264;
								assign node264 = (inp[5]) ? node270 : node265;
									assign node265 = (inp[11]) ? 3'b011 : node266;
										assign node266 = (inp[4]) ? 3'b011 : 3'b111;
									assign node270 = (inp[11]) ? 3'b101 : 3'b111;
								assign node273 = (inp[3]) ? 3'b001 : node274;
									assign node274 = (inp[2]) ? node278 : node275;
										assign node275 = (inp[11]) ? 3'b101 : 3'b011;
										assign node278 = (inp[11]) ? 3'b001 : 3'b101;
						assign node282 = (inp[10]) ? node284 : 3'b111;
							assign node284 = (inp[11]) ? node290 : node285;
								assign node285 = (inp[1]) ? node287 : 3'b111;
									assign node287 = (inp[2]) ? 3'b011 : 3'b111;
								assign node290 = (inp[1]) ? 3'b101 : 3'b111;
				assign node293 = (inp[7]) ? node367 : node294;
					assign node294 = (inp[10]) ? node338 : node295;
						assign node295 = (inp[2]) ? node317 : node296;
							assign node296 = (inp[1]) ? node308 : node297;
								assign node297 = (inp[4]) ? node303 : node298;
									assign node298 = (inp[5]) ? 3'b110 : node299;
										assign node299 = (inp[8]) ? 3'b101 : 3'b001;
									assign node303 = (inp[11]) ? 3'b001 : node304;
										assign node304 = (inp[8]) ? 3'b101 : 3'b001;
								assign node308 = (inp[11]) ? node312 : node309;
									assign node309 = (inp[8]) ? 3'b001 : 3'b110;
									assign node312 = (inp[8]) ? node314 : 3'b010;
										assign node314 = (inp[4]) ? 3'b010 : 3'b110;
							assign node317 = (inp[5]) ? node329 : node318;
								assign node318 = (inp[1]) ? node326 : node319;
									assign node319 = (inp[3]) ? node321 : 3'b110;
										assign node321 = (inp[8]) ? 3'b110 : node322;
											assign node322 = (inp[11]) ? 3'b010 : 3'b110;
									assign node326 = (inp[11]) ? 3'b100 : 3'b010;
								assign node329 = (inp[1]) ? node333 : node330;
									assign node330 = (inp[4]) ? 3'b110 : 3'b001;
									assign node333 = (inp[11]) ? 3'b010 : node334;
										assign node334 = (inp[8]) ? 3'b110 : 3'b010;
						assign node338 = (inp[2]) ? node352 : node339;
							assign node339 = (inp[11]) ? node345 : node340;
								assign node340 = (inp[5]) ? node342 : 3'b010;
									assign node342 = (inp[8]) ? 3'b110 : 3'b010;
								assign node345 = (inp[8]) ? node349 : node346;
									assign node346 = (inp[1]) ? 3'b000 : 3'b100;
									assign node349 = (inp[1]) ? 3'b100 : 3'b010;
							assign node352 = (inp[8]) ? node360 : node353;
								assign node353 = (inp[1]) ? 3'b000 : node354;
									assign node354 = (inp[3]) ? node356 : 3'b100;
										assign node356 = (inp[4]) ? 3'b000 : 3'b100;
								assign node360 = (inp[1]) ? node364 : node361;
									assign node361 = (inp[4]) ? 3'b100 : 3'b010;
									assign node364 = (inp[11]) ? 3'b000 : 3'b100;
					assign node367 = (inp[10]) ? node407 : node368;
						assign node368 = (inp[1]) ? node384 : node369;
							assign node369 = (inp[11]) ? node377 : node370;
								assign node370 = (inp[8]) ? 3'b111 : node371;
									assign node371 = (inp[4]) ? 3'b011 : node372;
										assign node372 = (inp[2]) ? 3'b011 : 3'b111;
								assign node377 = (inp[8]) ? 3'b011 : node378;
									assign node378 = (inp[4]) ? node380 : 3'b101;
										assign node380 = (inp[2]) ? 3'b001 : 3'b101;
							assign node384 = (inp[8]) ? node396 : node385;
								assign node385 = (inp[11]) ? node393 : node386;
									assign node386 = (inp[2]) ? node388 : 3'b101;
										assign node388 = (inp[5]) ? node390 : 3'b001;
											assign node390 = (inp[4]) ? 3'b001 : 3'b101;
									assign node393 = (inp[2]) ? 3'b110 : 3'b001;
								assign node396 = (inp[2]) ? node400 : node397;
									assign node397 = (inp[11]) ? 3'b101 : 3'b011;
									assign node400 = (inp[11]) ? node402 : 3'b101;
										assign node402 = (inp[4]) ? 3'b001 : node403;
											assign node403 = (inp[3]) ? 3'b001 : 3'b101;
						assign node407 = (inp[1]) ? node431 : node408;
							assign node408 = (inp[2]) ? node426 : node409;
								assign node409 = (inp[8]) ? node417 : node410;
									assign node410 = (inp[5]) ? 3'b001 : node411;
										assign node411 = (inp[4]) ? 3'b110 : node412;
											assign node412 = (inp[11]) ? 3'b001 : 3'b101;
									assign node417 = (inp[4]) ? node423 : node418;
										assign node418 = (inp[3]) ? 3'b101 : node419;
											assign node419 = (inp[11]) ? 3'b101 : 3'b011;
										assign node423 = (inp[11]) ? 3'b001 : 3'b101;
								assign node426 = (inp[8]) ? node428 : 3'b110;
									assign node428 = (inp[4]) ? 3'b001 : 3'b101;
							assign node431 = (inp[3]) ? node447 : node432;
								assign node432 = (inp[2]) ? node434 : 3'b110;
									assign node434 = (inp[8]) ? node444 : node435;
										assign node435 = (inp[5]) ? node441 : node436;
											assign node436 = (inp[11]) ? 3'b010 : node437;
												assign node437 = (inp[4]) ? 3'b010 : 3'b110;
											assign node441 = (inp[4]) ? 3'b100 : 3'b010;
										assign node444 = (inp[11]) ? 3'b110 : 3'b001;
								assign node447 = (inp[2]) ? node451 : node448;
									assign node448 = (inp[8]) ? 3'b001 : 3'b010;
									assign node451 = (inp[8]) ? node453 : 3'b100;
										assign node453 = (inp[11]) ? 3'b010 : 3'b110;
			assign node456 = (inp[0]) ? node584 : node457;
				assign node457 = (inp[7]) ? node513 : node458;
					assign node458 = (inp[10]) ? node498 : node459;
						assign node459 = (inp[11]) ? node479 : node460;
							assign node460 = (inp[1]) ? node468 : node461;
								assign node461 = (inp[2]) ? node465 : node462;
									assign node462 = (inp[8]) ? 3'b001 : 3'b110;
									assign node465 = (inp[8]) ? 3'b110 : 3'b010;
								assign node468 = (inp[2]) ? node476 : node469;
									assign node469 = (inp[5]) ? 3'b010 : node470;
										assign node470 = (inp[8]) ? node472 : 3'b010;
											assign node472 = (inp[3]) ? 3'b010 : 3'b110;
									assign node476 = (inp[8]) ? 3'b010 : 3'b100;
							assign node479 = (inp[1]) ? node491 : node480;
								assign node480 = (inp[8]) ? node486 : node481;
									assign node481 = (inp[2]) ? 3'b100 : node482;
										assign node482 = (inp[4]) ? 3'b100 : 3'b010;
									assign node486 = (inp[4]) ? 3'b010 : node487;
										assign node487 = (inp[3]) ? 3'b010 : 3'b110;
								assign node491 = (inp[8]) ? 3'b100 : node492;
									assign node492 = (inp[3]) ? 3'b000 : node493;
										assign node493 = (inp[5]) ? 3'b000 : 3'b100;
						assign node498 = (inp[8]) ? node500 : 3'b000;
							assign node500 = (inp[4]) ? node506 : node501;
								assign node501 = (inp[11]) ? 3'b000 : node502;
									assign node502 = (inp[1]) ? 3'b100 : 3'b010;
								assign node506 = (inp[1]) ? node508 : 3'b100;
									assign node508 = (inp[5]) ? 3'b000 : node509;
										assign node509 = (inp[2]) ? 3'b000 : 3'b100;
					assign node513 = (inp[8]) ? node547 : node514;
						assign node514 = (inp[10]) ? node528 : node515;
							assign node515 = (inp[1]) ? node517 : 3'b001;
								assign node517 = (inp[11]) ? node523 : node518;
									assign node518 = (inp[2]) ? 3'b110 : node519;
										assign node519 = (inp[3]) ? 3'b110 : 3'b001;
									assign node523 = (inp[3]) ? 3'b010 : node524;
										assign node524 = (inp[2]) ? 3'b010 : 3'b110;
							assign node528 = (inp[2]) ? node536 : node529;
								assign node529 = (inp[1]) ? node531 : 3'b110;
									assign node531 = (inp[4]) ? node533 : 3'b010;
										assign node533 = (inp[5]) ? 3'b100 : 3'b010;
								assign node536 = (inp[1]) ? node544 : node537;
									assign node537 = (inp[11]) ? node539 : 3'b010;
										assign node539 = (inp[5]) ? node541 : 3'b100;
											assign node541 = (inp[3]) ? 3'b100 : 3'b010;
									assign node544 = (inp[3]) ? 3'b100 : 3'b000;
						assign node547 = (inp[10]) ? node569 : node548;
							assign node548 = (inp[2]) ? node560 : node549;
								assign node549 = (inp[4]) ? node555 : node550;
									assign node550 = (inp[3]) ? node552 : 3'b101;
										assign node552 = (inp[5]) ? 3'b001 : 3'b101;
									assign node555 = (inp[11]) ? 3'b101 : node556;
										assign node556 = (inp[1]) ? 3'b101 : 3'b011;
								assign node560 = (inp[1]) ? node566 : node561;
									assign node561 = (inp[4]) ? node563 : 3'b101;
										assign node563 = (inp[11]) ? 3'b001 : 3'b101;
									assign node566 = (inp[11]) ? 3'b110 : 3'b001;
							assign node569 = (inp[11]) ? node579 : node570;
								assign node570 = (inp[1]) ? node576 : node571;
									assign node571 = (inp[3]) ? node573 : 3'b001;
										assign node573 = (inp[2]) ? 3'b110 : 3'b001;
									assign node576 = (inp[2]) ? 3'b010 : 3'b110;
								assign node579 = (inp[4]) ? node581 : 3'b100;
									assign node581 = (inp[2]) ? 3'b010 : 3'b110;
				assign node584 = (inp[7]) ? node594 : node585;
					assign node585 = (inp[10]) ? 3'b000 : node586;
						assign node586 = (inp[8]) ? node588 : 3'b000;
							assign node588 = (inp[5]) ? 3'b000 : node589;
								assign node589 = (inp[11]) ? 3'b000 : 3'b100;
					assign node594 = (inp[10]) ? node634 : node595;
						assign node595 = (inp[11]) ? node619 : node596;
							assign node596 = (inp[1]) ? node610 : node597;
								assign node597 = (inp[8]) ? node605 : node598;
									assign node598 = (inp[3]) ? node600 : 3'b010;
										assign node600 = (inp[2]) ? node602 : 3'b010;
											assign node602 = (inp[4]) ? 3'b100 : 3'b010;
									assign node605 = (inp[3]) ? 3'b110 : node606;
										assign node606 = (inp[5]) ? 3'b110 : 3'b001;
								assign node610 = (inp[8]) ? node614 : node611;
									assign node611 = (inp[2]) ? 3'b000 : 3'b100;
									assign node614 = (inp[2]) ? node616 : 3'b010;
										assign node616 = (inp[3]) ? 3'b100 : 3'b010;
							assign node619 = (inp[3]) ? node625 : node620;
								assign node620 = (inp[2]) ? 3'b100 : node621;
									assign node621 = (inp[8]) ? 3'b100 : 3'b000;
								assign node625 = (inp[2]) ? node629 : node626;
									assign node626 = (inp[5]) ? 3'b100 : 3'b000;
									assign node629 = (inp[1]) ? 3'b000 : node630;
										assign node630 = (inp[8]) ? 3'b010 : 3'b000;
						assign node634 = (inp[1]) ? 3'b000 : node635;
							assign node635 = (inp[11]) ? 3'b000 : node636;
								assign node636 = (inp[2]) ? 3'b100 : node637;
									assign node637 = (inp[3]) ? 3'b000 : node638;
										assign node638 = (inp[5]) ? 3'b000 : 3'b100;

endmodule