module dtc_split75_bm81 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node7;
	wire [3-1:0] node8;
	wire [3-1:0] node10;
	wire [3-1:0] node11;
	wire [3-1:0] node12;
	wire [3-1:0] node13;
	wire [3-1:0] node20;
	wire [3-1:0] node21;
	wire [3-1:0] node22;
	wire [3-1:0] node23;
	wire [3-1:0] node24;
	wire [3-1:0] node26;
	wire [3-1:0] node29;
	wire [3-1:0] node32;
	wire [3-1:0] node34;
	wire [3-1:0] node37;
	wire [3-1:0] node38;
	wire [3-1:0] node40;
	wire [3-1:0] node42;
	wire [3-1:0] node46;
	wire [3-1:0] node47;
	wire [3-1:0] node48;
	wire [3-1:0] node49;
	wire [3-1:0] node52;
	wire [3-1:0] node55;
	wire [3-1:0] node57;
	wire [3-1:0] node58;
	wire [3-1:0] node62;
	wire [3-1:0] node63;
	wire [3-1:0] node65;
	wire [3-1:0] node68;
	wire [3-1:0] node69;
	wire [3-1:0] node70;
	wire [3-1:0] node71;
	wire [3-1:0] node75;
	wire [3-1:0] node77;
	wire [3-1:0] node81;
	wire [3-1:0] node82;
	wire [3-1:0] node83;
	wire [3-1:0] node84;
	wire [3-1:0] node85;
	wire [3-1:0] node86;
	wire [3-1:0] node89;
	wire [3-1:0] node90;
	wire [3-1:0] node91;
	wire [3-1:0] node96;
	wire [3-1:0] node97;
	wire [3-1:0] node98;
	wire [3-1:0] node99;
	wire [3-1:0] node104;
	wire [3-1:0] node105;
	wire [3-1:0] node108;
	wire [3-1:0] node111;
	wire [3-1:0] node112;
	wire [3-1:0] node113;
	wire [3-1:0] node114;
	wire [3-1:0] node118;
	wire [3-1:0] node119;
	wire [3-1:0] node123;
	wire [3-1:0] node124;
	wire [3-1:0] node127;
	wire [3-1:0] node128;
	wire [3-1:0] node130;
	wire [3-1:0] node134;
	wire [3-1:0] node135;
	wire [3-1:0] node136;
	wire [3-1:0] node138;
	wire [3-1:0] node139;
	wire [3-1:0] node143;
	wire [3-1:0] node144;
	wire [3-1:0] node145;
	wire [3-1:0] node149;
	wire [3-1:0] node150;
	wire [3-1:0] node154;
	wire [3-1:0] node155;
	wire [3-1:0] node156;
	wire [3-1:0] node157;
	wire [3-1:0] node161;
	wire [3-1:0] node162;
	wire [3-1:0] node164;
	wire [3-1:0] node168;
	wire [3-1:0] node169;
	wire [3-1:0] node170;
	wire [3-1:0] node174;
	wire [3-1:0] node175;
	wire [3-1:0] node177;
	wire [3-1:0] node181;
	wire [3-1:0] node182;
	wire [3-1:0] node183;
	wire [3-1:0] node184;
	wire [3-1:0] node188;
	wire [3-1:0] node189;
	wire [3-1:0] node190;
	wire [3-1:0] node193;
	wire [3-1:0] node196;
	wire [3-1:0] node197;
	wire [3-1:0] node201;
	wire [3-1:0] node202;
	wire [3-1:0] node203;
	wire [3-1:0] node206;
	wire [3-1:0] node208;
	wire [3-1:0] node209;
	wire [3-1:0] node210;
	wire [3-1:0] node215;
	wire [3-1:0] node216;
	wire [3-1:0] node219;
	wire [3-1:0] node220;
	wire [3-1:0] node221;
	wire [3-1:0] node225;
	wire [3-1:0] node226;
	wire [3-1:0] node227;
	wire [3-1:0] node232;
	wire [3-1:0] node233;
	wire [3-1:0] node234;
	wire [3-1:0] node235;
	wire [3-1:0] node236;
	wire [3-1:0] node237;
	wire [3-1:0] node238;
	wire [3-1:0] node239;
	wire [3-1:0] node243;
	wire [3-1:0] node244;
	wire [3-1:0] node248;
	wire [3-1:0] node249;
	wire [3-1:0] node250;
	wire [3-1:0] node252;
	wire [3-1:0] node257;
	wire [3-1:0] node258;
	wire [3-1:0] node259;
	wire [3-1:0] node260;
	wire [3-1:0] node265;
	wire [3-1:0] node266;
	wire [3-1:0] node267;
	wire [3-1:0] node269;
	wire [3-1:0] node273;
	wire [3-1:0] node276;
	wire [3-1:0] node277;
	wire [3-1:0] node278;
	wire [3-1:0] node279;
	wire [3-1:0] node282;
	wire [3-1:0] node284;
	wire [3-1:0] node287;
	wire [3-1:0] node288;
	wire [3-1:0] node291;
	wire [3-1:0] node292;
	wire [3-1:0] node296;
	wire [3-1:0] node297;
	wire [3-1:0] node298;
	wire [3-1:0] node300;
	wire [3-1:0] node303;
	wire [3-1:0] node306;
	wire [3-1:0] node307;
	wire [3-1:0] node311;
	wire [3-1:0] node313;
	wire [3-1:0] node314;
	wire [3-1:0] node315;
	wire [3-1:0] node319;
	wire [3-1:0] node320;
	wire [3-1:0] node323;
	wire [3-1:0] node326;
	wire [3-1:0] node327;
	wire [3-1:0] node329;
	wire [3-1:0] node330;
	wire [3-1:0] node331;
	wire [3-1:0] node335;
	wire [3-1:0] node336;
	wire [3-1:0] node338;
	wire [3-1:0] node339;
	wire [3-1:0] node343;
	wire [3-1:0] node344;
	wire [3-1:0] node345;
	wire [3-1:0] node346;
	wire [3-1:0] node351;
	wire [3-1:0] node352;
	wire [3-1:0] node353;
	wire [3-1:0] node359;
	wire [3-1:0] node360;
	wire [3-1:0] node361;
	wire [3-1:0] node362;
	wire [3-1:0] node363;
	wire [3-1:0] node364;
	wire [3-1:0] node365;
	wire [3-1:0] node368;
	wire [3-1:0] node371;
	wire [3-1:0] node372;
	wire [3-1:0] node378;
	wire [3-1:0] node379;
	wire [3-1:0] node380;
	wire [3-1:0] node381;
	wire [3-1:0] node382;
	wire [3-1:0] node385;
	wire [3-1:0] node388;
	wire [3-1:0] node389;
	wire [3-1:0] node391;
	wire [3-1:0] node392;
	wire [3-1:0] node393;
	wire [3-1:0] node398;
	wire [3-1:0] node399;
	wire [3-1:0] node400;
	wire [3-1:0] node401;
	wire [3-1:0] node406;
	wire [3-1:0] node407;
	wire [3-1:0] node411;
	wire [3-1:0] node412;
	wire [3-1:0] node413;
	wire [3-1:0] node416;
	wire [3-1:0] node419;
	wire [3-1:0] node421;
	wire [3-1:0] node424;
	wire [3-1:0] node425;
	wire [3-1:0] node426;
	wire [3-1:0] node427;
	wire [3-1:0] node430;
	wire [3-1:0] node433;
	wire [3-1:0] node435;
	wire [3-1:0] node440;
	wire [3-1:0] node441;
	wire [3-1:0] node442;
	wire [3-1:0] node443;
	wire [3-1:0] node444;
	wire [3-1:0] node446;
	wire [3-1:0] node447;
	wire [3-1:0] node448;
	wire [3-1:0] node449;
	wire [3-1:0] node451;
	wire [3-1:0] node453;
	wire [3-1:0] node456;
	wire [3-1:0] node459;
	wire [3-1:0] node460;
	wire [3-1:0] node461;
	wire [3-1:0] node464;
	wire [3-1:0] node467;
	wire [3-1:0] node468;
	wire [3-1:0] node471;
	wire [3-1:0] node474;
	wire [3-1:0] node475;
	wire [3-1:0] node476;
	wire [3-1:0] node479;
	wire [3-1:0] node482;
	wire [3-1:0] node483;
	wire [3-1:0] node486;
	wire [3-1:0] node489;
	wire [3-1:0] node490;
	wire [3-1:0] node491;
	wire [3-1:0] node492;
	wire [3-1:0] node493;
	wire [3-1:0] node496;
	wire [3-1:0] node498;
	wire [3-1:0] node499;
	wire [3-1:0] node503;
	wire [3-1:0] node504;
	wire [3-1:0] node507;
	wire [3-1:0] node509;
	wire [3-1:0] node512;
	wire [3-1:0] node513;
	wire [3-1:0] node514;
	wire [3-1:0] node517;
	wire [3-1:0] node518;
	wire [3-1:0] node522;
	wire [3-1:0] node523;
	wire [3-1:0] node525;
	wire [3-1:0] node528;
	wire [3-1:0] node530;
	wire [3-1:0] node533;
	wire [3-1:0] node534;
	wire [3-1:0] node535;
	wire [3-1:0] node538;
	wire [3-1:0] node541;
	wire [3-1:0] node542;
	wire [3-1:0] node544;
	wire [3-1:0] node545;
	wire [3-1:0] node549;
	wire [3-1:0] node550;
	wire [3-1:0] node551;
	wire [3-1:0] node552;
	wire [3-1:0] node557;
	wire [3-1:0] node558;
	wire [3-1:0] node559;
	wire [3-1:0] node564;
	wire [3-1:0] node566;
	wire [3-1:0] node568;
	wire [3-1:0] node569;
	wire [3-1:0] node571;
	wire [3-1:0] node572;
	wire [3-1:0] node573;
	wire [3-1:0] node578;
	wire [3-1:0] node579;
	wire [3-1:0] node580;
	wire [3-1:0] node581;
	wire [3-1:0] node585;
	wire [3-1:0] node586;
	wire [3-1:0] node588;
	wire [3-1:0] node592;
	wire [3-1:0] node594;
	wire [3-1:0] node597;
	wire [3-1:0] node598;
	wire [3-1:0] node599;
	wire [3-1:0] node600;
	wire [3-1:0] node601;
	wire [3-1:0] node602;
	wire [3-1:0] node605;
	wire [3-1:0] node608;
	wire [3-1:0] node609;
	wire [3-1:0] node612;
	wire [3-1:0] node614;
	wire [3-1:0] node617;
	wire [3-1:0] node618;
	wire [3-1:0] node619;
	wire [3-1:0] node621;
	wire [3-1:0] node622;
	wire [3-1:0] node626;
	wire [3-1:0] node627;
	wire [3-1:0] node628;
	wire [3-1:0] node632;
	wire [3-1:0] node633;
	wire [3-1:0] node637;
	wire [3-1:0] node638;
	wire [3-1:0] node639;
	wire [3-1:0] node640;
	wire [3-1:0] node641;
	wire [3-1:0] node646;
	wire [3-1:0] node647;
	wire [3-1:0] node651;
	wire [3-1:0] node652;
	wire [3-1:0] node653;
	wire [3-1:0] node657;
	wire [3-1:0] node658;
	wire [3-1:0] node660;
	wire [3-1:0] node664;
	wire [3-1:0] node665;
	wire [3-1:0] node666;
	wire [3-1:0] node667;
	wire [3-1:0] node670;
	wire [3-1:0] node671;
	wire [3-1:0] node672;
	wire [3-1:0] node676;
	wire [3-1:0] node677;
	wire [3-1:0] node681;
	wire [3-1:0] node682;
	wire [3-1:0] node684;
	wire [3-1:0] node685;
	wire [3-1:0] node686;
	wire [3-1:0] node691;
	wire [3-1:0] node693;
	wire [3-1:0] node694;
	wire [3-1:0] node698;
	wire [3-1:0] node699;
	wire [3-1:0] node700;
	wire [3-1:0] node701;
	wire [3-1:0] node702;
	wire [3-1:0] node706;
	wire [3-1:0] node707;
	wire [3-1:0] node708;
	wire [3-1:0] node713;
	wire [3-1:0] node714;
	wire [3-1:0] node716;
	wire [3-1:0] node720;
	wire [3-1:0] node721;
	wire [3-1:0] node722;
	wire [3-1:0] node723;
	wire [3-1:0] node727;
	wire [3-1:0] node728;
	wire [3-1:0] node729;
	wire [3-1:0] node733;
	wire [3-1:0] node736;
	wire [3-1:0] node737;
	wire [3-1:0] node738;
	wire [3-1:0] node740;
	wire [3-1:0] node744;
	wire [3-1:0] node745;
	wire [3-1:0] node749;
	wire [3-1:0] node750;
	wire [3-1:0] node751;
	wire [3-1:0] node752;
	wire [3-1:0] node753;
	wire [3-1:0] node755;
	wire [3-1:0] node756;
	wire [3-1:0] node760;
	wire [3-1:0] node761;
	wire [3-1:0] node762;
	wire [3-1:0] node764;
	wire [3-1:0] node768;
	wire [3-1:0] node769;
	wire [3-1:0] node771;
	wire [3-1:0] node775;
	wire [3-1:0] node777;
	wire [3-1:0] node779;
	wire [3-1:0] node782;
	wire [3-1:0] node783;
	wire [3-1:0] node784;
	wire [3-1:0] node785;
	wire [3-1:0] node786;
	wire [3-1:0] node788;
	wire [3-1:0] node792;
	wire [3-1:0] node793;
	wire [3-1:0] node797;
	wire [3-1:0] node798;
	wire [3-1:0] node801;
	wire [3-1:0] node804;
	wire [3-1:0] node805;
	wire [3-1:0] node806;
	wire [3-1:0] node809;
	wire [3-1:0] node812;
	wire [3-1:0] node813;
	wire [3-1:0] node814;
	wire [3-1:0] node817;
	wire [3-1:0] node819;
	wire [3-1:0] node822;
	wire [3-1:0] node824;
	wire [3-1:0] node827;
	wire [3-1:0] node828;
	wire [3-1:0] node829;
	wire [3-1:0] node830;
	wire [3-1:0] node831;
	wire [3-1:0] node832;
	wire [3-1:0] node834;
	wire [3-1:0] node837;
	wire [3-1:0] node840;
	wire [3-1:0] node841;
	wire [3-1:0] node843;
	wire [3-1:0] node847;
	wire [3-1:0] node848;
	wire [3-1:0] node849;
	wire [3-1:0] node853;
	wire [3-1:0] node854;
	wire [3-1:0] node858;
	wire [3-1:0] node859;
	wire [3-1:0] node860;
	wire [3-1:0] node863;
	wire [3-1:0] node866;
	wire [3-1:0] node867;
	wire [3-1:0] node870;
	wire [3-1:0] node873;
	wire [3-1:0] node874;
	wire [3-1:0] node875;
	wire [3-1:0] node876;
	wire [3-1:0] node877;
	wire [3-1:0] node880;
	wire [3-1:0] node884;
	wire [3-1:0] node885;
	wire [3-1:0] node886;
	wire [3-1:0] node890;
	wire [3-1:0] node891;
	wire [3-1:0] node894;
	wire [3-1:0] node897;
	wire [3-1:0] node898;
	wire [3-1:0] node899;
	wire [3-1:0] node902;
	wire [3-1:0] node904;
	wire [3-1:0] node907;
	wire [3-1:0] node908;
	wire [3-1:0] node910;
	wire [3-1:0] node911;
	wire [3-1:0] node915;
	wire [3-1:0] node917;
	wire [3-1:0] node920;
	wire [3-1:0] node921;
	wire [3-1:0] node922;
	wire [3-1:0] node923;
	wire [3-1:0] node924;
	wire [3-1:0] node925;
	wire [3-1:0] node926;
	wire [3-1:0] node927;
	wire [3-1:0] node928;
	wire [3-1:0] node932;
	wire [3-1:0] node933;
	wire [3-1:0] node935;
	wire [3-1:0] node939;
	wire [3-1:0] node940;
	wire [3-1:0] node941;
	wire [3-1:0] node945;
	wire [3-1:0] node946;
	wire [3-1:0] node950;
	wire [3-1:0] node951;
	wire [3-1:0] node952;
	wire [3-1:0] node955;
	wire [3-1:0] node957;
	wire [3-1:0] node960;
	wire [3-1:0] node961;
	wire [3-1:0] node963;
	wire [3-1:0] node964;
	wire [3-1:0] node968;
	wire [3-1:0] node970;
	wire [3-1:0] node971;
	wire [3-1:0] node975;
	wire [3-1:0] node976;
	wire [3-1:0] node977;
	wire [3-1:0] node978;
	wire [3-1:0] node979;
	wire [3-1:0] node983;
	wire [3-1:0] node984;
	wire [3-1:0] node988;
	wire [3-1:0] node989;
	wire [3-1:0] node990;
	wire [3-1:0] node994;
	wire [3-1:0] node995;
	wire [3-1:0] node997;
	wire [3-1:0] node1001;
	wire [3-1:0] node1002;
	wire [3-1:0] node1003;
	wire [3-1:0] node1004;
	wire [3-1:0] node1006;
	wire [3-1:0] node1010;
	wire [3-1:0] node1013;
	wire [3-1:0] node1014;
	wire [3-1:0] node1017;
	wire [3-1:0] node1020;
	wire [3-1:0] node1021;
	wire [3-1:0] node1022;
	wire [3-1:0] node1023;
	wire [3-1:0] node1025;
	wire [3-1:0] node1026;
	wire [3-1:0] node1030;
	wire [3-1:0] node1031;
	wire [3-1:0] node1032;
	wire [3-1:0] node1036;
	wire [3-1:0] node1037;
	wire [3-1:0] node1039;
	wire [3-1:0] node1043;
	wire [3-1:0] node1044;
	wire [3-1:0] node1045;
	wire [3-1:0] node1046;
	wire [3-1:0] node1050;
	wire [3-1:0] node1051;
	wire [3-1:0] node1055;
	wire [3-1:0] node1056;
	wire [3-1:0] node1057;
	wire [3-1:0] node1059;
	wire [3-1:0] node1063;
	wire [3-1:0] node1064;
	wire [3-1:0] node1066;
	wire [3-1:0] node1070;
	wire [3-1:0] node1071;
	wire [3-1:0] node1072;
	wire [3-1:0] node1073;
	wire [3-1:0] node1075;
	wire [3-1:0] node1076;
	wire [3-1:0] node1080;
	wire [3-1:0] node1081;
	wire [3-1:0] node1082;
	wire [3-1:0] node1086;
	wire [3-1:0] node1087;
	wire [3-1:0] node1091;
	wire [3-1:0] node1092;
	wire [3-1:0] node1096;
	wire [3-1:0] node1097;
	wire [3-1:0] node1098;
	wire [3-1:0] node1099;
	wire [3-1:0] node1101;
	wire [3-1:0] node1105;
	wire [3-1:0] node1108;
	wire [3-1:0] node1109;
	wire [3-1:0] node1112;
	wire [3-1:0] node1115;
	wire [3-1:0] node1116;
	wire [3-1:0] node1117;
	wire [3-1:0] node1118;
	wire [3-1:0] node1119;
	wire [3-1:0] node1120;
	wire [3-1:0] node1122;
	wire [3-1:0] node1123;
	wire [3-1:0] node1126;
	wire [3-1:0] node1129;
	wire [3-1:0] node1131;
	wire [3-1:0] node1134;
	wire [3-1:0] node1135;
	wire [3-1:0] node1136;
	wire [3-1:0] node1137;
	wire [3-1:0] node1141;
	wire [3-1:0] node1144;
	wire [3-1:0] node1145;
	wire [3-1:0] node1147;
	wire [3-1:0] node1150;
	wire [3-1:0] node1153;
	wire [3-1:0] node1155;
	wire [3-1:0] node1157;
	wire [3-1:0] node1158;
	wire [3-1:0] node1162;
	wire [3-1:0] node1163;
	wire [3-1:0] node1164;
	wire [3-1:0] node1165;
	wire [3-1:0] node1166;
	wire [3-1:0] node1169;
	wire [3-1:0] node1172;
	wire [3-1:0] node1173;
	wire [3-1:0] node1176;
	wire [3-1:0] node1179;
	wire [3-1:0] node1180;
	wire [3-1:0] node1183;
	wire [3-1:0] node1184;
	wire [3-1:0] node1187;
	wire [3-1:0] node1188;
	wire [3-1:0] node1192;
	wire [3-1:0] node1193;
	wire [3-1:0] node1194;
	wire [3-1:0] node1197;
	wire [3-1:0] node1200;
	wire [3-1:0] node1201;
	wire [3-1:0] node1204;
	wire [3-1:0] node1206;
	wire [3-1:0] node1209;
	wire [3-1:0] node1210;
	wire [3-1:0] node1211;
	wire [3-1:0] node1212;
	wire [3-1:0] node1213;
	wire [3-1:0] node1216;
	wire [3-1:0] node1218;
	wire [3-1:0] node1221;
	wire [3-1:0] node1222;
	wire [3-1:0] node1223;
	wire [3-1:0] node1227;
	wire [3-1:0] node1228;
	wire [3-1:0] node1230;
	wire [3-1:0] node1234;
	wire [3-1:0] node1235;
	wire [3-1:0] node1236;
	wire [3-1:0] node1238;
	wire [3-1:0] node1242;
	wire [3-1:0] node1243;
	wire [3-1:0] node1245;
	wire [3-1:0] node1248;
	wire [3-1:0] node1250;
	wire [3-1:0] node1253;
	wire [3-1:0] node1254;
	wire [3-1:0] node1255;
	wire [3-1:0] node1256;
	wire [3-1:0] node1258;
	wire [3-1:0] node1259;
	wire [3-1:0] node1263;
	wire [3-1:0] node1266;
	wire [3-1:0] node1267;
	wire [3-1:0] node1269;
	wire [3-1:0] node1270;
	wire [3-1:0] node1274;
	wire [3-1:0] node1276;
	wire [3-1:0] node1279;
	wire [3-1:0] node1280;
	wire [3-1:0] node1281;
	wire [3-1:0] node1283;
	wire [3-1:0] node1287;
	wire [3-1:0] node1288;
	wire [3-1:0] node1290;
	wire [3-1:0] node1294;
	wire [3-1:0] node1295;
	wire [3-1:0] node1296;
	wire [3-1:0] node1297;
	wire [3-1:0] node1298;
	wire [3-1:0] node1299;
	wire [3-1:0] node1300;
	wire [3-1:0] node1301;
	wire [3-1:0] node1305;
	wire [3-1:0] node1306;
	wire [3-1:0] node1310;
	wire [3-1:0] node1311;
	wire [3-1:0] node1312;
	wire [3-1:0] node1317;
	wire [3-1:0] node1318;
	wire [3-1:0] node1319;
	wire [3-1:0] node1321;
	wire [3-1:0] node1322;
	wire [3-1:0] node1325;
	wire [3-1:0] node1328;
	wire [3-1:0] node1329;
	wire [3-1:0] node1332;
	wire [3-1:0] node1333;
	wire [3-1:0] node1337;
	wire [3-1:0] node1338;
	wire [3-1:0] node1339;
	wire [3-1:0] node1341;
	wire [3-1:0] node1345;
	wire [3-1:0] node1348;
	wire [3-1:0] node1350;
	wire [3-1:0] node1351;
	wire [3-1:0] node1352;
	wire [3-1:0] node1357;
	wire [3-1:0] node1358;
	wire [3-1:0] node1359;
	wire [3-1:0] node1360;
	wire [3-1:0] node1362;
	wire [3-1:0] node1368;
	wire [3-1:0] node1369;
	wire [3-1:0] node1370;
	wire [3-1:0] node1371;
	wire [3-1:0] node1372;
	wire [3-1:0] node1373;
	wire [3-1:0] node1376;
	wire [3-1:0] node1379;
	wire [3-1:0] node1380;
	wire [3-1:0] node1383;
	wire [3-1:0] node1384;
	wire [3-1:0] node1385;
	wire [3-1:0] node1389;
	wire [3-1:0] node1390;
	wire [3-1:0] node1394;
	wire [3-1:0] node1395;
	wire [3-1:0] node1396;
	wire [3-1:0] node1398;
	wire [3-1:0] node1401;
	wire [3-1:0] node1403;
	wire [3-1:0] node1406;
	wire [3-1:0] node1407;
	wire [3-1:0] node1410;
	wire [3-1:0] node1412;
	wire [3-1:0] node1415;
	wire [3-1:0] node1416;
	wire [3-1:0] node1417;
	wire [3-1:0] node1418;
	wire [3-1:0] node1420;
	wire [3-1:0] node1421;
	wire [3-1:0] node1425;
	wire [3-1:0] node1427;
	wire [3-1:0] node1430;
	wire [3-1:0] node1432;
	wire [3-1:0] node1434;
	wire [3-1:0] node1436;
	wire [3-1:0] node1439;
	wire [3-1:0] node1440;
	wire [3-1:0] node1441;
	wire [3-1:0] node1443;
	wire [3-1:0] node1447;
	wire [3-1:0] node1448;
	wire [3-1:0] node1450;
	wire [3-1:0] node1454;
	wire [3-1:0] node1455;
	wire [3-1:0] node1456;
	wire [3-1:0] node1457;
	wire [3-1:0] node1458;
	wire [3-1:0] node1460;
	wire [3-1:0] node1463;
	wire [3-1:0] node1465;
	wire [3-1:0] node1468;
	wire [3-1:0] node1469;
	wire [3-1:0] node1471;
	wire [3-1:0] node1472;
	wire [3-1:0] node1477;
	wire [3-1:0] node1478;
	wire [3-1:0] node1479;
	wire [3-1:0] node1481;
	wire [3-1:0] node1485;
	wire [3-1:0] node1486;
	wire [3-1:0] node1488;
	wire [3-1:0] node1492;
	wire [3-1:0] node1494;
	wire [3-1:0] node1495;
	wire [3-1:0] node1496;
	wire [3-1:0] node1498;
	wire [3-1:0] node1500;

	assign outp = (inp[9]) ? node440 : node1;
		assign node1 = (inp[3]) ? node359 : node2;
			assign node2 = (inp[6]) ? node232 : node3;
				assign node3 = (inp[4]) ? node81 : node4;
					assign node4 = (inp[7]) ? node20 : node5;
						assign node5 = (inp[5]) ? node7 : 3'b001;
							assign node7 = (inp[11]) ? 3'b001 : node8;
								assign node8 = (inp[8]) ? node10 : 3'b001;
									assign node10 = (inp[10]) ? 3'b001 : node11;
										assign node11 = (inp[1]) ? 3'b000 : node12;
											assign node12 = (inp[0]) ? 3'b000 : node13;
												assign node13 = (inp[2]) ? 3'b000 : 3'b001;
						assign node20 = (inp[10]) ? node46 : node21;
							assign node21 = (inp[8]) ? node37 : node22;
								assign node22 = (inp[5]) ? node32 : node23;
									assign node23 = (inp[11]) ? node29 : node24;
										assign node24 = (inp[1]) ? node26 : 3'b100;
											assign node26 = (inp[0]) ? 3'b000 : 3'b100;
										assign node29 = (inp[0]) ? 3'b001 : 3'b101;
									assign node32 = (inp[1]) ? node34 : 3'b000;
										assign node34 = (inp[0]) ? 3'b100 : 3'b000;
								assign node37 = (inp[5]) ? 3'b100 : node38;
									assign node38 = (inp[1]) ? node40 : 3'b000;
										assign node40 = (inp[0]) ? node42 : 3'b000;
											assign node42 = (inp[2]) ? 3'b100 : 3'b000;
							assign node46 = (inp[5]) ? node62 : node47;
								assign node47 = (inp[8]) ? node55 : node48;
									assign node48 = (inp[11]) ? node52 : node49;
										assign node49 = (inp[1]) ? 3'b001 : 3'b101;
										assign node52 = (inp[0]) ? 3'b000 : 3'b100;
									assign node55 = (inp[11]) ? node57 : 3'b001;
										assign node57 = (inp[0]) ? 3'b001 : node58;
											assign node58 = (inp[1]) ? 3'b001 : 3'b000;
								assign node62 = (inp[8]) ? node68 : node63;
									assign node63 = (inp[0]) ? node65 : 3'b001;
										assign node65 = (inp[1]) ? 3'b101 : 3'b001;
									assign node68 = (inp[11]) ? 3'b101 : node69;
										assign node69 = (inp[1]) ? node75 : node70;
											assign node70 = (inp[2]) ? 3'b100 : node71;
												assign node71 = (inp[0]) ? 3'b100 : 3'b101;
											assign node75 = (inp[0]) ? node77 : 3'b100;
												assign node77 = (inp[2]) ? 3'b000 : 3'b100;
					assign node81 = (inp[7]) ? node181 : node82;
						assign node82 = (inp[10]) ? node134 : node83;
							assign node83 = (inp[5]) ? node111 : node84;
								assign node84 = (inp[11]) ? node96 : node85;
									assign node85 = (inp[8]) ? node89 : node86;
										assign node86 = (inp[0]) ? 3'b110 : 3'b100;
										assign node89 = (inp[1]) ? 3'b010 : node90;
											assign node90 = (inp[2]) ? 3'b010 : node91;
												assign node91 = (inp[0]) ? 3'b010 : 3'b110;
									assign node96 = (inp[8]) ? node104 : node97;
										assign node97 = (inp[0]) ? 3'b001 : node98;
											assign node98 = (inp[1]) ? 3'b001 : node99;
												assign node99 = (inp[2]) ? 3'b101 : 3'b100;
										assign node104 = (inp[1]) ? node108 : node105;
											assign node105 = (inp[0]) ? 3'b100 : 3'b001;
											assign node108 = (inp[0]) ? 3'b110 : 3'b100;
								assign node111 = (inp[8]) ? node123 : node112;
									assign node112 = (inp[11]) ? node118 : node113;
										assign node113 = (inp[2]) ? 3'b010 : node114;
											assign node114 = (inp[1]) ? 3'b010 : 3'b110;
										assign node118 = (inp[0]) ? 3'b110 : node119;
											assign node119 = (inp[1]) ? 3'b100 : 3'b000;
									assign node123 = (inp[11]) ? node127 : node124;
										assign node124 = (inp[0]) ? 3'b100 : 3'b110;
										assign node127 = (inp[0]) ? 3'b010 : node128;
											assign node128 = (inp[2]) ? node130 : 3'b110;
												assign node130 = (inp[1]) ? 3'b010 : 3'b110;
							assign node134 = (inp[8]) ? node154 : node135;
								assign node135 = (inp[11]) ? node143 : node136;
									assign node136 = (inp[5]) ? node138 : 3'b101;
										assign node138 = (inp[0]) ? 3'b001 : node139;
											assign node139 = (inp[1]) ? 3'b001 : 3'b101;
									assign node143 = (inp[5]) ? node149 : node144;
										assign node144 = (inp[0]) ? 3'b011 : node145;
											assign node145 = (inp[1]) ? 3'b011 : 3'b111;
										assign node149 = (inp[0]) ? 3'b101 : node150;
											assign node150 = (inp[2]) ? 3'b101 : 3'b001;
								assign node154 = (inp[11]) ? node168 : node155;
									assign node155 = (inp[5]) ? node161 : node156;
										assign node156 = (inp[1]) ? 3'b001 : node157;
											assign node157 = (inp[2]) ? 3'b000 : 3'b101;
										assign node161 = (inp[0]) ? 3'b110 : node162;
											assign node162 = (inp[2]) ? node164 : 3'b111;
												assign node164 = (inp[1]) ? 3'b110 : 3'b111;
									assign node168 = (inp[5]) ? node174 : node169;
										assign node169 = (inp[0]) ? 3'b101 : node170;
											assign node170 = (inp[1]) ? 3'b101 : 3'b011;
										assign node174 = (inp[0]) ? 3'b001 : node175;
											assign node175 = (inp[1]) ? node177 : 3'b101;
												assign node177 = (inp[2]) ? 3'b001 : 3'b101;
						assign node181 = (inp[10]) ? node201 : node182;
							assign node182 = (inp[11]) ? node188 : node183;
								assign node183 = (inp[5]) ? 3'b000 : node184;
									assign node184 = (inp[8]) ? 3'b000 : 3'b100;
								assign node188 = (inp[1]) ? node196 : node189;
									assign node189 = (inp[5]) ? node193 : node190;
										assign node190 = (inp[8]) ? 3'b100 : 3'b010;
										assign node193 = (inp[8]) ? 3'b000 : 3'b100;
									assign node196 = (inp[2]) ? 3'b100 : node197;
										assign node197 = (inp[5]) ? 3'b000 : 3'b100;
							assign node201 = (inp[5]) ? node215 : node202;
								assign node202 = (inp[11]) ? node206 : node203;
									assign node203 = (inp[8]) ? 3'b010 : 3'b110;
									assign node206 = (inp[8]) ? node208 : 3'b001;
										assign node208 = (inp[0]) ? 3'b110 : node209;
											assign node209 = (inp[1]) ? 3'b110 : node210;
												assign node210 = (inp[2]) ? 3'b100 : 3'b000;
								assign node215 = (inp[8]) ? node219 : node216;
									assign node216 = (inp[11]) ? 3'b110 : 3'b010;
									assign node219 = (inp[11]) ? node225 : node220;
										assign node220 = (inp[2]) ? 3'b100 : node221;
											assign node221 = (inp[0]) ? 3'b100 : 3'b110;
										assign node225 = (inp[0]) ? 3'b010 : node226;
											assign node226 = (inp[1]) ? 3'b010 : node227;
												assign node227 = (inp[2]) ? 3'b010 : 3'b110;
				assign node232 = (inp[4]) ? node326 : node233;
					assign node233 = (inp[7]) ? node311 : node234;
						assign node234 = (inp[10]) ? node276 : node235;
							assign node235 = (inp[5]) ? node257 : node236;
								assign node236 = (inp[11]) ? node248 : node237;
									assign node237 = (inp[8]) ? node243 : node238;
										assign node238 = (inp[0]) ? 3'b100 : node239;
											assign node239 = (inp[1]) ? 3'b100 : 3'b000;
										assign node243 = (inp[0]) ? 3'b000 : node244;
											assign node244 = (inp[1]) ? 3'b000 : 3'b100;
									assign node248 = (inp[8]) ? 3'b100 : node249;
										assign node249 = (inp[0]) ? 3'b010 : node250;
											assign node250 = (inp[2]) ? node252 : 3'b110;
												assign node252 = (inp[1]) ? 3'b010 : 3'b110;
								assign node257 = (inp[11]) ? node265 : node258;
									assign node258 = (inp[1]) ? 3'b000 : node259;
										assign node259 = (inp[0]) ? 3'b000 : node260;
											assign node260 = (inp[8]) ? 3'b000 : 3'b100;
									assign node265 = (inp[8]) ? node273 : node266;
										assign node266 = (inp[0]) ? 3'b100 : node267;
											assign node267 = (inp[1]) ? node269 : 3'b000;
												assign node269 = (inp[2]) ? 3'b100 : 3'b000;
										assign node273 = (inp[0]) ? 3'b000 : 3'b100;
							assign node276 = (inp[11]) ? node296 : node277;
								assign node277 = (inp[5]) ? node287 : node278;
									assign node278 = (inp[8]) ? node282 : node279;
										assign node279 = (inp[0]) ? 3'b110 : 3'b011;
										assign node282 = (inp[2]) ? node284 : 3'b110;
											assign node284 = (inp[0]) ? 3'b010 : 3'b110;
									assign node287 = (inp[8]) ? node291 : node288;
										assign node288 = (inp[0]) ? 3'b010 : 3'b110;
										assign node291 = (inp[0]) ? 3'b100 : node292;
											assign node292 = (inp[1]) ? 3'b000 : 3'b010;
								assign node296 = (inp[1]) ? node306 : node297;
									assign node297 = (inp[5]) ? node303 : node298;
										assign node298 = (inp[8]) ? node300 : 3'b101;
											assign node300 = (inp[0]) ? 3'b011 : 3'b001;
										assign node303 = (inp[8]) ? 3'b110 : 3'b011;
									assign node306 = (inp[0]) ? 3'b110 : node307;
										assign node307 = (inp[8]) ? 3'b110 : 3'b011;
						assign node311 = (inp[10]) ? node313 : 3'b000;
							assign node313 = (inp[11]) ? node319 : node314;
								assign node314 = (inp[8]) ? 3'b000 : node315;
									assign node315 = (inp[5]) ? 3'b000 : 3'b100;
								assign node319 = (inp[8]) ? node323 : node320;
									assign node320 = (inp[5]) ? 3'b100 : 3'b010;
									assign node323 = (inp[5]) ? 3'b000 : 3'b100;
					assign node326 = (inp[7]) ? 3'b000 : node327;
						assign node327 = (inp[10]) ? node329 : 3'b000;
							assign node329 = (inp[11]) ? node335 : node330;
								assign node330 = (inp[5]) ? 3'b000 : node331;
									assign node331 = (inp[8]) ? 3'b000 : 3'b100;
								assign node335 = (inp[5]) ? node343 : node336;
									assign node336 = (inp[8]) ? node338 : 3'b010;
										assign node338 = (inp[2]) ? 3'b100 : node339;
											assign node339 = (inp[0]) ? 3'b100 : 3'b000;
									assign node343 = (inp[8]) ? node351 : node344;
										assign node344 = (inp[0]) ? 3'b100 : node345;
											assign node345 = (inp[2]) ? 3'b100 : node346;
												assign node346 = (inp[1]) ? 3'b100 : 3'b000;
										assign node351 = (inp[2]) ? 3'b000 : node352;
											assign node352 = (inp[1]) ? 3'b000 : node353;
												assign node353 = (inp[0]) ? 3'b000 : 3'b100;
			assign node359 = (inp[6]) ? 3'b000 : node360;
				assign node360 = (inp[10]) ? node378 : node361;
					assign node361 = (inp[4]) ? 3'b000 : node362;
						assign node362 = (inp[7]) ? 3'b000 : node363;
							assign node363 = (inp[5]) ? node371 : node364;
								assign node364 = (inp[8]) ? node368 : node365;
									assign node365 = (inp[11]) ? 3'b010 : 3'b100;
									assign node368 = (inp[11]) ? 3'b100 : 3'b000;
								assign node371 = (inp[8]) ? 3'b000 : node372;
									assign node372 = (inp[11]) ? 3'b100 : 3'b000;
					assign node378 = (inp[7]) ? node424 : node379;
						assign node379 = (inp[4]) ? node411 : node380;
							assign node380 = (inp[11]) ? node388 : node381;
								assign node381 = (inp[5]) ? node385 : node382;
									assign node382 = (inp[8]) ? 3'b010 : 3'b110;
									assign node385 = (inp[8]) ? 3'b100 : 3'b010;
								assign node388 = (inp[5]) ? node398 : node389;
									assign node389 = (inp[8]) ? node391 : 3'b001;
										assign node391 = (inp[1]) ? 3'b110 : node392;
											assign node392 = (inp[0]) ? 3'b110 : node393;
												assign node393 = (inp[2]) ? 3'b100 : 3'b000;
									assign node398 = (inp[8]) ? node406 : node399;
										assign node399 = (inp[2]) ? 3'b110 : node400;
											assign node400 = (inp[0]) ? 3'b110 : node401;
												assign node401 = (inp[1]) ? 3'b110 : 3'b010;
										assign node406 = (inp[0]) ? 3'b010 : node407;
											assign node407 = (inp[2]) ? 3'b010 : 3'b110;
							assign node411 = (inp[8]) ? node419 : node412;
								assign node412 = (inp[5]) ? node416 : node413;
									assign node413 = (inp[11]) ? 3'b010 : 3'b100;
									assign node416 = (inp[11]) ? 3'b100 : 3'b000;
								assign node419 = (inp[11]) ? node421 : 3'b000;
									assign node421 = (inp[5]) ? 3'b000 : 3'b100;
						assign node424 = (inp[4]) ? 3'b000 : node425;
							assign node425 = (inp[8]) ? node433 : node426;
								assign node426 = (inp[5]) ? node430 : node427;
									assign node427 = (inp[11]) ? 3'b010 : 3'b100;
									assign node430 = (inp[11]) ? 3'b100 : 3'b000;
								assign node433 = (inp[11]) ? node435 : 3'b000;
									assign node435 = (inp[5]) ? 3'b000 : 3'b100;
		assign node440 = (inp[6]) ? node920 : node441;
			assign node441 = (inp[3]) ? node597 : node442;
				assign node442 = (inp[10]) ? node564 : node443;
					assign node443 = (inp[7]) ? node489 : node444;
						assign node444 = (inp[4]) ? node446 : 3'b111;
							assign node446 = (inp[1]) ? node474 : node447;
								assign node447 = (inp[0]) ? node459 : node448;
									assign node448 = (inp[11]) ? node456 : node449;
										assign node449 = (inp[2]) ? node451 : 3'b111;
											assign node451 = (inp[8]) ? node453 : 3'b011;
												assign node453 = (inp[5]) ? 3'b101 : 3'b011;
										assign node456 = (inp[8]) ? 3'b001 : 3'b101;
									assign node459 = (inp[8]) ? node467 : node460;
										assign node460 = (inp[11]) ? node464 : node461;
											assign node461 = (inp[5]) ? 3'b011 : 3'b111;
											assign node464 = (inp[5]) ? 3'b111 : 3'b001;
										assign node467 = (inp[5]) ? node471 : node468;
											assign node468 = (inp[11]) ? 3'b111 : 3'b011;
											assign node471 = (inp[11]) ? 3'b011 : 3'b101;
								assign node474 = (inp[5]) ? node482 : node475;
									assign node475 = (inp[11]) ? node479 : node476;
										assign node476 = (inp[8]) ? 3'b011 : 3'b111;
										assign node479 = (inp[8]) ? 3'b111 : 3'b001;
									assign node482 = (inp[11]) ? node486 : node483;
										assign node483 = (inp[8]) ? 3'b101 : 3'b011;
										assign node486 = (inp[8]) ? 3'b011 : 3'b111;
						assign node489 = (inp[4]) ? node533 : node490;
							assign node490 = (inp[11]) ? node512 : node491;
								assign node491 = (inp[5]) ? node503 : node492;
									assign node492 = (inp[8]) ? node496 : node493;
										assign node493 = (inp[0]) ? 3'b111 : 3'b001;
										assign node496 = (inp[0]) ? node498 : 3'b111;
											assign node498 = (inp[1]) ? 3'b011 : node499;
												assign node499 = (inp[2]) ? 3'b011 : 3'b111;
									assign node503 = (inp[8]) ? node507 : node504;
										assign node504 = (inp[0]) ? 3'b011 : 3'b111;
										assign node507 = (inp[0]) ? node509 : 3'b011;
											assign node509 = (inp[1]) ? 3'b101 : 3'b011;
								assign node512 = (inp[5]) ? node522 : node513;
									assign node513 = (inp[0]) ? node517 : node514;
										assign node514 = (inp[8]) ? 3'b001 : 3'b101;
										assign node517 = (inp[8]) ? 3'b111 : node518;
											assign node518 = (inp[1]) ? 3'b001 : 3'b101;
									assign node522 = (inp[8]) ? node528 : node523;
										assign node523 = (inp[0]) ? node525 : 3'b001;
											assign node525 = (inp[1]) ? 3'b111 : 3'b001;
										assign node528 = (inp[0]) ? node530 : 3'b111;
											assign node530 = (inp[1]) ? 3'b011 : 3'b111;
							assign node533 = (inp[8]) ? node541 : node534;
								assign node534 = (inp[5]) ? node538 : node535;
									assign node535 = (inp[11]) ? 3'b011 : 3'b101;
									assign node538 = (inp[11]) ? 3'b101 : 3'b001;
								assign node541 = (inp[11]) ? node549 : node542;
									assign node542 = (inp[5]) ? node544 : 3'b001;
										assign node544 = (inp[1]) ? 3'b110 : node545;
											assign node545 = (inp[0]) ? 3'b110 : 3'b101;
									assign node549 = (inp[5]) ? node557 : node550;
										assign node550 = (inp[2]) ? 3'b101 : node551;
											assign node551 = (inp[1]) ? 3'b101 : node552;
												assign node552 = (inp[0]) ? 3'b101 : 3'b001;
										assign node557 = (inp[0]) ? 3'b001 : node558;
											assign node558 = (inp[2]) ? 3'b001 : node559;
												assign node559 = (inp[1]) ? 3'b001 : 3'b101;
					assign node564 = (inp[4]) ? node566 : 3'b111;
						assign node566 = (inp[7]) ? node568 : 3'b111;
							assign node568 = (inp[5]) ? node578 : node569;
								assign node569 = (inp[8]) ? node571 : 3'b111;
									assign node571 = (inp[11]) ? 3'b111 : node572;
										assign node572 = (inp[0]) ? 3'b011 : node573;
											assign node573 = (inp[1]) ? 3'b011 : 3'b101;
								assign node578 = (inp[11]) ? node592 : node579;
									assign node579 = (inp[8]) ? node585 : node580;
										assign node580 = (inp[0]) ? 3'b011 : node581;
											assign node581 = (inp[1]) ? 3'b011 : 3'b111;
										assign node585 = (inp[0]) ? 3'b101 : node586;
											assign node586 = (inp[2]) ? node588 : 3'b011;
												assign node588 = (inp[1]) ? 3'b101 : 3'b011;
									assign node592 = (inp[0]) ? node594 : 3'b111;
										assign node594 = (inp[8]) ? 3'b011 : 3'b111;
				assign node597 = (inp[10]) ? node749 : node598;
					assign node598 = (inp[4]) ? node664 : node599;
						assign node599 = (inp[7]) ? node617 : node600;
							assign node600 = (inp[8]) ? node608 : node601;
								assign node601 = (inp[11]) ? node605 : node602;
									assign node602 = (inp[5]) ? 3'b001 : 3'b101;
									assign node605 = (inp[5]) ? 3'b101 : 3'b011;
								assign node608 = (inp[5]) ? node612 : node609;
									assign node609 = (inp[11]) ? 3'b101 : 3'b001;
									assign node612 = (inp[11]) ? node614 : 3'b110;
										assign node614 = (inp[1]) ? 3'b001 : 3'b101;
							assign node617 = (inp[5]) ? node637 : node618;
								assign node618 = (inp[11]) ? node626 : node619;
									assign node619 = (inp[8]) ? node621 : 3'b110;
										assign node621 = (inp[2]) ? 3'b010 : node622;
											assign node622 = (inp[0]) ? 3'b010 : 3'b110;
									assign node626 = (inp[8]) ? node632 : node627;
										assign node627 = (inp[1]) ? 3'b001 : node628;
											assign node628 = (inp[0]) ? 3'b001 : 3'b101;
										assign node632 = (inp[1]) ? 3'b110 : node633;
											assign node633 = (inp[0]) ? 3'b110 : 3'b001;
								assign node637 = (inp[8]) ? node651 : node638;
									assign node638 = (inp[11]) ? node646 : node639;
										assign node639 = (inp[2]) ? 3'b010 : node640;
											assign node640 = (inp[1]) ? 3'b010 : node641;
												assign node641 = (inp[0]) ? 3'b010 : 3'b110;
										assign node646 = (inp[0]) ? 3'b110 : node647;
											assign node647 = (inp[1]) ? 3'b110 : 3'b010;
									assign node651 = (inp[11]) ? node657 : node652;
										assign node652 = (inp[2]) ? 3'b100 : node653;
											assign node653 = (inp[0]) ? 3'b100 : 3'b010;
										assign node657 = (inp[0]) ? 3'b010 : node658;
											assign node658 = (inp[1]) ? node660 : 3'b110;
												assign node660 = (inp[2]) ? 3'b010 : 3'b110;
						assign node664 = (inp[7]) ? node698 : node665;
							assign node665 = (inp[5]) ? node681 : node666;
								assign node666 = (inp[11]) ? node670 : node667;
									assign node667 = (inp[8]) ? 3'b010 : 3'b110;
									assign node670 = (inp[8]) ? node676 : node671;
										assign node671 = (inp[0]) ? 3'b001 : node672;
											assign node672 = (inp[2]) ? 3'b001 : 3'b110;
										assign node676 = (inp[1]) ? 3'b110 : node677;
											assign node677 = (inp[0]) ? 3'b110 : 3'b001;
								assign node681 = (inp[11]) ? node691 : node682;
									assign node682 = (inp[8]) ? node684 : 3'b010;
										assign node684 = (inp[1]) ? 3'b100 : node685;
											assign node685 = (inp[2]) ? 3'b100 : node686;
												assign node686 = (inp[0]) ? 3'b100 : 3'b010;
									assign node691 = (inp[8]) ? node693 : 3'b110;
										assign node693 = (inp[0]) ? 3'b010 : node694;
											assign node694 = (inp[1]) ? 3'b010 : 3'b110;
							assign node698 = (inp[11]) ? node720 : node699;
								assign node699 = (inp[8]) ? node713 : node700;
									assign node700 = (inp[5]) ? node706 : node701;
										assign node701 = (inp[2]) ? 3'b100 : node702;
											assign node702 = (inp[1]) ? 3'b100 : 3'b000;
										assign node706 = (inp[0]) ? 3'b000 : node707;
											assign node707 = (inp[1]) ? 3'b000 : node708;
												assign node708 = (inp[2]) ? 3'b000 : 3'b100;
									assign node713 = (inp[0]) ? 3'b000 : node714;
										assign node714 = (inp[2]) ? node716 : 3'b000;
											assign node716 = (inp[5]) ? 3'b000 : 3'b100;
								assign node720 = (inp[5]) ? node736 : node721;
									assign node721 = (inp[2]) ? node727 : node722;
										assign node722 = (inp[8]) ? 3'b010 : node723;
											assign node723 = (inp[0]) ? 3'b010 : 3'b110;
										assign node727 = (inp[0]) ? node733 : node728;
											assign node728 = (inp[1]) ? 3'b100 : node729;
												assign node729 = (inp[8]) ? 3'b010 : 3'b100;
											assign node733 = (inp[1]) ? 3'b010 : 3'b100;
									assign node736 = (inp[8]) ? node744 : node737;
										assign node737 = (inp[0]) ? 3'b100 : node738;
											assign node738 = (inp[2]) ? node740 : 3'b010;
												assign node740 = (inp[1]) ? 3'b100 : 3'b010;
										assign node744 = (inp[0]) ? 3'b000 : node745;
											assign node745 = (inp[1]) ? 3'b000 : 3'b100;
					assign node749 = (inp[4]) ? node827 : node750;
						assign node750 = (inp[7]) ? node782 : node751;
							assign node751 = (inp[11]) ? node775 : node752;
								assign node752 = (inp[8]) ? node760 : node753;
									assign node753 = (inp[5]) ? node755 : 3'b111;
										assign node755 = (inp[1]) ? 3'b011 : node756;
											assign node756 = (inp[0]) ? 3'b011 : 3'b111;
									assign node760 = (inp[5]) ? node768 : node761;
										assign node761 = (inp[0]) ? 3'b011 : node762;
											assign node762 = (inp[1]) ? node764 : 3'b101;
												assign node764 = (inp[2]) ? 3'b011 : 3'b111;
										assign node768 = (inp[0]) ? 3'b101 : node769;
											assign node769 = (inp[2]) ? node771 : 3'b011;
												assign node771 = (inp[1]) ? 3'b101 : 3'b011;
								assign node775 = (inp[0]) ? node777 : 3'b111;
									assign node777 = (inp[5]) ? node779 : 3'b111;
										assign node779 = (inp[8]) ? 3'b011 : 3'b111;
							assign node782 = (inp[0]) ? node804 : node783;
								assign node783 = (inp[8]) ? node797 : node784;
									assign node784 = (inp[5]) ? node792 : node785;
										assign node785 = (inp[11]) ? 3'b111 : node786;
											assign node786 = (inp[2]) ? node788 : 3'b011;
												assign node788 = (inp[1]) ? 3'b111 : 3'b011;
										assign node792 = (inp[11]) ? 3'b011 : node793;
											assign node793 = (inp[2]) ? 3'b001 : 3'b101;
									assign node797 = (inp[5]) ? node801 : node798;
										assign node798 = (inp[11]) ? 3'b011 : 3'b101;
										assign node801 = (inp[11]) ? 3'b101 : 3'b001;
								assign node804 = (inp[8]) ? node812 : node805;
									assign node805 = (inp[11]) ? node809 : node806;
										assign node806 = (inp[5]) ? 3'b001 : 3'b101;
										assign node809 = (inp[5]) ? 3'b101 : 3'b011;
									assign node812 = (inp[2]) ? node822 : node813;
										assign node813 = (inp[5]) ? node817 : node814;
											assign node814 = (inp[11]) ? 3'b011 : 3'b001;
											assign node817 = (inp[11]) ? node819 : 3'b110;
												assign node819 = (inp[1]) ? 3'b001 : 3'b101;
										assign node822 = (inp[11]) ? node824 : 3'b001;
											assign node824 = (inp[5]) ? 3'b001 : 3'b101;
						assign node827 = (inp[7]) ? node873 : node828;
							assign node828 = (inp[0]) ? node858 : node829;
								assign node829 = (inp[5]) ? node847 : node830;
									assign node830 = (inp[11]) ? node840 : node831;
										assign node831 = (inp[8]) ? node837 : node832;
											assign node832 = (inp[1]) ? node834 : 3'b001;
												assign node834 = (inp[2]) ? 3'b101 : 3'b001;
											assign node837 = (inp[2]) ? 3'b110 : 3'b111;
										assign node840 = (inp[8]) ? 3'b011 : node841;
											assign node841 = (inp[2]) ? node843 : 3'b111;
												assign node843 = (inp[1]) ? 3'b011 : 3'b111;
									assign node847 = (inp[8]) ? node853 : node848;
										assign node848 = (inp[11]) ? 3'b011 : node849;
											assign node849 = (inp[1]) ? 3'b001 : 3'b101;
										assign node853 = (inp[11]) ? 3'b101 : node854;
											assign node854 = (inp[1]) ? 3'b110 : 3'b001;
								assign node858 = (inp[11]) ? node866 : node859;
									assign node859 = (inp[5]) ? node863 : node860;
										assign node860 = (inp[8]) ? 3'b001 : 3'b101;
										assign node863 = (inp[8]) ? 3'b110 : 3'b001;
									assign node866 = (inp[8]) ? node870 : node867;
										assign node867 = (inp[5]) ? 3'b101 : 3'b011;
										assign node870 = (inp[5]) ? 3'b001 : 3'b101;
							assign node873 = (inp[11]) ? node897 : node874;
								assign node874 = (inp[1]) ? node884 : node875;
									assign node875 = (inp[0]) ? 3'b010 : node876;
										assign node876 = (inp[5]) ? node880 : node877;
											assign node877 = (inp[8]) ? 3'b100 : 3'b001;
											assign node880 = (inp[8]) ? 3'b010 : 3'b110;
									assign node884 = (inp[8]) ? node890 : node885;
										assign node885 = (inp[5]) ? 3'b110 : node886;
											assign node886 = (inp[0]) ? 3'b110 : 3'b001;
										assign node890 = (inp[0]) ? node894 : node891;
											assign node891 = (inp[5]) ? 3'b010 : 3'b110;
											assign node894 = (inp[5]) ? 3'b100 : 3'b010;
								assign node897 = (inp[8]) ? node907 : node898;
									assign node898 = (inp[5]) ? node902 : node899;
										assign node899 = (inp[1]) ? 3'b001 : 3'b101;
										assign node902 = (inp[0]) ? node904 : 3'b001;
											assign node904 = (inp[2]) ? 3'b110 : 3'b001;
									assign node907 = (inp[5]) ? node915 : node908;
										assign node908 = (inp[0]) ? node910 : 3'b001;
											assign node910 = (inp[2]) ? 3'b110 : node911;
												assign node911 = (inp[1]) ? 3'b110 : 3'b001;
										assign node915 = (inp[1]) ? node917 : 3'b110;
											assign node917 = (inp[2]) ? 3'b110 : 3'b010;
			assign node920 = (inp[3]) ? node1294 : node921;
				assign node921 = (inp[10]) ? node1115 : node922;
					assign node922 = (inp[4]) ? node1020 : node923;
						assign node923 = (inp[7]) ? node975 : node924;
							assign node924 = (inp[11]) ? node950 : node925;
								assign node925 = (inp[5]) ? node939 : node926;
									assign node926 = (inp[8]) ? node932 : node927;
										assign node927 = (inp[0]) ? 3'b101 : node928;
											assign node928 = (inp[1]) ? 3'b100 : 3'b000;
										assign node932 = (inp[0]) ? 3'b001 : node933;
											assign node933 = (inp[2]) ? node935 : 3'b101;
												assign node935 = (inp[1]) ? 3'b001 : 3'b101;
									assign node939 = (inp[8]) ? node945 : node940;
										assign node940 = (inp[0]) ? 3'b001 : node941;
											assign node941 = (inp[1]) ? 3'b001 : 3'b101;
										assign node945 = (inp[0]) ? 3'b110 : node946;
											assign node946 = (inp[1]) ? 3'b011 : 3'b001;
								assign node950 = (inp[8]) ? node960 : node951;
									assign node951 = (inp[5]) ? node955 : node952;
										assign node952 = (inp[0]) ? 3'b010 : 3'b110;
										assign node955 = (inp[0]) ? node957 : 3'b000;
											assign node957 = (inp[1]) ? 3'b101 : 3'b100;
									assign node960 = (inp[5]) ? node968 : node961;
										assign node961 = (inp[0]) ? node963 : 3'b000;
											assign node963 = (inp[1]) ? 3'b101 : node964;
												assign node964 = (inp[2]) ? 3'b100 : 3'b000;
										assign node968 = (inp[0]) ? node970 : 3'b101;
											assign node970 = (inp[1]) ? 3'b001 : node971;
												assign node971 = (inp[2]) ? 3'b001 : 3'b101;
							assign node975 = (inp[11]) ? node1001 : node976;
								assign node976 = (inp[8]) ? node988 : node977;
									assign node977 = (inp[5]) ? node983 : node978;
										assign node978 = (inp[0]) ? 3'b110 : node979;
											assign node979 = (inp[1]) ? 3'b110 : 3'b010;
										assign node983 = (inp[1]) ? 3'b010 : node984;
											assign node984 = (inp[0]) ? 3'b010 : 3'b110;
									assign node988 = (inp[5]) ? node994 : node989;
										assign node989 = (inp[0]) ? 3'b010 : node990;
											assign node990 = (inp[1]) ? 3'b010 : 3'b110;
										assign node994 = (inp[0]) ? 3'b100 : node995;
											assign node995 = (inp[2]) ? node997 : 3'b010;
												assign node997 = (inp[1]) ? 3'b100 : 3'b010;
								assign node1001 = (inp[8]) ? node1013 : node1002;
									assign node1002 = (inp[0]) ? node1010 : node1003;
										assign node1003 = (inp[5]) ? 3'b001 : node1004;
											assign node1004 = (inp[2]) ? node1006 : 3'b101;
												assign node1006 = (inp[1]) ? 3'b001 : 3'b101;
										assign node1010 = (inp[5]) ? 3'b110 : 3'b001;
									assign node1013 = (inp[5]) ? node1017 : node1014;
										assign node1014 = (inp[0]) ? 3'b110 : 3'b001;
										assign node1017 = (inp[0]) ? 3'b010 : 3'b110;
						assign node1020 = (inp[7]) ? node1070 : node1021;
							assign node1021 = (inp[5]) ? node1043 : node1022;
								assign node1022 = (inp[11]) ? node1030 : node1023;
									assign node1023 = (inp[8]) ? node1025 : 3'b110;
										assign node1025 = (inp[0]) ? 3'b010 : node1026;
											assign node1026 = (inp[1]) ? 3'b010 : 3'b100;
									assign node1030 = (inp[8]) ? node1036 : node1031;
										assign node1031 = (inp[0]) ? 3'b001 : node1032;
											assign node1032 = (inp[2]) ? 3'b110 : 3'b111;
										assign node1036 = (inp[0]) ? 3'b110 : node1037;
											assign node1037 = (inp[2]) ? node1039 : 3'b001;
												assign node1039 = (inp[1]) ? 3'b110 : 3'b001;
								assign node1043 = (inp[11]) ? node1055 : node1044;
									assign node1044 = (inp[8]) ? node1050 : node1045;
										assign node1045 = (inp[0]) ? 3'b010 : node1046;
											assign node1046 = (inp[1]) ? 3'b010 : 3'b110;
										assign node1050 = (inp[1]) ? 3'b100 : node1051;
											assign node1051 = (inp[0]) ? 3'b100 : 3'b010;
									assign node1055 = (inp[8]) ? node1063 : node1056;
										assign node1056 = (inp[0]) ? 3'b110 : node1057;
											assign node1057 = (inp[1]) ? node1059 : 3'b001;
												assign node1059 = (inp[2]) ? 3'b110 : 3'b001;
										assign node1063 = (inp[0]) ? 3'b010 : node1064;
											assign node1064 = (inp[2]) ? node1066 : 3'b110;
												assign node1066 = (inp[1]) ? 3'b010 : 3'b110;
							assign node1070 = (inp[11]) ? node1096 : node1071;
								assign node1071 = (inp[0]) ? node1091 : node1072;
									assign node1072 = (inp[1]) ? node1080 : node1073;
										assign node1073 = (inp[2]) ? node1075 : 3'b100;
											assign node1075 = (inp[8]) ? 3'b100 : node1076;
												assign node1076 = (inp[5]) ? 3'b100 : 3'b000;
										assign node1080 = (inp[2]) ? node1086 : node1081;
											assign node1081 = (inp[5]) ? 3'b100 : node1082;
												assign node1082 = (inp[8]) ? 3'b100 : 3'b000;
											assign node1086 = (inp[8]) ? 3'b000 : node1087;
												assign node1087 = (inp[5]) ? 3'b000 : 3'b100;
									assign node1091 = (inp[5]) ? 3'b000 : node1092;
										assign node1092 = (inp[8]) ? 3'b000 : 3'b100;
								assign node1096 = (inp[5]) ? node1108 : node1097;
									assign node1097 = (inp[8]) ? node1105 : node1098;
										assign node1098 = (inp[0]) ? 3'b010 : node1099;
											assign node1099 = (inp[1]) ? node1101 : 3'b110;
												assign node1101 = (inp[2]) ? 3'b010 : 3'b110;
										assign node1105 = (inp[0]) ? 3'b100 : 3'b010;
									assign node1108 = (inp[8]) ? node1112 : node1109;
										assign node1109 = (inp[0]) ? 3'b100 : 3'b010;
										assign node1112 = (inp[0]) ? 3'b000 : 3'b100;
					assign node1115 = (inp[7]) ? node1209 : node1116;
						assign node1116 = (inp[4]) ? node1162 : node1117;
							assign node1117 = (inp[11]) ? node1153 : node1118;
								assign node1118 = (inp[8]) ? node1134 : node1119;
									assign node1119 = (inp[2]) ? node1129 : node1120;
										assign node1120 = (inp[0]) ? node1122 : 3'b011;
											assign node1122 = (inp[1]) ? node1126 : node1123;
												assign node1123 = (inp[5]) ? 3'b111 : 3'b011;
												assign node1126 = (inp[5]) ? 3'b011 : 3'b111;
										assign node1129 = (inp[1]) ? node1131 : 3'b111;
											assign node1131 = (inp[5]) ? 3'b011 : 3'b111;
									assign node1134 = (inp[5]) ? node1144 : node1135;
										assign node1135 = (inp[0]) ? node1141 : node1136;
											assign node1136 = (inp[1]) ? 3'b111 : node1137;
												assign node1137 = (inp[2]) ? 3'b101 : 3'b111;
											assign node1141 = (inp[1]) ? 3'b011 : 3'b111;
										assign node1144 = (inp[0]) ? node1150 : node1145;
											assign node1145 = (inp[2]) ? node1147 : 3'b011;
												assign node1147 = (inp[1]) ? 3'b001 : 3'b011;
											assign node1150 = (inp[1]) ? 3'b101 : 3'b001;
								assign node1153 = (inp[8]) ? node1155 : 3'b111;
									assign node1155 = (inp[2]) ? node1157 : 3'b111;
										assign node1157 = (inp[5]) ? 3'b011 : node1158;
											assign node1158 = (inp[0]) ? 3'b111 : 3'b011;
							assign node1162 = (inp[5]) ? node1192 : node1163;
								assign node1163 = (inp[0]) ? node1179 : node1164;
									assign node1164 = (inp[1]) ? node1172 : node1165;
										assign node1165 = (inp[8]) ? node1169 : node1166;
											assign node1166 = (inp[11]) ? 3'b111 : 3'b011;
											assign node1169 = (inp[11]) ? 3'b011 : 3'b111;
										assign node1172 = (inp[11]) ? node1176 : node1173;
											assign node1173 = (inp[8]) ? 3'b101 : 3'b011;
											assign node1176 = (inp[8]) ? 3'b011 : 3'b111;
									assign node1179 = (inp[11]) ? node1183 : node1180;
										assign node1180 = (inp[8]) ? 3'b001 : 3'b101;
										assign node1183 = (inp[8]) ? node1187 : node1184;
											assign node1184 = (inp[2]) ? 3'b011 : 3'b111;
											assign node1187 = (inp[1]) ? 3'b101 : node1188;
												assign node1188 = (inp[2]) ? 3'b101 : 3'b011;
								assign node1192 = (inp[8]) ? node1200 : node1193;
									assign node1193 = (inp[11]) ? node1197 : node1194;
										assign node1194 = (inp[0]) ? 3'b001 : 3'b101;
										assign node1197 = (inp[0]) ? 3'b101 : 3'b011;
									assign node1200 = (inp[0]) ? node1204 : node1201;
										assign node1201 = (inp[11]) ? 3'b101 : 3'b001;
										assign node1204 = (inp[11]) ? node1206 : 3'b110;
											assign node1206 = (inp[1]) ? 3'b001 : 3'b101;
						assign node1209 = (inp[4]) ? node1253 : node1210;
							assign node1210 = (inp[11]) ? node1234 : node1211;
								assign node1211 = (inp[5]) ? node1221 : node1212;
									assign node1212 = (inp[0]) ? node1216 : node1213;
										assign node1213 = (inp[8]) ? 3'b101 : 3'b010;
										assign node1216 = (inp[8]) ? node1218 : 3'b101;
											assign node1218 = (inp[2]) ? 3'b001 : 3'b101;
									assign node1221 = (inp[2]) ? node1227 : node1222;
										assign node1222 = (inp[0]) ? 3'b001 : node1223;
											assign node1223 = (inp[8]) ? 3'b001 : 3'b101;
										assign node1227 = (inp[1]) ? 3'b001 : node1228;
											assign node1228 = (inp[8]) ? node1230 : 3'b001;
												assign node1230 = (inp[0]) ? 3'b110 : 3'b001;
								assign node1234 = (inp[8]) ? node1242 : node1235;
									assign node1235 = (inp[5]) ? 3'b011 : node1236;
										assign node1236 = (inp[0]) ? node1238 : 3'b111;
											assign node1238 = (inp[1]) ? 3'b011 : 3'b111;
									assign node1242 = (inp[5]) ? node1248 : node1243;
										assign node1243 = (inp[0]) ? node1245 : 3'b011;
											assign node1245 = (inp[1]) ? 3'b101 : 3'b011;
										assign node1248 = (inp[1]) ? node1250 : 3'b101;
											assign node1250 = (inp[0]) ? 3'b001 : 3'b101;
							assign node1253 = (inp[11]) ? node1279 : node1254;
								assign node1254 = (inp[5]) ? node1266 : node1255;
									assign node1255 = (inp[8]) ? node1263 : node1256;
										assign node1256 = (inp[0]) ? node1258 : 3'b001;
											assign node1258 = (inp[2]) ? 3'b110 : node1259;
												assign node1259 = (inp[1]) ? 3'b110 : 3'b001;
										assign node1263 = (inp[0]) ? 3'b010 : 3'b110;
									assign node1266 = (inp[8]) ? node1274 : node1267;
										assign node1267 = (inp[0]) ? node1269 : 3'b110;
											assign node1269 = (inp[2]) ? 3'b010 : node1270;
												assign node1270 = (inp[1]) ? 3'b010 : 3'b110;
										assign node1274 = (inp[1]) ? node1276 : 3'b010;
											assign node1276 = (inp[0]) ? 3'b100 : 3'b010;
								assign node1279 = (inp[5]) ? node1287 : node1280;
									assign node1280 = (inp[8]) ? 3'b001 : node1281;
										assign node1281 = (inp[0]) ? node1283 : 3'b101;
											assign node1283 = (inp[1]) ? 3'b001 : 3'b101;
									assign node1287 = (inp[8]) ? 3'b110 : node1288;
										assign node1288 = (inp[0]) ? node1290 : 3'b001;
											assign node1290 = (inp[1]) ? 3'b110 : 3'b001;
				assign node1294 = (inp[10]) ? node1368 : node1295;
					assign node1295 = (inp[4]) ? node1357 : node1296;
						assign node1296 = (inp[7]) ? node1348 : node1297;
							assign node1297 = (inp[11]) ? node1317 : node1298;
								assign node1298 = (inp[5]) ? node1310 : node1299;
									assign node1299 = (inp[8]) ? node1305 : node1300;
										assign node1300 = (inp[0]) ? 3'b100 : node1301;
											assign node1301 = (inp[1]) ? 3'b100 : 3'b010;
										assign node1305 = (inp[0]) ? 3'b000 : node1306;
											assign node1306 = (inp[1]) ? 3'b000 : 3'b100;
									assign node1310 = (inp[1]) ? 3'b000 : node1311;
										assign node1311 = (inp[8]) ? 3'b000 : node1312;
											assign node1312 = (inp[0]) ? 3'b000 : 3'b100;
								assign node1317 = (inp[8]) ? node1337 : node1318;
									assign node1318 = (inp[1]) ? node1328 : node1319;
										assign node1319 = (inp[2]) ? node1321 : 3'b010;
											assign node1321 = (inp[5]) ? node1325 : node1322;
												assign node1322 = (inp[0]) ? 3'b010 : 3'b110;
												assign node1325 = (inp[0]) ? 3'b110 : 3'b010;
										assign node1328 = (inp[5]) ? node1332 : node1329;
											assign node1329 = (inp[2]) ? 3'b010 : 3'b110;
											assign node1332 = (inp[2]) ? 3'b100 : node1333;
												assign node1333 = (inp[0]) ? 3'b100 : 3'b010;
									assign node1337 = (inp[5]) ? node1345 : node1338;
										assign node1338 = (inp[0]) ? 3'b100 : node1339;
											assign node1339 = (inp[2]) ? node1341 : 3'b010;
												assign node1341 = (inp[1]) ? 3'b100 : 3'b010;
										assign node1345 = (inp[0]) ? 3'b000 : 3'b100;
							assign node1348 = (inp[11]) ? node1350 : 3'b000;
								assign node1350 = (inp[8]) ? 3'b000 : node1351;
									assign node1351 = (inp[5]) ? 3'b000 : node1352;
										assign node1352 = (inp[0]) ? 3'b000 : 3'b100;
						assign node1357 = (inp[0]) ? 3'b000 : node1358;
							assign node1358 = (inp[5]) ? 3'b000 : node1359;
								assign node1359 = (inp[8]) ? 3'b000 : node1360;
									assign node1360 = (inp[11]) ? node1362 : 3'b000;
										assign node1362 = (inp[7]) ? 3'b000 : 3'b100;
					assign node1368 = (inp[4]) ? node1454 : node1369;
						assign node1369 = (inp[7]) ? node1415 : node1370;
							assign node1370 = (inp[11]) ? node1394 : node1371;
								assign node1371 = (inp[8]) ? node1379 : node1372;
									assign node1372 = (inp[5]) ? node1376 : node1373;
										assign node1373 = (inp[0]) ? 3'b110 : 3'b001;
										assign node1376 = (inp[0]) ? 3'b010 : 3'b110;
									assign node1379 = (inp[0]) ? node1383 : node1380;
										assign node1380 = (inp[5]) ? 3'b010 : 3'b110;
										assign node1383 = (inp[5]) ? node1389 : node1384;
											assign node1384 = (inp[2]) ? 3'b010 : node1385;
												assign node1385 = (inp[1]) ? 3'b010 : 3'b110;
											assign node1389 = (inp[1]) ? 3'b100 : node1390;
												assign node1390 = (inp[2]) ? 3'b100 : 3'b010;
								assign node1394 = (inp[5]) ? node1406 : node1395;
									assign node1395 = (inp[8]) ? node1401 : node1396;
										assign node1396 = (inp[0]) ? node1398 : 3'b101;
											assign node1398 = (inp[2]) ? 3'b001 : 3'b101;
										assign node1401 = (inp[1]) ? node1403 : 3'b001;
											assign node1403 = (inp[0]) ? 3'b110 : 3'b001;
									assign node1406 = (inp[8]) ? node1410 : node1407;
										assign node1407 = (inp[0]) ? 3'b110 : 3'b001;
										assign node1410 = (inp[1]) ? node1412 : 3'b110;
											assign node1412 = (inp[0]) ? 3'b010 : 3'b110;
							assign node1415 = (inp[8]) ? node1439 : node1416;
								assign node1416 = (inp[11]) ? node1430 : node1417;
									assign node1417 = (inp[5]) ? node1425 : node1418;
										assign node1418 = (inp[0]) ? node1420 : 3'b010;
											assign node1420 = (inp[1]) ? 3'b100 : node1421;
												assign node1421 = (inp[2]) ? 3'b100 : 3'b010;
										assign node1425 = (inp[0]) ? node1427 : 3'b100;
											assign node1427 = (inp[1]) ? 3'b000 : 3'b100;
									assign node1430 = (inp[5]) ? node1432 : 3'b110;
										assign node1432 = (inp[0]) ? node1434 : 3'b010;
											assign node1434 = (inp[2]) ? node1436 : 3'b010;
												assign node1436 = (inp[1]) ? 3'b100 : 3'b010;
								assign node1439 = (inp[11]) ? node1447 : node1440;
									assign node1440 = (inp[5]) ? 3'b000 : node1441;
										assign node1441 = (inp[1]) ? node1443 : 3'b100;
											assign node1443 = (inp[0]) ? 3'b000 : 3'b100;
									assign node1447 = (inp[5]) ? 3'b100 : node1448;
										assign node1448 = (inp[1]) ? node1450 : 3'b010;
											assign node1450 = (inp[0]) ? 3'b100 : 3'b010;
						assign node1454 = (inp[7]) ? node1492 : node1455;
							assign node1455 = (inp[11]) ? node1477 : node1456;
								assign node1456 = (inp[5]) ? node1468 : node1457;
									assign node1457 = (inp[8]) ? node1463 : node1458;
										assign node1458 = (inp[2]) ? node1460 : 3'b010;
											assign node1460 = (inp[0]) ? 3'b100 : 3'b010;
										assign node1463 = (inp[0]) ? node1465 : 3'b100;
											assign node1465 = (inp[1]) ? 3'b000 : 3'b100;
									assign node1468 = (inp[8]) ? 3'b000 : node1469;
										assign node1469 = (inp[0]) ? node1471 : 3'b100;
											assign node1471 = (inp[2]) ? 3'b000 : node1472;
												assign node1472 = (inp[1]) ? 3'b000 : 3'b100;
								assign node1477 = (inp[5]) ? node1485 : node1478;
									assign node1478 = (inp[8]) ? 3'b010 : node1479;
										assign node1479 = (inp[1]) ? node1481 : 3'b110;
											assign node1481 = (inp[0]) ? 3'b010 : 3'b110;
									assign node1485 = (inp[8]) ? 3'b100 : node1486;
										assign node1486 = (inp[0]) ? node1488 : 3'b010;
											assign node1488 = (inp[1]) ? 3'b100 : 3'b010;
							assign node1492 = (inp[11]) ? node1494 : 3'b000;
								assign node1494 = (inp[8]) ? 3'b000 : node1495;
									assign node1495 = (inp[5]) ? 3'b000 : node1496;
										assign node1496 = (inp[0]) ? node1498 : 3'b100;
											assign node1498 = (inp[2]) ? node1500 : 3'b100;
												assign node1500 = (inp[1]) ? 3'b000 : 3'b100;

endmodule