module dtc_split66_bm88 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node8;
	wire [3-1:0] node9;
	wire [3-1:0] node10;
	wire [3-1:0] node15;
	wire [3-1:0] node16;
	wire [3-1:0] node18;
	wire [3-1:0] node20;
	wire [3-1:0] node23;
	wire [3-1:0] node26;
	wire [3-1:0] node28;
	wire [3-1:0] node29;
	wire [3-1:0] node31;
	wire [3-1:0] node32;
	wire [3-1:0] node35;
	wire [3-1:0] node36;
	wire [3-1:0] node41;
	wire [3-1:0] node43;
	wire [3-1:0] node44;
	wire [3-1:0] node45;
	wire [3-1:0] node46;
	wire [3-1:0] node47;
	wire [3-1:0] node51;
	wire [3-1:0] node54;
	wire [3-1:0] node56;
	wire [3-1:0] node57;
	wire [3-1:0] node62;
	wire [3-1:0] node63;
	wire [3-1:0] node64;
	wire [3-1:0] node65;
	wire [3-1:0] node66;
	wire [3-1:0] node67;
	wire [3-1:0] node69;
	wire [3-1:0] node70;
	wire [3-1:0] node71;
	wire [3-1:0] node75;
	wire [3-1:0] node78;
	wire [3-1:0] node79;
	wire [3-1:0] node81;
	wire [3-1:0] node84;
	wire [3-1:0] node85;
	wire [3-1:0] node89;
	wire [3-1:0] node90;
	wire [3-1:0] node91;
	wire [3-1:0] node92;
	wire [3-1:0] node96;
	wire [3-1:0] node97;
	wire [3-1:0] node101;
	wire [3-1:0] node102;
	wire [3-1:0] node103;
	wire [3-1:0] node104;
	wire [3-1:0] node108;
	wire [3-1:0] node109;
	wire [3-1:0] node112;
	wire [3-1:0] node115;
	wire [3-1:0] node117;
	wire [3-1:0] node120;
	wire [3-1:0] node121;
	wire [3-1:0] node122;
	wire [3-1:0] node124;
	wire [3-1:0] node126;
	wire [3-1:0] node129;
	wire [3-1:0] node130;
	wire [3-1:0] node132;
	wire [3-1:0] node135;
	wire [3-1:0] node136;
	wire [3-1:0] node140;
	wire [3-1:0] node142;
	wire [3-1:0] node143;
	wire [3-1:0] node145;
	wire [3-1:0] node149;
	wire [3-1:0] node150;
	wire [3-1:0] node151;
	wire [3-1:0] node153;
	wire [3-1:0] node154;
	wire [3-1:0] node158;
	wire [3-1:0] node159;
	wire [3-1:0] node160;
	wire [3-1:0] node164;
	wire [3-1:0] node165;
	wire [3-1:0] node167;
	wire [3-1:0] node169;
	wire [3-1:0] node172;
	wire [3-1:0] node175;
	wire [3-1:0] node177;
	wire [3-1:0] node178;
	wire [3-1:0] node179;
	wire [3-1:0] node181;
	wire [3-1:0] node186;
	wire [3-1:0] node187;
	wire [3-1:0] node188;
	wire [3-1:0] node189;
	wire [3-1:0] node190;
	wire [3-1:0] node191;
	wire [3-1:0] node193;
	wire [3-1:0] node196;
	wire [3-1:0] node198;
	wire [3-1:0] node201;
	wire [3-1:0] node202;
	wire [3-1:0] node205;
	wire [3-1:0] node206;
	wire [3-1:0] node210;
	wire [3-1:0] node211;
	wire [3-1:0] node213;
	wire [3-1:0] node215;
	wire [3-1:0] node218;
	wire [3-1:0] node221;
	wire [3-1:0] node222;
	wire [3-1:0] node223;
	wire [3-1:0] node224;
	wire [3-1:0] node225;
	wire [3-1:0] node228;
	wire [3-1:0] node231;
	wire [3-1:0] node232;
	wire [3-1:0] node236;
	wire [3-1:0] node238;
	wire [3-1:0] node241;
	wire [3-1:0] node242;
	wire [3-1:0] node243;
	wire [3-1:0] node244;
	wire [3-1:0] node247;
	wire [3-1:0] node250;
	wire [3-1:0] node251;
	wire [3-1:0] node254;
	wire [3-1:0] node257;
	wire [3-1:0] node258;
	wire [3-1:0] node259;
	wire [3-1:0] node260;
	wire [3-1:0] node263;
	wire [3-1:0] node266;
	wire [3-1:0] node267;
	wire [3-1:0] node270;
	wire [3-1:0] node273;
	wire [3-1:0] node274;
	wire [3-1:0] node277;
	wire [3-1:0] node280;
	wire [3-1:0] node281;
	wire [3-1:0] node282;
	wire [3-1:0] node283;
	wire [3-1:0] node284;
	wire [3-1:0] node285;
	wire [3-1:0] node288;
	wire [3-1:0] node289;
	wire [3-1:0] node293;
	wire [3-1:0] node294;
	wire [3-1:0] node297;
	wire [3-1:0] node300;
	wire [3-1:0] node301;
	wire [3-1:0] node303;
	wire [3-1:0] node305;
	wire [3-1:0] node308;
	wire [3-1:0] node311;
	wire [3-1:0] node312;
	wire [3-1:0] node313;
	wire [3-1:0] node316;
	wire [3-1:0] node318;
	wire [3-1:0] node319;
	wire [3-1:0] node323;
	wire [3-1:0] node325;
	wire [3-1:0] node326;
	wire [3-1:0] node329;
	wire [3-1:0] node332;
	wire [3-1:0] node333;
	wire [3-1:0] node334;
	wire [3-1:0] node335;
	wire [3-1:0] node338;
	wire [3-1:0] node339;
	wire [3-1:0] node343;
	wire [3-1:0] node344;
	wire [3-1:0] node346;
	wire [3-1:0] node350;
	wire [3-1:0] node351;
	wire [3-1:0] node352;
	wire [3-1:0] node356;
	wire [3-1:0] node357;
	wire [3-1:0] node359;
	wire [3-1:0] node360;
	wire [3-1:0] node365;
	wire [3-1:0] node366;
	wire [3-1:0] node367;
	wire [3-1:0] node368;
	wire [3-1:0] node369;
	wire [3-1:0] node370;
	wire [3-1:0] node371;
	wire [3-1:0] node372;
	wire [3-1:0] node373;
	wire [3-1:0] node377;
	wire [3-1:0] node380;
	wire [3-1:0] node382;
	wire [3-1:0] node384;
	wire [3-1:0] node387;
	wire [3-1:0] node388;
	wire [3-1:0] node389;
	wire [3-1:0] node390;
	wire [3-1:0] node399;
	wire [3-1:0] node400;
	wire [3-1:0] node401;
	wire [3-1:0] node402;
	wire [3-1:0] node403;
	wire [3-1:0] node404;
	wire [3-1:0] node405;
	wire [3-1:0] node407;
	wire [3-1:0] node409;
	wire [3-1:0] node412;
	wire [3-1:0] node413;
	wire [3-1:0] node416;
	wire [3-1:0] node419;
	wire [3-1:0] node421;
	wire [3-1:0] node422;
	wire [3-1:0] node426;
	wire [3-1:0] node427;
	wire [3-1:0] node429;
	wire [3-1:0] node433;
	wire [3-1:0] node434;
	wire [3-1:0] node435;
	wire [3-1:0] node437;
	wire [3-1:0] node440;
	wire [3-1:0] node441;
	wire [3-1:0] node446;
	wire [3-1:0] node447;
	wire [3-1:0] node449;
	wire [3-1:0] node450;
	wire [3-1:0] node451;
	wire [3-1:0] node454;
	wire [3-1:0] node457;
	wire [3-1:0] node458;
	wire [3-1:0] node459;
	wire [3-1:0] node462;
	wire [3-1:0] node465;
	wire [3-1:0] node466;
	wire [3-1:0] node469;
	wire [3-1:0] node472;
	wire [3-1:0] node473;
	wire [3-1:0] node474;
	wire [3-1:0] node475;
	wire [3-1:0] node477;
	wire [3-1:0] node481;
	wire [3-1:0] node482;
	wire [3-1:0] node483;
	wire [3-1:0] node486;
	wire [3-1:0] node489;
	wire [3-1:0] node491;
	wire [3-1:0] node494;
	wire [3-1:0] node495;
	wire [3-1:0] node496;
	wire [3-1:0] node501;
	wire [3-1:0] node502;
	wire [3-1:0] node503;
	wire [3-1:0] node505;
	wire [3-1:0] node506;
	wire [3-1:0] node507;
	wire [3-1:0] node509;
	wire [3-1:0] node512;
	wire [3-1:0] node513;
	wire [3-1:0] node517;
	wire [3-1:0] node518;
	wire [3-1:0] node521;
	wire [3-1:0] node522;
	wire [3-1:0] node524;
	wire [3-1:0] node527;
	wire [3-1:0] node528;
	wire [3-1:0] node531;
	wire [3-1:0] node535;
	wire [3-1:0] node536;
	wire [3-1:0] node537;
	wire [3-1:0] node538;
	wire [3-1:0] node539;
	wire [3-1:0] node546;
	wire [3-1:0] node547;
	wire [3-1:0] node548;
	wire [3-1:0] node549;
	wire [3-1:0] node550;
	wire [3-1:0] node552;
	wire [3-1:0] node554;
	wire [3-1:0] node558;
	wire [3-1:0] node559;
	wire [3-1:0] node560;
	wire [3-1:0] node562;
	wire [3-1:0] node563;
	wire [3-1:0] node565;
	wire [3-1:0] node569;
	wire [3-1:0] node570;
	wire [3-1:0] node571;
	wire [3-1:0] node572;
	wire [3-1:0] node576;
	wire [3-1:0] node577;
	wire [3-1:0] node578;
	wire [3-1:0] node581;
	wire [3-1:0] node584;
	wire [3-1:0] node585;
	wire [3-1:0] node589;
	wire [3-1:0] node590;
	wire [3-1:0] node591;
	wire [3-1:0] node592;
	wire [3-1:0] node596;
	wire [3-1:0] node597;
	wire [3-1:0] node601;
	wire [3-1:0] node602;
	wire [3-1:0] node603;
	wire [3-1:0] node607;
	wire [3-1:0] node609;
	wire [3-1:0] node610;
	wire [3-1:0] node613;
	wire [3-1:0] node616;
	wire [3-1:0] node618;
	wire [3-1:0] node619;
	wire [3-1:0] node621;
	wire [3-1:0] node622;
	wire [3-1:0] node623;
	wire [3-1:0] node626;
	wire [3-1:0] node629;
	wire [3-1:0] node632;
	wire [3-1:0] node633;
	wire [3-1:0] node634;
	wire [3-1:0] node636;
	wire [3-1:0] node640;
	wire [3-1:0] node641;
	wire [3-1:0] node645;
	wire [3-1:0] node646;
	wire [3-1:0] node647;
	wire [3-1:0] node648;
	wire [3-1:0] node649;
	wire [3-1:0] node650;
	wire [3-1:0] node653;
	wire [3-1:0] node654;
	wire [3-1:0] node655;
	wire [3-1:0] node660;
	wire [3-1:0] node661;
	wire [3-1:0] node663;
	wire [3-1:0] node666;
	wire [3-1:0] node667;
	wire [3-1:0] node670;
	wire [3-1:0] node671;
	wire [3-1:0] node675;
	wire [3-1:0] node676;
	wire [3-1:0] node677;
	wire [3-1:0] node679;
	wire [3-1:0] node682;
	wire [3-1:0] node684;
	wire [3-1:0] node686;
	wire [3-1:0] node689;
	wire [3-1:0] node691;
	wire [3-1:0] node692;
	wire [3-1:0] node695;
	wire [3-1:0] node697;
	wire [3-1:0] node700;
	wire [3-1:0] node701;
	wire [3-1:0] node702;
	wire [3-1:0] node703;
	wire [3-1:0] node706;
	wire [3-1:0] node707;
	wire [3-1:0] node708;
	wire [3-1:0] node709;
	wire [3-1:0] node713;
	wire [3-1:0] node717;
	wire [3-1:0] node718;
	wire [3-1:0] node719;
	wire [3-1:0] node721;
	wire [3-1:0] node722;
	wire [3-1:0] node726;
	wire [3-1:0] node727;
	wire [3-1:0] node729;
	wire [3-1:0] node733;
	wire [3-1:0] node736;
	wire [3-1:0] node737;
	wire [3-1:0] node738;
	wire [3-1:0] node741;
	wire [3-1:0] node742;
	wire [3-1:0] node743;
	wire [3-1:0] node748;
	wire [3-1:0] node749;
	wire [3-1:0] node750;
	wire [3-1:0] node751;
	wire [3-1:0] node752;
	wire [3-1:0] node755;
	wire [3-1:0] node759;
	wire [3-1:0] node760;
	wire [3-1:0] node763;
	wire [3-1:0] node766;
	wire [3-1:0] node768;
	wire [3-1:0] node770;
	wire [3-1:0] node771;
	wire [3-1:0] node775;
	wire [3-1:0] node776;
	wire [3-1:0] node777;
	wire [3-1:0] node778;
	wire [3-1:0] node779;
	wire [3-1:0] node783;
	wire [3-1:0] node784;
	wire [3-1:0] node785;
	wire [3-1:0] node789;
	wire [3-1:0] node792;
	wire [3-1:0] node794;
	wire [3-1:0] node795;
	wire [3-1:0] node799;
	wire [3-1:0] node800;
	wire [3-1:0] node801;
	wire [3-1:0] node802;
	wire [3-1:0] node804;
	wire [3-1:0] node806;
	wire [3-1:0] node807;
	wire [3-1:0] node811;
	wire [3-1:0] node812;
	wire [3-1:0] node814;
	wire [3-1:0] node817;
	wire [3-1:0] node819;
	wire [3-1:0] node822;
	wire [3-1:0] node823;
	wire [3-1:0] node824;
	wire [3-1:0] node826;
	wire [3-1:0] node830;
	wire [3-1:0] node831;
	wire [3-1:0] node834;
	wire [3-1:0] node835;
	wire [3-1:0] node838;
	wire [3-1:0] node841;
	wire [3-1:0] node842;
	wire [3-1:0] node843;
	wire [3-1:0] node845;
	wire [3-1:0] node848;
	wire [3-1:0] node849;
	wire [3-1:0] node850;
	wire [3-1:0] node853;
	wire [3-1:0] node856;
	wire [3-1:0] node859;
	wire [3-1:0] node860;
	wire [3-1:0] node862;
	wire [3-1:0] node865;
	wire [3-1:0] node866;
	wire [3-1:0] node869;
	wire [3-1:0] node870;
	wire [3-1:0] node873;
	wire [3-1:0] node876;
	wire [3-1:0] node877;
	wire [3-1:0] node878;
	wire [3-1:0] node879;
	wire [3-1:0] node880;
	wire [3-1:0] node881;
	wire [3-1:0] node884;
	wire [3-1:0] node885;
	wire [3-1:0] node886;
	wire [3-1:0] node888;
	wire [3-1:0] node893;
	wire [3-1:0] node894;
	wire [3-1:0] node896;
	wire [3-1:0] node898;
	wire [3-1:0] node900;
	wire [3-1:0] node903;
	wire [3-1:0] node906;
	wire [3-1:0] node907;
	wire [3-1:0] node908;
	wire [3-1:0] node910;
	wire [3-1:0] node911;
	wire [3-1:0] node913;
	wire [3-1:0] node915;
	wire [3-1:0] node919;
	wire [3-1:0] node922;
	wire [3-1:0] node923;
	wire [3-1:0] node926;
	wire [3-1:0] node927;
	wire [3-1:0] node928;
	wire [3-1:0] node933;
	wire [3-1:0] node934;
	wire [3-1:0] node935;
	wire [3-1:0] node936;
	wire [3-1:0] node937;
	wire [3-1:0] node938;
	wire [3-1:0] node940;
	wire [3-1:0] node942;
	wire [3-1:0] node945;
	wire [3-1:0] node946;
	wire [3-1:0] node949;
	wire [3-1:0] node950;
	wire [3-1:0] node954;
	wire [3-1:0] node955;
	wire [3-1:0] node957;
	wire [3-1:0] node958;
	wire [3-1:0] node961;
	wire [3-1:0] node965;
	wire [3-1:0] node966;
	wire [3-1:0] node967;
	wire [3-1:0] node968;
	wire [3-1:0] node971;
	wire [3-1:0] node975;
	wire [3-1:0] node976;
	wire [3-1:0] node977;
	wire [3-1:0] node980;
	wire [3-1:0] node981;
	wire [3-1:0] node985;
	wire [3-1:0] node986;
	wire [3-1:0] node987;
	wire [3-1:0] node991;
	wire [3-1:0] node994;
	wire [3-1:0] node995;
	wire [3-1:0] node996;
	wire [3-1:0] node997;
	wire [3-1:0] node998;
	wire [3-1:0] node1001;
	wire [3-1:0] node1004;
	wire [3-1:0] node1005;
	wire [3-1:0] node1008;
	wire [3-1:0] node1011;
	wire [3-1:0] node1012;
	wire [3-1:0] node1013;
	wire [3-1:0] node1016;
	wire [3-1:0] node1019;
	wire [3-1:0] node1020;
	wire [3-1:0] node1024;
	wire [3-1:0] node1025;
	wire [3-1:0] node1026;
	wire [3-1:0] node1028;
	wire [3-1:0] node1031;
	wire [3-1:0] node1032;
	wire [3-1:0] node1035;
	wire [3-1:0] node1038;
	wire [3-1:0] node1039;
	wire [3-1:0] node1040;
	wire [3-1:0] node1041;
	wire [3-1:0] node1045;
	wire [3-1:0] node1047;
	wire [3-1:0] node1051;
	wire [3-1:0] node1052;
	wire [3-1:0] node1054;
	wire [3-1:0] node1055;
	wire [3-1:0] node1056;
	wire [3-1:0] node1061;
	wire [3-1:0] node1062;
	wire [3-1:0] node1063;
	wire [3-1:0] node1065;
	wire [3-1:0] node1067;
	wire [3-1:0] node1070;
	wire [3-1:0] node1072;
	wire [3-1:0] node1076;
	wire [3-1:0] node1077;
	wire [3-1:0] node1078;
	wire [3-1:0] node1079;
	wire [3-1:0] node1080;
	wire [3-1:0] node1081;
	wire [3-1:0] node1083;
	wire [3-1:0] node1084;
	wire [3-1:0] node1088;
	wire [3-1:0] node1089;
	wire [3-1:0] node1090;
	wire [3-1:0] node1094;
	wire [3-1:0] node1097;
	wire [3-1:0] node1098;
	wire [3-1:0] node1099;
	wire [3-1:0] node1101;
	wire [3-1:0] node1104;
	wire [3-1:0] node1105;
	wire [3-1:0] node1109;
	wire [3-1:0] node1110;
	wire [3-1:0] node1111;
	wire [3-1:0] node1114;
	wire [3-1:0] node1117;
	wire [3-1:0] node1118;
	wire [3-1:0] node1122;
	wire [3-1:0] node1123;
	wire [3-1:0] node1124;
	wire [3-1:0] node1125;
	wire [3-1:0] node1126;
	wire [3-1:0] node1128;
	wire [3-1:0] node1131;
	wire [3-1:0] node1134;
	wire [3-1:0] node1136;
	wire [3-1:0] node1138;
	wire [3-1:0] node1141;
	wire [3-1:0] node1142;
	wire [3-1:0] node1143;
	wire [3-1:0] node1147;
	wire [3-1:0] node1149;
	wire [3-1:0] node1152;
	wire [3-1:0] node1153;
	wire [3-1:0] node1154;
	wire [3-1:0] node1157;
	wire [3-1:0] node1158;
	wire [3-1:0] node1159;
	wire [3-1:0] node1164;
	wire [3-1:0] node1166;
	wire [3-1:0] node1167;
	wire [3-1:0] node1168;
	wire [3-1:0] node1173;
	wire [3-1:0] node1174;
	wire [3-1:0] node1175;
	wire [3-1:0] node1176;
	wire [3-1:0] node1177;
	wire [3-1:0] node1180;
	wire [3-1:0] node1183;
	wire [3-1:0] node1184;
	wire [3-1:0] node1188;
	wire [3-1:0] node1189;
	wire [3-1:0] node1190;
	wire [3-1:0] node1191;
	wire [3-1:0] node1195;
	wire [3-1:0] node1198;
	wire [3-1:0] node1199;
	wire [3-1:0] node1200;
	wire [3-1:0] node1204;
	wire [3-1:0] node1207;
	wire [3-1:0] node1208;
	wire [3-1:0] node1209;
	wire [3-1:0] node1211;
	wire [3-1:0] node1212;
	wire [3-1:0] node1214;
	wire [3-1:0] node1218;
	wire [3-1:0] node1219;
	wire [3-1:0] node1221;
	wire [3-1:0] node1223;
	wire [3-1:0] node1226;
	wire [3-1:0] node1227;
	wire [3-1:0] node1230;
	wire [3-1:0] node1233;
	wire [3-1:0] node1234;
	wire [3-1:0] node1235;
	wire [3-1:0] node1236;
	wire [3-1:0] node1240;
	wire [3-1:0] node1241;
	wire [3-1:0] node1245;
	wire [3-1:0] node1247;
	wire [3-1:0] node1248;
	wire [3-1:0] node1252;
	wire [3-1:0] node1253;
	wire [3-1:0] node1254;
	wire [3-1:0] node1255;
	wire [3-1:0] node1256;
	wire [3-1:0] node1257;
	wire [3-1:0] node1260;
	wire [3-1:0] node1263;
	wire [3-1:0] node1264;
	wire [3-1:0] node1265;
	wire [3-1:0] node1270;
	wire [3-1:0] node1271;
	wire [3-1:0] node1272;
	wire [3-1:0] node1275;
	wire [3-1:0] node1276;
	wire [3-1:0] node1280;
	wire [3-1:0] node1281;
	wire [3-1:0] node1284;
	wire [3-1:0] node1285;
	wire [3-1:0] node1289;
	wire [3-1:0] node1290;
	wire [3-1:0] node1291;
	wire [3-1:0] node1292;
	wire [3-1:0] node1293;
	wire [3-1:0] node1296;
	wire [3-1:0] node1299;
	wire [3-1:0] node1300;
	wire [3-1:0] node1303;
	wire [3-1:0] node1304;
	wire [3-1:0] node1308;
	wire [3-1:0] node1309;
	wire [3-1:0] node1310;
	wire [3-1:0] node1311;
	wire [3-1:0] node1315;
	wire [3-1:0] node1318;
	wire [3-1:0] node1320;
	wire [3-1:0] node1321;
	wire [3-1:0] node1325;
	wire [3-1:0] node1326;
	wire [3-1:0] node1327;
	wire [3-1:0] node1329;
	wire [3-1:0] node1333;
	wire [3-1:0] node1334;
	wire [3-1:0] node1335;
	wire [3-1:0] node1339;
	wire [3-1:0] node1340;
	wire [3-1:0] node1344;
	wire [3-1:0] node1345;
	wire [3-1:0] node1346;
	wire [3-1:0] node1347;
	wire [3-1:0] node1348;
	wire [3-1:0] node1351;
	wire [3-1:0] node1354;
	wire [3-1:0] node1355;
	wire [3-1:0] node1358;
	wire [3-1:0] node1359;
	wire [3-1:0] node1363;
	wire [3-1:0] node1365;
	wire [3-1:0] node1366;
	wire [3-1:0] node1369;
	wire [3-1:0] node1372;
	wire [3-1:0] node1373;
	wire [3-1:0] node1374;
	wire [3-1:0] node1375;
	wire [3-1:0] node1380;
	wire [3-1:0] node1381;
	wire [3-1:0] node1382;
	wire [3-1:0] node1383;
	wire [3-1:0] node1386;
	wire [3-1:0] node1389;
	wire [3-1:0] node1391;
	wire [3-1:0] node1394;
	wire [3-1:0] node1395;
	wire [3-1:0] node1397;
	wire [3-1:0] node1399;

	assign outp = (inp[6]) ? node546 : node1;
		assign node1 = (inp[3]) ? node365 : node2;
			assign node2 = (inp[0]) ? node62 : node3;
				assign node3 = (inp[9]) ? node41 : node4;
					assign node4 = (inp[7]) ? node26 : node5;
						assign node5 = (inp[10]) ? node15 : node6;
							assign node6 = (inp[5]) ? node8 : 3'b000;
								assign node8 = (inp[8]) ? 3'b000 : node9;
									assign node9 = (inp[4]) ? 3'b010 : node10;
										assign node10 = (inp[11]) ? 3'b000 : 3'b010;
							assign node15 = (inp[8]) ? node23 : node16;
								assign node16 = (inp[5]) ? node18 : 3'b010;
									assign node18 = (inp[11]) ? node20 : 3'b100;
										assign node20 = (inp[4]) ? 3'b100 : 3'b110;
								assign node23 = (inp[5]) ? 3'b010 : 3'b000;
						assign node26 = (inp[5]) ? node28 : 3'b000;
							assign node28 = (inp[8]) ? 3'b000 : node29;
								assign node29 = (inp[2]) ? node31 : 3'b000;
									assign node31 = (inp[4]) ? node35 : node32;
										assign node32 = (inp[10]) ? 3'b010 : 3'b000;
										assign node35 = (inp[10]) ? 3'b000 : node36;
											assign node36 = (inp[11]) ? 3'b000 : 3'b010;
					assign node41 = (inp[5]) ? node43 : 3'b000;
						assign node43 = (inp[8]) ? 3'b000 : node44;
							assign node44 = (inp[4]) ? node54 : node45;
								assign node45 = (inp[10]) ? node51 : node46;
									assign node46 = (inp[7]) ? 3'b000 : node47;
										assign node47 = (inp[1]) ? 3'b010 : 3'b000;
									assign node51 = (inp[7]) ? 3'b010 : 3'b000;
								assign node54 = (inp[7]) ? node56 : 3'b000;
									assign node56 = (inp[11]) ? 3'b000 : node57;
										assign node57 = (inp[10]) ? 3'b000 : 3'b010;
				assign node62 = (inp[7]) ? node186 : node63;
					assign node63 = (inp[9]) ? node149 : node64;
						assign node64 = (inp[10]) ? node120 : node65;
							assign node65 = (inp[4]) ? node89 : node66;
								assign node66 = (inp[11]) ? node78 : node67;
									assign node67 = (inp[2]) ? node69 : 3'b110;
										assign node69 = (inp[5]) ? node75 : node70;
											assign node70 = (inp[1]) ? 3'b110 : node71;
												assign node71 = (inp[8]) ? 3'b100 : 3'b110;
											assign node75 = (inp[1]) ? 3'b100 : 3'b000;
									assign node78 = (inp[5]) ? node84 : node79;
										assign node79 = (inp[8]) ? node81 : 3'b010;
											assign node81 = (inp[1]) ? 3'b110 : 3'b100;
										assign node84 = (inp[8]) ? 3'b010 : node85;
											assign node85 = (inp[1]) ? 3'b100 : 3'b000;
								assign node89 = (inp[11]) ? node101 : node90;
									assign node90 = (inp[8]) ? node96 : node91;
										assign node91 = (inp[1]) ? 3'b100 : node92;
											assign node92 = (inp[5]) ? 3'b000 : 3'b110;
										assign node96 = (inp[5]) ? 3'b110 : node97;
											assign node97 = (inp[1]) ? 3'b010 : 3'b000;
									assign node101 = (inp[2]) ? node115 : node102;
										assign node102 = (inp[1]) ? node108 : node103;
											assign node103 = (inp[8]) ? 3'b000 : node104;
												assign node104 = (inp[5]) ? 3'b000 : 3'b110;
											assign node108 = (inp[8]) ? node112 : node109;
												assign node109 = (inp[5]) ? 3'b000 : 3'b100;
												assign node112 = (inp[5]) ? 3'b100 : 3'b000;
										assign node115 = (inp[5]) ? node117 : 3'b100;
											assign node117 = (inp[8]) ? 3'b100 : 3'b000;
							assign node120 = (inp[4]) ? node140 : node121;
								assign node121 = (inp[11]) ? node129 : node122;
									assign node122 = (inp[1]) ? node124 : 3'b000;
										assign node124 = (inp[5]) ? node126 : 3'b010;
											assign node126 = (inp[8]) ? 3'b010 : 3'b100;
									assign node129 = (inp[8]) ? node135 : node130;
										assign node130 = (inp[5]) ? node132 : 3'b100;
											assign node132 = (inp[1]) ? 3'b100 : 3'b000;
										assign node135 = (inp[5]) ? 3'b100 : node136;
											assign node136 = (inp[1]) ? 3'b010 : 3'b000;
								assign node140 = (inp[8]) ? node142 : 3'b000;
									assign node142 = (inp[5]) ? 3'b000 : node143;
										assign node143 = (inp[2]) ? node145 : 3'b000;
											assign node145 = (inp[11]) ? 3'b000 : 3'b100;
						assign node149 = (inp[5]) ? node175 : node150;
							assign node150 = (inp[8]) ? node158 : node151;
								assign node151 = (inp[1]) ? node153 : 3'b000;
									assign node153 = (inp[10]) ? 3'b000 : node154;
										assign node154 = (inp[4]) ? 3'b000 : 3'b100;
								assign node158 = (inp[2]) ? node164 : node159;
									assign node159 = (inp[4]) ? 3'b000 : node160;
										assign node160 = (inp[10]) ? 3'b000 : 3'b100;
									assign node164 = (inp[10]) ? node172 : node165;
										assign node165 = (inp[1]) ? node167 : 3'b100;
											assign node167 = (inp[4]) ? node169 : 3'b100;
												assign node169 = (inp[11]) ? 3'b100 : 3'b000;
										assign node172 = (inp[11]) ? 3'b000 : 3'b100;
							assign node175 = (inp[8]) ? node177 : 3'b000;
								assign node177 = (inp[10]) ? 3'b000 : node178;
									assign node178 = (inp[4]) ? 3'b000 : node179;
										assign node179 = (inp[1]) ? node181 : 3'b000;
											assign node181 = (inp[11]) ? 3'b000 : 3'b100;
					assign node186 = (inp[4]) ? node280 : node187;
						assign node187 = (inp[10]) ? node221 : node188;
							assign node188 = (inp[9]) ? node210 : node189;
								assign node189 = (inp[5]) ? node201 : node190;
									assign node190 = (inp[8]) ? node196 : node191;
										assign node191 = (inp[11]) ? node193 : 3'b001;
											assign node193 = (inp[1]) ? 3'b001 : 3'b000;
										assign node196 = (inp[1]) ? node198 : 3'b010;
											assign node198 = (inp[11]) ? 3'b000 : 3'b100;
									assign node201 = (inp[8]) ? node205 : node202;
										assign node202 = (inp[1]) ? 3'b110 : 3'b100;
										assign node205 = (inp[1]) ? 3'b001 : node206;
											assign node206 = (inp[2]) ? 3'b001 : 3'b000;
								assign node210 = (inp[5]) ? node218 : node211;
									assign node211 = (inp[8]) ? node213 : 3'b010;
										assign node213 = (inp[1]) ? node215 : 3'b000;
											assign node215 = (inp[11]) ? 3'b010 : 3'b110;
									assign node218 = (inp[8]) ? 3'b010 : 3'b100;
							assign node221 = (inp[8]) ? node241 : node222;
								assign node222 = (inp[5]) ? node236 : node223;
									assign node223 = (inp[11]) ? node231 : node224;
										assign node224 = (inp[1]) ? node228 : node225;
											assign node225 = (inp[9]) ? 3'b110 : 3'b100;
											assign node228 = (inp[9]) ? 3'b100 : 3'b110;
										assign node231 = (inp[9]) ? 3'b100 : node232;
											assign node232 = (inp[1]) ? 3'b110 : 3'b100;
									assign node236 = (inp[1]) ? node238 : 3'b000;
										assign node238 = (inp[9]) ? 3'b000 : 3'b010;
								assign node241 = (inp[5]) ? node257 : node242;
									assign node242 = (inp[11]) ? node250 : node243;
										assign node243 = (inp[9]) ? node247 : node244;
											assign node244 = (inp[1]) ? 3'b000 : 3'b100;
											assign node247 = (inp[1]) ? 3'b010 : 3'b110;
										assign node250 = (inp[9]) ? node254 : node251;
											assign node251 = (inp[1]) ? 3'b110 : 3'b100;
											assign node254 = (inp[1]) ? 3'b100 : 3'b110;
									assign node257 = (inp[2]) ? node273 : node258;
										assign node258 = (inp[11]) ? node266 : node259;
											assign node259 = (inp[1]) ? node263 : node260;
												assign node260 = (inp[9]) ? 3'b110 : 3'b100;
												assign node263 = (inp[9]) ? 3'b100 : 3'b110;
											assign node266 = (inp[1]) ? node270 : node267;
												assign node267 = (inp[9]) ? 3'b110 : 3'b100;
												assign node270 = (inp[9]) ? 3'b100 : 3'b110;
										assign node273 = (inp[1]) ? node277 : node274;
											assign node274 = (inp[9]) ? 3'b110 : 3'b100;
											assign node277 = (inp[9]) ? 3'b100 : 3'b110;
						assign node280 = (inp[9]) ? node332 : node281;
							assign node281 = (inp[1]) ? node311 : node282;
								assign node282 = (inp[11]) ? node300 : node283;
									assign node283 = (inp[10]) ? node293 : node284;
										assign node284 = (inp[8]) ? node288 : node285;
											assign node285 = (inp[2]) ? 3'b111 : 3'b001;
											assign node288 = (inp[5]) ? 3'b001 : node289;
												assign node289 = (inp[2]) ? 3'b000 : 3'b100;
										assign node293 = (inp[8]) ? node297 : node294;
											assign node294 = (inp[2]) ? 3'b100 : 3'b010;
											assign node297 = (inp[5]) ? 3'b010 : 3'b000;
									assign node300 = (inp[8]) ? node308 : node301;
										assign node301 = (inp[5]) ? node303 : 3'b010;
											assign node303 = (inp[2]) ? node305 : 3'b000;
												assign node305 = (inp[10]) ? 3'b000 : 3'b100;
										assign node308 = (inp[5]) ? 3'b010 : 3'b110;
								assign node311 = (inp[10]) ? node323 : node312;
									assign node312 = (inp[5]) ? node316 : node313;
										assign node313 = (inp[8]) ? 3'b110 : 3'b010;
										assign node316 = (inp[2]) ? node318 : 3'b010;
											assign node318 = (inp[11]) ? 3'b010 : node319;
												assign node319 = (inp[8]) ? 3'b110 : 3'b010;
									assign node323 = (inp[5]) ? node325 : 3'b010;
										assign node325 = (inp[8]) ? node329 : node326;
											assign node326 = (inp[2]) ? 3'b100 : 3'b000;
											assign node329 = (inp[11]) ? 3'b000 : 3'b010;
							assign node332 = (inp[10]) ? node350 : node333;
								assign node333 = (inp[11]) ? node343 : node334;
									assign node334 = (inp[8]) ? node338 : node335;
										assign node335 = (inp[5]) ? 3'b000 : 3'b100;
										assign node338 = (inp[1]) ? 3'b100 : node339;
											assign node339 = (inp[5]) ? 3'b100 : 3'b010;
									assign node343 = (inp[2]) ? 3'b000 : node344;
										assign node344 = (inp[8]) ? node346 : 3'b000;
											assign node346 = (inp[5]) ? 3'b000 : 3'b100;
								assign node350 = (inp[1]) ? node356 : node351;
									assign node351 = (inp[5]) ? 3'b000 : node352;
										assign node352 = (inp[11]) ? 3'b000 : 3'b010;
									assign node356 = (inp[8]) ? 3'b000 : node357;
										assign node357 = (inp[2]) ? node359 : 3'b000;
											assign node359 = (inp[11]) ? 3'b000 : node360;
												assign node360 = (inp[5]) ? 3'b100 : 3'b000;
			assign node365 = (inp[7]) ? node399 : node366;
				assign node366 = (inp[4]) ? 3'b000 : node367;
					assign node367 = (inp[5]) ? 3'b000 : node368;
						assign node368 = (inp[9]) ? 3'b000 : node369;
							assign node369 = (inp[11]) ? node387 : node370;
								assign node370 = (inp[10]) ? node380 : node371;
									assign node371 = (inp[8]) ? node377 : node372;
										assign node372 = (inp[0]) ? 3'b000 : node373;
											assign node373 = (inp[1]) ? 3'b100 : 3'b000;
										assign node377 = (inp[0]) ? 3'b100 : 3'b000;
									assign node380 = (inp[1]) ? node382 : 3'b000;
										assign node382 = (inp[2]) ? node384 : 3'b000;
											assign node384 = (inp[8]) ? 3'b000 : 3'b100;
								assign node387 = (inp[10]) ? 3'b000 : node388;
									assign node388 = (inp[8]) ? 3'b000 : node389;
										assign node389 = (inp[0]) ? 3'b000 : node390;
											assign node390 = (inp[1]) ? 3'b100 : 3'b000;
				assign node399 = (inp[9]) ? node501 : node400;
					assign node400 = (inp[8]) ? node446 : node401;
						assign node401 = (inp[10]) ? node433 : node402;
							assign node402 = (inp[0]) ? node426 : node403;
								assign node403 = (inp[11]) ? node419 : node404;
									assign node404 = (inp[4]) ? node412 : node405;
										assign node405 = (inp[2]) ? node407 : 3'b010;
											assign node407 = (inp[1]) ? node409 : 3'b010;
												assign node409 = (inp[5]) ? 3'b110 : 3'b010;
										assign node412 = (inp[1]) ? node416 : node413;
											assign node413 = (inp[5]) ? 3'b010 : 3'b000;
											assign node416 = (inp[5]) ? 3'b100 : 3'b010;
									assign node419 = (inp[1]) ? node421 : 3'b000;
										assign node421 = (inp[4]) ? 3'b000 : node422;
											assign node422 = (inp[5]) ? 3'b110 : 3'b010;
								assign node426 = (inp[5]) ? 3'b000 : node427;
									assign node427 = (inp[4]) ? node429 : 3'b100;
										assign node429 = (inp[11]) ? 3'b000 : 3'b100;
							assign node433 = (inp[4]) ? 3'b000 : node434;
								assign node434 = (inp[5]) ? node440 : node435;
									assign node435 = (inp[1]) ? node437 : 3'b000;
										assign node437 = (inp[0]) ? 3'b000 : 3'b010;
									assign node440 = (inp[11]) ? 3'b000 : node441;
										assign node441 = (inp[1]) ? 3'b100 : 3'b000;
						assign node446 = (inp[0]) ? node472 : node447;
							assign node447 = (inp[5]) ? node449 : 3'b100;
								assign node449 = (inp[1]) ? node457 : node450;
									assign node450 = (inp[10]) ? node454 : node451;
										assign node451 = (inp[11]) ? 3'b100 : 3'b000;
										assign node454 = (inp[11]) ? 3'b000 : 3'b100;
									assign node457 = (inp[4]) ? node465 : node458;
										assign node458 = (inp[11]) ? node462 : node459;
											assign node459 = (inp[10]) ? 3'b110 : 3'b010;
											assign node462 = (inp[10]) ? 3'b010 : 3'b110;
										assign node465 = (inp[11]) ? node469 : node466;
											assign node466 = (inp[10]) ? 3'b100 : 3'b010;
											assign node469 = (inp[10]) ? 3'b000 : 3'b100;
							assign node472 = (inp[4]) ? node494 : node473;
								assign node473 = (inp[1]) ? node481 : node474;
									assign node474 = (inp[10]) ? 3'b000 : node475;
										assign node475 = (inp[5]) ? node477 : 3'b100;
											assign node477 = (inp[11]) ? 3'b000 : 3'b100;
									assign node481 = (inp[11]) ? node489 : node482;
										assign node482 = (inp[10]) ? node486 : node483;
											assign node483 = (inp[5]) ? 3'b100 : 3'b010;
											assign node486 = (inp[5]) ? 3'b000 : 3'b100;
										assign node489 = (inp[5]) ? node491 : 3'b100;
											assign node491 = (inp[10]) ? 3'b000 : 3'b100;
								assign node494 = (inp[10]) ? 3'b000 : node495;
									assign node495 = (inp[1]) ? 3'b000 : node496;
										assign node496 = (inp[5]) ? 3'b000 : 3'b100;
					assign node501 = (inp[0]) ? node535 : node502;
						assign node502 = (inp[5]) ? 3'b000 : node503;
							assign node503 = (inp[8]) ? node505 : 3'b000;
								assign node505 = (inp[11]) ? node517 : node506;
									assign node506 = (inp[4]) ? node512 : node507;
										assign node507 = (inp[10]) ? node509 : 3'b100;
											assign node509 = (inp[1]) ? 3'b100 : 3'b000;
										assign node512 = (inp[10]) ? 3'b100 : node513;
											assign node513 = (inp[1]) ? 3'b000 : 3'b100;
									assign node517 = (inp[1]) ? node521 : node518;
										assign node518 = (inp[10]) ? 3'b000 : 3'b100;
										assign node521 = (inp[2]) ? node527 : node522;
											assign node522 = (inp[10]) ? node524 : 3'b000;
												assign node524 = (inp[4]) ? 3'b100 : 3'b000;
											assign node527 = (inp[4]) ? node531 : node528;
												assign node528 = (inp[10]) ? 3'b000 : 3'b100;
												assign node531 = (inp[10]) ? 3'b100 : 3'b000;
						assign node535 = (inp[11]) ? 3'b000 : node536;
							assign node536 = (inp[10]) ? 3'b000 : node537;
								assign node537 = (inp[4]) ? 3'b000 : node538;
									assign node538 = (inp[5]) ? 3'b000 : node539;
										assign node539 = (inp[8]) ? 3'b010 : 3'b000;
		assign node546 = (inp[3]) ? node876 : node547;
			assign node547 = (inp[0]) ? node645 : node548;
				assign node548 = (inp[7]) ? node558 : node549;
					assign node549 = (inp[8]) ? 3'b001 : node550;
						assign node550 = (inp[5]) ? node552 : 3'b001;
							assign node552 = (inp[10]) ? node554 : 3'b000;
								assign node554 = (inp[9]) ? 3'b000 : 3'b001;
					assign node558 = (inp[5]) ? node616 : node559;
						assign node559 = (inp[9]) ? node569 : node560;
							assign node560 = (inp[1]) ? node562 : 3'b111;
								assign node562 = (inp[8]) ? 3'b111 : node563;
									assign node563 = (inp[10]) ? node565 : 3'b111;
										assign node565 = (inp[2]) ? 3'b111 : 3'b011;
							assign node569 = (inp[4]) ? node589 : node570;
								assign node570 = (inp[10]) ? node576 : node571;
									assign node571 = (inp[1]) ? 3'b111 : node572;
										assign node572 = (inp[11]) ? 3'b111 : 3'b011;
									assign node576 = (inp[11]) ? node584 : node577;
										assign node577 = (inp[1]) ? node581 : node578;
											assign node578 = (inp[8]) ? 3'b011 : 3'b111;
											assign node581 = (inp[8]) ? 3'b111 : 3'b011;
										assign node584 = (inp[8]) ? 3'b011 : node585;
											assign node585 = (inp[1]) ? 3'b011 : 3'b111;
								assign node589 = (inp[1]) ? node601 : node590;
									assign node590 = (inp[10]) ? node596 : node591;
										assign node591 = (inp[8]) ? 3'b111 : node592;
											assign node592 = (inp[11]) ? 3'b011 : 3'b111;
										assign node596 = (inp[8]) ? 3'b011 : node597;
											assign node597 = (inp[11]) ? 3'b101 : 3'b111;
									assign node601 = (inp[11]) ? node607 : node602;
										assign node602 = (inp[10]) ? 3'b101 : node603;
											assign node603 = (inp[2]) ? 3'b111 : 3'b011;
										assign node607 = (inp[2]) ? node609 : 3'b101;
											assign node609 = (inp[8]) ? node613 : node610;
												assign node610 = (inp[10]) ? 3'b001 : 3'b101;
												assign node613 = (inp[10]) ? 3'b101 : 3'b001;
						assign node616 = (inp[8]) ? node618 : 3'b000;
							assign node618 = (inp[1]) ? node632 : node619;
								assign node619 = (inp[9]) ? node621 : 3'b111;
									assign node621 = (inp[10]) ? node629 : node622;
										assign node622 = (inp[11]) ? node626 : node623;
											assign node623 = (inp[4]) ? 3'b111 : 3'b011;
											assign node626 = (inp[4]) ? 3'b011 : 3'b111;
										assign node629 = (inp[4]) ? 3'b101 : 3'b111;
								assign node632 = (inp[10]) ? node640 : node633;
									assign node633 = (inp[2]) ? 3'b111 : node634;
										assign node634 = (inp[4]) ? node636 : 3'b111;
											assign node636 = (inp[9]) ? 3'b101 : 3'b111;
									assign node640 = (inp[11]) ? 3'b011 : node641;
										assign node641 = (inp[9]) ? 3'b011 : 3'b111;
				assign node645 = (inp[10]) ? node775 : node646;
					assign node646 = (inp[4]) ? node700 : node647;
						assign node647 = (inp[8]) ? node675 : node648;
							assign node648 = (inp[7]) ? node660 : node649;
								assign node649 = (inp[5]) ? node653 : node650;
									assign node650 = (inp[11]) ? 3'b111 : 3'b011;
									assign node653 = (inp[9]) ? 3'b101 : node654;
										assign node654 = (inp[11]) ? 3'b001 : node655;
											assign node655 = (inp[1]) ? 3'b101 : 3'b001;
								assign node660 = (inp[1]) ? node666 : node661;
									assign node661 = (inp[9]) ? node663 : 3'b111;
										assign node663 = (inp[5]) ? 3'b111 : 3'b011;
									assign node666 = (inp[9]) ? node670 : node667;
										assign node667 = (inp[5]) ? 3'b011 : 3'b111;
										assign node670 = (inp[5]) ? 3'b111 : node671;
											assign node671 = (inp[11]) ? 3'b110 : 3'b101;
							assign node675 = (inp[11]) ? node689 : node676;
								assign node676 = (inp[5]) ? node682 : node677;
									assign node677 = (inp[1]) ? node679 : 3'b111;
										assign node679 = (inp[7]) ? 3'b011 : 3'b111;
									assign node682 = (inp[7]) ? node684 : 3'b011;
										assign node684 = (inp[9]) ? node686 : 3'b111;
											assign node686 = (inp[2]) ? 3'b101 : 3'b011;
								assign node689 = (inp[7]) ? node691 : 3'b111;
									assign node691 = (inp[9]) ? node695 : node692;
										assign node692 = (inp[1]) ? 3'b011 : 3'b111;
										assign node695 = (inp[5]) ? node697 : 3'b111;
											assign node697 = (inp[1]) ? 3'b110 : 3'b011;
						assign node700 = (inp[11]) ? node736 : node701;
							assign node701 = (inp[7]) ? node717 : node702;
								assign node702 = (inp[5]) ? node706 : node703;
									assign node703 = (inp[8]) ? 3'b101 : 3'b001;
									assign node706 = (inp[8]) ? 3'b001 : node707;
										assign node707 = (inp[2]) ? node713 : node708;
											assign node708 = (inp[1]) ? 3'b100 : node709;
												assign node709 = (inp[9]) ? 3'b100 : 3'b000;
											assign node713 = (inp[9]) ? 3'b110 : 3'b010;
								assign node717 = (inp[9]) ? node733 : node718;
									assign node718 = (inp[1]) ? node726 : node719;
										assign node719 = (inp[5]) ? node721 : 3'b111;
											assign node721 = (inp[8]) ? 3'b111 : node722;
												assign node722 = (inp[2]) ? 3'b001 : 3'b011;
										assign node726 = (inp[2]) ? 3'b101 : node727;
											assign node727 = (inp[5]) ? node729 : 3'b101;
												assign node729 = (inp[8]) ? 3'b101 : 3'b111;
									assign node733 = (inp[5]) ? 3'b101 : 3'b001;
							assign node736 = (inp[7]) ? node748 : node737;
								assign node737 = (inp[5]) ? node741 : node738;
									assign node738 = (inp[8]) ? 3'b111 : 3'b011;
									assign node741 = (inp[8]) ? 3'b011 : node742;
										assign node742 = (inp[9]) ? 3'b110 : node743;
											assign node743 = (inp[1]) ? 3'b110 : 3'b010;
								assign node748 = (inp[1]) ? node766 : node749;
									assign node749 = (inp[9]) ? node759 : node750;
										assign node750 = (inp[2]) ? 3'b101 : node751;
											assign node751 = (inp[5]) ? node755 : node752;
												assign node752 = (inp[8]) ? 3'b111 : 3'b011;
												assign node755 = (inp[8]) ? 3'b011 : 3'b101;
										assign node759 = (inp[8]) ? node763 : node760;
											assign node760 = (inp[5]) ? 3'b101 : 3'b001;
											assign node763 = (inp[5]) ? 3'b001 : 3'b101;
									assign node766 = (inp[9]) ? node768 : 3'b101;
										assign node768 = (inp[2]) ? node770 : 3'b110;
											assign node770 = (inp[8]) ? 3'b110 : node771;
												assign node771 = (inp[5]) ? 3'b101 : 3'b110;
					assign node775 = (inp[7]) ? node799 : node776;
						assign node776 = (inp[4]) ? node792 : node777;
							assign node777 = (inp[5]) ? node783 : node778;
								assign node778 = (inp[8]) ? 3'b110 : node779;
									assign node779 = (inp[11]) ? 3'b010 : 3'b110;
								assign node783 = (inp[8]) ? node789 : node784;
									assign node784 = (inp[9]) ? 3'b100 : node785;
										assign node785 = (inp[1]) ? 3'b000 : 3'b100;
									assign node789 = (inp[11]) ? 3'b010 : 3'b110;
							assign node792 = (inp[11]) ? node794 : 3'b110;
								assign node794 = (inp[8]) ? 3'b100 : node795;
									assign node795 = (inp[5]) ? 3'b110 : 3'b100;
						assign node799 = (inp[5]) ? node841 : node800;
							assign node800 = (inp[1]) ? node822 : node801;
								assign node801 = (inp[9]) ? node811 : node802;
									assign node802 = (inp[4]) ? node804 : 3'b111;
										assign node804 = (inp[2]) ? node806 : 3'b101;
											assign node806 = (inp[11]) ? 3'b011 : node807;
												assign node807 = (inp[8]) ? 3'b111 : 3'b011;
									assign node811 = (inp[8]) ? node817 : node812;
										assign node812 = (inp[4]) ? node814 : 3'b101;
											assign node814 = (inp[11]) ? 3'b110 : 3'b001;
										assign node817 = (inp[4]) ? node819 : 3'b011;
											assign node819 = (inp[11]) ? 3'b001 : 3'b101;
								assign node822 = (inp[9]) ? node830 : node823;
									assign node823 = (inp[11]) ? 3'b101 : node824;
										assign node824 = (inp[4]) ? node826 : 3'b011;
											assign node826 = (inp[8]) ? 3'b101 : 3'b001;
									assign node830 = (inp[8]) ? node834 : node831;
										assign node831 = (inp[4]) ? 3'b010 : 3'b110;
										assign node834 = (inp[4]) ? node838 : node835;
											assign node835 = (inp[11]) ? 3'b001 : 3'b101;
											assign node838 = (inp[11]) ? 3'b110 : 3'b100;
							assign node841 = (inp[4]) ? node859 : node842;
								assign node842 = (inp[8]) ? node848 : node843;
									assign node843 = (inp[1]) ? node845 : 3'b110;
										assign node845 = (inp[9]) ? 3'b110 : 3'b010;
									assign node848 = (inp[9]) ? node856 : node849;
										assign node849 = (inp[11]) ? node853 : node850;
											assign node850 = (inp[1]) ? 3'b011 : 3'b111;
											assign node853 = (inp[1]) ? 3'b101 : 3'b111;
										assign node856 = (inp[1]) ? 3'b110 : 3'b101;
								assign node859 = (inp[8]) ? node865 : node860;
									assign node860 = (inp[1]) ? node862 : 3'b100;
										assign node862 = (inp[9]) ? 3'b100 : 3'b000;
									assign node865 = (inp[9]) ? node869 : node866;
										assign node866 = (inp[2]) ? 3'b101 : 3'b001;
										assign node869 = (inp[1]) ? node873 : node870;
											assign node870 = (inp[11]) ? 3'b110 : 3'b001;
											assign node873 = (inp[11]) ? 3'b010 : 3'b110;
			assign node876 = (inp[7]) ? node1076 : node877;
				assign node877 = (inp[0]) ? node933 : node878;
					assign node878 = (inp[10]) ? node906 : node879;
						assign node879 = (inp[11]) ? node893 : node880;
							assign node880 = (inp[5]) ? node884 : node881;
								assign node881 = (inp[8]) ? 3'b000 : 3'b110;
								assign node884 = (inp[8]) ? 3'b110 : node885;
									assign node885 = (inp[9]) ? 3'b000 : node886;
										assign node886 = (inp[1]) ? node888 : 3'b000;
											assign node888 = (inp[2]) ? 3'b010 : 3'b000;
							assign node893 = (inp[8]) ? node903 : node894;
								assign node894 = (inp[5]) ? node896 : 3'b010;
									assign node896 = (inp[1]) ? node898 : 3'b000;
										assign node898 = (inp[4]) ? node900 : 3'b000;
											assign node900 = (inp[9]) ? 3'b000 : 3'b010;
								assign node903 = (inp[5]) ? 3'b010 : 3'b000;
						assign node906 = (inp[11]) ? node922 : node907;
							assign node907 = (inp[8]) ? node919 : node908;
								assign node908 = (inp[5]) ? node910 : 3'b010;
									assign node910 = (inp[9]) ? 3'b100 : node911;
										assign node911 = (inp[1]) ? node913 : 3'b110;
											assign node913 = (inp[4]) ? node915 : 3'b100;
												assign node915 = (inp[2]) ? 3'b100 : 3'b110;
								assign node919 = (inp[5]) ? 3'b010 : 3'b000;
							assign node922 = (inp[5]) ? node926 : node923;
								assign node923 = (inp[8]) ? 3'b000 : 3'b100;
								assign node926 = (inp[8]) ? 3'b100 : node927;
									assign node927 = (inp[1]) ? 3'b100 : node928;
										assign node928 = (inp[9]) ? 3'b100 : 3'b110;
					assign node933 = (inp[9]) ? node1051 : node934;
						assign node934 = (inp[10]) ? node994 : node935;
							assign node935 = (inp[4]) ? node965 : node936;
								assign node936 = (inp[2]) ? node954 : node937;
									assign node937 = (inp[11]) ? node945 : node938;
										assign node938 = (inp[8]) ? node940 : 3'b010;
											assign node940 = (inp[5]) ? node942 : 3'b100;
												assign node942 = (inp[1]) ? 3'b110 : 3'b010;
										assign node945 = (inp[8]) ? node949 : node946;
											assign node946 = (inp[5]) ? 3'b100 : 3'b010;
											assign node949 = (inp[5]) ? 3'b010 : node950;
												assign node950 = (inp[1]) ? 3'b110 : 3'b100;
									assign node954 = (inp[11]) ? 3'b010 : node955;
										assign node955 = (inp[5]) ? node957 : 3'b110;
											assign node957 = (inp[8]) ? node961 : node958;
												assign node958 = (inp[1]) ? 3'b010 : 3'b110;
												assign node961 = (inp[1]) ? 3'b110 : 3'b010;
								assign node965 = (inp[11]) ? node975 : node966;
									assign node966 = (inp[8]) ? 3'b010 : node967;
										assign node967 = (inp[1]) ? node971 : node968;
											assign node968 = (inp[5]) ? 3'b100 : 3'b010;
											assign node971 = (inp[5]) ? 3'b000 : 3'b100;
									assign node975 = (inp[1]) ? node985 : node976;
										assign node976 = (inp[2]) ? node980 : node977;
											assign node977 = (inp[8]) ? 3'b010 : 3'b100;
											assign node980 = (inp[5]) ? 3'b100 : node981;
												assign node981 = (inp[8]) ? 3'b100 : 3'b010;
										assign node985 = (inp[2]) ? node991 : node986;
											assign node986 = (inp[5]) ? 3'b100 : node987;
												assign node987 = (inp[8]) ? 3'b000 : 3'b100;
											assign node991 = (inp[8]) ? 3'b100 : 3'b000;
							assign node994 = (inp[1]) ? node1024 : node995;
								assign node995 = (inp[4]) ? node1011 : node996;
									assign node996 = (inp[2]) ? node1004 : node997;
										assign node997 = (inp[5]) ? node1001 : node998;
											assign node998 = (inp[8]) ? 3'b000 : 3'b100;
											assign node1001 = (inp[8]) ? 3'b100 : 3'b000;
										assign node1004 = (inp[5]) ? node1008 : node1005;
											assign node1005 = (inp[8]) ? 3'b000 : 3'b100;
											assign node1008 = (inp[8]) ? 3'b100 : 3'b000;
									assign node1011 = (inp[2]) ? node1019 : node1012;
										assign node1012 = (inp[8]) ? node1016 : node1013;
											assign node1013 = (inp[5]) ? 3'b000 : 3'b100;
											assign node1016 = (inp[5]) ? 3'b100 : 3'b000;
										assign node1019 = (inp[8]) ? 3'b100 : node1020;
											assign node1020 = (inp[5]) ? 3'b000 : 3'b100;
								assign node1024 = (inp[4]) ? node1038 : node1025;
									assign node1025 = (inp[11]) ? node1031 : node1026;
										assign node1026 = (inp[5]) ? node1028 : 3'b010;
											assign node1028 = (inp[2]) ? 3'b100 : 3'b010;
										assign node1031 = (inp[5]) ? node1035 : node1032;
											assign node1032 = (inp[8]) ? 3'b010 : 3'b000;
											assign node1035 = (inp[8]) ? 3'b000 : 3'b100;
									assign node1038 = (inp[11]) ? 3'b000 : node1039;
										assign node1039 = (inp[5]) ? node1045 : node1040;
											assign node1040 = (inp[2]) ? 3'b100 : node1041;
												assign node1041 = (inp[8]) ? 3'b000 : 3'b100;
											assign node1045 = (inp[8]) ? node1047 : 3'b000;
												assign node1047 = (inp[2]) ? 3'b000 : 3'b100;
						assign node1051 = (inp[8]) ? node1061 : node1052;
							assign node1052 = (inp[5]) ? node1054 : 3'b000;
								assign node1054 = (inp[4]) ? 3'b000 : node1055;
									assign node1055 = (inp[10]) ? 3'b000 : node1056;
										assign node1056 = (inp[11]) ? 3'b000 : 3'b010;
							assign node1061 = (inp[5]) ? 3'b000 : node1062;
								assign node1062 = (inp[10]) ? node1070 : node1063;
									assign node1063 = (inp[4]) ? node1065 : 3'b100;
										assign node1065 = (inp[2]) ? node1067 : 3'b000;
											assign node1067 = (inp[11]) ? 3'b100 : 3'b000;
									assign node1070 = (inp[4]) ? node1072 : 3'b000;
										assign node1072 = (inp[11]) ? 3'b000 : 3'b100;
				assign node1076 = (inp[0]) ? node1252 : node1077;
					assign node1077 = (inp[9]) ? node1173 : node1078;
						assign node1078 = (inp[4]) ? node1122 : node1079;
							assign node1079 = (inp[1]) ? node1097 : node1080;
								assign node1080 = (inp[10]) ? node1088 : node1081;
									assign node1081 = (inp[5]) ? node1083 : 3'b111;
										assign node1083 = (inp[8]) ? 3'b111 : node1084;
											assign node1084 = (inp[11]) ? 3'b110 : 3'b000;
									assign node1088 = (inp[5]) ? node1094 : node1089;
										assign node1089 = (inp[11]) ? 3'b011 : node1090;
											assign node1090 = (inp[8]) ? 3'b111 : 3'b011;
										assign node1094 = (inp[8]) ? 3'b011 : 3'b110;
								assign node1097 = (inp[10]) ? node1109 : node1098;
									assign node1098 = (inp[5]) ? node1104 : node1099;
										assign node1099 = (inp[8]) ? node1101 : 3'b011;
											assign node1101 = (inp[11]) ? 3'b011 : 3'b111;
										assign node1104 = (inp[11]) ? 3'b111 : node1105;
											assign node1105 = (inp[8]) ? 3'b011 : 3'b001;
									assign node1109 = (inp[11]) ? node1117 : node1110;
										assign node1110 = (inp[8]) ? node1114 : node1111;
											assign node1111 = (inp[5]) ? 3'b111 : 3'b101;
											assign node1114 = (inp[5]) ? 3'b101 : 3'b011;
										assign node1117 = (inp[8]) ? 3'b101 : node1118;
											assign node1118 = (inp[5]) ? 3'b111 : 3'b101;
							assign node1122 = (inp[10]) ? node1152 : node1123;
								assign node1123 = (inp[11]) ? node1141 : node1124;
									assign node1124 = (inp[8]) ? node1134 : node1125;
										assign node1125 = (inp[5]) ? node1131 : node1126;
											assign node1126 = (inp[1]) ? node1128 : 3'b101;
												assign node1128 = (inp[2]) ? 3'b001 : 3'b101;
											assign node1131 = (inp[1]) ? 3'b001 : 3'b000;
										assign node1134 = (inp[5]) ? node1136 : 3'b011;
											assign node1136 = (inp[2]) ? node1138 : 3'b101;
												assign node1138 = (inp[1]) ? 3'b001 : 3'b101;
									assign node1141 = (inp[8]) ? node1147 : node1142;
										assign node1142 = (inp[5]) ? 3'b110 : node1143;
											assign node1143 = (inp[1]) ? 3'b001 : 3'b101;
										assign node1147 = (inp[5]) ? node1149 : 3'b111;
											assign node1149 = (inp[1]) ? 3'b001 : 3'b101;
								assign node1152 = (inp[5]) ? node1164 : node1153;
									assign node1153 = (inp[1]) ? node1157 : node1154;
										assign node1154 = (inp[11]) ? 3'b001 : 3'b101;
										assign node1157 = (inp[8]) ? 3'b101 : node1158;
											assign node1158 = (inp[11]) ? 3'b110 : node1159;
												assign node1159 = (inp[2]) ? 3'b110 : 3'b001;
									assign node1164 = (inp[8]) ? node1166 : 3'b110;
										assign node1166 = (inp[2]) ? 3'b110 : node1167;
											assign node1167 = (inp[1]) ? 3'b001 : node1168;
												assign node1168 = (inp[11]) ? 3'b001 : 3'b101;
						assign node1173 = (inp[4]) ? node1207 : node1174;
							assign node1174 = (inp[8]) ? node1188 : node1175;
								assign node1175 = (inp[5]) ? node1183 : node1176;
									assign node1176 = (inp[10]) ? node1180 : node1177;
										assign node1177 = (inp[1]) ? 3'b001 : 3'b101;
										assign node1180 = (inp[1]) ? 3'b110 : 3'b001;
									assign node1183 = (inp[11]) ? 3'b110 : node1184;
										assign node1184 = (inp[10]) ? 3'b110 : 3'b000;
								assign node1188 = (inp[10]) ? node1198 : node1189;
									assign node1189 = (inp[1]) ? node1195 : node1190;
										assign node1190 = (inp[5]) ? 3'b101 : node1191;
											assign node1191 = (inp[11]) ? 3'b101 : 3'b011;
										assign node1195 = (inp[5]) ? 3'b001 : 3'b101;
									assign node1198 = (inp[1]) ? node1204 : node1199;
										assign node1199 = (inp[11]) ? 3'b001 : node1200;
											assign node1200 = (inp[5]) ? 3'b001 : 3'b101;
										assign node1204 = (inp[5]) ? 3'b110 : 3'b001;
							assign node1207 = (inp[10]) ? node1233 : node1208;
								assign node1208 = (inp[1]) ? node1218 : node1209;
									assign node1209 = (inp[5]) ? node1211 : 3'b001;
										assign node1211 = (inp[11]) ? 3'b110 : node1212;
											assign node1212 = (inp[2]) ? node1214 : 3'b001;
												assign node1214 = (inp[8]) ? 3'b110 : 3'b000;
									assign node1218 = (inp[11]) ? node1226 : node1219;
										assign node1219 = (inp[5]) ? node1221 : 3'b110;
											assign node1221 = (inp[8]) ? node1223 : 3'b000;
												assign node1223 = (inp[2]) ? 3'b010 : 3'b110;
										assign node1226 = (inp[5]) ? node1230 : node1227;
											assign node1227 = (inp[8]) ? 3'b110 : 3'b010;
											assign node1230 = (inp[8]) ? 3'b010 : 3'b110;
								assign node1233 = (inp[5]) ? node1245 : node1234;
									assign node1234 = (inp[1]) ? node1240 : node1235;
										assign node1235 = (inp[8]) ? 3'b110 : node1236;
											assign node1236 = (inp[11]) ? 3'b010 : 3'b110;
										assign node1240 = (inp[8]) ? 3'b010 : node1241;
											assign node1241 = (inp[11]) ? 3'b100 : 3'b010;
									assign node1245 = (inp[8]) ? node1247 : 3'b110;
										assign node1247 = (inp[1]) ? 3'b100 : node1248;
											assign node1248 = (inp[11]) ? 3'b010 : 3'b110;
					assign node1252 = (inp[9]) ? node1344 : node1253;
						assign node1253 = (inp[4]) ? node1289 : node1254;
							assign node1254 = (inp[8]) ? node1270 : node1255;
								assign node1255 = (inp[5]) ? node1263 : node1256;
									assign node1256 = (inp[10]) ? node1260 : node1257;
										assign node1257 = (inp[1]) ? 3'b001 : 3'b101;
										assign node1260 = (inp[1]) ? 3'b110 : 3'b001;
									assign node1263 = (inp[1]) ? 3'b110 : node1264;
										assign node1264 = (inp[11]) ? 3'b010 : node1265;
											assign node1265 = (inp[10]) ? 3'b010 : 3'b110;
								assign node1270 = (inp[10]) ? node1280 : node1271;
									assign node1271 = (inp[1]) ? node1275 : node1272;
										assign node1272 = (inp[5]) ? 3'b101 : 3'b011;
										assign node1275 = (inp[11]) ? 3'b001 : node1276;
											assign node1276 = (inp[5]) ? 3'b001 : 3'b101;
									assign node1280 = (inp[1]) ? node1284 : node1281;
										assign node1281 = (inp[5]) ? 3'b001 : 3'b101;
										assign node1284 = (inp[5]) ? 3'b110 : node1285;
											assign node1285 = (inp[11]) ? 3'b110 : 3'b001;
							assign node1289 = (inp[1]) ? node1325 : node1290;
								assign node1290 = (inp[10]) ? node1308 : node1291;
									assign node1291 = (inp[5]) ? node1299 : node1292;
										assign node1292 = (inp[8]) ? node1296 : node1293;
											assign node1293 = (inp[11]) ? 3'b110 : 3'b001;
											assign node1296 = (inp[11]) ? 3'b001 : 3'b101;
										assign node1299 = (inp[8]) ? node1303 : node1300;
											assign node1300 = (inp[11]) ? 3'b010 : 3'b110;
											assign node1303 = (inp[2]) ? 3'b110 : node1304;
												assign node1304 = (inp[11]) ? 3'b110 : 3'b001;
									assign node1308 = (inp[5]) ? node1318 : node1309;
										assign node1309 = (inp[8]) ? node1315 : node1310;
											assign node1310 = (inp[2]) ? 3'b010 : node1311;
												assign node1311 = (inp[11]) ? 3'b010 : 3'b110;
											assign node1315 = (inp[11]) ? 3'b110 : 3'b001;
										assign node1318 = (inp[8]) ? node1320 : 3'b010;
											assign node1320 = (inp[11]) ? 3'b010 : node1321;
												assign node1321 = (inp[2]) ? 3'b010 : 3'b110;
								assign node1325 = (inp[10]) ? node1333 : node1326;
									assign node1326 = (inp[8]) ? 3'b110 : node1327;
										assign node1327 = (inp[11]) ? node1329 : 3'b010;
											assign node1329 = (inp[2]) ? 3'b010 : 3'b110;
									assign node1333 = (inp[5]) ? node1339 : node1334;
										assign node1334 = (inp[8]) ? 3'b010 : node1335;
											assign node1335 = (inp[11]) ? 3'b100 : 3'b010;
										assign node1339 = (inp[11]) ? 3'b100 : node1340;
											assign node1340 = (inp[8]) ? 3'b110 : 3'b100;
						assign node1344 = (inp[4]) ? node1372 : node1345;
							assign node1345 = (inp[5]) ? node1363 : node1346;
								assign node1346 = (inp[8]) ? node1354 : node1347;
									assign node1347 = (inp[10]) ? node1351 : node1348;
										assign node1348 = (inp[1]) ? 3'b010 : 3'b110;
										assign node1351 = (inp[1]) ? 3'b100 : 3'b010;
									assign node1354 = (inp[1]) ? node1358 : node1355;
										assign node1355 = (inp[10]) ? 3'b110 : 3'b001;
										assign node1358 = (inp[11]) ? 3'b010 : node1359;
											assign node1359 = (inp[10]) ? 3'b010 : 3'b110;
								assign node1363 = (inp[8]) ? node1365 : 3'b000;
									assign node1365 = (inp[10]) ? node1369 : node1366;
										assign node1366 = (inp[1]) ? 3'b010 : 3'b110;
										assign node1369 = (inp[1]) ? 3'b100 : 3'b010;
							assign node1372 = (inp[8]) ? node1380 : node1373;
								assign node1373 = (inp[5]) ? 3'b000 : node1374;
									assign node1374 = (inp[1]) ? 3'b000 : node1375;
										assign node1375 = (inp[10]) ? 3'b000 : 3'b100;
								assign node1380 = (inp[1]) ? node1394 : node1381;
									assign node1381 = (inp[10]) ? node1389 : node1382;
										assign node1382 = (inp[5]) ? node1386 : node1383;
											assign node1383 = (inp[2]) ? 3'b011 : 3'b010;
											assign node1386 = (inp[11]) ? 3'b100 : 3'b010;
										assign node1389 = (inp[5]) ? node1391 : 3'b100;
											assign node1391 = (inp[11]) ? 3'b000 : 3'b100;
									assign node1394 = (inp[10]) ? 3'b000 : node1395;
										assign node1395 = (inp[5]) ? node1397 : 3'b100;
											assign node1397 = (inp[2]) ? node1399 : 3'b000;
												assign node1399 = (inp[11]) ? 3'b000 : 3'b100;

endmodule