module dtc_split125_bm75 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node9;
	wire [3-1:0] node12;
	wire [3-1:0] node13;
	wire [3-1:0] node16;
	wire [3-1:0] node19;
	wire [3-1:0] node21;
	wire [3-1:0] node23;
	wire [3-1:0] node26;
	wire [3-1:0] node27;
	wire [3-1:0] node28;
	wire [3-1:0] node29;
	wire [3-1:0] node32;
	wire [3-1:0] node35;
	wire [3-1:0] node36;
	wire [3-1:0] node39;
	wire [3-1:0] node42;
	wire [3-1:0] node43;
	wire [3-1:0] node44;
	wire [3-1:0] node47;
	wire [3-1:0] node50;
	wire [3-1:0] node51;
	wire [3-1:0] node54;
	wire [3-1:0] node57;
	wire [3-1:0] node58;
	wire [3-1:0] node59;
	wire [3-1:0] node60;
	wire [3-1:0] node61;
	wire [3-1:0] node64;
	wire [3-1:0] node67;
	wire [3-1:0] node68;
	wire [3-1:0] node71;
	wire [3-1:0] node74;
	wire [3-1:0] node75;
	wire [3-1:0] node76;
	wire [3-1:0] node79;
	wire [3-1:0] node82;
	wire [3-1:0] node83;
	wire [3-1:0] node86;
	wire [3-1:0] node89;
	wire [3-1:0] node90;
	wire [3-1:0] node91;
	wire [3-1:0] node92;
	wire [3-1:0] node95;
	wire [3-1:0] node98;
	wire [3-1:0] node99;
	wire [3-1:0] node102;
	wire [3-1:0] node105;
	wire [3-1:0] node106;
	wire [3-1:0] node107;
	wire [3-1:0] node110;
	wire [3-1:0] node113;
	wire [3-1:0] node114;
	wire [3-1:0] node117;
	wire [3-1:0] node120;
	wire [3-1:0] node121;
	wire [3-1:0] node122;
	wire [3-1:0] node123;
	wire [3-1:0] node124;
	wire [3-1:0] node125;
	wire [3-1:0] node128;
	wire [3-1:0] node131;
	wire [3-1:0] node132;
	wire [3-1:0] node135;
	wire [3-1:0] node138;
	wire [3-1:0] node139;
	wire [3-1:0] node140;
	wire [3-1:0] node143;
	wire [3-1:0] node146;
	wire [3-1:0] node147;
	wire [3-1:0] node150;
	wire [3-1:0] node153;
	wire [3-1:0] node154;
	wire [3-1:0] node155;
	wire [3-1:0] node157;
	wire [3-1:0] node160;
	wire [3-1:0] node161;
	wire [3-1:0] node164;
	wire [3-1:0] node167;
	wire [3-1:0] node168;
	wire [3-1:0] node169;
	wire [3-1:0] node172;
	wire [3-1:0] node175;
	wire [3-1:0] node176;
	wire [3-1:0] node179;
	wire [3-1:0] node182;
	wire [3-1:0] node183;
	wire [3-1:0] node184;
	wire [3-1:0] node185;
	wire [3-1:0] node186;
	wire [3-1:0] node190;
	wire [3-1:0] node191;
	wire [3-1:0] node195;
	wire [3-1:0] node196;
	wire [3-1:0] node197;
	wire [3-1:0] node200;
	wire [3-1:0] node203;
	wire [3-1:0] node204;
	wire [3-1:0] node207;
	wire [3-1:0] node210;
	wire [3-1:0] node212;
	wire [3-1:0] node214;
	wire [3-1:0] node215;
	wire [3-1:0] node218;

	assign outp = (inp[3]) ? node120 : node1;
		assign node1 = (inp[9]) ? node57 : node2;
			assign node2 = (inp[4]) ? node26 : node3;
				assign node3 = (inp[6]) ? node19 : node4;
					assign node4 = (inp[11]) ? node12 : node5;
						assign node5 = (inp[1]) ? node9 : node6;
							assign node6 = (inp[10]) ? 3'b011 : 3'b111;
							assign node9 = (inp[5]) ? 3'b111 : 3'b111;
						assign node12 = (inp[10]) ? node16 : node13;
							assign node13 = (inp[0]) ? 3'b111 : 3'b011;
							assign node16 = (inp[8]) ? 3'b101 : 3'b101;
					assign node19 = (inp[5]) ? node21 : 3'b111;
						assign node21 = (inp[1]) ? node23 : 3'b111;
							assign node23 = (inp[11]) ? 3'b011 : 3'b111;
				assign node26 = (inp[6]) ? node42 : node27;
					assign node27 = (inp[0]) ? node35 : node28;
						assign node28 = (inp[8]) ? node32 : node29;
							assign node29 = (inp[7]) ? 3'b110 : 3'b110;
							assign node32 = (inp[7]) ? 3'b001 : 3'b010;
						assign node35 = (inp[7]) ? node39 : node36;
							assign node36 = (inp[10]) ? 3'b101 : 3'b001;
							assign node39 = (inp[5]) ? 3'b101 : 3'b101;
					assign node42 = (inp[0]) ? node50 : node43;
						assign node43 = (inp[8]) ? node47 : node44;
							assign node44 = (inp[5]) ? 3'b001 : 3'b011;
							assign node47 = (inp[5]) ? 3'b101 : 3'b101;
						assign node50 = (inp[10]) ? node54 : node51;
							assign node51 = (inp[5]) ? 3'b011 : 3'b111;
							assign node54 = (inp[1]) ? 3'b011 : 3'b001;
			assign node57 = (inp[6]) ? node89 : node58;
				assign node58 = (inp[4]) ? node74 : node59;
					assign node59 = (inp[7]) ? node67 : node60;
						assign node60 = (inp[1]) ? node64 : node61;
							assign node61 = (inp[11]) ? 3'b010 : 3'b100;
							assign node64 = (inp[2]) ? 3'b001 : 3'b110;
						assign node67 = (inp[10]) ? node71 : node68;
							assign node68 = (inp[5]) ? 3'b101 : 3'b001;
							assign node71 = (inp[5]) ? 3'b010 : 3'b001;
					assign node74 = (inp[10]) ? node82 : node75;
						assign node75 = (inp[2]) ? node79 : node76;
							assign node76 = (inp[7]) ? 3'b001 : 3'b010;
							assign node79 = (inp[0]) ? 3'b110 : 3'b010;
						assign node82 = (inp[11]) ? node86 : node83;
							assign node83 = (inp[0]) ? 3'b010 : 3'b100;
							assign node86 = (inp[8]) ? 3'b100 : 3'b000;
				assign node89 = (inp[4]) ? node105 : node90;
					assign node90 = (inp[0]) ? node98 : node91;
						assign node91 = (inp[2]) ? node95 : node92;
							assign node92 = (inp[10]) ? 3'b001 : 3'b101;
							assign node95 = (inp[1]) ? 3'b011 : 3'b001;
						assign node98 = (inp[8]) ? node102 : node99;
							assign node99 = (inp[7]) ? 3'b111 : 3'b011;
							assign node102 = (inp[10]) ? 3'b101 : 3'b111;
					assign node105 = (inp[0]) ? node113 : node106;
						assign node106 = (inp[1]) ? node110 : node107;
							assign node107 = (inp[7]) ? 3'b010 : 3'b110;
							assign node110 = (inp[8]) ? 3'b101 : 3'b001;
						assign node113 = (inp[2]) ? node117 : node114;
							assign node114 = (inp[11]) ? 3'b001 : 3'b001;
							assign node117 = (inp[1]) ? 3'b001 : 3'b101;
		assign node120 = (inp[4]) ? node182 : node121;
			assign node121 = (inp[9]) ? node153 : node122;
				assign node122 = (inp[6]) ? node138 : node123;
					assign node123 = (inp[10]) ? node131 : node124;
						assign node124 = (inp[0]) ? node128 : node125;
							assign node125 = (inp[7]) ? 3'b010 : 3'b010;
							assign node128 = (inp[5]) ? 3'b110 : 3'b001;
						assign node131 = (inp[8]) ? node135 : node132;
							assign node132 = (inp[0]) ? 3'b010 : 3'b000;
							assign node135 = (inp[0]) ? 3'b010 : 3'b100;
					assign node138 = (inp[11]) ? node146 : node139;
						assign node139 = (inp[0]) ? node143 : node140;
							assign node140 = (inp[10]) ? 3'b110 : 3'b001;
							assign node143 = (inp[7]) ? 3'b011 : 3'b001;
						assign node146 = (inp[1]) ? node150 : node147;
							assign node147 = (inp[5]) ? 3'b110 : 3'b100;
							assign node150 = (inp[0]) ? 3'b101 : 3'b100;
				assign node153 = (inp[6]) ? node167 : node154;
					assign node154 = (inp[1]) ? node160 : node155;
						assign node155 = (inp[7]) ? node157 : 3'b000;
							assign node157 = (inp[0]) ? 3'b000 : 3'b000;
						assign node160 = (inp[2]) ? node164 : node161;
							assign node161 = (inp[0]) ? 3'b010 : 3'b000;
							assign node164 = (inp[8]) ? 3'b100 : 3'b000;
					assign node167 = (inp[10]) ? node175 : node168;
						assign node168 = (inp[2]) ? node172 : node169;
							assign node169 = (inp[1]) ? 3'b010 : 3'b000;
							assign node172 = (inp[0]) ? 3'b110 : 3'b100;
						assign node175 = (inp[7]) ? node179 : node176;
							assign node176 = (inp[2]) ? 3'b100 : 3'b000;
							assign node179 = (inp[0]) ? 3'b010 : 3'b100;
			assign node182 = (inp[9]) ? node210 : node183;
				assign node183 = (inp[6]) ? node195 : node184;
					assign node184 = (inp[0]) ? node190 : node185;
						assign node185 = (inp[5]) ? 3'b000 : node186;
							assign node186 = (inp[2]) ? 3'b000 : 3'b000;
						assign node190 = (inp[11]) ? 3'b000 : node191;
							assign node191 = (inp[10]) ? 3'b000 : 3'b100;
					assign node195 = (inp[11]) ? node203 : node196;
						assign node196 = (inp[0]) ? node200 : node197;
							assign node197 = (inp[5]) ? 3'b100 : 3'b010;
							assign node200 = (inp[1]) ? 3'b000 : 3'b110;
						assign node203 = (inp[5]) ? node207 : node204;
							assign node204 = (inp[0]) ? 3'b001 : 3'b000;
							assign node207 = (inp[8]) ? 3'b010 : 3'b000;
				assign node210 = (inp[0]) ? node212 : 3'b000;
					assign node212 = (inp[7]) ? node214 : 3'b000;
						assign node214 = (inp[2]) ? node218 : node215;
							assign node215 = (inp[5]) ? 3'b000 : 3'b000;
							assign node218 = (inp[6]) ? 3'b100 : 3'b000;

endmodule