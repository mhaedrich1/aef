module dtc_split75_bm57 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node7;
	wire [3-1:0] node8;
	wire [3-1:0] node9;
	wire [3-1:0] node10;
	wire [3-1:0] node11;
	wire [3-1:0] node14;
	wire [3-1:0] node17;
	wire [3-1:0] node19;
	wire [3-1:0] node22;
	wire [3-1:0] node23;
	wire [3-1:0] node25;
	wire [3-1:0] node29;
	wire [3-1:0] node30;
	wire [3-1:0] node31;
	wire [3-1:0] node33;
	wire [3-1:0] node36;
	wire [3-1:0] node38;
	wire [3-1:0] node41;
	wire [3-1:0] node43;
	wire [3-1:0] node44;
	wire [3-1:0] node48;
	wire [3-1:0] node49;
	wire [3-1:0] node50;
	wire [3-1:0] node51;
	wire [3-1:0] node55;
	wire [3-1:0] node56;
	wire [3-1:0] node58;
	wire [3-1:0] node61;
	wire [3-1:0] node62;
	wire [3-1:0] node66;
	wire [3-1:0] node67;
	wire [3-1:0] node68;
	wire [3-1:0] node69;
	wire [3-1:0] node73;
	wire [3-1:0] node74;
	wire [3-1:0] node77;
	wire [3-1:0] node80;
	wire [3-1:0] node81;
	wire [3-1:0] node84;
	wire [3-1:0] node87;
	wire [3-1:0] node88;
	wire [3-1:0] node89;
	wire [3-1:0] node91;
	wire [3-1:0] node92;
	wire [3-1:0] node93;
	wire [3-1:0] node96;
	wire [3-1:0] node99;
	wire [3-1:0] node101;
	wire [3-1:0] node104;
	wire [3-1:0] node105;
	wire [3-1:0] node106;
	wire [3-1:0] node109;
	wire [3-1:0] node112;
	wire [3-1:0] node113;
	wire [3-1:0] node114;
	wire [3-1:0] node117;
	wire [3-1:0] node120;
	wire [3-1:0] node121;
	wire [3-1:0] node124;
	wire [3-1:0] node127;
	wire [3-1:0] node128;
	wire [3-1:0] node129;
	wire [3-1:0] node131;
	wire [3-1:0] node134;
	wire [3-1:0] node135;
	wire [3-1:0] node136;
	wire [3-1:0] node139;
	wire [3-1:0] node142;
	wire [3-1:0] node144;
	wire [3-1:0] node147;
	wire [3-1:0] node148;
	wire [3-1:0] node150;
	wire [3-1:0] node153;
	wire [3-1:0] node155;
	wire [3-1:0] node158;
	wire [3-1:0] node159;
	wire [3-1:0] node160;
	wire [3-1:0] node161;
	wire [3-1:0] node163;
	wire [3-1:0] node164;
	wire [3-1:0] node165;
	wire [3-1:0] node168;
	wire [3-1:0] node171;
	wire [3-1:0] node172;
	wire [3-1:0] node175;
	wire [3-1:0] node178;
	wire [3-1:0] node180;
	wire [3-1:0] node182;
	wire [3-1:0] node185;
	wire [3-1:0] node186;
	wire [3-1:0] node187;
	wire [3-1:0] node189;
	wire [3-1:0] node192;
	wire [3-1:0] node193;
	wire [3-1:0] node194;
	wire [3-1:0] node197;
	wire [3-1:0] node201;
	wire [3-1:0] node202;
	wire [3-1:0] node203;
	wire [3-1:0] node206;
	wire [3-1:0] node209;
	wire [3-1:0] node210;
	wire [3-1:0] node211;
	wire [3-1:0] node214;
	wire [3-1:0] node217;
	wire [3-1:0] node218;
	wire [3-1:0] node221;
	wire [3-1:0] node224;
	wire [3-1:0] node225;
	wire [3-1:0] node226;
	wire [3-1:0] node227;
	wire [3-1:0] node229;
	wire [3-1:0] node230;
	wire [3-1:0] node234;
	wire [3-1:0] node235;
	wire [3-1:0] node236;
	wire [3-1:0] node239;
	wire [3-1:0] node242;
	wire [3-1:0] node243;
	wire [3-1:0] node246;
	wire [3-1:0] node249;
	wire [3-1:0] node250;
	wire [3-1:0] node251;
	wire [3-1:0] node254;
	wire [3-1:0] node257;
	wire [3-1:0] node258;
	wire [3-1:0] node259;
	wire [3-1:0] node262;
	wire [3-1:0] node265;
	wire [3-1:0] node266;
	wire [3-1:0] node270;
	wire [3-1:0] node271;
	wire [3-1:0] node272;
	wire [3-1:0] node273;
	wire [3-1:0] node274;
	wire [3-1:0] node279;
	wire [3-1:0] node281;
	wire [3-1:0] node284;
	wire [3-1:0] node285;
	wire [3-1:0] node286;
	wire [3-1:0] node287;
	wire [3-1:0] node290;
	wire [3-1:0] node293;
	wire [3-1:0] node295;
	wire [3-1:0] node298;
	wire [3-1:0] node300;
	wire [3-1:0] node301;
	wire [3-1:0] node305;
	wire [3-1:0] node306;
	wire [3-1:0] node307;
	wire [3-1:0] node308;
	wire [3-1:0] node309;
	wire [3-1:0] node310;
	wire [3-1:0] node313;
	wire [3-1:0] node315;
	wire [3-1:0] node318;
	wire [3-1:0] node319;
	wire [3-1:0] node320;
	wire [3-1:0] node325;
	wire [3-1:0] node326;
	wire [3-1:0] node327;
	wire [3-1:0] node329;
	wire [3-1:0] node330;
	wire [3-1:0] node333;
	wire [3-1:0] node336;
	wire [3-1:0] node337;
	wire [3-1:0] node338;
	wire [3-1:0] node341;
	wire [3-1:0] node344;
	wire [3-1:0] node346;
	wire [3-1:0] node349;
	wire [3-1:0] node350;
	wire [3-1:0] node351;
	wire [3-1:0] node355;
	wire [3-1:0] node356;
	wire [3-1:0] node357;
	wire [3-1:0] node362;
	wire [3-1:0] node363;
	wire [3-1:0] node364;
	wire [3-1:0] node365;
	wire [3-1:0] node366;
	wire [3-1:0] node370;
	wire [3-1:0] node371;
	wire [3-1:0] node373;
	wire [3-1:0] node377;
	wire [3-1:0] node378;
	wire [3-1:0] node380;
	wire [3-1:0] node381;
	wire [3-1:0] node384;
	wire [3-1:0] node387;
	wire [3-1:0] node388;
	wire [3-1:0] node392;
	wire [3-1:0] node393;
	wire [3-1:0] node394;
	wire [3-1:0] node396;
	wire [3-1:0] node399;
	wire [3-1:0] node400;
	wire [3-1:0] node404;
	wire [3-1:0] node405;
	wire [3-1:0] node407;
	wire [3-1:0] node410;
	wire [3-1:0] node411;
	wire [3-1:0] node415;
	wire [3-1:0] node416;
	wire [3-1:0] node417;
	wire [3-1:0] node418;
	wire [3-1:0] node419;
	wire [3-1:0] node420;
	wire [3-1:0] node423;
	wire [3-1:0] node426;
	wire [3-1:0] node427;
	wire [3-1:0] node430;
	wire [3-1:0] node433;
	wire [3-1:0] node435;
	wire [3-1:0] node436;
	wire [3-1:0] node437;
	wire [3-1:0] node440;
	wire [3-1:0] node444;
	wire [3-1:0] node445;
	wire [3-1:0] node446;
	wire [3-1:0] node447;
	wire [3-1:0] node449;
	wire [3-1:0] node452;
	wire [3-1:0] node453;
	wire [3-1:0] node456;
	wire [3-1:0] node459;
	wire [3-1:0] node460;
	wire [3-1:0] node463;
	wire [3-1:0] node466;
	wire [3-1:0] node467;
	wire [3-1:0] node468;
	wire [3-1:0] node471;
	wire [3-1:0] node474;
	wire [3-1:0] node475;
	wire [3-1:0] node476;
	wire [3-1:0] node481;
	wire [3-1:0] node482;
	wire [3-1:0] node483;
	wire [3-1:0] node484;
	wire [3-1:0] node485;
	wire [3-1:0] node488;
	wire [3-1:0] node491;
	wire [3-1:0] node493;
	wire [3-1:0] node494;
	wire [3-1:0] node498;
	wire [3-1:0] node499;
	wire [3-1:0] node500;
	wire [3-1:0] node503;
	wire [3-1:0] node506;
	wire [3-1:0] node507;
	wire [3-1:0] node509;
	wire [3-1:0] node512;
	wire [3-1:0] node513;
	wire [3-1:0] node516;
	wire [3-1:0] node519;
	wire [3-1:0] node520;
	wire [3-1:0] node521;
	wire [3-1:0] node524;
	wire [3-1:0] node527;
	wire [3-1:0] node528;
	wire [3-1:0] node530;
	wire [3-1:0] node532;
	wire [3-1:0] node535;
	wire [3-1:0] node536;
	wire [3-1:0] node537;
	wire [3-1:0] node540;
	wire [3-1:0] node543;
	wire [3-1:0] node545;
	wire [3-1:0] node548;
	wire [3-1:0] node549;
	wire [3-1:0] node550;
	wire [3-1:0] node551;
	wire [3-1:0] node552;
	wire [3-1:0] node553;
	wire [3-1:0] node554;
	wire [3-1:0] node557;
	wire [3-1:0] node558;
	wire [3-1:0] node560;
	wire [3-1:0] node563;
	wire [3-1:0] node566;
	wire [3-1:0] node567;
	wire [3-1:0] node568;
	wire [3-1:0] node569;
	wire [3-1:0] node572;
	wire [3-1:0] node575;
	wire [3-1:0] node576;
	wire [3-1:0] node579;
	wire [3-1:0] node582;
	wire [3-1:0] node583;
	wire [3-1:0] node584;
	wire [3-1:0] node588;
	wire [3-1:0] node589;
	wire [3-1:0] node592;
	wire [3-1:0] node595;
	wire [3-1:0] node596;
	wire [3-1:0] node597;
	wire [3-1:0] node598;
	wire [3-1:0] node601;
	wire [3-1:0] node604;
	wire [3-1:0] node605;
	wire [3-1:0] node606;
	wire [3-1:0] node610;
	wire [3-1:0] node611;
	wire [3-1:0] node614;
	wire [3-1:0] node617;
	wire [3-1:0] node618;
	wire [3-1:0] node619;
	wire [3-1:0] node622;
	wire [3-1:0] node624;
	wire [3-1:0] node627;
	wire [3-1:0] node628;
	wire [3-1:0] node629;
	wire [3-1:0] node633;
	wire [3-1:0] node635;
	wire [3-1:0] node638;
	wire [3-1:0] node639;
	wire [3-1:0] node640;
	wire [3-1:0] node641;
	wire [3-1:0] node643;
	wire [3-1:0] node644;
	wire [3-1:0] node647;
	wire [3-1:0] node650;
	wire [3-1:0] node651;
	wire [3-1:0] node654;
	wire [3-1:0] node655;
	wire [3-1:0] node659;
	wire [3-1:0] node660;
	wire [3-1:0] node661;
	wire [3-1:0] node662;
	wire [3-1:0] node666;
	wire [3-1:0] node668;
	wire [3-1:0] node671;
	wire [3-1:0] node673;
	wire [3-1:0] node675;
	wire [3-1:0] node678;
	wire [3-1:0] node679;
	wire [3-1:0] node680;
	wire [3-1:0] node682;
	wire [3-1:0] node685;
	wire [3-1:0] node686;
	wire [3-1:0] node688;
	wire [3-1:0] node691;
	wire [3-1:0] node692;
	wire [3-1:0] node695;
	wire [3-1:0] node698;
	wire [3-1:0] node699;
	wire [3-1:0] node701;
	wire [3-1:0] node702;
	wire [3-1:0] node706;
	wire [3-1:0] node709;
	wire [3-1:0] node710;
	wire [3-1:0] node711;
	wire [3-1:0] node712;
	wire [3-1:0] node713;
	wire [3-1:0] node716;
	wire [3-1:0] node717;
	wire [3-1:0] node719;
	wire [3-1:0] node722;
	wire [3-1:0] node723;
	wire [3-1:0] node727;
	wire [3-1:0] node728;
	wire [3-1:0] node731;
	wire [3-1:0] node732;
	wire [3-1:0] node734;
	wire [3-1:0] node737;
	wire [3-1:0] node738;
	wire [3-1:0] node742;
	wire [3-1:0] node743;
	wire [3-1:0] node744;
	wire [3-1:0] node747;
	wire [3-1:0] node748;
	wire [3-1:0] node751;
	wire [3-1:0] node754;
	wire [3-1:0] node755;
	wire [3-1:0] node757;
	wire [3-1:0] node758;
	wire [3-1:0] node761;
	wire [3-1:0] node764;
	wire [3-1:0] node765;
	wire [3-1:0] node766;
	wire [3-1:0] node769;
	wire [3-1:0] node772;
	wire [3-1:0] node773;
	wire [3-1:0] node777;
	wire [3-1:0] node778;
	wire [3-1:0] node779;
	wire [3-1:0] node780;
	wire [3-1:0] node781;
	wire [3-1:0] node782;
	wire [3-1:0] node787;
	wire [3-1:0] node789;
	wire [3-1:0] node790;
	wire [3-1:0] node794;
	wire [3-1:0] node795;
	wire [3-1:0] node796;
	wire [3-1:0] node799;
	wire [3-1:0] node802;
	wire [3-1:0] node803;
	wire [3-1:0] node804;
	wire [3-1:0] node807;
	wire [3-1:0] node811;
	wire [3-1:0] node812;
	wire [3-1:0] node813;
	wire [3-1:0] node814;
	wire [3-1:0] node815;
	wire [3-1:0] node818;
	wire [3-1:0] node821;
	wire [3-1:0] node823;
	wire [3-1:0] node826;
	wire [3-1:0] node827;
	wire [3-1:0] node828;
	wire [3-1:0] node832;
	wire [3-1:0] node834;
	wire [3-1:0] node837;
	wire [3-1:0] node838;
	wire [3-1:0] node840;
	wire [3-1:0] node842;
	wire [3-1:0] node845;
	wire [3-1:0] node846;
	wire [3-1:0] node848;
	wire [3-1:0] node851;
	wire [3-1:0] node852;
	wire [3-1:0] node855;
	wire [3-1:0] node858;
	wire [3-1:0] node859;
	wire [3-1:0] node860;
	wire [3-1:0] node861;
	wire [3-1:0] node862;
	wire [3-1:0] node863;
	wire [3-1:0] node864;
	wire [3-1:0] node867;
	wire [3-1:0] node870;
	wire [3-1:0] node871;
	wire [3-1:0] node874;
	wire [3-1:0] node877;
	wire [3-1:0] node878;
	wire [3-1:0] node880;
	wire [3-1:0] node884;
	wire [3-1:0] node885;
	wire [3-1:0] node886;
	wire [3-1:0] node887;
	wire [3-1:0] node891;
	wire [3-1:0] node892;
	wire [3-1:0] node896;
	wire [3-1:0] node897;
	wire [3-1:0] node899;
	wire [3-1:0] node903;
	wire [3-1:0] node904;
	wire [3-1:0] node905;
	wire [3-1:0] node906;
	wire [3-1:0] node907;
	wire [3-1:0] node908;
	wire [3-1:0] node911;
	wire [3-1:0] node914;
	wire [3-1:0] node915;
	wire [3-1:0] node918;
	wire [3-1:0] node921;
	wire [3-1:0] node922;
	wire [3-1:0] node925;
	wire [3-1:0] node928;
	wire [3-1:0] node929;
	wire [3-1:0] node931;
	wire [3-1:0] node934;
	wire [3-1:0] node936;
	wire [3-1:0] node939;
	wire [3-1:0] node940;
	wire [3-1:0] node941;
	wire [3-1:0] node942;
	wire [3-1:0] node945;
	wire [3-1:0] node948;
	wire [3-1:0] node949;
	wire [3-1:0] node952;
	wire [3-1:0] node955;
	wire [3-1:0] node956;
	wire [3-1:0] node959;
	wire [3-1:0] node960;
	wire [3-1:0] node964;
	wire [3-1:0] node965;
	wire [3-1:0] node966;
	wire [3-1:0] node967;
	wire [3-1:0] node968;
	wire [3-1:0] node970;
	wire [3-1:0] node973;
	wire [3-1:0] node974;
	wire [3-1:0] node978;
	wire [3-1:0] node981;
	wire [3-1:0] node982;
	wire [3-1:0] node983;
	wire [3-1:0] node985;
	wire [3-1:0] node988;
	wire [3-1:0] node989;
	wire [3-1:0] node993;
	wire [3-1:0] node996;
	wire [3-1:0] node997;
	wire [3-1:0] node998;
	wire [3-1:0] node999;
	wire [3-1:0] node1002;
	wire [3-1:0] node1003;
	wire [3-1:0] node1007;
	wire [3-1:0] node1010;
	wire [3-1:0] node1011;
	wire [3-1:0] node1012;
	wire [3-1:0] node1014;
	wire [3-1:0] node1017;
	wire [3-1:0] node1018;
	wire [3-1:0] node1022;
	wire [3-1:0] node1025;
	wire [3-1:0] node1026;
	wire [3-1:0] node1027;
	wire [3-1:0] node1028;
	wire [3-1:0] node1029;
	wire [3-1:0] node1030;
	wire [3-1:0] node1031;
	wire [3-1:0] node1033;
	wire [3-1:0] node1034;
	wire [3-1:0] node1035;
	wire [3-1:0] node1039;
	wire [3-1:0] node1040;
	wire [3-1:0] node1043;
	wire [3-1:0] node1046;
	wire [3-1:0] node1047;
	wire [3-1:0] node1050;
	wire [3-1:0] node1053;
	wire [3-1:0] node1054;
	wire [3-1:0] node1055;
	wire [3-1:0] node1057;
	wire [3-1:0] node1058;
	wire [3-1:0] node1061;
	wire [3-1:0] node1064;
	wire [3-1:0] node1065;
	wire [3-1:0] node1069;
	wire [3-1:0] node1070;
	wire [3-1:0] node1071;
	wire [3-1:0] node1072;
	wire [3-1:0] node1077;
	wire [3-1:0] node1079;
	wire [3-1:0] node1082;
	wire [3-1:0] node1083;
	wire [3-1:0] node1084;
	wire [3-1:0] node1085;
	wire [3-1:0] node1086;
	wire [3-1:0] node1089;
	wire [3-1:0] node1092;
	wire [3-1:0] node1094;
	wire [3-1:0] node1095;
	wire [3-1:0] node1098;
	wire [3-1:0] node1101;
	wire [3-1:0] node1102;
	wire [3-1:0] node1104;
	wire [3-1:0] node1105;
	wire [3-1:0] node1108;
	wire [3-1:0] node1111;
	wire [3-1:0] node1112;
	wire [3-1:0] node1113;
	wire [3-1:0] node1116;
	wire [3-1:0] node1119;
	wire [3-1:0] node1121;
	wire [3-1:0] node1124;
	wire [3-1:0] node1125;
	wire [3-1:0] node1126;
	wire [3-1:0] node1127;
	wire [3-1:0] node1128;
	wire [3-1:0] node1131;
	wire [3-1:0] node1134;
	wire [3-1:0] node1135;
	wire [3-1:0] node1138;
	wire [3-1:0] node1141;
	wire [3-1:0] node1142;
	wire [3-1:0] node1146;
	wire [3-1:0] node1147;
	wire [3-1:0] node1148;
	wire [3-1:0] node1151;
	wire [3-1:0] node1154;
	wire [3-1:0] node1155;
	wire [3-1:0] node1157;
	wire [3-1:0] node1161;
	wire [3-1:0] node1162;
	wire [3-1:0] node1163;
	wire [3-1:0] node1164;
	wire [3-1:0] node1165;
	wire [3-1:0] node1167;
	wire [3-1:0] node1169;
	wire [3-1:0] node1172;
	wire [3-1:0] node1175;
	wire [3-1:0] node1176;
	wire [3-1:0] node1178;
	wire [3-1:0] node1181;
	wire [3-1:0] node1183;
	wire [3-1:0] node1186;
	wire [3-1:0] node1187;
	wire [3-1:0] node1188;
	wire [3-1:0] node1189;
	wire [3-1:0] node1193;
	wire [3-1:0] node1195;
	wire [3-1:0] node1198;
	wire [3-1:0] node1199;
	wire [3-1:0] node1202;
	wire [3-1:0] node1203;
	wire [3-1:0] node1207;
	wire [3-1:0] node1208;
	wire [3-1:0] node1209;
	wire [3-1:0] node1210;
	wire [3-1:0] node1211;
	wire [3-1:0] node1214;
	wire [3-1:0] node1217;
	wire [3-1:0] node1218;
	wire [3-1:0] node1219;
	wire [3-1:0] node1222;
	wire [3-1:0] node1225;
	wire [3-1:0] node1226;
	wire [3-1:0] node1229;
	wire [3-1:0] node1232;
	wire [3-1:0] node1233;
	wire [3-1:0] node1235;
	wire [3-1:0] node1238;
	wire [3-1:0] node1239;
	wire [3-1:0] node1243;
	wire [3-1:0] node1244;
	wire [3-1:0] node1245;
	wire [3-1:0] node1246;
	wire [3-1:0] node1248;
	wire [3-1:0] node1252;
	wire [3-1:0] node1253;
	wire [3-1:0] node1256;
	wire [3-1:0] node1259;
	wire [3-1:0] node1260;
	wire [3-1:0] node1261;
	wire [3-1:0] node1262;
	wire [3-1:0] node1266;
	wire [3-1:0] node1268;
	wire [3-1:0] node1271;
	wire [3-1:0] node1272;
	wire [3-1:0] node1276;
	wire [3-1:0] node1277;
	wire [3-1:0] node1278;
	wire [3-1:0] node1279;
	wire [3-1:0] node1280;
	wire [3-1:0] node1282;
	wire [3-1:0] node1285;
	wire [3-1:0] node1287;
	wire [3-1:0] node1290;
	wire [3-1:0] node1291;
	wire [3-1:0] node1293;
	wire [3-1:0] node1296;
	wire [3-1:0] node1298;
	wire [3-1:0] node1301;
	wire [3-1:0] node1302;
	wire [3-1:0] node1303;
	wire [3-1:0] node1304;
	wire [3-1:0] node1306;
	wire [3-1:0] node1307;
	wire [3-1:0] node1310;
	wire [3-1:0] node1313;
	wire [3-1:0] node1314;
	wire [3-1:0] node1317;
	wire [3-1:0] node1320;
	wire [3-1:0] node1321;
	wire [3-1:0] node1323;
	wire [3-1:0] node1324;
	wire [3-1:0] node1327;
	wire [3-1:0] node1330;
	wire [3-1:0] node1332;
	wire [3-1:0] node1334;
	wire [3-1:0] node1337;
	wire [3-1:0] node1338;
	wire [3-1:0] node1341;
	wire [3-1:0] node1344;
	wire [3-1:0] node1345;
	wire [3-1:0] node1346;
	wire [3-1:0] node1347;
	wire [3-1:0] node1348;
	wire [3-1:0] node1349;
	wire [3-1:0] node1351;
	wire [3-1:0] node1355;
	wire [3-1:0] node1356;
	wire [3-1:0] node1359;
	wire [3-1:0] node1362;
	wire [3-1:0] node1363;
	wire [3-1:0] node1364;
	wire [3-1:0] node1367;
	wire [3-1:0] node1370;
	wire [3-1:0] node1371;
	wire [3-1:0] node1373;
	wire [3-1:0] node1376;
	wire [3-1:0] node1377;
	wire [3-1:0] node1380;
	wire [3-1:0] node1383;
	wire [3-1:0] node1384;
	wire [3-1:0] node1385;
	wire [3-1:0] node1386;
	wire [3-1:0] node1388;
	wire [3-1:0] node1391;
	wire [3-1:0] node1392;
	wire [3-1:0] node1395;
	wire [3-1:0] node1398;
	wire [3-1:0] node1399;
	wire [3-1:0] node1400;
	wire [3-1:0] node1404;
	wire [3-1:0] node1405;
	wire [3-1:0] node1408;
	wire [3-1:0] node1411;
	wire [3-1:0] node1412;
	wire [3-1:0] node1414;
	wire [3-1:0] node1416;
	wire [3-1:0] node1419;
	wire [3-1:0] node1420;
	wire [3-1:0] node1423;
	wire [3-1:0] node1426;
	wire [3-1:0] node1427;
	wire [3-1:0] node1430;
	wire [3-1:0] node1433;
	wire [3-1:0] node1434;
	wire [3-1:0] node1435;
	wire [3-1:0] node1436;
	wire [3-1:0] node1437;
	wire [3-1:0] node1438;
	wire [3-1:0] node1439;
	wire [3-1:0] node1440;
	wire [3-1:0] node1441;
	wire [3-1:0] node1444;
	wire [3-1:0] node1447;
	wire [3-1:0] node1448;
	wire [3-1:0] node1451;
	wire [3-1:0] node1454;
	wire [3-1:0] node1455;
	wire [3-1:0] node1456;
	wire [3-1:0] node1460;
	wire [3-1:0] node1462;
	wire [3-1:0] node1465;
	wire [3-1:0] node1466;
	wire [3-1:0] node1467;
	wire [3-1:0] node1469;
	wire [3-1:0] node1472;
	wire [3-1:0] node1474;
	wire [3-1:0] node1477;
	wire [3-1:0] node1478;
	wire [3-1:0] node1482;
	wire [3-1:0] node1483;
	wire [3-1:0] node1484;
	wire [3-1:0] node1485;
	wire [3-1:0] node1487;
	wire [3-1:0] node1490;
	wire [3-1:0] node1492;
	wire [3-1:0] node1495;
	wire [3-1:0] node1496;
	wire [3-1:0] node1500;
	wire [3-1:0] node1501;
	wire [3-1:0] node1502;
	wire [3-1:0] node1504;
	wire [3-1:0] node1507;
	wire [3-1:0] node1509;
	wire [3-1:0] node1512;
	wire [3-1:0] node1513;
	wire [3-1:0] node1517;
	wire [3-1:0] node1518;
	wire [3-1:0] node1519;
	wire [3-1:0] node1520;
	wire [3-1:0] node1521;
	wire [3-1:0] node1523;
	wire [3-1:0] node1526;
	wire [3-1:0] node1529;
	wire [3-1:0] node1532;
	wire [3-1:0] node1533;
	wire [3-1:0] node1534;
	wire [3-1:0] node1535;
	wire [3-1:0] node1540;
	wire [3-1:0] node1541;
	wire [3-1:0] node1543;
	wire [3-1:0] node1546;
	wire [3-1:0] node1548;
	wire [3-1:0] node1551;
	wire [3-1:0] node1552;
	wire [3-1:0] node1553;
	wire [3-1:0] node1554;
	wire [3-1:0] node1556;
	wire [3-1:0] node1560;
	wire [3-1:0] node1561;
	wire [3-1:0] node1564;
	wire [3-1:0] node1567;
	wire [3-1:0] node1568;
	wire [3-1:0] node1569;
	wire [3-1:0] node1570;
	wire [3-1:0] node1573;
	wire [3-1:0] node1577;
	wire [3-1:0] node1578;
	wire [3-1:0] node1579;
	wire [3-1:0] node1582;
	wire [3-1:0] node1585;
	wire [3-1:0] node1586;
	wire [3-1:0] node1589;
	wire [3-1:0] node1592;
	wire [3-1:0] node1593;
	wire [3-1:0] node1594;
	wire [3-1:0] node1595;
	wire [3-1:0] node1596;
	wire [3-1:0] node1601;
	wire [3-1:0] node1602;
	wire [3-1:0] node1603;
	wire [3-1:0] node1604;
	wire [3-1:0] node1605;
	wire [3-1:0] node1608;
	wire [3-1:0] node1611;
	wire [3-1:0] node1612;
	wire [3-1:0] node1615;
	wire [3-1:0] node1618;
	wire [3-1:0] node1619;
	wire [3-1:0] node1620;
	wire [3-1:0] node1624;
	wire [3-1:0] node1626;
	wire [3-1:0] node1630;
	wire [3-1:0] node1631;
	wire [3-1:0] node1632;
	wire [3-1:0] node1636;
	wire [3-1:0] node1637;
	wire [3-1:0] node1641;
	wire [3-1:0] node1642;
	wire [3-1:0] node1643;
	wire [3-1:0] node1644;
	wire [3-1:0] node1645;
	wire [3-1:0] node1646;
	wire [3-1:0] node1647;
	wire [3-1:0] node1648;
	wire [3-1:0] node1652;
	wire [3-1:0] node1653;
	wire [3-1:0] node1657;
	wire [3-1:0] node1660;
	wire [3-1:0] node1661;
	wire [3-1:0] node1662;
	wire [3-1:0] node1663;
	wire [3-1:0] node1666;
	wire [3-1:0] node1669;
	wire [3-1:0] node1671;
	wire [3-1:0] node1674;
	wire [3-1:0] node1675;
	wire [3-1:0] node1678;
	wire [3-1:0] node1681;
	wire [3-1:0] node1682;
	wire [3-1:0] node1683;
	wire [3-1:0] node1684;
	wire [3-1:0] node1685;
	wire [3-1:0] node1688;
	wire [3-1:0] node1691;
	wire [3-1:0] node1692;
	wire [3-1:0] node1695;
	wire [3-1:0] node1698;
	wire [3-1:0] node1699;
	wire [3-1:0] node1700;
	wire [3-1:0] node1703;
	wire [3-1:0] node1706;
	wire [3-1:0] node1708;
	wire [3-1:0] node1711;
	wire [3-1:0] node1712;
	wire [3-1:0] node1713;
	wire [3-1:0] node1714;
	wire [3-1:0] node1717;
	wire [3-1:0] node1721;
	wire [3-1:0] node1722;
	wire [3-1:0] node1723;
	wire [3-1:0] node1727;
	wire [3-1:0] node1728;
	wire [3-1:0] node1731;
	wire [3-1:0] node1734;
	wire [3-1:0] node1735;
	wire [3-1:0] node1736;
	wire [3-1:0] node1737;
	wire [3-1:0] node1738;
	wire [3-1:0] node1742;
	wire [3-1:0] node1743;
	wire [3-1:0] node1747;
	wire [3-1:0] node1748;
	wire [3-1:0] node1750;
	wire [3-1:0] node1751;
	wire [3-1:0] node1755;
	wire [3-1:0] node1756;
	wire [3-1:0] node1759;
	wire [3-1:0] node1762;
	wire [3-1:0] node1763;
	wire [3-1:0] node1764;
	wire [3-1:0] node1765;
	wire [3-1:0] node1769;
	wire [3-1:0] node1770;
	wire [3-1:0] node1774;
	wire [3-1:0] node1775;
	wire [3-1:0] node1776;
	wire [3-1:0] node1780;
	wire [3-1:0] node1781;
	wire [3-1:0] node1785;
	wire [3-1:0] node1786;
	wire [3-1:0] node1787;
	wire [3-1:0] node1788;
	wire [3-1:0] node1789;
	wire [3-1:0] node1793;
	wire [3-1:0] node1794;
	wire [3-1:0] node1799;
	wire [3-1:0] node1800;
	wire [3-1:0] node1801;
	wire [3-1:0] node1802;
	wire [3-1:0] node1806;
	wire [3-1:0] node1807;
	wire [3-1:0] node1812;
	wire [3-1:0] node1813;
	wire [3-1:0] node1814;
	wire [3-1:0] node1815;
	wire [3-1:0] node1816;
	wire [3-1:0] node1817;
	wire [3-1:0] node1818;
	wire [3-1:0] node1819;
	wire [3-1:0] node1820;
	wire [3-1:0] node1821;
	wire [3-1:0] node1825;
	wire [3-1:0] node1826;
	wire [3-1:0] node1830;
	wire [3-1:0] node1831;
	wire [3-1:0] node1835;
	wire [3-1:0] node1836;
	wire [3-1:0] node1837;
	wire [3-1:0] node1839;
	wire [3-1:0] node1842;
	wire [3-1:0] node1844;
	wire [3-1:0] node1847;
	wire [3-1:0] node1848;
	wire [3-1:0] node1850;
	wire [3-1:0] node1853;
	wire [3-1:0] node1855;
	wire [3-1:0] node1858;
	wire [3-1:0] node1859;
	wire [3-1:0] node1860;
	wire [3-1:0] node1861;
	wire [3-1:0] node1863;
	wire [3-1:0] node1865;
	wire [3-1:0] node1868;
	wire [3-1:0] node1869;
	wire [3-1:0] node1872;
	wire [3-1:0] node1875;
	wire [3-1:0] node1876;
	wire [3-1:0] node1878;
	wire [3-1:0] node1879;
	wire [3-1:0] node1883;
	wire [3-1:0] node1884;
	wire [3-1:0] node1886;
	wire [3-1:0] node1889;
	wire [3-1:0] node1891;
	wire [3-1:0] node1894;
	wire [3-1:0] node1895;
	wire [3-1:0] node1896;
	wire [3-1:0] node1897;
	wire [3-1:0] node1901;
	wire [3-1:0] node1902;
	wire [3-1:0] node1906;
	wire [3-1:0] node1907;
	wire [3-1:0] node1910;
	wire [3-1:0] node1911;
	wire [3-1:0] node1915;
	wire [3-1:0] node1916;
	wire [3-1:0] node1917;
	wire [3-1:0] node1918;
	wire [3-1:0] node1919;
	wire [3-1:0] node1920;
	wire [3-1:0] node1921;
	wire [3-1:0] node1924;
	wire [3-1:0] node1927;
	wire [3-1:0] node1928;
	wire [3-1:0] node1932;
	wire [3-1:0] node1933;
	wire [3-1:0] node1934;
	wire [3-1:0] node1937;
	wire [3-1:0] node1940;
	wire [3-1:0] node1941;
	wire [3-1:0] node1944;
	wire [3-1:0] node1947;
	wire [3-1:0] node1948;
	wire [3-1:0] node1949;
	wire [3-1:0] node1950;
	wire [3-1:0] node1953;
	wire [3-1:0] node1957;
	wire [3-1:0] node1959;
	wire [3-1:0] node1962;
	wire [3-1:0] node1963;
	wire [3-1:0] node1964;
	wire [3-1:0] node1965;
	wire [3-1:0] node1969;
	wire [3-1:0] node1971;
	wire [3-1:0] node1973;
	wire [3-1:0] node1976;
	wire [3-1:0] node1977;
	wire [3-1:0] node1979;
	wire [3-1:0] node1980;
	wire [3-1:0] node1983;
	wire [3-1:0] node1986;
	wire [3-1:0] node1987;
	wire [3-1:0] node1988;
	wire [3-1:0] node1991;
	wire [3-1:0] node1995;
	wire [3-1:0] node1996;
	wire [3-1:0] node1997;
	wire [3-1:0] node1998;
	wire [3-1:0] node1999;
	wire [3-1:0] node2001;
	wire [3-1:0] node2004;
	wire [3-1:0] node2007;
	wire [3-1:0] node2008;
	wire [3-1:0] node2009;
	wire [3-1:0] node2013;
	wire [3-1:0] node2016;
	wire [3-1:0] node2017;
	wire [3-1:0] node2020;
	wire [3-1:0] node2021;
	wire [3-1:0] node2023;
	wire [3-1:0] node2026;
	wire [3-1:0] node2029;
	wire [3-1:0] node2030;
	wire [3-1:0] node2031;
	wire [3-1:0] node2033;
	wire [3-1:0] node2034;
	wire [3-1:0] node2037;
	wire [3-1:0] node2040;
	wire [3-1:0] node2041;
	wire [3-1:0] node2045;
	wire [3-1:0] node2046;
	wire [3-1:0] node2048;
	wire [3-1:0] node2049;
	wire [3-1:0] node2052;
	wire [3-1:0] node2055;
	wire [3-1:0] node2056;
	wire [3-1:0] node2058;
	wire [3-1:0] node2061;
	wire [3-1:0] node2062;
	wire [3-1:0] node2065;
	wire [3-1:0] node2068;
	wire [3-1:0] node2069;
	wire [3-1:0] node2070;
	wire [3-1:0] node2071;
	wire [3-1:0] node2072;
	wire [3-1:0] node2073;
	wire [3-1:0] node2074;
	wire [3-1:0] node2075;
	wire [3-1:0] node2079;
	wire [3-1:0] node2081;
	wire [3-1:0] node2084;
	wire [3-1:0] node2086;
	wire [3-1:0] node2087;
	wire [3-1:0] node2090;
	wire [3-1:0] node2093;
	wire [3-1:0] node2094;
	wire [3-1:0] node2095;
	wire [3-1:0] node2096;
	wire [3-1:0] node2099;
	wire [3-1:0] node2102;
	wire [3-1:0] node2103;
	wire [3-1:0] node2107;
	wire [3-1:0] node2109;
	wire [3-1:0] node2110;
	wire [3-1:0] node2113;
	wire [3-1:0] node2116;
	wire [3-1:0] node2117;
	wire [3-1:0] node2118;
	wire [3-1:0] node2119;
	wire [3-1:0] node2120;
	wire [3-1:0] node2123;
	wire [3-1:0] node2126;
	wire [3-1:0] node2127;
	wire [3-1:0] node2131;
	wire [3-1:0] node2132;
	wire [3-1:0] node2133;
	wire [3-1:0] node2136;
	wire [3-1:0] node2139;
	wire [3-1:0] node2140;
	wire [3-1:0] node2143;
	wire [3-1:0] node2146;
	wire [3-1:0] node2147;
	wire [3-1:0] node2148;
	wire [3-1:0] node2149;
	wire [3-1:0] node2152;
	wire [3-1:0] node2155;
	wire [3-1:0] node2156;
	wire [3-1:0] node2160;
	wire [3-1:0] node2161;
	wire [3-1:0] node2163;
	wire [3-1:0] node2166;
	wire [3-1:0] node2168;
	wire [3-1:0] node2171;
	wire [3-1:0] node2172;
	wire [3-1:0] node2173;
	wire [3-1:0] node2175;
	wire [3-1:0] node2176;
	wire [3-1:0] node2177;
	wire [3-1:0] node2180;
	wire [3-1:0] node2183;
	wire [3-1:0] node2184;
	wire [3-1:0] node2187;
	wire [3-1:0] node2190;
	wire [3-1:0] node2191;
	wire [3-1:0] node2192;
	wire [3-1:0] node2194;
	wire [3-1:0] node2197;
	wire [3-1:0] node2198;
	wire [3-1:0] node2201;
	wire [3-1:0] node2204;
	wire [3-1:0] node2205;
	wire [3-1:0] node2208;
	wire [3-1:0] node2211;
	wire [3-1:0] node2212;
	wire [3-1:0] node2213;
	wire [3-1:0] node2214;
	wire [3-1:0] node2215;
	wire [3-1:0] node2218;
	wire [3-1:0] node2221;
	wire [3-1:0] node2222;
	wire [3-1:0] node2225;
	wire [3-1:0] node2228;
	wire [3-1:0] node2229;
	wire [3-1:0] node2232;
	wire [3-1:0] node2235;
	wire [3-1:0] node2236;
	wire [3-1:0] node2237;
	wire [3-1:0] node2238;
	wire [3-1:0] node2241;
	wire [3-1:0] node2244;
	wire [3-1:0] node2246;
	wire [3-1:0] node2249;
	wire [3-1:0] node2250;
	wire [3-1:0] node2251;
	wire [3-1:0] node2255;
	wire [3-1:0] node2258;
	wire [3-1:0] node2259;
	wire [3-1:0] node2260;
	wire [3-1:0] node2261;
	wire [3-1:0] node2262;
	wire [3-1:0] node2263;
	wire [3-1:0] node2266;
	wire [3-1:0] node2269;
	wire [3-1:0] node2271;
	wire [3-1:0] node2273;
	wire [3-1:0] node2276;
	wire [3-1:0] node2277;
	wire [3-1:0] node2279;
	wire [3-1:0] node2280;
	wire [3-1:0] node2283;
	wire [3-1:0] node2286;
	wire [3-1:0] node2288;
	wire [3-1:0] node2289;
	wire [3-1:0] node2292;
	wire [3-1:0] node2295;
	wire [3-1:0] node2296;
	wire [3-1:0] node2297;
	wire [3-1:0] node2298;
	wire [3-1:0] node2302;
	wire [3-1:0] node2303;
	wire [3-1:0] node2304;
	wire [3-1:0] node2307;
	wire [3-1:0] node2311;
	wire [3-1:0] node2312;
	wire [3-1:0] node2313;
	wire [3-1:0] node2317;
	wire [3-1:0] node2318;
	wire [3-1:0] node2320;
	wire [3-1:0] node2324;
	wire [3-1:0] node2325;
	wire [3-1:0] node2326;
	wire [3-1:0] node2327;
	wire [3-1:0] node2328;
	wire [3-1:0] node2332;
	wire [3-1:0] node2333;
	wire [3-1:0] node2337;
	wire [3-1:0] node2338;
	wire [3-1:0] node2340;
	wire [3-1:0] node2341;
	wire [3-1:0] node2345;
	wire [3-1:0] node2347;
	wire [3-1:0] node2350;
	wire [3-1:0] node2351;
	wire [3-1:0] node2352;
	wire [3-1:0] node2353;
	wire [3-1:0] node2354;
	wire [3-1:0] node2359;
	wire [3-1:0] node2360;
	wire [3-1:0] node2361;
	wire [3-1:0] node2366;
	wire [3-1:0] node2368;
	wire [3-1:0] node2369;
	wire [3-1:0] node2371;
	wire [3-1:0] node2375;
	wire [3-1:0] node2376;
	wire [3-1:0] node2377;
	wire [3-1:0] node2378;
	wire [3-1:0] node2379;
	wire [3-1:0] node2380;
	wire [3-1:0] node2382;
	wire [3-1:0] node2384;
	wire [3-1:0] node2387;
	wire [3-1:0] node2388;
	wire [3-1:0] node2390;
	wire [3-1:0] node2393;
	wire [3-1:0] node2396;
	wire [3-1:0] node2397;
	wire [3-1:0] node2398;
	wire [3-1:0] node2400;
	wire [3-1:0] node2403;
	wire [3-1:0] node2405;
	wire [3-1:0] node2408;
	wire [3-1:0] node2409;
	wire [3-1:0] node2411;
	wire [3-1:0] node2414;
	wire [3-1:0] node2416;
	wire [3-1:0] node2419;
	wire [3-1:0] node2420;
	wire [3-1:0] node2421;
	wire [3-1:0] node2424;
	wire [3-1:0] node2427;
	wire [3-1:0] node2428;
	wire [3-1:0] node2429;
	wire [3-1:0] node2432;
	wire [3-1:0] node2435;
	wire [3-1:0] node2436;
	wire [3-1:0] node2439;
	wire [3-1:0] node2442;
	wire [3-1:0] node2443;
	wire [3-1:0] node2444;
	wire [3-1:0] node2445;
	wire [3-1:0] node2446;
	wire [3-1:0] node2450;
	wire [3-1:0] node2453;
	wire [3-1:0] node2454;
	wire [3-1:0] node2456;
	wire [3-1:0] node2459;
	wire [3-1:0] node2460;
	wire [3-1:0] node2463;
	wire [3-1:0] node2466;
	wire [3-1:0] node2467;
	wire [3-1:0] node2468;
	wire [3-1:0] node2470;
	wire [3-1:0] node2473;
	wire [3-1:0] node2474;
	wire [3-1:0] node2478;
	wire [3-1:0] node2479;
	wire [3-1:0] node2482;
	wire [3-1:0] node2485;
	wire [3-1:0] node2486;
	wire [3-1:0] node2487;
	wire [3-1:0] node2488;
	wire [3-1:0] node2489;
	wire [3-1:0] node2491;
	wire [3-1:0] node2494;
	wire [3-1:0] node2495;
	wire [3-1:0] node2499;
	wire [3-1:0] node2500;
	wire [3-1:0] node2501;
	wire [3-1:0] node2505;
	wire [3-1:0] node2506;
	wire [3-1:0] node2510;
	wire [3-1:0] node2511;
	wire [3-1:0] node2512;
	wire [3-1:0] node2515;
	wire [3-1:0] node2518;
	wire [3-1:0] node2519;
	wire [3-1:0] node2520;
	wire [3-1:0] node2523;
	wire [3-1:0] node2526;
	wire [3-1:0] node2527;
	wire [3-1:0] node2530;
	wire [3-1:0] node2533;
	wire [3-1:0] node2534;
	wire [3-1:0] node2535;
	wire [3-1:0] node2536;
	wire [3-1:0] node2537;
	wire [3-1:0] node2541;
	wire [3-1:0] node2542;
	wire [3-1:0] node2547;
	wire [3-1:0] node2548;
	wire [3-1:0] node2549;
	wire [3-1:0] node2550;
	wire [3-1:0] node2554;
	wire [3-1:0] node2555;
	wire [3-1:0] node2560;
	wire [3-1:0] node2561;
	wire [3-1:0] node2562;
	wire [3-1:0] node2563;
	wire [3-1:0] node2564;
	wire [3-1:0] node2565;
	wire [3-1:0] node2566;
	wire [3-1:0] node2567;
	wire [3-1:0] node2570;
	wire [3-1:0] node2573;
	wire [3-1:0] node2574;
	wire [3-1:0] node2575;
	wire [3-1:0] node2576;
	wire [3-1:0] node2579;
	wire [3-1:0] node2583;
	wire [3-1:0] node2584;
	wire [3-1:0] node2585;
	wire [3-1:0] node2588;
	wire [3-1:0] node2591;
	wire [3-1:0] node2592;
	wire [3-1:0] node2595;
	wire [3-1:0] node2598;
	wire [3-1:0] node2599;
	wire [3-1:0] node2600;
	wire [3-1:0] node2602;
	wire [3-1:0] node2605;
	wire [3-1:0] node2606;
	wire [3-1:0] node2607;
	wire [3-1:0] node2610;
	wire [3-1:0] node2613;
	wire [3-1:0] node2614;
	wire [3-1:0] node2617;
	wire [3-1:0] node2620;
	wire [3-1:0] node2621;
	wire [3-1:0] node2623;
	wire [3-1:0] node2625;
	wire [3-1:0] node2628;
	wire [3-1:0] node2629;
	wire [3-1:0] node2632;
	wire [3-1:0] node2635;
	wire [3-1:0] node2636;
	wire [3-1:0] node2637;
	wire [3-1:0] node2639;
	wire [3-1:0] node2642;
	wire [3-1:0] node2643;
	wire [3-1:0] node2644;
	wire [3-1:0] node2648;
	wire [3-1:0] node2649;
	wire [3-1:0] node2652;
	wire [3-1:0] node2655;
	wire [3-1:0] node2656;
	wire [3-1:0] node2657;
	wire [3-1:0] node2660;
	wire [3-1:0] node2663;
	wire [3-1:0] node2664;
	wire [3-1:0] node2665;
	wire [3-1:0] node2668;
	wire [3-1:0] node2672;
	wire [3-1:0] node2673;
	wire [3-1:0] node2674;
	wire [3-1:0] node2675;
	wire [3-1:0] node2676;
	wire [3-1:0] node2677;
	wire [3-1:0] node2680;
	wire [3-1:0] node2684;
	wire [3-1:0] node2685;
	wire [3-1:0] node2686;
	wire [3-1:0] node2687;
	wire [3-1:0] node2690;
	wire [3-1:0] node2693;
	wire [3-1:0] node2695;
	wire [3-1:0] node2699;
	wire [3-1:0] node2700;
	wire [3-1:0] node2701;
	wire [3-1:0] node2705;
	wire [3-1:0] node2706;
	wire [3-1:0] node2710;
	wire [3-1:0] node2711;
	wire [3-1:0] node2712;
	wire [3-1:0] node2713;
	wire [3-1:0] node2714;
	wire [3-1:0] node2717;
	wire [3-1:0] node2721;
	wire [3-1:0] node2722;
	wire [3-1:0] node2726;
	wire [3-1:0] node2727;
	wire [3-1:0] node2728;
	wire [3-1:0] node2729;
	wire [3-1:0] node2732;
	wire [3-1:0] node2736;
	wire [3-1:0] node2737;
	wire [3-1:0] node2741;
	wire [3-1:0] node2742;
	wire [3-1:0] node2743;
	wire [3-1:0] node2744;
	wire [3-1:0] node2745;
	wire [3-1:0] node2746;
	wire [3-1:0] node2748;
	wire [3-1:0] node2751;
	wire [3-1:0] node2752;
	wire [3-1:0] node2756;
	wire [3-1:0] node2757;
	wire [3-1:0] node2758;
	wire [3-1:0] node2759;
	wire [3-1:0] node2762;
	wire [3-1:0] node2766;
	wire [3-1:0] node2767;
	wire [3-1:0] node2770;
	wire [3-1:0] node2773;
	wire [3-1:0] node2774;
	wire [3-1:0] node2775;
	wire [3-1:0] node2776;
	wire [3-1:0] node2777;
	wire [3-1:0] node2782;
	wire [3-1:0] node2783;
	wire [3-1:0] node2785;
	wire [3-1:0] node2788;
	wire [3-1:0] node2789;
	wire [3-1:0] node2792;
	wire [3-1:0] node2795;
	wire [3-1:0] node2796;
	wire [3-1:0] node2797;
	wire [3-1:0] node2801;
	wire [3-1:0] node2802;
	wire [3-1:0] node2805;
	wire [3-1:0] node2808;
	wire [3-1:0] node2809;
	wire [3-1:0] node2810;
	wire [3-1:0] node2813;
	wire [3-1:0] node2816;
	wire [3-1:0] node2817;
	wire [3-1:0] node2820;
	wire [3-1:0] node2823;
	wire [3-1:0] node2824;
	wire [3-1:0] node2825;
	wire [3-1:0] node2829;
	wire [3-1:0] node2830;
	wire [3-1:0] node2834;
	wire [3-1:0] node2835;
	wire [3-1:0] node2836;
	wire [3-1:0] node2837;
	wire [3-1:0] node2838;
	wire [3-1:0] node2839;
	wire [3-1:0] node2841;
	wire [3-1:0] node2844;
	wire [3-1:0] node2846;
	wire [3-1:0] node2849;
	wire [3-1:0] node2850;
	wire [3-1:0] node2851;
	wire [3-1:0] node2855;
	wire [3-1:0] node2856;
	wire [3-1:0] node2860;
	wire [3-1:0] node2861;
	wire [3-1:0] node2862;
	wire [3-1:0] node2863;
	wire [3-1:0] node2864;
	wire [3-1:0] node2865;
	wire [3-1:0] node2868;
	wire [3-1:0] node2871;
	wire [3-1:0] node2873;
	wire [3-1:0] node2876;
	wire [3-1:0] node2877;
	wire [3-1:0] node2880;
	wire [3-1:0] node2883;
	wire [3-1:0] node2884;
	wire [3-1:0] node2886;
	wire [3-1:0] node2887;
	wire [3-1:0] node2891;
	wire [3-1:0] node2892;
	wire [3-1:0] node2893;
	wire [3-1:0] node2896;
	wire [3-1:0] node2899;
	wire [3-1:0] node2901;
	wire [3-1:0] node2904;
	wire [3-1:0] node2905;
	wire [3-1:0] node2908;
	wire [3-1:0] node2911;
	wire [3-1:0] node2912;
	wire [3-1:0] node2913;
	wire [3-1:0] node2914;
	wire [3-1:0] node2915;
	wire [3-1:0] node2919;
	wire [3-1:0] node2920;
	wire [3-1:0] node2925;
	wire [3-1:0] node2926;
	wire [3-1:0] node2927;
	wire [3-1:0] node2928;
	wire [3-1:0] node2932;
	wire [3-1:0] node2933;
	wire [3-1:0] node2938;
	wire [3-1:0] node2939;
	wire [3-1:0] node2940;
	wire [3-1:0] node2941;
	wire [3-1:0] node2945;
	wire [3-1:0] node2946;
	wire [3-1:0] node2950;
	wire [3-1:0] node2951;

	assign outp = (inp[4]) ? node1812 : node1;
		assign node1 = (inp[6]) ? node1025 : node2;
			assign node2 = (inp[8]) ? node548 : node3;
				assign node3 = (inp[5]) ? node305 : node4;
					assign node4 = (inp[3]) ? node158 : node5;
						assign node5 = (inp[10]) ? node87 : node6;
							assign node6 = (inp[7]) ? node48 : node7;
								assign node7 = (inp[11]) ? node29 : node8;
									assign node8 = (inp[1]) ? node22 : node9;
										assign node9 = (inp[2]) ? node17 : node10;
											assign node10 = (inp[9]) ? node14 : node11;
												assign node11 = (inp[0]) ? 3'b001 : 3'b000;
												assign node14 = (inp[0]) ? 3'b000 : 3'b001;
											assign node17 = (inp[9]) ? node19 : 3'b000;
												assign node19 = (inp[0]) ? 3'b000 : 3'b001;
										assign node22 = (inp[0]) ? 3'b000 : node23;
											assign node23 = (inp[2]) ? node25 : 3'b000;
												assign node25 = (inp[9]) ? 3'b000 : 3'b001;
									assign node29 = (inp[0]) ? node41 : node30;
										assign node30 = (inp[9]) ? node36 : node31;
											assign node31 = (inp[2]) ? node33 : 3'b000;
												assign node33 = (inp[1]) ? 3'b001 : 3'b000;
											assign node36 = (inp[2]) ? node38 : 3'b001;
												assign node38 = (inp[1]) ? 3'b000 : 3'b001;
										assign node41 = (inp[2]) ? node43 : 3'b001;
											assign node43 = (inp[9]) ? 3'b001 : node44;
												assign node44 = (inp[1]) ? 3'b000 : 3'b001;
								assign node48 = (inp[11]) ? node66 : node49;
									assign node49 = (inp[2]) ? node55 : node50;
										assign node50 = (inp[9]) ? 3'b001 : node51;
											assign node51 = (inp[0]) ? 3'b001 : 3'b000;
										assign node55 = (inp[0]) ? node61 : node56;
											assign node56 = (inp[1]) ? node58 : 3'b000;
												assign node58 = (inp[9]) ? 3'b000 : 3'b001;
											assign node61 = (inp[9]) ? 3'b001 : node62;
												assign node62 = (inp[1]) ? 3'b000 : 3'b001;
									assign node66 = (inp[1]) ? node80 : node67;
										assign node67 = (inp[9]) ? node73 : node68;
											assign node68 = (inp[0]) ? 3'b011 : node69;
												assign node69 = (inp[2]) ? 3'b011 : 3'b010;
											assign node73 = (inp[0]) ? node77 : node74;
												assign node74 = (inp[2]) ? 3'b010 : 3'b011;
												assign node77 = (inp[2]) ? 3'b011 : 3'b010;
										assign node80 = (inp[9]) ? node84 : node81;
											assign node81 = (inp[0]) ? 3'b010 : 3'b011;
											assign node84 = (inp[0]) ? 3'b011 : 3'b010;
							assign node87 = (inp[7]) ? node127 : node88;
								assign node88 = (inp[11]) ? node104 : node89;
									assign node89 = (inp[1]) ? node91 : 3'b011;
										assign node91 = (inp[0]) ? node99 : node92;
											assign node92 = (inp[9]) ? node96 : node93;
												assign node93 = (inp[2]) ? 3'b011 : 3'b010;
												assign node96 = (inp[2]) ? 3'b010 : 3'b011;
											assign node99 = (inp[9]) ? node101 : 3'b011;
												assign node101 = (inp[2]) ? 3'b011 : 3'b010;
									assign node104 = (inp[2]) ? node112 : node105;
										assign node105 = (inp[9]) ? node109 : node106;
											assign node106 = (inp[0]) ? 3'b010 : 3'b011;
											assign node109 = (inp[0]) ? 3'b011 : 3'b010;
										assign node112 = (inp[1]) ? node120 : node113;
											assign node113 = (inp[0]) ? node117 : node114;
												assign node114 = (inp[9]) ? 3'b010 : 3'b011;
												assign node117 = (inp[9]) ? 3'b011 : 3'b010;
											assign node120 = (inp[9]) ? node124 : node121;
												assign node121 = (inp[0]) ? 3'b011 : 3'b010;
												assign node124 = (inp[0]) ? 3'b010 : 3'b011;
								assign node127 = (inp[11]) ? node147 : node128;
									assign node128 = (inp[1]) ? node134 : node129;
										assign node129 = (inp[9]) ? node131 : 3'b011;
											assign node131 = (inp[0]) ? 3'b010 : 3'b011;
										assign node134 = (inp[9]) ? node142 : node135;
											assign node135 = (inp[0]) ? node139 : node136;
												assign node136 = (inp[2]) ? 3'b011 : 3'b010;
												assign node139 = (inp[2]) ? 3'b010 : 3'b011;
											assign node142 = (inp[0]) ? node144 : 3'b010;
												assign node144 = (inp[2]) ? 3'b011 : 3'b010;
									assign node147 = (inp[9]) ? node153 : node148;
										assign node148 = (inp[0]) ? node150 : 3'b000;
											assign node150 = (inp[1]) ? 3'b000 : 3'b001;
										assign node153 = (inp[0]) ? node155 : 3'b001;
											assign node155 = (inp[1]) ? 3'b001 : 3'b000;
						assign node158 = (inp[10]) ? node224 : node159;
							assign node159 = (inp[7]) ? node185 : node160;
								assign node160 = (inp[9]) ? node178 : node161;
									assign node161 = (inp[1]) ? node163 : 3'b010;
										assign node163 = (inp[11]) ? node171 : node164;
											assign node164 = (inp[2]) ? node168 : node165;
												assign node165 = (inp[0]) ? 3'b011 : 3'b010;
												assign node168 = (inp[0]) ? 3'b010 : 3'b011;
											assign node171 = (inp[2]) ? node175 : node172;
												assign node172 = (inp[0]) ? 3'b011 : 3'b010;
												assign node175 = (inp[0]) ? 3'b010 : 3'b011;
									assign node178 = (inp[0]) ? node180 : 3'b011;
										assign node180 = (inp[2]) ? node182 : 3'b010;
											assign node182 = (inp[1]) ? 3'b011 : 3'b010;
								assign node185 = (inp[11]) ? node201 : node186;
									assign node186 = (inp[2]) ? node192 : node187;
										assign node187 = (inp[9]) ? node189 : 3'b010;
											assign node189 = (inp[1]) ? 3'b010 : 3'b011;
										assign node192 = (inp[9]) ? 3'b011 : node193;
											assign node193 = (inp[0]) ? node197 : node194;
												assign node194 = (inp[1]) ? 3'b010 : 3'b011;
												assign node197 = (inp[1]) ? 3'b011 : 3'b010;
									assign node201 = (inp[1]) ? node209 : node202;
										assign node202 = (inp[0]) ? node206 : node203;
											assign node203 = (inp[9]) ? 3'b001 : 3'b000;
											assign node206 = (inp[9]) ? 3'b000 : 3'b001;
										assign node209 = (inp[2]) ? node217 : node210;
											assign node210 = (inp[9]) ? node214 : node211;
												assign node211 = (inp[0]) ? 3'b001 : 3'b000;
												assign node214 = (inp[0]) ? 3'b000 : 3'b001;
											assign node217 = (inp[9]) ? node221 : node218;
												assign node218 = (inp[0]) ? 3'b000 : 3'b001;
												assign node221 = (inp[0]) ? 3'b001 : 3'b000;
							assign node224 = (inp[11]) ? node270 : node225;
								assign node225 = (inp[2]) ? node249 : node226;
									assign node226 = (inp[1]) ? node234 : node227;
										assign node227 = (inp[7]) ? node229 : 3'b000;
											assign node229 = (inp[9]) ? 3'b000 : node230;
												assign node230 = (inp[0]) ? 3'b000 : 3'b001;
										assign node234 = (inp[7]) ? node242 : node235;
											assign node235 = (inp[0]) ? node239 : node236;
												assign node236 = (inp[9]) ? 3'b000 : 3'b001;
												assign node239 = (inp[9]) ? 3'b001 : 3'b000;
											assign node242 = (inp[9]) ? node246 : node243;
												assign node243 = (inp[0]) ? 3'b001 : 3'b000;
												assign node246 = (inp[0]) ? 3'b000 : 3'b001;
									assign node249 = (inp[9]) ? node257 : node250;
										assign node250 = (inp[7]) ? node254 : node251;
											assign node251 = (inp[0]) ? 3'b000 : 3'b001;
											assign node254 = (inp[0]) ? 3'b001 : 3'b000;
										assign node257 = (inp[1]) ? node265 : node258;
											assign node258 = (inp[0]) ? node262 : node259;
												assign node259 = (inp[7]) ? 3'b001 : 3'b000;
												assign node262 = (inp[7]) ? 3'b000 : 3'b001;
											assign node265 = (inp[0]) ? 3'b001 : node266;
												assign node266 = (inp[7]) ? 3'b001 : 3'b000;
								assign node270 = (inp[7]) ? node284 : node271;
									assign node271 = (inp[2]) ? node279 : node272;
										assign node272 = (inp[0]) ? 3'b000 : node273;
											assign node273 = (inp[9]) ? 3'b000 : node274;
												assign node274 = (inp[1]) ? 3'b000 : 3'b001;
										assign node279 = (inp[0]) ? node281 : 3'b001;
											assign node281 = (inp[9]) ? 3'b000 : 3'b001;
									assign node284 = (inp[1]) ? node298 : node285;
										assign node285 = (inp[2]) ? node293 : node286;
											assign node286 = (inp[9]) ? node290 : node287;
												assign node287 = (inp[0]) ? 3'b010 : 3'b011;
												assign node290 = (inp[0]) ? 3'b011 : 3'b010;
											assign node293 = (inp[0]) ? node295 : 3'b010;
												assign node295 = (inp[9]) ? 3'b011 : 3'b010;
										assign node298 = (inp[9]) ? node300 : 3'b010;
											assign node300 = (inp[0]) ? 3'b010 : node301;
												assign node301 = (inp[2]) ? 3'b011 : 3'b010;
					assign node305 = (inp[3]) ? node415 : node306;
						assign node306 = (inp[10]) ? node362 : node307;
							assign node307 = (inp[11]) ? node325 : node308;
								assign node308 = (inp[0]) ? node318 : node309;
									assign node309 = (inp[9]) ? node313 : node310;
										assign node310 = (inp[1]) ? 3'b100 : 3'b101;
										assign node313 = (inp[2]) ? node315 : 3'b101;
											assign node315 = (inp[1]) ? 3'b101 : 3'b100;
									assign node318 = (inp[9]) ? 3'b100 : node319;
										assign node319 = (inp[1]) ? 3'b101 : node320;
											assign node320 = (inp[2]) ? 3'b100 : 3'b101;
								assign node325 = (inp[7]) ? node349 : node326;
									assign node326 = (inp[2]) ? node336 : node327;
										assign node327 = (inp[1]) ? node329 : 3'b110;
											assign node329 = (inp[0]) ? node333 : node330;
												assign node330 = (inp[9]) ? 3'b111 : 3'b110;
												assign node333 = (inp[9]) ? 3'b110 : 3'b111;
										assign node336 = (inp[1]) ? node344 : node337;
											assign node337 = (inp[9]) ? node341 : node338;
												assign node338 = (inp[0]) ? 3'b110 : 3'b111;
												assign node341 = (inp[0]) ? 3'b111 : 3'b110;
											assign node344 = (inp[0]) ? node346 : 3'b111;
												assign node346 = (inp[9]) ? 3'b110 : 3'b111;
									assign node349 = (inp[9]) ? node355 : node350;
										assign node350 = (inp[0]) ? 3'b100 : node351;
											assign node351 = (inp[1]) ? 3'b101 : 3'b100;
										assign node355 = (inp[0]) ? 3'b101 : node356;
											assign node356 = (inp[1]) ? 3'b100 : node357;
												assign node357 = (inp[2]) ? 3'b101 : 3'b100;
							assign node362 = (inp[7]) ? node392 : node363;
								assign node363 = (inp[11]) ? node377 : node364;
									assign node364 = (inp[2]) ? node370 : node365;
										assign node365 = (inp[0]) ? 3'b111 : node366;
											assign node366 = (inp[9]) ? 3'b111 : 3'b110;
										assign node370 = (inp[0]) ? 3'b110 : node371;
											assign node371 = (inp[1]) ? node373 : 3'b110;
												assign node373 = (inp[9]) ? 3'b111 : 3'b110;
									assign node377 = (inp[2]) ? node387 : node378;
										assign node378 = (inp[0]) ? node380 : 3'b101;
											assign node380 = (inp[1]) ? node384 : node381;
												assign node381 = (inp[9]) ? 3'b101 : 3'b100;
												assign node384 = (inp[9]) ? 3'b100 : 3'b101;
										assign node387 = (inp[9]) ? 3'b100 : node388;
											assign node388 = (inp[1]) ? 3'b100 : 3'b101;
								assign node392 = (inp[0]) ? node404 : node393;
									assign node393 = (inp[9]) ? node399 : node394;
										assign node394 = (inp[2]) ? node396 : 3'b110;
											assign node396 = (inp[1]) ? 3'b110 : 3'b111;
										assign node399 = (inp[1]) ? 3'b111 : node400;
											assign node400 = (inp[2]) ? 3'b110 : 3'b111;
									assign node404 = (inp[9]) ? node410 : node405;
										assign node405 = (inp[2]) ? node407 : 3'b111;
											assign node407 = (inp[1]) ? 3'b111 : 3'b110;
										assign node410 = (inp[1]) ? 3'b110 : node411;
											assign node411 = (inp[2]) ? 3'b111 : 3'b110;
						assign node415 = (inp[10]) ? node481 : node416;
							assign node416 = (inp[11]) ? node444 : node417;
								assign node417 = (inp[1]) ? node433 : node418;
									assign node418 = (inp[7]) ? node426 : node419;
										assign node419 = (inp[9]) ? node423 : node420;
											assign node420 = (inp[0]) ? 3'b111 : 3'b110;
											assign node423 = (inp[0]) ? 3'b110 : 3'b111;
										assign node426 = (inp[9]) ? node430 : node427;
											assign node427 = (inp[0]) ? 3'b110 : 3'b111;
											assign node430 = (inp[0]) ? 3'b111 : 3'b110;
									assign node433 = (inp[0]) ? node435 : 3'b111;
										assign node435 = (inp[9]) ? 3'b111 : node436;
											assign node436 = (inp[2]) ? node440 : node437;
												assign node437 = (inp[7]) ? 3'b111 : 3'b110;
												assign node440 = (inp[7]) ? 3'b110 : 3'b111;
								assign node444 = (inp[7]) ? node466 : node445;
									assign node445 = (inp[1]) ? node459 : node446;
										assign node446 = (inp[0]) ? node452 : node447;
											assign node447 = (inp[2]) ? node449 : 3'b100;
												assign node449 = (inp[9]) ? 3'b101 : 3'b100;
											assign node452 = (inp[9]) ? node456 : node453;
												assign node453 = (inp[2]) ? 3'b101 : 3'b100;
												assign node456 = (inp[2]) ? 3'b100 : 3'b101;
										assign node459 = (inp[9]) ? node463 : node460;
											assign node460 = (inp[0]) ? 3'b100 : 3'b101;
											assign node463 = (inp[0]) ? 3'b101 : 3'b100;
									assign node466 = (inp[1]) ? node474 : node467;
										assign node467 = (inp[0]) ? node471 : node468;
											assign node468 = (inp[9]) ? 3'b111 : 3'b110;
											assign node471 = (inp[9]) ? 3'b110 : 3'b111;
										assign node474 = (inp[9]) ? 3'b110 : node475;
											assign node475 = (inp[0]) ? 3'b111 : node476;
												assign node476 = (inp[2]) ? 3'b110 : 3'b111;
							assign node481 = (inp[7]) ? node519 : node482;
								assign node482 = (inp[11]) ? node498 : node483;
									assign node483 = (inp[2]) ? node491 : node484;
										assign node484 = (inp[9]) ? node488 : node485;
											assign node485 = (inp[0]) ? 3'b100 : 3'b101;
											assign node488 = (inp[0]) ? 3'b101 : 3'b100;
										assign node491 = (inp[9]) ? node493 : 3'b101;
											assign node493 = (inp[0]) ? 3'b101 : node494;
												assign node494 = (inp[1]) ? 3'b100 : 3'b101;
									assign node498 = (inp[2]) ? node506 : node499;
										assign node499 = (inp[9]) ? node503 : node500;
											assign node500 = (inp[0]) ? 3'b111 : 3'b110;
											assign node503 = (inp[0]) ? 3'b110 : 3'b111;
										assign node506 = (inp[0]) ? node512 : node507;
											assign node507 = (inp[1]) ? node509 : 3'b110;
												assign node509 = (inp[9]) ? 3'b111 : 3'b110;
											assign node512 = (inp[9]) ? node516 : node513;
												assign node513 = (inp[1]) ? 3'b111 : 3'b110;
												assign node516 = (inp[1]) ? 3'b110 : 3'b111;
								assign node519 = (inp[2]) ? node527 : node520;
									assign node520 = (inp[9]) ? node524 : node521;
										assign node521 = (inp[0]) ? 3'b101 : 3'b100;
										assign node524 = (inp[0]) ? 3'b100 : 3'b101;
									assign node527 = (inp[11]) ? node535 : node528;
										assign node528 = (inp[1]) ? node530 : 3'b101;
											assign node530 = (inp[0]) ? node532 : 3'b101;
												assign node532 = (inp[9]) ? 3'b100 : 3'b101;
										assign node535 = (inp[1]) ? node543 : node536;
											assign node536 = (inp[9]) ? node540 : node537;
												assign node537 = (inp[0]) ? 3'b100 : 3'b101;
												assign node540 = (inp[0]) ? 3'b101 : 3'b100;
											assign node543 = (inp[0]) ? node545 : 3'b101;
												assign node545 = (inp[9]) ? 3'b100 : 3'b101;
				assign node548 = (inp[2]) ? node858 : node549;
					assign node549 = (inp[0]) ? node709 : node550;
						assign node550 = (inp[10]) ? node638 : node551;
							assign node551 = (inp[9]) ? node595 : node552;
								assign node552 = (inp[1]) ? node566 : node553;
									assign node553 = (inp[3]) ? node557 : node554;
										assign node554 = (inp[7]) ? 3'b110 : 3'b100;
										assign node557 = (inp[7]) ? node563 : node558;
											assign node558 = (inp[5]) ? node560 : 3'b110;
												assign node560 = (inp[11]) ? 3'b111 : 3'b110;
											assign node563 = (inp[11]) ? 3'b100 : 3'b101;
									assign node566 = (inp[11]) ? node582 : node567;
										assign node567 = (inp[5]) ? node575 : node568;
											assign node568 = (inp[3]) ? node572 : node569;
												assign node569 = (inp[7]) ? 3'b111 : 3'b101;
												assign node572 = (inp[7]) ? 3'b100 : 3'b111;
											assign node575 = (inp[7]) ? node579 : node576;
												assign node576 = (inp[3]) ? 3'b111 : 3'b101;
												assign node579 = (inp[3]) ? 3'b101 : 3'b111;
										assign node582 = (inp[5]) ? node588 : node583;
											assign node583 = (inp[3]) ? 3'b101 : node584;
												assign node584 = (inp[7]) ? 3'b111 : 3'b101;
											assign node588 = (inp[7]) ? node592 : node589;
												assign node589 = (inp[3]) ? 3'b110 : 3'b101;
												assign node592 = (inp[3]) ? 3'b100 : 3'b110;
								assign node595 = (inp[1]) ? node617 : node596;
									assign node596 = (inp[5]) ? node604 : node597;
										assign node597 = (inp[3]) ? node601 : node598;
											assign node598 = (inp[7]) ? 3'b111 : 3'b101;
											assign node601 = (inp[7]) ? 3'b101 : 3'b111;
										assign node604 = (inp[11]) ? node610 : node605;
											assign node605 = (inp[7]) ? 3'b111 : node606;
												assign node606 = (inp[3]) ? 3'b111 : 3'b101;
											assign node610 = (inp[7]) ? node614 : node611;
												assign node611 = (inp[3]) ? 3'b110 : 3'b101;
												assign node614 = (inp[3]) ? 3'b100 : 3'b110;
									assign node617 = (inp[11]) ? node627 : node618;
										assign node618 = (inp[7]) ? node622 : node619;
											assign node619 = (inp[3]) ? 3'b110 : 3'b100;
											assign node622 = (inp[3]) ? node624 : 3'b110;
												assign node624 = (inp[5]) ? 3'b100 : 3'b101;
										assign node627 = (inp[5]) ? node633 : node628;
											assign node628 = (inp[7]) ? 3'b110 : node629;
												assign node629 = (inp[3]) ? 3'b110 : 3'b100;
											assign node633 = (inp[3]) ? node635 : 3'b111;
												assign node635 = (inp[7]) ? 3'b101 : 3'b111;
							assign node638 = (inp[1]) ? node678 : node639;
								assign node639 = (inp[9]) ? node659 : node640;
									assign node640 = (inp[5]) ? node650 : node641;
										assign node641 = (inp[11]) ? node643 : 3'b100;
											assign node643 = (inp[3]) ? node647 : node644;
												assign node644 = (inp[7]) ? 3'b110 : 3'b101;
												assign node647 = (inp[7]) ? 3'b101 : 3'b111;
										assign node650 = (inp[3]) ? node654 : node651;
											assign node651 = (inp[7]) ? 3'b110 : 3'b100;
											assign node654 = (inp[7]) ? 3'b100 : node655;
												assign node655 = (inp[11]) ? 3'b110 : 3'b111;
									assign node659 = (inp[7]) ? node671 : node660;
										assign node660 = (inp[3]) ? node666 : node661;
											assign node661 = (inp[5]) ? 3'b101 : node662;
												assign node662 = (inp[11]) ? 3'b100 : 3'b101;
											assign node666 = (inp[11]) ? node668 : 3'b110;
												assign node668 = (inp[5]) ? 3'b111 : 3'b110;
										assign node671 = (inp[3]) ? node673 : 3'b111;
											assign node673 = (inp[11]) ? node675 : 3'b101;
												assign node675 = (inp[5]) ? 3'b101 : 3'b100;
								assign node678 = (inp[9]) ? node698 : node679;
									assign node679 = (inp[11]) ? node685 : node680;
										assign node680 = (inp[3]) ? node682 : 3'b111;
											assign node682 = (inp[7]) ? 3'b101 : 3'b111;
										assign node685 = (inp[5]) ? node691 : node686;
											assign node686 = (inp[3]) ? node688 : 3'b100;
												assign node688 = (inp[7]) ? 3'b100 : 3'b110;
											assign node691 = (inp[3]) ? node695 : node692;
												assign node692 = (inp[7]) ? 3'b111 : 3'b101;
												assign node695 = (inp[7]) ? 3'b101 : 3'b111;
									assign node698 = (inp[7]) ? node706 : node699;
										assign node699 = (inp[3]) ? node701 : 3'b100;
											assign node701 = (inp[11]) ? 3'b110 : node702;
												assign node702 = (inp[5]) ? 3'b111 : 3'b110;
										assign node706 = (inp[3]) ? 3'b100 : 3'b110;
						assign node709 = (inp[11]) ? node777 : node710;
							assign node710 = (inp[9]) ? node742 : node711;
								assign node711 = (inp[1]) ? node727 : node712;
									assign node712 = (inp[3]) ? node716 : node713;
										assign node713 = (inp[7]) ? 3'b110 : 3'b100;
										assign node716 = (inp[7]) ? node722 : node717;
											assign node717 = (inp[5]) ? node719 : 3'b110;
												assign node719 = (inp[10]) ? 3'b111 : 3'b110;
											assign node722 = (inp[5]) ? 3'b100 : node723;
												assign node723 = (inp[10]) ? 3'b100 : 3'b101;
									assign node727 = (inp[3]) ? node731 : node728;
										assign node728 = (inp[7]) ? 3'b111 : 3'b101;
										assign node731 = (inp[7]) ? node737 : node732;
											assign node732 = (inp[10]) ? node734 : 3'b111;
												assign node734 = (inp[5]) ? 3'b110 : 3'b111;
											assign node737 = (inp[10]) ? 3'b101 : node738;
												assign node738 = (inp[5]) ? 3'b101 : 3'b100;
								assign node742 = (inp[1]) ? node754 : node743;
									assign node743 = (inp[3]) ? node747 : node744;
										assign node744 = (inp[7]) ? 3'b111 : 3'b101;
										assign node747 = (inp[7]) ? node751 : node748;
											assign node748 = (inp[10]) ? 3'b110 : 3'b111;
											assign node751 = (inp[5]) ? 3'b101 : 3'b100;
									assign node754 = (inp[10]) ? node764 : node755;
										assign node755 = (inp[5]) ? node757 : 3'b110;
											assign node757 = (inp[3]) ? node761 : node758;
												assign node758 = (inp[7]) ? 3'b110 : 3'b100;
												assign node761 = (inp[7]) ? 3'b100 : 3'b110;
										assign node764 = (inp[5]) ? node772 : node765;
											assign node765 = (inp[3]) ? node769 : node766;
												assign node766 = (inp[7]) ? 3'b110 : 3'b100;
												assign node769 = (inp[7]) ? 3'b100 : 3'b110;
											assign node772 = (inp[7]) ? 3'b100 : node773;
												assign node773 = (inp[3]) ? 3'b111 : 3'b100;
							assign node777 = (inp[5]) ? node811 : node778;
								assign node778 = (inp[7]) ? node794 : node779;
									assign node779 = (inp[3]) ? node787 : node780;
										assign node780 = (inp[10]) ? 3'b101 : node781;
											assign node781 = (inp[9]) ? 3'b101 : node782;
												assign node782 = (inp[1]) ? 3'b101 : 3'b100;
										assign node787 = (inp[1]) ? node789 : 3'b111;
											assign node789 = (inp[10]) ? 3'b111 : node790;
												assign node790 = (inp[9]) ? 3'b110 : 3'b111;
									assign node794 = (inp[3]) ? node802 : node795;
										assign node795 = (inp[9]) ? node799 : node796;
											assign node796 = (inp[1]) ? 3'b111 : 3'b110;
											assign node799 = (inp[1]) ? 3'b110 : 3'b111;
										assign node802 = (inp[1]) ? 3'b101 : node803;
											assign node803 = (inp[9]) ? node807 : node804;
												assign node804 = (inp[10]) ? 3'b101 : 3'b100;
												assign node807 = (inp[10]) ? 3'b100 : 3'b101;
								assign node811 = (inp[9]) ? node837 : node812;
									assign node812 = (inp[1]) ? node826 : node813;
										assign node813 = (inp[10]) ? node821 : node814;
											assign node814 = (inp[3]) ? node818 : node815;
												assign node815 = (inp[7]) ? 3'b111 : 3'b100;
												assign node818 = (inp[7]) ? 3'b101 : 3'b111;
											assign node821 = (inp[3]) ? node823 : 3'b110;
												assign node823 = (inp[7]) ? 3'b100 : 3'b110;
										assign node826 = (inp[10]) ? node832 : node827;
											assign node827 = (inp[7]) ? 3'b110 : node828;
												assign node828 = (inp[3]) ? 3'b110 : 3'b101;
											assign node832 = (inp[3]) ? node834 : 3'b101;
												assign node834 = (inp[7]) ? 3'b101 : 3'b111;
									assign node837 = (inp[1]) ? node845 : node838;
										assign node838 = (inp[3]) ? node840 : 3'b101;
											assign node840 = (inp[10]) ? node842 : 3'b110;
												assign node842 = (inp[7]) ? 3'b101 : 3'b111;
										assign node845 = (inp[10]) ? node851 : node846;
											assign node846 = (inp[7]) ? node848 : 3'b100;
												assign node848 = (inp[3]) ? 3'b101 : 3'b111;
											assign node851 = (inp[3]) ? node855 : node852;
												assign node852 = (inp[7]) ? 3'b110 : 3'b100;
												assign node855 = (inp[7]) ? 3'b100 : 3'b110;
					assign node858 = (inp[11]) ? node964 : node859;
						assign node859 = (inp[9]) ? node903 : node860;
							assign node860 = (inp[1]) ? node884 : node861;
								assign node861 = (inp[3]) ? node877 : node862;
									assign node862 = (inp[7]) ? node870 : node863;
										assign node863 = (inp[5]) ? node867 : node864;
											assign node864 = (inp[10]) ? 3'b101 : 3'b100;
											assign node867 = (inp[10]) ? 3'b100 : 3'b101;
										assign node870 = (inp[5]) ? node874 : node871;
											assign node871 = (inp[10]) ? 3'b111 : 3'b110;
											assign node874 = (inp[10]) ? 3'b110 : 3'b111;
									assign node877 = (inp[7]) ? 3'b100 : node878;
										assign node878 = (inp[10]) ? node880 : 3'b110;
											assign node880 = (inp[5]) ? 3'b110 : 3'b111;
								assign node884 = (inp[3]) ? node896 : node885;
									assign node885 = (inp[7]) ? node891 : node886;
										assign node886 = (inp[5]) ? 3'b100 : node887;
											assign node887 = (inp[10]) ? 3'b100 : 3'b101;
										assign node891 = (inp[5]) ? 3'b110 : node892;
											assign node892 = (inp[10]) ? 3'b110 : 3'b111;
									assign node896 = (inp[7]) ? 3'b101 : node897;
										assign node897 = (inp[10]) ? node899 : 3'b111;
											assign node899 = (inp[5]) ? 3'b111 : 3'b110;
							assign node903 = (inp[1]) ? node939 : node904;
								assign node904 = (inp[3]) ? node928 : node905;
									assign node905 = (inp[7]) ? node921 : node906;
										assign node906 = (inp[0]) ? node914 : node907;
											assign node907 = (inp[10]) ? node911 : node908;
												assign node908 = (inp[5]) ? 3'b100 : 3'b101;
												assign node911 = (inp[5]) ? 3'b101 : 3'b100;
											assign node914 = (inp[5]) ? node918 : node915;
												assign node915 = (inp[10]) ? 3'b100 : 3'b101;
												assign node918 = (inp[10]) ? 3'b101 : 3'b100;
										assign node921 = (inp[10]) ? node925 : node922;
											assign node922 = (inp[5]) ? 3'b110 : 3'b111;
											assign node925 = (inp[5]) ? 3'b111 : 3'b110;
									assign node928 = (inp[7]) ? node934 : node929;
										assign node929 = (inp[10]) ? node931 : 3'b111;
											assign node931 = (inp[5]) ? 3'b111 : 3'b110;
										assign node934 = (inp[5]) ? node936 : 3'b101;
											assign node936 = (inp[10]) ? 3'b101 : 3'b100;
								assign node939 = (inp[3]) ? node955 : node940;
									assign node940 = (inp[7]) ? node948 : node941;
										assign node941 = (inp[5]) ? node945 : node942;
											assign node942 = (inp[10]) ? 3'b101 : 3'b100;
											assign node945 = (inp[10]) ? 3'b100 : 3'b101;
										assign node948 = (inp[10]) ? node952 : node949;
											assign node949 = (inp[5]) ? 3'b111 : 3'b110;
											assign node952 = (inp[5]) ? 3'b110 : 3'b111;
									assign node955 = (inp[7]) ? node959 : node956;
										assign node956 = (inp[10]) ? 3'b111 : 3'b110;
										assign node959 = (inp[10]) ? 3'b100 : node960;
											assign node960 = (inp[5]) ? 3'b101 : 3'b100;
						assign node964 = (inp[9]) ? node996 : node965;
							assign node965 = (inp[1]) ? node981 : node966;
								assign node966 = (inp[3]) ? node978 : node967;
									assign node967 = (inp[7]) ? node973 : node968;
										assign node968 = (inp[10]) ? node970 : 3'b100;
											assign node970 = (inp[5]) ? 3'b101 : 3'b100;
										assign node973 = (inp[10]) ? 3'b110 : node974;
											assign node974 = (inp[5]) ? 3'b110 : 3'b111;
									assign node978 = (inp[7]) ? 3'b100 : 3'b110;
								assign node981 = (inp[3]) ? node993 : node982;
									assign node982 = (inp[7]) ? node988 : node983;
										assign node983 = (inp[10]) ? node985 : 3'b101;
											assign node985 = (inp[5]) ? 3'b100 : 3'b101;
										assign node988 = (inp[5]) ? 3'b111 : node989;
											assign node989 = (inp[10]) ? 3'b111 : 3'b110;
									assign node993 = (inp[7]) ? 3'b101 : 3'b111;
							assign node996 = (inp[1]) ? node1010 : node997;
								assign node997 = (inp[3]) ? node1007 : node998;
									assign node998 = (inp[7]) ? node1002 : node999;
										assign node999 = (inp[10]) ? 3'b100 : 3'b101;
										assign node1002 = (inp[5]) ? 3'b111 : node1003;
											assign node1003 = (inp[10]) ? 3'b111 : 3'b110;
									assign node1007 = (inp[7]) ? 3'b101 : 3'b111;
								assign node1010 = (inp[3]) ? node1022 : node1011;
									assign node1011 = (inp[7]) ? node1017 : node1012;
										assign node1012 = (inp[5]) ? node1014 : 3'b100;
											assign node1014 = (inp[0]) ? 3'b101 : 3'b100;
										assign node1017 = (inp[5]) ? 3'b110 : node1018;
											assign node1018 = (inp[10]) ? 3'b110 : 3'b111;
									assign node1022 = (inp[7]) ? 3'b100 : 3'b110;
			assign node1025 = (inp[5]) ? node1433 : node1026;
				assign node1026 = (inp[8]) ? node1276 : node1027;
					assign node1027 = (inp[3]) ? node1161 : node1028;
						assign node1028 = (inp[10]) ? node1082 : node1029;
							assign node1029 = (inp[7]) ? node1053 : node1030;
								assign node1030 = (inp[2]) ? node1046 : node1031;
									assign node1031 = (inp[1]) ? node1033 : 3'b101;
										assign node1033 = (inp[11]) ? node1039 : node1034;
											assign node1034 = (inp[9]) ? 3'b101 : node1035;
												assign node1035 = (inp[0]) ? 3'b100 : 3'b101;
											assign node1039 = (inp[9]) ? node1043 : node1040;
												assign node1040 = (inp[0]) ? 3'b100 : 3'b101;
												assign node1043 = (inp[0]) ? 3'b101 : 3'b100;
									assign node1046 = (inp[9]) ? node1050 : node1047;
										assign node1047 = (inp[0]) ? 3'b101 : 3'b100;
										assign node1050 = (inp[0]) ? 3'b100 : 3'b101;
								assign node1053 = (inp[11]) ? node1069 : node1054;
									assign node1054 = (inp[0]) ? node1064 : node1055;
										assign node1055 = (inp[1]) ? node1057 : 3'b110;
											assign node1057 = (inp[2]) ? node1061 : node1058;
												assign node1058 = (inp[9]) ? 3'b110 : 3'b111;
												assign node1061 = (inp[9]) ? 3'b111 : 3'b110;
										assign node1064 = (inp[2]) ? 3'b111 : node1065;
											assign node1065 = (inp[9]) ? 3'b111 : 3'b110;
									assign node1069 = (inp[1]) ? node1077 : node1070;
										assign node1070 = (inp[2]) ? 3'b100 : node1071;
											assign node1071 = (inp[0]) ? 3'b101 : node1072;
												assign node1072 = (inp[9]) ? 3'b100 : 3'b101;
										assign node1077 = (inp[9]) ? node1079 : 3'b101;
											assign node1079 = (inp[2]) ? 3'b101 : 3'b100;
							assign node1082 = (inp[7]) ? node1124 : node1083;
								assign node1083 = (inp[0]) ? node1101 : node1084;
									assign node1084 = (inp[2]) ? node1092 : node1085;
										assign node1085 = (inp[9]) ? node1089 : node1086;
											assign node1086 = (inp[11]) ? 3'b111 : 3'b110;
											assign node1089 = (inp[11]) ? 3'b110 : 3'b111;
										assign node1092 = (inp[9]) ? node1094 : 3'b111;
											assign node1094 = (inp[11]) ? node1098 : node1095;
												assign node1095 = (inp[1]) ? 3'b111 : 3'b110;
												assign node1098 = (inp[1]) ? 3'b110 : 3'b111;
									assign node1101 = (inp[1]) ? node1111 : node1102;
										assign node1102 = (inp[2]) ? node1104 : 3'b111;
											assign node1104 = (inp[9]) ? node1108 : node1105;
												assign node1105 = (inp[11]) ? 3'b111 : 3'b110;
												assign node1108 = (inp[11]) ? 3'b110 : 3'b111;
										assign node1111 = (inp[2]) ? node1119 : node1112;
											assign node1112 = (inp[9]) ? node1116 : node1113;
												assign node1113 = (inp[11]) ? 3'b110 : 3'b111;
												assign node1116 = (inp[11]) ? 3'b111 : 3'b110;
											assign node1119 = (inp[11]) ? node1121 : 3'b111;
												assign node1121 = (inp[9]) ? 3'b111 : 3'b110;
								assign node1124 = (inp[11]) ? node1146 : node1125;
									assign node1125 = (inp[2]) ? node1141 : node1126;
										assign node1126 = (inp[9]) ? node1134 : node1127;
											assign node1127 = (inp[1]) ? node1131 : node1128;
												assign node1128 = (inp[0]) ? 3'b100 : 3'b101;
												assign node1131 = (inp[0]) ? 3'b101 : 3'b100;
											assign node1134 = (inp[0]) ? node1138 : node1135;
												assign node1135 = (inp[1]) ? 3'b101 : 3'b100;
												assign node1138 = (inp[1]) ? 3'b100 : 3'b101;
										assign node1141 = (inp[9]) ? 3'b101 : node1142;
											assign node1142 = (inp[0]) ? 3'b100 : 3'b101;
									assign node1146 = (inp[2]) ? node1154 : node1147;
										assign node1147 = (inp[9]) ? node1151 : node1148;
											assign node1148 = (inp[1]) ? 3'b110 : 3'b111;
											assign node1151 = (inp[0]) ? 3'b110 : 3'b111;
										assign node1154 = (inp[9]) ? 3'b111 : node1155;
											assign node1155 = (inp[1]) ? node1157 : 3'b111;
												assign node1157 = (inp[0]) ? 3'b111 : 3'b110;
						assign node1161 = (inp[10]) ? node1207 : node1162;
							assign node1162 = (inp[11]) ? node1186 : node1163;
								assign node1163 = (inp[7]) ? node1175 : node1164;
									assign node1164 = (inp[9]) ? node1172 : node1165;
										assign node1165 = (inp[0]) ? node1167 : 3'b110;
											assign node1167 = (inp[1]) ? node1169 : 3'b111;
												assign node1169 = (inp[2]) ? 3'b111 : 3'b110;
										assign node1172 = (inp[0]) ? 3'b110 : 3'b111;
									assign node1175 = (inp[9]) ? node1181 : node1176;
										assign node1176 = (inp[1]) ? node1178 : 3'b101;
											assign node1178 = (inp[0]) ? 3'b100 : 3'b101;
										assign node1181 = (inp[0]) ? node1183 : 3'b100;
											assign node1183 = (inp[2]) ? 3'b100 : 3'b101;
								assign node1186 = (inp[0]) ? node1198 : node1187;
									assign node1187 = (inp[9]) ? node1193 : node1188;
										assign node1188 = (inp[2]) ? 3'b110 : node1189;
											assign node1189 = (inp[1]) ? 3'b111 : 3'b110;
										assign node1193 = (inp[1]) ? node1195 : 3'b111;
											assign node1195 = (inp[2]) ? 3'b111 : 3'b110;
									assign node1198 = (inp[9]) ? node1202 : node1199;
										assign node1199 = (inp[2]) ? 3'b111 : 3'b110;
										assign node1202 = (inp[2]) ? 3'b110 : node1203;
											assign node1203 = (inp[1]) ? 3'b111 : 3'b110;
							assign node1207 = (inp[7]) ? node1243 : node1208;
								assign node1208 = (inp[9]) ? node1232 : node1209;
									assign node1209 = (inp[1]) ? node1217 : node1210;
										assign node1210 = (inp[0]) ? node1214 : node1211;
											assign node1211 = (inp[11]) ? 3'b100 : 3'b101;
											assign node1214 = (inp[11]) ? 3'b101 : 3'b100;
										assign node1217 = (inp[2]) ? node1225 : node1218;
											assign node1218 = (inp[0]) ? node1222 : node1219;
												assign node1219 = (inp[11]) ? 3'b101 : 3'b100;
												assign node1222 = (inp[11]) ? 3'b100 : 3'b101;
											assign node1225 = (inp[0]) ? node1229 : node1226;
												assign node1226 = (inp[11]) ? 3'b100 : 3'b101;
												assign node1229 = (inp[11]) ? 3'b101 : 3'b100;
									assign node1232 = (inp[11]) ? node1238 : node1233;
										assign node1233 = (inp[0]) ? node1235 : 3'b100;
											assign node1235 = (inp[2]) ? 3'b101 : 3'b100;
										assign node1238 = (inp[0]) ? 3'b100 : node1239;
											assign node1239 = (inp[1]) ? 3'b100 : 3'b101;
								assign node1243 = (inp[11]) ? node1259 : node1244;
									assign node1244 = (inp[2]) ? node1252 : node1245;
										assign node1245 = (inp[1]) ? 3'b110 : node1246;
											assign node1246 = (inp[0]) ? node1248 : 3'b110;
												assign node1248 = (inp[9]) ? 3'b110 : 3'b111;
										assign node1252 = (inp[0]) ? node1256 : node1253;
											assign node1253 = (inp[9]) ? 3'b111 : 3'b110;
											assign node1256 = (inp[9]) ? 3'b110 : 3'b111;
									assign node1259 = (inp[0]) ? node1271 : node1260;
										assign node1260 = (inp[9]) ? node1266 : node1261;
											assign node1261 = (inp[2]) ? 3'b100 : node1262;
												assign node1262 = (inp[1]) ? 3'b101 : 3'b100;
											assign node1266 = (inp[1]) ? node1268 : 3'b101;
												assign node1268 = (inp[2]) ? 3'b101 : 3'b100;
										assign node1271 = (inp[9]) ? 3'b100 : node1272;
											assign node1272 = (inp[1]) ? 3'b100 : 3'b101;
					assign node1276 = (inp[11]) ? node1344 : node1277;
						assign node1277 = (inp[3]) ? node1301 : node1278;
							assign node1278 = (inp[10]) ? node1290 : node1279;
								assign node1279 = (inp[9]) ? node1285 : node1280;
									assign node1280 = (inp[7]) ? node1282 : 3'b000;
										assign node1282 = (inp[2]) ? 3'b001 : 3'b000;
									assign node1285 = (inp[7]) ? node1287 : 3'b001;
										assign node1287 = (inp[2]) ? 3'b000 : 3'b001;
								assign node1290 = (inp[9]) ? node1296 : node1291;
									assign node1291 = (inp[7]) ? node1293 : 3'b001;
										assign node1293 = (inp[2]) ? 3'b000 : 3'b001;
									assign node1296 = (inp[2]) ? node1298 : 3'b000;
										assign node1298 = (inp[7]) ? 3'b001 : 3'b000;
							assign node1301 = (inp[2]) ? node1337 : node1302;
								assign node1302 = (inp[0]) ? node1320 : node1303;
									assign node1303 = (inp[10]) ? node1313 : node1304;
										assign node1304 = (inp[1]) ? node1306 : 3'b011;
											assign node1306 = (inp[9]) ? node1310 : node1307;
												assign node1307 = (inp[7]) ? 3'b011 : 3'b010;
												assign node1310 = (inp[7]) ? 3'b010 : 3'b011;
										assign node1313 = (inp[9]) ? node1317 : node1314;
											assign node1314 = (inp[7]) ? 3'b010 : 3'b011;
											assign node1317 = (inp[7]) ? 3'b011 : 3'b010;
									assign node1320 = (inp[1]) ? node1330 : node1321;
										assign node1321 = (inp[9]) ? node1323 : 3'b011;
											assign node1323 = (inp[7]) ? node1327 : node1324;
												assign node1324 = (inp[10]) ? 3'b010 : 3'b011;
												assign node1327 = (inp[10]) ? 3'b011 : 3'b010;
										assign node1330 = (inp[7]) ? node1332 : 3'b011;
											assign node1332 = (inp[10]) ? node1334 : 3'b011;
												assign node1334 = (inp[9]) ? 3'b011 : 3'b010;
								assign node1337 = (inp[10]) ? node1341 : node1338;
									assign node1338 = (inp[9]) ? 3'b011 : 3'b010;
									assign node1341 = (inp[9]) ? 3'b010 : 3'b011;
						assign node1344 = (inp[3]) ? node1426 : node1345;
							assign node1345 = (inp[10]) ? node1383 : node1346;
								assign node1346 = (inp[2]) ? node1362 : node1347;
									assign node1347 = (inp[0]) ? node1355 : node1348;
										assign node1348 = (inp[1]) ? 3'b010 : node1349;
											assign node1349 = (inp[7]) ? node1351 : 3'b010;
												assign node1351 = (inp[9]) ? 3'b010 : 3'b011;
										assign node1355 = (inp[9]) ? node1359 : node1356;
											assign node1356 = (inp[7]) ? 3'b011 : 3'b010;
											assign node1359 = (inp[1]) ? 3'b011 : 3'b010;
									assign node1362 = (inp[0]) ? node1370 : node1363;
										assign node1363 = (inp[9]) ? node1367 : node1364;
											assign node1364 = (inp[7]) ? 3'b011 : 3'b010;
											assign node1367 = (inp[7]) ? 3'b010 : 3'b011;
										assign node1370 = (inp[1]) ? node1376 : node1371;
											assign node1371 = (inp[9]) ? node1373 : 3'b010;
												assign node1373 = (inp[7]) ? 3'b010 : 3'b011;
											assign node1376 = (inp[9]) ? node1380 : node1377;
												assign node1377 = (inp[7]) ? 3'b011 : 3'b010;
												assign node1380 = (inp[7]) ? 3'b010 : 3'b011;
								assign node1383 = (inp[2]) ? node1411 : node1384;
									assign node1384 = (inp[0]) ? node1398 : node1385;
										assign node1385 = (inp[1]) ? node1391 : node1386;
											assign node1386 = (inp[7]) ? node1388 : 3'b010;
												assign node1388 = (inp[9]) ? 3'b010 : 3'b011;
											assign node1391 = (inp[7]) ? node1395 : node1392;
												assign node1392 = (inp[9]) ? 3'b011 : 3'b010;
												assign node1395 = (inp[9]) ? 3'b010 : 3'b011;
										assign node1398 = (inp[1]) ? node1404 : node1399;
											assign node1399 = (inp[7]) ? 3'b011 : node1400;
												assign node1400 = (inp[9]) ? 3'b011 : 3'b010;
											assign node1404 = (inp[9]) ? node1408 : node1405;
												assign node1405 = (inp[7]) ? 3'b011 : 3'b010;
												assign node1408 = (inp[7]) ? 3'b010 : 3'b011;
									assign node1411 = (inp[0]) ? node1419 : node1412;
										assign node1412 = (inp[1]) ? node1414 : 3'b011;
											assign node1414 = (inp[7]) ? node1416 : 3'b011;
												assign node1416 = (inp[9]) ? 3'b010 : 3'b011;
										assign node1419 = (inp[7]) ? node1423 : node1420;
											assign node1420 = (inp[9]) ? 3'b011 : 3'b010;
											assign node1423 = (inp[9]) ? 3'b010 : 3'b011;
							assign node1426 = (inp[9]) ? node1430 : node1427;
								assign node1427 = (inp[2]) ? 3'b001 : 3'b000;
								assign node1430 = (inp[2]) ? 3'b000 : 3'b001;
				assign node1433 = (inp[3]) ? node1641 : node1434;
					assign node1434 = (inp[8]) ? node1592 : node1435;
						assign node1435 = (inp[10]) ? node1517 : node1436;
							assign node1436 = (inp[7]) ? node1482 : node1437;
								assign node1437 = (inp[11]) ? node1465 : node1438;
									assign node1438 = (inp[2]) ? node1454 : node1439;
										assign node1439 = (inp[1]) ? node1447 : node1440;
											assign node1440 = (inp[9]) ? node1444 : node1441;
												assign node1441 = (inp[0]) ? 3'b011 : 3'b010;
												assign node1444 = (inp[0]) ? 3'b010 : 3'b011;
											assign node1447 = (inp[0]) ? node1451 : node1448;
												assign node1448 = (inp[9]) ? 3'b010 : 3'b011;
												assign node1451 = (inp[9]) ? 3'b011 : 3'b010;
										assign node1454 = (inp[1]) ? node1460 : node1455;
											assign node1455 = (inp[0]) ? 3'b010 : node1456;
												assign node1456 = (inp[9]) ? 3'b010 : 3'b011;
											assign node1460 = (inp[0]) ? node1462 : 3'b010;
												assign node1462 = (inp[9]) ? 3'b011 : 3'b010;
									assign node1465 = (inp[0]) ? node1477 : node1466;
										assign node1466 = (inp[9]) ? node1472 : node1467;
											assign node1467 = (inp[1]) ? node1469 : 3'b000;
												assign node1469 = (inp[2]) ? 3'b001 : 3'b000;
											assign node1472 = (inp[2]) ? node1474 : 3'b001;
												assign node1474 = (inp[1]) ? 3'b000 : 3'b001;
										assign node1477 = (inp[9]) ? 3'b000 : node1478;
											assign node1478 = (inp[2]) ? 3'b000 : 3'b001;
								assign node1482 = (inp[11]) ? node1500 : node1483;
									assign node1483 = (inp[9]) ? node1495 : node1484;
										assign node1484 = (inp[0]) ? node1490 : node1485;
											assign node1485 = (inp[2]) ? node1487 : 3'b000;
												assign node1487 = (inp[1]) ? 3'b001 : 3'b000;
											assign node1490 = (inp[1]) ? node1492 : 3'b001;
												assign node1492 = (inp[2]) ? 3'b000 : 3'b001;
										assign node1495 = (inp[0]) ? 3'b000 : node1496;
											assign node1496 = (inp[2]) ? 3'b000 : 3'b001;
									assign node1500 = (inp[9]) ? node1512 : node1501;
										assign node1501 = (inp[0]) ? node1507 : node1502;
											assign node1502 = (inp[1]) ? node1504 : 3'b001;
												assign node1504 = (inp[2]) ? 3'b000 : 3'b001;
											assign node1507 = (inp[1]) ? node1509 : 3'b000;
												assign node1509 = (inp[2]) ? 3'b001 : 3'b000;
										assign node1512 = (inp[2]) ? 3'b001 : node1513;
											assign node1513 = (inp[0]) ? 3'b001 : 3'b000;
							assign node1517 = (inp[11]) ? node1551 : node1518;
								assign node1518 = (inp[7]) ? node1532 : node1519;
									assign node1519 = (inp[9]) ? node1529 : node1520;
										assign node1520 = (inp[1]) ? node1526 : node1521;
											assign node1521 = (inp[0]) ? node1523 : 3'b001;
												assign node1523 = (inp[2]) ? 3'b001 : 3'b000;
											assign node1526 = (inp[0]) ? 3'b001 : 3'b000;
										assign node1529 = (inp[0]) ? 3'b000 : 3'b001;
									assign node1532 = (inp[2]) ? node1540 : node1533;
										assign node1533 = (inp[0]) ? 3'b011 : node1534;
											assign node1534 = (inp[1]) ? 3'b010 : node1535;
												assign node1535 = (inp[9]) ? 3'b010 : 3'b011;
										assign node1540 = (inp[1]) ? node1546 : node1541;
											assign node1541 = (inp[9]) ? node1543 : 3'b010;
												assign node1543 = (inp[0]) ? 3'b010 : 3'b011;
											assign node1546 = (inp[0]) ? node1548 : 3'b010;
												assign node1548 = (inp[9]) ? 3'b010 : 3'b011;
								assign node1551 = (inp[7]) ? node1567 : node1552;
									assign node1552 = (inp[1]) ? node1560 : node1553;
										assign node1553 = (inp[0]) ? 3'b010 : node1554;
											assign node1554 = (inp[9]) ? node1556 : 3'b010;
												assign node1556 = (inp[2]) ? 3'b010 : 3'b011;
										assign node1560 = (inp[0]) ? node1564 : node1561;
											assign node1561 = (inp[9]) ? 3'b010 : 3'b011;
											assign node1564 = (inp[9]) ? 3'b011 : 3'b010;
									assign node1567 = (inp[1]) ? node1577 : node1568;
										assign node1568 = (inp[9]) ? 3'b011 : node1569;
											assign node1569 = (inp[2]) ? node1573 : node1570;
												assign node1570 = (inp[0]) ? 3'b010 : 3'b011;
												assign node1573 = (inp[0]) ? 3'b011 : 3'b010;
										assign node1577 = (inp[2]) ? node1585 : node1578;
											assign node1578 = (inp[9]) ? node1582 : node1579;
												assign node1579 = (inp[0]) ? 3'b011 : 3'b010;
												assign node1582 = (inp[0]) ? 3'b010 : 3'b011;
											assign node1585 = (inp[0]) ? node1589 : node1586;
												assign node1586 = (inp[9]) ? 3'b011 : 3'b010;
												assign node1589 = (inp[9]) ? 3'b010 : 3'b011;
						assign node1592 = (inp[7]) ? node1630 : node1593;
							assign node1593 = (inp[9]) ? node1601 : node1594;
								assign node1594 = (inp[11]) ? 3'b010 : node1595;
									assign node1595 = (inp[2]) ? 3'b010 : node1596;
										assign node1596 = (inp[10]) ? 3'b011 : 3'b010;
								assign node1601 = (inp[11]) ? 3'b011 : node1602;
									assign node1602 = (inp[0]) ? node1618 : node1603;
										assign node1603 = (inp[1]) ? node1611 : node1604;
											assign node1604 = (inp[2]) ? node1608 : node1605;
												assign node1605 = (inp[10]) ? 3'b010 : 3'b011;
												assign node1608 = (inp[10]) ? 3'b011 : 3'b010;
											assign node1611 = (inp[2]) ? node1615 : node1612;
												assign node1612 = (inp[10]) ? 3'b010 : 3'b011;
												assign node1615 = (inp[10]) ? 3'b011 : 3'b010;
										assign node1618 = (inp[1]) ? node1624 : node1619;
											assign node1619 = (inp[2]) ? 3'b010 : node1620;
												assign node1620 = (inp[10]) ? 3'b010 : 3'b011;
											assign node1624 = (inp[10]) ? node1626 : 3'b010;
												assign node1626 = (inp[2]) ? 3'b011 : 3'b010;
							assign node1630 = (inp[9]) ? node1636 : node1631;
								assign node1631 = (inp[11]) ? 3'b011 : node1632;
									assign node1632 = (inp[10]) ? 3'b011 : 3'b010;
								assign node1636 = (inp[10]) ? 3'b010 : node1637;
									assign node1637 = (inp[11]) ? 3'b010 : 3'b011;
					assign node1641 = (inp[8]) ? node1785 : node1642;
						assign node1642 = (inp[10]) ? node1734 : node1643;
							assign node1643 = (inp[7]) ? node1681 : node1644;
								assign node1644 = (inp[11]) ? node1660 : node1645;
									assign node1645 = (inp[0]) ? node1657 : node1646;
										assign node1646 = (inp[9]) ? node1652 : node1647;
											assign node1647 = (inp[2]) ? 3'b000 : node1648;
												assign node1648 = (inp[1]) ? 3'b000 : 3'b001;
											assign node1652 = (inp[1]) ? 3'b001 : node1653;
												assign node1653 = (inp[2]) ? 3'b001 : 3'b000;
										assign node1657 = (inp[9]) ? 3'b000 : 3'b001;
									assign node1660 = (inp[1]) ? node1674 : node1661;
										assign node1661 = (inp[0]) ? node1669 : node1662;
											assign node1662 = (inp[9]) ? node1666 : node1663;
												assign node1663 = (inp[2]) ? 3'b010 : 3'b011;
												assign node1666 = (inp[2]) ? 3'b011 : 3'b010;
											assign node1669 = (inp[2]) ? node1671 : 3'b010;
												assign node1671 = (inp[9]) ? 3'b010 : 3'b011;
										assign node1674 = (inp[0]) ? node1678 : node1675;
											assign node1675 = (inp[9]) ? 3'b011 : 3'b010;
											assign node1678 = (inp[9]) ? 3'b010 : 3'b011;
								assign node1681 = (inp[2]) ? node1711 : node1682;
									assign node1682 = (inp[11]) ? node1698 : node1683;
										assign node1683 = (inp[1]) ? node1691 : node1684;
											assign node1684 = (inp[0]) ? node1688 : node1685;
												assign node1685 = (inp[9]) ? 3'b011 : 3'b010;
												assign node1688 = (inp[9]) ? 3'b010 : 3'b011;
											assign node1691 = (inp[0]) ? node1695 : node1692;
												assign node1692 = (inp[9]) ? 3'b010 : 3'b011;
												assign node1695 = (inp[9]) ? 3'b011 : 3'b010;
										assign node1698 = (inp[0]) ? node1706 : node1699;
											assign node1699 = (inp[1]) ? node1703 : node1700;
												assign node1700 = (inp[9]) ? 3'b010 : 3'b011;
												assign node1703 = (inp[9]) ? 3'b011 : 3'b010;
											assign node1706 = (inp[9]) ? node1708 : 3'b010;
												assign node1708 = (inp[1]) ? 3'b010 : 3'b011;
									assign node1711 = (inp[1]) ? node1721 : node1712;
										assign node1712 = (inp[11]) ? 3'b011 : node1713;
											assign node1713 = (inp[9]) ? node1717 : node1714;
												assign node1714 = (inp[0]) ? 3'b010 : 3'b011;
												assign node1717 = (inp[0]) ? 3'b011 : 3'b010;
										assign node1721 = (inp[0]) ? node1727 : node1722;
											assign node1722 = (inp[9]) ? 3'b011 : node1723;
												assign node1723 = (inp[11]) ? 3'b010 : 3'b011;
											assign node1727 = (inp[9]) ? node1731 : node1728;
												assign node1728 = (inp[11]) ? 3'b011 : 3'b010;
												assign node1731 = (inp[11]) ? 3'b010 : 3'b011;
							assign node1734 = (inp[7]) ? node1762 : node1735;
								assign node1735 = (inp[11]) ? node1747 : node1736;
									assign node1736 = (inp[9]) ? node1742 : node1737;
										assign node1737 = (inp[0]) ? 3'b010 : node1738;
											assign node1738 = (inp[1]) ? 3'b010 : 3'b011;
										assign node1742 = (inp[0]) ? 3'b011 : node1743;
											assign node1743 = (inp[2]) ? 3'b011 : 3'b010;
									assign node1747 = (inp[1]) ? node1755 : node1748;
										assign node1748 = (inp[0]) ? node1750 : 3'b000;
											assign node1750 = (inp[9]) ? 3'b000 : node1751;
												assign node1751 = (inp[2]) ? 3'b001 : 3'b000;
										assign node1755 = (inp[9]) ? node1759 : node1756;
											assign node1756 = (inp[0]) ? 3'b001 : 3'b000;
											assign node1759 = (inp[0]) ? 3'b000 : 3'b001;
								assign node1762 = (inp[0]) ? node1774 : node1763;
									assign node1763 = (inp[9]) ? node1769 : node1764;
										assign node1764 = (inp[1]) ? 3'b000 : node1765;
											assign node1765 = (inp[2]) ? 3'b000 : 3'b001;
										assign node1769 = (inp[1]) ? 3'b001 : node1770;
											assign node1770 = (inp[2]) ? 3'b001 : 3'b000;
									assign node1774 = (inp[9]) ? node1780 : node1775;
										assign node1775 = (inp[1]) ? 3'b001 : node1776;
											assign node1776 = (inp[2]) ? 3'b001 : 3'b000;
										assign node1780 = (inp[1]) ? 3'b000 : node1781;
											assign node1781 = (inp[2]) ? 3'b000 : 3'b001;
						assign node1785 = (inp[9]) ? node1799 : node1786;
							assign node1786 = (inp[11]) ? 3'b001 : node1787;
								assign node1787 = (inp[10]) ? node1793 : node1788;
									assign node1788 = (inp[7]) ? 3'b000 : node1789;
										assign node1789 = (inp[2]) ? 3'b000 : 3'b001;
									assign node1793 = (inp[7]) ? 3'b001 : node1794;
										assign node1794 = (inp[2]) ? 3'b001 : 3'b000;
							assign node1799 = (inp[11]) ? 3'b000 : node1800;
								assign node1800 = (inp[10]) ? node1806 : node1801;
									assign node1801 = (inp[2]) ? 3'b001 : node1802;
										assign node1802 = (inp[7]) ? 3'b001 : 3'b000;
									assign node1806 = (inp[7]) ? 3'b000 : node1807;
										assign node1807 = (inp[2]) ? 3'b000 : 3'b001;
		assign node1812 = (inp[8]) ? node2560 : node1813;
			assign node1813 = (inp[5]) ? node2375 : node1814;
				assign node1814 = (inp[6]) ? node2068 : node1815;
					assign node1815 = (inp[7]) ? node1915 : node1816;
						assign node1816 = (inp[11]) ? node1858 : node1817;
							assign node1817 = (inp[10]) ? node1835 : node1818;
								assign node1818 = (inp[2]) ? node1830 : node1819;
									assign node1819 = (inp[0]) ? node1825 : node1820;
										assign node1820 = (inp[9]) ? 3'b100 : node1821;
											assign node1821 = (inp[3]) ? 3'b101 : 3'b100;
										assign node1825 = (inp[9]) ? 3'b101 : node1826;
											assign node1826 = (inp[1]) ? 3'b100 : 3'b101;
									assign node1830 = (inp[0]) ? 3'b100 : node1831;
										assign node1831 = (inp[1]) ? 3'b100 : 3'b101;
								assign node1835 = (inp[2]) ? node1847 : node1836;
									assign node1836 = (inp[0]) ? node1842 : node1837;
										assign node1837 = (inp[3]) ? node1839 : 3'b110;
											assign node1839 = (inp[9]) ? 3'b110 : 3'b111;
										assign node1842 = (inp[3]) ? node1844 : 3'b111;
											assign node1844 = (inp[1]) ? 3'b110 : 3'b111;
									assign node1847 = (inp[0]) ? node1853 : node1848;
										assign node1848 = (inp[1]) ? node1850 : 3'b111;
											assign node1850 = (inp[3]) ? 3'b110 : 3'b111;
										assign node1853 = (inp[1]) ? node1855 : 3'b110;
											assign node1855 = (inp[3]) ? 3'b111 : 3'b110;
							assign node1858 = (inp[10]) ? node1894 : node1859;
								assign node1859 = (inp[9]) ? node1875 : node1860;
									assign node1860 = (inp[2]) ? node1868 : node1861;
										assign node1861 = (inp[1]) ? node1863 : 3'b111;
											assign node1863 = (inp[0]) ? node1865 : 3'b111;
												assign node1865 = (inp[3]) ? 3'b110 : 3'b111;
										assign node1868 = (inp[3]) ? node1872 : node1869;
											assign node1869 = (inp[0]) ? 3'b110 : 3'b111;
											assign node1872 = (inp[0]) ? 3'b111 : 3'b110;
									assign node1875 = (inp[2]) ? node1883 : node1876;
										assign node1876 = (inp[3]) ? node1878 : 3'b110;
											assign node1878 = (inp[0]) ? 3'b111 : node1879;
												assign node1879 = (inp[1]) ? 3'b111 : 3'b110;
										assign node1883 = (inp[0]) ? node1889 : node1884;
											assign node1884 = (inp[1]) ? node1886 : 3'b111;
												assign node1886 = (inp[3]) ? 3'b110 : 3'b111;
											assign node1889 = (inp[3]) ? node1891 : 3'b110;
												assign node1891 = (inp[1]) ? 3'b111 : 3'b110;
								assign node1894 = (inp[0]) ? node1906 : node1895;
									assign node1895 = (inp[2]) ? node1901 : node1896;
										assign node1896 = (inp[1]) ? 3'b100 : node1897;
											assign node1897 = (inp[3]) ? 3'b100 : 3'b101;
										assign node1901 = (inp[1]) ? 3'b101 : node1902;
											assign node1902 = (inp[3]) ? 3'b101 : 3'b100;
									assign node1906 = (inp[2]) ? node1910 : node1907;
										assign node1907 = (inp[3]) ? 3'b101 : 3'b100;
										assign node1910 = (inp[3]) ? 3'b100 : node1911;
											assign node1911 = (inp[1]) ? 3'b100 : 3'b101;
						assign node1915 = (inp[9]) ? node1995 : node1916;
							assign node1916 = (inp[10]) ? node1962 : node1917;
								assign node1917 = (inp[11]) ? node1947 : node1918;
									assign node1918 = (inp[1]) ? node1932 : node1919;
										assign node1919 = (inp[2]) ? node1927 : node1920;
											assign node1920 = (inp[0]) ? node1924 : node1921;
												assign node1921 = (inp[3]) ? 3'b101 : 3'b100;
												assign node1924 = (inp[3]) ? 3'b100 : 3'b101;
											assign node1927 = (inp[3]) ? 3'b100 : node1928;
												assign node1928 = (inp[0]) ? 3'b100 : 3'b101;
										assign node1932 = (inp[3]) ? node1940 : node1933;
											assign node1933 = (inp[0]) ? node1937 : node1934;
												assign node1934 = (inp[2]) ? 3'b101 : 3'b100;
												assign node1937 = (inp[2]) ? 3'b100 : 3'b101;
											assign node1940 = (inp[2]) ? node1944 : node1941;
												assign node1941 = (inp[0]) ? 3'b101 : 3'b100;
												assign node1944 = (inp[0]) ? 3'b100 : 3'b101;
									assign node1947 = (inp[3]) ? node1957 : node1948;
										assign node1948 = (inp[2]) ? 3'b110 : node1949;
											assign node1949 = (inp[1]) ? node1953 : node1950;
												assign node1950 = (inp[0]) ? 3'b111 : 3'b110;
												assign node1953 = (inp[0]) ? 3'b110 : 3'b111;
										assign node1957 = (inp[0]) ? node1959 : 3'b111;
											assign node1959 = (inp[2]) ? 3'b110 : 3'b111;
								assign node1962 = (inp[11]) ? node1976 : node1963;
									assign node1963 = (inp[0]) ? node1969 : node1964;
										assign node1964 = (inp[2]) ? 3'b111 : node1965;
											assign node1965 = (inp[3]) ? 3'b111 : 3'b110;
										assign node1969 = (inp[2]) ? node1971 : 3'b111;
											assign node1971 = (inp[3]) ? node1973 : 3'b110;
												assign node1973 = (inp[1]) ? 3'b110 : 3'b111;
									assign node1976 = (inp[3]) ? node1986 : node1977;
										assign node1977 = (inp[1]) ? node1979 : 3'b101;
											assign node1979 = (inp[2]) ? node1983 : node1980;
												assign node1980 = (inp[0]) ? 3'b101 : 3'b100;
												assign node1983 = (inp[0]) ? 3'b100 : 3'b101;
										assign node1986 = (inp[2]) ? 3'b100 : node1987;
											assign node1987 = (inp[1]) ? node1991 : node1988;
												assign node1988 = (inp[0]) ? 3'b100 : 3'b101;
												assign node1991 = (inp[0]) ? 3'b101 : 3'b100;
							assign node1995 = (inp[10]) ? node2029 : node1996;
								assign node1996 = (inp[11]) ? node2016 : node1997;
									assign node1997 = (inp[2]) ? node2007 : node1998;
										assign node1998 = (inp[1]) ? node2004 : node1999;
											assign node1999 = (inp[3]) ? node2001 : 3'b101;
												assign node2001 = (inp[0]) ? 3'b100 : 3'b101;
											assign node2004 = (inp[0]) ? 3'b101 : 3'b100;
										assign node2007 = (inp[0]) ? node2013 : node2008;
											assign node2008 = (inp[1]) ? 3'b101 : node2009;
												assign node2009 = (inp[3]) ? 3'b100 : 3'b101;
											assign node2013 = (inp[1]) ? 3'b100 : 3'b101;
									assign node2016 = (inp[2]) ? node2020 : node2017;
										assign node2017 = (inp[0]) ? 3'b111 : 3'b110;
										assign node2020 = (inp[0]) ? node2026 : node2021;
											assign node2021 = (inp[1]) ? node2023 : 3'b111;
												assign node2023 = (inp[3]) ? 3'b111 : 3'b110;
											assign node2026 = (inp[1]) ? 3'b111 : 3'b110;
								assign node2029 = (inp[11]) ? node2045 : node2030;
									assign node2030 = (inp[0]) ? node2040 : node2031;
										assign node2031 = (inp[3]) ? node2033 : 3'b111;
											assign node2033 = (inp[2]) ? node2037 : node2034;
												assign node2034 = (inp[1]) ? 3'b110 : 3'b111;
												assign node2037 = (inp[1]) ? 3'b111 : 3'b110;
										assign node2040 = (inp[2]) ? 3'b110 : node2041;
											assign node2041 = (inp[1]) ? 3'b111 : 3'b110;
									assign node2045 = (inp[1]) ? node2055 : node2046;
										assign node2046 = (inp[2]) ? node2048 : 3'b100;
											assign node2048 = (inp[3]) ? node2052 : node2049;
												assign node2049 = (inp[0]) ? 3'b100 : 3'b101;
												assign node2052 = (inp[0]) ? 3'b101 : 3'b100;
										assign node2055 = (inp[3]) ? node2061 : node2056;
											assign node2056 = (inp[2]) ? node2058 : 3'b101;
												assign node2058 = (inp[0]) ? 3'b100 : 3'b101;
											assign node2061 = (inp[0]) ? node2065 : node2062;
												assign node2062 = (inp[2]) ? 3'b101 : 3'b100;
												assign node2065 = (inp[2]) ? 3'b100 : 3'b101;
					assign node2068 = (inp[9]) ? node2258 : node2069;
						assign node2069 = (inp[3]) ? node2171 : node2070;
							assign node2070 = (inp[1]) ? node2116 : node2071;
								assign node2071 = (inp[10]) ? node2093 : node2072;
									assign node2072 = (inp[11]) ? node2084 : node2073;
										assign node2073 = (inp[7]) ? node2079 : node2074;
											assign node2074 = (inp[0]) ? 3'b100 : node2075;
												assign node2075 = (inp[2]) ? 3'b101 : 3'b100;
											assign node2079 = (inp[0]) ? node2081 : 3'b100;
												assign node2081 = (inp[2]) ? 3'b100 : 3'b101;
										assign node2084 = (inp[7]) ? node2086 : 3'b110;
											assign node2086 = (inp[0]) ? node2090 : node2087;
												assign node2087 = (inp[2]) ? 3'b110 : 3'b111;
												assign node2090 = (inp[2]) ? 3'b111 : 3'b110;
									assign node2093 = (inp[11]) ? node2107 : node2094;
										assign node2094 = (inp[7]) ? node2102 : node2095;
											assign node2095 = (inp[0]) ? node2099 : node2096;
												assign node2096 = (inp[2]) ? 3'b111 : 3'b110;
												assign node2099 = (inp[2]) ? 3'b110 : 3'b111;
											assign node2102 = (inp[0]) ? 3'b111 : node2103;
												assign node2103 = (inp[2]) ? 3'b110 : 3'b111;
										assign node2107 = (inp[2]) ? node2109 : 3'b100;
											assign node2109 = (inp[7]) ? node2113 : node2110;
												assign node2110 = (inp[0]) ? 3'b100 : 3'b101;
												assign node2113 = (inp[0]) ? 3'b101 : 3'b100;
								assign node2116 = (inp[7]) ? node2146 : node2117;
									assign node2117 = (inp[0]) ? node2131 : node2118;
										assign node2118 = (inp[2]) ? node2126 : node2119;
											assign node2119 = (inp[10]) ? node2123 : node2120;
												assign node2120 = (inp[11]) ? 3'b111 : 3'b101;
												assign node2123 = (inp[11]) ? 3'b101 : 3'b110;
											assign node2126 = (inp[10]) ? 3'b111 : node2127;
												assign node2127 = (inp[11]) ? 3'b110 : 3'b100;
										assign node2131 = (inp[2]) ? node2139 : node2132;
											assign node2132 = (inp[10]) ? node2136 : node2133;
												assign node2133 = (inp[11]) ? 3'b110 : 3'b100;
												assign node2136 = (inp[11]) ? 3'b100 : 3'b111;
											assign node2139 = (inp[10]) ? node2143 : node2140;
												assign node2140 = (inp[11]) ? 3'b111 : 3'b101;
												assign node2143 = (inp[11]) ? 3'b101 : 3'b110;
									assign node2146 = (inp[0]) ? node2160 : node2147;
										assign node2147 = (inp[2]) ? node2155 : node2148;
											assign node2148 = (inp[10]) ? node2152 : node2149;
												assign node2149 = (inp[11]) ? 3'b110 : 3'b100;
												assign node2152 = (inp[11]) ? 3'b100 : 3'b110;
											assign node2155 = (inp[11]) ? 3'b111 : node2156;
												assign node2156 = (inp[10]) ? 3'b111 : 3'b101;
										assign node2160 = (inp[2]) ? node2166 : node2161;
											assign node2161 = (inp[10]) ? node2163 : 3'b111;
												assign node2163 = (inp[11]) ? 3'b101 : 3'b111;
											assign node2166 = (inp[11]) ? node2168 : 3'b110;
												assign node2168 = (inp[10]) ? 3'b100 : 3'b110;
							assign node2171 = (inp[1]) ? node2211 : node2172;
								assign node2172 = (inp[10]) ? node2190 : node2173;
									assign node2173 = (inp[11]) ? node2175 : 3'b101;
										assign node2175 = (inp[7]) ? node2183 : node2176;
											assign node2176 = (inp[0]) ? node2180 : node2177;
												assign node2177 = (inp[2]) ? 3'b111 : 3'b110;
												assign node2180 = (inp[2]) ? 3'b110 : 3'b111;
											assign node2183 = (inp[0]) ? node2187 : node2184;
												assign node2184 = (inp[2]) ? 3'b111 : 3'b110;
												assign node2187 = (inp[2]) ? 3'b110 : 3'b111;
									assign node2190 = (inp[11]) ? node2204 : node2191;
										assign node2191 = (inp[7]) ? node2197 : node2192;
											assign node2192 = (inp[2]) ? node2194 : 3'b111;
												assign node2194 = (inp[0]) ? 3'b111 : 3'b110;
											assign node2197 = (inp[0]) ? node2201 : node2198;
												assign node2198 = (inp[2]) ? 3'b111 : 3'b110;
												assign node2201 = (inp[2]) ? 3'b110 : 3'b111;
										assign node2204 = (inp[0]) ? node2208 : node2205;
											assign node2205 = (inp[2]) ? 3'b101 : 3'b100;
											assign node2208 = (inp[2]) ? 3'b100 : 3'b101;
								assign node2211 = (inp[0]) ? node2235 : node2212;
									assign node2212 = (inp[2]) ? node2228 : node2213;
										assign node2213 = (inp[7]) ? node2221 : node2214;
											assign node2214 = (inp[10]) ? node2218 : node2215;
												assign node2215 = (inp[11]) ? 3'b110 : 3'b100;
												assign node2218 = (inp[11]) ? 3'b100 : 3'b110;
											assign node2221 = (inp[11]) ? node2225 : node2222;
												assign node2222 = (inp[10]) ? 3'b110 : 3'b101;
												assign node2225 = (inp[10]) ? 3'b100 : 3'b110;
										assign node2228 = (inp[11]) ? node2232 : node2229;
											assign node2229 = (inp[10]) ? 3'b111 : 3'b100;
											assign node2232 = (inp[10]) ? 3'b101 : 3'b111;
									assign node2235 = (inp[2]) ? node2249 : node2236;
										assign node2236 = (inp[7]) ? node2244 : node2237;
											assign node2237 = (inp[11]) ? node2241 : node2238;
												assign node2238 = (inp[10]) ? 3'b111 : 3'b101;
												assign node2241 = (inp[10]) ? 3'b101 : 3'b111;
											assign node2244 = (inp[10]) ? node2246 : 3'b100;
												assign node2246 = (inp[11]) ? 3'b101 : 3'b111;
										assign node2249 = (inp[11]) ? node2255 : node2250;
											assign node2250 = (inp[10]) ? 3'b110 : node2251;
												assign node2251 = (inp[7]) ? 3'b101 : 3'b100;
											assign node2255 = (inp[10]) ? 3'b100 : 3'b110;
						assign node2258 = (inp[10]) ? node2324 : node2259;
							assign node2259 = (inp[11]) ? node2295 : node2260;
								assign node2260 = (inp[3]) ? node2276 : node2261;
									assign node2261 = (inp[1]) ? node2269 : node2262;
										assign node2262 = (inp[2]) ? node2266 : node2263;
											assign node2263 = (inp[0]) ? 3'b101 : 3'b100;
											assign node2266 = (inp[0]) ? 3'b100 : 3'b101;
										assign node2269 = (inp[0]) ? node2271 : 3'b101;
											assign node2271 = (inp[2]) ? node2273 : 3'b101;
												assign node2273 = (inp[7]) ? 3'b100 : 3'b101;
									assign node2276 = (inp[7]) ? node2286 : node2277;
										assign node2277 = (inp[1]) ? node2279 : 3'b101;
											assign node2279 = (inp[0]) ? node2283 : node2280;
												assign node2280 = (inp[2]) ? 3'b101 : 3'b100;
												assign node2283 = (inp[2]) ? 3'b100 : 3'b101;
										assign node2286 = (inp[1]) ? node2288 : 3'b100;
											assign node2288 = (inp[0]) ? node2292 : node2289;
												assign node2289 = (inp[2]) ? 3'b100 : 3'b101;
												assign node2292 = (inp[2]) ? 3'b101 : 3'b100;
								assign node2295 = (inp[2]) ? node2311 : node2296;
									assign node2296 = (inp[0]) ? node2302 : node2297;
										assign node2297 = (inp[1]) ? 3'b110 : node2298;
											assign node2298 = (inp[7]) ? 3'b111 : 3'b110;
										assign node2302 = (inp[3]) ? 3'b111 : node2303;
											assign node2303 = (inp[7]) ? node2307 : node2304;
												assign node2304 = (inp[1]) ? 3'b110 : 3'b111;
												assign node2307 = (inp[1]) ? 3'b111 : 3'b110;
									assign node2311 = (inp[0]) ? node2317 : node2312;
										assign node2312 = (inp[1]) ? 3'b111 : node2313;
											assign node2313 = (inp[7]) ? 3'b110 : 3'b111;
										assign node2317 = (inp[3]) ? 3'b110 : node2318;
											assign node2318 = (inp[7]) ? node2320 : 3'b110;
												assign node2320 = (inp[1]) ? 3'b110 : 3'b111;
							assign node2324 = (inp[11]) ? node2350 : node2325;
								assign node2325 = (inp[7]) ? node2337 : node2326;
									assign node2326 = (inp[2]) ? node2332 : node2327;
										assign node2327 = (inp[0]) ? 3'b111 : node2328;
											assign node2328 = (inp[3]) ? 3'b111 : 3'b110;
										assign node2332 = (inp[0]) ? 3'b110 : node2333;
											assign node2333 = (inp[1]) ? 3'b111 : 3'b110;
									assign node2337 = (inp[2]) ? node2345 : node2338;
										assign node2338 = (inp[0]) ? node2340 : 3'b110;
											assign node2340 = (inp[1]) ? 3'b111 : node2341;
												assign node2341 = (inp[3]) ? 3'b111 : 3'b110;
										assign node2345 = (inp[0]) ? node2347 : 3'b111;
											assign node2347 = (inp[3]) ? 3'b110 : 3'b111;
								assign node2350 = (inp[0]) ? node2366 : node2351;
									assign node2351 = (inp[2]) ? node2359 : node2352;
										assign node2352 = (inp[3]) ? 3'b100 : node2353;
											assign node2353 = (inp[1]) ? 3'b100 : node2354;
												assign node2354 = (inp[7]) ? 3'b101 : 3'b100;
										assign node2359 = (inp[3]) ? 3'b101 : node2360;
											assign node2360 = (inp[7]) ? 3'b101 : node2361;
												assign node2361 = (inp[1]) ? 3'b100 : 3'b101;
									assign node2366 = (inp[2]) ? node2368 : 3'b101;
										assign node2368 = (inp[3]) ? 3'b100 : node2369;
											assign node2369 = (inp[1]) ? node2371 : 3'b101;
												assign node2371 = (inp[7]) ? 3'b100 : 3'b101;
				assign node2375 = (inp[10]) ? node2485 : node2376;
					assign node2376 = (inp[6]) ? node2442 : node2377;
						assign node2377 = (inp[7]) ? node2419 : node2378;
							assign node2378 = (inp[9]) ? node2396 : node2379;
								assign node2379 = (inp[0]) ? node2387 : node2380;
									assign node2380 = (inp[3]) ? node2382 : 3'b000;
										assign node2382 = (inp[11]) ? node2384 : 3'b001;
											assign node2384 = (inp[1]) ? 3'b000 : 3'b001;
									assign node2387 = (inp[3]) ? node2393 : node2388;
										assign node2388 = (inp[11]) ? node2390 : 3'b001;
											assign node2390 = (inp[1]) ? 3'b000 : 3'b001;
										assign node2393 = (inp[1]) ? 3'b001 : 3'b000;
								assign node2396 = (inp[0]) ? node2408 : node2397;
									assign node2397 = (inp[3]) ? node2403 : node2398;
										assign node2398 = (inp[1]) ? node2400 : 3'b000;
											assign node2400 = (inp[11]) ? 3'b001 : 3'b000;
										assign node2403 = (inp[11]) ? node2405 : 3'b001;
											assign node2405 = (inp[1]) ? 3'b000 : 3'b001;
									assign node2408 = (inp[3]) ? node2414 : node2409;
										assign node2409 = (inp[1]) ? node2411 : 3'b001;
											assign node2411 = (inp[11]) ? 3'b000 : 3'b001;
										assign node2414 = (inp[1]) ? node2416 : 3'b000;
											assign node2416 = (inp[11]) ? 3'b001 : 3'b000;
							assign node2419 = (inp[3]) ? node2427 : node2420;
								assign node2420 = (inp[11]) ? node2424 : node2421;
									assign node2421 = (inp[0]) ? 3'b011 : 3'b010;
									assign node2424 = (inp[0]) ? 3'b010 : 3'b011;
								assign node2427 = (inp[9]) ? node2435 : node2428;
									assign node2428 = (inp[0]) ? node2432 : node2429;
										assign node2429 = (inp[11]) ? 3'b011 : 3'b010;
										assign node2432 = (inp[11]) ? 3'b010 : 3'b011;
									assign node2435 = (inp[11]) ? node2439 : node2436;
										assign node2436 = (inp[0]) ? 3'b011 : 3'b010;
										assign node2439 = (inp[0]) ? 3'b010 : 3'b011;
						assign node2442 = (inp[3]) ? node2466 : node2443;
							assign node2443 = (inp[0]) ? node2453 : node2444;
								assign node2444 = (inp[7]) ? node2450 : node2445;
									assign node2445 = (inp[11]) ? 3'b010 : node2446;
										assign node2446 = (inp[1]) ? 3'b011 : 3'b010;
									assign node2450 = (inp[11]) ? 3'b011 : 3'b010;
								assign node2453 = (inp[1]) ? node2459 : node2454;
									assign node2454 = (inp[7]) ? node2456 : 3'b011;
										assign node2456 = (inp[11]) ? 3'b010 : 3'b011;
									assign node2459 = (inp[11]) ? node2463 : node2460;
										assign node2460 = (inp[7]) ? 3'b011 : 3'b010;
										assign node2463 = (inp[7]) ? 3'b010 : 3'b011;
							assign node2466 = (inp[7]) ? node2478 : node2467;
								assign node2467 = (inp[0]) ? node2473 : node2468;
									assign node2468 = (inp[1]) ? node2470 : 3'b011;
										assign node2470 = (inp[11]) ? 3'b011 : 3'b010;
									assign node2473 = (inp[11]) ? 3'b010 : node2474;
										assign node2474 = (inp[1]) ? 3'b011 : 3'b010;
								assign node2478 = (inp[0]) ? node2482 : node2479;
									assign node2479 = (inp[11]) ? 3'b011 : 3'b010;
									assign node2482 = (inp[11]) ? 3'b010 : 3'b011;
					assign node2485 = (inp[6]) ? node2533 : node2486;
						assign node2486 = (inp[7]) ? node2510 : node2487;
							assign node2487 = (inp[0]) ? node2499 : node2488;
								assign node2488 = (inp[3]) ? node2494 : node2489;
									assign node2489 = (inp[11]) ? node2491 : 3'b010;
										assign node2491 = (inp[1]) ? 3'b010 : 3'b011;
									assign node2494 = (inp[1]) ? 3'b011 : node2495;
										assign node2495 = (inp[11]) ? 3'b010 : 3'b011;
								assign node2499 = (inp[3]) ? node2505 : node2500;
									assign node2500 = (inp[1]) ? 3'b011 : node2501;
										assign node2501 = (inp[11]) ? 3'b010 : 3'b011;
									assign node2505 = (inp[1]) ? 3'b010 : node2506;
										assign node2506 = (inp[11]) ? 3'b011 : 3'b010;
							assign node2510 = (inp[2]) ? node2518 : node2511;
								assign node2511 = (inp[1]) ? node2515 : node2512;
									assign node2512 = (inp[0]) ? 3'b001 : 3'b000;
									assign node2515 = (inp[0]) ? 3'b000 : 3'b001;
								assign node2518 = (inp[11]) ? node2526 : node2519;
									assign node2519 = (inp[0]) ? node2523 : node2520;
										assign node2520 = (inp[1]) ? 3'b001 : 3'b000;
										assign node2523 = (inp[1]) ? 3'b000 : 3'b001;
									assign node2526 = (inp[0]) ? node2530 : node2527;
										assign node2527 = (inp[1]) ? 3'b001 : 3'b000;
										assign node2530 = (inp[1]) ? 3'b000 : 3'b001;
						assign node2533 = (inp[0]) ? node2547 : node2534;
							assign node2534 = (inp[7]) ? 3'b001 : node2535;
								assign node2535 = (inp[3]) ? node2541 : node2536;
									assign node2536 = (inp[1]) ? 3'b000 : node2537;
										assign node2537 = (inp[11]) ? 3'b000 : 3'b001;
									assign node2541 = (inp[1]) ? 3'b001 : node2542;
										assign node2542 = (inp[11]) ? 3'b001 : 3'b000;
							assign node2547 = (inp[7]) ? 3'b000 : node2548;
								assign node2548 = (inp[3]) ? node2554 : node2549;
									assign node2549 = (inp[11]) ? 3'b001 : node2550;
										assign node2550 = (inp[1]) ? 3'b001 : 3'b000;
									assign node2554 = (inp[1]) ? 3'b000 : node2555;
										assign node2555 = (inp[11]) ? 3'b000 : 3'b001;
			assign node2560 = (inp[7]) ? node2834 : node2561;
				assign node2561 = (inp[6]) ? node2741 : node2562;
					assign node2562 = (inp[11]) ? node2672 : node2563;
						assign node2563 = (inp[5]) ? node2635 : node2564;
							assign node2564 = (inp[0]) ? node2598 : node2565;
								assign node2565 = (inp[10]) ? node2573 : node2566;
									assign node2566 = (inp[1]) ? node2570 : node2567;
										assign node2567 = (inp[2]) ? 3'b001 : 3'b000;
										assign node2570 = (inp[2]) ? 3'b000 : 3'b001;
									assign node2573 = (inp[2]) ? node2583 : node2574;
										assign node2574 = (inp[9]) ? 3'b000 : node2575;
											assign node2575 = (inp[3]) ? node2579 : node2576;
												assign node2576 = (inp[1]) ? 3'b001 : 3'b000;
												assign node2579 = (inp[1]) ? 3'b000 : 3'b001;
										assign node2583 = (inp[9]) ? node2591 : node2584;
											assign node2584 = (inp[3]) ? node2588 : node2585;
												assign node2585 = (inp[1]) ? 3'b000 : 3'b001;
												assign node2588 = (inp[1]) ? 3'b001 : 3'b000;
											assign node2591 = (inp[1]) ? node2595 : node2592;
												assign node2592 = (inp[3]) ? 3'b000 : 3'b001;
												assign node2595 = (inp[3]) ? 3'b001 : 3'b000;
								assign node2598 = (inp[9]) ? node2620 : node2599;
									assign node2599 = (inp[3]) ? node2605 : node2600;
										assign node2600 = (inp[2]) ? node2602 : 3'b000;
											assign node2602 = (inp[1]) ? 3'b000 : 3'b001;
										assign node2605 = (inp[2]) ? node2613 : node2606;
											assign node2606 = (inp[10]) ? node2610 : node2607;
												assign node2607 = (inp[1]) ? 3'b001 : 3'b000;
												assign node2610 = (inp[1]) ? 3'b000 : 3'b001;
											assign node2613 = (inp[10]) ? node2617 : node2614;
												assign node2614 = (inp[1]) ? 3'b000 : 3'b001;
												assign node2617 = (inp[1]) ? 3'b001 : 3'b000;
									assign node2620 = (inp[2]) ? node2628 : node2621;
										assign node2621 = (inp[10]) ? node2623 : 3'b001;
											assign node2623 = (inp[3]) ? node2625 : 3'b001;
												assign node2625 = (inp[1]) ? 3'b000 : 3'b001;
										assign node2628 = (inp[1]) ? node2632 : node2629;
											assign node2629 = (inp[10]) ? 3'b000 : 3'b001;
											assign node2632 = (inp[10]) ? 3'b001 : 3'b000;
							assign node2635 = (inp[2]) ? node2655 : node2636;
								assign node2636 = (inp[0]) ? node2642 : node2637;
									assign node2637 = (inp[3]) ? node2639 : 3'b011;
										assign node2639 = (inp[1]) ? 3'b010 : 3'b011;
									assign node2642 = (inp[9]) ? node2648 : node2643;
										assign node2643 = (inp[3]) ? 3'b011 : node2644;
											assign node2644 = (inp[1]) ? 3'b011 : 3'b010;
										assign node2648 = (inp[1]) ? node2652 : node2649;
											assign node2649 = (inp[3]) ? 3'b011 : 3'b010;
											assign node2652 = (inp[3]) ? 3'b010 : 3'b011;
								assign node2655 = (inp[0]) ? node2663 : node2656;
									assign node2656 = (inp[3]) ? node2660 : node2657;
										assign node2657 = (inp[1]) ? 3'b011 : 3'b010;
										assign node2660 = (inp[1]) ? 3'b010 : 3'b011;
									assign node2663 = (inp[10]) ? 3'b010 : node2664;
										assign node2664 = (inp[3]) ? node2668 : node2665;
											assign node2665 = (inp[1]) ? 3'b011 : 3'b010;
											assign node2668 = (inp[1]) ? 3'b010 : 3'b011;
						assign node2672 = (inp[0]) ? node2710 : node2673;
							assign node2673 = (inp[3]) ? node2699 : node2674;
								assign node2674 = (inp[1]) ? node2684 : node2675;
									assign node2675 = (inp[5]) ? 3'b010 : node2676;
										assign node2676 = (inp[10]) ? node2680 : node2677;
											assign node2677 = (inp[2]) ? 3'b011 : 3'b010;
											assign node2680 = (inp[2]) ? 3'b010 : 3'b011;
									assign node2684 = (inp[5]) ? 3'b011 : node2685;
										assign node2685 = (inp[9]) ? node2693 : node2686;
											assign node2686 = (inp[2]) ? node2690 : node2687;
												assign node2687 = (inp[10]) ? 3'b010 : 3'b011;
												assign node2690 = (inp[10]) ? 3'b011 : 3'b010;
											assign node2693 = (inp[2]) ? node2695 : 3'b010;
												assign node2695 = (inp[10]) ? 3'b011 : 3'b010;
								assign node2699 = (inp[1]) ? node2705 : node2700;
									assign node2700 = (inp[5]) ? 3'b011 : node2701;
										assign node2701 = (inp[2]) ? 3'b011 : 3'b010;
									assign node2705 = (inp[2]) ? 3'b010 : node2706;
										assign node2706 = (inp[5]) ? 3'b010 : 3'b011;
							assign node2710 = (inp[1]) ? node2726 : node2711;
								assign node2711 = (inp[3]) ? node2721 : node2712;
									assign node2712 = (inp[5]) ? 3'b010 : node2713;
										assign node2713 = (inp[2]) ? node2717 : node2714;
											assign node2714 = (inp[10]) ? 3'b011 : 3'b010;
											assign node2717 = (inp[10]) ? 3'b010 : 3'b011;
									assign node2721 = (inp[5]) ? 3'b011 : node2722;
										assign node2722 = (inp[2]) ? 3'b011 : 3'b010;
								assign node2726 = (inp[3]) ? node2736 : node2727;
									assign node2727 = (inp[5]) ? 3'b011 : node2728;
										assign node2728 = (inp[2]) ? node2732 : node2729;
											assign node2729 = (inp[10]) ? 3'b010 : 3'b011;
											assign node2732 = (inp[10]) ? 3'b011 : 3'b010;
									assign node2736 = (inp[5]) ? 3'b010 : node2737;
										assign node2737 = (inp[2]) ? 3'b010 : 3'b011;
					assign node2741 = (inp[5]) ? node2823 : node2742;
						assign node2742 = (inp[11]) ? node2808 : node2743;
							assign node2743 = (inp[3]) ? node2773 : node2744;
								assign node2744 = (inp[9]) ? node2756 : node2745;
									assign node2745 = (inp[0]) ? node2751 : node2746;
										assign node2746 = (inp[2]) ? node2748 : 3'b010;
											assign node2748 = (inp[10]) ? 3'b010 : 3'b011;
										assign node2751 = (inp[2]) ? 3'b010 : node2752;
											assign node2752 = (inp[10]) ? 3'b011 : 3'b010;
									assign node2756 = (inp[0]) ? node2766 : node2757;
										assign node2757 = (inp[1]) ? 3'b011 : node2758;
											assign node2758 = (inp[2]) ? node2762 : node2759;
												assign node2759 = (inp[10]) ? 3'b011 : 3'b010;
												assign node2762 = (inp[10]) ? 3'b010 : 3'b011;
										assign node2766 = (inp[2]) ? node2770 : node2767;
											assign node2767 = (inp[10]) ? 3'b011 : 3'b010;
											assign node2770 = (inp[10]) ? 3'b010 : 3'b011;
								assign node2773 = (inp[9]) ? node2795 : node2774;
									assign node2774 = (inp[0]) ? node2782 : node2775;
										assign node2775 = (inp[1]) ? 3'b011 : node2776;
											assign node2776 = (inp[2]) ? 3'b011 : node2777;
												assign node2777 = (inp[10]) ? 3'b011 : 3'b010;
										assign node2782 = (inp[1]) ? node2788 : node2783;
											assign node2783 = (inp[2]) ? node2785 : 3'b011;
												assign node2785 = (inp[10]) ? 3'b010 : 3'b011;
											assign node2788 = (inp[2]) ? node2792 : node2789;
												assign node2789 = (inp[10]) ? 3'b011 : 3'b010;
												assign node2792 = (inp[10]) ? 3'b010 : 3'b011;
									assign node2795 = (inp[0]) ? node2801 : node2796;
										assign node2796 = (inp[10]) ? 3'b010 : node2797;
											assign node2797 = (inp[2]) ? 3'b011 : 3'b010;
										assign node2801 = (inp[2]) ? node2805 : node2802;
											assign node2802 = (inp[10]) ? 3'b011 : 3'b010;
											assign node2805 = (inp[10]) ? 3'b010 : 3'b011;
							assign node2808 = (inp[1]) ? node2816 : node2809;
								assign node2809 = (inp[2]) ? node2813 : node2810;
									assign node2810 = (inp[3]) ? 3'b001 : 3'b000;
									assign node2813 = (inp[3]) ? 3'b000 : 3'b001;
								assign node2816 = (inp[2]) ? node2820 : node2817;
									assign node2817 = (inp[3]) ? 3'b001 : 3'b000;
									assign node2820 = (inp[3]) ? 3'b000 : 3'b001;
						assign node2823 = (inp[3]) ? node2829 : node2824;
							assign node2824 = (inp[10]) ? 3'b001 : node2825;
								assign node2825 = (inp[11]) ? 3'b001 : 3'b000;
							assign node2829 = (inp[11]) ? 3'b000 : node2830;
								assign node2830 = (inp[10]) ? 3'b000 : 3'b001;
				assign node2834 = (inp[5]) ? node2938 : node2835;
					assign node2835 = (inp[11]) ? node2911 : node2836;
						assign node2836 = (inp[3]) ? node2860 : node2837;
							assign node2837 = (inp[1]) ? node2849 : node2838;
								assign node2838 = (inp[2]) ? node2844 : node2839;
									assign node2839 = (inp[6]) ? node2841 : 3'b010;
										assign node2841 = (inp[10]) ? 3'b011 : 3'b010;
									assign node2844 = (inp[6]) ? node2846 : 3'b011;
										assign node2846 = (inp[10]) ? 3'b010 : 3'b011;
								assign node2849 = (inp[2]) ? node2855 : node2850;
									assign node2850 = (inp[10]) ? 3'b011 : node2851;
										assign node2851 = (inp[6]) ? 3'b010 : 3'b011;
									assign node2855 = (inp[10]) ? 3'b010 : node2856;
										assign node2856 = (inp[6]) ? 3'b011 : 3'b010;
							assign node2860 = (inp[6]) ? node2904 : node2861;
								assign node2861 = (inp[0]) ? node2883 : node2862;
									assign node2862 = (inp[2]) ? node2876 : node2863;
										assign node2863 = (inp[9]) ? node2871 : node2864;
											assign node2864 = (inp[1]) ? node2868 : node2865;
												assign node2865 = (inp[10]) ? 3'b010 : 3'b011;
												assign node2868 = (inp[10]) ? 3'b011 : 3'b010;
											assign node2871 = (inp[1]) ? node2873 : 3'b011;
												assign node2873 = (inp[10]) ? 3'b011 : 3'b010;
										assign node2876 = (inp[10]) ? node2880 : node2877;
											assign node2877 = (inp[1]) ? 3'b011 : 3'b010;
											assign node2880 = (inp[1]) ? 3'b010 : 3'b011;
									assign node2883 = (inp[2]) ? node2891 : node2884;
										assign node2884 = (inp[9]) ? node2886 : 3'b010;
											assign node2886 = (inp[1]) ? 3'b010 : node2887;
												assign node2887 = (inp[10]) ? 3'b010 : 3'b011;
										assign node2891 = (inp[9]) ? node2899 : node2892;
											assign node2892 = (inp[10]) ? node2896 : node2893;
												assign node2893 = (inp[1]) ? 3'b011 : 3'b010;
												assign node2896 = (inp[1]) ? 3'b010 : 3'b011;
											assign node2899 = (inp[10]) ? node2901 : 3'b010;
												assign node2901 = (inp[1]) ? 3'b010 : 3'b011;
								assign node2904 = (inp[2]) ? node2908 : node2905;
									assign node2905 = (inp[10]) ? 3'b011 : 3'b010;
									assign node2908 = (inp[10]) ? 3'b010 : 3'b011;
						assign node2911 = (inp[2]) ? node2925 : node2912;
							assign node2912 = (inp[6]) ? 3'b001 : node2913;
								assign node2913 = (inp[1]) ? node2919 : node2914;
									assign node2914 = (inp[3]) ? 3'b000 : node2915;
										assign node2915 = (inp[10]) ? 3'b000 : 3'b001;
									assign node2919 = (inp[3]) ? 3'b001 : node2920;
										assign node2920 = (inp[10]) ? 3'b001 : 3'b000;
							assign node2925 = (inp[6]) ? 3'b000 : node2926;
								assign node2926 = (inp[1]) ? node2932 : node2927;
									assign node2927 = (inp[3]) ? 3'b001 : node2928;
										assign node2928 = (inp[10]) ? 3'b001 : 3'b000;
									assign node2932 = (inp[3]) ? 3'b000 : node2933;
										assign node2933 = (inp[10]) ? 3'b000 : 3'b001;
					assign node2938 = (inp[6]) ? node2950 : node2939;
						assign node2939 = (inp[1]) ? node2945 : node2940;
							assign node2940 = (inp[11]) ? 3'b001 : node2941;
								assign node2941 = (inp[10]) ? 3'b001 : 3'b000;
							assign node2945 = (inp[10]) ? 3'b000 : node2946;
								assign node2946 = (inp[11]) ? 3'b000 : 3'b001;
						assign node2950 = (inp[10]) ? 3'b000 : node2951;
							assign node2951 = (inp[11]) ? 3'b000 : 3'b001;

endmodule