module dtc_split25_bm15 (
	input  wire [15-1:0] inp,
	output wire [1-1:0] outp
);

	wire [1-1:0] node1;
	wire [1-1:0] node2;
	wire [1-1:0] node3;
	wire [1-1:0] node4;
	wire [1-1:0] node5;
	wire [1-1:0] node7;
	wire [1-1:0] node9;
	wire [1-1:0] node10;
	wire [1-1:0] node12;
	wire [1-1:0] node14;
	wire [1-1:0] node16;
	wire [1-1:0] node19;
	wire [1-1:0] node20;
	wire [1-1:0] node22;
	wire [1-1:0] node25;
	wire [1-1:0] node26;
	wire [1-1:0] node28;
	wire [1-1:0] node31;
	wire [1-1:0] node32;
	wire [1-1:0] node35;
	wire [1-1:0] node36;
	wire [1-1:0] node40;
	wire [1-1:0] node41;
	wire [1-1:0] node43;
	wire [1-1:0] node44;
	wire [1-1:0] node46;
	wire [1-1:0] node48;
	wire [1-1:0] node50;
	wire [1-1:0] node53;
	wire [1-1:0] node54;
	wire [1-1:0] node56;
	wire [1-1:0] node58;
	wire [1-1:0] node61;
	wire [1-1:0] node62;
	wire [1-1:0] node64;
	wire [1-1:0] node66;
	wire [1-1:0] node69;
	wire [1-1:0] node70;
	wire [1-1:0] node74;
	wire [1-1:0] node75;
	wire [1-1:0] node77;
	wire [1-1:0] node79;
	wire [1-1:0] node81;
	wire [1-1:0] node82;
	wire [1-1:0] node84;
	wire [1-1:0] node88;
	wire [1-1:0] node89;
	wire [1-1:0] node91;
	wire [1-1:0] node92;
	wire [1-1:0] node94;
	wire [1-1:0] node96;
	wire [1-1:0] node99;
	wire [1-1:0] node100;
	wire [1-1:0] node102;
	wire [1-1:0] node105;
	wire [1-1:0] node106;
	wire [1-1:0] node110;
	wire [1-1:0] node111;
	wire [1-1:0] node112;
	wire [1-1:0] node114;
	wire [1-1:0] node116;
	wire [1-1:0] node119;
	wire [1-1:0] node120;
	wire [1-1:0] node124;
	wire [1-1:0] node125;
	wire [1-1:0] node129;
	wire [1-1:0] node130;
	wire [1-1:0] node131;
	wire [1-1:0] node133;
	wire [1-1:0] node134;
	wire [1-1:0] node136;
	wire [1-1:0] node137;
	wire [1-1:0] node139;
	wire [1-1:0] node143;
	wire [1-1:0] node144;
	wire [1-1:0] node146;
	wire [1-1:0] node148;
	wire [1-1:0] node151;
	wire [1-1:0] node153;
	wire [1-1:0] node155;
	wire [1-1:0] node156;
	wire [1-1:0] node160;
	wire [1-1:0] node161;
	wire [1-1:0] node163;
	wire [1-1:0] node165;
	wire [1-1:0] node166;
	wire [1-1:0] node168;
	wire [1-1:0] node170;
	wire [1-1:0] node173;
	wire [1-1:0] node174;
	wire [1-1:0] node176;
	wire [1-1:0] node179;
	wire [1-1:0] node182;
	wire [1-1:0] node183;
	wire [1-1:0] node185;
	wire [1-1:0] node186;
	wire [1-1:0] node188;
	wire [1-1:0] node191;
	wire [1-1:0] node192;
	wire [1-1:0] node194;
	wire [1-1:0] node198;
	wire [1-1:0] node199;
	wire [1-1:0] node200;
	wire [1-1:0] node202;
	wire [1-1:0] node204;
	wire [1-1:0] node207;
	wire [1-1:0] node208;
	wire [1-1:0] node211;
	wire [1-1:0] node214;
	wire [1-1:0] node215;
	wire [1-1:0] node219;
	wire [1-1:0] node220;
	wire [1-1:0] node221;
	wire [1-1:0] node223;
	wire [1-1:0] node225;
	wire [1-1:0] node226;
	wire [1-1:0] node228;
	wire [1-1:0] node231;
	wire [1-1:0] node232;
	wire [1-1:0] node234;
	wire [1-1:0] node238;
	wire [1-1:0] node239;
	wire [1-1:0] node240;
	wire [1-1:0] node242;
	wire [1-1:0] node244;
	wire [1-1:0] node247;
	wire [1-1:0] node248;
	wire [1-1:0] node250;
	wire [1-1:0] node253;
	wire [1-1:0] node256;
	wire [1-1:0] node257;
	wire [1-1:0] node259;
	wire [1-1:0] node260;
	wire [1-1:0] node262;
	wire [1-1:0] node265;
	wire [1-1:0] node266;
	wire [1-1:0] node270;
	wire [1-1:0] node271;
	wire [1-1:0] node272;
	wire [1-1:0] node274;
	wire [1-1:0] node279;
	wire [1-1:0] node280;
	wire [1-1:0] node281;
	wire [1-1:0] node283;
	wire [1-1:0] node285;
	wire [1-1:0] node286;
	wire [1-1:0] node290;
	wire [1-1:0] node291;
	wire [1-1:0] node293;
	wire [1-1:0] node294;
	wire [1-1:0] node296;
	wire [1-1:0] node299;
	wire [1-1:0] node300;
	wire [1-1:0] node304;
	wire [1-1:0] node305;
	wire [1-1:0] node306;
	wire [1-1:0] node308;
	wire [1-1:0] node311;
	wire [1-1:0] node312;
	wire [1-1:0] node317;
	wire [1-1:0] node318;
	wire [1-1:0] node319;
	wire [1-1:0] node321;
	wire [1-1:0] node323;
	wire [1-1:0] node324;
	wire [1-1:0] node328;
	wire [1-1:0] node329;
	wire [1-1:0] node331;
	wire [1-1:0] node332;
	wire [1-1:0] node337;
	wire [1-1:0] node338;
	wire [1-1:0] node339;
	wire [1-1:0] node340;
	wire [1-1:0] node342;
	wire [1-1:0] node348;
	wire [1-1:0] node349;
	wire [1-1:0] node350;
	wire [1-1:0] node351;
	wire [1-1:0] node353;
	wire [1-1:0] node354;
	wire [1-1:0] node356;
	wire [1-1:0] node358;
	wire [1-1:0] node361;
	wire [1-1:0] node362;
	wire [1-1:0] node364;
	wire [1-1:0] node366;
	wire [1-1:0] node368;
	wire [1-1:0] node371;
	wire [1-1:0] node372;
	wire [1-1:0] node374;
	wire [1-1:0] node377;
	wire [1-1:0] node378;
	wire [1-1:0] node382;
	wire [1-1:0] node383;
	wire [1-1:0] node385;
	wire [1-1:0] node386;
	wire [1-1:0] node388;
	wire [1-1:0] node390;
	wire [1-1:0] node392;
	wire [1-1:0] node395;
	wire [1-1:0] node396;
	wire [1-1:0] node398;
	wire [1-1:0] node401;
	wire [1-1:0] node402;
	wire [1-1:0] node405;
	wire [1-1:0] node406;
	wire [1-1:0] node410;
	wire [1-1:0] node411;
	wire [1-1:0] node413;
	wire [1-1:0] node415;
	wire [1-1:0] node416;
	wire [1-1:0] node418;
	wire [1-1:0] node421;
	wire [1-1:0] node422;
	wire [1-1:0] node426;
	wire [1-1:0] node427;
	wire [1-1:0] node428;
	wire [1-1:0] node430;
	wire [1-1:0] node433;
	wire [1-1:0] node434;
	wire [1-1:0] node436;
	wire [1-1:0] node439;
	wire [1-1:0] node440;
	wire [1-1:0] node444;
	wire [1-1:0] node445;
	wire [1-1:0] node447;
	wire [1-1:0] node448;
	wire [1-1:0] node452;
	wire [1-1:0] node453;
	wire [1-1:0] node457;
	wire [1-1:0] node458;
	wire [1-1:0] node459;
	wire [1-1:0] node461;
	wire [1-1:0] node463;
	wire [1-1:0] node465;
	wire [1-1:0] node466;
	wire [1-1:0] node468;
	wire [1-1:0] node471;
	wire [1-1:0] node474;
	wire [1-1:0] node475;
	wire [1-1:0] node477;
	wire [1-1:0] node478;
	wire [1-1:0] node480;
	wire [1-1:0] node482;
	wire [1-1:0] node485;
	wire [1-1:0] node486;
	wire [1-1:0] node488;
	wire [1-1:0] node492;
	wire [1-1:0] node493;
	wire [1-1:0] node495;
	wire [1-1:0] node496;
	wire [1-1:0] node498;
	wire [1-1:0] node502;
	wire [1-1:0] node503;
	wire [1-1:0] node504;
	wire [1-1:0] node506;
	wire [1-1:0] node509;
	wire [1-1:0] node510;
	wire [1-1:0] node515;
	wire [1-1:0] node516;
	wire [1-1:0] node517;
	wire [1-1:0] node518;
	wire [1-1:0] node519;
	wire [1-1:0] node521;
	wire [1-1:0] node525;
	wire [1-1:0] node526;
	wire [1-1:0] node528;
	wire [1-1:0] node531;
	wire [1-1:0] node532;
	wire [1-1:0] node534;
	wire [1-1:0] node538;
	wire [1-1:0] node539;
	wire [1-1:0] node541;
	wire [1-1:0] node542;
	wire [1-1:0] node544;
	wire [1-1:0] node548;
	wire [1-1:0] node549;
	wire [1-1:0] node553;
	wire [1-1:0] node554;
	wire [1-1:0] node555;
	wire [1-1:0] node557;
	wire [1-1:0] node560;
	wire [1-1:0] node561;
	wire [1-1:0] node562;
	wire [1-1:0] node563;
	wire [1-1:0] node567;
	wire [1-1:0] node568;
	wire [1-1:0] node573;
	wire [1-1:0] node574;
	wire [1-1:0] node575;
	wire [1-1:0] node578;
	wire [1-1:0] node579;
	wire [1-1:0] node580;
	wire [1-1:0] node586;
	wire [1-1:0] node587;
	wire [1-1:0] node588;
	wire [1-1:0] node589;
	wire [1-1:0] node591;
	wire [1-1:0] node593;
	wire [1-1:0] node595;
	wire [1-1:0] node596;
	wire [1-1:0] node598;
	wire [1-1:0] node601;
	wire [1-1:0] node602;
	wire [1-1:0] node606;
	wire [1-1:0] node607;
	wire [1-1:0] node609;
	wire [1-1:0] node610;
	wire [1-1:0] node612;
	wire [1-1:0] node614;
	wire [1-1:0] node617;
	wire [1-1:0] node618;
	wire [1-1:0] node620;
	wire [1-1:0] node624;
	wire [1-1:0] node625;
	wire [1-1:0] node627;
	wire [1-1:0] node628;
	wire [1-1:0] node632;
	wire [1-1:0] node633;
	wire [1-1:0] node635;
	wire [1-1:0] node636;
	wire [1-1:0] node641;
	wire [1-1:0] node642;
	wire [1-1:0] node643;
	wire [1-1:0] node645;
	wire [1-1:0] node647;
	wire [1-1:0] node648;
	wire [1-1:0] node650;
	wire [1-1:0] node654;
	wire [1-1:0] node655;
	wire [1-1:0] node656;
	wire [1-1:0] node658;
	wire [1-1:0] node660;
	wire [1-1:0] node663;
	wire [1-1:0] node665;
	wire [1-1:0] node666;
	wire [1-1:0] node670;
	wire [1-1:0] node671;
	wire [1-1:0] node672;
	wire [1-1:0] node677;
	wire [1-1:0] node678;
	wire [1-1:0] node679;
	wire [1-1:0] node681;
	wire [1-1:0] node684;
	wire [1-1:0] node685;
	wire [1-1:0] node686;
	wire [1-1:0] node688;
	wire [1-1:0] node691;
	wire [1-1:0] node692;
	wire [1-1:0] node696;
	wire [1-1:0] node697;
	wire [1-1:0] node698;
	wire [1-1:0] node703;
	wire [1-1:0] node704;
	wire [1-1:0] node705;
	wire [1-1:0] node710;
	wire [1-1:0] node711;
	wire [1-1:0] node712;
	wire [1-1:0] node713;
	wire [1-1:0] node714;
	wire [1-1:0] node716;
	wire [1-1:0] node718;
	wire [1-1:0] node720;
	wire [1-1:0] node723;
	wire [1-1:0] node724;
	wire [1-1:0] node726;
	wire [1-1:0] node728;
	wire [1-1:0] node731;
	wire [1-1:0] node732;
	wire [1-1:0] node734;
	wire [1-1:0] node737;
	wire [1-1:0] node739;
	wire [1-1:0] node742;
	wire [1-1:0] node743;
	wire [1-1:0] node745;
	wire [1-1:0] node746;
	wire [1-1:0] node748;
	wire [1-1:0] node752;
	wire [1-1:0] node753;
	wire [1-1:0] node754;
	wire [1-1:0] node756;
	wire [1-1:0] node760;
	wire [1-1:0] node761;
	wire [1-1:0] node762;
	wire [1-1:0] node767;
	wire [1-1:0] node768;
	wire [1-1:0] node769;
	wire [1-1:0] node771;
	wire [1-1:0] node772;
	wire [1-1:0] node774;
	wire [1-1:0] node778;
	wire [1-1:0] node779;
	wire [1-1:0] node781;
	wire [1-1:0] node782;
	wire [1-1:0] node787;
	wire [1-1:0] node788;
	wire [1-1:0] node789;
	wire [1-1:0] node790;
	wire [1-1:0] node792;
	wire [1-1:0] node795;
	wire [1-1:0] node796;
	wire [1-1:0] node802;
	wire [1-1:0] node803;
	wire [1-1:0] node804;
	wire [1-1:0] node805;
	wire [1-1:0] node807;
	wire [1-1:0] node809;
	wire [1-1:0] node810;
	wire [1-1:0] node814;
	wire [1-1:0] node815;
	wire [1-1:0] node816;
	wire [1-1:0] node819;
	wire [1-1:0] node820;
	wire [1-1:0] node824;
	wire [1-1:0] node825;
	wire [1-1:0] node829;
	wire [1-1:0] node830;
	wire [1-1:0] node831;
	wire [1-1:0] node833;
	wire [1-1:0] node838;
	wire [1-1:0] node839;
	wire [1-1:0] node840;
	wire [1-1:0] node841;
	wire [1-1:0] node843;
	wire [1-1:0] node845;
	wire [1-1:0] node848;
	wire [1-1:0] node849;
	wire [1-1:0] node855;
	wire [1-1:0] node856;
	wire [1-1:0] node857;
	wire [1-1:0] node858;
	wire [1-1:0] node859;
	wire [1-1:0] node861;
	wire [1-1:0] node862;
	wire [1-1:0] node864;
	wire [1-1:0] node866;
	wire [1-1:0] node868;
	wire [1-1:0] node871;
	wire [1-1:0] node872;
	wire [1-1:0] node874;
	wire [1-1:0] node876;
	wire [1-1:0] node879;
	wire [1-1:0] node880;
	wire [1-1:0] node881;
	wire [1-1:0] node885;
	wire [1-1:0] node886;
	wire [1-1:0] node890;
	wire [1-1:0] node891;
	wire [1-1:0] node893;
	wire [1-1:0] node895;
	wire [1-1:0] node896;
	wire [1-1:0] node897;
	wire [1-1:0] node899;
	wire [1-1:0] node903;
	wire [1-1:0] node904;
	wire [1-1:0] node906;
	wire [1-1:0] node910;
	wire [1-1:0] node911;
	wire [1-1:0] node913;
	wire [1-1:0] node916;
	wire [1-1:0] node917;
	wire [1-1:0] node919;
	wire [1-1:0] node921;
	wire [1-1:0] node924;
	wire [1-1:0] node925;
	wire [1-1:0] node926;
	wire [1-1:0] node928;
	wire [1-1:0] node931;
	wire [1-1:0] node932;
	wire [1-1:0] node937;
	wire [1-1:0] node938;
	wire [1-1:0] node939;
	wire [1-1:0] node941;
	wire [1-1:0] node943;
	wire [1-1:0] node944;
	wire [1-1:0] node946;
	wire [1-1:0] node948;
	wire [1-1:0] node952;
	wire [1-1:0] node953;
	wire [1-1:0] node955;
	wire [1-1:0] node957;
	wire [1-1:0] node958;
	wire [1-1:0] node960;
	wire [1-1:0] node964;
	wire [1-1:0] node965;
	wire [1-1:0] node966;
	wire [1-1:0] node968;
	wire [1-1:0] node971;
	wire [1-1:0] node972;
	wire [1-1:0] node974;
	wire [1-1:0] node978;
	wire [1-1:0] node979;
	wire [1-1:0] node981;
	wire [1-1:0] node982;
	wire [1-1:0] node987;
	wire [1-1:0] node988;
	wire [1-1:0] node989;
	wire [1-1:0] node991;
	wire [1-1:0] node992;
	wire [1-1:0] node994;
	wire [1-1:0] node997;
	wire [1-1:0] node998;
	wire [1-1:0] node1000;
	wire [1-1:0] node1003;
	wire [1-1:0] node1004;
	wire [1-1:0] node1008;
	wire [1-1:0] node1009;
	wire [1-1:0] node1010;
	wire [1-1:0] node1012;
	wire [1-1:0] node1015;
	wire [1-1:0] node1016;
	wire [1-1:0] node1018;
	wire [1-1:0] node1022;
	wire [1-1:0] node1023;
	wire [1-1:0] node1024;
	wire [1-1:0] node1026;
	wire [1-1:0] node1031;
	wire [1-1:0] node1032;
	wire [1-1:0] node1033;
	wire [1-1:0] node1034;
	wire [1-1:0] node1036;
	wire [1-1:0] node1039;
	wire [1-1:0] node1040;
	wire [1-1:0] node1042;
	wire [1-1:0] node1046;
	wire [1-1:0] node1047;
	wire [1-1:0] node1049;
	wire [1-1:0] node1052;
	wire [1-1:0] node1053;
	wire [1-1:0] node1054;
	wire [1-1:0] node1059;
	wire [1-1:0] node1060;
	wire [1-1:0] node1061;
	wire [1-1:0] node1062;
	wire [1-1:0] node1064;
	wire [1-1:0] node1070;
	wire [1-1:0] node1071;
	wire [1-1:0] node1072;
	wire [1-1:0] node1073;
	wire [1-1:0] node1075;
	wire [1-1:0] node1076;
	wire [1-1:0] node1078;
	wire [1-1:0] node1080;
	wire [1-1:0] node1083;
	wire [1-1:0] node1084;
	wire [1-1:0] node1086;
	wire [1-1:0] node1089;
	wire [1-1:0] node1090;
	wire [1-1:0] node1094;
	wire [1-1:0] node1095;
	wire [1-1:0] node1096;
	wire [1-1:0] node1098;
	wire [1-1:0] node1100;
	wire [1-1:0] node1103;
	wire [1-1:0] node1104;
	wire [1-1:0] node1106;
	wire [1-1:0] node1109;
	wire [1-1:0] node1112;
	wire [1-1:0] node1113;
	wire [1-1:0] node1114;
	wire [1-1:0] node1116;
	wire [1-1:0] node1118;
	wire [1-1:0] node1121;
	wire [1-1:0] node1124;
	wire [1-1:0] node1125;
	wire [1-1:0] node1126;
	wire [1-1:0] node1128;
	wire [1-1:0] node1131;
	wire [1-1:0] node1132;
	wire [1-1:0] node1137;
	wire [1-1:0] node1138;
	wire [1-1:0] node1139;
	wire [1-1:0] node1140;
	wire [1-1:0] node1142;
	wire [1-1:0] node1144;
	wire [1-1:0] node1147;
	wire [1-1:0] node1148;
	wire [1-1:0] node1150;
	wire [1-1:0] node1153;
	wire [1-1:0] node1154;
	wire [1-1:0] node1156;
	wire [1-1:0] node1160;
	wire [1-1:0] node1161;
	wire [1-1:0] node1162;
	wire [1-1:0] node1164;
	wire [1-1:0] node1167;
	wire [1-1:0] node1168;
	wire [1-1:0] node1170;
	wire [1-1:0] node1174;
	wire [1-1:0] node1175;
	wire [1-1:0] node1177;
	wire [1-1:0] node1178;
	wire [1-1:0] node1183;
	wire [1-1:0] node1184;
	wire [1-1:0] node1185;
	wire [1-1:0] node1187;
	wire [1-1:0] node1189;
	wire [1-1:0] node1190;
	wire [1-1:0] node1194;
	wire [1-1:0] node1195;
	wire [1-1:0] node1197;
	wire [1-1:0] node1198;
	wire [1-1:0] node1203;
	wire [1-1:0] node1204;
	wire [1-1:0] node1205;
	wire [1-1:0] node1207;
	wire [1-1:0] node1208;
	wire [1-1:0] node1214;
	wire [1-1:0] node1215;
	wire [1-1:0] node1216;
	wire [1-1:0] node1217;
	wire [1-1:0] node1219;
	wire [1-1:0] node1221;
	wire [1-1:0] node1222;
	wire [1-1:0] node1224;
	wire [1-1:0] node1228;
	wire [1-1:0] node1229;
	wire [1-1:0] node1230;
	wire [1-1:0] node1232;
	wire [1-1:0] node1234;
	wire [1-1:0] node1237;
	wire [1-1:0] node1240;
	wire [1-1:0] node1241;
	wire [1-1:0] node1242;
	wire [1-1:0] node1244;
	wire [1-1:0] node1247;
	wire [1-1:0] node1248;
	wire [1-1:0] node1252;
	wire [1-1:0] node1253;
	wire [1-1:0] node1257;
	wire [1-1:0] node1258;
	wire [1-1:0] node1259;
	wire [1-1:0] node1260;
	wire [1-1:0] node1262;
	wire [1-1:0] node1264;
	wire [1-1:0] node1267;
	wire [1-1:0] node1268;
	wire [1-1:0] node1270;
	wire [1-1:0] node1273;
	wire [1-1:0] node1274;
	wire [1-1:0] node1278;
	wire [1-1:0] node1279;
	wire [1-1:0] node1281;
	wire [1-1:0] node1282;
	wire [1-1:0] node1286;
	wire [1-1:0] node1287;
	wire [1-1:0] node1289;
	wire [1-1:0] node1293;
	wire [1-1:0] node1294;
	wire [1-1:0] node1295;
	wire [1-1:0] node1296;
	wire [1-1:0] node1298;
	wire [1-1:0] node1301;
	wire [1-1:0] node1302;
	wire [1-1:0] node1308;
	wire [1-1:0] node1309;
	wire [1-1:0] node1310;
	wire [1-1:0] node1311;
	wire [1-1:0] node1313;
	wire [1-1:0] node1315;
	wire [1-1:0] node1316;
	wire [1-1:0] node1320;
	wire [1-1:0] node1321;
	wire [1-1:0] node1322;
	wire [1-1:0] node1324;
	wire [1-1:0] node1329;
	wire [1-1:0] node1330;
	wire [1-1:0] node1331;
	wire [1-1:0] node1333;
	wire [1-1:0] node1336;
	wire [1-1:0] node1337;
	wire [1-1:0] node1338;
	wire [1-1:0] node1344;
	wire [1-1:0] node1345;
	wire [1-1:0] node1346;
	wire [1-1:0] node1347;
	wire [1-1:0] node1349;
	wire [1-1:0] node1350;
	wire [1-1:0] node1355;
	wire [1-1:0] node1356;
	wire [1-1:0] node1357;
	wire [1-1:0] node1363;
	wire [1-1:0] node1364;
	wire [1-1:0] node1365;
	wire [1-1:0] node1366;
	wire [1-1:0] node1367;
	wire [1-1:0] node1369;
	wire [1-1:0] node1371;
	wire [1-1:0] node1373;
	wire [1-1:0] node1374;
	wire [1-1:0] node1378;
	wire [1-1:0] node1379;
	wire [1-1:0] node1381;
	wire [1-1:0] node1383;
	wire [1-1:0] node1386;
	wire [1-1:0] node1387;
	wire [1-1:0] node1389;
	wire [1-1:0] node1392;
	wire [1-1:0] node1393;
	wire [1-1:0] node1395;
	wire [1-1:0] node1399;
	wire [1-1:0] node1400;
	wire [1-1:0] node1401;
	wire [1-1:0] node1403;
	wire [1-1:0] node1404;
	wire [1-1:0] node1406;
	wire [1-1:0] node1408;
	wire [1-1:0] node1411;
	wire [1-1:0] node1412;
	wire [1-1:0] node1416;
	wire [1-1:0] node1417;
	wire [1-1:0] node1419;
	wire [1-1:0] node1420;
	wire [1-1:0] node1422;
	wire [1-1:0] node1426;
	wire [1-1:0] node1427;
	wire [1-1:0] node1428;
	wire [1-1:0] node1433;
	wire [1-1:0] node1434;
	wire [1-1:0] node1435;
	wire [1-1:0] node1436;
	wire [1-1:0] node1438;
	wire [1-1:0] node1440;
	wire [1-1:0] node1443;
	wire [1-1:0] node1444;
	wire [1-1:0] node1446;
	wire [1-1:0] node1449;
	wire [1-1:0] node1452;
	wire [1-1:0] node1453;
	wire [1-1:0] node1456;
	wire [1-1:0] node1457;
	wire [1-1:0] node1458;
	wire [1-1:0] node1463;
	wire [1-1:0] node1464;
	wire [1-1:0] node1465;
	wire [1-1:0] node1466;
	wire [1-1:0] node1468;
	wire [1-1:0] node1471;
	wire [1-1:0] node1474;
	wire [1-1:0] node1475;
	wire [1-1:0] node1476;
	wire [1-1:0] node1482;
	wire [1-1:0] node1483;
	wire [1-1:0] node1484;
	wire [1-1:0] node1485;
	wire [1-1:0] node1487;
	wire [1-1:0] node1489;
	wire [1-1:0] node1490;
	wire [1-1:0] node1492;
	wire [1-1:0] node1496;
	wire [1-1:0] node1497;
	wire [1-1:0] node1498;
	wire [1-1:0] node1500;
	wire [1-1:0] node1503;
	wire [1-1:0] node1505;
	wire [1-1:0] node1506;
	wire [1-1:0] node1510;
	wire [1-1:0] node1511;
	wire [1-1:0] node1512;
	wire [1-1:0] node1514;
	wire [1-1:0] node1519;
	wire [1-1:0] node1520;
	wire [1-1:0] node1521;
	wire [1-1:0] node1523;
	wire [1-1:0] node1524;
	wire [1-1:0] node1526;
	wire [1-1:0] node1530;
	wire [1-1:0] node1531;
	wire [1-1:0] node1532;
	wire [1-1:0] node1535;
	wire [1-1:0] node1536;
	wire [1-1:0] node1541;
	wire [1-1:0] node1542;
	wire [1-1:0] node1543;
	wire [1-1:0] node1545;
	wire [1-1:0] node1549;
	wire [1-1:0] node1550;
	wire [1-1:0] node1551;
	wire [1-1:0] node1556;
	wire [1-1:0] node1557;
	wire [1-1:0] node1558;
	wire [1-1:0] node1559;
	wire [1-1:0] node1561;
	wire [1-1:0] node1563;
	wire [1-1:0] node1566;
	wire [1-1:0] node1567;
	wire [1-1:0] node1571;
	wire [1-1:0] node1572;
	wire [1-1:0] node1573;
	wire [1-1:0] node1574;
	wire [1-1:0] node1576;
	wire [1-1:0] node1580;
	wire [1-1:0] node1581;
	wire [1-1:0] node1586;
	wire [1-1:0] node1587;
	wire [1-1:0] node1588;
	wire [1-1:0] node1589;
	wire [1-1:0] node1590;
	wire [1-1:0] node1592;
	wire [1-1:0] node1595;
	wire [1-1:0] node1596;
	wire [1-1:0] node1600;
	wire [1-1:0] node1601;
	wire [1-1:0] node1602;
	wire [1-1:0] node1607;
	wire [1-1:0] node1608;
	wire [1-1:0] node1609;
	wire [1-1:0] node1610;
	wire [1-1:0] node1617;
	wire [1-1:0] node1618;
	wire [1-1:0] node1619;
	wire [1-1:0] node1620;
	wire [1-1:0] node1621;
	wire [1-1:0] node1623;
	wire [1-1:0] node1625;
	wire [1-1:0] node1626;
	wire [1-1:0] node1628;
	wire [1-1:0] node1632;
	wire [1-1:0] node1633;
	wire [1-1:0] node1635;
	wire [1-1:0] node1636;
	wire [1-1:0] node1638;
	wire [1-1:0] node1641;
	wire [1-1:0] node1642;
	wire [1-1:0] node1646;
	wire [1-1:0] node1647;
	wire [1-1:0] node1648;
	wire [1-1:0] node1652;
	wire [1-1:0] node1653;
	wire [1-1:0] node1654;
	wire [1-1:0] node1659;
	wire [1-1:0] node1660;
	wire [1-1:0] node1661;
	wire [1-1:0] node1663;
	wire [1-1:0] node1665;
	wire [1-1:0] node1666;
	wire [1-1:0] node1670;
	wire [1-1:0] node1671;
	wire [1-1:0] node1675;
	wire [1-1:0] node1676;
	wire [1-1:0] node1677;
	wire [1-1:0] node1678;
	wire [1-1:0] node1680;
	wire [1-1:0] node1683;
	wire [1-1:0] node1684;
	wire [1-1:0] node1690;
	wire [1-1:0] node1691;
	wire [1-1:0] node1692;
	wire [1-1:0] node1693;
	wire [1-1:0] node1694;
	wire [1-1:0] node1696;
	wire [1-1:0] node1698;
	wire [1-1:0] node1701;
	wire [1-1:0] node1702;
	wire [1-1:0] node1704;
	wire [1-1:0] node1708;
	wire [1-1:0] node1709;
	wire [1-1:0] node1711;
	wire [1-1:0] node1712;
	wire [1-1:0] node1717;
	wire [1-1:0] node1718;
	wire [1-1:0] node1719;
	wire [1-1:0] node1720;
	wire [1-1:0] node1723;
	wire [1-1:0] node1726;
	wire [1-1:0] node1727;
	wire [1-1:0] node1731;
	wire [1-1:0] node1732;
	wire [1-1:0] node1733;
	wire [1-1:0] node1738;
	wire [1-1:0] node1739;
	wire [1-1:0] node1740;
	wire [1-1:0] node1741;
	wire [1-1:0] node1743;
	wire [1-1:0] node1745;
	wire [1-1:0] node1751;
	wire [1-1:0] node1752;
	wire [1-1:0] node1753;
	wire [1-1:0] node1754;
	wire [1-1:0] node1755;
	wire [1-1:0] node1757;
	wire [1-1:0] node1758;
	wire [1-1:0] node1762;
	wire [1-1:0] node1763;
	wire [1-1:0] node1765;
	wire [1-1:0] node1769;
	wire [1-1:0] node1770;
	wire [1-1:0] node1771;
	wire [1-1:0] node1772;
	wire [1-1:0] node1774;
	wire [1-1:0] node1777;
	wire [1-1:0] node1778;
	wire [1-1:0] node1784;
	wire [1-1:0] node1785;
	wire [1-1:0] node1786;
	wire [1-1:0] node1787;
	wire [1-1:0] node1789;
	wire [1-1:0] node1792;
	wire [1-1:0] node1793;
	wire [1-1:0] node1797;
	wire [1-1:0] node1798;
	wire [1-1:0] node1799;
	wire [1-1:0] node1805;
	wire [1-1:0] node1806;
	wire [1-1:0] node1807;
	wire [1-1:0] node1808;
	wire [1-1:0] node1809;
	wire [1-1:0] node1811;
	wire [1-1:0] node1814;
	wire [1-1:0] node1815;
	wire [1-1:0] node1822;
	wire [1-1:0] node1823;
	wire [1-1:0] node1824;
	wire [1-1:0] node1825;
	wire [1-1:0] node1826;
	wire [1-1:0] node1827;
	wire [1-1:0] node1829;
	wire [1-1:0] node1830;
	wire [1-1:0] node1832;
	wire [1-1:0] node1834;
	wire [1-1:0] node1836;
	wire [1-1:0] node1839;
	wire [1-1:0] node1841;
	wire [1-1:0] node1843;
	wire [1-1:0] node1844;
	wire [1-1:0] node1846;
	wire [1-1:0] node1850;
	wire [1-1:0] node1851;
	wire [1-1:0] node1853;
	wire [1-1:0] node1855;
	wire [1-1:0] node1857;
	wire [1-1:0] node1858;
	wire [1-1:0] node1860;
	wire [1-1:0] node1863;
	wire [1-1:0] node1864;
	wire [1-1:0] node1868;
	wire [1-1:0] node1869;
	wire [1-1:0] node1871;
	wire [1-1:0] node1872;
	wire [1-1:0] node1873;
	wire [1-1:0] node1875;
	wire [1-1:0] node1879;
	wire [1-1:0] node1880;
	wire [1-1:0] node1882;
	wire [1-1:0] node1885;
	wire [1-1:0] node1886;
	wire [1-1:0] node1890;
	wire [1-1:0] node1891;
	wire [1-1:0] node1893;
	wire [1-1:0] node1894;
	wire [1-1:0] node1898;
	wire [1-1:0] node1899;
	wire [1-1:0] node1900;
	wire [1-1:0] node1903;
	wire [1-1:0] node1904;
	wire [1-1:0] node1909;
	wire [1-1:0] node1910;
	wire [1-1:0] node1911;
	wire [1-1:0] node1913;
	wire [1-1:0] node1914;
	wire [1-1:0] node1916;
	wire [1-1:0] node1918;
	wire [1-1:0] node1921;
	wire [1-1:0] node1922;
	wire [1-1:0] node1924;
	wire [1-1:0] node1926;
	wire [1-1:0] node1929;
	wire [1-1:0] node1932;
	wire [1-1:0] node1933;
	wire [1-1:0] node1935;
	wire [1-1:0] node1937;
	wire [1-1:0] node1939;
	wire [1-1:0] node1942;
	wire [1-1:0] node1943;
	wire [1-1:0] node1944;
	wire [1-1:0] node1946;
	wire [1-1:0] node1948;
	wire [1-1:0] node1951;
	wire [1-1:0] node1952;
	wire [1-1:0] node1954;
	wire [1-1:0] node1957;
	wire [1-1:0] node1960;
	wire [1-1:0] node1961;
	wire [1-1:0] node1962;
	wire [1-1:0] node1964;
	wire [1-1:0] node1969;
	wire [1-1:0] node1970;
	wire [1-1:0] node1971;
	wire [1-1:0] node1973;
	wire [1-1:0] node1975;
	wire [1-1:0] node1977;
	wire [1-1:0] node1978;
	wire [1-1:0] node1982;
	wire [1-1:0] node1983;
	wire [1-1:0] node1985;
	wire [1-1:0] node1986;
	wire [1-1:0] node1988;
	wire [1-1:0] node1992;
	wire [1-1:0] node1993;
	wire [1-1:0] node1994;
	wire [1-1:0] node1997;
	wire [1-1:0] node1998;
	wire [1-1:0] node2003;
	wire [1-1:0] node2004;
	wire [1-1:0] node2005;
	wire [1-1:0] node2006;
	wire [1-1:0] node2008;
	wire [1-1:0] node2011;
	wire [1-1:0] node2012;
	wire [1-1:0] node2014;
	wire [1-1:0] node2017;
	wire [1-1:0] node2020;
	wire [1-1:0] node2021;
	wire [1-1:0] node2022;
	wire [1-1:0] node2027;
	wire [1-1:0] node2028;
	wire [1-1:0] node2029;
	wire [1-1:0] node2030;
	wire [1-1:0] node2032;
	wire [1-1:0] node2035;
	wire [1-1:0] node2040;
	wire [1-1:0] node2041;
	wire [1-1:0] node2042;
	wire [1-1:0] node2043;
	wire [1-1:0] node2044;
	wire [1-1:0] node2045;
	wire [1-1:0] node2047;
	wire [1-1:0] node2051;
	wire [1-1:0] node2052;
	wire [1-1:0] node2054;
	wire [1-1:0] node2056;
	wire [1-1:0] node2059;
	wire [1-1:0] node2061;
	wire [1-1:0] node2062;
	wire [1-1:0] node2064;
	wire [1-1:0] node2067;
	wire [1-1:0] node2068;
	wire [1-1:0] node2072;
	wire [1-1:0] node2073;
	wire [1-1:0] node2074;
	wire [1-1:0] node2076;
	wire [1-1:0] node2078;
	wire [1-1:0] node2080;
	wire [1-1:0] node2083;
	wire [1-1:0] node2084;
	wire [1-1:0] node2086;
	wire [1-1:0] node2089;
	wire [1-1:0] node2090;
	wire [1-1:0] node2094;
	wire [1-1:0] node2095;
	wire [1-1:0] node2097;
	wire [1-1:0] node2098;
	wire [1-1:0] node2100;
	wire [1-1:0] node2104;
	wire [1-1:0] node2105;
	wire [1-1:0] node2107;
	wire [1-1:0] node2109;
	wire [1-1:0] node2113;
	wire [1-1:0] node2114;
	wire [1-1:0] node2115;
	wire [1-1:0] node2117;
	wire [1-1:0] node2118;
	wire [1-1:0] node2120;
	wire [1-1:0] node2122;
	wire [1-1:0] node2125;
	wire [1-1:0] node2126;
	wire [1-1:0] node2130;
	wire [1-1:0] node2131;
	wire [1-1:0] node2133;
	wire [1-1:0] node2135;
	wire [1-1:0] node2136;
	wire [1-1:0] node2140;
	wire [1-1:0] node2141;
	wire [1-1:0] node2143;
	wire [1-1:0] node2144;
	wire [1-1:0] node2148;
	wire [1-1:0] node2150;
	wire [1-1:0] node2151;
	wire [1-1:0] node2155;
	wire [1-1:0] node2156;
	wire [1-1:0] node2157;
	wire [1-1:0] node2159;
	wire [1-1:0] node2162;
	wire [1-1:0] node2163;
	wire [1-1:0] node2165;
	wire [1-1:0] node2166;
	wire [1-1:0] node2171;
	wire [1-1:0] node2172;
	wire [1-1:0] node2173;
	wire [1-1:0] node2175;
	wire [1-1:0] node2176;
	wire [1-1:0] node2180;
	wire [1-1:0] node2181;
	wire [1-1:0] node2185;
	wire [1-1:0] node2186;
	wire [1-1:0] node2187;
	wire [1-1:0] node2192;
	wire [1-1:0] node2193;
	wire [1-1:0] node2194;
	wire [1-1:0] node2195;
	wire [1-1:0] node2197;
	wire [1-1:0] node2199;
	wire [1-1:0] node2201;
	wire [1-1:0] node2202;
	wire [1-1:0] node2206;
	wire [1-1:0] node2207;
	wire [1-1:0] node2208;
	wire [1-1:0] node2210;
	wire [1-1:0] node2211;
	wire [1-1:0] node2215;
	wire [1-1:0] node2216;
	wire [1-1:0] node2218;
	wire [1-1:0] node2222;
	wire [1-1:0] node2223;
	wire [1-1:0] node2224;
	wire [1-1:0] node2229;
	wire [1-1:0] node2230;
	wire [1-1:0] node2231;
	wire [1-1:0] node2232;
	wire [1-1:0] node2234;
	wire [1-1:0] node2236;
	wire [1-1:0] node2239;
	wire [1-1:0] node2240;
	wire [1-1:0] node2242;
	wire [1-1:0] node2246;
	wire [1-1:0] node2247;
	wire [1-1:0] node2251;
	wire [1-1:0] node2252;
	wire [1-1:0] node2253;
	wire [1-1:0] node2255;
	wire [1-1:0] node2260;
	wire [1-1:0] node2261;
	wire [1-1:0] node2262;
	wire [1-1:0] node2263;
	wire [1-1:0] node2265;
	wire [1-1:0] node2267;
	wire [1-1:0] node2269;
	wire [1-1:0] node2272;
	wire [1-1:0] node2273;
	wire [1-1:0] node2275;
	wire [1-1:0] node2279;
	wire [1-1:0] node2280;
	wire [1-1:0] node2281;
	wire [1-1:0] node2283;
	wire [1-1:0] node2286;
	wire [1-1:0] node2287;
	wire [1-1:0] node2288;
	wire [1-1:0] node2294;
	wire [1-1:0] node2295;
	wire [1-1:0] node2296;
	wire [1-1:0] node2297;
	wire [1-1:0] node2298;
	wire [1-1:0] node2300;
	wire [1-1:0] node2305;
	wire [1-1:0] node2306;
	wire [1-1:0] node2308;
	wire [1-1:0] node2313;
	wire [1-1:0] node2314;
	wire [1-1:0] node2315;
	wire [1-1:0] node2316;
	wire [1-1:0] node2317;
	wire [1-1:0] node2319;
	wire [1-1:0] node2320;
	wire [1-1:0] node2322;
	wire [1-1:0] node2324;
	wire [1-1:0] node2326;
	wire [1-1:0] node2329;
	wire [1-1:0] node2330;
	wire [1-1:0] node2332;
	wire [1-1:0] node2335;
	wire [1-1:0] node2337;
	wire [1-1:0] node2338;
	wire [1-1:0] node2342;
	wire [1-1:0] node2343;
	wire [1-1:0] node2345;
	wire [1-1:0] node2346;
	wire [1-1:0] node2348;
	wire [1-1:0] node2350;
	wire [1-1:0] node2353;
	wire [1-1:0] node2354;
	wire [1-1:0] node2356;
	wire [1-1:0] node2360;
	wire [1-1:0] node2361;
	wire [1-1:0] node2363;
	wire [1-1:0] node2364;
	wire [1-1:0] node2366;
	wire [1-1:0] node2369;
	wire [1-1:0] node2370;
	wire [1-1:0] node2374;
	wire [1-1:0] node2375;
	wire [1-1:0] node2379;
	wire [1-1:0] node2380;
	wire [1-1:0] node2381;
	wire [1-1:0] node2383;
	wire [1-1:0] node2385;
	wire [1-1:0] node2388;
	wire [1-1:0] node2389;
	wire [1-1:0] node2391;
	wire [1-1:0] node2392;
	wire [1-1:0] node2396;
	wire [1-1:0] node2397;
	wire [1-1:0] node2398;
	wire [1-1:0] node2400;
	wire [1-1:0] node2405;
	wire [1-1:0] node2406;
	wire [1-1:0] node2407;
	wire [1-1:0] node2408;
	wire [1-1:0] node2411;
	wire [1-1:0] node2412;
	wire [1-1:0] node2414;
	wire [1-1:0] node2418;
	wire [1-1:0] node2419;
	wire [1-1:0] node2421;
	wire [1-1:0] node2422;
	wire [1-1:0] node2426;
	wire [1-1:0] node2428;
	wire [1-1:0] node2429;
	wire [1-1:0] node2433;
	wire [1-1:0] node2434;
	wire [1-1:0] node2435;
	wire [1-1:0] node2437;
	wire [1-1:0] node2438;
	wire [1-1:0] node2444;
	wire [1-1:0] node2445;
	wire [1-1:0] node2446;
	wire [1-1:0] node2447;
	wire [1-1:0] node2448;
	wire [1-1:0] node2450;
	wire [1-1:0] node2452;
	wire [1-1:0] node2454;
	wire [1-1:0] node2457;
	wire [1-1:0] node2458;
	wire [1-1:0] node2460;
	wire [1-1:0] node2462;
	wire [1-1:0] node2465;
	wire [1-1:0] node2466;
	wire [1-1:0] node2469;
	wire [1-1:0] node2472;
	wire [1-1:0] node2473;
	wire [1-1:0] node2475;
	wire [1-1:0] node2477;
	wire [1-1:0] node2478;
	wire [1-1:0] node2482;
	wire [1-1:0] node2483;
	wire [1-1:0] node2484;
	wire [1-1:0] node2489;
	wire [1-1:0] node2490;
	wire [1-1:0] node2491;
	wire [1-1:0] node2493;
	wire [1-1:0] node2495;
	wire [1-1:0] node2498;
	wire [1-1:0] node2499;
	wire [1-1:0] node2501;
	wire [1-1:0] node2502;
	wire [1-1:0] node2506;
	wire [1-1:0] node2507;
	wire [1-1:0] node2511;
	wire [1-1:0] node2512;
	wire [1-1:0] node2513;
	wire [1-1:0] node2515;
	wire [1-1:0] node2518;
	wire [1-1:0] node2519;
	wire [1-1:0] node2524;
	wire [1-1:0] node2525;
	wire [1-1:0] node2526;
	wire [1-1:0] node2527;
	wire [1-1:0] node2529;
	wire [1-1:0] node2530;
	wire [1-1:0] node2532;
	wire [1-1:0] node2536;
	wire [1-1:0] node2537;
	wire [1-1:0] node2541;
	wire [1-1:0] node2542;
	wire [1-1:0] node2543;
	wire [1-1:0] node2544;
	wire [1-1:0] node2546;
	wire [1-1:0] node2549;
	wire [1-1:0] node2551;
	wire [1-1:0] node2554;
	wire [1-1:0] node2556;
	wire [1-1:0] node2560;
	wire [1-1:0] node2561;
	wire [1-1:0] node2562;
	wire [1-1:0] node2563;
	wire [1-1:0] node2564;
	wire [1-1:0] node2566;
	wire [1-1:0] node2570;
	wire [1-1:0] node2571;
	wire [1-1:0] node2572;
	wire [1-1:0] node2579;
	wire [1-1:0] node2580;
	wire [1-1:0] node2581;
	wire [1-1:0] node2582;
	wire [1-1:0] node2583;
	wire [1-1:0] node2585;
	wire [1-1:0] node2587;
	wire [1-1:0] node2588;
	wire [1-1:0] node2590;
	wire [1-1:0] node2594;
	wire [1-1:0] node2595;
	wire [1-1:0] node2596;
	wire [1-1:0] node2598;
	wire [1-1:0] node2600;
	wire [1-1:0] node2603;
	wire [1-1:0] node2604;
	wire [1-1:0] node2606;
	wire [1-1:0] node2610;
	wire [1-1:0] node2611;
	wire [1-1:0] node2612;
	wire [1-1:0] node2614;
	wire [1-1:0] node2617;
	wire [1-1:0] node2618;
	wire [1-1:0] node2623;
	wire [1-1:0] node2624;
	wire [1-1:0] node2625;
	wire [1-1:0] node2627;
	wire [1-1:0] node2630;
	wire [1-1:0] node2631;
	wire [1-1:0] node2633;
	wire [1-1:0] node2634;
	wire [1-1:0] node2639;
	wire [1-1:0] node2640;
	wire [1-1:0] node2641;
	wire [1-1:0] node2643;
	wire [1-1:0] node2644;
	wire [1-1:0] node2650;
	wire [1-1:0] node2651;
	wire [1-1:0] node2652;
	wire [1-1:0] node2653;
	wire [1-1:0] node2655;
	wire [1-1:0] node2658;
	wire [1-1:0] node2659;
	wire [1-1:0] node2660;
	wire [1-1:0] node2662;
	wire [1-1:0] node2665;
	wire [1-1:0] node2666;
	wire [1-1:0] node2671;
	wire [1-1:0] node2672;
	wire [1-1:0] node2673;
	wire [1-1:0] node2674;
	wire [1-1:0] node2676;
	wire [1-1:0] node2682;
	wire [1-1:0] node2683;
	wire [1-1:0] node2684;
	wire [1-1:0] node2685;
	wire [1-1:0] node2686;
	wire [1-1:0] node2688;
	wire [1-1:0] node2692;
	wire [1-1:0] node2693;
	wire [1-1:0] node2694;
	wire [1-1:0] node2699;
	wire [1-1:0] node2700;
	wire [1-1:0] node2701;
	wire [1-1:0] node2702;
	wire [1-1:0] node2709;
	wire [1-1:0] node2710;
	wire [1-1:0] node2711;
	wire [1-1:0] node2712;
	wire [1-1:0] node2713;
	wire [1-1:0] node2715;
	wire [1-1:0] node2718;
	wire [1-1:0] node2719;
	wire [1-1:0] node2721;
	wire [1-1:0] node2725;
	wire [1-1:0] node2726;
	wire [1-1:0] node2727;
	wire [1-1:0] node2729;
	wire [1-1:0] node2734;
	wire [1-1:0] node2735;
	wire [1-1:0] node2736;
	wire [1-1:0] node2737;
	wire [1-1:0] node2740;
	wire [1-1:0] node2741;
	wire [1-1:0] node2747;
	wire [1-1:0] node2748;
	wire [1-1:0] node2749;
	wire [1-1:0] node2750;
	wire [1-1:0] node2751;
	wire [1-1:0] node2755;
	wire [1-1:0] node2756;
	wire [1-1:0] node2757;
	wire [1-1:0] node2758;
	wire [1-1:0] node2766;
	wire [1-1:0] node2767;
	wire [1-1:0] node2768;
	wire [1-1:0] node2769;
	wire [1-1:0] node2770;
	wire [1-1:0] node2771;
	wire [1-1:0] node2773;
	wire [1-1:0] node2775;
	wire [1-1:0] node2777;
	wire [1-1:0] node2778;
	wire [1-1:0] node2780;
	wire [1-1:0] node2784;
	wire [1-1:0] node2785;
	wire [1-1:0] node2787;
	wire [1-1:0] node2788;
	wire [1-1:0] node2790;
	wire [1-1:0] node2793;
	wire [1-1:0] node2796;
	wire [1-1:0] node2797;
	wire [1-1:0] node2798;
	wire [1-1:0] node2800;
	wire [1-1:0] node2802;
	wire [1-1:0] node2805;
	wire [1-1:0] node2808;
	wire [1-1:0] node2809;
	wire [1-1:0] node2811;
	wire [1-1:0] node2814;
	wire [1-1:0] node2815;
	wire [1-1:0] node2816;
	wire [1-1:0] node2821;
	wire [1-1:0] node2822;
	wire [1-1:0] node2823;
	wire [1-1:0] node2825;
	wire [1-1:0] node2827;
	wire [1-1:0] node2829;
	wire [1-1:0] node2832;
	wire [1-1:0] node2833;
	wire [1-1:0] node2835;
	wire [1-1:0] node2836;
	wire [1-1:0] node2838;
	wire [1-1:0] node2842;
	wire [1-1:0] node2843;
	wire [1-1:0] node2847;
	wire [1-1:0] node2848;
	wire [1-1:0] node2849;
	wire [1-1:0] node2850;
	wire [1-1:0] node2852;
	wire [1-1:0] node2854;
	wire [1-1:0] node2857;
	wire [1-1:0] node2858;
	wire [1-1:0] node2860;
	wire [1-1:0] node2864;
	wire [1-1:0] node2865;
	wire [1-1:0] node2867;
	wire [1-1:0] node2869;
	wire [1-1:0] node2873;
	wire [1-1:0] node2874;
	wire [1-1:0] node2875;
	wire [1-1:0] node2877;
	wire [1-1:0] node2878;
	wire [1-1:0] node2882;
	wire [1-1:0] node2883;
	wire [1-1:0] node2884;
	wire [1-1:0] node2890;
	wire [1-1:0] node2891;
	wire [1-1:0] node2892;
	wire [1-1:0] node2893;
	wire [1-1:0] node2895;
	wire [1-1:0] node2896;
	wire [1-1:0] node2898;
	wire [1-1:0] node2901;
	wire [1-1:0] node2902;
	wire [1-1:0] node2904;
	wire [1-1:0] node2908;
	wire [1-1:0] node2909;
	wire [1-1:0] node2911;
	wire [1-1:0] node2912;
	wire [1-1:0] node2914;
	wire [1-1:0] node2917;
	wire [1-1:0] node2920;
	wire [1-1:0] node2921;
	wire [1-1:0] node2922;
	wire [1-1:0] node2924;
	wire [1-1:0] node2929;
	wire [1-1:0] node2930;
	wire [1-1:0] node2931;
	wire [1-1:0] node2933;
	wire [1-1:0] node2934;
	wire [1-1:0] node2936;
	wire [1-1:0] node2940;
	wire [1-1:0] node2941;
	wire [1-1:0] node2943;
	wire [1-1:0] node2944;
	wire [1-1:0] node2949;
	wire [1-1:0] node2950;
	wire [1-1:0] node2951;
	wire [1-1:0] node2953;
	wire [1-1:0] node2954;
	wire [1-1:0] node2958;
	wire [1-1:0] node2959;
	wire [1-1:0] node2964;
	wire [1-1:0] node2965;
	wire [1-1:0] node2966;
	wire [1-1:0] node2967;
	wire [1-1:0] node2969;
	wire [1-1:0] node2971;
	wire [1-1:0] node2972;
	wire [1-1:0] node2976;
	wire [1-1:0] node2977;
	wire [1-1:0] node2979;
	wire [1-1:0] node2980;
	wire [1-1:0] node2984;
	wire [1-1:0] node2985;
	wire [1-1:0] node2986;
	wire [1-1:0] node2991;
	wire [1-1:0] node2992;
	wire [1-1:0] node2993;
	wire [1-1:0] node2995;
	wire [1-1:0] node2996;
	wire [1-1:0] node3002;
	wire [1-1:0] node3003;
	wire [1-1:0] node3004;
	wire [1-1:0] node3005;
	wire [1-1:0] node3006;
	wire [1-1:0] node3008;
	wire [1-1:0] node3015;
	wire [1-1:0] node3016;
	wire [1-1:0] node3017;
	wire [1-1:0] node3018;
	wire [1-1:0] node3019;
	wire [1-1:0] node3021;
	wire [1-1:0] node3023;
	wire [1-1:0] node3024;
	wire [1-1:0] node3028;
	wire [1-1:0] node3029;
	wire [1-1:0] node3031;
	wire [1-1:0] node3033;
	wire [1-1:0] node3034;
	wire [1-1:0] node3038;
	wire [1-1:0] node3039;
	wire [1-1:0] node3043;
	wire [1-1:0] node3044;
	wire [1-1:0] node3045;
	wire [1-1:0] node3047;
	wire [1-1:0] node3050;
	wire [1-1:0] node3051;
	wire [1-1:0] node3052;
	wire [1-1:0] node3054;
	wire [1-1:0] node3057;
	wire [1-1:0] node3058;
	wire [1-1:0] node3063;
	wire [1-1:0] node3064;
	wire [1-1:0] node3065;
	wire [1-1:0] node3066;
	wire [1-1:0] node3068;
	wire [1-1:0] node3074;
	wire [1-1:0] node3075;
	wire [1-1:0] node3076;
	wire [1-1:0] node3077;
	wire [1-1:0] node3079;
	wire [1-1:0] node3082;
	wire [1-1:0] node3083;
	wire [1-1:0] node3087;
	wire [1-1:0] node3088;
	wire [1-1:0] node3089;
	wire [1-1:0] node3091;
	wire [1-1:0] node3092;
	wire [1-1:0] node3096;
	wire [1-1:0] node3097;
	wire [1-1:0] node3102;
	wire [1-1:0] node3103;
	wire [1-1:0] node3104;
	wire [1-1:0] node3105;
	wire [1-1:0] node3107;
	wire [1-1:0] node3108;
	wire [1-1:0] node3113;
	wire [1-1:0] node3114;
	wire [1-1:0] node3115;
	wire [1-1:0] node3121;
	wire [1-1:0] node3122;
	wire [1-1:0] node3123;
	wire [1-1:0] node3124;
	wire [1-1:0] node3125;
	wire [1-1:0] node3127;
	wire [1-1:0] node3128;
	wire [1-1:0] node3130;
	wire [1-1:0] node3133;
	wire [1-1:0] node3134;
	wire [1-1:0] node3138;
	wire [1-1:0] node3141;
	wire [1-1:0] node3142;
	wire [1-1:0] node3143;
	wire [1-1:0] node3144;
	wire [1-1:0] node3146;
	wire [1-1:0] node3149;
	wire [1-1:0] node3150;
	wire [1-1:0] node3154;
	wire [1-1:0] node3156;
	wire [1-1:0] node3157;
	wire [1-1:0] node3162;
	wire [1-1:0] node3163;
	wire [1-1:0] node3164;
	wire [1-1:0] node3165;
	wire [1-1:0] node3167;
	wire [1-1:0] node3168;
	wire [1-1:0] node3172;
	wire [1-1:0] node3173;
	wire [1-1:0] node3174;
	wire [1-1:0] node3181;
	wire [1-1:0] node3182;
	wire [1-1:0] node3183;
	wire [1-1:0] node3184;
	wire [1-1:0] node3185;
	wire [1-1:0] node3187;
	wire [1-1:0] node3189;
	wire [1-1:0] node3192;
	wire [1-1:0] node3193;
	wire [1-1:0] node3197;
	wire [1-1:0] node3198;
	wire [1-1:0] node3199;
	wire [1-1:0] node3206;
	wire [1-1:0] node3207;
	wire [1-1:0] node3208;
	wire [1-1:0] node3209;
	wire [1-1:0] node3210;
	wire [1-1:0] node3211;
	wire [1-1:0] node3213;
	wire [1-1:0] node3214;
	wire [1-1:0] node3216;
	wire [1-1:0] node3218;
	wire [1-1:0] node3221;
	wire [1-1:0] node3222;
	wire [1-1:0] node3224;
	wire [1-1:0] node3228;
	wire [1-1:0] node3229;
	wire [1-1:0] node3230;
	wire [1-1:0] node3232;
	wire [1-1:0] node3235;
	wire [1-1:0] node3236;
	wire [1-1:0] node3240;
	wire [1-1:0] node3241;
	wire [1-1:0] node3242;
	wire [1-1:0] node3243;
	wire [1-1:0] node3247;
	wire [1-1:0] node3248;
	wire [1-1:0] node3253;
	wire [1-1:0] node3254;
	wire [1-1:0] node3255;
	wire [1-1:0] node3257;
	wire [1-1:0] node3258;
	wire [1-1:0] node3260;
	wire [1-1:0] node3264;
	wire [1-1:0] node3265;
	wire [1-1:0] node3267;
	wire [1-1:0] node3268;
	wire [1-1:0] node3272;
	wire [1-1:0] node3273;
	wire [1-1:0] node3274;
	wire [1-1:0] node3279;
	wire [1-1:0] node3280;
	wire [1-1:0] node3281;
	wire [1-1:0] node3282;
	wire [1-1:0] node3284;
	wire [1-1:0] node3287;
	wire [1-1:0] node3288;
	wire [1-1:0] node3294;
	wire [1-1:0] node3295;
	wire [1-1:0] node3296;
	wire [1-1:0] node3297;
	wire [1-1:0] node3298;
	wire [1-1:0] node3300;
	wire [1-1:0] node3302;
	wire [1-1:0] node3305;
	wire [1-1:0] node3306;
	wire [1-1:0] node3308;
	wire [1-1:0] node3312;
	wire [1-1:0] node3313;
	wire [1-1:0] node3314;
	wire [1-1:0] node3316;
	wire [1-1:0] node3319;
	wire [1-1:0] node3320;
	wire [1-1:0] node3324;
	wire [1-1:0] node3325;
	wire [1-1:0] node3329;
	wire [1-1:0] node3330;
	wire [1-1:0] node3331;
	wire [1-1:0] node3333;
	wire [1-1:0] node3334;
	wire [1-1:0] node3340;
	wire [1-1:0] node3341;
	wire [1-1:0] node3342;
	wire [1-1:0] node3343;
	wire [1-1:0] node3345;
	wire [1-1:0] node3348;
	wire [1-1:0] node3349;
	wire [1-1:0] node3350;
	wire [1-1:0] node3357;
	wire [1-1:0] node3358;
	wire [1-1:0] node3359;
	wire [1-1:0] node3360;
	wire [1-1:0] node3361;
	wire [1-1:0] node3363;
	wire [1-1:0] node3364;
	wire [1-1:0] node3368;
	wire [1-1:0] node3369;
	wire [1-1:0] node3371;
	wire [1-1:0] node3372;
	wire [1-1:0] node3376;
	wire [1-1:0] node3377;
	wire [1-1:0] node3378;
	wire [1-1:0] node3383;
	wire [1-1:0] node3384;
	wire [1-1:0] node3385;
	wire [1-1:0] node3387;
	wire [1-1:0] node3388;
	wire [1-1:0] node3392;
	wire [1-1:0] node3393;
	wire [1-1:0] node3394;
	wire [1-1:0] node3400;
	wire [1-1:0] node3401;
	wire [1-1:0] node3402;
	wire [1-1:0] node3404;
	wire [1-1:0] node3405;
	wire [1-1:0] node3409;
	wire [1-1:0] node3410;
	wire [1-1:0] node3411;
	wire [1-1:0] node3412;
	wire [1-1:0] node3419;
	wire [1-1:0] node3420;
	wire [1-1:0] node3421;
	wire [1-1:0] node3422;
	wire [1-1:0] node3424;
	wire [1-1:0] node3425;
	wire [1-1:0] node3426;
	wire [1-1:0] node3431;
	wire [1-1:0] node3432;
	wire [1-1:0] node3433;
	wire [1-1:0] node3440;
	wire [1-1:0] node3441;
	wire [1-1:0] node3442;
	wire [1-1:0] node3443;
	wire [1-1:0] node3444;
	wire [1-1:0] node3445;
	wire [1-1:0] node3447;
	wire [1-1:0] node3448;
	wire [1-1:0] node3450;
	wire [1-1:0] node3454;
	wire [1-1:0] node3455;
	wire [1-1:0] node3457;
	wire [1-1:0] node3458;
	wire [1-1:0] node3463;
	wire [1-1:0] node3464;
	wire [1-1:0] node3465;
	wire [1-1:0] node3467;
	wire [1-1:0] node3468;
	wire [1-1:0] node3474;
	wire [1-1:0] node3475;
	wire [1-1:0] node3476;
	wire [1-1:0] node3477;
	wire [1-1:0] node3479;
	wire [1-1:0] node3480;
	wire [1-1:0] node3487;
	wire [1-1:0] node3488;
	wire [1-1:0] node3489;
	wire [1-1:0] node3490;
	wire [1-1:0] node3491;
	wire [1-1:0] node3495;
	wire [1-1:0] node3496;
	wire [1-1:0] node3497;
	wire [1-1:0] node3502;
	wire [1-1:0] node3503;
	wire [1-1:0] node3504;
	wire [1-1:0] node3505;
	wire [1-1:0] node3512;
	wire [1-1:0] node3513;
	wire [1-1:0] node3514;
	wire [1-1:0] node3515;
	wire [1-1:0] node3516;
	wire [1-1:0] node3517;
	wire [1-1:0] node3519;
	wire [1-1:0] node3523;
	wire [1-1:0] node3524;
	wire [1-1:0] node3525;
	wire [1-1:0] node3530;
	wire [1-1:0] node3531;
	wire [1-1:0] node3532;
	wire [1-1:0] node3533;
	wire [1-1:0] node3539;
	wire [1-1:0] node3540;
	wire [1-1:0] node3541;
	wire [1-1:0] node3542;
	wire [1-1:0] node3543;

	assign outp = (inp[4]) ? node1822 : node1;
		assign node1 = (inp[7]) ? node855 : node2;
			assign node2 = (inp[14]) ? node348 : node3;
				assign node3 = (inp[11]) ? node129 : node4;
					assign node4 = (inp[8]) ? node40 : node5;
						assign node5 = (inp[2]) ? node7 : 1'b1;
							assign node7 = (inp[5]) ? node9 : 1'b1;
								assign node9 = (inp[3]) ? node19 : node10;
									assign node10 = (inp[13]) ? node12 : 1'b1;
										assign node12 = (inp[1]) ? node14 : 1'b1;
											assign node14 = (inp[0]) ? node16 : 1'b1;
												assign node16 = (inp[9]) ? 1'b0 : 1'b1;
									assign node19 = (inp[1]) ? node25 : node20;
										assign node20 = (inp[13]) ? node22 : 1'b1;
											assign node22 = (inp[0]) ? 1'b0 : 1'b1;
										assign node25 = (inp[9]) ? node31 : node26;
											assign node26 = (inp[13]) ? node28 : 1'b1;
												assign node28 = (inp[0]) ? 1'b0 : 1'b1;
											assign node31 = (inp[10]) ? node35 : node32;
												assign node32 = (inp[12]) ? 1'b0 : 1'b1;
												assign node35 = (inp[6]) ? 1'b0 : node36;
													assign node36 = (inp[0]) ? 1'b0 : 1'b1;
						assign node40 = (inp[1]) ? node74 : node41;
							assign node41 = (inp[13]) ? node43 : 1'b1;
								assign node43 = (inp[0]) ? node53 : node44;
									assign node44 = (inp[5]) ? node46 : 1'b1;
										assign node46 = (inp[10]) ? node48 : 1'b1;
											assign node48 = (inp[12]) ? node50 : 1'b1;
												assign node50 = (inp[3]) ? 1'b0 : 1'b1;
									assign node53 = (inp[10]) ? node61 : node54;
										assign node54 = (inp[5]) ? node56 : 1'b1;
											assign node56 = (inp[3]) ? node58 : 1'b1;
												assign node58 = (inp[12]) ? 1'b0 : 1'b1;
										assign node61 = (inp[2]) ? node69 : node62;
											assign node62 = (inp[12]) ? node64 : 1'b1;
												assign node64 = (inp[3]) ? node66 : 1'b1;
													assign node66 = (inp[6]) ? 1'b0 : 1'b1;
											assign node69 = (inp[9]) ? 1'b0 : node70;
												assign node70 = (inp[6]) ? 1'b0 : 1'b1;
							assign node74 = (inp[3]) ? node88 : node75;
								assign node75 = (inp[10]) ? node77 : 1'b1;
									assign node77 = (inp[9]) ? node79 : 1'b1;
										assign node79 = (inp[13]) ? node81 : 1'b1;
											assign node81 = (inp[12]) ? 1'b0 : node82;
												assign node82 = (inp[5]) ? node84 : 1'b1;
													assign node84 = (inp[0]) ? 1'b0 : 1'b1;
								assign node88 = (inp[6]) ? node110 : node89;
									assign node89 = (inp[10]) ? node91 : 1'b1;
										assign node91 = (inp[12]) ? node99 : node92;
											assign node92 = (inp[13]) ? node94 : 1'b1;
												assign node94 = (inp[2]) ? node96 : 1'b1;
													assign node96 = (inp[5]) ? 1'b1 : 1'b0;
											assign node99 = (inp[5]) ? node105 : node100;
												assign node100 = (inp[0]) ? node102 : 1'b1;
													assign node102 = (inp[13]) ? 1'b0 : 1'b1;
												assign node105 = (inp[2]) ? 1'b0 : node106;
													assign node106 = (inp[0]) ? 1'b0 : 1'b1;
									assign node110 = (inp[5]) ? node124 : node111;
										assign node111 = (inp[2]) ? node119 : node112;
											assign node112 = (inp[12]) ? node114 : 1'b1;
												assign node114 = (inp[9]) ? node116 : 1'b1;
													assign node116 = (inp[0]) ? 1'b0 : 1'b1;
											assign node119 = (inp[12]) ? 1'b0 : node120;
												assign node120 = (inp[10]) ? 1'b0 : 1'b1;
										assign node124 = (inp[2]) ? 1'b0 : node125;
											assign node125 = (inp[10]) ? 1'b0 : 1'b1;
					assign node129 = (inp[12]) ? node219 : node130;
						assign node130 = (inp[13]) ? node160 : node131;
							assign node131 = (inp[9]) ? node133 : 1'b1;
								assign node133 = (inp[6]) ? node143 : node134;
									assign node134 = (inp[8]) ? node136 : 1'b1;
										assign node136 = (inp[3]) ? 1'b1 : node137;
											assign node137 = (inp[2]) ? node139 : 1'b1;
												assign node139 = (inp[10]) ? 1'b0 : 1'b1;
									assign node143 = (inp[0]) ? node151 : node144;
										assign node144 = (inp[10]) ? node146 : 1'b1;
											assign node146 = (inp[3]) ? node148 : 1'b1;
												assign node148 = (inp[5]) ? 1'b0 : 1'b1;
										assign node151 = (inp[1]) ? node153 : 1'b1;
											assign node153 = (inp[5]) ? node155 : 1'b1;
												assign node155 = (inp[2]) ? 1'b0 : node156;
													assign node156 = (inp[8]) ? 1'b0 : 1'b1;
							assign node160 = (inp[3]) ? node182 : node161;
								assign node161 = (inp[9]) ? node163 : 1'b1;
									assign node163 = (inp[6]) ? node165 : 1'b1;
										assign node165 = (inp[10]) ? node173 : node166;
											assign node166 = (inp[1]) ? node168 : 1'b1;
												assign node168 = (inp[2]) ? node170 : 1'b1;
													assign node170 = (inp[5]) ? 1'b0 : 1'b1;
											assign node173 = (inp[1]) ? node179 : node174;
												assign node174 = (inp[5]) ? node176 : 1'b1;
													assign node176 = (inp[2]) ? 1'b0 : 1'b1;
												assign node179 = (inp[8]) ? 1'b0 : 1'b1;
								assign node182 = (inp[0]) ? node198 : node183;
									assign node183 = (inp[2]) ? node185 : 1'b1;
										assign node185 = (inp[5]) ? node191 : node186;
											assign node186 = (inp[9]) ? node188 : 1'b1;
												assign node188 = (inp[6]) ? 1'b0 : 1'b1;
											assign node191 = (inp[8]) ? 1'b0 : node192;
												assign node192 = (inp[10]) ? node194 : 1'b1;
													assign node194 = (inp[1]) ? 1'b0 : 1'b1;
									assign node198 = (inp[8]) ? node214 : node199;
										assign node199 = (inp[2]) ? node207 : node200;
											assign node200 = (inp[5]) ? node202 : 1'b1;
												assign node202 = (inp[10]) ? node204 : 1'b1;
													assign node204 = (inp[1]) ? 1'b0 : 1'b0;
											assign node207 = (inp[10]) ? node211 : node208;
												assign node208 = (inp[5]) ? 1'b0 : 1'b1;
												assign node211 = (inp[9]) ? 1'b0 : 1'b1;
										assign node214 = (inp[6]) ? 1'b0 : node215;
											assign node215 = (inp[10]) ? 1'b0 : 1'b1;
						assign node219 = (inp[9]) ? node279 : node220;
							assign node220 = (inp[2]) ? node238 : node221;
								assign node221 = (inp[0]) ? node223 : 1'b1;
									assign node223 = (inp[13]) ? node225 : 1'b1;
										assign node225 = (inp[10]) ? node231 : node226;
											assign node226 = (inp[1]) ? node228 : 1'b1;
												assign node228 = (inp[6]) ? 1'b0 : 1'b1;
											assign node231 = (inp[8]) ? 1'b0 : node232;
												assign node232 = (inp[6]) ? node234 : 1'b1;
													assign node234 = (inp[1]) ? 1'b0 : 1'b1;
								assign node238 = (inp[0]) ? node256 : node239;
									assign node239 = (inp[3]) ? node247 : node240;
										assign node240 = (inp[5]) ? node242 : 1'b1;
											assign node242 = (inp[1]) ? node244 : 1'b1;
												assign node244 = (inp[13]) ? 1'b0 : 1'b1;
										assign node247 = (inp[13]) ? node253 : node248;
											assign node248 = (inp[5]) ? node250 : 1'b1;
												assign node250 = (inp[1]) ? 1'b0 : 1'b1;
											assign node253 = (inp[10]) ? 1'b0 : 1'b1;
									assign node256 = (inp[1]) ? node270 : node257;
										assign node257 = (inp[5]) ? node259 : 1'b1;
											assign node259 = (inp[8]) ? node265 : node260;
												assign node260 = (inp[6]) ? node262 : 1'b1;
													assign node262 = (inp[10]) ? 1'b0 : 1'b1;
												assign node265 = (inp[6]) ? 1'b0 : node266;
													assign node266 = (inp[3]) ? 1'b0 : 1'b0;
										assign node270 = (inp[3]) ? 1'b0 : node271;
											assign node271 = (inp[5]) ? 1'b0 : node272;
												assign node272 = (inp[6]) ? node274 : 1'b1;
													assign node274 = (inp[13]) ? 1'b0 : 1'b1;
							assign node279 = (inp[1]) ? node317 : node280;
								assign node280 = (inp[0]) ? node290 : node281;
									assign node281 = (inp[10]) ? node283 : 1'b1;
										assign node283 = (inp[2]) ? node285 : 1'b1;
											assign node285 = (inp[6]) ? 1'b0 : node286;
												assign node286 = (inp[8]) ? 1'b0 : 1'b1;
									assign node290 = (inp[5]) ? node304 : node291;
										assign node291 = (inp[3]) ? node293 : 1'b1;
											assign node293 = (inp[2]) ? node299 : node294;
												assign node294 = (inp[13]) ? node296 : 1'b1;
													assign node296 = (inp[10]) ? 1'b0 : 1'b1;
												assign node299 = (inp[8]) ? 1'b0 : node300;
													assign node300 = (inp[10]) ? 1'b0 : 1'b1;
										assign node304 = (inp[13]) ? 1'b0 : node305;
											assign node305 = (inp[2]) ? node311 : node306;
												assign node306 = (inp[6]) ? node308 : 1'b1;
													assign node308 = (inp[3]) ? 1'b0 : 1'b1;
												assign node311 = (inp[8]) ? 1'b0 : node312;
													assign node312 = (inp[3]) ? 1'b0 : 1'b1;
								assign node317 = (inp[10]) ? node337 : node318;
									assign node318 = (inp[6]) ? node328 : node319;
										assign node319 = (inp[5]) ? node321 : 1'b1;
											assign node321 = (inp[3]) ? node323 : 1'b1;
												assign node323 = (inp[2]) ? 1'b0 : node324;
													assign node324 = (inp[13]) ? 1'b0 : 1'b1;
										assign node328 = (inp[13]) ? 1'b0 : node329;
											assign node329 = (inp[2]) ? node331 : 1'b1;
												assign node331 = (inp[8]) ? 1'b0 : node332;
													assign node332 = (inp[5]) ? 1'b0 : 1'b1;
									assign node337 = (inp[5]) ? 1'b0 : node338;
										assign node338 = (inp[0]) ? 1'b0 : node339;
											assign node339 = (inp[13]) ? 1'b0 : node340;
												assign node340 = (inp[3]) ? node342 : 1'b1;
													assign node342 = (inp[8]) ? 1'b0 : 1'b1;
				assign node348 = (inp[0]) ? node586 : node349;
					assign node349 = (inp[2]) ? node457 : node350;
						assign node350 = (inp[12]) ? node382 : node351;
							assign node351 = (inp[10]) ? node353 : 1'b1;
								assign node353 = (inp[5]) ? node361 : node354;
									assign node354 = (inp[11]) ? node356 : 1'b1;
										assign node356 = (inp[9]) ? node358 : 1'b1;
											assign node358 = (inp[8]) ? 1'b0 : 1'b1;
									assign node361 = (inp[1]) ? node371 : node362;
										assign node362 = (inp[3]) ? node364 : 1'b1;
											assign node364 = (inp[8]) ? node366 : 1'b1;
												assign node366 = (inp[11]) ? node368 : 1'b1;
													assign node368 = (inp[13]) ? 1'b0 : 1'b1;
										assign node371 = (inp[9]) ? node377 : node372;
											assign node372 = (inp[8]) ? node374 : 1'b1;
												assign node374 = (inp[6]) ? 1'b0 : 1'b1;
											assign node377 = (inp[3]) ? 1'b0 : node378;
												assign node378 = (inp[6]) ? 1'b0 : 1'b1;
							assign node382 = (inp[3]) ? node410 : node383;
								assign node383 = (inp[6]) ? node385 : 1'b1;
									assign node385 = (inp[1]) ? node395 : node386;
										assign node386 = (inp[10]) ? node388 : 1'b1;
											assign node388 = (inp[8]) ? node390 : 1'b1;
												assign node390 = (inp[5]) ? node392 : 1'b1;
													assign node392 = (inp[13]) ? 1'b0 : 1'b1;
										assign node395 = (inp[8]) ? node401 : node396;
											assign node396 = (inp[10]) ? node398 : 1'b1;
												assign node398 = (inp[11]) ? 1'b0 : 1'b1;
											assign node401 = (inp[13]) ? node405 : node402;
												assign node402 = (inp[5]) ? 1'b0 : 1'b1;
												assign node405 = (inp[11]) ? 1'b0 : node406;
													assign node406 = (inp[10]) ? 1'b0 : 1'b1;
								assign node410 = (inp[9]) ? node426 : node411;
									assign node411 = (inp[10]) ? node413 : 1'b1;
										assign node413 = (inp[6]) ? node415 : 1'b1;
											assign node415 = (inp[11]) ? node421 : node416;
												assign node416 = (inp[13]) ? node418 : 1'b1;
													assign node418 = (inp[1]) ? 1'b0 : 1'b1;
												assign node421 = (inp[1]) ? 1'b0 : node422;
													assign node422 = (inp[13]) ? 1'b0 : 1'b1;
									assign node426 = (inp[5]) ? node444 : node427;
										assign node427 = (inp[10]) ? node433 : node428;
											assign node428 = (inp[8]) ? node430 : 1'b1;
												assign node430 = (inp[6]) ? 1'b0 : 1'b1;
											assign node433 = (inp[13]) ? node439 : node434;
												assign node434 = (inp[1]) ? node436 : 1'b1;
													assign node436 = (inp[6]) ? 1'b0 : 1'b1;
												assign node439 = (inp[6]) ? 1'b0 : node440;
													assign node440 = (inp[8]) ? 1'b0 : 1'b1;
										assign node444 = (inp[11]) ? node452 : node445;
											assign node445 = (inp[8]) ? node447 : 1'b1;
												assign node447 = (inp[10]) ? 1'b0 : node448;
													assign node448 = (inp[6]) ? 1'b0 : 1'b1;
											assign node452 = (inp[1]) ? 1'b0 : node453;
												assign node453 = (inp[10]) ? 1'b0 : 1'b1;
						assign node457 = (inp[6]) ? node515 : node458;
							assign node458 = (inp[8]) ? node474 : node459;
								assign node459 = (inp[10]) ? node461 : 1'b1;
									assign node461 = (inp[12]) ? node463 : 1'b1;
										assign node463 = (inp[11]) ? node465 : 1'b1;
											assign node465 = (inp[1]) ? node471 : node466;
												assign node466 = (inp[13]) ? node468 : 1'b1;
													assign node468 = (inp[3]) ? 1'b0 : 1'b1;
												assign node471 = (inp[5]) ? 1'b0 : 1'b1;
								assign node474 = (inp[9]) ? node492 : node475;
									assign node475 = (inp[3]) ? node477 : 1'b1;
										assign node477 = (inp[1]) ? node485 : node478;
											assign node478 = (inp[5]) ? node480 : 1'b1;
												assign node480 = (inp[13]) ? node482 : 1'b1;
													assign node482 = (inp[12]) ? 1'b0 : 1'b1;
											assign node485 = (inp[12]) ? 1'b0 : node486;
												assign node486 = (inp[11]) ? node488 : 1'b1;
													assign node488 = (inp[10]) ? 1'b0 : 1'b1;
									assign node492 = (inp[11]) ? node502 : node493;
										assign node493 = (inp[10]) ? node495 : 1'b1;
											assign node495 = (inp[3]) ? 1'b0 : node496;
												assign node496 = (inp[13]) ? node498 : 1'b1;
													assign node498 = (inp[12]) ? 1'b0 : 1'b0;
										assign node502 = (inp[1]) ? 1'b0 : node503;
											assign node503 = (inp[5]) ? node509 : node504;
												assign node504 = (inp[12]) ? node506 : 1'b1;
													assign node506 = (inp[10]) ? 1'b0 : 1'b1;
												assign node509 = (inp[13]) ? 1'b0 : node510;
													assign node510 = (inp[3]) ? 1'b0 : 1'b1;
							assign node515 = (inp[11]) ? node553 : node516;
								assign node516 = (inp[10]) ? node538 : node517;
									assign node517 = (inp[3]) ? node525 : node518;
										assign node518 = (inp[9]) ? 1'b1 : node519;
											assign node519 = (inp[13]) ? node521 : 1'b1;
												assign node521 = (inp[8]) ? 1'b0 : 1'b1;
										assign node525 = (inp[8]) ? node531 : node526;
											assign node526 = (inp[5]) ? node528 : 1'b1;
												assign node528 = (inp[9]) ? 1'b0 : 1'b1;
											assign node531 = (inp[13]) ? 1'b0 : node532;
												assign node532 = (inp[12]) ? node534 : 1'b1;
													assign node534 = (inp[5]) ? 1'b0 : 1'b1;
									assign node538 = (inp[12]) ? node548 : node539;
										assign node539 = (inp[3]) ? node541 : 1'b1;
											assign node541 = (inp[8]) ? 1'b0 : node542;
												assign node542 = (inp[13]) ? node544 : 1'b1;
													assign node544 = (inp[5]) ? 1'b0 : 1'b1;
										assign node548 = (inp[8]) ? 1'b0 : node549;
											assign node549 = (inp[13]) ? 1'b0 : 1'b1;
								assign node553 = (inp[8]) ? node573 : node554;
									assign node554 = (inp[9]) ? node560 : node555;
										assign node555 = (inp[5]) ? node557 : 1'b1;
											assign node557 = (inp[12]) ? 1'b0 : 1'b1;
										assign node560 = (inp[12]) ? 1'b0 : node561;
											assign node561 = (inp[1]) ? node567 : node562;
												assign node562 = (inp[3]) ? 1'b1 : node563;
													assign node563 = (inp[10]) ? 1'b0 : 1'b1;
												assign node567 = (inp[3]) ? 1'b0 : node568;
													assign node568 = (inp[10]) ? 1'b0 : 1'b1;
									assign node573 = (inp[10]) ? 1'b0 : node574;
										assign node574 = (inp[3]) ? node578 : node575;
											assign node575 = (inp[12]) ? 1'b0 : 1'b1;
											assign node578 = (inp[13]) ? 1'b0 : node579;
												assign node579 = (inp[1]) ? 1'b0 : node580;
													assign node580 = (inp[9]) ? 1'b0 : 1'b1;
					assign node586 = (inp[1]) ? node710 : node587;
						assign node587 = (inp[9]) ? node641 : node588;
							assign node588 = (inp[5]) ? node606 : node589;
								assign node589 = (inp[10]) ? node591 : 1'b1;
									assign node591 = (inp[13]) ? node593 : 1'b1;
										assign node593 = (inp[8]) ? node595 : 1'b1;
											assign node595 = (inp[12]) ? node601 : node596;
												assign node596 = (inp[6]) ? node598 : 1'b1;
													assign node598 = (inp[3]) ? 1'b0 : 1'b1;
												assign node601 = (inp[2]) ? 1'b0 : node602;
													assign node602 = (inp[11]) ? 1'b0 : 1'b1;
								assign node606 = (inp[8]) ? node624 : node607;
									assign node607 = (inp[11]) ? node609 : 1'b1;
										assign node609 = (inp[3]) ? node617 : node610;
											assign node610 = (inp[13]) ? node612 : 1'b1;
												assign node612 = (inp[6]) ? node614 : 1'b1;
													assign node614 = (inp[10]) ? 1'b0 : 1'b1;
											assign node617 = (inp[10]) ? 1'b0 : node618;
												assign node618 = (inp[2]) ? node620 : 1'b1;
													assign node620 = (inp[6]) ? 1'b0 : 1'b1;
									assign node624 = (inp[2]) ? node632 : node625;
										assign node625 = (inp[6]) ? node627 : 1'b1;
											assign node627 = (inp[12]) ? 1'b0 : node628;
												assign node628 = (inp[10]) ? 1'b0 : 1'b1;
										assign node632 = (inp[13]) ? 1'b0 : node633;
											assign node633 = (inp[12]) ? node635 : 1'b1;
												assign node635 = (inp[6]) ? 1'b0 : node636;
													assign node636 = (inp[10]) ? 1'b0 : 1'b0;
							assign node641 = (inp[8]) ? node677 : node642;
								assign node642 = (inp[3]) ? node654 : node643;
									assign node643 = (inp[10]) ? node645 : 1'b1;
										assign node645 = (inp[12]) ? node647 : 1'b1;
											assign node647 = (inp[5]) ? 1'b0 : node648;
												assign node648 = (inp[6]) ? node650 : 1'b1;
													assign node650 = (inp[2]) ? 1'b0 : 1'b1;
									assign node654 = (inp[12]) ? node670 : node655;
										assign node655 = (inp[10]) ? node663 : node656;
											assign node656 = (inp[11]) ? node658 : 1'b1;
												assign node658 = (inp[6]) ? node660 : 1'b1;
													assign node660 = (inp[13]) ? 1'b0 : 1'b1;
											assign node663 = (inp[6]) ? node665 : 1'b1;
												assign node665 = (inp[13]) ? 1'b0 : node666;
													assign node666 = (inp[2]) ? 1'b0 : 1'b1;
										assign node670 = (inp[6]) ? 1'b0 : node671;
											assign node671 = (inp[11]) ? 1'b0 : node672;
												assign node672 = (inp[10]) ? 1'b0 : 1'b1;
								assign node677 = (inp[5]) ? node703 : node678;
									assign node678 = (inp[10]) ? node684 : node679;
										assign node679 = (inp[2]) ? node681 : 1'b1;
											assign node681 = (inp[12]) ? 1'b0 : 1'b1;
										assign node684 = (inp[6]) ? node696 : node685;
											assign node685 = (inp[12]) ? node691 : node686;
												assign node686 = (inp[2]) ? node688 : 1'b1;
													assign node688 = (inp[11]) ? 1'b0 : 1'b1;
												assign node691 = (inp[13]) ? 1'b0 : node692;
													assign node692 = (inp[3]) ? 1'b0 : 1'b1;
											assign node696 = (inp[11]) ? 1'b0 : node697;
												assign node697 = (inp[12]) ? 1'b0 : node698;
													assign node698 = (inp[3]) ? 1'b0 : 1'b0;
									assign node703 = (inp[6]) ? 1'b0 : node704;
										assign node704 = (inp[3]) ? 1'b0 : node705;
											assign node705 = (inp[10]) ? 1'b0 : 1'b1;
						assign node710 = (inp[2]) ? node802 : node711;
							assign node711 = (inp[3]) ? node767 : node712;
								assign node712 = (inp[9]) ? node742 : node713;
									assign node713 = (inp[12]) ? node723 : node714;
										assign node714 = (inp[11]) ? node716 : 1'b1;
											assign node716 = (inp[8]) ? node718 : 1'b1;
												assign node718 = (inp[5]) ? node720 : 1'b1;
													assign node720 = (inp[10]) ? 1'b0 : 1'b1;
										assign node723 = (inp[6]) ? node731 : node724;
											assign node724 = (inp[5]) ? node726 : 1'b1;
												assign node726 = (inp[13]) ? node728 : 1'b1;
													assign node728 = (inp[10]) ? 1'b0 : 1'b1;
											assign node731 = (inp[11]) ? node737 : node732;
												assign node732 = (inp[10]) ? node734 : 1'b1;
													assign node734 = (inp[13]) ? 1'b0 : 1'b1;
												assign node737 = (inp[5]) ? node739 : 1'b0;
													assign node739 = (inp[13]) ? 1'b0 : 1'b1;
									assign node742 = (inp[10]) ? node752 : node743;
										assign node743 = (inp[8]) ? node745 : 1'b1;
											assign node745 = (inp[13]) ? 1'b0 : node746;
												assign node746 = (inp[6]) ? node748 : 1'b1;
													assign node748 = (inp[5]) ? 1'b0 : 1'b1;
										assign node752 = (inp[6]) ? node760 : node753;
											assign node753 = (inp[12]) ? 1'b0 : node754;
												assign node754 = (inp[8]) ? node756 : 1'b1;
													assign node756 = (inp[5]) ? 1'b0 : 1'b1;
											assign node760 = (inp[13]) ? 1'b0 : node761;
												assign node761 = (inp[5]) ? 1'b0 : node762;
													assign node762 = (inp[12]) ? 1'b0 : 1'b1;
								assign node767 = (inp[10]) ? node787 : node768;
									assign node768 = (inp[12]) ? node778 : node769;
										assign node769 = (inp[5]) ? node771 : 1'b1;
											assign node771 = (inp[6]) ? 1'b0 : node772;
												assign node772 = (inp[11]) ? node774 : 1'b1;
													assign node774 = (inp[9]) ? 1'b0 : 1'b0;
										assign node778 = (inp[13]) ? 1'b0 : node779;
											assign node779 = (inp[9]) ? node781 : 1'b1;
												assign node781 = (inp[8]) ? 1'b0 : node782;
													assign node782 = (inp[6]) ? 1'b0 : 1'b1;
									assign node787 = (inp[13]) ? 1'b0 : node788;
										assign node788 = (inp[9]) ? 1'b0 : node789;
											assign node789 = (inp[11]) ? node795 : node790;
												assign node790 = (inp[5]) ? node792 : 1'b1;
													assign node792 = (inp[12]) ? 1'b0 : 1'b1;
												assign node795 = (inp[12]) ? 1'b0 : node796;
													assign node796 = (inp[5]) ? 1'b0 : 1'b1;
							assign node802 = (inp[13]) ? node838 : node803;
								assign node803 = (inp[12]) ? node829 : node804;
									assign node804 = (inp[8]) ? node814 : node805;
										assign node805 = (inp[6]) ? node807 : 1'b1;
											assign node807 = (inp[3]) ? node809 : 1'b1;
												assign node809 = (inp[11]) ? 1'b0 : node810;
													assign node810 = (inp[10]) ? 1'b0 : 1'b1;
										assign node814 = (inp[9]) ? node824 : node815;
											assign node815 = (inp[11]) ? node819 : node816;
												assign node816 = (inp[3]) ? 1'b0 : 1'b1;
												assign node819 = (inp[5]) ? 1'b0 : node820;
													assign node820 = (inp[6]) ? 1'b0 : 1'b1;
											assign node824 = (inp[5]) ? 1'b0 : node825;
												assign node825 = (inp[6]) ? 1'b0 : 1'b1;
									assign node829 = (inp[9]) ? 1'b0 : node830;
										assign node830 = (inp[5]) ? 1'b0 : node831;
											assign node831 = (inp[6]) ? node833 : 1'b1;
												assign node833 = (inp[11]) ? 1'b0 : 1'b1;
								assign node838 = (inp[9]) ? 1'b0 : node839;
									assign node839 = (inp[6]) ? 1'b0 : node840;
										assign node840 = (inp[10]) ? node848 : node841;
											assign node841 = (inp[12]) ? node843 : 1'b0;
												assign node843 = (inp[3]) ? node845 : 1'b1;
													assign node845 = (inp[5]) ? 1'b0 : 1'b1;
											assign node848 = (inp[12]) ? 1'b0 : node849;
												assign node849 = (inp[8]) ? 1'b0 : 1'b1;
			assign node855 = (inp[2]) ? node1363 : node856;
				assign node856 = (inp[14]) ? node1070 : node857;
					assign node857 = (inp[3]) ? node937 : node858;
						assign node858 = (inp[1]) ? node890 : node859;
							assign node859 = (inp[9]) ? node861 : 1'b1;
								assign node861 = (inp[13]) ? node871 : node862;
									assign node862 = (inp[10]) ? node864 : 1'b1;
										assign node864 = (inp[6]) ? node866 : 1'b1;
											assign node866 = (inp[11]) ? node868 : 1'b1;
												assign node868 = (inp[8]) ? 1'b0 : 1'b1;
									assign node871 = (inp[6]) ? node879 : node872;
										assign node872 = (inp[8]) ? node874 : 1'b1;
											assign node874 = (inp[12]) ? node876 : 1'b1;
												assign node876 = (inp[0]) ? 1'b0 : 1'b1;
										assign node879 = (inp[10]) ? node885 : node880;
											assign node880 = (inp[0]) ? 1'b1 : node881;
												assign node881 = (inp[5]) ? 1'b0 : 1'b1;
											assign node885 = (inp[11]) ? 1'b0 : node886;
												assign node886 = (inp[8]) ? 1'b0 : 1'b1;
							assign node890 = (inp[13]) ? node910 : node891;
								assign node891 = (inp[10]) ? node893 : 1'b1;
									assign node893 = (inp[12]) ? node895 : 1'b1;
										assign node895 = (inp[5]) ? node903 : node896;
											assign node896 = (inp[9]) ? 1'b1 : node897;
												assign node897 = (inp[6]) ? node899 : 1'b1;
													assign node899 = (inp[11]) ? 1'b0 : 1'b1;
											assign node903 = (inp[9]) ? 1'b0 : node904;
												assign node904 = (inp[6]) ? node906 : 1'b1;
													assign node906 = (inp[8]) ? 1'b0 : 1'b1;
								assign node910 = (inp[0]) ? node916 : node911;
									assign node911 = (inp[12]) ? node913 : 1'b1;
										assign node913 = (inp[6]) ? 1'b0 : 1'b1;
									assign node916 = (inp[5]) ? node924 : node917;
										assign node917 = (inp[10]) ? node919 : 1'b1;
											assign node919 = (inp[6]) ? node921 : 1'b1;
												assign node921 = (inp[11]) ? 1'b0 : 1'b1;
										assign node924 = (inp[6]) ? 1'b0 : node925;
											assign node925 = (inp[11]) ? node931 : node926;
												assign node926 = (inp[12]) ? node928 : 1'b1;
													assign node928 = (inp[8]) ? 1'b0 : 1'b1;
												assign node931 = (inp[8]) ? 1'b0 : node932;
													assign node932 = (inp[12]) ? 1'b0 : 1'b1;
						assign node937 = (inp[9]) ? node987 : node938;
							assign node938 = (inp[0]) ? node952 : node939;
								assign node939 = (inp[10]) ? node941 : 1'b1;
									assign node941 = (inp[5]) ? node943 : 1'b1;
										assign node943 = (inp[13]) ? 1'b0 : node944;
											assign node944 = (inp[8]) ? node946 : 1'b1;
												assign node946 = (inp[6]) ? node948 : 1'b1;
													assign node948 = (inp[11]) ? 1'b0 : 1'b1;
								assign node952 = (inp[12]) ? node964 : node953;
									assign node953 = (inp[10]) ? node955 : 1'b1;
										assign node955 = (inp[13]) ? node957 : 1'b1;
											assign node957 = (inp[8]) ? 1'b0 : node958;
												assign node958 = (inp[11]) ? node960 : 1'b1;
													assign node960 = (inp[6]) ? 1'b0 : 1'b1;
									assign node964 = (inp[8]) ? node978 : node965;
										assign node965 = (inp[11]) ? node971 : node966;
											assign node966 = (inp[10]) ? node968 : 1'b1;
												assign node968 = (inp[1]) ? 1'b0 : 1'b1;
											assign node971 = (inp[1]) ? 1'b0 : node972;
												assign node972 = (inp[13]) ? node974 : 1'b1;
													assign node974 = (inp[5]) ? 1'b0 : 1'b0;
										assign node978 = (inp[13]) ? 1'b0 : node979;
											assign node979 = (inp[11]) ? node981 : 1'b1;
												assign node981 = (inp[6]) ? 1'b0 : node982;
													assign node982 = (inp[10]) ? 1'b0 : 1'b1;
							assign node987 = (inp[0]) ? node1031 : node988;
								assign node988 = (inp[12]) ? node1008 : node989;
									assign node989 = (inp[1]) ? node991 : 1'b1;
										assign node991 = (inp[5]) ? node997 : node992;
											assign node992 = (inp[6]) ? node994 : 1'b1;
												assign node994 = (inp[8]) ? 1'b0 : 1'b1;
											assign node997 = (inp[13]) ? node1003 : node998;
												assign node998 = (inp[11]) ? node1000 : 1'b1;
													assign node1000 = (inp[6]) ? 1'b0 : 1'b1;
												assign node1003 = (inp[8]) ? 1'b0 : node1004;
													assign node1004 = (inp[10]) ? 1'b0 : 1'b0;
									assign node1008 = (inp[13]) ? node1022 : node1009;
										assign node1009 = (inp[11]) ? node1015 : node1010;
											assign node1010 = (inp[6]) ? node1012 : 1'b1;
												assign node1012 = (inp[5]) ? 1'b0 : 1'b1;
											assign node1015 = (inp[8]) ? 1'b0 : node1016;
												assign node1016 = (inp[10]) ? node1018 : 1'b1;
													assign node1018 = (inp[1]) ? 1'b0 : 1'b1;
										assign node1022 = (inp[1]) ? 1'b0 : node1023;
											assign node1023 = (inp[8]) ? 1'b0 : node1024;
												assign node1024 = (inp[6]) ? node1026 : 1'b1;
													assign node1026 = (inp[11]) ? 1'b0 : 1'b1;
								assign node1031 = (inp[10]) ? node1059 : node1032;
									assign node1032 = (inp[6]) ? node1046 : node1033;
										assign node1033 = (inp[13]) ? node1039 : node1034;
											assign node1034 = (inp[5]) ? node1036 : 1'b1;
												assign node1036 = (inp[12]) ? 1'b0 : 1'b1;
											assign node1039 = (inp[11]) ? 1'b0 : node1040;
												assign node1040 = (inp[1]) ? node1042 : 1'b1;
													assign node1042 = (inp[8]) ? 1'b0 : 1'b1;
										assign node1046 = (inp[1]) ? node1052 : node1047;
											assign node1047 = (inp[8]) ? node1049 : 1'b1;
												assign node1049 = (inp[12]) ? 1'b0 : 1'b1;
											assign node1052 = (inp[13]) ? 1'b0 : node1053;
												assign node1053 = (inp[5]) ? 1'b0 : node1054;
													assign node1054 = (inp[12]) ? 1'b0 : 1'b1;
									assign node1059 = (inp[6]) ? 1'b0 : node1060;
										assign node1060 = (inp[11]) ? 1'b0 : node1061;
											assign node1061 = (inp[5]) ? 1'b0 : node1062;
												assign node1062 = (inp[12]) ? node1064 : 1'b1;
													assign node1064 = (inp[8]) ? 1'b0 : 1'b1;
					assign node1070 = (inp[10]) ? node1214 : node1071;
						assign node1071 = (inp[5]) ? node1137 : node1072;
							assign node1072 = (inp[0]) ? node1094 : node1073;
								assign node1073 = (inp[6]) ? node1075 : 1'b1;
									assign node1075 = (inp[11]) ? node1083 : node1076;
										assign node1076 = (inp[9]) ? node1078 : 1'b1;
											assign node1078 = (inp[8]) ? node1080 : 1'b1;
												assign node1080 = (inp[12]) ? 1'b0 : 1'b1;
										assign node1083 = (inp[3]) ? node1089 : node1084;
											assign node1084 = (inp[1]) ? node1086 : 1'b1;
												assign node1086 = (inp[12]) ? 1'b0 : 1'b1;
											assign node1089 = (inp[8]) ? 1'b0 : node1090;
												assign node1090 = (inp[12]) ? 1'b0 : 1'b1;
								assign node1094 = (inp[8]) ? node1112 : node1095;
									assign node1095 = (inp[11]) ? node1103 : node1096;
										assign node1096 = (inp[12]) ? node1098 : 1'b1;
											assign node1098 = (inp[9]) ? node1100 : 1'b1;
												assign node1100 = (inp[1]) ? 1'b0 : 1'b1;
										assign node1103 = (inp[3]) ? node1109 : node1104;
											assign node1104 = (inp[12]) ? node1106 : 1'b1;
												assign node1106 = (inp[6]) ? 1'b0 : 1'b1;
											assign node1109 = (inp[6]) ? 1'b0 : 1'b1;
									assign node1112 = (inp[13]) ? node1124 : node1113;
										assign node1113 = (inp[9]) ? node1121 : node1114;
											assign node1114 = (inp[3]) ? node1116 : 1'b1;
												assign node1116 = (inp[11]) ? node1118 : 1'b1;
													assign node1118 = (inp[6]) ? 1'b0 : 1'b1;
											assign node1121 = (inp[1]) ? 1'b0 : 1'b1;
										assign node1124 = (inp[12]) ? 1'b0 : node1125;
											assign node1125 = (inp[11]) ? node1131 : node1126;
												assign node1126 = (inp[3]) ? node1128 : 1'b1;
													assign node1128 = (inp[1]) ? 1'b0 : 1'b1;
												assign node1131 = (inp[6]) ? 1'b0 : node1132;
													assign node1132 = (inp[9]) ? 1'b0 : 1'b1;
							assign node1137 = (inp[12]) ? node1183 : node1138;
								assign node1138 = (inp[3]) ? node1160 : node1139;
									assign node1139 = (inp[1]) ? node1147 : node1140;
										assign node1140 = (inp[13]) ? node1142 : 1'b1;
											assign node1142 = (inp[0]) ? node1144 : 1'b1;
												assign node1144 = (inp[11]) ? 1'b0 : 1'b1;
										assign node1147 = (inp[11]) ? node1153 : node1148;
											assign node1148 = (inp[9]) ? node1150 : 1'b1;
												assign node1150 = (inp[6]) ? 1'b0 : 1'b1;
											assign node1153 = (inp[0]) ? 1'b0 : node1154;
												assign node1154 = (inp[6]) ? node1156 : 1'b1;
													assign node1156 = (inp[13]) ? 1'b0 : 1'b1;
									assign node1160 = (inp[11]) ? node1174 : node1161;
										assign node1161 = (inp[9]) ? node1167 : node1162;
											assign node1162 = (inp[13]) ? node1164 : 1'b1;
												assign node1164 = (inp[0]) ? 1'b0 : 1'b1;
											assign node1167 = (inp[1]) ? 1'b0 : node1168;
												assign node1168 = (inp[6]) ? node1170 : 1'b1;
													assign node1170 = (inp[0]) ? 1'b0 : 1'b1;
										assign node1174 = (inp[13]) ? 1'b0 : node1175;
											assign node1175 = (inp[6]) ? node1177 : 1'b1;
												assign node1177 = (inp[0]) ? 1'b0 : node1178;
													assign node1178 = (inp[9]) ? 1'b0 : 1'b1;
								assign node1183 = (inp[6]) ? node1203 : node1184;
									assign node1184 = (inp[8]) ? node1194 : node1185;
										assign node1185 = (inp[0]) ? node1187 : 1'b1;
											assign node1187 = (inp[1]) ? node1189 : 1'b1;
												assign node1189 = (inp[13]) ? 1'b0 : node1190;
													assign node1190 = (inp[3]) ? 1'b0 : 1'b1;
										assign node1194 = (inp[11]) ? 1'b0 : node1195;
											assign node1195 = (inp[1]) ? node1197 : 1'b1;
												assign node1197 = (inp[3]) ? 1'b0 : node1198;
													assign node1198 = (inp[9]) ? 1'b0 : 1'b1;
									assign node1203 = (inp[3]) ? 1'b0 : node1204;
										assign node1204 = (inp[13]) ? 1'b0 : node1205;
											assign node1205 = (inp[0]) ? node1207 : 1'b1;
												assign node1207 = (inp[9]) ? 1'b0 : node1208;
													assign node1208 = (inp[11]) ? 1'b0 : 1'b1;
						assign node1214 = (inp[5]) ? node1308 : node1215;
							assign node1215 = (inp[8]) ? node1257 : node1216;
								assign node1216 = (inp[12]) ? node1228 : node1217;
									assign node1217 = (inp[13]) ? node1219 : 1'b1;
										assign node1219 = (inp[1]) ? node1221 : 1'b1;
											assign node1221 = (inp[0]) ? 1'b0 : node1222;
												assign node1222 = (inp[11]) ? node1224 : 1'b1;
													assign node1224 = (inp[6]) ? 1'b0 : 1'b1;
									assign node1228 = (inp[3]) ? node1240 : node1229;
										assign node1229 = (inp[9]) ? node1237 : node1230;
											assign node1230 = (inp[1]) ? node1232 : 1'b1;
												assign node1232 = (inp[0]) ? node1234 : 1'b1;
													assign node1234 = (inp[6]) ? 1'b0 : 1'b1;
											assign node1237 = (inp[13]) ? 1'b0 : 1'b1;
										assign node1240 = (inp[1]) ? node1252 : node1241;
											assign node1241 = (inp[9]) ? node1247 : node1242;
												assign node1242 = (inp[13]) ? node1244 : 1'b1;
													assign node1244 = (inp[11]) ? 1'b0 : 1'b1;
												assign node1247 = (inp[0]) ? 1'b0 : node1248;
													assign node1248 = (inp[13]) ? 1'b0 : 1'b1;
											assign node1252 = (inp[13]) ? 1'b0 : node1253;
												assign node1253 = (inp[0]) ? 1'b0 : 1'b1;
								assign node1257 = (inp[6]) ? node1293 : node1258;
									assign node1258 = (inp[3]) ? node1278 : node1259;
										assign node1259 = (inp[0]) ? node1267 : node1260;
											assign node1260 = (inp[11]) ? node1262 : 1'b1;
												assign node1262 = (inp[12]) ? node1264 : 1'b1;
													assign node1264 = (inp[9]) ? 1'b0 : 1'b1;
											assign node1267 = (inp[11]) ? node1273 : node1268;
												assign node1268 = (inp[13]) ? node1270 : 1'b1;
													assign node1270 = (inp[12]) ? 1'b0 : 1'b1;
												assign node1273 = (inp[9]) ? 1'b0 : node1274;
													assign node1274 = (inp[1]) ? 1'b0 : 1'b1;
										assign node1278 = (inp[9]) ? node1286 : node1279;
											assign node1279 = (inp[13]) ? node1281 : 1'b1;
												assign node1281 = (inp[12]) ? 1'b0 : node1282;
													assign node1282 = (inp[11]) ? 1'b0 : 1'b1;
											assign node1286 = (inp[0]) ? 1'b0 : node1287;
												assign node1287 = (inp[12]) ? node1289 : 1'b1;
													assign node1289 = (inp[1]) ? 1'b0 : 1'b0;
									assign node1293 = (inp[1]) ? 1'b0 : node1294;
										assign node1294 = (inp[11]) ? 1'b0 : node1295;
											assign node1295 = (inp[0]) ? node1301 : node1296;
												assign node1296 = (inp[3]) ? node1298 : 1'b1;
													assign node1298 = (inp[12]) ? 1'b0 : 1'b1;
												assign node1301 = (inp[13]) ? 1'b0 : node1302;
													assign node1302 = (inp[3]) ? 1'b0 : 1'b1;
							assign node1308 = (inp[6]) ? node1344 : node1309;
								assign node1309 = (inp[0]) ? node1329 : node1310;
									assign node1310 = (inp[8]) ? node1320 : node1311;
										assign node1311 = (inp[3]) ? node1313 : 1'b1;
											assign node1313 = (inp[13]) ? node1315 : 1'b1;
												assign node1315 = (inp[1]) ? 1'b0 : node1316;
													assign node1316 = (inp[9]) ? 1'b0 : 1'b1;
										assign node1320 = (inp[11]) ? 1'b0 : node1321;
											assign node1321 = (inp[13]) ? 1'b0 : node1322;
												assign node1322 = (inp[1]) ? node1324 : 1'b1;
													assign node1324 = (inp[3]) ? 1'b0 : 1'b1;
									assign node1329 = (inp[13]) ? 1'b0 : node1330;
										assign node1330 = (inp[8]) ? node1336 : node1331;
											assign node1331 = (inp[9]) ? node1333 : 1'b1;
												assign node1333 = (inp[3]) ? 1'b0 : 1'b1;
											assign node1336 = (inp[11]) ? 1'b0 : node1337;
												assign node1337 = (inp[3]) ? 1'b0 : node1338;
													assign node1338 = (inp[1]) ? 1'b0 : 1'b0;
								assign node1344 = (inp[1]) ? 1'b0 : node1345;
									assign node1345 = (inp[9]) ? node1355 : node1346;
										assign node1346 = (inp[8]) ? 1'b0 : node1347;
											assign node1347 = (inp[12]) ? node1349 : 1'b1;
												assign node1349 = (inp[11]) ? 1'b0 : node1350;
													assign node1350 = (inp[13]) ? 1'b0 : 1'b1;
										assign node1355 = (inp[11]) ? 1'b0 : node1356;
											assign node1356 = (inp[8]) ? 1'b0 : node1357;
												assign node1357 = (inp[0]) ? 1'b0 : 1'b1;
				assign node1363 = (inp[5]) ? node1617 : node1364;
					assign node1364 = (inp[1]) ? node1482 : node1365;
						assign node1365 = (inp[8]) ? node1399 : node1366;
							assign node1366 = (inp[6]) ? node1378 : node1367;
								assign node1367 = (inp[10]) ? node1369 : 1'b1;
									assign node1369 = (inp[11]) ? node1371 : 1'b1;
										assign node1371 = (inp[3]) ? node1373 : 1'b1;
											assign node1373 = (inp[14]) ? 1'b0 : node1374;
												assign node1374 = (inp[9]) ? 1'b1 : 1'b0;
								assign node1378 = (inp[10]) ? node1386 : node1379;
									assign node1379 = (inp[13]) ? node1381 : 1'b1;
										assign node1381 = (inp[9]) ? node1383 : 1'b1;
											assign node1383 = (inp[11]) ? 1'b0 : 1'b1;
									assign node1386 = (inp[12]) ? node1392 : node1387;
										assign node1387 = (inp[0]) ? node1389 : 1'b1;
											assign node1389 = (inp[9]) ? 1'b0 : 1'b1;
										assign node1392 = (inp[0]) ? 1'b0 : node1393;
											assign node1393 = (inp[9]) ? node1395 : 1'b0;
												assign node1395 = (inp[3]) ? 1'b0 : 1'b1;
							assign node1399 = (inp[11]) ? node1433 : node1400;
								assign node1400 = (inp[6]) ? node1416 : node1401;
									assign node1401 = (inp[10]) ? node1403 : 1'b1;
										assign node1403 = (inp[0]) ? node1411 : node1404;
											assign node1404 = (inp[14]) ? node1406 : 1'b1;
												assign node1406 = (inp[3]) ? node1408 : 1'b1;
													assign node1408 = (inp[13]) ? 1'b0 : 1'b1;
											assign node1411 = (inp[12]) ? 1'b0 : node1412;
												assign node1412 = (inp[14]) ? 1'b0 : 1'b1;
									assign node1416 = (inp[13]) ? node1426 : node1417;
										assign node1417 = (inp[9]) ? node1419 : 1'b1;
											assign node1419 = (inp[10]) ? 1'b0 : node1420;
												assign node1420 = (inp[3]) ? node1422 : 1'b1;
													assign node1422 = (inp[0]) ? 1'b0 : 1'b1;
										assign node1426 = (inp[10]) ? 1'b0 : node1427;
											assign node1427 = (inp[0]) ? 1'b0 : node1428;
												assign node1428 = (inp[9]) ? 1'b0 : 1'b1;
								assign node1433 = (inp[3]) ? node1463 : node1434;
									assign node1434 = (inp[12]) ? node1452 : node1435;
										assign node1435 = (inp[13]) ? node1443 : node1436;
											assign node1436 = (inp[14]) ? node1438 : 1'b1;
												assign node1438 = (inp[6]) ? node1440 : 1'b1;
													assign node1440 = (inp[0]) ? 1'b0 : 1'b1;
											assign node1443 = (inp[10]) ? node1449 : node1444;
												assign node1444 = (inp[0]) ? node1446 : 1'b1;
													assign node1446 = (inp[14]) ? 1'b0 : 1'b1;
												assign node1449 = (inp[6]) ? 1'b0 : 1'b1;
										assign node1452 = (inp[14]) ? node1456 : node1453;
											assign node1453 = (inp[6]) ? 1'b0 : 1'b1;
											assign node1456 = (inp[6]) ? 1'b0 : node1457;
												assign node1457 = (inp[0]) ? 1'b0 : node1458;
													assign node1458 = (inp[9]) ? 1'b0 : 1'b1;
									assign node1463 = (inp[14]) ? 1'b0 : node1464;
										assign node1464 = (inp[9]) ? node1474 : node1465;
											assign node1465 = (inp[0]) ? node1471 : node1466;
												assign node1466 = (inp[10]) ? node1468 : 1'b1;
													assign node1468 = (inp[6]) ? 1'b0 : 1'b1;
												assign node1471 = (inp[6]) ? 1'b0 : 1'b1;
											assign node1474 = (inp[13]) ? 1'b0 : node1475;
												assign node1475 = (inp[12]) ? 1'b0 : node1476;
													assign node1476 = (inp[10]) ? 1'b0 : 1'b1;
						assign node1482 = (inp[12]) ? node1556 : node1483;
							assign node1483 = (inp[8]) ? node1519 : node1484;
								assign node1484 = (inp[11]) ? node1496 : node1485;
									assign node1485 = (inp[0]) ? node1487 : 1'b1;
										assign node1487 = (inp[10]) ? node1489 : 1'b1;
											assign node1489 = (inp[14]) ? 1'b0 : node1490;
												assign node1490 = (inp[9]) ? node1492 : 1'b1;
													assign node1492 = (inp[13]) ? 1'b0 : 1'b1;
									assign node1496 = (inp[10]) ? node1510 : node1497;
										assign node1497 = (inp[0]) ? node1503 : node1498;
											assign node1498 = (inp[9]) ? node1500 : 1'b1;
												assign node1500 = (inp[14]) ? 1'b0 : 1'b1;
											assign node1503 = (inp[6]) ? node1505 : 1'b1;
												assign node1505 = (inp[3]) ? 1'b0 : node1506;
													assign node1506 = (inp[14]) ? 1'b0 : 1'b1;
										assign node1510 = (inp[9]) ? 1'b0 : node1511;
											assign node1511 = (inp[14]) ? 1'b0 : node1512;
												assign node1512 = (inp[3]) ? node1514 : 1'b1;
													assign node1514 = (inp[6]) ? 1'b0 : 1'b1;
								assign node1519 = (inp[3]) ? node1541 : node1520;
									assign node1520 = (inp[11]) ? node1530 : node1521;
										assign node1521 = (inp[10]) ? node1523 : 1'b1;
											assign node1523 = (inp[14]) ? 1'b0 : node1524;
												assign node1524 = (inp[6]) ? node1526 : 1'b1;
													assign node1526 = (inp[13]) ? 1'b0 : 1'b1;
										assign node1530 = (inp[13]) ? 1'b0 : node1531;
											assign node1531 = (inp[6]) ? node1535 : node1532;
												assign node1532 = (inp[9]) ? 1'b0 : 1'b1;
												assign node1535 = (inp[14]) ? 1'b0 : node1536;
													assign node1536 = (inp[10]) ? 1'b0 : 1'b1;
									assign node1541 = (inp[0]) ? node1549 : node1542;
										assign node1542 = (inp[10]) ? 1'b0 : node1543;
											assign node1543 = (inp[9]) ? node1545 : 1'b1;
												assign node1545 = (inp[14]) ? 1'b0 : 1'b1;
										assign node1549 = (inp[14]) ? 1'b0 : node1550;
											assign node1550 = (inp[6]) ? 1'b0 : node1551;
												assign node1551 = (inp[13]) ? 1'b0 : 1'b1;
							assign node1556 = (inp[9]) ? node1586 : node1557;
								assign node1557 = (inp[10]) ? node1571 : node1558;
									assign node1558 = (inp[6]) ? node1566 : node1559;
										assign node1559 = (inp[13]) ? node1561 : 1'b1;
											assign node1561 = (inp[14]) ? node1563 : 1'b1;
												assign node1563 = (inp[11]) ? 1'b0 : 1'b1;
										assign node1566 = (inp[11]) ? 1'b0 : node1567;
											assign node1567 = (inp[0]) ? 1'b0 : 1'b1;
									assign node1571 = (inp[3]) ? 1'b0 : node1572;
										assign node1572 = (inp[14]) ? node1580 : node1573;
											assign node1573 = (inp[13]) ? 1'b0 : node1574;
												assign node1574 = (inp[0]) ? node1576 : 1'b1;
													assign node1576 = (inp[8]) ? 1'b0 : 1'b1;
											assign node1580 = (inp[6]) ? 1'b0 : node1581;
												assign node1581 = (inp[11]) ? 1'b0 : 1'b1;
								assign node1586 = (inp[14]) ? 1'b0 : node1587;
									assign node1587 = (inp[0]) ? node1607 : node1588;
										assign node1588 = (inp[13]) ? node1600 : node1589;
											assign node1589 = (inp[6]) ? node1595 : node1590;
												assign node1590 = (inp[10]) ? node1592 : 1'b1;
													assign node1592 = (inp[8]) ? 1'b0 : 1'b1;
												assign node1595 = (inp[8]) ? 1'b0 : node1596;
													assign node1596 = (inp[3]) ? 1'b0 : 1'b1;
											assign node1600 = (inp[11]) ? 1'b0 : node1601;
												assign node1601 = (inp[3]) ? 1'b0 : node1602;
													assign node1602 = (inp[6]) ? 1'b0 : 1'b1;
										assign node1607 = (inp[8]) ? 1'b0 : node1608;
											assign node1608 = (inp[11]) ? 1'b0 : node1609;
												assign node1609 = (inp[3]) ? 1'b0 : node1610;
													assign node1610 = (inp[6]) ? 1'b0 : 1'b1;
					assign node1617 = (inp[0]) ? node1751 : node1618;
						assign node1618 = (inp[14]) ? node1690 : node1619;
							assign node1619 = (inp[10]) ? node1659 : node1620;
								assign node1620 = (inp[9]) ? node1632 : node1621;
									assign node1621 = (inp[13]) ? node1623 : 1'b1;
										assign node1623 = (inp[3]) ? node1625 : 1'b1;
											assign node1625 = (inp[11]) ? 1'b0 : node1626;
												assign node1626 = (inp[8]) ? node1628 : 1'b1;
													assign node1628 = (inp[12]) ? 1'b0 : 1'b1;
									assign node1632 = (inp[1]) ? node1646 : node1633;
										assign node1633 = (inp[13]) ? node1635 : 1'b1;
											assign node1635 = (inp[12]) ? node1641 : node1636;
												assign node1636 = (inp[3]) ? node1638 : 1'b1;
													assign node1638 = (inp[11]) ? 1'b0 : 1'b1;
												assign node1641 = (inp[6]) ? 1'b0 : node1642;
													assign node1642 = (inp[11]) ? 1'b0 : 1'b1;
										assign node1646 = (inp[6]) ? node1652 : node1647;
											assign node1647 = (inp[3]) ? 1'b1 : node1648;
												assign node1648 = (inp[11]) ? 1'b0 : 1'b1;
											assign node1652 = (inp[3]) ? 1'b0 : node1653;
												assign node1653 = (inp[13]) ? 1'b0 : node1654;
													assign node1654 = (inp[8]) ? 1'b0 : 1'b1;
								assign node1659 = (inp[6]) ? node1675 : node1660;
									assign node1660 = (inp[3]) ? node1670 : node1661;
										assign node1661 = (inp[8]) ? node1663 : 1'b1;
											assign node1663 = (inp[12]) ? node1665 : 1'b1;
												assign node1665 = (inp[1]) ? 1'b0 : node1666;
													assign node1666 = (inp[9]) ? 1'b0 : 1'b1;
										assign node1670 = (inp[12]) ? 1'b0 : node1671;
											assign node1671 = (inp[13]) ? 1'b0 : 1'b1;
									assign node1675 = (inp[13]) ? 1'b0 : node1676;
										assign node1676 = (inp[8]) ? 1'b0 : node1677;
											assign node1677 = (inp[9]) ? node1683 : node1678;
												assign node1678 = (inp[3]) ? node1680 : 1'b1;
													assign node1680 = (inp[1]) ? 1'b0 : 1'b1;
												assign node1683 = (inp[11]) ? 1'b0 : node1684;
													assign node1684 = (inp[12]) ? 1'b0 : 1'b1;
							assign node1690 = (inp[11]) ? node1738 : node1691;
								assign node1691 = (inp[13]) ? node1717 : node1692;
									assign node1692 = (inp[9]) ? node1708 : node1693;
										assign node1693 = (inp[3]) ? node1701 : node1694;
											assign node1694 = (inp[10]) ? node1696 : 1'b1;
												assign node1696 = (inp[12]) ? node1698 : 1'b1;
													assign node1698 = (inp[1]) ? 1'b0 : 1'b1;
											assign node1701 = (inp[1]) ? 1'b0 : node1702;
												assign node1702 = (inp[10]) ? node1704 : 1'b1;
													assign node1704 = (inp[6]) ? 1'b0 : 1'b1;
										assign node1708 = (inp[6]) ? 1'b0 : node1709;
											assign node1709 = (inp[8]) ? node1711 : 1'b1;
												assign node1711 = (inp[10]) ? 1'b0 : node1712;
													assign node1712 = (inp[12]) ? 1'b0 : 1'b1;
									assign node1717 = (inp[1]) ? node1731 : node1718;
										assign node1718 = (inp[8]) ? node1726 : node1719;
											assign node1719 = (inp[12]) ? node1723 : node1720;
												assign node1720 = (inp[6]) ? 1'b0 : 1'b1;
												assign node1723 = (inp[10]) ? 1'b0 : 1'b1;
											assign node1726 = (inp[6]) ? 1'b0 : node1727;
												assign node1727 = (inp[12]) ? 1'b0 : 1'b1;
										assign node1731 = (inp[3]) ? 1'b0 : node1732;
											assign node1732 = (inp[6]) ? 1'b0 : node1733;
												assign node1733 = (inp[10]) ? 1'b0 : 1'b1;
								assign node1738 = (inp[6]) ? 1'b0 : node1739;
									assign node1739 = (inp[12]) ? 1'b0 : node1740;
										assign node1740 = (inp[9]) ? 1'b0 : node1741;
											assign node1741 = (inp[3]) ? node1743 : 1'b1;
												assign node1743 = (inp[10]) ? node1745 : 1'b0;
													assign node1745 = (inp[1]) ? 1'b0 : 1'b1;
						assign node1751 = (inp[11]) ? node1805 : node1752;
							assign node1752 = (inp[8]) ? node1784 : node1753;
								assign node1753 = (inp[1]) ? node1769 : node1754;
									assign node1754 = (inp[14]) ? node1762 : node1755;
										assign node1755 = (inp[6]) ? node1757 : 1'b1;
											assign node1757 = (inp[9]) ? 1'b1 : node1758;
												assign node1758 = (inp[12]) ? 1'b0 : 1'b1;
										assign node1762 = (inp[12]) ? 1'b0 : node1763;
											assign node1763 = (inp[9]) ? node1765 : 1'b1;
												assign node1765 = (inp[3]) ? 1'b0 : 1'b1;
									assign node1769 = (inp[6]) ? 1'b0 : node1770;
										assign node1770 = (inp[14]) ? 1'b0 : node1771;
											assign node1771 = (inp[3]) ? node1777 : node1772;
												assign node1772 = (inp[13]) ? node1774 : 1'b1;
													assign node1774 = (inp[9]) ? 1'b0 : 1'b1;
												assign node1777 = (inp[10]) ? 1'b0 : node1778;
													assign node1778 = (inp[13]) ? 1'b0 : 1'b1;
								assign node1784 = (inp[3]) ? 1'b0 : node1785;
									assign node1785 = (inp[13]) ? node1797 : node1786;
										assign node1786 = (inp[6]) ? node1792 : node1787;
											assign node1787 = (inp[1]) ? node1789 : 1'b1;
												assign node1789 = (inp[14]) ? 1'b0 : 1'b1;
											assign node1792 = (inp[14]) ? 1'b0 : node1793;
												assign node1793 = (inp[12]) ? 1'b0 : 1'b1;
										assign node1797 = (inp[9]) ? 1'b0 : node1798;
											assign node1798 = (inp[14]) ? 1'b0 : node1799;
												assign node1799 = (inp[1]) ? 1'b0 : 1'b1;
							assign node1805 = (inp[9]) ? 1'b0 : node1806;
								assign node1806 = (inp[8]) ? 1'b0 : node1807;
									assign node1807 = (inp[14]) ? 1'b0 : node1808;
										assign node1808 = (inp[12]) ? node1814 : node1809;
											assign node1809 = (inp[3]) ? node1811 : 1'b1;
												assign node1811 = (inp[6]) ? 1'b0 : 1'b1;
											assign node1814 = (inp[6]) ? 1'b0 : node1815;
												assign node1815 = (inp[1]) ? 1'b0 : 1'b1;
		assign node1822 = (inp[3]) ? node2766 : node1823;
			assign node1823 = (inp[12]) ? node2313 : node1824;
				assign node1824 = (inp[6]) ? node2040 : node1825;
					assign node1825 = (inp[0]) ? node1909 : node1826;
						assign node1826 = (inp[11]) ? node1850 : node1827;
							assign node1827 = (inp[1]) ? node1829 : 1'b1;
								assign node1829 = (inp[9]) ? node1839 : node1830;
									assign node1830 = (inp[8]) ? node1832 : 1'b1;
										assign node1832 = (inp[2]) ? node1834 : 1'b1;
											assign node1834 = (inp[14]) ? node1836 : 1'b1;
												assign node1836 = (inp[5]) ? 1'b0 : 1'b1;
									assign node1839 = (inp[14]) ? node1841 : 1'b1;
										assign node1841 = (inp[13]) ? node1843 : 1'b1;
											assign node1843 = (inp[7]) ? 1'b0 : node1844;
												assign node1844 = (inp[10]) ? node1846 : 1'b1;
													assign node1846 = (inp[5]) ? 1'b0 : 1'b0;
							assign node1850 = (inp[7]) ? node1868 : node1851;
								assign node1851 = (inp[14]) ? node1853 : 1'b1;
									assign node1853 = (inp[5]) ? node1855 : 1'b1;
										assign node1855 = (inp[9]) ? node1857 : 1'b1;
											assign node1857 = (inp[8]) ? node1863 : node1858;
												assign node1858 = (inp[1]) ? node1860 : 1'b1;
													assign node1860 = (inp[2]) ? 1'b0 : 1'b1;
												assign node1863 = (inp[13]) ? 1'b0 : node1864;
													assign node1864 = (inp[2]) ? 1'b0 : 1'b1;
								assign node1868 = (inp[2]) ? node1890 : node1869;
									assign node1869 = (inp[14]) ? node1871 : 1'b1;
										assign node1871 = (inp[1]) ? node1879 : node1872;
											assign node1872 = (inp[10]) ? 1'b1 : node1873;
												assign node1873 = (inp[9]) ? node1875 : 1'b1;
													assign node1875 = (inp[5]) ? 1'b0 : 1'b1;
											assign node1879 = (inp[10]) ? node1885 : node1880;
												assign node1880 = (inp[8]) ? node1882 : 1'b1;
													assign node1882 = (inp[5]) ? 1'b0 : 1'b1;
												assign node1885 = (inp[13]) ? 1'b0 : node1886;
													assign node1886 = (inp[5]) ? 1'b0 : 1'b1;
									assign node1890 = (inp[8]) ? node1898 : node1891;
										assign node1891 = (inp[10]) ? node1893 : 1'b1;
											assign node1893 = (inp[14]) ? 1'b0 : node1894;
												assign node1894 = (inp[13]) ? 1'b0 : 1'b1;
										assign node1898 = (inp[14]) ? 1'b0 : node1899;
											assign node1899 = (inp[13]) ? node1903 : node1900;
												assign node1900 = (inp[1]) ? 1'b0 : 1'b1;
												assign node1903 = (inp[9]) ? 1'b0 : node1904;
													assign node1904 = (inp[10]) ? 1'b0 : 1'b1;
						assign node1909 = (inp[14]) ? node1969 : node1910;
							assign node1910 = (inp[1]) ? node1932 : node1911;
								assign node1911 = (inp[5]) ? node1913 : 1'b1;
									assign node1913 = (inp[7]) ? node1921 : node1914;
										assign node1914 = (inp[8]) ? node1916 : 1'b1;
											assign node1916 = (inp[13]) ? node1918 : 1'b1;
												assign node1918 = (inp[11]) ? 1'b0 : 1'b1;
										assign node1921 = (inp[2]) ? node1929 : node1922;
											assign node1922 = (inp[9]) ? node1924 : 1'b1;
												assign node1924 = (inp[13]) ? node1926 : 1'b1;
													assign node1926 = (inp[11]) ? 1'b0 : 1'b1;
											assign node1929 = (inp[8]) ? 1'b0 : 1'b1;
								assign node1932 = (inp[13]) ? node1942 : node1933;
									assign node1933 = (inp[2]) ? node1935 : 1'b1;
										assign node1935 = (inp[5]) ? node1937 : 1'b1;
											assign node1937 = (inp[10]) ? node1939 : 1'b1;
												assign node1939 = (inp[7]) ? 1'b0 : 1'b1;
									assign node1942 = (inp[2]) ? node1960 : node1943;
										assign node1943 = (inp[10]) ? node1951 : node1944;
											assign node1944 = (inp[5]) ? node1946 : 1'b1;
												assign node1946 = (inp[9]) ? node1948 : 1'b1;
													assign node1948 = (inp[7]) ? 1'b0 : 1'b1;
											assign node1951 = (inp[11]) ? node1957 : node1952;
												assign node1952 = (inp[7]) ? node1954 : 1'b1;
													assign node1954 = (inp[8]) ? 1'b0 : 1'b1;
												assign node1957 = (inp[9]) ? 1'b0 : 1'b1;
										assign node1960 = (inp[11]) ? 1'b0 : node1961;
											assign node1961 = (inp[9]) ? 1'b0 : node1962;
												assign node1962 = (inp[5]) ? node1964 : 1'b1;
													assign node1964 = (inp[7]) ? 1'b0 : 1'b0;
							assign node1969 = (inp[8]) ? node2003 : node1970;
								assign node1970 = (inp[13]) ? node1982 : node1971;
									assign node1971 = (inp[9]) ? node1973 : 1'b1;
										assign node1973 = (inp[2]) ? node1975 : 1'b1;
											assign node1975 = (inp[10]) ? node1977 : 1'b1;
												assign node1977 = (inp[1]) ? 1'b0 : node1978;
													assign node1978 = (inp[7]) ? 1'b0 : 1'b0;
									assign node1982 = (inp[9]) ? node1992 : node1983;
										assign node1983 = (inp[11]) ? node1985 : 1'b1;
											assign node1985 = (inp[2]) ? 1'b0 : node1986;
												assign node1986 = (inp[7]) ? node1988 : 1'b1;
													assign node1988 = (inp[5]) ? 1'b0 : 1'b1;
										assign node1992 = (inp[11]) ? 1'b0 : node1993;
											assign node1993 = (inp[10]) ? node1997 : node1994;
												assign node1994 = (inp[5]) ? 1'b0 : 1'b1;
												assign node1997 = (inp[7]) ? 1'b0 : node1998;
													assign node1998 = (inp[1]) ? 1'b0 : 1'b1;
								assign node2003 = (inp[10]) ? node2027 : node2004;
									assign node2004 = (inp[9]) ? node2020 : node2005;
										assign node2005 = (inp[5]) ? node2011 : node2006;
											assign node2006 = (inp[2]) ? node2008 : 1'b1;
												assign node2008 = (inp[13]) ? 1'b0 : 1'b1;
											assign node2011 = (inp[7]) ? node2017 : node2012;
												assign node2012 = (inp[1]) ? node2014 : 1'b1;
													assign node2014 = (inp[2]) ? 1'b0 : 1'b1;
												assign node2017 = (inp[11]) ? 1'b0 : 1'b1;
										assign node2020 = (inp[11]) ? 1'b0 : node2021;
											assign node2021 = (inp[2]) ? 1'b0 : node2022;
												assign node2022 = (inp[13]) ? 1'b0 : 1'b1;
									assign node2027 = (inp[1]) ? 1'b0 : node2028;
										assign node2028 = (inp[11]) ? 1'b0 : node2029;
											assign node2029 = (inp[5]) ? node2035 : node2030;
												assign node2030 = (inp[9]) ? node2032 : 1'b1;
													assign node2032 = (inp[7]) ? 1'b0 : 1'b1;
												assign node2035 = (inp[13]) ? 1'b0 : 1'b1;
					assign node2040 = (inp[10]) ? node2192 : node2041;
						assign node2041 = (inp[13]) ? node2113 : node2042;
							assign node2042 = (inp[9]) ? node2072 : node2043;
								assign node2043 = (inp[5]) ? node2051 : node2044;
									assign node2044 = (inp[0]) ? 1'b1 : node2045;
										assign node2045 = (inp[1]) ? node2047 : 1'b1;
											assign node2047 = (inp[7]) ? 1'b0 : 1'b1;
									assign node2051 = (inp[14]) ? node2059 : node2052;
										assign node2052 = (inp[8]) ? node2054 : 1'b1;
											assign node2054 = (inp[0]) ? node2056 : 1'b1;
												assign node2056 = (inp[1]) ? 1'b0 : 1'b1;
										assign node2059 = (inp[11]) ? node2061 : 1'b1;
											assign node2061 = (inp[0]) ? node2067 : node2062;
												assign node2062 = (inp[8]) ? node2064 : 1'b1;
													assign node2064 = (inp[1]) ? 1'b0 : 1'b1;
												assign node2067 = (inp[1]) ? 1'b0 : node2068;
													assign node2068 = (inp[2]) ? 1'b0 : 1'b1;
								assign node2072 = (inp[8]) ? node2094 : node2073;
									assign node2073 = (inp[5]) ? node2083 : node2074;
										assign node2074 = (inp[1]) ? node2076 : 1'b1;
											assign node2076 = (inp[7]) ? node2078 : 1'b1;
												assign node2078 = (inp[11]) ? node2080 : 1'b1;
													assign node2080 = (inp[2]) ? 1'b0 : 1'b1;
										assign node2083 = (inp[0]) ? node2089 : node2084;
											assign node2084 = (inp[2]) ? node2086 : 1'b1;
												assign node2086 = (inp[11]) ? 1'b0 : 1'b1;
											assign node2089 = (inp[1]) ? 1'b0 : node2090;
												assign node2090 = (inp[11]) ? 1'b0 : 1'b1;
									assign node2094 = (inp[1]) ? node2104 : node2095;
										assign node2095 = (inp[7]) ? node2097 : 1'b1;
											assign node2097 = (inp[5]) ? 1'b0 : node2098;
												assign node2098 = (inp[11]) ? node2100 : 1'b1;
													assign node2100 = (inp[2]) ? 1'b0 : 1'b0;
										assign node2104 = (inp[2]) ? 1'b0 : node2105;
											assign node2105 = (inp[0]) ? node2107 : 1'b1;
												assign node2107 = (inp[7]) ? node2109 : 1'b0;
													assign node2109 = (inp[14]) ? 1'b0 : 1'b1;
							assign node2113 = (inp[8]) ? node2155 : node2114;
								assign node2114 = (inp[9]) ? node2130 : node2115;
									assign node2115 = (inp[1]) ? node2117 : 1'b1;
										assign node2117 = (inp[14]) ? node2125 : node2118;
											assign node2118 = (inp[2]) ? node2120 : 1'b1;
												assign node2120 = (inp[0]) ? node2122 : 1'b1;
													assign node2122 = (inp[5]) ? 1'b0 : 1'b1;
											assign node2125 = (inp[11]) ? 1'b0 : node2126;
												assign node2126 = (inp[2]) ? 1'b0 : 1'b1;
									assign node2130 = (inp[5]) ? node2140 : node2131;
										assign node2131 = (inp[7]) ? node2133 : 1'b1;
											assign node2133 = (inp[1]) ? node2135 : 1'b1;
												assign node2135 = (inp[14]) ? 1'b0 : node2136;
													assign node2136 = (inp[2]) ? 1'b0 : 1'b1;
										assign node2140 = (inp[11]) ? node2148 : node2141;
											assign node2141 = (inp[0]) ? node2143 : 1'b1;
												assign node2143 = (inp[1]) ? 1'b0 : node2144;
													assign node2144 = (inp[2]) ? 1'b0 : 1'b1;
											assign node2148 = (inp[0]) ? node2150 : 1'b0;
												assign node2150 = (inp[1]) ? 1'b0 : node2151;
													assign node2151 = (inp[7]) ? 1'b0 : 1'b0;
								assign node2155 = (inp[5]) ? node2171 : node2156;
									assign node2156 = (inp[14]) ? node2162 : node2157;
										assign node2157 = (inp[7]) ? node2159 : 1'b1;
											assign node2159 = (inp[11]) ? 1'b0 : 1'b1;
										assign node2162 = (inp[2]) ? 1'b0 : node2163;
											assign node2163 = (inp[11]) ? node2165 : 1'b1;
												assign node2165 = (inp[7]) ? 1'b0 : node2166;
													assign node2166 = (inp[9]) ? 1'b0 : 1'b1;
									assign node2171 = (inp[1]) ? node2185 : node2172;
										assign node2172 = (inp[7]) ? node2180 : node2173;
											assign node2173 = (inp[9]) ? node2175 : 1'b1;
												assign node2175 = (inp[0]) ? 1'b0 : node2176;
													assign node2176 = (inp[11]) ? 1'b0 : 1'b1;
											assign node2180 = (inp[14]) ? 1'b0 : node2181;
												assign node2181 = (inp[2]) ? 1'b0 : 1'b1;
										assign node2185 = (inp[0]) ? 1'b0 : node2186;
											assign node2186 = (inp[14]) ? 1'b0 : node2187;
												assign node2187 = (inp[9]) ? 1'b0 : 1'b1;
						assign node2192 = (inp[7]) ? node2260 : node2193;
							assign node2193 = (inp[1]) ? node2229 : node2194;
								assign node2194 = (inp[5]) ? node2206 : node2195;
									assign node2195 = (inp[0]) ? node2197 : 1'b1;
										assign node2197 = (inp[14]) ? node2199 : 1'b1;
											assign node2199 = (inp[2]) ? node2201 : 1'b1;
												assign node2201 = (inp[11]) ? 1'b0 : node2202;
													assign node2202 = (inp[9]) ? 1'b0 : 1'b1;
									assign node2206 = (inp[9]) ? node2222 : node2207;
										assign node2207 = (inp[8]) ? node2215 : node2208;
											assign node2208 = (inp[13]) ? node2210 : 1'b1;
												assign node2210 = (inp[0]) ? 1'b1 : node2211;
													assign node2211 = (inp[14]) ? 1'b0 : 1'b1;
											assign node2215 = (inp[0]) ? 1'b0 : node2216;
												assign node2216 = (inp[11]) ? node2218 : 1'b1;
													assign node2218 = (inp[14]) ? 1'b0 : 1'b1;
										assign node2222 = (inp[8]) ? 1'b0 : node2223;
											assign node2223 = (inp[13]) ? 1'b0 : node2224;
												assign node2224 = (inp[11]) ? 1'b0 : 1'b1;
								assign node2229 = (inp[13]) ? node2251 : node2230;
									assign node2230 = (inp[2]) ? node2246 : node2231;
										assign node2231 = (inp[9]) ? node2239 : node2232;
											assign node2232 = (inp[8]) ? node2234 : 1'b1;
												assign node2234 = (inp[0]) ? node2236 : 1'b1;
													assign node2236 = (inp[11]) ? 1'b0 : 1'b1;
											assign node2239 = (inp[8]) ? 1'b0 : node2240;
												assign node2240 = (inp[14]) ? node2242 : 1'b1;
													assign node2242 = (inp[5]) ? 1'b0 : 1'b1;
										assign node2246 = (inp[0]) ? 1'b0 : node2247;
											assign node2247 = (inp[11]) ? 1'b0 : 1'b1;
									assign node2251 = (inp[8]) ? 1'b0 : node2252;
										assign node2252 = (inp[14]) ? 1'b0 : node2253;
											assign node2253 = (inp[9]) ? node2255 : 1'b1;
												assign node2255 = (inp[11]) ? 1'b0 : 1'b1;
							assign node2260 = (inp[2]) ? node2294 : node2261;
								assign node2261 = (inp[5]) ? node2279 : node2262;
									assign node2262 = (inp[11]) ? node2272 : node2263;
										assign node2263 = (inp[14]) ? node2265 : 1'b1;
											assign node2265 = (inp[8]) ? node2267 : 1'b1;
												assign node2267 = (inp[13]) ? node2269 : 1'b1;
													assign node2269 = (inp[9]) ? 1'b0 : 1'b0;
										assign node2272 = (inp[0]) ? 1'b0 : node2273;
											assign node2273 = (inp[9]) ? node2275 : 1'b1;
												assign node2275 = (inp[14]) ? 1'b0 : 1'b1;
									assign node2279 = (inp[14]) ? 1'b0 : node2280;
										assign node2280 = (inp[8]) ? node2286 : node2281;
											assign node2281 = (inp[0]) ? node2283 : 1'b1;
												assign node2283 = (inp[13]) ? 1'b0 : 1'b1;
											assign node2286 = (inp[0]) ? 1'b0 : node2287;
												assign node2287 = (inp[1]) ? 1'b0 : node2288;
													assign node2288 = (inp[13]) ? 1'b0 : 1'b1;
								assign node2294 = (inp[0]) ? 1'b0 : node2295;
									assign node2295 = (inp[14]) ? node2305 : node2296;
										assign node2296 = (inp[5]) ? 1'b0 : node2297;
											assign node2297 = (inp[13]) ? 1'b0 : node2298;
												assign node2298 = (inp[11]) ? node2300 : 1'b1;
													assign node2300 = (inp[1]) ? 1'b0 : 1'b1;
										assign node2305 = (inp[9]) ? 1'b0 : node2306;
											assign node2306 = (inp[5]) ? node2308 : 1'b0;
												assign node2308 = (inp[11]) ? 1'b0 : 1'b1;
				assign node2313 = (inp[5]) ? node2579 : node2314;
					assign node2314 = (inp[8]) ? node2444 : node2315;
						assign node2315 = (inp[2]) ? node2379 : node2316;
							assign node2316 = (inp[11]) ? node2342 : node2317;
								assign node2317 = (inp[1]) ? node2319 : 1'b1;
									assign node2319 = (inp[13]) ? node2329 : node2320;
										assign node2320 = (inp[9]) ? node2322 : 1'b1;
											assign node2322 = (inp[7]) ? node2324 : 1'b1;
												assign node2324 = (inp[6]) ? node2326 : 1'b1;
													assign node2326 = (inp[10]) ? 1'b0 : 1'b1;
										assign node2329 = (inp[7]) ? node2335 : node2330;
											assign node2330 = (inp[9]) ? node2332 : 1'b1;
												assign node2332 = (inp[14]) ? 1'b0 : 1'b1;
											assign node2335 = (inp[0]) ? node2337 : 1'b1;
												assign node2337 = (inp[10]) ? 1'b0 : node2338;
													assign node2338 = (inp[6]) ? 1'b0 : 1'b1;
								assign node2342 = (inp[14]) ? node2360 : node2343;
									assign node2343 = (inp[9]) ? node2345 : 1'b1;
										assign node2345 = (inp[7]) ? node2353 : node2346;
											assign node2346 = (inp[0]) ? node2348 : 1'b1;
												assign node2348 = (inp[13]) ? node2350 : 1'b1;
													assign node2350 = (inp[1]) ? 1'b0 : 1'b1;
											assign node2353 = (inp[6]) ? 1'b0 : node2354;
												assign node2354 = (inp[1]) ? node2356 : 1'b1;
													assign node2356 = (inp[10]) ? 1'b0 : 1'b1;
									assign node2360 = (inp[10]) ? node2374 : node2361;
										assign node2361 = (inp[0]) ? node2363 : 1'b1;
											assign node2363 = (inp[1]) ? node2369 : node2364;
												assign node2364 = (inp[9]) ? node2366 : 1'b1;
													assign node2366 = (inp[6]) ? 1'b0 : 1'b1;
												assign node2369 = (inp[13]) ? 1'b0 : node2370;
													assign node2370 = (inp[6]) ? 1'b0 : 1'b1;
										assign node2374 = (inp[1]) ? 1'b0 : node2375;
											assign node2375 = (inp[6]) ? 1'b0 : 1'b1;
							assign node2379 = (inp[6]) ? node2405 : node2380;
								assign node2380 = (inp[13]) ? node2388 : node2381;
									assign node2381 = (inp[10]) ? node2383 : 1'b1;
										assign node2383 = (inp[9]) ? node2385 : 1'b1;
											assign node2385 = (inp[11]) ? 1'b0 : 1'b1;
									assign node2388 = (inp[9]) ? node2396 : node2389;
										assign node2389 = (inp[11]) ? node2391 : 1'b1;
											assign node2391 = (inp[1]) ? 1'b0 : node2392;
												assign node2392 = (inp[14]) ? 1'b0 : 1'b1;
										assign node2396 = (inp[0]) ? 1'b0 : node2397;
											assign node2397 = (inp[11]) ? 1'b0 : node2398;
												assign node2398 = (inp[14]) ? node2400 : 1'b1;
													assign node2400 = (inp[7]) ? 1'b0 : 1'b1;
								assign node2405 = (inp[11]) ? node2433 : node2406;
									assign node2406 = (inp[1]) ? node2418 : node2407;
										assign node2407 = (inp[0]) ? node2411 : node2408;
											assign node2408 = (inp[10]) ? 1'b0 : 1'b1;
											assign node2411 = (inp[9]) ? 1'b0 : node2412;
												assign node2412 = (inp[14]) ? node2414 : 1'b1;
													assign node2414 = (inp[7]) ? 1'b0 : 1'b1;
										assign node2418 = (inp[9]) ? node2426 : node2419;
											assign node2419 = (inp[0]) ? node2421 : 1'b1;
												assign node2421 = (inp[7]) ? 1'b0 : node2422;
													assign node2422 = (inp[13]) ? 1'b0 : 1'b1;
											assign node2426 = (inp[7]) ? node2428 : 1'b0;
												assign node2428 = (inp[14]) ? 1'b0 : node2429;
													assign node2429 = (inp[13]) ? 1'b0 : 1'b1;
									assign node2433 = (inp[14]) ? 1'b0 : node2434;
										assign node2434 = (inp[9]) ? 1'b0 : node2435;
											assign node2435 = (inp[1]) ? node2437 : 1'b1;
												assign node2437 = (inp[0]) ? 1'b0 : node2438;
													assign node2438 = (inp[13]) ? 1'b0 : 1'b1;
						assign node2444 = (inp[1]) ? node2524 : node2445;
							assign node2445 = (inp[13]) ? node2489 : node2446;
								assign node2446 = (inp[11]) ? node2472 : node2447;
									assign node2447 = (inp[6]) ? node2457 : node2448;
										assign node2448 = (inp[2]) ? node2450 : 1'b1;
											assign node2450 = (inp[7]) ? node2452 : 1'b1;
												assign node2452 = (inp[14]) ? node2454 : 1'b1;
													assign node2454 = (inp[9]) ? 1'b0 : 1'b1;
										assign node2457 = (inp[7]) ? node2465 : node2458;
											assign node2458 = (inp[2]) ? node2460 : 1'b1;
												assign node2460 = (inp[9]) ? node2462 : 1'b1;
													assign node2462 = (inp[10]) ? 1'b0 : 1'b1;
											assign node2465 = (inp[9]) ? node2469 : node2466;
												assign node2466 = (inp[2]) ? 1'b0 : 1'b1;
												assign node2469 = (inp[14]) ? 1'b0 : 1'b1;
									assign node2472 = (inp[14]) ? node2482 : node2473;
										assign node2473 = (inp[6]) ? node2475 : 1'b1;
											assign node2475 = (inp[10]) ? node2477 : 1'b1;
												assign node2477 = (inp[2]) ? 1'b0 : node2478;
													assign node2478 = (inp[9]) ? 1'b0 : 1'b1;
										assign node2482 = (inp[6]) ? 1'b0 : node2483;
											assign node2483 = (inp[7]) ? 1'b0 : node2484;
												assign node2484 = (inp[2]) ? 1'b0 : 1'b1;
								assign node2489 = (inp[2]) ? node2511 : node2490;
									assign node2490 = (inp[10]) ? node2498 : node2491;
										assign node2491 = (inp[14]) ? node2493 : 1'b1;
											assign node2493 = (inp[0]) ? node2495 : 1'b1;
												assign node2495 = (inp[6]) ? 1'b0 : 1'b1;
										assign node2498 = (inp[9]) ? node2506 : node2499;
											assign node2499 = (inp[14]) ? node2501 : 1'b1;
												assign node2501 = (inp[11]) ? 1'b0 : node2502;
													assign node2502 = (inp[7]) ? 1'b0 : 1'b1;
											assign node2506 = (inp[0]) ? 1'b0 : node2507;
												assign node2507 = (inp[6]) ? 1'b1 : 1'b0;
									assign node2511 = (inp[6]) ? 1'b0 : node2512;
										assign node2512 = (inp[11]) ? node2518 : node2513;
											assign node2513 = (inp[9]) ? node2515 : 1'b1;
												assign node2515 = (inp[10]) ? 1'b0 : 1'b1;
											assign node2518 = (inp[10]) ? 1'b0 : node2519;
												assign node2519 = (inp[9]) ? 1'b0 : 1'b1;
							assign node2524 = (inp[9]) ? node2560 : node2525;
								assign node2525 = (inp[0]) ? node2541 : node2526;
									assign node2526 = (inp[2]) ? node2536 : node2527;
										assign node2527 = (inp[11]) ? node2529 : 1'b1;
											assign node2529 = (inp[6]) ? 1'b0 : node2530;
												assign node2530 = (inp[14]) ? node2532 : 1'b1;
													assign node2532 = (inp[10]) ? 1'b0 : 1'b1;
										assign node2536 = (inp[10]) ? 1'b0 : node2537;
											assign node2537 = (inp[6]) ? 1'b0 : 1'b1;
									assign node2541 = (inp[11]) ? 1'b0 : node2542;
										assign node2542 = (inp[13]) ? node2554 : node2543;
											assign node2543 = (inp[14]) ? node2549 : node2544;
												assign node2544 = (inp[2]) ? node2546 : 1'b1;
													assign node2546 = (inp[10]) ? 1'b0 : 1'b1;
												assign node2549 = (inp[6]) ? node2551 : 1'b0;
													assign node2551 = (inp[10]) ? 1'b0 : 1'b0;
											assign node2554 = (inp[14]) ? node2556 : 1'b0;
												assign node2556 = (inp[6]) ? 1'b0 : 1'b1;
								assign node2560 = (inp[0]) ? 1'b0 : node2561;
									assign node2561 = (inp[14]) ? 1'b0 : node2562;
										assign node2562 = (inp[10]) ? node2570 : node2563;
											assign node2563 = (inp[11]) ? 1'b0 : node2564;
												assign node2564 = (inp[6]) ? node2566 : 1'b1;
													assign node2566 = (inp[7]) ? 1'b0 : 1'b1;
											assign node2570 = (inp[2]) ? 1'b0 : node2571;
												assign node2571 = (inp[13]) ? 1'b0 : node2572;
													assign node2572 = (inp[6]) ? 1'b0 : 1'b1;
					assign node2579 = (inp[7]) ? node2709 : node2580;
						assign node2580 = (inp[1]) ? node2650 : node2581;
							assign node2581 = (inp[0]) ? node2623 : node2582;
								assign node2582 = (inp[13]) ? node2594 : node2583;
									assign node2583 = (inp[11]) ? node2585 : 1'b1;
										assign node2585 = (inp[8]) ? node2587 : 1'b1;
											assign node2587 = (inp[6]) ? 1'b0 : node2588;
												assign node2588 = (inp[9]) ? node2590 : 1'b1;
													assign node2590 = (inp[2]) ? 1'b0 : 1'b1;
									assign node2594 = (inp[9]) ? node2610 : node2595;
										assign node2595 = (inp[11]) ? node2603 : node2596;
											assign node2596 = (inp[10]) ? node2598 : 1'b1;
												assign node2598 = (inp[14]) ? node2600 : 1'b1;
													assign node2600 = (inp[6]) ? 1'b0 : 1'b1;
											assign node2603 = (inp[6]) ? 1'b0 : node2604;
												assign node2604 = (inp[2]) ? node2606 : 1'b1;
													assign node2606 = (inp[8]) ? 1'b0 : 1'b0;
										assign node2610 = (inp[10]) ? 1'b0 : node2611;
											assign node2611 = (inp[8]) ? node2617 : node2612;
												assign node2612 = (inp[6]) ? node2614 : 1'b1;
													assign node2614 = (inp[14]) ? 1'b0 : 1'b1;
												assign node2617 = (inp[14]) ? 1'b0 : node2618;
													assign node2618 = (inp[11]) ? 1'b0 : 1'b0;
								assign node2623 = (inp[14]) ? node2639 : node2624;
									assign node2624 = (inp[11]) ? node2630 : node2625;
										assign node2625 = (inp[10]) ? node2627 : 1'b1;
											assign node2627 = (inp[6]) ? 1'b0 : 1'b1;
										assign node2630 = (inp[9]) ? 1'b0 : node2631;
											assign node2631 = (inp[13]) ? node2633 : 1'b1;
												assign node2633 = (inp[2]) ? 1'b0 : node2634;
													assign node2634 = (inp[8]) ? 1'b0 : 1'b1;
									assign node2639 = (inp[8]) ? 1'b0 : node2640;
										assign node2640 = (inp[6]) ? 1'b0 : node2641;
											assign node2641 = (inp[11]) ? node2643 : 1'b1;
												assign node2643 = (inp[2]) ? 1'b0 : node2644;
													assign node2644 = (inp[13]) ? 1'b0 : 1'b1;
							assign node2650 = (inp[9]) ? node2682 : node2651;
								assign node2651 = (inp[10]) ? node2671 : node2652;
									assign node2652 = (inp[6]) ? node2658 : node2653;
										assign node2653 = (inp[0]) ? node2655 : 1'b1;
											assign node2655 = (inp[2]) ? 1'b0 : 1'b1;
										assign node2658 = (inp[13]) ? 1'b0 : node2659;
											assign node2659 = (inp[8]) ? node2665 : node2660;
												assign node2660 = (inp[2]) ? node2662 : 1'b1;
													assign node2662 = (inp[11]) ? 1'b0 : 1'b1;
												assign node2665 = (inp[11]) ? 1'b0 : node2666;
													assign node2666 = (inp[14]) ? 1'b0 : 1'b0;
									assign node2671 = (inp[14]) ? 1'b0 : node2672;
										assign node2672 = (inp[0]) ? 1'b0 : node2673;
											assign node2673 = (inp[2]) ? 1'b0 : node2674;
												assign node2674 = (inp[8]) ? node2676 : 1'b1;
													assign node2676 = (inp[6]) ? 1'b0 : 1'b1;
								assign node2682 = (inp[11]) ? 1'b0 : node2683;
									assign node2683 = (inp[2]) ? node2699 : node2684;
										assign node2684 = (inp[8]) ? node2692 : node2685;
											assign node2685 = (inp[6]) ? 1'b0 : node2686;
												assign node2686 = (inp[10]) ? node2688 : 1'b1;
													assign node2688 = (inp[13]) ? 1'b0 : 1'b1;
											assign node2692 = (inp[0]) ? 1'b0 : node2693;
												assign node2693 = (inp[14]) ? 1'b0 : node2694;
													assign node2694 = (inp[13]) ? 1'b0 : 1'b1;
										assign node2699 = (inp[0]) ? 1'b0 : node2700;
											assign node2700 = (inp[8]) ? 1'b0 : node2701;
												assign node2701 = (inp[13]) ? 1'b0 : node2702;
													assign node2702 = (inp[6]) ? 1'b0 : 1'b1;
						assign node2709 = (inp[8]) ? node2747 : node2710;
							assign node2710 = (inp[9]) ? node2734 : node2711;
								assign node2711 = (inp[14]) ? node2725 : node2712;
									assign node2712 = (inp[11]) ? node2718 : node2713;
										assign node2713 = (inp[10]) ? node2715 : 1'b1;
											assign node2715 = (inp[0]) ? 1'b0 : 1'b1;
										assign node2718 = (inp[2]) ? 1'b0 : node2719;
											assign node2719 = (inp[10]) ? node2721 : 1'b1;
												assign node2721 = (inp[1]) ? 1'b0 : 1'b1;
									assign node2725 = (inp[0]) ? 1'b0 : node2726;
										assign node2726 = (inp[13]) ? 1'b0 : node2727;
											assign node2727 = (inp[6]) ? node2729 : 1'b1;
												assign node2729 = (inp[10]) ? 1'b0 : 1'b1;
								assign node2734 = (inp[14]) ? 1'b0 : node2735;
									assign node2735 = (inp[1]) ? 1'b0 : node2736;
										assign node2736 = (inp[6]) ? node2740 : node2737;
											assign node2737 = (inp[2]) ? 1'b0 : 1'b1;
											assign node2740 = (inp[13]) ? 1'b0 : node2741;
												assign node2741 = (inp[10]) ? 1'b0 : 1'b1;
							assign node2747 = (inp[1]) ? 1'b0 : node2748;
								assign node2748 = (inp[10]) ? 1'b0 : node2749;
									assign node2749 = (inp[13]) ? node2755 : node2750;
										assign node2750 = (inp[11]) ? 1'b0 : node2751;
											assign node2751 = (inp[9]) ? 1'b0 : 1'b1;
										assign node2755 = (inp[0]) ? 1'b0 : node2756;
											assign node2756 = (inp[2]) ? 1'b0 : node2757;
												assign node2757 = (inp[9]) ? 1'b0 : node2758;
													assign node2758 = (inp[6]) ? 1'b0 : 1'b1;
			assign node2766 = (inp[10]) ? node3206 : node2767;
				assign node2767 = (inp[0]) ? node3015 : node2768;
					assign node2768 = (inp[11]) ? node2890 : node2769;
						assign node2769 = (inp[2]) ? node2821 : node2770;
							assign node2770 = (inp[9]) ? node2784 : node2771;
								assign node2771 = (inp[13]) ? node2773 : 1'b1;
									assign node2773 = (inp[8]) ? node2775 : 1'b1;
										assign node2775 = (inp[12]) ? node2777 : 1'b1;
											assign node2777 = (inp[5]) ? 1'b0 : node2778;
												assign node2778 = (inp[1]) ? node2780 : 1'b1;
													assign node2780 = (inp[7]) ? 1'b0 : 1'b1;
								assign node2784 = (inp[8]) ? node2796 : node2785;
									assign node2785 = (inp[5]) ? node2787 : 1'b1;
										assign node2787 = (inp[14]) ? node2793 : node2788;
											assign node2788 = (inp[6]) ? node2790 : 1'b1;
												assign node2790 = (inp[12]) ? 1'b0 : 1'b1;
											assign node2793 = (inp[6]) ? 1'b1 : 1'b0;
									assign node2796 = (inp[5]) ? node2808 : node2797;
										assign node2797 = (inp[12]) ? node2805 : node2798;
											assign node2798 = (inp[14]) ? node2800 : 1'b1;
												assign node2800 = (inp[7]) ? node2802 : 1'b1;
													assign node2802 = (inp[1]) ? 1'b0 : 1'b1;
											assign node2805 = (inp[13]) ? 1'b0 : 1'b1;
										assign node2808 = (inp[6]) ? node2814 : node2809;
											assign node2809 = (inp[13]) ? node2811 : 1'b1;
												assign node2811 = (inp[1]) ? 1'b0 : 1'b1;
											assign node2814 = (inp[12]) ? 1'b0 : node2815;
												assign node2815 = (inp[13]) ? 1'b0 : node2816;
													assign node2816 = (inp[1]) ? 1'b0 : 1'b1;
							assign node2821 = (inp[13]) ? node2847 : node2822;
								assign node2822 = (inp[9]) ? node2832 : node2823;
									assign node2823 = (inp[1]) ? node2825 : 1'b1;
										assign node2825 = (inp[5]) ? node2827 : 1'b1;
											assign node2827 = (inp[8]) ? node2829 : 1'b1;
												assign node2829 = (inp[14]) ? 1'b0 : 1'b1;
									assign node2832 = (inp[1]) ? node2842 : node2833;
										assign node2833 = (inp[6]) ? node2835 : 1'b1;
											assign node2835 = (inp[7]) ? 1'b0 : node2836;
												assign node2836 = (inp[8]) ? node2838 : 1'b1;
													assign node2838 = (inp[14]) ? 1'b0 : 1'b1;
										assign node2842 = (inp[8]) ? 1'b0 : node2843;
											assign node2843 = (inp[6]) ? 1'b0 : 1'b1;
								assign node2847 = (inp[6]) ? node2873 : node2848;
									assign node2848 = (inp[9]) ? node2864 : node2849;
										assign node2849 = (inp[5]) ? node2857 : node2850;
											assign node2850 = (inp[14]) ? node2852 : 1'b1;
												assign node2852 = (inp[7]) ? node2854 : 1'b1;
													assign node2854 = (inp[1]) ? 1'b0 : 1'b1;
											assign node2857 = (inp[12]) ? 1'b0 : node2858;
												assign node2858 = (inp[1]) ? node2860 : 1'b1;
													assign node2860 = (inp[8]) ? 1'b0 : 1'b1;
										assign node2864 = (inp[14]) ? 1'b0 : node2865;
											assign node2865 = (inp[5]) ? node2867 : 1'b0;
												assign node2867 = (inp[7]) ? node2869 : 1'b1;
													assign node2869 = (inp[8]) ? 1'b0 : 1'b1;
									assign node2873 = (inp[1]) ? 1'b0 : node2874;
										assign node2874 = (inp[5]) ? node2882 : node2875;
											assign node2875 = (inp[8]) ? node2877 : 1'b1;
												assign node2877 = (inp[14]) ? 1'b0 : node2878;
													assign node2878 = (inp[12]) ? 1'b0 : 1'b1;
											assign node2882 = (inp[8]) ? 1'b0 : node2883;
												assign node2883 = (inp[7]) ? 1'b0 : node2884;
													assign node2884 = (inp[12]) ? 1'b0 : 1'b1;
						assign node2890 = (inp[7]) ? node2964 : node2891;
							assign node2891 = (inp[9]) ? node2929 : node2892;
								assign node2892 = (inp[6]) ? node2908 : node2893;
									assign node2893 = (inp[2]) ? node2895 : 1'b1;
										assign node2895 = (inp[5]) ? node2901 : node2896;
											assign node2896 = (inp[13]) ? node2898 : 1'b1;
												assign node2898 = (inp[8]) ? 1'b0 : 1'b1;
											assign node2901 = (inp[8]) ? 1'b0 : node2902;
												assign node2902 = (inp[1]) ? node2904 : 1'b1;
													assign node2904 = (inp[14]) ? 1'b0 : 1'b1;
									assign node2908 = (inp[1]) ? node2920 : node2909;
										assign node2909 = (inp[5]) ? node2911 : 1'b1;
											assign node2911 = (inp[2]) ? node2917 : node2912;
												assign node2912 = (inp[14]) ? node2914 : 1'b1;
													assign node2914 = (inp[8]) ? 1'b0 : 1'b1;
												assign node2917 = (inp[13]) ? 1'b0 : 1'b1;
										assign node2920 = (inp[5]) ? 1'b0 : node2921;
											assign node2921 = (inp[12]) ? 1'b0 : node2922;
												assign node2922 = (inp[2]) ? node2924 : 1'b1;
													assign node2924 = (inp[13]) ? 1'b0 : 1'b1;
								assign node2929 = (inp[14]) ? node2949 : node2930;
									assign node2930 = (inp[1]) ? node2940 : node2931;
										assign node2931 = (inp[6]) ? node2933 : 1'b1;
											assign node2933 = (inp[5]) ? 1'b0 : node2934;
												assign node2934 = (inp[13]) ? node2936 : 1'b1;
													assign node2936 = (inp[8]) ? 1'b0 : 1'b1;
										assign node2940 = (inp[8]) ? 1'b0 : node2941;
											assign node2941 = (inp[12]) ? node2943 : 1'b1;
												assign node2943 = (inp[5]) ? 1'b0 : node2944;
													assign node2944 = (inp[13]) ? 1'b0 : 1'b1;
									assign node2949 = (inp[8]) ? 1'b0 : node2950;
										assign node2950 = (inp[13]) ? node2958 : node2951;
											assign node2951 = (inp[5]) ? node2953 : 1'b1;
												assign node2953 = (inp[6]) ? 1'b0 : node2954;
													assign node2954 = (inp[12]) ? 1'b0 : 1'b1;
											assign node2958 = (inp[12]) ? 1'b0 : node2959;
												assign node2959 = (inp[6]) ? 1'b0 : 1'b1;
							assign node2964 = (inp[14]) ? node3002 : node2965;
								assign node2965 = (inp[1]) ? node2991 : node2966;
									assign node2966 = (inp[5]) ? node2976 : node2967;
										assign node2967 = (inp[12]) ? node2969 : 1'b1;
											assign node2969 = (inp[2]) ? node2971 : 1'b1;
												assign node2971 = (inp[9]) ? 1'b0 : node2972;
													assign node2972 = (inp[13]) ? 1'b0 : 1'b1;
										assign node2976 = (inp[6]) ? node2984 : node2977;
											assign node2977 = (inp[2]) ? node2979 : 1'b1;
												assign node2979 = (inp[13]) ? 1'b0 : node2980;
													assign node2980 = (inp[9]) ? 1'b0 : 1'b1;
											assign node2984 = (inp[12]) ? 1'b0 : node2985;
												assign node2985 = (inp[2]) ? 1'b0 : node2986;
													assign node2986 = (inp[9]) ? 1'b0 : 1'b1;
									assign node2991 = (inp[13]) ? 1'b0 : node2992;
										assign node2992 = (inp[9]) ? 1'b0 : node2993;
											assign node2993 = (inp[12]) ? node2995 : 1'b1;
												assign node2995 = (inp[2]) ? 1'b0 : node2996;
													assign node2996 = (inp[6]) ? 1'b0 : 1'b1;
								assign node3002 = (inp[5]) ? 1'b0 : node3003;
									assign node3003 = (inp[1]) ? 1'b0 : node3004;
										assign node3004 = (inp[12]) ? 1'b0 : node3005;
											assign node3005 = (inp[8]) ? 1'b0 : node3006;
												assign node3006 = (inp[9]) ? node3008 : 1'b1;
													assign node3008 = (inp[13]) ? 1'b0 : 1'b1;
					assign node3015 = (inp[8]) ? node3121 : node3016;
						assign node3016 = (inp[7]) ? node3074 : node3017;
							assign node3017 = (inp[2]) ? node3043 : node3018;
								assign node3018 = (inp[1]) ? node3028 : node3019;
									assign node3019 = (inp[6]) ? node3021 : 1'b1;
										assign node3021 = (inp[5]) ? node3023 : 1'b1;
											assign node3023 = (inp[9]) ? 1'b0 : node3024;
												assign node3024 = (inp[13]) ? 1'b0 : 1'b1;
									assign node3028 = (inp[9]) ? node3038 : node3029;
										assign node3029 = (inp[5]) ? node3031 : 1'b1;
											assign node3031 = (inp[14]) ? node3033 : 1'b1;
												assign node3033 = (inp[11]) ? 1'b0 : node3034;
													assign node3034 = (inp[13]) ? 1'b0 : 1'b1;
										assign node3038 = (inp[11]) ? 1'b0 : node3039;
											assign node3039 = (inp[12]) ? 1'b0 : 1'b1;
								assign node3043 = (inp[11]) ? node3063 : node3044;
									assign node3044 = (inp[5]) ? node3050 : node3045;
										assign node3045 = (inp[14]) ? node3047 : 1'b1;
											assign node3047 = (inp[12]) ? 1'b0 : 1'b1;
										assign node3050 = (inp[6]) ? 1'b0 : node3051;
											assign node3051 = (inp[12]) ? node3057 : node3052;
												assign node3052 = (inp[14]) ? node3054 : 1'b1;
													assign node3054 = (inp[9]) ? 1'b0 : 1'b1;
												assign node3057 = (inp[9]) ? 1'b0 : node3058;
													assign node3058 = (inp[1]) ? 1'b0 : 1'b1;
									assign node3063 = (inp[12]) ? 1'b0 : node3064;
										assign node3064 = (inp[13]) ? 1'b0 : node3065;
											assign node3065 = (inp[9]) ? 1'b0 : node3066;
												assign node3066 = (inp[1]) ? node3068 : 1'b1;
													assign node3068 = (inp[6]) ? 1'b0 : 1'b1;
							assign node3074 = (inp[13]) ? node3102 : node3075;
								assign node3075 = (inp[1]) ? node3087 : node3076;
									assign node3076 = (inp[6]) ? node3082 : node3077;
										assign node3077 = (inp[2]) ? node3079 : 1'b1;
											assign node3079 = (inp[11]) ? 1'b0 : 1'b1;
										assign node3082 = (inp[14]) ? 1'b0 : node3083;
											assign node3083 = (inp[11]) ? 1'b0 : 1'b1;
									assign node3087 = (inp[5]) ? 1'b0 : node3088;
										assign node3088 = (inp[11]) ? node3096 : node3089;
											assign node3089 = (inp[14]) ? node3091 : 1'b1;
												assign node3091 = (inp[12]) ? 1'b0 : node3092;
													assign node3092 = (inp[2]) ? 1'b0 : 1'b1;
											assign node3096 = (inp[2]) ? 1'b0 : node3097;
												assign node3097 = (inp[12]) ? 1'b0 : 1'b1;
								assign node3102 = (inp[12]) ? 1'b0 : node3103;
									assign node3103 = (inp[5]) ? node3113 : node3104;
										assign node3104 = (inp[11]) ? 1'b0 : node3105;
											assign node3105 = (inp[1]) ? node3107 : 1'b1;
												assign node3107 = (inp[6]) ? 1'b0 : node3108;
													assign node3108 = (inp[2]) ? 1'b0 : 1'b1;
										assign node3113 = (inp[1]) ? 1'b0 : node3114;
											assign node3114 = (inp[2]) ? 1'b0 : node3115;
												assign node3115 = (inp[6]) ? 1'b0 : 1'b1;
						assign node3121 = (inp[5]) ? node3181 : node3122;
							assign node3122 = (inp[13]) ? node3162 : node3123;
								assign node3123 = (inp[2]) ? node3141 : node3124;
									assign node3124 = (inp[9]) ? node3138 : node3125;
										assign node3125 = (inp[11]) ? node3127 : 1'b1;
											assign node3127 = (inp[12]) ? node3133 : node3128;
												assign node3128 = (inp[7]) ? node3130 : 1'b1;
													assign node3130 = (inp[1]) ? 1'b0 : 1'b1;
												assign node3133 = (inp[1]) ? 1'b0 : node3134;
													assign node3134 = (inp[7]) ? 1'b0 : 1'b1;
										assign node3138 = (inp[7]) ? 1'b0 : 1'b1;
									assign node3141 = (inp[7]) ? 1'b0 : node3142;
										assign node3142 = (inp[6]) ? node3154 : node3143;
											assign node3143 = (inp[11]) ? node3149 : node3144;
												assign node3144 = (inp[14]) ? node3146 : 1'b1;
													assign node3146 = (inp[1]) ? 1'b0 : 1'b1;
												assign node3149 = (inp[12]) ? 1'b0 : node3150;
													assign node3150 = (inp[9]) ? 1'b0 : 1'b1;
											assign node3154 = (inp[11]) ? node3156 : 1'b0;
												assign node3156 = (inp[12]) ? 1'b0 : node3157;
													assign node3157 = (inp[9]) ? 1'b0 : 1'b1;
								assign node3162 = (inp[14]) ? 1'b0 : node3163;
									assign node3163 = (inp[6]) ? 1'b0 : node3164;
										assign node3164 = (inp[1]) ? node3172 : node3165;
											assign node3165 = (inp[9]) ? node3167 : 1'b1;
												assign node3167 = (inp[2]) ? 1'b0 : node3168;
													assign node3168 = (inp[11]) ? 1'b0 : 1'b1;
											assign node3172 = (inp[2]) ? 1'b0 : node3173;
												assign node3173 = (inp[12]) ? 1'b0 : node3174;
													assign node3174 = (inp[11]) ? 1'b0 : 1'b1;
							assign node3181 = (inp[13]) ? 1'b0 : node3182;
								assign node3182 = (inp[11]) ? 1'b0 : node3183;
									assign node3183 = (inp[1]) ? node3197 : node3184;
										assign node3184 = (inp[9]) ? node3192 : node3185;
											assign node3185 = (inp[14]) ? node3187 : 1'b1;
												assign node3187 = (inp[2]) ? node3189 : 1'b0;
													assign node3189 = (inp[7]) ? 1'b0 : 1'b1;
											assign node3192 = (inp[12]) ? 1'b0 : node3193;
												assign node3193 = (inp[14]) ? 1'b0 : 1'b1;
										assign node3197 = (inp[2]) ? 1'b0 : node3198;
											assign node3198 = (inp[6]) ? 1'b0 : node3199;
												assign node3199 = (inp[12]) ? 1'b0 : 1'b1;
				assign node3206 = (inp[1]) ? node3440 : node3207;
					assign node3207 = (inp[8]) ? node3357 : node3208;
						assign node3208 = (inp[11]) ? node3294 : node3209;
							assign node3209 = (inp[9]) ? node3253 : node3210;
								assign node3210 = (inp[13]) ? node3228 : node3211;
									assign node3211 = (inp[0]) ? node3213 : 1'b1;
										assign node3213 = (inp[6]) ? node3221 : node3214;
											assign node3214 = (inp[12]) ? node3216 : 1'b1;
												assign node3216 = (inp[14]) ? node3218 : 1'b1;
													assign node3218 = (inp[7]) ? 1'b0 : 1'b1;
											assign node3221 = (inp[2]) ? 1'b0 : node3222;
												assign node3222 = (inp[7]) ? node3224 : 1'b1;
													assign node3224 = (inp[5]) ? 1'b0 : 1'b1;
									assign node3228 = (inp[5]) ? node3240 : node3229;
										assign node3229 = (inp[6]) ? node3235 : node3230;
											assign node3230 = (inp[12]) ? node3232 : 1'b1;
												assign node3232 = (inp[7]) ? 1'b0 : 1'b1;
											assign node3235 = (inp[0]) ? 1'b0 : node3236;
												assign node3236 = (inp[14]) ? 1'b0 : 1'b1;
										assign node3240 = (inp[14]) ? 1'b0 : node3241;
											assign node3241 = (inp[7]) ? node3247 : node3242;
												assign node3242 = (inp[2]) ? 1'b0 : node3243;
													assign node3243 = (inp[12]) ? 1'b0 : 1'b1;
												assign node3247 = (inp[0]) ? 1'b0 : node3248;
													assign node3248 = (inp[6]) ? 1'b0 : 1'b1;
								assign node3253 = (inp[7]) ? node3279 : node3254;
									assign node3254 = (inp[12]) ? node3264 : node3255;
										assign node3255 = (inp[14]) ? node3257 : 1'b1;
											assign node3257 = (inp[0]) ? 1'b0 : node3258;
												assign node3258 = (inp[2]) ? node3260 : 1'b1;
													assign node3260 = (inp[6]) ? 1'b0 : 1'b1;
										assign node3264 = (inp[2]) ? node3272 : node3265;
											assign node3265 = (inp[14]) ? node3267 : 1'b1;
												assign node3267 = (inp[13]) ? 1'b0 : node3268;
													assign node3268 = (inp[0]) ? 1'b0 : 1'b1;
											assign node3272 = (inp[13]) ? 1'b0 : node3273;
												assign node3273 = (inp[5]) ? 1'b0 : node3274;
													assign node3274 = (inp[6]) ? 1'b0 : 1'b1;
									assign node3279 = (inp[0]) ? 1'b0 : node3280;
										assign node3280 = (inp[2]) ? 1'b0 : node3281;
											assign node3281 = (inp[13]) ? node3287 : node3282;
												assign node3282 = (inp[5]) ? node3284 : 1'b1;
													assign node3284 = (inp[12]) ? 1'b0 : 1'b1;
												assign node3287 = (inp[6]) ? 1'b0 : node3288;
													assign node3288 = (inp[5]) ? 1'b0 : 1'b1;
							assign node3294 = (inp[7]) ? node3340 : node3295;
								assign node3295 = (inp[5]) ? node3329 : node3296;
									assign node3296 = (inp[9]) ? node3312 : node3297;
										assign node3297 = (inp[13]) ? node3305 : node3298;
											assign node3298 = (inp[2]) ? node3300 : 1'b1;
												assign node3300 = (inp[0]) ? node3302 : 1'b1;
													assign node3302 = (inp[14]) ? 1'b0 : 1'b1;
											assign node3305 = (inp[12]) ? 1'b0 : node3306;
												assign node3306 = (inp[14]) ? node3308 : 1'b1;
													assign node3308 = (inp[2]) ? 1'b0 : 1'b1;
										assign node3312 = (inp[14]) ? node3324 : node3313;
											assign node3313 = (inp[13]) ? node3319 : node3314;
												assign node3314 = (inp[12]) ? node3316 : 1'b1;
													assign node3316 = (inp[6]) ? 1'b0 : 1'b1;
												assign node3319 = (inp[0]) ? 1'b0 : node3320;
													assign node3320 = (inp[6]) ? 1'b0 : 1'b1;
											assign node3324 = (inp[12]) ? 1'b0 : node3325;
												assign node3325 = (inp[0]) ? 1'b0 : 1'b1;
									assign node3329 = (inp[0]) ? 1'b0 : node3330;
										assign node3330 = (inp[12]) ? 1'b0 : node3331;
											assign node3331 = (inp[2]) ? node3333 : 1'b1;
												assign node3333 = (inp[9]) ? 1'b0 : node3334;
													assign node3334 = (inp[6]) ? 1'b0 : 1'b1;
								assign node3340 = (inp[0]) ? 1'b0 : node3341;
									assign node3341 = (inp[13]) ? 1'b0 : node3342;
										assign node3342 = (inp[14]) ? node3348 : node3343;
											assign node3343 = (inp[12]) ? node3345 : 1'b1;
												assign node3345 = (inp[6]) ? 1'b0 : 1'b1;
											assign node3348 = (inp[12]) ? 1'b0 : node3349;
												assign node3349 = (inp[9]) ? 1'b0 : node3350;
													assign node3350 = (inp[5]) ? 1'b0 : 1'b1;
						assign node3357 = (inp[5]) ? node3419 : node3358;
							assign node3358 = (inp[12]) ? node3400 : node3359;
								assign node3359 = (inp[2]) ? node3383 : node3360;
									assign node3360 = (inp[0]) ? node3368 : node3361;
										assign node3361 = (inp[13]) ? node3363 : 1'b1;
											assign node3363 = (inp[9]) ? 1'b0 : node3364;
												assign node3364 = (inp[14]) ? 1'b0 : 1'b1;
										assign node3368 = (inp[6]) ? node3376 : node3369;
											assign node3369 = (inp[13]) ? node3371 : 1'b1;
												assign node3371 = (inp[7]) ? 1'b0 : node3372;
													assign node3372 = (inp[14]) ? 1'b0 : 1'b1;
											assign node3376 = (inp[9]) ? 1'b0 : node3377;
												assign node3377 = (inp[14]) ? 1'b0 : node3378;
													assign node3378 = (inp[7]) ? 1'b0 : 1'b1;
									assign node3383 = (inp[0]) ? 1'b0 : node3384;
										assign node3384 = (inp[11]) ? node3392 : node3385;
											assign node3385 = (inp[7]) ? node3387 : 1'b1;
												assign node3387 = (inp[6]) ? 1'b0 : node3388;
													assign node3388 = (inp[9]) ? 1'b0 : 1'b1;
											assign node3392 = (inp[6]) ? 1'b0 : node3393;
												assign node3393 = (inp[7]) ? 1'b0 : node3394;
													assign node3394 = (inp[9]) ? 1'b0 : 1'b1;
								assign node3400 = (inp[7]) ? 1'b0 : node3401;
									assign node3401 = (inp[14]) ? node3409 : node3402;
										assign node3402 = (inp[0]) ? node3404 : 1'b1;
											assign node3404 = (inp[13]) ? 1'b0 : node3405;
												assign node3405 = (inp[6]) ? 1'b0 : 1'b1;
										assign node3409 = (inp[9]) ? 1'b0 : node3410;
											assign node3410 = (inp[11]) ? 1'b0 : node3411;
												assign node3411 = (inp[0]) ? 1'b0 : node3412;
													assign node3412 = (inp[2]) ? 1'b0 : 1'b1;
							assign node3419 = (inp[12]) ? 1'b0 : node3420;
								assign node3420 = (inp[11]) ? 1'b0 : node3421;
									assign node3421 = (inp[14]) ? node3431 : node3422;
										assign node3422 = (inp[7]) ? node3424 : 1'b1;
											assign node3424 = (inp[9]) ? 1'b0 : node3425;
												assign node3425 = (inp[2]) ? 1'b0 : node3426;
													assign node3426 = (inp[13]) ? 1'b0 : 1'b1;
										assign node3431 = (inp[2]) ? 1'b0 : node3432;
											assign node3432 = (inp[9]) ? 1'b0 : node3433;
												assign node3433 = (inp[6]) ? 1'b0 : 1'b1;
					assign node3440 = (inp[5]) ? node3512 : node3441;
						assign node3441 = (inp[14]) ? node3487 : node3442;
							assign node3442 = (inp[0]) ? node3474 : node3443;
								assign node3443 = (inp[11]) ? node3463 : node3444;
									assign node3444 = (inp[7]) ? node3454 : node3445;
										assign node3445 = (inp[2]) ? node3447 : 1'b1;
											assign node3447 = (inp[9]) ? 1'b0 : node3448;
												assign node3448 = (inp[12]) ? node3450 : 1'b1;
													assign node3450 = (inp[6]) ? 1'b0 : 1'b1;
										assign node3454 = (inp[12]) ? 1'b0 : node3455;
											assign node3455 = (inp[8]) ? node3457 : 1'b1;
												assign node3457 = (inp[6]) ? 1'b0 : node3458;
													assign node3458 = (inp[2]) ? 1'b0 : 1'b1;
									assign node3463 = (inp[9]) ? 1'b0 : node3464;
										assign node3464 = (inp[6]) ? 1'b0 : node3465;
											assign node3465 = (inp[2]) ? node3467 : 1'b1;
												assign node3467 = (inp[8]) ? 1'b0 : node3468;
													assign node3468 = (inp[7]) ? 1'b0 : 1'b1;
								assign node3474 = (inp[13]) ? 1'b0 : node3475;
									assign node3475 = (inp[2]) ? 1'b0 : node3476;
										assign node3476 = (inp[7]) ? 1'b0 : node3477;
											assign node3477 = (inp[6]) ? node3479 : 1'b1;
												assign node3479 = (inp[9]) ? 1'b0 : node3480;
													assign node3480 = (inp[12]) ? 1'b0 : 1'b1;
							assign node3487 = (inp[7]) ? 1'b0 : node3488;
								assign node3488 = (inp[13]) ? node3502 : node3489;
									assign node3489 = (inp[11]) ? node3495 : node3490;
										assign node3490 = (inp[12]) ? 1'b0 : node3491;
											assign node3491 = (inp[2]) ? 1'b0 : 1'b1;
										assign node3495 = (inp[8]) ? 1'b0 : node3496;
											assign node3496 = (inp[6]) ? 1'b0 : node3497;
												assign node3497 = (inp[9]) ? 1'b0 : 1'b1;
									assign node3502 = (inp[0]) ? 1'b0 : node3503;
										assign node3503 = (inp[9]) ? 1'b0 : node3504;
											assign node3504 = (inp[12]) ? 1'b0 : node3505;
												assign node3505 = (inp[6]) ? 1'b0 : 1'b1;
						assign node3512 = (inp[13]) ? 1'b0 : node3513;
							assign node3513 = (inp[0]) ? node3539 : node3514;
								assign node3514 = (inp[9]) ? node3530 : node3515;
									assign node3515 = (inp[12]) ? node3523 : node3516;
										assign node3516 = (inp[8]) ? 1'b0 : node3517;
											assign node3517 = (inp[6]) ? node3519 : 1'b1;
												assign node3519 = (inp[14]) ? 1'b0 : 1'b1;
										assign node3523 = (inp[14]) ? 1'b0 : node3524;
											assign node3524 = (inp[7]) ? 1'b0 : node3525;
												assign node3525 = (inp[6]) ? 1'b0 : 1'b1;
									assign node3530 = (inp[2]) ? 1'b0 : node3531;
										assign node3531 = (inp[11]) ? 1'b0 : node3532;
											assign node3532 = (inp[8]) ? 1'b0 : node3533;
												assign node3533 = (inp[7]) ? 1'b0 : 1'b1;
								assign node3539 = (inp[6]) ? 1'b0 : node3540;
									assign node3540 = (inp[9]) ? 1'b0 : node3541;
										assign node3541 = (inp[7]) ? 1'b0 : node3542;
											assign node3542 = (inp[11]) ? 1'b0 : node3543;
												assign node3543 = (inp[8]) ? 1'b0 : 1'b1;

endmodule