module dtc_split75_bm45 (
	input  wire [16-1:0] inp,
	output wire [46-1:0] outp
);

	wire [46-1:0] node1;
	wire [46-1:0] node2;
	wire [46-1:0] node5;
	wire [46-1:0] node6;
	wire [46-1:0] node8;
	wire [46-1:0] node10;
	wire [46-1:0] node11;
	wire [46-1:0] node13;
	wire [46-1:0] node15;
	wire [46-1:0] node16;
	wire [46-1:0] node18;
	wire [46-1:0] node19;
	wire [46-1:0] node24;
	wire [46-1:0] node26;
	wire [46-1:0] node27;
	wire [46-1:0] node28;
	wire [46-1:0] node30;
	wire [46-1:0] node32;
	wire [46-1:0] node34;
	wire [46-1:0] node36;
	wire [46-1:0] node40;
	wire [46-1:0] node41;
	wire [46-1:0] node43;
	wire [46-1:0] node45;
	wire [46-1:0] node47;
	wire [46-1:0] node49;
	wire [46-1:0] node52;
	wire [46-1:0] node54;
	wire [46-1:0] node56;
	wire [46-1:0] node58;
	wire [46-1:0] node60;
	wire [46-1:0] node63;
	wire [46-1:0] node64;
	wire [46-1:0] node65;
	wire [46-1:0] node66;
	wire [46-1:0] node67;
	wire [46-1:0] node71;
	wire [46-1:0] node72;
	wire [46-1:0] node74;
	wire [46-1:0] node76;
	wire [46-1:0] node78;
	wire [46-1:0] node79;
	wire [46-1:0] node80;
	wire [46-1:0] node82;
	wire [46-1:0] node85;
	wire [46-1:0] node86;
	wire [46-1:0] node90;
	wire [46-1:0] node91;
	wire [46-1:0] node93;
	wire [46-1:0] node96;
	wire [46-1:0] node97;
	wire [46-1:0] node100;
	wire [46-1:0] node104;
	wire [46-1:0] node105;
	wire [46-1:0] node106;
	wire [46-1:0] node110;
	wire [46-1:0] node111;
	wire [46-1:0] node114;
	wire [46-1:0] node117;
	wire [46-1:0] node118;
	wire [46-1:0] node119;
	wire [46-1:0] node120;
	wire [46-1:0] node123;
	wire [46-1:0] node125;
	wire [46-1:0] node127;
	wire [46-1:0] node128;
	wire [46-1:0] node130;
	wire [46-1:0] node132;
	wire [46-1:0] node134;
	wire [46-1:0] node137;
	wire [46-1:0] node138;
	wire [46-1:0] node139;
	wire [46-1:0] node140;
	wire [46-1:0] node143;
	wire [46-1:0] node146;
	wire [46-1:0] node147;
	wire [46-1:0] node151;
	wire [46-1:0] node152;
	wire [46-1:0] node154;
	wire [46-1:0] node157;
	wire [46-1:0] node158;
	wire [46-1:0] node161;
	wire [46-1:0] node164;
	wire [46-1:0] node165;
	wire [46-1:0] node167;
	wire [46-1:0] node169;
	wire [46-1:0] node171;
	wire [46-1:0] node173;
	wire [46-1:0] node174;
	wire [46-1:0] node175;
	wire [46-1:0] node178;
	wire [46-1:0] node181;
	wire [46-1:0] node182;
	wire [46-1:0] node186;
	wire [46-1:0] node188;
	wire [46-1:0] node190;
	wire [46-1:0] node192;
	wire [46-1:0] node193;
	wire [46-1:0] node195;
	wire [46-1:0] node197;
	wire [46-1:0] node200;
	wire [46-1:0] node201;
	wire [46-1:0] node202;
	wire [46-1:0] node205;
	wire [46-1:0] node208;
	wire [46-1:0] node209;
	wire [46-1:0] node213;
	wire [46-1:0] node215;
	wire [46-1:0] node217;
	wire [46-1:0] node219;
	wire [46-1:0] node220;
	wire [46-1:0] node222;
	wire [46-1:0] node224;
	wire [46-1:0] node226;
	wire [46-1:0] node228;
	wire [46-1:0] node231;
	wire [46-1:0] node232;
	wire [46-1:0] node234;
	wire [46-1:0] node236;
	wire [46-1:0] node237;
	wire [46-1:0] node240;
	wire [46-1:0] node243;
	wire [46-1:0] node244;
	wire [46-1:0] node245;
	wire [46-1:0] node246;
	wire [46-1:0] node249;
	wire [46-1:0] node253;
	wire [46-1:0] node254;
	wire [46-1:0] node256;
	wire [46-1:0] node259;
	wire [46-1:0] node260;
	wire [46-1:0] node264;
	wire [46-1:0] node265;
	wire [46-1:0] node266;
	wire [46-1:0] node269;
	wire [46-1:0] node270;
	wire [46-1:0] node271;
	wire [46-1:0] node272;
	wire [46-1:0] node273;
	wire [46-1:0] node276;
	wire [46-1:0] node279;
	wire [46-1:0] node280;
	wire [46-1:0] node283;
	wire [46-1:0] node286;
	wire [46-1:0] node287;
	wire [46-1:0] node288;
	wire [46-1:0] node291;
	wire [46-1:0] node294;
	wire [46-1:0] node295;
	wire [46-1:0] node298;
	wire [46-1:0] node301;
	wire [46-1:0] node302;
	wire [46-1:0] node303;
	wire [46-1:0] node304;
	wire [46-1:0] node307;
	wire [46-1:0] node310;
	wire [46-1:0] node311;
	wire [46-1:0] node314;
	wire [46-1:0] node317;
	wire [46-1:0] node318;
	wire [46-1:0] node319;
	wire [46-1:0] node322;
	wire [46-1:0] node325;
	wire [46-1:0] node326;
	wire [46-1:0] node329;
	wire [46-1:0] node332;
	wire [46-1:0] node333;
	wire [46-1:0] node336;
	wire [46-1:0] node338;
	wire [46-1:0] node339;
	wire [46-1:0] node340;
	wire [46-1:0] node341;
	wire [46-1:0] node342;
	wire [46-1:0] node343;
	wire [46-1:0] node344;
	wire [46-1:0] node345;
	wire [46-1:0] node346;
	wire [46-1:0] node347;
	wire [46-1:0] node350;
	wire [46-1:0] node353;
	wire [46-1:0] node354;
	wire [46-1:0] node357;
	wire [46-1:0] node360;
	wire [46-1:0] node361;
	wire [46-1:0] node362;
	wire [46-1:0] node365;
	wire [46-1:0] node368;
	wire [46-1:0] node369;
	wire [46-1:0] node372;
	wire [46-1:0] node375;
	wire [46-1:0] node376;
	wire [46-1:0] node377;
	wire [46-1:0] node378;
	wire [46-1:0] node381;
	wire [46-1:0] node384;
	wire [46-1:0] node385;
	wire [46-1:0] node388;
	wire [46-1:0] node391;
	wire [46-1:0] node392;
	wire [46-1:0] node393;
	wire [46-1:0] node396;
	wire [46-1:0] node399;
	wire [46-1:0] node400;
	wire [46-1:0] node403;
	wire [46-1:0] node406;
	wire [46-1:0] node407;
	wire [46-1:0] node408;
	wire [46-1:0] node409;
	wire [46-1:0] node410;
	wire [46-1:0] node413;
	wire [46-1:0] node416;
	wire [46-1:0] node417;
	wire [46-1:0] node420;
	wire [46-1:0] node423;
	wire [46-1:0] node424;
	wire [46-1:0] node425;
	wire [46-1:0] node428;
	wire [46-1:0] node431;
	wire [46-1:0] node432;
	wire [46-1:0] node435;
	wire [46-1:0] node438;
	wire [46-1:0] node439;
	wire [46-1:0] node440;
	wire [46-1:0] node441;
	wire [46-1:0] node444;
	wire [46-1:0] node447;
	wire [46-1:0] node448;
	wire [46-1:0] node451;
	wire [46-1:0] node454;
	wire [46-1:0] node455;
	wire [46-1:0] node456;
	wire [46-1:0] node459;
	wire [46-1:0] node462;
	wire [46-1:0] node463;
	wire [46-1:0] node466;
	wire [46-1:0] node469;
	wire [46-1:0] node470;
	wire [46-1:0] node471;
	wire [46-1:0] node472;
	wire [46-1:0] node473;
	wire [46-1:0] node474;
	wire [46-1:0] node477;
	wire [46-1:0] node480;
	wire [46-1:0] node481;
	wire [46-1:0] node484;
	wire [46-1:0] node487;
	wire [46-1:0] node488;
	wire [46-1:0] node489;
	wire [46-1:0] node492;
	wire [46-1:0] node495;
	wire [46-1:0] node496;
	wire [46-1:0] node499;
	wire [46-1:0] node502;
	wire [46-1:0] node503;
	wire [46-1:0] node504;
	wire [46-1:0] node505;
	wire [46-1:0] node508;
	wire [46-1:0] node511;
	wire [46-1:0] node512;
	wire [46-1:0] node515;
	wire [46-1:0] node518;
	wire [46-1:0] node519;
	wire [46-1:0] node520;
	wire [46-1:0] node523;
	wire [46-1:0] node526;
	wire [46-1:0] node527;
	wire [46-1:0] node530;
	wire [46-1:0] node533;
	wire [46-1:0] node534;
	wire [46-1:0] node535;
	wire [46-1:0] node536;
	wire [46-1:0] node537;
	wire [46-1:0] node540;
	wire [46-1:0] node543;
	wire [46-1:0] node544;
	wire [46-1:0] node547;
	wire [46-1:0] node550;
	wire [46-1:0] node551;
	wire [46-1:0] node552;
	wire [46-1:0] node555;
	wire [46-1:0] node558;
	wire [46-1:0] node559;
	wire [46-1:0] node562;
	wire [46-1:0] node565;
	wire [46-1:0] node566;
	wire [46-1:0] node567;
	wire [46-1:0] node568;
	wire [46-1:0] node571;
	wire [46-1:0] node574;
	wire [46-1:0] node575;
	wire [46-1:0] node578;
	wire [46-1:0] node581;
	wire [46-1:0] node582;
	wire [46-1:0] node583;
	wire [46-1:0] node586;
	wire [46-1:0] node589;
	wire [46-1:0] node590;
	wire [46-1:0] node593;
	wire [46-1:0] node596;
	wire [46-1:0] node597;
	wire [46-1:0] node599;
	wire [46-1:0] node601;
	wire [46-1:0] node602;
	wire [46-1:0] node604;
	wire [46-1:0] node605;
	wire [46-1:0] node608;
	wire [46-1:0] node611;
	wire [46-1:0] node612;
	wire [46-1:0] node613;
	wire [46-1:0] node616;
	wire [46-1:0] node620;
	wire [46-1:0] node621;
	wire [46-1:0] node622;
	wire [46-1:0] node623;
	wire [46-1:0] node624;
	wire [46-1:0] node625;
	wire [46-1:0] node628;
	wire [46-1:0] node631;
	wire [46-1:0] node632;
	wire [46-1:0] node635;
	wire [46-1:0] node638;
	wire [46-1:0] node639;
	wire [46-1:0] node640;
	wire [46-1:0] node643;
	wire [46-1:0] node646;
	wire [46-1:0] node647;
	wire [46-1:0] node650;
	wire [46-1:0] node653;
	wire [46-1:0] node654;
	wire [46-1:0] node655;
	wire [46-1:0] node656;
	wire [46-1:0] node659;
	wire [46-1:0] node662;
	wire [46-1:0] node663;
	wire [46-1:0] node666;
	wire [46-1:0] node669;
	wire [46-1:0] node670;
	wire [46-1:0] node671;
	wire [46-1:0] node674;
	wire [46-1:0] node677;
	wire [46-1:0] node678;
	wire [46-1:0] node681;
	wire [46-1:0] node684;
	wire [46-1:0] node685;
	wire [46-1:0] node686;
	wire [46-1:0] node687;
	wire [46-1:0] node688;
	wire [46-1:0] node691;
	wire [46-1:0] node694;
	wire [46-1:0] node695;
	wire [46-1:0] node698;
	wire [46-1:0] node701;
	wire [46-1:0] node702;
	wire [46-1:0] node703;
	wire [46-1:0] node706;
	wire [46-1:0] node709;
	wire [46-1:0] node710;
	wire [46-1:0] node713;
	wire [46-1:0] node716;
	wire [46-1:0] node717;
	wire [46-1:0] node718;
	wire [46-1:0] node719;
	wire [46-1:0] node722;
	wire [46-1:0] node725;
	wire [46-1:0] node726;
	wire [46-1:0] node729;
	wire [46-1:0] node732;
	wire [46-1:0] node733;
	wire [46-1:0] node734;
	wire [46-1:0] node737;
	wire [46-1:0] node740;
	wire [46-1:0] node741;
	wire [46-1:0] node744;
	wire [46-1:0] node747;
	wire [46-1:0] node748;
	wire [46-1:0] node749;
	wire [46-1:0] node750;
	wire [46-1:0] node752;
	wire [46-1:0] node753;
	wire [46-1:0] node754;
	wire [46-1:0] node755;
	wire [46-1:0] node758;
	wire [46-1:0] node761;
	wire [46-1:0] node762;
	wire [46-1:0] node766;
	wire [46-1:0] node767;
	wire [46-1:0] node768;
	wire [46-1:0] node773;
	wire [46-1:0] node774;
	wire [46-1:0] node775;
	wire [46-1:0] node776;
	wire [46-1:0] node778;
	wire [46-1:0] node782;
	wire [46-1:0] node783;
	wire [46-1:0] node784;
	wire [46-1:0] node787;
	wire [46-1:0] node790;
	wire [46-1:0] node792;
	wire [46-1:0] node797;
	wire [46-1:0] node798;
	wire [46-1:0] node799;
	wire [46-1:0] node800;
	wire [46-1:0] node801;
	wire [46-1:0] node802;
	wire [46-1:0] node803;
	wire [46-1:0] node806;
	wire [46-1:0] node809;
	wire [46-1:0] node810;
	wire [46-1:0] node813;
	wire [46-1:0] node816;
	wire [46-1:0] node817;
	wire [46-1:0] node818;
	wire [46-1:0] node821;
	wire [46-1:0] node824;
	wire [46-1:0] node825;
	wire [46-1:0] node828;
	wire [46-1:0] node831;
	wire [46-1:0] node832;
	wire [46-1:0] node833;
	wire [46-1:0] node834;
	wire [46-1:0] node837;
	wire [46-1:0] node840;
	wire [46-1:0] node841;
	wire [46-1:0] node844;
	wire [46-1:0] node847;
	wire [46-1:0] node848;
	wire [46-1:0] node849;
	wire [46-1:0] node852;
	wire [46-1:0] node855;
	wire [46-1:0] node856;
	wire [46-1:0] node859;
	wire [46-1:0] node862;
	wire [46-1:0] node863;
	wire [46-1:0] node864;
	wire [46-1:0] node865;
	wire [46-1:0] node866;
	wire [46-1:0] node869;
	wire [46-1:0] node872;
	wire [46-1:0] node873;
	wire [46-1:0] node876;
	wire [46-1:0] node879;
	wire [46-1:0] node880;
	wire [46-1:0] node881;
	wire [46-1:0] node884;
	wire [46-1:0] node887;
	wire [46-1:0] node888;
	wire [46-1:0] node891;
	wire [46-1:0] node894;
	wire [46-1:0] node895;
	wire [46-1:0] node896;
	wire [46-1:0] node897;
	wire [46-1:0] node900;
	wire [46-1:0] node903;
	wire [46-1:0] node904;
	wire [46-1:0] node907;
	wire [46-1:0] node910;
	wire [46-1:0] node911;
	wire [46-1:0] node912;
	wire [46-1:0] node915;
	wire [46-1:0] node918;
	wire [46-1:0] node919;
	wire [46-1:0] node922;
	wire [46-1:0] node925;
	wire [46-1:0] node926;
	wire [46-1:0] node927;
	wire [46-1:0] node928;
	wire [46-1:0] node929;
	wire [46-1:0] node930;
	wire [46-1:0] node933;
	wire [46-1:0] node936;
	wire [46-1:0] node937;
	wire [46-1:0] node940;
	wire [46-1:0] node943;
	wire [46-1:0] node944;
	wire [46-1:0] node945;
	wire [46-1:0] node948;
	wire [46-1:0] node951;
	wire [46-1:0] node952;
	wire [46-1:0] node955;
	wire [46-1:0] node958;
	wire [46-1:0] node959;
	wire [46-1:0] node960;
	wire [46-1:0] node961;
	wire [46-1:0] node964;
	wire [46-1:0] node967;
	wire [46-1:0] node968;
	wire [46-1:0] node971;
	wire [46-1:0] node974;
	wire [46-1:0] node975;
	wire [46-1:0] node976;
	wire [46-1:0] node979;
	wire [46-1:0] node982;
	wire [46-1:0] node983;
	wire [46-1:0] node986;
	wire [46-1:0] node989;
	wire [46-1:0] node990;
	wire [46-1:0] node991;
	wire [46-1:0] node992;
	wire [46-1:0] node993;
	wire [46-1:0] node996;
	wire [46-1:0] node999;
	wire [46-1:0] node1000;
	wire [46-1:0] node1003;
	wire [46-1:0] node1006;
	wire [46-1:0] node1007;
	wire [46-1:0] node1008;
	wire [46-1:0] node1011;
	wire [46-1:0] node1014;
	wire [46-1:0] node1015;
	wire [46-1:0] node1018;
	wire [46-1:0] node1021;
	wire [46-1:0] node1022;
	wire [46-1:0] node1023;
	wire [46-1:0] node1024;
	wire [46-1:0] node1027;
	wire [46-1:0] node1030;
	wire [46-1:0] node1031;
	wire [46-1:0] node1034;
	wire [46-1:0] node1037;
	wire [46-1:0] node1038;
	wire [46-1:0] node1039;
	wire [46-1:0] node1042;
	wire [46-1:0] node1045;
	wire [46-1:0] node1046;
	wire [46-1:0] node1049;
	wire [46-1:0] node1052;
	wire [46-1:0] node1053;
	wire [46-1:0] node1054;
	wire [46-1:0] node1055;
	wire [46-1:0] node1057;
	wire [46-1:0] node1059;
	wire [46-1:0] node1061;
	wire [46-1:0] node1063;
	wire [46-1:0] node1064;
	wire [46-1:0] node1067;
	wire [46-1:0] node1070;
	wire [46-1:0] node1071;
	wire [46-1:0] node1073;
	wire [46-1:0] node1075;
	wire [46-1:0] node1077;
	wire [46-1:0] node1078;
	wire [46-1:0] node1081;
	wire [46-1:0] node1084;
	wire [46-1:0] node1085;
	wire [46-1:0] node1086;
	wire [46-1:0] node1087;
	wire [46-1:0] node1088;
	wire [46-1:0] node1091;
	wire [46-1:0] node1094;
	wire [46-1:0] node1095;
	wire [46-1:0] node1098;
	wire [46-1:0] node1101;
	wire [46-1:0] node1102;
	wire [46-1:0] node1103;
	wire [46-1:0] node1106;
	wire [46-1:0] node1109;
	wire [46-1:0] node1110;
	wire [46-1:0] node1113;
	wire [46-1:0] node1116;
	wire [46-1:0] node1117;
	wire [46-1:0] node1119;
	wire [46-1:0] node1120;
	wire [46-1:0] node1123;
	wire [46-1:0] node1126;
	wire [46-1:0] node1127;
	wire [46-1:0] node1128;
	wire [46-1:0] node1131;
	wire [46-1:0] node1135;
	wire [46-1:0] node1136;
	wire [46-1:0] node1137;
	wire [46-1:0] node1138;
	wire [46-1:0] node1139;
	wire [46-1:0] node1140;
	wire [46-1:0] node1141;
	wire [46-1:0] node1144;
	wire [46-1:0] node1147;
	wire [46-1:0] node1148;
	wire [46-1:0] node1151;
	wire [46-1:0] node1154;
	wire [46-1:0] node1155;
	wire [46-1:0] node1156;
	wire [46-1:0] node1159;
	wire [46-1:0] node1162;
	wire [46-1:0] node1163;
	wire [46-1:0] node1166;
	wire [46-1:0] node1169;
	wire [46-1:0] node1170;
	wire [46-1:0] node1171;
	wire [46-1:0] node1172;
	wire [46-1:0] node1175;
	wire [46-1:0] node1178;
	wire [46-1:0] node1179;
	wire [46-1:0] node1182;
	wire [46-1:0] node1185;
	wire [46-1:0] node1186;
	wire [46-1:0] node1187;
	wire [46-1:0] node1190;
	wire [46-1:0] node1193;
	wire [46-1:0] node1194;
	wire [46-1:0] node1197;
	wire [46-1:0] node1200;
	wire [46-1:0] node1201;
	wire [46-1:0] node1202;
	wire [46-1:0] node1203;
	wire [46-1:0] node1204;
	wire [46-1:0] node1207;
	wire [46-1:0] node1210;
	wire [46-1:0] node1211;
	wire [46-1:0] node1214;
	wire [46-1:0] node1217;
	wire [46-1:0] node1218;
	wire [46-1:0] node1219;
	wire [46-1:0] node1222;
	wire [46-1:0] node1225;
	wire [46-1:0] node1226;
	wire [46-1:0] node1229;
	wire [46-1:0] node1232;
	wire [46-1:0] node1233;
	wire [46-1:0] node1234;
	wire [46-1:0] node1235;
	wire [46-1:0] node1238;
	wire [46-1:0] node1241;
	wire [46-1:0] node1242;
	wire [46-1:0] node1245;
	wire [46-1:0] node1248;
	wire [46-1:0] node1249;
	wire [46-1:0] node1250;
	wire [46-1:0] node1253;
	wire [46-1:0] node1256;
	wire [46-1:0] node1257;
	wire [46-1:0] node1260;
	wire [46-1:0] node1263;
	wire [46-1:0] node1264;
	wire [46-1:0] node1265;
	wire [46-1:0] node1266;
	wire [46-1:0] node1267;
	wire [46-1:0] node1268;
	wire [46-1:0] node1271;
	wire [46-1:0] node1274;
	wire [46-1:0] node1275;
	wire [46-1:0] node1278;
	wire [46-1:0] node1281;
	wire [46-1:0] node1282;
	wire [46-1:0] node1283;
	wire [46-1:0] node1286;
	wire [46-1:0] node1289;
	wire [46-1:0] node1290;
	wire [46-1:0] node1293;
	wire [46-1:0] node1296;
	wire [46-1:0] node1297;
	wire [46-1:0] node1298;
	wire [46-1:0] node1299;
	wire [46-1:0] node1302;
	wire [46-1:0] node1305;
	wire [46-1:0] node1306;
	wire [46-1:0] node1309;
	wire [46-1:0] node1312;
	wire [46-1:0] node1313;
	wire [46-1:0] node1314;
	wire [46-1:0] node1317;
	wire [46-1:0] node1320;
	wire [46-1:0] node1321;
	wire [46-1:0] node1324;
	wire [46-1:0] node1327;
	wire [46-1:0] node1328;
	wire [46-1:0] node1329;
	wire [46-1:0] node1330;
	wire [46-1:0] node1331;
	wire [46-1:0] node1334;
	wire [46-1:0] node1337;
	wire [46-1:0] node1338;
	wire [46-1:0] node1341;
	wire [46-1:0] node1344;
	wire [46-1:0] node1345;
	wire [46-1:0] node1346;
	wire [46-1:0] node1349;
	wire [46-1:0] node1352;
	wire [46-1:0] node1353;
	wire [46-1:0] node1356;
	wire [46-1:0] node1359;
	wire [46-1:0] node1360;
	wire [46-1:0] node1361;
	wire [46-1:0] node1362;
	wire [46-1:0] node1365;
	wire [46-1:0] node1368;
	wire [46-1:0] node1369;
	wire [46-1:0] node1372;
	wire [46-1:0] node1375;
	wire [46-1:0] node1376;
	wire [46-1:0] node1377;
	wire [46-1:0] node1380;
	wire [46-1:0] node1383;
	wire [46-1:0] node1384;
	wire [46-1:0] node1387;
	wire [46-1:0] node1390;
	wire [46-1:0] node1391;
	wire [46-1:0] node1392;
	wire [46-1:0] node1393;
	wire [46-1:0] node1394;
	wire [46-1:0] node1395;
	wire [46-1:0] node1398;
	wire [46-1:0] node1403;
	wire [46-1:0] node1404;
	wire [46-1:0] node1405;
	wire [46-1:0] node1406;
	wire [46-1:0] node1409;
	wire [46-1:0] node1412;
	wire [46-1:0] node1413;
	wire [46-1:0] node1416;
	wire [46-1:0] node1419;
	wire [46-1:0] node1420;
	wire [46-1:0] node1421;
	wire [46-1:0] node1424;
	wire [46-1:0] node1428;
	wire [46-1:0] node1429;
	wire [46-1:0] node1430;
	wire [46-1:0] node1431;
	wire [46-1:0] node1432;
	wire [46-1:0] node1435;
	wire [46-1:0] node1438;
	wire [46-1:0] node1439;
	wire [46-1:0] node1442;
	wire [46-1:0] node1445;
	wire [46-1:0] node1446;
	wire [46-1:0] node1447;
	wire [46-1:0] node1450;
	wire [46-1:0] node1454;
	wire [46-1:0] node1455;
	wire [46-1:0] node1456;
	wire [46-1:0] node1457;
	wire [46-1:0] node1460;

	assign outp = (inp[1]) ? node264 : node1;
		assign node1 = (inp[3]) ? node5 : node2;
			assign node2 = (inp[15]) ? 46'b0000000000000000000000000000001000000000000000 : 46'b0000000000000000000000000000000000000000000000;
			assign node5 = (inp[15]) ? node63 : node6;
				assign node6 = (inp[7]) ? node8 : 46'b0000000000000000000000000000000000000000000000;
					assign node8 = (inp[5]) ? node10 : 46'b0000000000000000000000000000000000000000000000;
						assign node10 = (inp[9]) ? node24 : node11;
							assign node11 = (inp[6]) ? node13 : 46'b0000000000000000000000000000000000000000000000;
								assign node13 = (inp[13]) ? node15 : 46'b0000000000000000000000000000000000000000000000;
									assign node15 = (inp[11]) ? 46'b0000000000000000000000000000000000000000000000 : node16;
										assign node16 = (inp[2]) ? node18 : 46'b0000000000000000000000000000000000000000000000;
											assign node18 = (inp[0]) ? 46'b0000000000000000000000000000000000000000000000 : node19;
												assign node19 = (inp[12]) ? 46'b0000000000000000000000000000000000000100000000 : 46'b0000000000000000000000000000000000000000000000;
							assign node24 = (inp[12]) ? node26 : 46'b0000000000000000000000000000000000000000000000;
								assign node26 = (inp[2]) ? node40 : node27;
									assign node27 = (inp[13]) ? 46'b0000000000000000000000000000000000000000000000 : node28;
										assign node28 = (inp[0]) ? node30 : 46'b0000000000000000000000000000000000000000000000;
											assign node30 = (inp[6]) ? node32 : 46'b0000000000000000000000000000000000000000000000;
												assign node32 = (inp[11]) ? node34 : 46'b0000000000000000000000000000000000000000000000;
													assign node34 = (inp[14]) ? node36 : 46'b0000000000000000000000000000000000000000000000;
														assign node36 = (inp[10]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0000000000000000000000000000000000000000000000;
									assign node40 = (inp[13]) ? node52 : node41;
										assign node41 = (inp[14]) ? node43 : 46'b0000000000000000000000000000000000000000000000;
											assign node43 = (inp[10]) ? node45 : 46'b0000000000000000000000000000000000000000000000;
												assign node45 = (inp[8]) ? node47 : 46'b0000000000000000000000000000000000000000000000;
													assign node47 = (inp[6]) ? node49 : 46'b0000000000000000000000000000000000000000000000;
														assign node49 = (inp[11]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0000000000000000000000000000000000000000000000;
										assign node52 = (inp[8]) ? node54 : 46'b0000000000000000000000000000000000000000000000;
											assign node54 = (inp[10]) ? node56 : 46'b0000000000000000000000000000000000000000000000;
												assign node56 = (inp[6]) ? node58 : 46'b0000000000000000000000000000000000000000000000;
													assign node58 = (inp[0]) ? node60 : 46'b0000000000000000000000000000000000000000000000;
														assign node60 = (inp[4]) ? 46'b0000100001000000000000000000000000000000000000 : 46'b0000000000000000000000000000000000000000000000;
				assign node63 = (inp[9]) ? node117 : node64;
					assign node64 = (inp[11]) ? node104 : node65;
						assign node65 = (inp[13]) ? node71 : node66;
							assign node66 = (inp[2]) ? 46'b0000000000000000000000000000000000000000000000 : node67;
								assign node67 = (inp[0]) ? 46'b0000000000001000000000000010000000000000000000 : 46'b0000001000001000000000000000000000000000000000;
							assign node71 = (inp[0]) ? 46'b0000000000000000000000000000000000000000000000 : node72;
								assign node72 = (inp[6]) ? node74 : 46'b0000000000000000000000000000000000000000000000;
									assign node74 = (inp[14]) ? node76 : 46'b0000000000000000000000000000000000000000000000;
										assign node76 = (inp[5]) ? node78 : 46'b0000000000000000000000000000000000000000000000;
											assign node78 = (inp[2]) ? node90 : node79;
												assign node79 = (inp[12]) ? node85 : node80;
													assign node80 = (inp[7]) ? node82 : 46'b0000000000000000000000000000000000000000000000;
														assign node82 = (inp[8]) ? 46'b0000000000001000010100000000000000000000010000 : 46'b0000000000000000000000000000000000000000000000;
													assign node85 = (inp[7]) ? 46'b0000000000000000000000000000000000000000000000 : node86;
														assign node86 = (inp[4]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0000000000000000000000000000000000000000000000;
												assign node90 = (inp[10]) ? node96 : node91;
													assign node91 = (inp[4]) ? node93 : 46'b0000000000000000000000000000000000000000000000;
														assign node93 = (inp[7]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0000000000000000000000000000000000000000000000;
													assign node96 = (inp[12]) ? node100 : node97;
														assign node97 = (inp[7]) ? 46'b0000000000001000010000000000000001000010000000 : 46'b0000000000000000000000000000000000000000000000;
														assign node100 = (inp[7]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0000010000000000010000000000000001000010000000;
						assign node104 = (inp[13]) ? node110 : node105;
							assign node105 = (inp[2]) ? 46'b0000000000000000000000000000000000000000000000 : node106;
								assign node106 = (inp[0]) ? 46'b0000010000000000000000000010000000000000000000 : 46'b0000011000000000000000000000000000000000000000;
							assign node110 = (inp[2]) ? node114 : node111;
								assign node111 = (inp[0]) ? 46'b0000001000000000011000000100000000000000010000 : 46'b0000001000000000010000000100000000000000010010;
								assign node114 = (inp[0]) ? 46'b0000001000000000010010000000010000000010000000 : 46'b0000001000000000010010100000000000000010000000;
					assign node117 = (inp[2]) ? node213 : node118;
						assign node118 = (inp[0]) ? node164 : node119;
							assign node119 = (inp[13]) ? node123 : node120;
								assign node120 = (inp[11]) ? 46'b0000010100000000000000000000000000000000000000 : 46'b0000000100001000000000000000000000000000000000;
								assign node123 = (inp[14]) ? node125 : 46'b0000000000000000000000000000000000000000000000;
									assign node125 = (inp[5]) ? node127 : 46'b0000000000000000000000000000000000000000000000;
										assign node127 = (inp[6]) ? node137 : node128;
											assign node128 = (inp[4]) ? node130 : 46'b0000000000000000000000000000000000000000000000;
												assign node130 = (inp[11]) ? node132 : 46'b0000000000000000000000000000000000000000000000;
													assign node132 = (inp[8]) ? node134 : 46'b0000000000000000000000000000000000000000000000;
														assign node134 = (inp[10]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0000000000000000000000000000000000000000000000;
											assign node137 = (inp[11]) ? node151 : node138;
												assign node138 = (inp[7]) ? node146 : node139;
													assign node139 = (inp[12]) ? node143 : node140;
														assign node140 = (inp[10]) ? 46'b0010000000000000000000000000000000000000010000 : 46'b0000000000000000000000000000000000000000000000;
														assign node143 = (inp[8]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0000000000000000000000000000000000000000000000;
													assign node146 = (inp[12]) ? 46'b0000000000000000000000000000000000000000000000 : node147;
														assign node147 = (inp[4]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0000000000000000000000000000000000000000000000;
												assign node151 = (inp[8]) ? node157 : node152;
													assign node152 = (inp[4]) ? node154 : 46'b0000000000000000000000000000000000000000000000;
														assign node154 = (inp[10]) ? 46'b0000000000010000010000000100000000000000010010 : 46'b0000000000000000000000000000000000000000000000;
													assign node157 = (inp[12]) ? node161 : node158;
														assign node158 = (inp[7]) ? 46'b0000000000001000010000000100000000000000010010 : 46'b0000000000000000000000000000000000000000000000;
														assign node161 = (inp[7]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0000000000000000000000000000000000000000000000;
							assign node164 = (inp[11]) ? node186 : node165;
								assign node165 = (inp[13]) ? node167 : 46'b0010001000000000000000000000000000000000010000;
									assign node167 = (inp[6]) ? node169 : 46'b0000000000000000000000000000000000000000000000;
										assign node169 = (inp[14]) ? node171 : 46'b0000000000000000000000000000000000000000000000;
											assign node171 = (inp[5]) ? node173 : 46'b0000000000000000000000000000000000000000000000;
												assign node173 = (inp[7]) ? node181 : node174;
													assign node174 = (inp[12]) ? node178 : node175;
														assign node175 = (inp[4]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0000000000000000000000000000000000000000000000;
														assign node178 = (inp[8]) ? 46'b0000010000000000010000000000000000000000010100 : 46'b0000000000000000000000000000000000000000000000;
													assign node181 = (inp[12]) ? 46'b0000000000000000000000000000000000000000000000 : node182;
														assign node182 = (inp[10]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0000000000000000000000000000000000000000000000;
								assign node186 = (inp[14]) ? node188 : 46'b0000000000000000000000000000000000000000000000;
									assign node188 = (inp[13]) ? node190 : 46'b0000000000000000000000000000000000000000000000;
										assign node190 = (inp[5]) ? node192 : 46'b0000000000000000000000000000000000000000000000;
											assign node192 = (inp[6]) ? node200 : node193;
												assign node193 = (inp[10]) ? node195 : 46'b0000000000000000000000000000000000000000000000;
													assign node195 = (inp[4]) ? node197 : 46'b0000000000000000000000000000000000000000000000;
														assign node197 = (inp[8]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0000000000000000000000000000000000000000000000;
												assign node200 = (inp[12]) ? node208 : node201;
													assign node201 = (inp[8]) ? node205 : node202;
														assign node202 = (inp[4]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0000000000000000000000000000000000000000000000;
														assign node205 = (inp[4]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0000000000000000001000010100000000000000010000;
													assign node208 = (inp[7]) ? 46'b0000000000000000000000000000000000000000000000 : node209;
														assign node209 = (inp[4]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0000000000000000000000000000000000000000000000;
						assign node213 = (inp[14]) ? node215 : 46'b0000000000000000000000000000000000000000000000;
							assign node215 = (inp[5]) ? node217 : 46'b0000000000000000000000000000000000000000000000;
								assign node217 = (inp[13]) ? node219 : 46'b0000000000000000000000000000000000000000000000;
									assign node219 = (inp[6]) ? node231 : node220;
										assign node220 = (inp[4]) ? node222 : 46'b0000000000000000000000000000000000000000000000;
											assign node222 = (inp[11]) ? node224 : 46'b0000000000000000000000000000000000000000000000;
												assign node224 = (inp[10]) ? node226 : 46'b0000000000000000000000000000000000000000000000;
													assign node226 = (inp[8]) ? node228 : 46'b0000000000000000000000000000000000000000000000;
														assign node228 = (inp[7]) ? 46'b0000000000000000000010000000010000000000000000 : 46'b0000000000000000000110000000010000000000000000;
										assign node231 = (inp[8]) ? node243 : node232;
											assign node232 = (inp[10]) ? node234 : 46'b0000000000000000000000000000000000000000000000;
												assign node234 = (inp[4]) ? node236 : 46'b0000000000000000000000000000000000000000000000;
													assign node236 = (inp[12]) ? node240 : node237;
														assign node237 = (inp[11]) ? 46'b0010000000010000000010000000000000000010000000 : 46'b0000000000000000000000000000000000000000000000;
														assign node240 = (inp[7]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0000000000000000000000000000000000000000000000;
											assign node243 = (inp[11]) ? node253 : node244;
												assign node244 = (inp[0]) ? 46'b0000000000000000000000000000000000000000000000 : node245;
													assign node245 = (inp[7]) ? node249 : node246;
														assign node246 = (inp[12]) ? 46'b0000010000000000010000000000000100000010000000 : 46'b0010000000000000000000000000000000000010000000;
														assign node249 = (inp[12]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0000000000000000000000000000000000000000000000;
												assign node253 = (inp[10]) ? node259 : node254;
													assign node254 = (inp[4]) ? node256 : 46'b0000000000000000000000000000000000000000000000;
														assign node256 = (inp[12]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0000000000001000010010000000000100000010000000;
													assign node259 = (inp[4]) ? 46'b0000000000000000000000000000000000000000000000 : node260;
														assign node260 = (inp[0]) ? 46'b0000000000000000010010010000010000000010000000 : 46'b0000000000000000010010110000000000000010000000;
		assign node264 = (inp[15]) ? node332 : node265;
			assign node265 = (inp[13]) ? node269 : node266;
				assign node266 = (inp[3]) ? 46'b0000100000000000000000000000001000000000000000 : 46'b0000100000000000000000000000000000000000000000;
				assign node269 = (inp[2]) ? node301 : node270;
					assign node270 = (inp[9]) ? node286 : node271;
						assign node271 = (inp[11]) ? node279 : node272;
							assign node272 = (inp[0]) ? node276 : node273;
								assign node273 = (inp[3]) ? 46'b0000100000001000010000010100001000000000010010 : 46'b0000100000001000010000010100000000000000010010;
								assign node276 = (inp[3]) ? 46'b0000100000001000010000000100001100000000010010 : 46'b0000100000001000010000000100000100000000010010;
							assign node279 = (inp[0]) ? node283 : node280;
								assign node280 = (inp[3]) ? 46'b0000100000001000011000010100001000000000010000 : 46'b0000100000001000011000010100000000000000010000;
								assign node283 = (inp[3]) ? 46'b0000100000001000011000000100001100000000010000 : 46'b0000100000001000011000000100000100000000010000;
						assign node286 = (inp[0]) ? node294 : node287;
							assign node287 = (inp[11]) ? node291 : node288;
								assign node288 = (inp[3]) ? 46'b0000110000000000010000010100001000000000010010 : 46'b0000110000000000010000010100000000000000010010;
								assign node291 = (inp[3]) ? 46'b0000110000000000011000010100001000000000010000 : 46'b0000110000000000011000010100000000000000010000;
							assign node294 = (inp[11]) ? node298 : node295;
								assign node295 = (inp[3]) ? 46'b0000110000000000010000000100001100000000010010 : 46'b0000110000000000010000000100000100000000010010;
								assign node298 = (inp[3]) ? 46'b0000110000000000011000000100001100000000010000 : 46'b0000110000000000011000000100000100000000010000;
					assign node301 = (inp[0]) ? node317 : node302;
						assign node302 = (inp[11]) ? node310 : node303;
							assign node303 = (inp[9]) ? node307 : node304;
								assign node304 = (inp[3]) ? 46'b0000100000001000010010110000001000000010000000 : 46'b0000100000001000010010110000000000000010000000;
								assign node307 = (inp[3]) ? 46'b0000110000000000010010110000001000000010000000 : 46'b0000110000000000010010110000000000000010000000;
							assign node310 = (inp[9]) ? node314 : node311;
								assign node311 = (inp[3]) ? 46'b0000100000001000010010010000011000000010000000 : 46'b0000100000001000010010010000010000000010000000;
								assign node314 = (inp[3]) ? 46'b0000110000000000010010010000011000000010000000 : 46'b0000110000000000010010010000010000000010000000;
						assign node317 = (inp[11]) ? node325 : node318;
							assign node318 = (inp[9]) ? node322 : node319;
								assign node319 = (inp[3]) ? 46'b0000100000001000010010100000001100000010000000 : 46'b0000100000001000010010100000000100000010000000;
								assign node322 = (inp[3]) ? 46'b0000110000000000010010100000001100000010000000 : 46'b0000110000000000010010100000000100000010000000;
							assign node325 = (inp[9]) ? node329 : node326;
								assign node326 = (inp[3]) ? 46'b0000100000001000010010000000011100000010000000 : 46'b0000100000001000010010000000010100000010000000;
								assign node329 = (inp[3]) ? 46'b0000110000000000010010000000011100000010000000 : 46'b0000110000000000010010000000010100000010000000;
			assign node332 = (inp[13]) ? node336 : node333;
				assign node333 = (inp[3]) ? 46'b0000000000000000000000000000000000000000001000 : 46'b0000000000000000000000000000001000000000001000;
				assign node336 = (inp[3]) ? node338 : 46'b0000000000000000000000000000001000000000000000;
					assign node338 = (inp[2]) ? node1052 : node339;
						assign node339 = (inp[9]) ? node747 : node340;
							assign node340 = (inp[11]) ? node596 : node341;
								assign node341 = (inp[0]) ? node469 : node342;
									assign node342 = (inp[5]) ? node406 : node343;
										assign node343 = (inp[12]) ? node375 : node344;
											assign node344 = (inp[6]) ? node360 : node345;
												assign node345 = (inp[7]) ? node353 : node346;
													assign node346 = (inp[10]) ? node350 : node347;
														assign node347 = (inp[4]) ? 46'b0011000000000000001000010001100010110001010000 : 46'b0011000000000100000000010000100010110001010000;
														assign node350 = (inp[4]) ? 46'b0011000000000010000000010000100010110001010000 : 46'b0011000000000000000000010001100010110001010010;
													assign node353 = (inp[14]) ? node357 : node354;
														assign node354 = (inp[4]) ? 46'b0011000000000100001000010001000010110001010000 : 46'b0011000000000100000000010001000010110001010010;
														assign node357 = (inp[8]) ? 46'b0011000000000010000000010000000010110001010000 : 46'b0011000000000000001000010001000010110001010000;
												assign node360 = (inp[7]) ? node368 : node361;
													assign node361 = (inp[4]) ? node365 : node362;
														assign node362 = (inp[10]) ? 46'b0011000000000000000000010001100010010001010010 : 46'b0011000000000100000000010000100010010001010000;
														assign node365 = (inp[10]) ? 46'b0011000000000010000000010000100010010001010000 : 46'b0011000000000000001000010001100010010001010000;
													assign node368 = (inp[8]) ? node372 : node369;
														assign node369 = (inp[14]) ? 46'b0011000000000000001000010001000010010001010000 : 46'b0011000000000100000000010000000010010001010000;
														assign node372 = (inp[14]) ? 46'b0011000000000010000000010000000010010001010000 : 46'b0011000000000000000000010001000010010001010010;
											assign node375 = (inp[7]) ? node391 : node376;
												assign node376 = (inp[6]) ? node384 : node377;
													assign node377 = (inp[8]) ? node381 : node378;
														assign node378 = (inp[14]) ? 46'b0011000000000000001000010001100000110001010000 : 46'b0011000000000100000000010000100000110001010000;
														assign node381 = (inp[14]) ? 46'b0011000000000010000000010001100000110001010000 : 46'b0011000000000000000000010001100000110001010010;
													assign node384 = (inp[4]) ? node388 : node385;
														assign node385 = (inp[10]) ? 46'b0011000000000000000000010001100000010001010010 : 46'b0011000000000100000000010000100000010001010000;
														assign node388 = (inp[10]) ? 46'b0011000000000010000000010001100000010001010000 : 46'b0011000000000000001000010001100000010001010000;
												assign node391 = (inp[6]) ? node399 : node392;
													assign node392 = (inp[14]) ? node396 : node393;
														assign node393 = (inp[8]) ? 46'b0011000000000000000000010001000000110001010010 : 46'b0011000000000100000000010000000000110001010000;
														assign node396 = (inp[8]) ? 46'b0011000000000010000000010000000000110001010000 : 46'b0011000000000000001000010001000000110001010000;
													assign node399 = (inp[14]) ? node403 : node400;
														assign node400 = (inp[10]) ? 46'b0011000000000010000000010000000000010001010000 : 46'b0011000000000100001000010001000000010001010010;
														assign node403 = (inp[4]) ? 46'b0011000000000000001000010001000000010001010000 : 46'b0011000000000000001000010001000000010001010010;
										assign node406 = (inp[12]) ? node438 : node407;
											assign node407 = (inp[6]) ? node423 : node408;
												assign node408 = (inp[7]) ? node416 : node409;
													assign node409 = (inp[10]) ? node413 : node410;
														assign node410 = (inp[4]) ? 46'b0010000000000000001000010001100010110001010000 : 46'b0010000000000100000000010000100010110001010000;
														assign node413 = (inp[4]) ? 46'b0010000000000010000000010000100010110001010000 : 46'b0010000000000000000000010001100010110001010010;
													assign node416 = (inp[14]) ? node420 : node417;
														assign node417 = (inp[8]) ? 46'b0010000000000000000000010001000010110001010010 : 46'b0010000000000100000000010000000010110001010000;
														assign node420 = (inp[4]) ? 46'b0010000000000010001000010001000010110001010000 : 46'b0010000000000000000000010001000010110001010010;
												assign node423 = (inp[7]) ? node431 : node424;
													assign node424 = (inp[4]) ? node428 : node425;
														assign node425 = (inp[10]) ? 46'b0010000000000000000000010001100010010001010010 : 46'b0010000000000100000000010000100010010001010000;
														assign node428 = (inp[10]) ? 46'b0010000000000010000000010000100010010001010000 : 46'b0010000000000000001000010001100010010001010000;
													assign node431 = (inp[4]) ? node435 : node432;
														assign node432 = (inp[10]) ? 46'b0010000000000000000000010001000010010001010010 : 46'b0010000000000100000000010000000010010001010000;
														assign node435 = (inp[10]) ? 46'b0010000000000010000000010000000010010001010000 : 46'b0010000000000000001000010001000010010001010000;
											assign node438 = (inp[7]) ? node454 : node439;
												assign node439 = (inp[6]) ? node447 : node440;
													assign node440 = (inp[4]) ? node444 : node441;
														assign node441 = (inp[10]) ? 46'b0010000000000000000000010001100000110001010010 : 46'b0010000000000100000000010001100000110001010000;
														assign node444 = (inp[10]) ? 46'b0010000000000010000000010000100000110001010000 : 46'b0010000000000000001000010001100000110001010000;
													assign node447 = (inp[8]) ? node451 : node448;
														assign node448 = (inp[14]) ? 46'b0010000000000000001000010001100000010001010000 : 46'b0010000000000100000000010000100000010001010000;
														assign node451 = (inp[14]) ? 46'b0010000000000010000000010000100000010001010000 : 46'b0010000000000000000000010001100000010001010010;
												assign node454 = (inp[6]) ? node462 : node455;
													assign node455 = (inp[4]) ? node459 : node456;
														assign node456 = (inp[10]) ? 46'b0010000000000000000000010001000000110001010010 : 46'b0010000000000100000000010000000000110001010000;
														assign node459 = (inp[14]) ? 46'b0010000000000000001000010001000000110001010000 : 46'b0010000000000100001000010001000000110001010000;
													assign node462 = (inp[4]) ? node466 : node463;
														assign node463 = (inp[10]) ? 46'b0010000000000000000000010001000000010001010010 : 46'b0010000000000100000000010000000000010001010000;
														assign node466 = (inp[10]) ? 46'b0010000000000010000000010000000000010001010000 : 46'b0010000000000000001000010001000000010001010000;
									assign node469 = (inp[5]) ? node533 : node470;
										assign node470 = (inp[6]) ? node502 : node471;
											assign node471 = (inp[12]) ? node487 : node472;
												assign node472 = (inp[7]) ? node480 : node473;
													assign node473 = (inp[4]) ? node477 : node474;
														assign node474 = (inp[10]) ? 46'b0011000000000000000000010001100010110000010010 : 46'b0011000000000100000000010001100010110000010000;
														assign node477 = (inp[10]) ? 46'b0011000000000010000000010000100010110000010000 : 46'b0011000000000000001000010001100010110000010000;
													assign node480 = (inp[4]) ? node484 : node481;
														assign node481 = (inp[10]) ? 46'b0011000000000000000000010001000010110000010010 : 46'b0011000000000100000000010000000010110000010000;
														assign node484 = (inp[10]) ? 46'b0011000000000010000000010000000010110000010000 : 46'b0011000000000000001000010001000010110000010000;
												assign node487 = (inp[7]) ? node495 : node488;
													assign node488 = (inp[8]) ? node492 : node489;
														assign node489 = (inp[14]) ? 46'b0011000000000000001000010001100000110000010000 : 46'b0011000000000100000000010001100000110000010000;
														assign node492 = (inp[14]) ? 46'b0011000000000010000000010000100000110000010000 : 46'b0011000000000100000000010001100000110000010010;
													assign node495 = (inp[8]) ? node499 : node496;
														assign node496 = (inp[14]) ? 46'b0011000000000000001000010001000000110000010000 : 46'b0011000000000100000000010001000000110000010000;
														assign node499 = (inp[4]) ? 46'b0011000000000010001000010001000000110000010010 : 46'b0011000000000110000000010001000000110000010010;
											assign node502 = (inp[12]) ? node518 : node503;
												assign node503 = (inp[7]) ? node511 : node504;
													assign node504 = (inp[10]) ? node508 : node505;
														assign node505 = (inp[4]) ? 46'b0011000000000000001000010001100010010000010000 : 46'b0011000000000100000000010001100010010000010000;
														assign node508 = (inp[4]) ? 46'b0011000000000010000000010000100010010000010000 : 46'b0011000000000000000000010001100010010000010010;
													assign node511 = (inp[8]) ? node515 : node512;
														assign node512 = (inp[14]) ? 46'b0011000000000000001000010001000010010000010000 : 46'b0011000000000100000000010000000010010000010000;
														assign node515 = (inp[10]) ? 46'b0011000000000010000000010001000010010000010010 : 46'b0011000000000000001000010001000010010000010000;
												assign node518 = (inp[7]) ? node526 : node519;
													assign node519 = (inp[10]) ? node523 : node520;
														assign node520 = (inp[4]) ? 46'b0011000000000000001000010001100000010000010000 : 46'b0011000000000100000000010000100000010000010000;
														assign node523 = (inp[4]) ? 46'b0011000000000010000000010000100000010000010000 : 46'b0011000000000000000000010001100000010000010010;
													assign node526 = (inp[4]) ? node530 : node527;
														assign node527 = (inp[10]) ? 46'b0011000000000000000000010001000000010000010010 : 46'b0011000000000100000000010000000000010000010000;
														assign node530 = (inp[8]) ? 46'b0011000000000000001000010001000000010000010000 : 46'b0011000000000100001000010001000000010000010000;
										assign node533 = (inp[6]) ? node565 : node534;
											assign node534 = (inp[12]) ? node550 : node535;
												assign node535 = (inp[7]) ? node543 : node536;
													assign node536 = (inp[10]) ? node540 : node537;
														assign node537 = (inp[4]) ? 46'b0010000000000000001000010001100010110000010000 : 46'b0010000000000100000000010000100010110000010000;
														assign node540 = (inp[4]) ? 46'b0010000000000010000000010000100010110000010000 : 46'b0010000000000000000000010001100010110000010010;
													assign node543 = (inp[10]) ? node547 : node544;
														assign node544 = (inp[8]) ? 46'b0010000000000000001000010001000010110000010010 : 46'b0010000000000100001000010001000010110000010000;
														assign node547 = (inp[4]) ? 46'b0010000000000010000000010000000010110000010000 : 46'b0010000000000000000000010001000010110000010010;
												assign node550 = (inp[7]) ? node558 : node551;
													assign node551 = (inp[10]) ? node555 : node552;
														assign node552 = (inp[4]) ? 46'b0010000000000000001000010001100000110000010000 : 46'b0010000000000100000000010000100000110000010000;
														assign node555 = (inp[4]) ? 46'b0010000000000010000000010001100000110000010000 : 46'b0010000000000000000000010001100000110000010010;
													assign node558 = (inp[4]) ? node562 : node559;
														assign node559 = (inp[10]) ? 46'b0010000000000000000000010001000000110000010010 : 46'b0010000000000100001000010001000000110000010000;
														assign node562 = (inp[14]) ? 46'b0010000000000010001000010001000000110000010000 : 46'b0010000000000100000000010000000000110000010000;
											assign node565 = (inp[12]) ? node581 : node566;
												assign node566 = (inp[7]) ? node574 : node567;
													assign node567 = (inp[8]) ? node571 : node568;
														assign node568 = (inp[14]) ? 46'b0010000000000000001000010001100010010000010000 : 46'b0010000000000100000000010001100010010000010000;
														assign node571 = (inp[14]) ? 46'b0010000000000010000000010000100010010000010000 : 46'b0010000000000000000000010001100010010000010010;
													assign node574 = (inp[14]) ? node578 : node575;
														assign node575 = (inp[8]) ? 46'b0010000000000000000000010001000010010000010010 : 46'b0010000000000100000000010001000010010000010000;
														assign node578 = (inp[8]) ? 46'b0010000000000010000000010000000010010000010000 : 46'b0010000000000000001000010001000010010000010000;
												assign node581 = (inp[7]) ? node589 : node582;
													assign node582 = (inp[14]) ? node586 : node583;
														assign node583 = (inp[8]) ? 46'b0010000000000000000000010001100000010000010010 : 46'b0010000000000100000000010000100000010000010000;
														assign node586 = (inp[8]) ? 46'b0010000000000010000000010001100000010000010000 : 46'b0010000000000000001000010001100000010000010000;
													assign node589 = (inp[10]) ? node593 : node590;
														assign node590 = (inp[4]) ? 46'b0010000000000000001000010001000000010000010000 : 46'b0010000000000100000000010000000000010000010000;
														assign node593 = (inp[4]) ? 46'b0010000000000010000000010000000000010000010000 : 46'b0010000000000000000000010001000000010000010010;
								assign node596 = (inp[0]) ? node620 : node597;
									assign node597 = (inp[7]) ? node599 : 46'b0000000000000000000000000000000000000000000000;
										assign node599 = (inp[5]) ? node601 : 46'b0000000000000000000000000000000000000000000000;
											assign node601 = (inp[6]) ? node611 : node602;
												assign node602 = (inp[12]) ? node604 : 46'b0000000000000000000000000000000000000000000000;
													assign node604 = (inp[8]) ? node608 : node605;
														assign node605 = (inp[14]) ? 46'b0000000000000000001001000001000000100000000000 : 46'b0000000000000100000001000000000000100000000000;
														assign node608 = (inp[14]) ? 46'b0000000000000010000001000000000000100000000000 : 46'b0000000000000000000001000001000000100000000010;
												assign node611 = (inp[12]) ? 46'b0000000000000000000000000000000000000000000000 : node612;
													assign node612 = (inp[10]) ? node616 : node613;
														assign node613 = (inp[4]) ? 46'b0000000000000000001001000001000010000000000000 : 46'b0000000000000100000001000001000010000000000000;
														assign node616 = (inp[4]) ? 46'b0000000000000010000001000000000010000000000000 : 46'b0000000000000000000001000001000010000000000010;
									assign node620 = (inp[6]) ? node684 : node621;
										assign node621 = (inp[7]) ? node653 : node622;
											assign node622 = (inp[12]) ? node638 : node623;
												assign node623 = (inp[5]) ? node631 : node624;
													assign node624 = (inp[14]) ? node628 : node625;
														assign node625 = (inp[8]) ? 46'b0101000000000000000000000001100010100000000010 : 46'b0101000000000100000000000000100010100000000000;
														assign node628 = (inp[8]) ? 46'b0101000000000010000000000000100010100000000000 : 46'b0101000000000000001000000001100010100000000000;
													assign node631 = (inp[4]) ? node635 : node632;
														assign node632 = (inp[10]) ? 46'b0100000000000000000000000001100010100000000010 : 46'b0100000000000100000000000000100010100000000000;
														assign node635 = (inp[10]) ? 46'b0100000000000010000000000000100010100000000000 : 46'b0100000000000000001000000001100010100000000000;
												assign node638 = (inp[5]) ? node646 : node639;
													assign node639 = (inp[14]) ? node643 : node640;
														assign node640 = (inp[8]) ? 46'b0101000000000000000000000001100000100000000010 : 46'b0101000000000100000000000001100000100000000000;
														assign node643 = (inp[8]) ? 46'b0101000000000010000000000000100000100000000000 : 46'b0101000000000000001000000001100000100000000000;
													assign node646 = (inp[8]) ? node650 : node647;
														assign node647 = (inp[14]) ? 46'b0100000000000000001000000001100000100000000000 : 46'b0100000000000100000000000000100000100000000000;
														assign node650 = (inp[14]) ? 46'b0100000000000010000000000000100000100000000000 : 46'b0100000000000000000000000001100000100000000010;
											assign node653 = (inp[5]) ? node669 : node654;
												assign node654 = (inp[12]) ? node662 : node655;
													assign node655 = (inp[10]) ? node659 : node656;
														assign node656 = (inp[4]) ? 46'b0101000000000000001000000001000010100000000000 : 46'b0101000000000100000000000000000010100000000000;
														assign node659 = (inp[4]) ? 46'b0101000000000010000000000001000010100000000000 : 46'b0101000000000000000000000001000010100000000010;
													assign node662 = (inp[10]) ? node666 : node663;
														assign node663 = (inp[8]) ? 46'b0101000000000000000000000001000000100000000010 : 46'b0101000000000100001000000001000000100000000000;
														assign node666 = (inp[4]) ? 46'b0101000000000010000000000000000000100000000000 : 46'b0101000000000000000000000001000000100000000010;
												assign node669 = (inp[12]) ? node677 : node670;
													assign node670 = (inp[10]) ? node674 : node671;
														assign node671 = (inp[4]) ? 46'b0100000000000000001000000001000010100000000000 : 46'b0100000000000100000000000000000010100000000000;
														assign node674 = (inp[8]) ? 46'b0100000000000010000000000001000010100000000010 : 46'b0100000000000000000000000001000010100000000010;
													assign node677 = (inp[14]) ? node681 : node678;
														assign node678 = (inp[8]) ? 46'b0100000000000000000000000001000000100000000010 : 46'b0100000000000100000000000001000000100000000000;
														assign node681 = (inp[8]) ? 46'b0100000000000010000000000000000000100000000000 : 46'b0100000000000000001000000001000000100000000000;
										assign node684 = (inp[5]) ? node716 : node685;
											assign node685 = (inp[7]) ? node701 : node686;
												assign node686 = (inp[12]) ? node694 : node687;
													assign node687 = (inp[4]) ? node691 : node688;
														assign node688 = (inp[10]) ? 46'b0101000000000000000000000001100010000000000010 : 46'b0101000000000100000000000000100010000000000000;
														assign node691 = (inp[10]) ? 46'b0101000000000010000000000000100010000000000000 : 46'b0101000000000010001000000001100010000000000000;
													assign node694 = (inp[14]) ? node698 : node695;
														assign node695 = (inp[8]) ? 46'b0101000000000000000000000001100000000000000010 : 46'b0101000000000100000000000000100000000000000000;
														assign node698 = (inp[8]) ? 46'b0101000000000010000000000000100000000000000000 : 46'b0101000000000000001000000001100000000000000000;
												assign node701 = (inp[12]) ? node709 : node702;
													assign node702 = (inp[8]) ? node706 : node703;
														assign node703 = (inp[14]) ? 46'b0101000000000000001000000001000010000000000000 : 46'b0101000000000100000000000000000010000000000000;
														assign node706 = (inp[14]) ? 46'b0101000000000010000000000000000010000000000000 : 46'b0101000000000000000000000001000010000000000010;
													assign node709 = (inp[4]) ? node713 : node710;
														assign node710 = (inp[14]) ? 46'b0101000000000000001000000001000000000000000000 : 46'b0101000000000100000000000001000000000000000010;
														assign node713 = (inp[10]) ? 46'b0101000000000010000000000000000000000000000000 : 46'b0101000000000000001000000001000000000000000000;
											assign node716 = (inp[12]) ? node732 : node717;
												assign node717 = (inp[8]) ? node725 : node718;
													assign node718 = (inp[14]) ? node722 : node719;
														assign node719 = (inp[7]) ? 46'b0100000000000100000000000001000010000000000000 : 46'b0100000000000100000000000000100010000000000000;
														assign node722 = (inp[7]) ? 46'b0100000000000000001000000001000010000000000000 : 46'b0100000000000000001000000001100010000000000000;
													assign node725 = (inp[7]) ? node729 : node726;
														assign node726 = (inp[14]) ? 46'b0100000000000010000000000000100010000000000000 : 46'b0100000000000010000000000001100010000000000010;
														assign node729 = (inp[14]) ? 46'b0100000000000010000000000000000010000000000000 : 46'b0100000000000000000000000001000010000000000010;
												assign node732 = (inp[7]) ? node740 : node733;
													assign node733 = (inp[4]) ? node737 : node734;
														assign node734 = (inp[14]) ? 46'b0100000000000110000000000000100000000000000000 : 46'b0100000000000100000000000001100000000000000010;
														assign node737 = (inp[10]) ? 46'b0100000000000010000000000000100000000000000000 : 46'b0100000000000000001000000001100000000000000000;
													assign node740 = (inp[14]) ? node744 : node741;
														assign node741 = (inp[8]) ? 46'b0100000000000000000000000001000000000000000010 : 46'b0100000000000100000000000000000000000000000000;
														assign node744 = (inp[8]) ? 46'b0100000000000010000000000000000000000000000000 : 46'b0100000000000000001000000001000000000000000000;
							assign node747 = (inp[11]) ? node797 : node748;
								assign node748 = (inp[0]) ? 46'b0000000000000000000000000000000000000000000000 : node749;
									assign node749 = (inp[5]) ? node773 : node750;
										assign node750 = (inp[7]) ? node752 : 46'b0000000000000000000000000000000000000000000000;
											assign node752 = (inp[4]) ? node766 : node753;
												assign node753 = (inp[10]) ? node761 : node754;
													assign node754 = (inp[12]) ? node758 : node755;
														assign node755 = (inp[6]) ? 46'b0001000000000100000000001000000010000000000000 : 46'b0001000000000100000000001001000010100000000000;
														assign node758 = (inp[6]) ? 46'b0001000000000100000000001000000000000000000000 : 46'b0001000000000100000000001000000000100000000000;
													assign node761 = (inp[14]) ? 46'b0000000000000000000000000000000000000000000000 : node762;
														assign node762 = (inp[8]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0001000000000100000000001001000010100000000010;
												assign node766 = (inp[8]) ? 46'b0000000000000000000000000000000000000000000000 : node767;
													assign node767 = (inp[14]) ? 46'b0000000000000000000000000000000000000000000000 : node768;
														assign node768 = (inp[12]) ? 46'b0001000000000100001000001001000000000000000000 : 46'b0001000000000110000000001000000010000000000000;
										assign node773 = (inp[7]) ? 46'b0000000000000000000000000000000000000000000000 : node774;
											assign node774 = (inp[10]) ? node782 : node775;
												assign node775 = (inp[14]) ? 46'b0000000000000000000000000000000000000000000000 : node776;
													assign node776 = (inp[8]) ? node778 : 46'b0000000000000000000000000000000000000000000000;
														assign node778 = (inp[4]) ? 46'b0000000000000000001000001001100000000000000010 : 46'b0000000000000100000000001001100000000000000010;
												assign node782 = (inp[4]) ? node790 : node783;
													assign node783 = (inp[6]) ? node787 : node784;
														assign node784 = (inp[8]) ? 46'b0000000000000010000000001001100000100000000010 : 46'b0000000000000000000000001001100010100000000010;
														assign node787 = (inp[12]) ? 46'b0000000000000000000000001001100000000000000010 : 46'b0000000000000000000000001001100010000000000010;
													assign node790 = (inp[8]) ? node792 : 46'b0000000000000000000000000000000000000000000000;
														assign node792 = (inp[14]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0000000000000010000000001001100010000000000010;
								assign node797 = (inp[0]) ? node925 : node798;
									assign node798 = (inp[7]) ? node862 : node799;
										assign node799 = (inp[6]) ? node831 : node800;
											assign node800 = (inp[12]) ? node816 : node801;
												assign node801 = (inp[5]) ? node809 : node802;
													assign node802 = (inp[8]) ? node806 : node803;
														assign node803 = (inp[14]) ? 46'b1001000000000000001000000001100010100000000000 : 46'b1001000000000100000000000000100010100000000000;
														assign node806 = (inp[14]) ? 46'b1001000000000010000000000000100010100000000000 : 46'b1001000000000000000000000001100010100000000010;
													assign node809 = (inp[14]) ? node813 : node810;
														assign node810 = (inp[8]) ? 46'b1000000000000000000000000001100010100000000010 : 46'b1000000000000100000000000000100010100000000000;
														assign node813 = (inp[8]) ? 46'b1000000000000010000000000000100010100000000000 : 46'b1000000000000000001000000001100010100000000000;
												assign node816 = (inp[5]) ? node824 : node817;
													assign node817 = (inp[8]) ? node821 : node818;
														assign node818 = (inp[10]) ? 46'b1001000000000110000000000001100000100000000000 : 46'b1001000000000100001000000001100000100000000000;
														assign node821 = (inp[10]) ? 46'b1001000000000010000000000001100000100000000010 : 46'b1001000000000110000000000000100000100000000000;
													assign node824 = (inp[10]) ? node828 : node825;
														assign node825 = (inp[4]) ? 46'b1000000000000000001000000001100000100000000000 : 46'b1000000000000100000000000000100000100000000000;
														assign node828 = (inp[4]) ? 46'b1000000000000010000000000000100000100000000000 : 46'b1000000000000000000000000001100000100000000010;
											assign node831 = (inp[12]) ? node847 : node832;
												assign node832 = (inp[5]) ? node840 : node833;
													assign node833 = (inp[8]) ? node837 : node834;
														assign node834 = (inp[14]) ? 46'b1001000000000000001000000001100010000000000000 : 46'b1001000000000100000000000000100010000000000000;
														assign node837 = (inp[14]) ? 46'b1001000000000010000000000000100010000000000000 : 46'b1001000000000000000000000001100010000000000010;
													assign node840 = (inp[14]) ? node844 : node841;
														assign node841 = (inp[8]) ? 46'b1000000000000000000000000001100010000000000010 : 46'b1000000000000100000000000000100010000000000000;
														assign node844 = (inp[8]) ? 46'b1000000000000010000000000000100010000000000000 : 46'b1000000000000000001000000001100010000000000000;
												assign node847 = (inp[5]) ? node855 : node848;
													assign node848 = (inp[4]) ? node852 : node849;
														assign node849 = (inp[10]) ? 46'b1001000000000000000000000001100000000000000010 : 46'b1001000000000100000000000000100000000000000000;
														assign node852 = (inp[10]) ? 46'b1001000000000010000000000000100000000000000000 : 46'b1001000000000000001000000001100000000000000000;
													assign node855 = (inp[14]) ? node859 : node856;
														assign node856 = (inp[8]) ? 46'b1000000000000000000000000001100000000000000010 : 46'b1000000000000100000000000000100000000000000000;
														assign node859 = (inp[10]) ? 46'b1000000000000010000000000001100000000000000000 : 46'b1000000000000000001000000001100000000000000000;
										assign node862 = (inp[12]) ? node894 : node863;
											assign node863 = (inp[6]) ? node879 : node864;
												assign node864 = (inp[5]) ? node872 : node865;
													assign node865 = (inp[10]) ? node869 : node866;
														assign node866 = (inp[14]) ? 46'b1001000000000000001000000001000010100000000000 : 46'b1001000000000100000000000001000010100000000000;
														assign node869 = (inp[4]) ? 46'b1001000000000010000000000000000010100000000000 : 46'b1001000000000000000000000001000010100000000010;
													assign node872 = (inp[10]) ? node876 : node873;
														assign node873 = (inp[4]) ? 46'b1000000000000000001000000001000010100000000000 : 46'b1000000000000100000000000000000010100000000000;
														assign node876 = (inp[4]) ? 46'b1000000000000010000000000001000010100000000000 : 46'b1000000000000000000000000001000010100000000010;
												assign node879 = (inp[4]) ? node887 : node880;
													assign node880 = (inp[10]) ? node884 : node881;
														assign node881 = (inp[5]) ? 46'b1000000000000100000000000000000010000000000000 : 46'b1001000000000100000000000000000010000000000000;
														assign node884 = (inp[5]) ? 46'b1000000000000000000000000001000010000000000010 : 46'b1001000000000000000000000001000010000000000010;
													assign node887 = (inp[10]) ? node891 : node888;
														assign node888 = (inp[14]) ? 46'b1000000000000000001000000001000010000000000000 : 46'b1000000000000000001000000001000010000000000010;
														assign node891 = (inp[5]) ? 46'b1000000000000010000000000000000010000000000000 : 46'b1001000000000010000000000001000010000000000000;
											assign node894 = (inp[6]) ? node910 : node895;
												assign node895 = (inp[5]) ? node903 : node896;
													assign node896 = (inp[4]) ? node900 : node897;
														assign node897 = (inp[10]) ? 46'b1001000000000000000000000001000000100000000010 : 46'b1001000000000100000000000000000000100000000000;
														assign node900 = (inp[10]) ? 46'b1001000000000010000000000000000000100000000000 : 46'b1001000000000000001000000001000000100000000000;
													assign node903 = (inp[4]) ? node907 : node904;
														assign node904 = (inp[14]) ? 46'b1000000000000000001000000001000000100000000000 : 46'b1000000000000100000000000001000000100000000010;
														assign node907 = (inp[14]) ? 46'b1000000000000010000000000000000000100000000000 : 46'b1000000000000010000000000000000000100000000000;
												assign node910 = (inp[5]) ? node918 : node911;
													assign node911 = (inp[8]) ? node915 : node912;
														assign node912 = (inp[14]) ? 46'b1001000000000000001000000001000000000000000000 : 46'b1001000000000100000000000000000000000000000000;
														assign node915 = (inp[14]) ? 46'b1001000000000010000000000001000000000000000000 : 46'b1001000000000000000000000001000000000000000010;
													assign node918 = (inp[8]) ? node922 : node919;
														assign node919 = (inp[14]) ? 46'b1000000000000000001000000001000000000000000000 : 46'b1000000000000100000000000000000000000000000000;
														assign node922 = (inp[14]) ? 46'b1000000000000010000000000001000000000000000000 : 46'b1000000000000000000000000001000000000000000010;
									assign node925 = (inp[5]) ? node989 : node926;
										assign node926 = (inp[6]) ? node958 : node927;
											assign node927 = (inp[7]) ? node943 : node928;
												assign node928 = (inp[12]) ? node936 : node929;
													assign node929 = (inp[14]) ? node933 : node930;
														assign node930 = (inp[4]) ? 46'b0001000000000110000000000000100010101000000000 : 46'b0001000000000100000000000000100010101000000000;
														assign node933 = (inp[8]) ? 46'b0001000000000010000000000000100010101000000000 : 46'b0001000000000000001000000001100010101000000000;
													assign node936 = (inp[4]) ? node940 : node937;
														assign node937 = (inp[10]) ? 46'b0001000000000000000000000001100000101000000010 : 46'b0001000000000100000000000000100000101000000000;
														assign node940 = (inp[10]) ? 46'b0001000000000010000000000000100000101000000000 : 46'b0001000000000000001000000001100000101000000000;
												assign node943 = (inp[12]) ? node951 : node944;
													assign node944 = (inp[10]) ? node948 : node945;
														assign node945 = (inp[4]) ? 46'b0001000000000000001000000001000010101000000000 : 46'b0001000000000100000000000000000010101000000000;
														assign node948 = (inp[4]) ? 46'b0001000000000010000000000000000010101000000000 : 46'b0001000000000000000000000001000010101000000010;
													assign node951 = (inp[10]) ? node955 : node952;
														assign node952 = (inp[4]) ? 46'b0001000000000000001000000001000000101000000000 : 46'b0001000000000100000000000000000000101000000000;
														assign node955 = (inp[8]) ? 46'b0001000000000010000000000001000000101000000010 : 46'b0001000000000000001000000001000000101000000000;
											assign node958 = (inp[7]) ? node974 : node959;
												assign node959 = (inp[12]) ? node967 : node960;
													assign node960 = (inp[10]) ? node964 : node961;
														assign node961 = (inp[4]) ? 46'b0001000000000000001000000001100010001000000000 : 46'b0001000000000100000000000000100010001000000000;
														assign node964 = (inp[4]) ? 46'b0001000000000010000000000000100010001000000000 : 46'b0001000000000000000000000001100010001000000010;
													assign node967 = (inp[14]) ? node971 : node968;
														assign node968 = (inp[4]) ? 46'b0001000000000000001000000001100000001000000010 : 46'b0001000000000100000000000001100000001000000010;
														assign node971 = (inp[8]) ? 46'b0001000000000010000000000001100000001000000000 : 46'b0001000000000000001000000001100000001000000000;
												assign node974 = (inp[12]) ? node982 : node975;
													assign node975 = (inp[14]) ? node979 : node976;
														assign node976 = (inp[10]) ? 46'b0001000000000110000000000000000010001000000000 : 46'b0001000000000100000000000001000010001000000000;
														assign node979 = (inp[8]) ? 46'b0001000000000010000000000000000010001000000000 : 46'b0001000000000000001000000001000010001000000000;
													assign node982 = (inp[10]) ? node986 : node983;
														assign node983 = (inp[4]) ? 46'b0001000000000000001000000001000000001000000000 : 46'b0001000000000100000000000000000000001000000000;
														assign node986 = (inp[4]) ? 46'b0001000000000010000000000000000000001000000000 : 46'b0001000000000010000000000001000000001000000010;
										assign node989 = (inp[7]) ? node1021 : node990;
											assign node990 = (inp[6]) ? node1006 : node991;
												assign node991 = (inp[12]) ? node999 : node992;
													assign node992 = (inp[4]) ? node996 : node993;
														assign node993 = (inp[10]) ? 46'b0000000000000000000000000001100010101000000010 : 46'b0000000000000100000000000000100010101000000000;
														assign node996 = (inp[14]) ? 46'b0000000000000010001000000001100010101000000000 : 46'b0000000000000100000000000000100010101000000000;
													assign node999 = (inp[14]) ? node1003 : node1000;
														assign node1000 = (inp[8]) ? 46'b0000000000000000000000000001100000101000000010 : 46'b0000000000000100000000000000100000101000000000;
														assign node1003 = (inp[8]) ? 46'b0000000000000010000000000000100000101000000000 : 46'b0000000000000000001000000001100000101000000000;
												assign node1006 = (inp[12]) ? node1014 : node1007;
													assign node1007 = (inp[14]) ? node1011 : node1008;
														assign node1008 = (inp[8]) ? 46'b0000000000000000000000000001100010001000000010 : 46'b0000000000000100000000000001100010001000000010;
														assign node1011 = (inp[8]) ? 46'b0000000000000010000000000000100010001000000000 : 46'b0000000000000000001000000001100010001000000000;
													assign node1014 = (inp[10]) ? node1018 : node1015;
														assign node1015 = (inp[4]) ? 46'b0000000000000000001000000001100000001000000000 : 46'b0000000000000100000000000000100000001000000000;
														assign node1018 = (inp[4]) ? 46'b0000000000000010000000000000100000001000000000 : 46'b0000000000000000000000000001100000001000000010;
											assign node1021 = (inp[12]) ? node1037 : node1022;
												assign node1022 = (inp[14]) ? node1030 : node1023;
													assign node1023 = (inp[6]) ? node1027 : node1024;
														assign node1024 = (inp[8]) ? 46'b0000000000000000000000000001000010101000000010 : 46'b0000000000000100000000000000000010101000000000;
														assign node1027 = (inp[4]) ? 46'b0000000000000100001000000001000010001000000000 : 46'b0000000000000100000000000001000010001000000010;
													assign node1030 = (inp[8]) ? node1034 : node1031;
														assign node1031 = (inp[6]) ? 46'b0000000000000000001000000001000010001000000000 : 46'b0000000000000000001000000001000010101000000000;
														assign node1034 = (inp[4]) ? 46'b0000000000000010000000000000000010001000000000 : 46'b0000000000000110000000000000000010001000000000;
												assign node1037 = (inp[6]) ? node1045 : node1038;
													assign node1038 = (inp[8]) ? node1042 : node1039;
														assign node1039 = (inp[14]) ? 46'b0000000000000000001000000001000000101000000000 : 46'b0000000000000100000000000001000000101000000000;
														assign node1042 = (inp[14]) ? 46'b0000000000000010000000000000000000101000000000 : 46'b0000000000000000000000000001000000101000000010;
													assign node1045 = (inp[10]) ? node1049 : node1046;
														assign node1046 = (inp[4]) ? 46'b0000000000000000001000000001000000001000000000 : 46'b0000000000000100000000000000000000001000000000;
														assign node1049 = (inp[4]) ? 46'b0000000000000010000000000000000000001000000000 : 46'b0000000000000000000000000001000000001000000010;
						assign node1052 = (inp[11]) ? node1390 : node1053;
							assign node1053 = (inp[9]) ? node1135 : node1054;
								assign node1054 = (inp[7]) ? node1070 : node1055;
									assign node1055 = (inp[12]) ? node1057 : 46'b0000000000000000000000000000000000000000000000;
										assign node1057 = (inp[5]) ? node1059 : 46'b0000000000000000000000000000000000000000000000;
											assign node1059 = (inp[6]) ? node1061 : 46'b0000000000000000000000000000000000000000000000;
												assign node1061 = (inp[0]) ? node1063 : 46'b0000000000000000000000000000000000000000000000;
													assign node1063 = (inp[8]) ? node1067 : node1064;
														assign node1064 = (inp[14]) ? 46'b0000000000000001001000000001100000000000100010 : 46'b0000000000000101000000000000100000000000100000;
														assign node1067 = (inp[14]) ? 46'b0000000000000011000000000001100000000000100000 : 46'b0000000000000001000000000001100000000000100010;
									assign node1070 = (inp[5]) ? node1084 : node1071;
										assign node1071 = (inp[0]) ? node1073 : 46'b0000000000000000000000000000000000000000000000;
											assign node1073 = (inp[6]) ? node1075 : 46'b0000000000000000000000000000000000000000000000;
												assign node1075 = (inp[12]) ? node1077 : 46'b0000000000000000000000000000000000000000000000;
													assign node1077 = (inp[8]) ? node1081 : node1078;
														assign node1078 = (inp[14]) ? 46'b0001000000000001001000000001000000000000100000 : 46'b0001000000000101000000000000000000000000100000;
														assign node1081 = (inp[14]) ? 46'b0001000000000011000000000000000000000000100000 : 46'b0001000000000001000000000001000000000000100010;
										assign node1084 = (inp[0]) ? node1116 : node1085;
											assign node1085 = (inp[6]) ? node1101 : node1086;
												assign node1086 = (inp[12]) ? node1094 : node1087;
													assign node1087 = (inp[8]) ? node1091 : node1088;
														assign node1088 = (inp[14]) ? 46'b0000000000100000001001000001000010100000000000 : 46'b0000000000100100000001000000000010100000000000;
														assign node1091 = (inp[14]) ? 46'b0000000000100010000001000000000010100000000000 : 46'b0000000000100000000001000001000010100000000010;
													assign node1094 = (inp[14]) ? node1098 : node1095;
														assign node1095 = (inp[8]) ? 46'b0000000000100000000001000001000000100000000010 : 46'b0000000000100100000001000000000000100000000000;
														assign node1098 = (inp[4]) ? 46'b0000000000100010001001000001000000100000000000 : 46'b0000000000100000001001000001000000100000000010;
												assign node1101 = (inp[12]) ? node1109 : node1102;
													assign node1102 = (inp[14]) ? node1106 : node1103;
														assign node1103 = (inp[4]) ? 46'b0000000000100000001001000001000010000000000000 : 46'b0000000000100100000001000001000010000000000010;
														assign node1106 = (inp[4]) ? 46'b0000000000100010001001000001000010000000000000 : 46'b0000000000100000001001000001000010000000000000;
													assign node1109 = (inp[8]) ? node1113 : node1110;
														assign node1110 = (inp[14]) ? 46'b0000000000100000001001000001000000000000000000 : 46'b0000000000100100000001000000000000000000000000;
														assign node1113 = (inp[14]) ? 46'b0000000000100010000001000001000000000000000000 : 46'b0000000000100000000001000001000000000000000010;
											assign node1116 = (inp[12]) ? node1126 : node1117;
												assign node1117 = (inp[6]) ? node1119 : 46'b0000000000000000000000000000000000000000000000;
													assign node1119 = (inp[8]) ? node1123 : node1120;
														assign node1120 = (inp[10]) ? 46'b0000000000000001000000000001000010000000100010 : 46'b0000000000000101001000000001000010000000100000;
														assign node1123 = (inp[14]) ? 46'b0000000000000011000000000000000010000000100000 : 46'b0000000000000001000000000001000010000000100010;
												assign node1126 = (inp[6]) ? 46'b0000000000000000000000000000000000000000000000 : node1127;
													assign node1127 = (inp[14]) ? node1131 : node1128;
														assign node1128 = (inp[8]) ? 46'b0000000000000001000000000001000000100000100010 : 46'b0000000000000101000000000000000000100000100000;
														assign node1131 = (inp[4]) ? 46'b0000000000000011001000000001000000100000100000 : 46'b0000000000000101001000000001000000100000100000;
								assign node1135 = (inp[7]) ? node1263 : node1136;
									assign node1136 = (inp[6]) ? node1200 : node1137;
										assign node1137 = (inp[12]) ? node1169 : node1138;
											assign node1138 = (inp[0]) ? node1154 : node1139;
												assign node1139 = (inp[5]) ? node1147 : node1140;
													assign node1140 = (inp[10]) ? node1144 : node1141;
														assign node1141 = (inp[4]) ? 46'b0001000000100000001000000001100010100000100000 : 46'b0001000000100100000000000000100010100000100000;
														assign node1144 = (inp[4]) ? 46'b0001000000100010000000000001100010100000100000 : 46'b0001000000100000000000000001100010100000100010;
													assign node1147 = (inp[4]) ? node1151 : node1148;
														assign node1148 = (inp[10]) ? 46'b0000000000100000000000000001100010100000100010 : 46'b0000000000100100000000000000100010100000100000;
														assign node1151 = (inp[10]) ? 46'b0000000000100010000000000000100010100000100000 : 46'b0000000000100000001000000001100010100000100000;
												assign node1154 = (inp[5]) ? node1162 : node1155;
													assign node1155 = (inp[4]) ? node1159 : node1156;
														assign node1156 = (inp[10]) ? 46'b0001000000000000000000000001100010100000100010 : 46'b0001000000000100000000000000100010100000100000;
														assign node1159 = (inp[14]) ? 46'b0001000000000010001000000001100010100000100000 : 46'b0001000000000100000000000000100010100000100000;
													assign node1162 = (inp[14]) ? node1166 : node1163;
														assign node1163 = (inp[8]) ? 46'b0000000000000000000000000001100010100000100010 : 46'b0000000000000100000000000000100010100000100000;
														assign node1166 = (inp[8]) ? 46'b0000000000000010000000000000100010100000100000 : 46'b0000000000000000001000000001100010100000100000;
											assign node1169 = (inp[5]) ? node1185 : node1170;
												assign node1170 = (inp[0]) ? node1178 : node1171;
													assign node1171 = (inp[14]) ? node1175 : node1172;
														assign node1172 = (inp[8]) ? 46'b0001000000100000000000000001100000100000100010 : 46'b0001000000100100000000000001100000100000100000;
														assign node1175 = (inp[8]) ? 46'b0001000000100010000000000000100000100000100000 : 46'b0001000000100000001000000001100000100000100000;
													assign node1178 = (inp[4]) ? node1182 : node1179;
														assign node1179 = (inp[10]) ? 46'b0001000000000000000000000001100000100000100010 : 46'b0001000000000100000000000000100000100000100000;
														assign node1182 = (inp[14]) ? 46'b0001000000000010001000000001100000100000100000 : 46'b0001000000000110000000000000100000100000100000;
												assign node1185 = (inp[0]) ? node1193 : node1186;
													assign node1186 = (inp[10]) ? node1190 : node1187;
														assign node1187 = (inp[4]) ? 46'b0000000000100000001000000001100000100000100000 : 46'b0000000000100100000000000000100000100000100000;
														assign node1190 = (inp[4]) ? 46'b0000000000100010000000000001100000100000100000 : 46'b0000000000100000000000000001100000100000100010;
													assign node1193 = (inp[10]) ? node1197 : node1194;
														assign node1194 = (inp[4]) ? 46'b0000000000000000001000000001100000100000100000 : 46'b0000000000000100000000000000100000100000100000;
														assign node1197 = (inp[4]) ? 46'b0000000000000010000000000001100000100000100000 : 46'b0000000000000000000000000001100000100000100010;
										assign node1200 = (inp[5]) ? node1232 : node1201;
											assign node1201 = (inp[12]) ? node1217 : node1202;
												assign node1202 = (inp[0]) ? node1210 : node1203;
													assign node1203 = (inp[4]) ? node1207 : node1204;
														assign node1204 = (inp[10]) ? 46'b0001000000100000000000000001100010000000100010 : 46'b0001000000100100000000000001100010000000100000;
														assign node1207 = (inp[10]) ? 46'b0001000000100010000000000000100010000000100000 : 46'b0001000000100000001000000001100010000000100000;
													assign node1210 = (inp[10]) ? node1214 : node1211;
														assign node1211 = (inp[4]) ? 46'b0001000000000000001000000001100010000000100000 : 46'b0001000000000100000000000000100010000000100000;
														assign node1214 = (inp[4]) ? 46'b0001000000000010000000000001100010000000100000 : 46'b0001000000000000000000000001100010000000100010;
												assign node1217 = (inp[0]) ? node1225 : node1218;
													assign node1218 = (inp[8]) ? node1222 : node1219;
														assign node1219 = (inp[14]) ? 46'b0001000000100000001000000001100000000000100000 : 46'b0001000000100100000000000001100000000000100000;
														assign node1222 = (inp[14]) ? 46'b0001000000100010000000000000100000000000100000 : 46'b0001000000100000000000000001100000000000100010;
													assign node1225 = (inp[14]) ? node1229 : node1226;
														assign node1226 = (inp[4]) ? 46'b0001000000000000001000000001100000000000100010 : 46'b0001000000000100000000000001100000000000100010;
														assign node1229 = (inp[8]) ? 46'b0001000000000010000000000000100000000000100000 : 46'b0001000000000000001000000001100000000000100000;
											assign node1232 = (inp[0]) ? node1248 : node1233;
												assign node1233 = (inp[12]) ? node1241 : node1234;
													assign node1234 = (inp[10]) ? node1238 : node1235;
														assign node1235 = (inp[8]) ? 46'b0000000000100000000000000001100010000000100010 : 46'b0000000000100100001000000001100010000000100000;
														assign node1238 = (inp[4]) ? 46'b0000000000100010000000000000100010000000100000 : 46'b0000000000100000000000000001100010000000100010;
													assign node1241 = (inp[14]) ? node1245 : node1242;
														assign node1242 = (inp[8]) ? 46'b0000000000100000000000000001100000000000100010 : 46'b0000000000100100000000000000100000000000100000;
														assign node1245 = (inp[4]) ? 46'b0000000000100010001000000001100000000000100000 : 46'b0000000000100000000000000001100000000000100010;
												assign node1248 = (inp[12]) ? node1256 : node1249;
													assign node1249 = (inp[8]) ? node1253 : node1250;
														assign node1250 = (inp[14]) ? 46'b0000000000000000001000000001100010000000100000 : 46'b0000000000000100000000000000100010000000100000;
														assign node1253 = (inp[14]) ? 46'b0000000000000010000000000001100010000000100000 : 46'b0000000000000000000000000001100010000000100010;
													assign node1256 = (inp[8]) ? node1260 : node1257;
														assign node1257 = (inp[14]) ? 46'b0000000000000000001000000001100000000000100000 : 46'b0000000000000100000000000000100000000000100000;
														assign node1260 = (inp[10]) ? 46'b0000000000000010000000000001100000000000100010 : 46'b0000000000000000000000000001100000000000100010;
									assign node1263 = (inp[12]) ? node1327 : node1264;
										assign node1264 = (inp[0]) ? node1296 : node1265;
											assign node1265 = (inp[6]) ? node1281 : node1266;
												assign node1266 = (inp[5]) ? node1274 : node1267;
													assign node1267 = (inp[14]) ? node1271 : node1268;
														assign node1268 = (inp[4]) ? 46'b0001000000100000001000000001000010100000100000 : 46'b0001000000100100000000000001000010100000100010;
														assign node1271 = (inp[8]) ? 46'b0001000000100010000000000000000010100000100000 : 46'b0001000000100000001000000001000010100000100000;
													assign node1274 = (inp[14]) ? node1278 : node1275;
														assign node1275 = (inp[8]) ? 46'b0000000000100000000000000001000010100000100010 : 46'b0000000000100100000000000001000010100000100000;
														assign node1278 = (inp[8]) ? 46'b0000000000100010000000000000000010100000100000 : 46'b0000000000100000001000000001000010100000100000;
												assign node1281 = (inp[5]) ? node1289 : node1282;
													assign node1282 = (inp[14]) ? node1286 : node1283;
														assign node1283 = (inp[8]) ? 46'b0001000000100000000000000001000010000000100010 : 46'b0001000000100100000000000000000010000000100000;
														assign node1286 = (inp[8]) ? 46'b0001000000100010000000000000000010000000100000 : 46'b0001000000100000001000000001000010000000100000;
													assign node1289 = (inp[10]) ? node1293 : node1290;
														assign node1290 = (inp[8]) ? 46'b0000000000100000001000000001000010000000100000 : 46'b0000000000100100001000000001000010000000100000;
														assign node1293 = (inp[4]) ? 46'b0000000000100010000000000000000010000000100000 : 46'b0000000000100000000000000001000010000000100010;
											assign node1296 = (inp[5]) ? node1312 : node1297;
												assign node1297 = (inp[6]) ? node1305 : node1298;
													assign node1298 = (inp[14]) ? node1302 : node1299;
														assign node1299 = (inp[8]) ? 46'b0001000000000000000000000001000010100000100010 : 46'b0001000000000100000000000000000010100000100000;
														assign node1302 = (inp[8]) ? 46'b0001000000000010000000000000000010100000100000 : 46'b0001000000000000001000000001000010100000100000;
													assign node1305 = (inp[4]) ? node1309 : node1306;
														assign node1306 = (inp[14]) ? 46'b0001000000000000000000000001000010000000100010 : 46'b0001000000000100000000000001000010000000100010;
														assign node1309 = (inp[8]) ? 46'b0001000000000000001000000001000010000000100000 : 46'b0001000000000010000000000000000010000000100000;
												assign node1312 = (inp[6]) ? node1320 : node1313;
													assign node1313 = (inp[10]) ? node1317 : node1314;
														assign node1314 = (inp[4]) ? 46'b0000000000000000001000000001000010100000100000 : 46'b0000000000000100000000000000000010100000100000;
														assign node1317 = (inp[4]) ? 46'b0000000000000010000000000000000010100000100000 : 46'b0000000000000000001000000001000010100000100010;
													assign node1320 = (inp[4]) ? node1324 : node1321;
														assign node1321 = (inp[10]) ? 46'b0000000000000000000000000001000010000000100010 : 46'b0000000000000100000000000000000010000000100000;
														assign node1324 = (inp[8]) ? 46'b0000000000000010000000000001000010000000100000 : 46'b0000000000000110000000000000000010000000100000;
										assign node1327 = (inp[0]) ? node1359 : node1328;
											assign node1328 = (inp[6]) ? node1344 : node1329;
												assign node1329 = (inp[5]) ? node1337 : node1330;
													assign node1330 = (inp[10]) ? node1334 : node1331;
														assign node1331 = (inp[4]) ? 46'b0001000000100000001000000001000000100000100000 : 46'b0001000000100100000000000000000000100000100000;
														assign node1334 = (inp[8]) ? 46'b0001000000100010000000000001000000100000100010 : 46'b0001000000100100000000000001000000100000100010;
													assign node1337 = (inp[4]) ? node1341 : node1338;
														assign node1338 = (inp[14]) ? 46'b0000000000100000001000000001000000100000100000 : 46'b0000000000100100000000000001000000100000100010;
														assign node1341 = (inp[10]) ? 46'b0000000000100010000000000000000000100000100000 : 46'b0000000000100000001000000001000000100000100000;
												assign node1344 = (inp[5]) ? node1352 : node1345;
													assign node1345 = (inp[10]) ? node1349 : node1346;
														assign node1346 = (inp[8]) ? 46'b0001000000100100000000000000000000000000100000 : 46'b0001000000100100001000000001000000000000100000;
														assign node1349 = (inp[4]) ? 46'b0001000000100010000000000000000000000000100000 : 46'b0001000000100000000000000001000000000000100010;
													assign node1352 = (inp[10]) ? node1356 : node1353;
														assign node1353 = (inp[4]) ? 46'b0000000000100100001000000001000000000000100000 : 46'b0000000000100100000000000000000000000000100000;
														assign node1356 = (inp[8]) ? 46'b0000000000100010000000000001000000000000100010 : 46'b0000000000100110000000000001000000000000100000;
											assign node1359 = (inp[5]) ? node1375 : node1360;
												assign node1360 = (inp[6]) ? node1368 : node1361;
													assign node1361 = (inp[4]) ? node1365 : node1362;
														assign node1362 = (inp[10]) ? 46'b0001000000000000000000000001000000100000100010 : 46'b0001000000000100000000000000000000100000100000;
														assign node1365 = (inp[10]) ? 46'b0001000000000010000000000000000000100000100000 : 46'b0001000000000000001000000001000000100000100000;
													assign node1368 = (inp[4]) ? node1372 : node1369;
														assign node1369 = (inp[10]) ? 46'b0001000000000000000000000001000000000000100010 : 46'b0001000000000100000000000000000000000000100000;
														assign node1372 = (inp[10]) ? 46'b0001000000000010000000000000000000000000100000 : 46'b0001000000000000001000000001000000000000100000;
												assign node1375 = (inp[6]) ? node1383 : node1376;
													assign node1376 = (inp[10]) ? node1380 : node1377;
														assign node1377 = (inp[4]) ? 46'b0000000000000000001000000001000000100000100000 : 46'b0000000000000100000000000000000000100000100000;
														assign node1380 = (inp[4]) ? 46'b0000000000000010000000000001000000100000100000 : 46'b0000000000000000000000000001000000100000100010;
													assign node1383 = (inp[8]) ? node1387 : node1384;
														assign node1384 = (inp[14]) ? 46'b0000000000000000001000000001000000000000100000 : 46'b0000000000000100000000000000000000000000100000;
														assign node1387 = (inp[14]) ? 46'b0000000000000010000000000000000000000000100000 : 46'b0000000000000000000000000001000000000000100010;
							assign node1390 = (inp[7]) ? node1428 : node1391;
								assign node1391 = (inp[5]) ? node1403 : node1392;
									assign node1392 = (inp[0]) ? 46'b0000000000000000000000000000000000000000000000 : node1393;
										assign node1393 = (inp[9]) ? 46'b0000000000000000000000000000000000000000000000 : node1394;
											assign node1394 = (inp[6]) ? node1398 : node1395;
												assign node1395 = (inp[12]) ? 46'b0001000000100000001000000001100000100000100000 : 46'b0000000000000000000000000000000000000000000000;
												assign node1398 = (inp[12]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0001000000100010000000000000100010000000100000;
									assign node1403 = (inp[0]) ? node1419 : node1404;
										assign node1404 = (inp[9]) ? node1412 : node1405;
											assign node1405 = (inp[6]) ? node1409 : node1406;
												assign node1406 = (inp[12]) ? 46'b0000000000100000001000000001100000100000100000 : 46'b0000000000000000000000000000000000000000000000;
												assign node1409 = (inp[12]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0000000000100010000000000000100010000000100000;
											assign node1412 = (inp[12]) ? node1416 : node1413;
												assign node1413 = (inp[6]) ? 46'b0000000010000000000000000001100010000001000010 : 46'b0000000010000000000000000001100010100001000010;
												assign node1416 = (inp[6]) ? 46'b0000000010000000000000000001100000000001000010 : 46'b0000000010000000000000000001100000100001000010;
										assign node1419 = (inp[9]) ? 46'b0000000000000000000000000000000000000000000000 : node1420;
											assign node1420 = (inp[6]) ? node1424 : node1421;
												assign node1421 = (inp[12]) ? 46'b0000000010000000000000000001100000100000000010 : 46'b0000000010000000000000000001100010100000000010;
												assign node1424 = (inp[12]) ? 46'b0000000010000000000000000001100000000000000010 : 46'b0000000010000000000000000001100010000000000010;
								assign node1428 = (inp[5]) ? node1454 : node1429;
									assign node1429 = (inp[0]) ? node1445 : node1430;
										assign node1430 = (inp[9]) ? node1438 : node1431;
											assign node1431 = (inp[6]) ? node1435 : node1432;
												assign node1432 = (inp[12]) ? 46'b0001000000100000001000000001000000100000100000 : 46'b0000000000000000000000000000000000000000000000;
												assign node1435 = (inp[12]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0001000000100010000000000000000010000000100000;
											assign node1438 = (inp[12]) ? node1442 : node1439;
												assign node1439 = (inp[6]) ? 46'b0001000010000100000000000000000010000001000000 : 46'b0001000010000100000000000000000010100001000000;
												assign node1442 = (inp[6]) ? 46'b0001000010000100000000000000000000000001000000 : 46'b0001000010000100000000000000000000100001000000;
										assign node1445 = (inp[9]) ? 46'b0000000000000000000000000000000000000000000000 : node1446;
											assign node1446 = (inp[12]) ? node1450 : node1447;
												assign node1447 = (inp[6]) ? 46'b0001000010000100000000000000000010000000000000 : 46'b0001000010000100000000000000000010100000000000;
												assign node1450 = (inp[6]) ? 46'b0001000010000100000000000000000000000000000000 : 46'b0001000010000100000000000000000000100000000000;
									assign node1454 = (inp[0]) ? 46'b0000000000000000000000000000000000000000000000 : node1455;
										assign node1455 = (inp[9]) ? 46'b0000000000000000000000000000000000000000000000 : node1456;
											assign node1456 = (inp[6]) ? node1460 : node1457;
												assign node1457 = (inp[12]) ? 46'b0000000000100000001000000001000000100000100000 : 46'b0000000000000000000000000000000000000000000000;
												assign node1460 = (inp[12]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0000000000100010000000000000000010000000100000;

endmodule