module dtc_split875_bm71 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node7;
	wire [3-1:0] node8;
	wire [3-1:0] node9;
	wire [3-1:0] node10;
	wire [3-1:0] node14;
	wire [3-1:0] node17;
	wire [3-1:0] node19;
	wire [3-1:0] node21;
	wire [3-1:0] node22;
	wire [3-1:0] node26;
	wire [3-1:0] node27;
	wire [3-1:0] node28;
	wire [3-1:0] node29;
	wire [3-1:0] node30;
	wire [3-1:0] node35;
	wire [3-1:0] node37;
	wire [3-1:0] node40;
	wire [3-1:0] node41;
	wire [3-1:0] node42;
	wire [3-1:0] node46;
	wire [3-1:0] node48;
	wire [3-1:0] node51;
	wire [3-1:0] node52;
	wire [3-1:0] node53;
	wire [3-1:0] node55;
	wire [3-1:0] node56;
	wire [3-1:0] node60;
	wire [3-1:0] node62;
	wire [3-1:0] node63;
	wire [3-1:0] node65;
	wire [3-1:0] node69;
	wire [3-1:0] node71;
	wire [3-1:0] node73;
	wire [3-1:0] node74;
	wire [3-1:0] node76;
	wire [3-1:0] node80;
	wire [3-1:0] node81;
	wire [3-1:0] node82;
	wire [3-1:0] node83;
	wire [3-1:0] node84;
	wire [3-1:0] node85;
	wire [3-1:0] node91;
	wire [3-1:0] node92;
	wire [3-1:0] node93;
	wire [3-1:0] node94;
	wire [3-1:0] node98;
	wire [3-1:0] node100;
	wire [3-1:0] node103;
	wire [3-1:0] node104;
	wire [3-1:0] node105;
	wire [3-1:0] node107;
	wire [3-1:0] node113;
	wire [3-1:0] node114;
	wire [3-1:0] node115;
	wire [3-1:0] node116;
	wire [3-1:0] node117;
	wire [3-1:0] node118;
	wire [3-1:0] node119;
	wire [3-1:0] node123;
	wire [3-1:0] node125;
	wire [3-1:0] node128;
	wire [3-1:0] node129;
	wire [3-1:0] node132;
	wire [3-1:0] node134;
	wire [3-1:0] node137;
	wire [3-1:0] node138;
	wire [3-1:0] node139;
	wire [3-1:0] node140;
	wire [3-1:0] node144;
	wire [3-1:0] node146;
	wire [3-1:0] node148;
	wire [3-1:0] node151;
	wire [3-1:0] node152;
	wire [3-1:0] node155;
	wire [3-1:0] node157;
	wire [3-1:0] node159;
	wire [3-1:0] node162;
	wire [3-1:0] node163;
	wire [3-1:0] node164;
	wire [3-1:0] node166;
	wire [3-1:0] node167;
	wire [3-1:0] node169;
	wire [3-1:0] node173;
	wire [3-1:0] node175;
	wire [3-1:0] node178;
	wire [3-1:0] node179;
	wire [3-1:0] node180;
	wire [3-1:0] node181;
	wire [3-1:0] node182;
	wire [3-1:0] node187;
	wire [3-1:0] node190;
	wire [3-1:0] node191;
	wire [3-1:0] node192;
	wire [3-1:0] node193;
	wire [3-1:0] node198;
	wire [3-1:0] node200;
	wire [3-1:0] node201;
	wire [3-1:0] node205;
	wire [3-1:0] node206;
	wire [3-1:0] node207;
	wire [3-1:0] node208;
	wire [3-1:0] node209;
	wire [3-1:0] node210;
	wire [3-1:0] node212;
	wire [3-1:0] node216;
	wire [3-1:0] node218;
	wire [3-1:0] node220;
	wire [3-1:0] node223;
	wire [3-1:0] node224;
	wire [3-1:0] node227;
	wire [3-1:0] node229;
	wire [3-1:0] node231;
	wire [3-1:0] node234;
	wire [3-1:0] node235;
	wire [3-1:0] node236;
	wire [3-1:0] node240;
	wire [3-1:0] node241;
	wire [3-1:0] node245;
	wire [3-1:0] node246;
	wire [3-1:0] node247;
	wire [3-1:0] node249;
	wire [3-1:0] node253;
	wire [3-1:0] node254;
	wire [3-1:0] node255;
	wire [3-1:0] node256;
	wire [3-1:0] node257;
	wire [3-1:0] node262;
	wire [3-1:0] node264;
	wire [3-1:0] node265;
	wire [3-1:0] node269;
	wire [3-1:0] node270;
	wire [3-1:0] node271;
	wire [3-1:0] node275;
	wire [3-1:0] node277;
	wire [3-1:0] node278;
	wire [3-1:0] node282;
	wire [3-1:0] node283;
	wire [3-1:0] node284;
	wire [3-1:0] node285;
	wire [3-1:0] node286;
	wire [3-1:0] node288;
	wire [3-1:0] node289;
	wire [3-1:0] node291;
	wire [3-1:0] node298;
	wire [3-1:0] node299;
	wire [3-1:0] node300;
	wire [3-1:0] node301;
	wire [3-1:0] node302;
	wire [3-1:0] node303;
	wire [3-1:0] node305;
	wire [3-1:0] node308;
	wire [3-1:0] node309;
	wire [3-1:0] node310;
	wire [3-1:0] node315;
	wire [3-1:0] node317;
	wire [3-1:0] node318;
	wire [3-1:0] node322;
	wire [3-1:0] node323;
	wire [3-1:0] node325;
	wire [3-1:0] node326;
	wire [3-1:0] node330;
	wire [3-1:0] node332;
	wire [3-1:0] node333;
	wire [3-1:0] node337;
	wire [3-1:0] node338;
	wire [3-1:0] node339;
	wire [3-1:0] node340;
	wire [3-1:0] node345;
	wire [3-1:0] node346;
	wire [3-1:0] node347;
	wire [3-1:0] node349;
	wire [3-1:0] node353;
	wire [3-1:0] node354;
	wire [3-1:0] node356;
	wire [3-1:0] node360;
	wire [3-1:0] node362;
	wire [3-1:0] node363;
	wire [3-1:0] node364;
	wire [3-1:0] node366;
	wire [3-1:0] node367;
	wire [3-1:0] node373;
	wire [3-1:0] node374;
	wire [3-1:0] node376;
	wire [3-1:0] node377;
	wire [3-1:0] node378;
	wire [3-1:0] node379;
	wire [3-1:0] node380;
	wire [3-1:0] node381;
	wire [3-1:0] node386;
	wire [3-1:0] node387;
	wire [3-1:0] node388;
	wire [3-1:0] node390;
	wire [3-1:0] node391;
	wire [3-1:0] node396;
	wire [3-1:0] node397;
	wire [3-1:0] node399;
	wire [3-1:0] node403;
	wire [3-1:0] node404;
	wire [3-1:0] node405;
	wire [3-1:0] node407;
	wire [3-1:0] node408;
	wire [3-1:0] node416;
	wire [3-1:0] node417;
	wire [3-1:0] node418;
	wire [3-1:0] node419;
	wire [3-1:0] node420;
	wire [3-1:0] node421;
	wire [3-1:0] node422;
	wire [3-1:0] node423;
	wire [3-1:0] node424;
	wire [3-1:0] node428;
	wire [3-1:0] node429;
	wire [3-1:0] node431;
	wire [3-1:0] node435;
	wire [3-1:0] node437;
	wire [3-1:0] node438;
	wire [3-1:0] node440;
	wire [3-1:0] node444;
	wire [3-1:0] node445;
	wire [3-1:0] node446;
	wire [3-1:0] node447;
	wire [3-1:0] node448;
	wire [3-1:0] node449;
	wire [3-1:0] node454;
	wire [3-1:0] node456;
	wire [3-1:0] node457;
	wire [3-1:0] node461;
	wire [3-1:0] node462;
	wire [3-1:0] node463;
	wire [3-1:0] node467;
	wire [3-1:0] node469;
	wire [3-1:0] node472;
	wire [3-1:0] node473;
	wire [3-1:0] node474;
	wire [3-1:0] node475;
	wire [3-1:0] node479;
	wire [3-1:0] node481;
	wire [3-1:0] node484;
	wire [3-1:0] node485;
	wire [3-1:0] node486;
	wire [3-1:0] node490;
	wire [3-1:0] node492;
	wire [3-1:0] node495;
	wire [3-1:0] node496;
	wire [3-1:0] node497;
	wire [3-1:0] node498;
	wire [3-1:0] node499;
	wire [3-1:0] node501;
	wire [3-1:0] node502;
	wire [3-1:0] node507;
	wire [3-1:0] node508;
	wire [3-1:0] node510;
	wire [3-1:0] node514;
	wire [3-1:0] node515;
	wire [3-1:0] node516;
	wire [3-1:0] node518;
	wire [3-1:0] node519;
	wire [3-1:0] node524;
	wire [3-1:0] node525;
	wire [3-1:0] node527;
	wire [3-1:0] node531;
	wire [3-1:0] node532;
	wire [3-1:0] node533;
	wire [3-1:0] node534;
	wire [3-1:0] node535;
	wire [3-1:0] node539;
	wire [3-1:0] node541;
	wire [3-1:0] node544;
	wire [3-1:0] node545;
	wire [3-1:0] node546;
	wire [3-1:0] node548;
	wire [3-1:0] node552;
	wire [3-1:0] node554;
	wire [3-1:0] node557;
	wire [3-1:0] node558;
	wire [3-1:0] node559;
	wire [3-1:0] node560;
	wire [3-1:0] node562;
	wire [3-1:0] node566;
	wire [3-1:0] node568;
	wire [3-1:0] node571;
	wire [3-1:0] node572;
	wire [3-1:0] node575;
	wire [3-1:0] node577;
	wire [3-1:0] node579;
	wire [3-1:0] node582;
	wire [3-1:0] node583;
	wire [3-1:0] node584;
	wire [3-1:0] node586;
	wire [3-1:0] node587;
	wire [3-1:0] node589;
	wire [3-1:0] node591;
	wire [3-1:0] node593;
	wire [3-1:0] node596;
	wire [3-1:0] node597;
	wire [3-1:0] node602;
	wire [3-1:0] node603;
	wire [3-1:0] node604;
	wire [3-1:0] node605;
	wire [3-1:0] node606;
	wire [3-1:0] node608;
	wire [3-1:0] node610;
	wire [3-1:0] node614;
	wire [3-1:0] node615;
	wire [3-1:0] node617;
	wire [3-1:0] node620;
	wire [3-1:0] node621;
	wire [3-1:0] node622;
	wire [3-1:0] node627;
	wire [3-1:0] node629;
	wire [3-1:0] node631;
	wire [3-1:0] node632;
	wire [3-1:0] node636;
	wire [3-1:0] node637;
	wire [3-1:0] node638;
	wire [3-1:0] node639;
	wire [3-1:0] node643;
	wire [3-1:0] node644;
	wire [3-1:0] node648;
	wire [3-1:0] node649;
	wire [3-1:0] node650;
	wire [3-1:0] node654;
	wire [3-1:0] node655;
	wire [3-1:0] node657;
	wire [3-1:0] node658;
	wire [3-1:0] node663;
	wire [3-1:0] node664;
	wire [3-1:0] node665;
	wire [3-1:0] node666;
	wire [3-1:0] node667;
	wire [3-1:0] node668;
	wire [3-1:0] node670;
	wire [3-1:0] node671;
	wire [3-1:0] node675;
	wire [3-1:0] node677;
	wire [3-1:0] node678;
	wire [3-1:0] node682;
	wire [3-1:0] node683;
	wire [3-1:0] node685;
	wire [3-1:0] node686;
	wire [3-1:0] node688;
	wire [3-1:0] node692;
	wire [3-1:0] node694;
	wire [3-1:0] node697;
	wire [3-1:0] node698;
	wire [3-1:0] node699;
	wire [3-1:0] node700;
	wire [3-1:0] node702;
	wire [3-1:0] node706;
	wire [3-1:0] node707;
	wire [3-1:0] node709;
	wire [3-1:0] node712;
	wire [3-1:0] node713;
	wire [3-1:0] node717;
	wire [3-1:0] node718;
	wire [3-1:0] node719;
	wire [3-1:0] node721;
	wire [3-1:0] node725;
	wire [3-1:0] node726;
	wire [3-1:0] node728;
	wire [3-1:0] node730;
	wire [3-1:0] node733;
	wire [3-1:0] node734;
	wire [3-1:0] node735;
	wire [3-1:0] node740;
	wire [3-1:0] node741;
	wire [3-1:0] node742;
	wire [3-1:0] node743;
	wire [3-1:0] node745;
	wire [3-1:0] node746;
	wire [3-1:0] node748;
	wire [3-1:0] node752;
	wire [3-1:0] node754;
	wire [3-1:0] node757;
	wire [3-1:0] node758;
	wire [3-1:0] node760;
	wire [3-1:0] node763;
	wire [3-1:0] node764;
	wire [3-1:0] node765;
	wire [3-1:0] node766;
	wire [3-1:0] node771;
	wire [3-1:0] node773;
	wire [3-1:0] node774;
	wire [3-1:0] node778;
	wire [3-1:0] node779;
	wire [3-1:0] node780;
	wire [3-1:0] node781;
	wire [3-1:0] node783;
	wire [3-1:0] node785;
	wire [3-1:0] node788;
	wire [3-1:0] node789;
	wire [3-1:0] node790;
	wire [3-1:0] node796;
	wire [3-1:0] node797;
	wire [3-1:0] node799;
	wire [3-1:0] node800;
	wire [3-1:0] node801;
	wire [3-1:0] node806;
	wire [3-1:0] node808;
	wire [3-1:0] node809;
	wire [3-1:0] node813;
	wire [3-1:0] node814;
	wire [3-1:0] node815;
	wire [3-1:0] node816;
	wire [3-1:0] node817;
	wire [3-1:0] node818;
	wire [3-1:0] node819;
	wire [3-1:0] node820;
	wire [3-1:0] node825;
	wire [3-1:0] node828;
	wire [3-1:0] node829;
	wire [3-1:0] node830;
	wire [3-1:0] node831;
	wire [3-1:0] node836;
	wire [3-1:0] node838;
	wire [3-1:0] node839;
	wire [3-1:0] node843;
	wire [3-1:0] node844;
	wire [3-1:0] node846;
	wire [3-1:0] node848;
	wire [3-1:0] node849;
	wire [3-1:0] node853;
	wire [3-1:0] node854;
	wire [3-1:0] node855;
	wire [3-1:0] node859;
	wire [3-1:0] node861;
	wire [3-1:0] node864;
	wire [3-1:0] node865;
	wire [3-1:0] node866;
	wire [3-1:0] node868;
	wire [3-1:0] node869;
	wire [3-1:0] node873;
	wire [3-1:0] node875;
	wire [3-1:0] node876;
	wire [3-1:0] node880;
	wire [3-1:0] node881;
	wire [3-1:0] node883;
	wire [3-1:0] node884;
	wire [3-1:0] node888;
	wire [3-1:0] node890;
	wire [3-1:0] node891;
	wire [3-1:0] node895;
	wire [3-1:0] node896;
	wire [3-1:0] node897;
	wire [3-1:0] node898;
	wire [3-1:0] node899;
	wire [3-1:0] node900;
	wire [3-1:0] node901;
	wire [3-1:0] node906;
	wire [3-1:0] node909;
	wire [3-1:0] node910;
	wire [3-1:0] node912;
	wire [3-1:0] node914;
	wire [3-1:0] node917;
	wire [3-1:0] node918;
	wire [3-1:0] node920;
	wire [3-1:0] node924;
	wire [3-1:0] node925;
	wire [3-1:0] node926;
	wire [3-1:0] node929;
	wire [3-1:0] node931;
	wire [3-1:0] node934;
	wire [3-1:0] node935;
	wire [3-1:0] node936;
	wire [3-1:0] node940;
	wire [3-1:0] node942;
	wire [3-1:0] node945;
	wire [3-1:0] node946;
	wire [3-1:0] node947;
	wire [3-1:0] node949;
	wire [3-1:0] node950;
	wire [3-1:0] node954;
	wire [3-1:0] node956;
	wire [3-1:0] node959;
	wire [3-1:0] node960;
	wire [3-1:0] node962;
	wire [3-1:0] node963;
	wire [3-1:0] node965;
	wire [3-1:0] node969;
	wire [3-1:0] node971;
	wire [3-1:0] node974;
	wire [3-1:0] node975;
	wire [3-1:0] node976;
	wire [3-1:0] node977;
	wire [3-1:0] node978;
	wire [3-1:0] node979;
	wire [3-1:0] node980;
	wire [3-1:0] node981;
	wire [3-1:0] node983;
	wire [3-1:0] node987;
	wire [3-1:0] node988;
	wire [3-1:0] node990;
	wire [3-1:0] node994;
	wire [3-1:0] node995;
	wire [3-1:0] node996;
	wire [3-1:0] node998;
	wire [3-1:0] node1000;
	wire [3-1:0] node1004;
	wire [3-1:0] node1005;
	wire [3-1:0] node1007;
	wire [3-1:0] node1009;
	wire [3-1:0] node1012;
	wire [3-1:0] node1013;
	wire [3-1:0] node1014;
	wire [3-1:0] node1019;
	wire [3-1:0] node1020;
	wire [3-1:0] node1021;
	wire [3-1:0] node1022;
	wire [3-1:0] node1023;
	wire [3-1:0] node1025;
	wire [3-1:0] node1029;
	wire [3-1:0] node1031;
	wire [3-1:0] node1033;
	wire [3-1:0] node1036;
	wire [3-1:0] node1037;
	wire [3-1:0] node1038;
	wire [3-1:0] node1040;
	wire [3-1:0] node1045;
	wire [3-1:0] node1046;
	wire [3-1:0] node1047;
	wire [3-1:0] node1051;
	wire [3-1:0] node1052;
	wire [3-1:0] node1056;
	wire [3-1:0] node1057;
	wire [3-1:0] node1058;
	wire [3-1:0] node1059;
	wire [3-1:0] node1063;
	wire [3-1:0] node1064;
	wire [3-1:0] node1066;
	wire [3-1:0] node1067;
	wire [3-1:0] node1068;
	wire [3-1:0] node1073;
	wire [3-1:0] node1076;
	wire [3-1:0] node1078;
	wire [3-1:0] node1079;
	wire [3-1:0] node1080;
	wire [3-1:0] node1082;
	wire [3-1:0] node1083;
	wire [3-1:0] node1089;
	wire [3-1:0] node1090;
	wire [3-1:0] node1091;
	wire [3-1:0] node1092;
	wire [3-1:0] node1093;
	wire [3-1:0] node1094;
	wire [3-1:0] node1096;
	wire [3-1:0] node1098;
	wire [3-1:0] node1101;
	wire [3-1:0] node1102;
	wire [3-1:0] node1103;
	wire [3-1:0] node1108;
	wire [3-1:0] node1110;
	wire [3-1:0] node1111;
	wire [3-1:0] node1115;
	wire [3-1:0] node1116;
	wire [3-1:0] node1118;
	wire [3-1:0] node1119;
	wire [3-1:0] node1120;
	wire [3-1:0] node1125;
	wire [3-1:0] node1127;
	wire [3-1:0] node1128;
	wire [3-1:0] node1132;
	wire [3-1:0] node1133;
	wire [3-1:0] node1134;
	wire [3-1:0] node1135;
	wire [3-1:0] node1137;
	wire [3-1:0] node1138;
	wire [3-1:0] node1143;
	wire [3-1:0] node1144;
	wire [3-1:0] node1146;
	wire [3-1:0] node1147;
	wire [3-1:0] node1152;
	wire [3-1:0] node1153;
	wire [3-1:0] node1154;
	wire [3-1:0] node1156;
	wire [3-1:0] node1160;
	wire [3-1:0] node1161;
	wire [3-1:0] node1163;
	wire [3-1:0] node1167;
	wire [3-1:0] node1168;
	wire [3-1:0] node1169;
	wire [3-1:0] node1170;
	wire [3-1:0] node1172;
	wire [3-1:0] node1173;
	wire [3-1:0] node1177;
	wire [3-1:0] node1179;
	wire [3-1:0] node1180;
	wire [3-1:0] node1184;
	wire [3-1:0] node1185;
	wire [3-1:0] node1187;
	wire [3-1:0] node1188;
	wire [3-1:0] node1190;
	wire [3-1:0] node1194;
	wire [3-1:0] node1196;
	wire [3-1:0] node1197;
	wire [3-1:0] node1199;
	wire [3-1:0] node1203;
	wire [3-1:0] node1204;
	wire [3-1:0] node1205;
	wire [3-1:0] node1206;
	wire [3-1:0] node1208;
	wire [3-1:0] node1212;
	wire [3-1:0] node1213;
	wire [3-1:0] node1215;
	wire [3-1:0] node1219;
	wire [3-1:0] node1220;
	wire [3-1:0] node1221;
	wire [3-1:0] node1223;
	wire [3-1:0] node1227;
	wire [3-1:0] node1228;
	wire [3-1:0] node1230;
	wire [3-1:0] node1232;
	wire [3-1:0] node1236;
	wire [3-1:0] node1237;
	wire [3-1:0] node1239;
	wire [3-1:0] node1240;
	wire [3-1:0] node1241;
	wire [3-1:0] node1242;
	wire [3-1:0] node1243;
	wire [3-1:0] node1244;
	wire [3-1:0] node1245;
	wire [3-1:0] node1250;
	wire [3-1:0] node1252;
	wire [3-1:0] node1255;
	wire [3-1:0] node1256;
	wire [3-1:0] node1257;
	wire [3-1:0] node1264;
	wire [3-1:0] node1265;
	wire [3-1:0] node1266;
	wire [3-1:0] node1267;
	wire [3-1:0] node1268;
	wire [3-1:0] node1269;
	wire [3-1:0] node1270;
	wire [3-1:0] node1274;
	wire [3-1:0] node1276;
	wire [3-1:0] node1279;
	wire [3-1:0] node1280;
	wire [3-1:0] node1281;
	wire [3-1:0] node1283;
	wire [3-1:0] node1287;
	wire [3-1:0] node1289;
	wire [3-1:0] node1291;
	wire [3-1:0] node1294;
	wire [3-1:0] node1295;
	wire [3-1:0] node1296;
	wire [3-1:0] node1297;
	wire [3-1:0] node1299;
	wire [3-1:0] node1303;
	wire [3-1:0] node1305;
	wire [3-1:0] node1308;
	wire [3-1:0] node1309;
	wire [3-1:0] node1310;
	wire [3-1:0] node1312;
	wire [3-1:0] node1316;
	wire [3-1:0] node1318;
	wire [3-1:0] node1321;
	wire [3-1:0] node1322;
	wire [3-1:0] node1323;
	wire [3-1:0] node1325;
	wire [3-1:0] node1326;
	wire [3-1:0] node1331;
	wire [3-1:0] node1332;
	wire [3-1:0] node1334;
	wire [3-1:0] node1337;
	wire [3-1:0] node1338;
	wire [3-1:0] node1339;
	wire [3-1:0] node1343;
	wire [3-1:0] node1346;
	wire [3-1:0] node1347;
	wire [3-1:0] node1348;
	wire [3-1:0] node1349;
	wire [3-1:0] node1350;
	wire [3-1:0] node1351;
	wire [3-1:0] node1353;
	wire [3-1:0] node1359;
	wire [3-1:0] node1360;
	wire [3-1:0] node1361;
	wire [3-1:0] node1365;
	wire [3-1:0] node1366;

	assign outp = (inp[6]) ? node416 : node1;
		assign node1 = (inp[9]) ? node373 : node2;
			assign node2 = (inp[0]) ? node282 : node3;
				assign node3 = (inp[7]) ? node113 : node4;
					assign node4 = (inp[10]) ? node80 : node5;
						assign node5 = (inp[1]) ? node51 : node6;
							assign node6 = (inp[8]) ? node26 : node7;
								assign node7 = (inp[11]) ? node17 : node8;
									assign node8 = (inp[3]) ? node14 : node9;
										assign node9 = (inp[2]) ? 3'b010 : node10;
											assign node10 = (inp[5]) ? 3'b010 : 3'b110;
										assign node14 = (inp[2]) ? 3'b100 : 3'b010;
									assign node17 = (inp[2]) ? node19 : 3'b100;
										assign node19 = (inp[3]) ? node21 : 3'b100;
											assign node21 = (inp[4]) ? 3'b000 : node22;
												assign node22 = (inp[5]) ? 3'b000 : 3'b100;
								assign node26 = (inp[11]) ? node40 : node27;
									assign node27 = (inp[2]) ? node35 : node28;
										assign node28 = (inp[3]) ? 3'b110 : node29;
											assign node29 = (inp[4]) ? 3'b110 : node30;
												assign node30 = (inp[5]) ? 3'b110 : 3'b001;
										assign node35 = (inp[3]) ? node37 : 3'b110;
											assign node37 = (inp[4]) ? 3'b010 : 3'b110;
									assign node40 = (inp[4]) ? node46 : node41;
										assign node41 = (inp[2]) ? 3'b010 : node42;
											assign node42 = (inp[3]) ? 3'b010 : 3'b110;
										assign node46 = (inp[2]) ? node48 : 3'b010;
											assign node48 = (inp[3]) ? 3'b100 : 3'b010;
							assign node51 = (inp[11]) ? node69 : node52;
								assign node52 = (inp[8]) ? node60 : node53;
									assign node53 = (inp[2]) ? node55 : 3'b100;
										assign node55 = (inp[3]) ? 3'b000 : node56;
											assign node56 = (inp[4]) ? 3'b000 : 3'b100;
									assign node60 = (inp[2]) ? node62 : 3'b010;
										assign node62 = (inp[3]) ? 3'b100 : node63;
											assign node63 = (inp[4]) ? node65 : 3'b010;
												assign node65 = (inp[5]) ? 3'b100 : 3'b010;
								assign node69 = (inp[8]) ? node71 : 3'b000;
									assign node71 = (inp[2]) ? node73 : 3'b100;
										assign node73 = (inp[3]) ? 3'b000 : node74;
											assign node74 = (inp[4]) ? node76 : 3'b100;
												assign node76 = (inp[5]) ? 3'b000 : 3'b100;
						assign node80 = (inp[1]) ? 3'b000 : node81;
							assign node81 = (inp[8]) ? node91 : node82;
								assign node82 = (inp[5]) ? 3'b000 : node83;
									assign node83 = (inp[4]) ? 3'b000 : node84;
										assign node84 = (inp[11]) ? 3'b000 : node85;
											assign node85 = (inp[3]) ? 3'b000 : 3'b100;
								assign node91 = (inp[11]) ? node103 : node92;
									assign node92 = (inp[2]) ? node98 : node93;
										assign node93 = (inp[4]) ? 3'b100 : node94;
											assign node94 = (inp[3]) ? 3'b100 : 3'b010;
										assign node98 = (inp[3]) ? node100 : 3'b100;
											assign node100 = (inp[4]) ? 3'b000 : 3'b100;
									assign node103 = (inp[2]) ? 3'b000 : node104;
										assign node104 = (inp[3]) ? 3'b000 : node105;
											assign node105 = (inp[5]) ? node107 : 3'b100;
												assign node107 = (inp[4]) ? 3'b000 : 3'b100;
					assign node113 = (inp[10]) ? node205 : node114;
						assign node114 = (inp[1]) ? node162 : node115;
							assign node115 = (inp[8]) ? node137 : node116;
								assign node116 = (inp[11]) ? node128 : node117;
									assign node117 = (inp[3]) ? node123 : node118;
										assign node118 = (inp[2]) ? 3'b001 : node119;
											assign node119 = (inp[4]) ? 3'b001 : 3'b101;
										assign node123 = (inp[2]) ? node125 : 3'b001;
											assign node125 = (inp[4]) ? 3'b110 : 3'b001;
									assign node128 = (inp[2]) ? node132 : node129;
										assign node129 = (inp[3]) ? 3'b110 : 3'b001;
										assign node132 = (inp[3]) ? node134 : 3'b110;
											assign node134 = (inp[4]) ? 3'b010 : 3'b110;
								assign node137 = (inp[11]) ? node151 : node138;
									assign node138 = (inp[3]) ? node144 : node139;
										assign node139 = (inp[2]) ? 3'b101 : node140;
											assign node140 = (inp[5]) ? 3'b101 : 3'b011;
										assign node144 = (inp[4]) ? node146 : 3'b101;
											assign node146 = (inp[5]) ? node148 : 3'b101;
												assign node148 = (inp[2]) ? 3'b001 : 3'b101;
									assign node151 = (inp[3]) ? node155 : node152;
										assign node152 = (inp[2]) ? 3'b001 : 3'b101;
										assign node155 = (inp[5]) ? node157 : 3'b001;
											assign node157 = (inp[4]) ? node159 : 3'b001;
												assign node159 = (inp[2]) ? 3'b110 : 3'b001;
							assign node162 = (inp[8]) ? node178 : node163;
								assign node163 = (inp[11]) ? node173 : node164;
									assign node164 = (inp[2]) ? node166 : 3'b110;
										assign node166 = (inp[3]) ? 3'b010 : node167;
											assign node167 = (inp[5]) ? node169 : 3'b110;
												assign node169 = (inp[4]) ? 3'b010 : 3'b110;
									assign node173 = (inp[2]) ? node175 : 3'b010;
										assign node175 = (inp[3]) ? 3'b100 : 3'b010;
								assign node178 = (inp[11]) ? node190 : node179;
									assign node179 = (inp[2]) ? node187 : node180;
										assign node180 = (inp[4]) ? 3'b001 : node181;
											assign node181 = (inp[5]) ? 3'b001 : node182;
												assign node182 = (inp[3]) ? 3'b001 : 3'b101;
										assign node187 = (inp[3]) ? 3'b110 : 3'b001;
									assign node190 = (inp[2]) ? node198 : node191;
										assign node191 = (inp[5]) ? 3'b110 : node192;
											assign node192 = (inp[4]) ? 3'b110 : node193;
												assign node193 = (inp[3]) ? 3'b110 : 3'b001;
										assign node198 = (inp[3]) ? node200 : 3'b110;
											assign node200 = (inp[4]) ? 3'b010 : node201;
												assign node201 = (inp[5]) ? 3'b010 : 3'b110;
						assign node205 = (inp[1]) ? node245 : node206;
							assign node206 = (inp[8]) ? node234 : node207;
								assign node207 = (inp[11]) ? node223 : node208;
									assign node208 = (inp[2]) ? node216 : node209;
										assign node209 = (inp[3]) ? 3'b010 : node210;
											assign node210 = (inp[4]) ? node212 : 3'b110;
												assign node212 = (inp[5]) ? 3'b010 : 3'b110;
										assign node216 = (inp[4]) ? node218 : 3'b010;
											assign node218 = (inp[5]) ? node220 : 3'b010;
												assign node220 = (inp[3]) ? 3'b100 : 3'b010;
									assign node223 = (inp[3]) ? node227 : node224;
										assign node224 = (inp[2]) ? 3'b100 : 3'b010;
										assign node227 = (inp[2]) ? node229 : 3'b100;
											assign node229 = (inp[5]) ? node231 : 3'b100;
												assign node231 = (inp[4]) ? 3'b000 : 3'b100;
								assign node234 = (inp[11]) ? node240 : node235;
									assign node235 = (inp[2]) ? 3'b110 : node236;
										assign node236 = (inp[3]) ? 3'b110 : 3'b001;
									assign node240 = (inp[2]) ? 3'b010 : node241;
										assign node241 = (inp[3]) ? 3'b010 : 3'b110;
							assign node245 = (inp[8]) ? node253 : node246;
								assign node246 = (inp[11]) ? 3'b000 : node247;
									assign node247 = (inp[3]) ? node249 : 3'b100;
										assign node249 = (inp[2]) ? 3'b000 : 3'b100;
								assign node253 = (inp[11]) ? node269 : node254;
									assign node254 = (inp[3]) ? node262 : node255;
										assign node255 = (inp[2]) ? 3'b010 : node256;
											assign node256 = (inp[5]) ? 3'b010 : node257;
												assign node257 = (inp[4]) ? 3'b010 : 3'b110;
										assign node262 = (inp[2]) ? node264 : 3'b010;
											assign node264 = (inp[5]) ? 3'b100 : node265;
												assign node265 = (inp[4]) ? 3'b100 : 3'b010;
									assign node269 = (inp[3]) ? node275 : node270;
										assign node270 = (inp[2]) ? 3'b100 : node271;
											assign node271 = (inp[4]) ? 3'b100 : 3'b010;
										assign node275 = (inp[2]) ? node277 : 3'b100;
											assign node277 = (inp[4]) ? 3'b000 : node278;
												assign node278 = (inp[5]) ? 3'b000 : 3'b100;
				assign node282 = (inp[7]) ? node298 : node283;
					assign node283 = (inp[11]) ? 3'b000 : node284;
						assign node284 = (inp[1]) ? 3'b000 : node285;
							assign node285 = (inp[10]) ? 3'b000 : node286;
								assign node286 = (inp[8]) ? node288 : 3'b000;
									assign node288 = (inp[2]) ? 3'b000 : node289;
										assign node289 = (inp[4]) ? node291 : 3'b100;
											assign node291 = (inp[3]) ? 3'b000 : 3'b100;
					assign node298 = (inp[10]) ? node360 : node299;
						assign node299 = (inp[1]) ? node337 : node300;
							assign node300 = (inp[8]) ? node322 : node301;
								assign node301 = (inp[11]) ? node315 : node302;
									assign node302 = (inp[2]) ? node308 : node303;
										assign node303 = (inp[4]) ? node305 : 3'b010;
											assign node305 = (inp[5]) ? 3'b100 : 3'b010;
										assign node308 = (inp[3]) ? 3'b100 : node309;
											assign node309 = (inp[5]) ? 3'b100 : node310;
												assign node310 = (inp[4]) ? 3'b100 : 3'b010;
									assign node315 = (inp[2]) ? node317 : 3'b100;
										assign node317 = (inp[3]) ? 3'b000 : node318;
											assign node318 = (inp[4]) ? 3'b000 : 3'b100;
								assign node322 = (inp[11]) ? node330 : node323;
									assign node323 = (inp[2]) ? node325 : 3'b110;
										assign node325 = (inp[4]) ? 3'b010 : node326;
											assign node326 = (inp[3]) ? 3'b010 : 3'b110;
									assign node330 = (inp[2]) ? node332 : 3'b010;
										assign node332 = (inp[3]) ? 3'b100 : node333;
											assign node333 = (inp[4]) ? 3'b100 : 3'b010;
							assign node337 = (inp[8]) ? node345 : node338;
								assign node338 = (inp[11]) ? 3'b000 : node339;
									assign node339 = (inp[3]) ? 3'b000 : node340;
										assign node340 = (inp[2]) ? 3'b000 : 3'b100;
								assign node345 = (inp[11]) ? node353 : node346;
									assign node346 = (inp[2]) ? 3'b100 : node347;
										assign node347 = (inp[3]) ? node349 : 3'b010;
											assign node349 = (inp[4]) ? 3'b100 : 3'b010;
									assign node353 = (inp[2]) ? 3'b000 : node354;
										assign node354 = (inp[3]) ? node356 : 3'b100;
											assign node356 = (inp[4]) ? 3'b000 : 3'b100;
						assign node360 = (inp[8]) ? node362 : 3'b000;
							assign node362 = (inp[11]) ? 3'b000 : node363;
								assign node363 = (inp[1]) ? 3'b000 : node364;
									assign node364 = (inp[2]) ? node366 : 3'b100;
										assign node366 = (inp[4]) ? 3'b000 : node367;
											assign node367 = (inp[3]) ? 3'b000 : 3'b100;
			assign node373 = (inp[10]) ? 3'b000 : node374;
				assign node374 = (inp[7]) ? node376 : 3'b000;
					assign node376 = (inp[0]) ? 3'b000 : node377;
						assign node377 = (inp[1]) ? node403 : node378;
							assign node378 = (inp[8]) ? node386 : node379;
								assign node379 = (inp[11]) ? 3'b000 : node380;
									assign node380 = (inp[3]) ? 3'b000 : node381;
										assign node381 = (inp[2]) ? 3'b000 : 3'b100;
								assign node386 = (inp[11]) ? node396 : node387;
									assign node387 = (inp[2]) ? 3'b100 : node388;
										assign node388 = (inp[3]) ? node390 : 3'b010;
											assign node390 = (inp[5]) ? 3'b100 : node391;
												assign node391 = (inp[4]) ? 3'b100 : 3'b010;
									assign node396 = (inp[2]) ? 3'b000 : node397;
										assign node397 = (inp[3]) ? node399 : 3'b100;
											assign node399 = (inp[4]) ? 3'b000 : 3'b100;
							assign node403 = (inp[4]) ? 3'b000 : node404;
								assign node404 = (inp[11]) ? 3'b000 : node405;
									assign node405 = (inp[8]) ? node407 : 3'b000;
										assign node407 = (inp[3]) ? 3'b000 : node408;
											assign node408 = (inp[2]) ? 3'b000 : 3'b100;
		assign node416 = (inp[9]) ? node974 : node417;
			assign node417 = (inp[0]) ? node663 : node418;
				assign node418 = (inp[7]) ? node582 : node419;
					assign node419 = (inp[10]) ? node495 : node420;
						assign node420 = (inp[1]) ? node444 : node421;
							assign node421 = (inp[8]) ? node435 : node422;
								assign node422 = (inp[11]) ? node428 : node423;
									assign node423 = (inp[2]) ? 3'b011 : node424;
										assign node424 = (inp[3]) ? 3'b011 : 3'b111;
									assign node428 = (inp[2]) ? 3'b101 : node429;
										assign node429 = (inp[3]) ? node431 : 3'b011;
											assign node431 = (inp[5]) ? 3'b101 : 3'b011;
								assign node435 = (inp[11]) ? node437 : 3'b111;
									assign node437 = (inp[2]) ? 3'b011 : node438;
										assign node438 = (inp[3]) ? node440 : 3'b111;
											assign node440 = (inp[5]) ? 3'b011 : 3'b111;
							assign node444 = (inp[8]) ? node472 : node445;
								assign node445 = (inp[11]) ? node461 : node446;
									assign node446 = (inp[2]) ? node454 : node447;
										assign node447 = (inp[5]) ? 3'b101 : node448;
											assign node448 = (inp[3]) ? 3'b101 : node449;
												assign node449 = (inp[4]) ? 3'b101 : 3'b011;
										assign node454 = (inp[3]) ? node456 : 3'b101;
											assign node456 = (inp[4]) ? 3'b001 : node457;
												assign node457 = (inp[5]) ? 3'b001 : 3'b101;
									assign node461 = (inp[4]) ? node467 : node462;
										assign node462 = (inp[2]) ? 3'b001 : node463;
											assign node463 = (inp[3]) ? 3'b001 : 3'b101;
										assign node467 = (inp[2]) ? node469 : 3'b001;
											assign node469 = (inp[3]) ? 3'b110 : 3'b001;
								assign node472 = (inp[11]) ? node484 : node473;
									assign node473 = (inp[3]) ? node479 : node474;
										assign node474 = (inp[2]) ? 3'b011 : node475;
											assign node475 = (inp[4]) ? 3'b011 : 3'b111;
										assign node479 = (inp[2]) ? node481 : 3'b011;
											assign node481 = (inp[4]) ? 3'b101 : 3'b011;
									assign node484 = (inp[2]) ? node490 : node485;
										assign node485 = (inp[3]) ? 3'b101 : node486;
											assign node486 = (inp[4]) ? 3'b101 : 3'b011;
										assign node490 = (inp[3]) ? node492 : 3'b101;
											assign node492 = (inp[4]) ? 3'b001 : 3'b101;
						assign node495 = (inp[1]) ? node531 : node496;
							assign node496 = (inp[11]) ? node514 : node497;
								assign node497 = (inp[8]) ? node507 : node498;
									assign node498 = (inp[2]) ? 3'b001 : node499;
										assign node499 = (inp[3]) ? node501 : 3'b101;
											assign node501 = (inp[4]) ? 3'b001 : node502;
												assign node502 = (inp[5]) ? 3'b001 : 3'b101;
									assign node507 = (inp[2]) ? 3'b101 : node508;
										assign node508 = (inp[4]) ? node510 : 3'b011;
											assign node510 = (inp[3]) ? 3'b101 : 3'b011;
								assign node514 = (inp[8]) ? node524 : node515;
									assign node515 = (inp[2]) ? 3'b110 : node516;
										assign node516 = (inp[3]) ? node518 : 3'b001;
											assign node518 = (inp[4]) ? 3'b110 : node519;
												assign node519 = (inp[5]) ? 3'b110 : 3'b001;
									assign node524 = (inp[2]) ? 3'b001 : node525;
										assign node525 = (inp[4]) ? node527 : 3'b101;
											assign node527 = (inp[3]) ? 3'b001 : 3'b101;
							assign node531 = (inp[8]) ? node557 : node532;
								assign node532 = (inp[11]) ? node544 : node533;
									assign node533 = (inp[3]) ? node539 : node534;
										assign node534 = (inp[4]) ? 3'b110 : node535;
											assign node535 = (inp[2]) ? 3'b110 : 3'b001;
										assign node539 = (inp[4]) ? node541 : 3'b110;
											assign node541 = (inp[2]) ? 3'b010 : 3'b110;
									assign node544 = (inp[3]) ? node552 : node545;
										assign node545 = (inp[2]) ? 3'b010 : node546;
											assign node546 = (inp[4]) ? node548 : 3'b110;
												assign node548 = (inp[5]) ? 3'b010 : 3'b110;
										assign node552 = (inp[2]) ? node554 : 3'b010;
											assign node554 = (inp[4]) ? 3'b100 : 3'b010;
								assign node557 = (inp[11]) ? node571 : node558;
									assign node558 = (inp[2]) ? node566 : node559;
										assign node559 = (inp[3]) ? 3'b001 : node560;
											assign node560 = (inp[5]) ? node562 : 3'b101;
												assign node562 = (inp[4]) ? 3'b001 : 3'b101;
										assign node566 = (inp[4]) ? node568 : 3'b001;
											assign node568 = (inp[3]) ? 3'b110 : 3'b001;
									assign node571 = (inp[2]) ? node575 : node572;
										assign node572 = (inp[3]) ? 3'b110 : 3'b001;
										assign node575 = (inp[3]) ? node577 : 3'b110;
											assign node577 = (inp[4]) ? node579 : 3'b110;
												assign node579 = (inp[5]) ? 3'b010 : 3'b110;
					assign node582 = (inp[10]) ? node602 : node583;
						assign node583 = (inp[8]) ? 3'b111 : node584;
							assign node584 = (inp[1]) ? node586 : 3'b111;
								assign node586 = (inp[11]) ? node596 : node587;
									assign node587 = (inp[4]) ? node589 : 3'b111;
										assign node589 = (inp[3]) ? node591 : 3'b111;
											assign node591 = (inp[2]) ? node593 : 3'b111;
												assign node593 = (inp[5]) ? 3'b011 : 3'b111;
									assign node596 = (inp[2]) ? 3'b011 : node597;
										assign node597 = (inp[3]) ? 3'b011 : 3'b111;
						assign node602 = (inp[1]) ? node636 : node603;
							assign node603 = (inp[8]) ? node627 : node604;
								assign node604 = (inp[11]) ? node614 : node605;
									assign node605 = (inp[2]) ? 3'b011 : node606;
										assign node606 = (inp[4]) ? node608 : 3'b111;
											assign node608 = (inp[5]) ? node610 : 3'b111;
												assign node610 = (inp[3]) ? 3'b011 : 3'b111;
									assign node614 = (inp[2]) ? node620 : node615;
										assign node615 = (inp[4]) ? node617 : 3'b011;
											assign node617 = (inp[3]) ? 3'b101 : 3'b011;
										assign node620 = (inp[5]) ? 3'b101 : node621;
											assign node621 = (inp[3]) ? 3'b101 : node622;
												assign node622 = (inp[4]) ? 3'b101 : 3'b011;
								assign node627 = (inp[2]) ? node629 : 3'b111;
									assign node629 = (inp[11]) ? node631 : 3'b111;
										assign node631 = (inp[4]) ? 3'b011 : node632;
											assign node632 = (inp[3]) ? 3'b011 : 3'b111;
							assign node636 = (inp[8]) ? node648 : node637;
								assign node637 = (inp[11]) ? node643 : node638;
									assign node638 = (inp[3]) ? 3'b101 : node639;
										assign node639 = (inp[2]) ? 3'b101 : 3'b011;
									assign node643 = (inp[2]) ? 3'b001 : node644;
										assign node644 = (inp[3]) ? 3'b001 : 3'b101;
								assign node648 = (inp[11]) ? node654 : node649;
									assign node649 = (inp[2]) ? 3'b011 : node650;
										assign node650 = (inp[3]) ? 3'b011 : 3'b111;
									assign node654 = (inp[2]) ? 3'b101 : node655;
										assign node655 = (inp[3]) ? node657 : 3'b011;
											assign node657 = (inp[5]) ? 3'b101 : node658;
												assign node658 = (inp[4]) ? 3'b101 : 3'b011;
				assign node663 = (inp[7]) ? node813 : node664;
					assign node664 = (inp[10]) ? node740 : node665;
						assign node665 = (inp[1]) ? node697 : node666;
							assign node666 = (inp[8]) ? node682 : node667;
								assign node667 = (inp[11]) ? node675 : node668;
									assign node668 = (inp[2]) ? node670 : 3'b001;
										assign node670 = (inp[3]) ? 3'b110 : node671;
											assign node671 = (inp[4]) ? 3'b110 : 3'b001;
									assign node675 = (inp[2]) ? node677 : 3'b110;
										assign node677 = (inp[3]) ? 3'b010 : node678;
											assign node678 = (inp[5]) ? 3'b010 : 3'b110;
								assign node682 = (inp[11]) ? node692 : node683;
									assign node683 = (inp[2]) ? node685 : 3'b101;
										assign node685 = (inp[3]) ? 3'b001 : node686;
											assign node686 = (inp[5]) ? node688 : 3'b101;
												assign node688 = (inp[4]) ? 3'b001 : 3'b101;
									assign node692 = (inp[2]) ? node694 : 3'b001;
										assign node694 = (inp[3]) ? 3'b110 : 3'b001;
							assign node697 = (inp[11]) ? node717 : node698;
								assign node698 = (inp[8]) ? node706 : node699;
									assign node699 = (inp[2]) ? 3'b010 : node700;
										assign node700 = (inp[4]) ? node702 : 3'b110;
											assign node702 = (inp[3]) ? 3'b010 : 3'b110;
									assign node706 = (inp[2]) ? node712 : node707;
										assign node707 = (inp[4]) ? node709 : 3'b001;
											assign node709 = (inp[5]) ? 3'b110 : 3'b001;
										assign node712 = (inp[3]) ? 3'b110 : node713;
											assign node713 = (inp[4]) ? 3'b110 : 3'b001;
								assign node717 = (inp[8]) ? node725 : node718;
									assign node718 = (inp[2]) ? 3'b100 : node719;
										assign node719 = (inp[5]) ? node721 : 3'b010;
											assign node721 = (inp[4]) ? 3'b100 : 3'b010;
									assign node725 = (inp[2]) ? node733 : node726;
										assign node726 = (inp[4]) ? node728 : 3'b110;
											assign node728 = (inp[3]) ? node730 : 3'b110;
												assign node730 = (inp[5]) ? 3'b010 : 3'b110;
										assign node733 = (inp[5]) ? 3'b010 : node734;
											assign node734 = (inp[3]) ? 3'b010 : node735;
												assign node735 = (inp[4]) ? 3'b010 : 3'b110;
						assign node740 = (inp[1]) ? node778 : node741;
							assign node741 = (inp[8]) ? node757 : node742;
								assign node742 = (inp[11]) ? node752 : node743;
									assign node743 = (inp[2]) ? node745 : 3'b010;
										assign node745 = (inp[3]) ? 3'b100 : node746;
											assign node746 = (inp[5]) ? node748 : 3'b010;
												assign node748 = (inp[4]) ? 3'b100 : 3'b010;
									assign node752 = (inp[2]) ? node754 : 3'b100;
										assign node754 = (inp[3]) ? 3'b000 : 3'b100;
								assign node757 = (inp[11]) ? node763 : node758;
									assign node758 = (inp[3]) ? node760 : 3'b110;
										assign node760 = (inp[2]) ? 3'b010 : 3'b110;
									assign node763 = (inp[2]) ? node771 : node764;
										assign node764 = (inp[5]) ? 3'b010 : node765;
											assign node765 = (inp[3]) ? 3'b010 : node766;
												assign node766 = (inp[4]) ? 3'b010 : 3'b110;
										assign node771 = (inp[3]) ? node773 : 3'b010;
											assign node773 = (inp[4]) ? 3'b100 : node774;
												assign node774 = (inp[5]) ? 3'b100 : 3'b010;
							assign node778 = (inp[8]) ? node796 : node779;
								assign node779 = (inp[11]) ? 3'b000 : node780;
									assign node780 = (inp[2]) ? node788 : node781;
										assign node781 = (inp[4]) ? node783 : 3'b100;
											assign node783 = (inp[3]) ? node785 : 3'b100;
												assign node785 = (inp[5]) ? 3'b000 : 3'b100;
										assign node788 = (inp[3]) ? 3'b000 : node789;
											assign node789 = (inp[5]) ? 3'b000 : node790;
												assign node790 = (inp[4]) ? 3'b000 : 3'b100;
								assign node796 = (inp[11]) ? node806 : node797;
									assign node797 = (inp[2]) ? node799 : 3'b010;
										assign node799 = (inp[4]) ? 3'b100 : node800;
											assign node800 = (inp[5]) ? 3'b100 : node801;
												assign node801 = (inp[3]) ? 3'b100 : 3'b010;
									assign node806 = (inp[2]) ? node808 : 3'b100;
										assign node808 = (inp[4]) ? 3'b000 : node809;
											assign node809 = (inp[3]) ? 3'b000 : 3'b100;
					assign node813 = (inp[10]) ? node895 : node814;
						assign node814 = (inp[1]) ? node864 : node815;
							assign node815 = (inp[8]) ? node843 : node816;
								assign node816 = (inp[11]) ? node828 : node817;
									assign node817 = (inp[3]) ? node825 : node818;
										assign node818 = (inp[5]) ? 3'b011 : node819;
											assign node819 = (inp[2]) ? 3'b011 : node820;
												assign node820 = (inp[4]) ? 3'b011 : 3'b111;
										assign node825 = (inp[2]) ? 3'b101 : 3'b011;
									assign node828 = (inp[2]) ? node836 : node829;
										assign node829 = (inp[5]) ? 3'b101 : node830;
											assign node830 = (inp[4]) ? 3'b101 : node831;
												assign node831 = (inp[3]) ? 3'b101 : 3'b011;
										assign node836 = (inp[3]) ? node838 : 3'b101;
											assign node838 = (inp[5]) ? 3'b001 : node839;
												assign node839 = (inp[4]) ? 3'b001 : 3'b101;
								assign node843 = (inp[11]) ? node853 : node844;
									assign node844 = (inp[3]) ? node846 : 3'b111;
										assign node846 = (inp[2]) ? node848 : 3'b111;
											assign node848 = (inp[5]) ? 3'b011 : node849;
												assign node849 = (inp[4]) ? 3'b011 : 3'b111;
									assign node853 = (inp[4]) ? node859 : node854;
										assign node854 = (inp[3]) ? 3'b011 : node855;
											assign node855 = (inp[2]) ? 3'b011 : 3'b111;
										assign node859 = (inp[2]) ? node861 : 3'b011;
											assign node861 = (inp[3]) ? 3'b101 : 3'b011;
							assign node864 = (inp[11]) ? node880 : node865;
								assign node865 = (inp[8]) ? node873 : node866;
									assign node866 = (inp[2]) ? node868 : 3'b101;
										assign node868 = (inp[4]) ? 3'b001 : node869;
											assign node869 = (inp[3]) ? 3'b001 : 3'b101;
									assign node873 = (inp[2]) ? node875 : 3'b011;
										assign node875 = (inp[3]) ? 3'b101 : node876;
											assign node876 = (inp[4]) ? 3'b101 : 3'b011;
								assign node880 = (inp[8]) ? node888 : node881;
									assign node881 = (inp[2]) ? node883 : 3'b001;
										assign node883 = (inp[4]) ? 3'b110 : node884;
											assign node884 = (inp[3]) ? 3'b110 : 3'b001;
									assign node888 = (inp[2]) ? node890 : 3'b101;
										assign node890 = (inp[3]) ? 3'b001 : node891;
											assign node891 = (inp[5]) ? 3'b001 : 3'b101;
						assign node895 = (inp[1]) ? node945 : node896;
							assign node896 = (inp[8]) ? node924 : node897;
								assign node897 = (inp[11]) ? node909 : node898;
									assign node898 = (inp[3]) ? node906 : node899;
										assign node899 = (inp[2]) ? 3'b001 : node900;
											assign node900 = (inp[4]) ? 3'b001 : node901;
												assign node901 = (inp[5]) ? 3'b001 : 3'b101;
										assign node906 = (inp[2]) ? 3'b110 : 3'b001;
									assign node909 = (inp[5]) ? node917 : node910;
										assign node910 = (inp[4]) ? node912 : 3'b110;
											assign node912 = (inp[3]) ? node914 : 3'b110;
												assign node914 = (inp[2]) ? 3'b010 : 3'b110;
										assign node917 = (inp[4]) ? 3'b110 : node918;
											assign node918 = (inp[2]) ? node920 : 3'b001;
												assign node920 = (inp[3]) ? 3'b010 : 3'b110;
								assign node924 = (inp[11]) ? node934 : node925;
									assign node925 = (inp[3]) ? node929 : node926;
										assign node926 = (inp[4]) ? 3'b101 : 3'b011;
										assign node929 = (inp[4]) ? node931 : 3'b101;
											assign node931 = (inp[2]) ? 3'b001 : 3'b101;
									assign node934 = (inp[2]) ? node940 : node935;
										assign node935 = (inp[3]) ? 3'b001 : node936;
											assign node936 = (inp[4]) ? 3'b001 : 3'b101;
										assign node940 = (inp[4]) ? node942 : 3'b001;
											assign node942 = (inp[3]) ? 3'b110 : 3'b001;
							assign node945 = (inp[11]) ? node959 : node946;
								assign node946 = (inp[8]) ? node954 : node947;
									assign node947 = (inp[2]) ? node949 : 3'b110;
										assign node949 = (inp[3]) ? 3'b010 : node950;
											assign node950 = (inp[4]) ? 3'b010 : 3'b110;
									assign node954 = (inp[2]) ? node956 : 3'b001;
										assign node956 = (inp[3]) ? 3'b110 : 3'b001;
								assign node959 = (inp[8]) ? node969 : node960;
									assign node960 = (inp[2]) ? node962 : 3'b010;
										assign node962 = (inp[3]) ? 3'b100 : node963;
											assign node963 = (inp[5]) ? node965 : 3'b010;
												assign node965 = (inp[4]) ? 3'b100 : 3'b010;
									assign node969 = (inp[3]) ? node971 : 3'b110;
										assign node971 = (inp[2]) ? 3'b010 : 3'b110;
			assign node974 = (inp[0]) ? node1236 : node975;
				assign node975 = (inp[7]) ? node1089 : node976;
					assign node976 = (inp[10]) ? node1056 : node977;
						assign node977 = (inp[1]) ? node1019 : node978;
							assign node978 = (inp[8]) ? node994 : node979;
								assign node979 = (inp[11]) ? node987 : node980;
									assign node980 = (inp[2]) ? 3'b010 : node981;
										assign node981 = (inp[3]) ? node983 : 3'b110;
											assign node983 = (inp[4]) ? 3'b010 : 3'b110;
									assign node987 = (inp[2]) ? 3'b100 : node988;
										assign node988 = (inp[3]) ? node990 : 3'b010;
											assign node990 = (inp[4]) ? 3'b100 : 3'b010;
								assign node994 = (inp[11]) ? node1004 : node995;
									assign node995 = (inp[2]) ? 3'b110 : node996;
										assign node996 = (inp[5]) ? node998 : 3'b001;
											assign node998 = (inp[4]) ? node1000 : 3'b001;
												assign node1000 = (inp[3]) ? 3'b110 : 3'b001;
									assign node1004 = (inp[2]) ? node1012 : node1005;
										assign node1005 = (inp[3]) ? node1007 : 3'b110;
											assign node1007 = (inp[5]) ? node1009 : 3'b110;
												assign node1009 = (inp[4]) ? 3'b010 : 3'b110;
										assign node1012 = (inp[4]) ? 3'b010 : node1013;
											assign node1013 = (inp[5]) ? 3'b010 : node1014;
												assign node1014 = (inp[3]) ? 3'b010 : 3'b110;
							assign node1019 = (inp[8]) ? node1045 : node1020;
								assign node1020 = (inp[11]) ? node1036 : node1021;
									assign node1021 = (inp[2]) ? node1029 : node1022;
										assign node1022 = (inp[3]) ? 3'b100 : node1023;
											assign node1023 = (inp[4]) ? node1025 : 3'b010;
												assign node1025 = (inp[5]) ? 3'b100 : 3'b010;
										assign node1029 = (inp[3]) ? node1031 : 3'b100;
											assign node1031 = (inp[4]) ? node1033 : 3'b100;
												assign node1033 = (inp[5]) ? 3'b000 : 3'b100;
									assign node1036 = (inp[3]) ? 3'b000 : node1037;
										assign node1037 = (inp[2]) ? 3'b000 : node1038;
											assign node1038 = (inp[4]) ? node1040 : 3'b100;
												assign node1040 = (inp[5]) ? 3'b000 : 3'b100;
								assign node1045 = (inp[11]) ? node1051 : node1046;
									assign node1046 = (inp[2]) ? 3'b010 : node1047;
										assign node1047 = (inp[3]) ? 3'b010 : 3'b110;
									assign node1051 = (inp[2]) ? 3'b100 : node1052;
										assign node1052 = (inp[3]) ? 3'b100 : 3'b010;
						assign node1056 = (inp[1]) ? node1076 : node1057;
							assign node1057 = (inp[8]) ? node1063 : node1058;
								assign node1058 = (inp[11]) ? 3'b000 : node1059;
									assign node1059 = (inp[2]) ? 3'b000 : 3'b100;
								assign node1063 = (inp[11]) ? node1073 : node1064;
									assign node1064 = (inp[2]) ? node1066 : 3'b010;
										assign node1066 = (inp[3]) ? 3'b100 : node1067;
											assign node1067 = (inp[4]) ? 3'b100 : node1068;
												assign node1068 = (inp[5]) ? 3'b100 : 3'b010;
									assign node1073 = (inp[2]) ? 3'b000 : 3'b100;
							assign node1076 = (inp[8]) ? node1078 : 3'b000;
								assign node1078 = (inp[11]) ? 3'b000 : node1079;
									assign node1079 = (inp[2]) ? 3'b000 : node1080;
										assign node1080 = (inp[3]) ? node1082 : 3'b100;
											assign node1082 = (inp[4]) ? 3'b000 : node1083;
												assign node1083 = (inp[5]) ? 3'b000 : 3'b100;
					assign node1089 = (inp[10]) ? node1167 : node1090;
						assign node1090 = (inp[1]) ? node1132 : node1091;
							assign node1091 = (inp[11]) ? node1115 : node1092;
								assign node1092 = (inp[8]) ? node1108 : node1093;
									assign node1093 = (inp[2]) ? node1101 : node1094;
										assign node1094 = (inp[5]) ? node1096 : 3'b101;
											assign node1096 = (inp[3]) ? node1098 : 3'b101;
												assign node1098 = (inp[4]) ? 3'b001 : 3'b101;
										assign node1101 = (inp[5]) ? 3'b001 : node1102;
											assign node1102 = (inp[3]) ? 3'b001 : node1103;
												assign node1103 = (inp[4]) ? 3'b001 : 3'b101;
									assign node1108 = (inp[2]) ? node1110 : 3'b011;
										assign node1110 = (inp[4]) ? 3'b101 : node1111;
											assign node1111 = (inp[3]) ? 3'b101 : 3'b011;
								assign node1115 = (inp[8]) ? node1125 : node1116;
									assign node1116 = (inp[2]) ? node1118 : 3'b001;
										assign node1118 = (inp[3]) ? 3'b110 : node1119;
											assign node1119 = (inp[5]) ? 3'b110 : node1120;
												assign node1120 = (inp[4]) ? 3'b110 : 3'b001;
									assign node1125 = (inp[2]) ? node1127 : 3'b101;
										assign node1127 = (inp[4]) ? 3'b001 : node1128;
											assign node1128 = (inp[3]) ? 3'b001 : 3'b101;
							assign node1132 = (inp[8]) ? node1152 : node1133;
								assign node1133 = (inp[11]) ? node1143 : node1134;
									assign node1134 = (inp[2]) ? 3'b110 : node1135;
										assign node1135 = (inp[3]) ? node1137 : 3'b001;
											assign node1137 = (inp[4]) ? 3'b110 : node1138;
												assign node1138 = (inp[5]) ? 3'b110 : 3'b001;
									assign node1143 = (inp[2]) ? 3'b010 : node1144;
										assign node1144 = (inp[3]) ? node1146 : 3'b110;
											assign node1146 = (inp[5]) ? 3'b010 : node1147;
												assign node1147 = (inp[4]) ? 3'b010 : 3'b110;
								assign node1152 = (inp[11]) ? node1160 : node1153;
									assign node1153 = (inp[2]) ? 3'b001 : node1154;
										assign node1154 = (inp[4]) ? node1156 : 3'b101;
											assign node1156 = (inp[3]) ? 3'b001 : 3'b101;
									assign node1160 = (inp[2]) ? 3'b110 : node1161;
										assign node1161 = (inp[4]) ? node1163 : 3'b001;
											assign node1163 = (inp[3]) ? 3'b110 : 3'b001;
						assign node1167 = (inp[1]) ? node1203 : node1168;
							assign node1168 = (inp[8]) ? node1184 : node1169;
								assign node1169 = (inp[11]) ? node1177 : node1170;
									assign node1170 = (inp[2]) ? node1172 : 3'b110;
										assign node1172 = (inp[3]) ? 3'b010 : node1173;
											assign node1173 = (inp[4]) ? 3'b010 : 3'b110;
									assign node1177 = (inp[2]) ? node1179 : 3'b010;
										assign node1179 = (inp[4]) ? 3'b100 : node1180;
											assign node1180 = (inp[3]) ? 3'b100 : 3'b010;
								assign node1184 = (inp[11]) ? node1194 : node1185;
									assign node1185 = (inp[2]) ? node1187 : 3'b001;
										assign node1187 = (inp[3]) ? 3'b110 : node1188;
											assign node1188 = (inp[4]) ? node1190 : 3'b001;
												assign node1190 = (inp[5]) ? 3'b110 : 3'b001;
									assign node1194 = (inp[2]) ? node1196 : 3'b110;
										assign node1196 = (inp[3]) ? 3'b010 : node1197;
											assign node1197 = (inp[5]) ? node1199 : 3'b110;
												assign node1199 = (inp[4]) ? 3'b010 : 3'b110;
							assign node1203 = (inp[8]) ? node1219 : node1204;
								assign node1204 = (inp[11]) ? node1212 : node1205;
									assign node1205 = (inp[2]) ? 3'b100 : node1206;
										assign node1206 = (inp[4]) ? node1208 : 3'b010;
											assign node1208 = (inp[3]) ? 3'b100 : 3'b010;
									assign node1212 = (inp[2]) ? 3'b000 : node1213;
										assign node1213 = (inp[3]) ? node1215 : 3'b100;
											assign node1215 = (inp[4]) ? 3'b000 : 3'b100;
								assign node1219 = (inp[11]) ? node1227 : node1220;
									assign node1220 = (inp[2]) ? 3'b010 : node1221;
										assign node1221 = (inp[4]) ? node1223 : 3'b110;
											assign node1223 = (inp[3]) ? 3'b010 : 3'b110;
									assign node1227 = (inp[2]) ? 3'b100 : node1228;
										assign node1228 = (inp[4]) ? node1230 : 3'b010;
											assign node1230 = (inp[3]) ? node1232 : 3'b010;
												assign node1232 = (inp[5]) ? 3'b100 : 3'b010;
				assign node1236 = (inp[7]) ? node1264 : node1237;
					assign node1237 = (inp[8]) ? node1239 : 3'b000;
						assign node1239 = (inp[10]) ? 3'b000 : node1240;
							assign node1240 = (inp[1]) ? 3'b000 : node1241;
								assign node1241 = (inp[11]) ? node1255 : node1242;
									assign node1242 = (inp[2]) ? node1250 : node1243;
										assign node1243 = (inp[3]) ? 3'b100 : node1244;
											assign node1244 = (inp[4]) ? 3'b100 : node1245;
												assign node1245 = (inp[5]) ? 3'b100 : 3'b010;
										assign node1250 = (inp[4]) ? node1252 : 3'b100;
											assign node1252 = (inp[3]) ? 3'b000 : 3'b100;
									assign node1255 = (inp[3]) ? 3'b000 : node1256;
										assign node1256 = (inp[4]) ? 3'b000 : node1257;
											assign node1257 = (inp[2]) ? 3'b000 : 3'b100;
					assign node1264 = (inp[10]) ? node1346 : node1265;
						assign node1265 = (inp[1]) ? node1321 : node1266;
							assign node1266 = (inp[11]) ? node1294 : node1267;
								assign node1267 = (inp[8]) ? node1279 : node1268;
									assign node1268 = (inp[3]) ? node1274 : node1269;
										assign node1269 = (inp[4]) ? 3'b010 : node1270;
											assign node1270 = (inp[2]) ? 3'b010 : 3'b110;
										assign node1274 = (inp[2]) ? node1276 : 3'b010;
											assign node1276 = (inp[4]) ? 3'b100 : 3'b010;
									assign node1279 = (inp[2]) ? node1287 : node1280;
										assign node1280 = (inp[3]) ? 3'b110 : node1281;
											assign node1281 = (inp[5]) ? node1283 : 3'b001;
												assign node1283 = (inp[4]) ? 3'b110 : 3'b001;
										assign node1287 = (inp[4]) ? node1289 : 3'b110;
											assign node1289 = (inp[5]) ? node1291 : 3'b110;
												assign node1291 = (inp[3]) ? 3'b010 : 3'b110;
								assign node1294 = (inp[8]) ? node1308 : node1295;
									assign node1295 = (inp[3]) ? node1303 : node1296;
										assign node1296 = (inp[2]) ? 3'b100 : node1297;
											assign node1297 = (inp[5]) ? node1299 : 3'b010;
												assign node1299 = (inp[4]) ? 3'b100 : 3'b010;
										assign node1303 = (inp[4]) ? node1305 : 3'b100;
											assign node1305 = (inp[2]) ? 3'b000 : 3'b100;
									assign node1308 = (inp[2]) ? node1316 : node1309;
										assign node1309 = (inp[3]) ? 3'b010 : node1310;
											assign node1310 = (inp[5]) ? node1312 : 3'b110;
												assign node1312 = (inp[4]) ? 3'b010 : 3'b110;
										assign node1316 = (inp[5]) ? node1318 : 3'b010;
											assign node1318 = (inp[3]) ? 3'b100 : 3'b010;
							assign node1321 = (inp[8]) ? node1331 : node1322;
								assign node1322 = (inp[11]) ? 3'b000 : node1323;
									assign node1323 = (inp[2]) ? node1325 : 3'b100;
										assign node1325 = (inp[3]) ? 3'b000 : node1326;
											assign node1326 = (inp[4]) ? 3'b000 : 3'b100;
								assign node1331 = (inp[11]) ? node1337 : node1332;
									assign node1332 = (inp[3]) ? node1334 : 3'b010;
										assign node1334 = (inp[2]) ? 3'b100 : 3'b010;
									assign node1337 = (inp[2]) ? node1343 : node1338;
										assign node1338 = (inp[3]) ? 3'b100 : node1339;
											assign node1339 = (inp[4]) ? 3'b100 : 3'b010;
										assign node1343 = (inp[3]) ? 3'b000 : 3'b100;
						assign node1346 = (inp[1]) ? 3'b000 : node1347;
							assign node1347 = (inp[8]) ? node1359 : node1348;
								assign node1348 = (inp[11]) ? 3'b000 : node1349;
									assign node1349 = (inp[2]) ? 3'b000 : node1350;
										assign node1350 = (inp[3]) ? 3'b000 : node1351;
											assign node1351 = (inp[4]) ? node1353 : 3'b100;
												assign node1353 = (inp[5]) ? 3'b000 : 3'b100;
								assign node1359 = (inp[11]) ? node1365 : node1360;
									assign node1360 = (inp[3]) ? 3'b100 : node1361;
										assign node1361 = (inp[2]) ? 3'b100 : 3'b010;
									assign node1365 = (inp[3]) ? 3'b000 : node1366;
										assign node1366 = (inp[2]) ? 3'b000 : 3'b100;

endmodule