module dtc_split25_bm65 (
	input  wire [16-1:0] inp,
	output wire [4-1:0] outp
);

	wire [4-1:0] node1;
	wire [4-1:0] node2;
	wire [4-1:0] node3;
	wire [4-1:0] node4;
	wire [4-1:0] node5;
	wire [4-1:0] node6;
	wire [4-1:0] node7;
	wire [4-1:0] node8;
	wire [4-1:0] node9;
	wire [4-1:0] node10;
	wire [4-1:0] node11;
	wire [4-1:0] node12;
	wire [4-1:0] node16;
	wire [4-1:0] node18;
	wire [4-1:0] node21;
	wire [4-1:0] node22;
	wire [4-1:0] node25;
	wire [4-1:0] node27;
	wire [4-1:0] node29;
	wire [4-1:0] node32;
	wire [4-1:0] node33;
	wire [4-1:0] node34;
	wire [4-1:0] node35;
	wire [4-1:0] node37;
	wire [4-1:0] node41;
	wire [4-1:0] node42;
	wire [4-1:0] node44;
	wire [4-1:0] node47;
	wire [4-1:0] node49;
	wire [4-1:0] node50;
	wire [4-1:0] node54;
	wire [4-1:0] node55;
	wire [4-1:0] node56;
	wire [4-1:0] node57;
	wire [4-1:0] node59;
	wire [4-1:0] node64;
	wire [4-1:0] node65;
	wire [4-1:0] node66;
	wire [4-1:0] node70;
	wire [4-1:0] node73;
	wire [4-1:0] node74;
	wire [4-1:0] node75;
	wire [4-1:0] node76;
	wire [4-1:0] node77;
	wire [4-1:0] node78;
	wire [4-1:0] node84;
	wire [4-1:0] node85;
	wire [4-1:0] node86;
	wire [4-1:0] node87;
	wire [4-1:0] node89;
	wire [4-1:0] node93;
	wire [4-1:0] node96;
	wire [4-1:0] node97;
	wire [4-1:0] node98;
	wire [4-1:0] node102;
	wire [4-1:0] node103;
	wire [4-1:0] node107;
	wire [4-1:0] node108;
	wire [4-1:0] node109;
	wire [4-1:0] node110;
	wire [4-1:0] node112;
	wire [4-1:0] node115;
	wire [4-1:0] node117;
	wire [4-1:0] node120;
	wire [4-1:0] node121;
	wire [4-1:0] node123;
	wire [4-1:0] node126;
	wire [4-1:0] node127;
	wire [4-1:0] node131;
	wire [4-1:0] node132;
	wire [4-1:0] node133;
	wire [4-1:0] node136;
	wire [4-1:0] node138;
	wire [4-1:0] node141;
	wire [4-1:0] node143;
	wire [4-1:0] node145;
	wire [4-1:0] node149;
	wire [4-1:0] node150;
	wire [4-1:0] node151;
	wire [4-1:0] node152;
	wire [4-1:0] node153;
	wire [4-1:0] node154;
	wire [4-1:0] node155;
	wire [4-1:0] node156;
	wire [4-1:0] node160;
	wire [4-1:0] node163;
	wire [4-1:0] node164;
	wire [4-1:0] node168;
	wire [4-1:0] node169;
	wire [4-1:0] node170;
	wire [4-1:0] node172;
	wire [4-1:0] node176;
	wire [4-1:0] node178;
	wire [4-1:0] node181;
	wire [4-1:0] node182;
	wire [4-1:0] node183;
	wire [4-1:0] node186;
	wire [4-1:0] node189;
	wire [4-1:0] node190;
	wire [4-1:0] node191;
	wire [4-1:0] node194;
	wire [4-1:0] node195;
	wire [4-1:0] node197;
	wire [4-1:0] node201;
	wire [4-1:0] node204;
	wire [4-1:0] node205;
	wire [4-1:0] node206;
	wire [4-1:0] node207;
	wire [4-1:0] node209;
	wire [4-1:0] node210;
	wire [4-1:0] node214;
	wire [4-1:0] node215;
	wire [4-1:0] node217;
	wire [4-1:0] node220;
	wire [4-1:0] node222;
	wire [4-1:0] node225;
	wire [4-1:0] node226;
	wire [4-1:0] node227;
	wire [4-1:0] node229;
	wire [4-1:0] node232;
	wire [4-1:0] node233;
	wire [4-1:0] node234;
	wire [4-1:0] node239;
	wire [4-1:0] node240;
	wire [4-1:0] node242;
	wire [4-1:0] node244;
	wire [4-1:0] node247;
	wire [4-1:0] node250;
	wire [4-1:0] node251;
	wire [4-1:0] node252;
	wire [4-1:0] node253;
	wire [4-1:0] node254;
	wire [4-1:0] node258;
	wire [4-1:0] node260;
	wire [4-1:0] node263;
	wire [4-1:0] node264;
	wire [4-1:0] node265;
	wire [4-1:0] node266;
	wire [4-1:0] node272;
	wire [4-1:0] node273;
	wire [4-1:0] node274;
	wire [4-1:0] node275;
	wire [4-1:0] node279;
	wire [4-1:0] node280;
	wire [4-1:0] node281;
	wire [4-1:0] node286;
	wire [4-1:0] node288;
	wire [4-1:0] node291;
	wire [4-1:0] node292;
	wire [4-1:0] node293;
	wire [4-1:0] node294;
	wire [4-1:0] node295;
	wire [4-1:0] node296;
	wire [4-1:0] node297;
	wire [4-1:0] node302;
	wire [4-1:0] node304;
	wire [4-1:0] node305;
	wire [4-1:0] node309;
	wire [4-1:0] node310;
	wire [4-1:0] node312;
	wire [4-1:0] node315;
	wire [4-1:0] node316;
	wire [4-1:0] node318;
	wire [4-1:0] node322;
	wire [4-1:0] node323;
	wire [4-1:0] node324;
	wire [4-1:0] node326;
	wire [4-1:0] node329;
	wire [4-1:0] node330;
	wire [4-1:0] node333;
	wire [4-1:0] node336;
	wire [4-1:0] node337;
	wire [4-1:0] node338;
	wire [4-1:0] node342;
	wire [4-1:0] node343;
	wire [4-1:0] node344;
	wire [4-1:0] node349;
	wire [4-1:0] node350;
	wire [4-1:0] node351;
	wire [4-1:0] node352;
	wire [4-1:0] node353;
	wire [4-1:0] node357;
	wire [4-1:0] node359;
	wire [4-1:0] node362;
	wire [4-1:0] node363;
	wire [4-1:0] node364;
	wire [4-1:0] node366;
	wire [4-1:0] node367;
	wire [4-1:0] node371;
	wire [4-1:0] node374;
	wire [4-1:0] node376;
	wire [4-1:0] node379;
	wire [4-1:0] node380;
	wire [4-1:0] node381;
	wire [4-1:0] node382;
	wire [4-1:0] node386;
	wire [4-1:0] node389;
	wire [4-1:0] node390;
	wire [4-1:0] node392;
	wire [4-1:0] node393;
	wire [4-1:0] node396;
	wire [4-1:0] node399;
	wire [4-1:0] node400;
	wire [4-1:0] node403;
	wire [4-1:0] node404;
	wire [4-1:0] node409;
	wire [4-1:0] node410;
	wire [4-1:0] node411;
	wire [4-1:0] node413;
	wire [4-1:0] node414;
	wire [4-1:0] node415;
	wire [4-1:0] node416;
	wire [4-1:0] node417;
	wire [4-1:0] node418;
	wire [4-1:0] node419;
	wire [4-1:0] node423;
	wire [4-1:0] node426;
	wire [4-1:0] node428;
	wire [4-1:0] node430;
	wire [4-1:0] node434;
	wire [4-1:0] node435;
	wire [4-1:0] node436;
	wire [4-1:0] node438;
	wire [4-1:0] node440;
	wire [4-1:0] node443;
	wire [4-1:0] node444;
	wire [4-1:0] node446;
	wire [4-1:0] node448;
	wire [4-1:0] node451;
	wire [4-1:0] node454;
	wire [4-1:0] node455;
	wire [4-1:0] node456;
	wire [4-1:0] node459;
	wire [4-1:0] node460;
	wire [4-1:0] node462;
	wire [4-1:0] node466;
	wire [4-1:0] node467;
	wire [4-1:0] node469;
	wire [4-1:0] node472;
	wire [4-1:0] node476;
	wire [4-1:0] node477;
	wire [4-1:0] node478;
	wire [4-1:0] node479;
	wire [4-1:0] node480;
	wire [4-1:0] node481;
	wire [4-1:0] node482;
	wire [4-1:0] node483;
	wire [4-1:0] node487;
	wire [4-1:0] node490;
	wire [4-1:0] node492;
	wire [4-1:0] node495;
	wire [4-1:0] node496;
	wire [4-1:0] node497;
	wire [4-1:0] node499;
	wire [4-1:0] node503;
	wire [4-1:0] node504;
	wire [4-1:0] node505;
	wire [4-1:0] node506;
	wire [4-1:0] node510;
	wire [4-1:0] node513;
	wire [4-1:0] node516;
	wire [4-1:0] node517;
	wire [4-1:0] node518;
	wire [4-1:0] node519;
	wire [4-1:0] node521;
	wire [4-1:0] node522;
	wire [4-1:0] node525;
	wire [4-1:0] node528;
	wire [4-1:0] node529;
	wire [4-1:0] node533;
	wire [4-1:0] node534;
	wire [4-1:0] node538;
	wire [4-1:0] node539;
	wire [4-1:0] node540;
	wire [4-1:0] node541;
	wire [4-1:0] node544;
	wire [4-1:0] node547;
	wire [4-1:0] node549;
	wire [4-1:0] node551;
	wire [4-1:0] node554;
	wire [4-1:0] node555;
	wire [4-1:0] node558;
	wire [4-1:0] node560;
	wire [4-1:0] node563;
	wire [4-1:0] node564;
	wire [4-1:0] node565;
	wire [4-1:0] node566;
	wire [4-1:0] node567;
	wire [4-1:0] node568;
	wire [4-1:0] node569;
	wire [4-1:0] node575;
	wire [4-1:0] node576;
	wire [4-1:0] node577;
	wire [4-1:0] node579;
	wire [4-1:0] node582;
	wire [4-1:0] node586;
	wire [4-1:0] node587;
	wire [4-1:0] node588;
	wire [4-1:0] node589;
	wire [4-1:0] node593;
	wire [4-1:0] node594;
	wire [4-1:0] node598;
	wire [4-1:0] node599;
	wire [4-1:0] node601;
	wire [4-1:0] node605;
	wire [4-1:0] node606;
	wire [4-1:0] node607;
	wire [4-1:0] node608;
	wire [4-1:0] node611;
	wire [4-1:0] node612;
	wire [4-1:0] node616;
	wire [4-1:0] node617;
	wire [4-1:0] node621;
	wire [4-1:0] node622;
	wire [4-1:0] node623;
	wire [4-1:0] node624;
	wire [4-1:0] node629;
	wire [4-1:0] node630;
	wire [4-1:0] node633;
	wire [4-1:0] node634;
	wire [4-1:0] node635;
	wire [4-1:0] node640;
	wire [4-1:0] node642;
	wire [4-1:0] node643;
	wire [4-1:0] node644;
	wire [4-1:0] node645;
	wire [4-1:0] node646;
	wire [4-1:0] node648;
	wire [4-1:0] node651;
	wire [4-1:0] node652;
	wire [4-1:0] node656;
	wire [4-1:0] node660;
	wire [4-1:0] node661;
	wire [4-1:0] node662;
	wire [4-1:0] node663;
	wire [4-1:0] node665;
	wire [4-1:0] node669;
	wire [4-1:0] node670;
	wire [4-1:0] node672;
	wire [4-1:0] node676;
	wire [4-1:0] node677;
	wire [4-1:0] node679;
	wire [4-1:0] node681;
	wire [4-1:0] node684;
	wire [4-1:0] node685;
	wire [4-1:0] node687;
	wire [4-1:0] node690;
	wire [4-1:0] node694;
	wire [4-1:0] node695;
	wire [4-1:0] node696;
	wire [4-1:0] node697;
	wire [4-1:0] node698;
	wire [4-1:0] node699;
	wire [4-1:0] node700;
	wire [4-1:0] node701;
	wire [4-1:0] node702;
	wire [4-1:0] node703;
	wire [4-1:0] node705;
	wire [4-1:0] node708;
	wire [4-1:0] node710;
	wire [4-1:0] node713;
	wire [4-1:0] node714;
	wire [4-1:0] node717;
	wire [4-1:0] node719;
	wire [4-1:0] node722;
	wire [4-1:0] node723;
	wire [4-1:0] node724;
	wire [4-1:0] node726;
	wire [4-1:0] node727;
	wire [4-1:0] node731;
	wire [4-1:0] node734;
	wire [4-1:0] node735;
	wire [4-1:0] node736;
	wire [4-1:0] node741;
	wire [4-1:0] node742;
	wire [4-1:0] node743;
	wire [4-1:0] node744;
	wire [4-1:0] node745;
	wire [4-1:0] node749;
	wire [4-1:0] node752;
	wire [4-1:0] node754;
	wire [4-1:0] node755;
	wire [4-1:0] node759;
	wire [4-1:0] node760;
	wire [4-1:0] node762;
	wire [4-1:0] node763;
	wire [4-1:0] node765;
	wire [4-1:0] node768;
	wire [4-1:0] node770;
	wire [4-1:0] node774;
	wire [4-1:0] node775;
	wire [4-1:0] node776;
	wire [4-1:0] node777;
	wire [4-1:0] node778;
	wire [4-1:0] node779;
	wire [4-1:0] node780;
	wire [4-1:0] node783;
	wire [4-1:0] node787;
	wire [4-1:0] node788;
	wire [4-1:0] node791;
	wire [4-1:0] node794;
	wire [4-1:0] node797;
	wire [4-1:0] node798;
	wire [4-1:0] node799;
	wire [4-1:0] node801;
	wire [4-1:0] node803;
	wire [4-1:0] node806;
	wire [4-1:0] node808;
	wire [4-1:0] node811;
	wire [4-1:0] node812;
	wire [4-1:0] node815;
	wire [4-1:0] node818;
	wire [4-1:0] node819;
	wire [4-1:0] node820;
	wire [4-1:0] node821;
	wire [4-1:0] node822;
	wire [4-1:0] node824;
	wire [4-1:0] node827;
	wire [4-1:0] node830;
	wire [4-1:0] node831;
	wire [4-1:0] node835;
	wire [4-1:0] node836;
	wire [4-1:0] node837;
	wire [4-1:0] node839;
	wire [4-1:0] node842;
	wire [4-1:0] node843;
	wire [4-1:0] node846;
	wire [4-1:0] node849;
	wire [4-1:0] node850;
	wire [4-1:0] node854;
	wire [4-1:0] node855;
	wire [4-1:0] node856;
	wire [4-1:0] node858;
	wire [4-1:0] node861;
	wire [4-1:0] node864;
	wire [4-1:0] node866;
	wire [4-1:0] node867;
	wire [4-1:0] node870;
	wire [4-1:0] node873;
	wire [4-1:0] node874;
	wire [4-1:0] node875;
	wire [4-1:0] node876;
	wire [4-1:0] node877;
	wire [4-1:0] node878;
	wire [4-1:0] node881;
	wire [4-1:0] node882;
	wire [4-1:0] node886;
	wire [4-1:0] node888;
	wire [4-1:0] node889;
	wire [4-1:0] node892;
	wire [4-1:0] node895;
	wire [4-1:0] node896;
	wire [4-1:0] node898;
	wire [4-1:0] node901;
	wire [4-1:0] node903;
	wire [4-1:0] node904;
	wire [4-1:0] node906;
	wire [4-1:0] node909;
	wire [4-1:0] node912;
	wire [4-1:0] node913;
	wire [4-1:0] node914;
	wire [4-1:0] node915;
	wire [4-1:0] node919;
	wire [4-1:0] node920;
	wire [4-1:0] node922;
	wire [4-1:0] node924;
	wire [4-1:0] node927;
	wire [4-1:0] node928;
	wire [4-1:0] node930;
	wire [4-1:0] node933;
	wire [4-1:0] node934;
	wire [4-1:0] node938;
	wire [4-1:0] node939;
	wire [4-1:0] node940;
	wire [4-1:0] node943;
	wire [4-1:0] node946;
	wire [4-1:0] node947;
	wire [4-1:0] node950;
	wire [4-1:0] node952;
	wire [4-1:0] node955;
	wire [4-1:0] node956;
	wire [4-1:0] node957;
	wire [4-1:0] node958;
	wire [4-1:0] node959;
	wire [4-1:0] node963;
	wire [4-1:0] node965;
	wire [4-1:0] node966;
	wire [4-1:0] node969;
	wire [4-1:0] node970;
	wire [4-1:0] node972;
	wire [4-1:0] node975;
	wire [4-1:0] node978;
	wire [4-1:0] node979;
	wire [4-1:0] node981;
	wire [4-1:0] node983;
	wire [4-1:0] node986;
	wire [4-1:0] node987;
	wire [4-1:0] node988;
	wire [4-1:0] node992;
	wire [4-1:0] node995;
	wire [4-1:0] node996;
	wire [4-1:0] node997;
	wire [4-1:0] node998;
	wire [4-1:0] node1000;
	wire [4-1:0] node1003;
	wire [4-1:0] node1006;
	wire [4-1:0] node1007;
	wire [4-1:0] node1010;
	wire [4-1:0] node1012;
	wire [4-1:0] node1014;
	wire [4-1:0] node1015;
	wire [4-1:0] node1019;
	wire [4-1:0] node1020;
	wire [4-1:0] node1022;
	wire [4-1:0] node1023;
	wire [4-1:0] node1024;
	wire [4-1:0] node1028;
	wire [4-1:0] node1031;
	wire [4-1:0] node1034;
	wire [4-1:0] node1035;
	wire [4-1:0] node1036;
	wire [4-1:0] node1037;
	wire [4-1:0] node1038;
	wire [4-1:0] node1039;
	wire [4-1:0] node1040;
	wire [4-1:0] node1041;
	wire [4-1:0] node1045;
	wire [4-1:0] node1047;
	wire [4-1:0] node1050;
	wire [4-1:0] node1051;
	wire [4-1:0] node1052;
	wire [4-1:0] node1056;
	wire [4-1:0] node1059;
	wire [4-1:0] node1060;
	wire [4-1:0] node1061;
	wire [4-1:0] node1064;
	wire [4-1:0] node1067;
	wire [4-1:0] node1068;
	wire [4-1:0] node1071;
	wire [4-1:0] node1072;
	wire [4-1:0] node1075;
	wire [4-1:0] node1078;
	wire [4-1:0] node1079;
	wire [4-1:0] node1080;
	wire [4-1:0] node1082;
	wire [4-1:0] node1083;
	wire [4-1:0] node1087;
	wire [4-1:0] node1088;
	wire [4-1:0] node1090;
	wire [4-1:0] node1093;
	wire [4-1:0] node1094;
	wire [4-1:0] node1098;
	wire [4-1:0] node1099;
	wire [4-1:0] node1101;
	wire [4-1:0] node1103;
	wire [4-1:0] node1106;
	wire [4-1:0] node1108;
	wire [4-1:0] node1111;
	wire [4-1:0] node1112;
	wire [4-1:0] node1113;
	wire [4-1:0] node1114;
	wire [4-1:0] node1115;
	wire [4-1:0] node1116;
	wire [4-1:0] node1117;
	wire [4-1:0] node1120;
	wire [4-1:0] node1122;
	wire [4-1:0] node1125;
	wire [4-1:0] node1128;
	wire [4-1:0] node1130;
	wire [4-1:0] node1133;
	wire [4-1:0] node1134;
	wire [4-1:0] node1138;
	wire [4-1:0] node1139;
	wire [4-1:0] node1141;
	wire [4-1:0] node1142;
	wire [4-1:0] node1146;
	wire [4-1:0] node1147;
	wire [4-1:0] node1149;
	wire [4-1:0] node1152;
	wire [4-1:0] node1153;
	wire [4-1:0] node1157;
	wire [4-1:0] node1158;
	wire [4-1:0] node1159;
	wire [4-1:0] node1160;
	wire [4-1:0] node1163;
	wire [4-1:0] node1166;
	wire [4-1:0] node1167;
	wire [4-1:0] node1168;
	wire [4-1:0] node1171;
	wire [4-1:0] node1173;
	wire [4-1:0] node1176;
	wire [4-1:0] node1179;
	wire [4-1:0] node1180;
	wire [4-1:0] node1181;
	wire [4-1:0] node1184;
	wire [4-1:0] node1187;
	wire [4-1:0] node1189;
	wire [4-1:0] node1190;
	wire [4-1:0] node1192;
	wire [4-1:0] node1196;
	wire [4-1:0] node1197;
	wire [4-1:0] node1198;
	wire [4-1:0] node1199;
	wire [4-1:0] node1201;
	wire [4-1:0] node1202;
	wire [4-1:0] node1206;
	wire [4-1:0] node1207;
	wire [4-1:0] node1208;
	wire [4-1:0] node1211;
	wire [4-1:0] node1212;
	wire [4-1:0] node1216;
	wire [4-1:0] node1218;
	wire [4-1:0] node1219;
	wire [4-1:0] node1222;
	wire [4-1:0] node1224;
	wire [4-1:0] node1227;
	wire [4-1:0] node1228;
	wire [4-1:0] node1229;
	wire [4-1:0] node1230;
	wire [4-1:0] node1233;
	wire [4-1:0] node1234;
	wire [4-1:0] node1238;
	wire [4-1:0] node1239;
	wire [4-1:0] node1240;
	wire [4-1:0] node1244;
	wire [4-1:0] node1245;
	wire [4-1:0] node1246;
	wire [4-1:0] node1250;
	wire [4-1:0] node1253;
	wire [4-1:0] node1254;
	wire [4-1:0] node1255;
	wire [4-1:0] node1256;
	wire [4-1:0] node1258;
	wire [4-1:0] node1263;
	wire [4-1:0] node1264;
	wire [4-1:0] node1265;
	wire [4-1:0] node1267;
	wire [4-1:0] node1271;
	wire [4-1:0] node1272;
	wire [4-1:0] node1275;
	wire [4-1:0] node1277;
	wire [4-1:0] node1280;
	wire [4-1:0] node1281;
	wire [4-1:0] node1282;
	wire [4-1:0] node1283;
	wire [4-1:0] node1284;
	wire [4-1:0] node1285;
	wire [4-1:0] node1288;
	wire [4-1:0] node1291;
	wire [4-1:0] node1294;
	wire [4-1:0] node1295;
	wire [4-1:0] node1296;
	wire [4-1:0] node1299;
	wire [4-1:0] node1300;
	wire [4-1:0] node1304;
	wire [4-1:0] node1305;
	wire [4-1:0] node1308;
	wire [4-1:0] node1309;
	wire [4-1:0] node1313;
	wire [4-1:0] node1314;
	wire [4-1:0] node1317;
	wire [4-1:0] node1318;
	wire [4-1:0] node1321;
	wire [4-1:0] node1322;
	wire [4-1:0] node1325;
	wire [4-1:0] node1328;
	wire [4-1:0] node1329;
	wire [4-1:0] node1331;
	wire [4-1:0] node1332;
	wire [4-1:0] node1333;
	wire [4-1:0] node1337;
	wire [4-1:0] node1340;
	wire [4-1:0] node1341;
	wire [4-1:0] node1342;
	wire [4-1:0] node1344;
	wire [4-1:0] node1347;
	wire [4-1:0] node1350;
	wire [4-1:0] node1351;
	wire [4-1:0] node1355;
	wire [4-1:0] node1356;
	wire [4-1:0] node1357;
	wire [4-1:0] node1358;
	wire [4-1:0] node1359;
	wire [4-1:0] node1360;
	wire [4-1:0] node1361;
	wire [4-1:0] node1363;
	wire [4-1:0] node1364;
	wire [4-1:0] node1366;
	wire [4-1:0] node1369;
	wire [4-1:0] node1370;
	wire [4-1:0] node1373;
	wire [4-1:0] node1376;
	wire [4-1:0] node1378;
	wire [4-1:0] node1381;
	wire [4-1:0] node1382;
	wire [4-1:0] node1383;
	wire [4-1:0] node1386;
	wire [4-1:0] node1387;
	wire [4-1:0] node1391;
	wire [4-1:0] node1392;
	wire [4-1:0] node1393;
	wire [4-1:0] node1397;
	wire [4-1:0] node1398;
	wire [4-1:0] node1400;
	wire [4-1:0] node1402;
	wire [4-1:0] node1406;
	wire [4-1:0] node1407;
	wire [4-1:0] node1408;
	wire [4-1:0] node1409;
	wire [4-1:0] node1413;
	wire [4-1:0] node1414;
	wire [4-1:0] node1418;
	wire [4-1:0] node1419;
	wire [4-1:0] node1421;
	wire [4-1:0] node1424;
	wire [4-1:0] node1425;
	wire [4-1:0] node1428;
	wire [4-1:0] node1429;
	wire [4-1:0] node1433;
	wire [4-1:0] node1434;
	wire [4-1:0] node1435;
	wire [4-1:0] node1436;
	wire [4-1:0] node1437;
	wire [4-1:0] node1439;
	wire [4-1:0] node1442;
	wire [4-1:0] node1446;
	wire [4-1:0] node1447;
	wire [4-1:0] node1448;
	wire [4-1:0] node1450;
	wire [4-1:0] node1454;
	wire [4-1:0] node1455;
	wire [4-1:0] node1456;
	wire [4-1:0] node1460;
	wire [4-1:0] node1461;
	wire [4-1:0] node1465;
	wire [4-1:0] node1466;
	wire [4-1:0] node1467;
	wire [4-1:0] node1468;
	wire [4-1:0] node1470;
	wire [4-1:0] node1472;
	wire [4-1:0] node1475;
	wire [4-1:0] node1476;
	wire [4-1:0] node1480;
	wire [4-1:0] node1482;
	wire [4-1:0] node1483;
	wire [4-1:0] node1484;
	wire [4-1:0] node1489;
	wire [4-1:0] node1490;
	wire [4-1:0] node1492;
	wire [4-1:0] node1493;
	wire [4-1:0] node1497;
	wire [4-1:0] node1498;
	wire [4-1:0] node1499;
	wire [4-1:0] node1502;
	wire [4-1:0] node1507;
	wire [4-1:0] node1508;
	wire [4-1:0] node1510;
	wire [4-1:0] node1511;
	wire [4-1:0] node1512;
	wire [4-1:0] node1513;
	wire [4-1:0] node1515;
	wire [4-1:0] node1518;
	wire [4-1:0] node1519;
	wire [4-1:0] node1524;
	wire [4-1:0] node1525;
	wire [4-1:0] node1526;
	wire [4-1:0] node1527;
	wire [4-1:0] node1530;
	wire [4-1:0] node1533;
	wire [4-1:0] node1535;
	wire [4-1:0] node1538;
	wire [4-1:0] node1539;
	wire [4-1:0] node1541;
	wire [4-1:0] node1543;
	wire [4-1:0] node1544;
	wire [4-1:0] node1548;
	wire [4-1:0] node1549;
	wire [4-1:0] node1552;
	wire [4-1:0] node1554;
	wire [4-1:0] node1558;
	wire [4-1:0] node1559;
	wire [4-1:0] node1560;
	wire [4-1:0] node1561;
	wire [4-1:0] node1562;
	wire [4-1:0] node1563;
	wire [4-1:0] node1564;
	wire [4-1:0] node1565;
	wire [4-1:0] node1566;
	wire [4-1:0] node1567;
	wire [4-1:0] node1569;
	wire [4-1:0] node1571;
	wire [4-1:0] node1574;
	wire [4-1:0] node1577;
	wire [4-1:0] node1579;
	wire [4-1:0] node1582;
	wire [4-1:0] node1583;
	wire [4-1:0] node1586;
	wire [4-1:0] node1587;
	wire [4-1:0] node1591;
	wire [4-1:0] node1592;
	wire [4-1:0] node1593;
	wire [4-1:0] node1596;
	wire [4-1:0] node1597;
	wire [4-1:0] node1598;
	wire [4-1:0] node1603;
	wire [4-1:0] node1604;
	wire [4-1:0] node1605;
	wire [4-1:0] node1607;
	wire [4-1:0] node1610;
	wire [4-1:0] node1612;
	wire [4-1:0] node1615;
	wire [4-1:0] node1617;
	wire [4-1:0] node1620;
	wire [4-1:0] node1621;
	wire [4-1:0] node1622;
	wire [4-1:0] node1623;
	wire [4-1:0] node1625;
	wire [4-1:0] node1628;
	wire [4-1:0] node1631;
	wire [4-1:0] node1633;
	wire [4-1:0] node1636;
	wire [4-1:0] node1637;
	wire [4-1:0] node1638;
	wire [4-1:0] node1639;
	wire [4-1:0] node1644;
	wire [4-1:0] node1645;
	wire [4-1:0] node1646;
	wire [4-1:0] node1650;
	wire [4-1:0] node1653;
	wire [4-1:0] node1654;
	wire [4-1:0] node1655;
	wire [4-1:0] node1656;
	wire [4-1:0] node1658;
	wire [4-1:0] node1659;
	wire [4-1:0] node1662;
	wire [4-1:0] node1665;
	wire [4-1:0] node1667;
	wire [4-1:0] node1669;
	wire [4-1:0] node1672;
	wire [4-1:0] node1673;
	wire [4-1:0] node1674;
	wire [4-1:0] node1678;
	wire [4-1:0] node1679;
	wire [4-1:0] node1682;
	wire [4-1:0] node1684;
	wire [4-1:0] node1686;
	wire [4-1:0] node1689;
	wire [4-1:0] node1690;
	wire [4-1:0] node1691;
	wire [4-1:0] node1693;
	wire [4-1:0] node1695;
	wire [4-1:0] node1696;
	wire [4-1:0] node1698;
	wire [4-1:0] node1702;
	wire [4-1:0] node1703;
	wire [4-1:0] node1706;
	wire [4-1:0] node1709;
	wire [4-1:0] node1710;
	wire [4-1:0] node1712;
	wire [4-1:0] node1714;
	wire [4-1:0] node1717;
	wire [4-1:0] node1718;
	wire [4-1:0] node1720;
	wire [4-1:0] node1723;
	wire [4-1:0] node1726;
	wire [4-1:0] node1727;
	wire [4-1:0] node1728;
	wire [4-1:0] node1729;
	wire [4-1:0] node1730;
	wire [4-1:0] node1731;
	wire [4-1:0] node1732;
	wire [4-1:0] node1733;
	wire [4-1:0] node1738;
	wire [4-1:0] node1740;
	wire [4-1:0] node1743;
	wire [4-1:0] node1745;
	wire [4-1:0] node1746;
	wire [4-1:0] node1747;
	wire [4-1:0] node1750;
	wire [4-1:0] node1754;
	wire [4-1:0] node1755;
	wire [4-1:0] node1756;
	wire [4-1:0] node1757;
	wire [4-1:0] node1758;
	wire [4-1:0] node1762;
	wire [4-1:0] node1763;
	wire [4-1:0] node1767;
	wire [4-1:0] node1768;
	wire [4-1:0] node1772;
	wire [4-1:0] node1774;
	wire [4-1:0] node1776;
	wire [4-1:0] node1779;
	wire [4-1:0] node1780;
	wire [4-1:0] node1781;
	wire [4-1:0] node1782;
	wire [4-1:0] node1783;
	wire [4-1:0] node1786;
	wire [4-1:0] node1789;
	wire [4-1:0] node1791;
	wire [4-1:0] node1794;
	wire [4-1:0] node1795;
	wire [4-1:0] node1798;
	wire [4-1:0] node1799;
	wire [4-1:0] node1802;
	wire [4-1:0] node1805;
	wire [4-1:0] node1806;
	wire [4-1:0] node1810;
	wire [4-1:0] node1811;
	wire [4-1:0] node1812;
	wire [4-1:0] node1813;
	wire [4-1:0] node1815;
	wire [4-1:0] node1816;
	wire [4-1:0] node1818;
	wire [4-1:0] node1819;
	wire [4-1:0] node1824;
	wire [4-1:0] node1825;
	wire [4-1:0] node1826;
	wire [4-1:0] node1833;
	wire [4-1:0] node1834;
	wire [4-1:0] node1835;
	wire [4-1:0] node1836;
	wire [4-1:0] node1837;
	wire [4-1:0] node1838;
	wire [4-1:0] node1839;
	wire [4-1:0] node1841;
	wire [4-1:0] node1844;
	wire [4-1:0] node1846;
	wire [4-1:0] node1847;
	wire [4-1:0] node1851;
	wire [4-1:0] node1852;
	wire [4-1:0] node1854;
	wire [4-1:0] node1855;
	wire [4-1:0] node1859;
	wire [4-1:0] node1861;
	wire [4-1:0] node1863;
	wire [4-1:0] node1866;
	wire [4-1:0] node1867;
	wire [4-1:0] node1868;
	wire [4-1:0] node1869;
	wire [4-1:0] node1873;
	wire [4-1:0] node1876;
	wire [4-1:0] node1878;
	wire [4-1:0] node1879;
	wire [4-1:0] node1880;
	wire [4-1:0] node1884;
	wire [4-1:0] node1887;
	wire [4-1:0] node1888;
	wire [4-1:0] node1889;
	wire [4-1:0] node1890;
	wire [4-1:0] node1894;
	wire [4-1:0] node1895;
	wire [4-1:0] node1897;
	wire [4-1:0] node1898;
	wire [4-1:0] node1901;
	wire [4-1:0] node1904;
	wire [4-1:0] node1905;
	wire [4-1:0] node1906;
	wire [4-1:0] node1907;
	wire [4-1:0] node1913;
	wire [4-1:0] node1914;
	wire [4-1:0] node1915;
	wire [4-1:0] node1916;
	wire [4-1:0] node1919;
	wire [4-1:0] node1920;
	wire [4-1:0] node1924;
	wire [4-1:0] node1925;
	wire [4-1:0] node1926;
	wire [4-1:0] node1929;
	wire [4-1:0] node1933;
	wire [4-1:0] node1934;
	wire [4-1:0] node1938;
	wire [4-1:0] node1939;
	wire [4-1:0] node1940;
	wire [4-1:0] node1941;
	wire [4-1:0] node1943;
	wire [4-1:0] node1944;
	wire [4-1:0] node1945;
	wire [4-1:0] node1949;
	wire [4-1:0] node1952;
	wire [4-1:0] node1953;
	wire [4-1:0] node1954;
	wire [4-1:0] node1957;
	wire [4-1:0] node1961;
	wire [4-1:0] node1962;
	wire [4-1:0] node1963;
	wire [4-1:0] node1964;
	wire [4-1:0] node1967;
	wire [4-1:0] node1970;
	wire [4-1:0] node1972;
	wire [4-1:0] node1975;
	wire [4-1:0] node1977;
	wire [4-1:0] node1978;
	wire [4-1:0] node1982;
	wire [4-1:0] node1983;
	wire [4-1:0] node1984;
	wire [4-1:0] node1985;
	wire [4-1:0] node1986;
	wire [4-1:0] node1990;
	wire [4-1:0] node1991;
	wire [4-1:0] node1996;
	wire [4-1:0] node1997;
	wire [4-1:0] node1999;
	wire [4-1:0] node2000;
	wire [4-1:0] node2003;
	wire [4-1:0] node2007;
	wire [4-1:0] node2008;
	wire [4-1:0] node2009;
	wire [4-1:0] node2010;
	wire [4-1:0] node2011;
	wire [4-1:0] node2012;
	wire [4-1:0] node2013;
	wire [4-1:0] node2017;
	wire [4-1:0] node2020;
	wire [4-1:0] node2021;
	wire [4-1:0] node2023;
	wire [4-1:0] node2025;
	wire [4-1:0] node2028;
	wire [4-1:0] node2031;
	wire [4-1:0] node2032;
	wire [4-1:0] node2033;
	wire [4-1:0] node2034;
	wire [4-1:0] node2038;
	wire [4-1:0] node2040;
	wire [4-1:0] node2043;
	wire [4-1:0] node2045;
	wire [4-1:0] node2048;
	wire [4-1:0] node2049;
	wire [4-1:0] node2050;
	wire [4-1:0] node2052;
	wire [4-1:0] node2054;
	wire [4-1:0] node2057;
	wire [4-1:0] node2058;
	wire [4-1:0] node2061;
	wire [4-1:0] node2064;
	wire [4-1:0] node2065;
	wire [4-1:0] node2066;
	wire [4-1:0] node2070;
	wire [4-1:0] node2071;
	wire [4-1:0] node2072;
	wire [4-1:0] node2076;
	wire [4-1:0] node2077;
	wire [4-1:0] node2081;
	wire [4-1:0] node2082;
	wire [4-1:0] node2083;
	wire [4-1:0] node2084;
	wire [4-1:0] node2085;
	wire [4-1:0] node2086;
	wire [4-1:0] node2087;
	wire [4-1:0] node2089;
	wire [4-1:0] node2094;
	wire [4-1:0] node2095;
	wire [4-1:0] node2099;
	wire [4-1:0] node2100;
	wire [4-1:0] node2104;
	wire [4-1:0] node2105;
	wire [4-1:0] node2106;
	wire [4-1:0] node2109;
	wire [4-1:0] node2111;
	wire [4-1:0] node2114;
	wire [4-1:0] node2115;
	wire [4-1:0] node2120;
	wire [4-1:0] node2121;
	wire [4-1:0] node2122;
	wire [4-1:0] node2123;
	wire [4-1:0] node2124;
	wire [4-1:0] node2125;
	wire [4-1:0] node2126;
	wire [4-1:0] node2127;
	wire [4-1:0] node2130;
	wire [4-1:0] node2131;
	wire [4-1:0] node2133;
	wire [4-1:0] node2137;
	wire [4-1:0] node2138;
	wire [4-1:0] node2139;
	wire [4-1:0] node2141;
	wire [4-1:0] node2144;
	wire [4-1:0] node2146;
	wire [4-1:0] node2149;
	wire [4-1:0] node2151;
	wire [4-1:0] node2154;
	wire [4-1:0] node2155;
	wire [4-1:0] node2157;
	wire [4-1:0] node2159;
	wire [4-1:0] node2162;
	wire [4-1:0] node2165;
	wire [4-1:0] node2166;
	wire [4-1:0] node2167;
	wire [4-1:0] node2170;
	wire [4-1:0] node2171;
	wire [4-1:0] node2173;
	wire [4-1:0] node2176;
	wire [4-1:0] node2178;
	wire [4-1:0] node2181;
	wire [4-1:0] node2182;
	wire [4-1:0] node2183;
	wire [4-1:0] node2184;
	wire [4-1:0] node2187;
	wire [4-1:0] node2190;
	wire [4-1:0] node2192;
	wire [4-1:0] node2194;
	wire [4-1:0] node2197;
	wire [4-1:0] node2198;
	wire [4-1:0] node2202;
	wire [4-1:0] node2203;
	wire [4-1:0] node2204;
	wire [4-1:0] node2205;
	wire [4-1:0] node2206;
	wire [4-1:0] node2207;
	wire [4-1:0] node2211;
	wire [4-1:0] node2212;
	wire [4-1:0] node2213;
	wire [4-1:0] node2218;
	wire [4-1:0] node2220;
	wire [4-1:0] node2221;
	wire [4-1:0] node2225;
	wire [4-1:0] node2226;
	wire [4-1:0] node2227;
	wire [4-1:0] node2228;
	wire [4-1:0] node2230;
	wire [4-1:0] node2233;
	wire [4-1:0] node2234;
	wire [4-1:0] node2238;
	wire [4-1:0] node2239;
	wire [4-1:0] node2243;
	wire [4-1:0] node2246;
	wire [4-1:0] node2247;
	wire [4-1:0] node2248;
	wire [4-1:0] node2250;
	wire [4-1:0] node2251;
	wire [4-1:0] node2252;
	wire [4-1:0] node2255;
	wire [4-1:0] node2256;
	wire [4-1:0] node2260;
	wire [4-1:0] node2263;
	wire [4-1:0] node2264;
	wire [4-1:0] node2265;
	wire [4-1:0] node2267;
	wire [4-1:0] node2270;
	wire [4-1:0] node2273;
	wire [4-1:0] node2275;
	wire [4-1:0] node2276;
	wire [4-1:0] node2280;
	wire [4-1:0] node2281;
	wire [4-1:0] node2283;
	wire [4-1:0] node2284;
	wire [4-1:0] node2287;
	wire [4-1:0] node2290;
	wire [4-1:0] node2291;
	wire [4-1:0] node2292;
	wire [4-1:0] node2297;
	wire [4-1:0] node2298;
	wire [4-1:0] node2299;
	wire [4-1:0] node2300;
	wire [4-1:0] node2301;
	wire [4-1:0] node2302;
	wire [4-1:0] node2304;
	wire [4-1:0] node2307;
	wire [4-1:0] node2309;
	wire [4-1:0] node2310;
	wire [4-1:0] node2312;
	wire [4-1:0] node2315;
	wire [4-1:0] node2318;
	wire [4-1:0] node2319;
	wire [4-1:0] node2322;
	wire [4-1:0] node2324;
	wire [4-1:0] node2326;
	wire [4-1:0] node2329;
	wire [4-1:0] node2330;
	wire [4-1:0] node2331;
	wire [4-1:0] node2332;
	wire [4-1:0] node2336;
	wire [4-1:0] node2337;
	wire [4-1:0] node2342;
	wire [4-1:0] node2343;
	wire [4-1:0] node2344;
	wire [4-1:0] node2345;
	wire [4-1:0] node2346;
	wire [4-1:0] node2349;
	wire [4-1:0] node2353;
	wire [4-1:0] node2355;
	wire [4-1:0] node2358;
	wire [4-1:0] node2359;
	wire [4-1:0] node2360;
	wire [4-1:0] node2362;
	wire [4-1:0] node2365;
	wire [4-1:0] node2368;
	wire [4-1:0] node2369;
	wire [4-1:0] node2370;
	wire [4-1:0] node2371;
	wire [4-1:0] node2375;
	wire [4-1:0] node2377;
	wire [4-1:0] node2380;
	wire [4-1:0] node2381;
	wire [4-1:0] node2382;
	wire [4-1:0] node2383;
	wire [4-1:0] node2389;
	wire [4-1:0] node2390;
	wire [4-1:0] node2391;
	wire [4-1:0] node2392;
	wire [4-1:0] node2395;
	wire [4-1:0] node2396;
	wire [4-1:0] node2398;
	wire [4-1:0] node2402;
	wire [4-1:0] node2403;
	wire [4-1:0] node2404;
	wire [4-1:0] node2408;
	wire [4-1:0] node2409;
	wire [4-1:0] node2410;
	wire [4-1:0] node2414;
	wire [4-1:0] node2417;
	wire [4-1:0] node2418;
	wire [4-1:0] node2419;
	wire [4-1:0] node2420;
	wire [4-1:0] node2421;
	wire [4-1:0] node2422;
	wire [4-1:0] node2428;
	wire [4-1:0] node2429;
	wire [4-1:0] node2430;
	wire [4-1:0] node2434;
	wire [4-1:0] node2435;
	wire [4-1:0] node2440;
	wire [4-1:0] node2441;
	wire [4-1:0] node2442;
	wire [4-1:0] node2443;
	wire [4-1:0] node2444;
	wire [4-1:0] node2445;
	wire [4-1:0] node2446;
	wire [4-1:0] node2448;
	wire [4-1:0] node2449;
	wire [4-1:0] node2453;
	wire [4-1:0] node2454;
	wire [4-1:0] node2457;
	wire [4-1:0] node2459;
	wire [4-1:0] node2462;
	wire [4-1:0] node2463;
	wire [4-1:0] node2465;
	wire [4-1:0] node2468;
	wire [4-1:0] node2469;
	wire [4-1:0] node2471;
	wire [4-1:0] node2474;
	wire [4-1:0] node2475;
	wire [4-1:0] node2479;
	wire [4-1:0] node2480;
	wire [4-1:0] node2482;
	wire [4-1:0] node2483;
	wire [4-1:0] node2485;
	wire [4-1:0] node2489;
	wire [4-1:0] node2490;
	wire [4-1:0] node2491;
	wire [4-1:0] node2494;
	wire [4-1:0] node2498;
	wire [4-1:0] node2499;
	wire [4-1:0] node2500;
	wire [4-1:0] node2501;
	wire [4-1:0] node2503;
	wire [4-1:0] node2506;
	wire [4-1:0] node2509;
	wire [4-1:0] node2510;
	wire [4-1:0] node2512;
	wire [4-1:0] node2513;
	wire [4-1:0] node2518;
	wire [4-1:0] node2519;
	wire [4-1:0] node2520;
	wire [4-1:0] node2523;
	wire [4-1:0] node2526;
	wire [4-1:0] node2527;
	wire [4-1:0] node2528;
	wire [4-1:0] node2530;
	wire [4-1:0] node2533;
	wire [4-1:0] node2536;
	wire [4-1:0] node2537;
	wire [4-1:0] node2541;
	wire [4-1:0] node2542;
	wire [4-1:0] node2543;
	wire [4-1:0] node2544;
	wire [4-1:0] node2545;
	wire [4-1:0] node2547;
	wire [4-1:0] node2549;
	wire [4-1:0] node2553;
	wire [4-1:0] node2554;
	wire [4-1:0] node2555;
	wire [4-1:0] node2556;
	wire [4-1:0] node2562;
	wire [4-1:0] node2563;
	wire [4-1:0] node2565;
	wire [4-1:0] node2568;
	wire [4-1:0] node2569;
	wire [4-1:0] node2570;
	wire [4-1:0] node2571;
	wire [4-1:0] node2572;
	wire [4-1:0] node2578;
	wire [4-1:0] node2581;
	wire [4-1:0] node2582;
	wire [4-1:0] node2583;
	wire [4-1:0] node2584;
	wire [4-1:0] node2585;
	wire [4-1:0] node2590;
	wire [4-1:0] node2591;
	wire [4-1:0] node2596;
	wire [4-1:0] node2597;
	wire [4-1:0] node2598;
	wire [4-1:0] node2599;
	wire [4-1:0] node2600;
	wire [4-1:0] node2602;
	wire [4-1:0] node2605;
	wire [4-1:0] node2607;
	wire [4-1:0] node2610;
	wire [4-1:0] node2612;
	wire [4-1:0] node2615;
	wire [4-1:0] node2616;
	wire [4-1:0] node2617;
	wire [4-1:0] node2618;
	wire [4-1:0] node2620;
	wire [4-1:0] node2623;
	wire [4-1:0] node2625;
	wire [4-1:0] node2628;
	wire [4-1:0] node2629;
	wire [4-1:0] node2631;
	wire [4-1:0] node2636;
	wire [4-1:0] node2638;
	wire [4-1:0] node2639;
	wire [4-1:0] node2641;
	wire [4-1:0] node2645;
	wire [4-1:0] node2646;
	wire [4-1:0] node2647;
	wire [4-1:0] node2648;
	wire [4-1:0] node2649;
	wire [4-1:0] node2650;
	wire [4-1:0] node2651;
	wire [4-1:0] node2652;
	wire [4-1:0] node2653;
	wire [4-1:0] node2655;
	wire [4-1:0] node2656;
	wire [4-1:0] node2657;
	wire [4-1:0] node2663;
	wire [4-1:0] node2664;
	wire [4-1:0] node2665;
	wire [4-1:0] node2666;
	wire [4-1:0] node2668;
	wire [4-1:0] node2671;
	wire [4-1:0] node2673;
	wire [4-1:0] node2675;
	wire [4-1:0] node2678;
	wire [4-1:0] node2679;
	wire [4-1:0] node2681;
	wire [4-1:0] node2684;
	wire [4-1:0] node2686;
	wire [4-1:0] node2689;
	wire [4-1:0] node2691;
	wire [4-1:0] node2692;
	wire [4-1:0] node2693;
	wire [4-1:0] node2697;
	wire [4-1:0] node2698;
	wire [4-1:0] node2699;
	wire [4-1:0] node2702;
	wire [4-1:0] node2706;
	wire [4-1:0] node2707;
	wire [4-1:0] node2708;
	wire [4-1:0] node2709;
	wire [4-1:0] node2711;
	wire [4-1:0] node2713;
	wire [4-1:0] node2716;
	wire [4-1:0] node2718;
	wire [4-1:0] node2721;
	wire [4-1:0] node2722;
	wire [4-1:0] node2724;
	wire [4-1:0] node2727;
	wire [4-1:0] node2728;
	wire [4-1:0] node2731;
	wire [4-1:0] node2732;
	wire [4-1:0] node2734;
	wire [4-1:0] node2737;
	wire [4-1:0] node2740;
	wire [4-1:0] node2741;
	wire [4-1:0] node2742;
	wire [4-1:0] node2744;
	wire [4-1:0] node2747;
	wire [4-1:0] node2749;
	wire [4-1:0] node2752;
	wire [4-1:0] node2753;
	wire [4-1:0] node2754;
	wire [4-1:0] node2755;
	wire [4-1:0] node2759;
	wire [4-1:0] node2760;
	wire [4-1:0] node2761;
	wire [4-1:0] node2766;
	wire [4-1:0] node2767;
	wire [4-1:0] node2769;
	wire [4-1:0] node2772;
	wire [4-1:0] node2774;
	wire [4-1:0] node2775;
	wire [4-1:0] node2780;
	wire [4-1:0] node2781;
	wire [4-1:0] node2782;
	wire [4-1:0] node2783;
	wire [4-1:0] node2784;
	wire [4-1:0] node2785;
	wire [4-1:0] node2786;
	wire [4-1:0] node2788;
	wire [4-1:0] node2791;
	wire [4-1:0] node2792;
	wire [4-1:0] node2796;
	wire [4-1:0] node2797;
	wire [4-1:0] node2798;
	wire [4-1:0] node2801;
	wire [4-1:0] node2804;
	wire [4-1:0] node2807;
	wire [4-1:0] node2808;
	wire [4-1:0] node2810;
	wire [4-1:0] node2813;
	wire [4-1:0] node2814;
	wire [4-1:0] node2818;
	wire [4-1:0] node2819;
	wire [4-1:0] node2821;
	wire [4-1:0] node2823;
	wire [4-1:0] node2825;
	wire [4-1:0] node2828;
	wire [4-1:0] node2829;
	wire [4-1:0] node2830;
	wire [4-1:0] node2832;
	wire [4-1:0] node2834;
	wire [4-1:0] node2837;
	wire [4-1:0] node2840;
	wire [4-1:0] node2842;
	wire [4-1:0] node2845;
	wire [4-1:0] node2846;
	wire [4-1:0] node2847;
	wire [4-1:0] node2849;
	wire [4-1:0] node2850;
	wire [4-1:0] node2851;
	wire [4-1:0] node2856;
	wire [4-1:0] node2857;
	wire [4-1:0] node2858;
	wire [4-1:0] node2862;
	wire [4-1:0] node2863;
	wire [4-1:0] node2865;
	wire [4-1:0] node2869;
	wire [4-1:0] node2870;
	wire [4-1:0] node2871;
	wire [4-1:0] node2872;
	wire [4-1:0] node2873;
	wire [4-1:0] node2878;
	wire [4-1:0] node2879;
	wire [4-1:0] node2883;
	wire [4-1:0] node2884;
	wire [4-1:0] node2885;
	wire [4-1:0] node2887;
	wire [4-1:0] node2891;
	wire [4-1:0] node2893;
	wire [4-1:0] node2896;
	wire [4-1:0] node2897;
	wire [4-1:0] node2898;
	wire [4-1:0] node2899;
	wire [4-1:0] node2900;
	wire [4-1:0] node2901;
	wire [4-1:0] node2904;
	wire [4-1:0] node2907;
	wire [4-1:0] node2908;
	wire [4-1:0] node2909;
	wire [4-1:0] node2913;
	wire [4-1:0] node2916;
	wire [4-1:0] node2918;
	wire [4-1:0] node2919;
	wire [4-1:0] node2923;
	wire [4-1:0] node2924;
	wire [4-1:0] node2925;
	wire [4-1:0] node2927;
	wire [4-1:0] node2930;
	wire [4-1:0] node2932;
	wire [4-1:0] node2935;
	wire [4-1:0] node2936;
	wire [4-1:0] node2937;
	wire [4-1:0] node2939;
	wire [4-1:0] node2942;
	wire [4-1:0] node2945;
	wire [4-1:0] node2946;
	wire [4-1:0] node2947;
	wire [4-1:0] node2951;
	wire [4-1:0] node2954;
	wire [4-1:0] node2955;
	wire [4-1:0] node2956;
	wire [4-1:0] node2957;
	wire [4-1:0] node2959;
	wire [4-1:0] node2962;
	wire [4-1:0] node2964;
	wire [4-1:0] node2967;
	wire [4-1:0] node2968;
	wire [4-1:0] node2969;
	wire [4-1:0] node2973;
	wire [4-1:0] node2974;
	wire [4-1:0] node2978;
	wire [4-1:0] node2979;
	wire [4-1:0] node2980;
	wire [4-1:0] node2981;
	wire [4-1:0] node2984;
	wire [4-1:0] node2986;
	wire [4-1:0] node2989;
	wire [4-1:0] node2990;
	wire [4-1:0] node2993;
	wire [4-1:0] node2995;
	wire [4-1:0] node2998;
	wire [4-1:0] node2999;
	wire [4-1:0] node3000;
	wire [4-1:0] node3001;
	wire [4-1:0] node3003;
	wire [4-1:0] node3004;
	wire [4-1:0] node3007;
	wire [4-1:0] node3011;
	wire [4-1:0] node3014;
	wire [4-1:0] node3015;
	wire [4-1:0] node3018;
	wire [4-1:0] node3022;
	wire [4-1:0] node3023;
	wire [4-1:0] node3024;
	wire [4-1:0] node3025;
	wire [4-1:0] node3026;
	wire [4-1:0] node3027;
	wire [4-1:0] node3028;
	wire [4-1:0] node3029;
	wire [4-1:0] node3030;
	wire [4-1:0] node3032;
	wire [4-1:0] node3035;
	wire [4-1:0] node3038;
	wire [4-1:0] node3039;
	wire [4-1:0] node3040;
	wire [4-1:0] node3042;
	wire [4-1:0] node3043;
	wire [4-1:0] node3049;
	wire [4-1:0] node3050;
	wire [4-1:0] node3051;
	wire [4-1:0] node3054;
	wire [4-1:0] node3056;
	wire [4-1:0] node3058;
	wire [4-1:0] node3061;
	wire [4-1:0] node3062;
	wire [4-1:0] node3064;
	wire [4-1:0] node3067;
	wire [4-1:0] node3070;
	wire [4-1:0] node3071;
	wire [4-1:0] node3072;
	wire [4-1:0] node3075;
	wire [4-1:0] node3076;
	wire [4-1:0] node3077;
	wire [4-1:0] node3081;
	wire [4-1:0] node3082;
	wire [4-1:0] node3084;
	wire [4-1:0] node3088;
	wire [4-1:0] node3089;
	wire [4-1:0] node3090;
	wire [4-1:0] node3092;
	wire [4-1:0] node3095;
	wire [4-1:0] node3098;
	wire [4-1:0] node3099;
	wire [4-1:0] node3100;
	wire [4-1:0] node3102;
	wire [4-1:0] node3107;
	wire [4-1:0] node3108;
	wire [4-1:0] node3109;
	wire [4-1:0] node3110;
	wire [4-1:0] node3111;
	wire [4-1:0] node3113;
	wire [4-1:0] node3116;
	wire [4-1:0] node3119;
	wire [4-1:0] node3120;
	wire [4-1:0] node3121;
	wire [4-1:0] node3124;
	wire [4-1:0] node3127;
	wire [4-1:0] node3128;
	wire [4-1:0] node3129;
	wire [4-1:0] node3132;
	wire [4-1:0] node3135;
	wire [4-1:0] node3138;
	wire [4-1:0] node3139;
	wire [4-1:0] node3140;
	wire [4-1:0] node3142;
	wire [4-1:0] node3145;
	wire [4-1:0] node3147;
	wire [4-1:0] node3150;
	wire [4-1:0] node3151;
	wire [4-1:0] node3154;
	wire [4-1:0] node3155;
	wire [4-1:0] node3159;
	wire [4-1:0] node3160;
	wire [4-1:0] node3161;
	wire [4-1:0] node3163;
	wire [4-1:0] node3164;
	wire [4-1:0] node3168;
	wire [4-1:0] node3170;
	wire [4-1:0] node3172;
	wire [4-1:0] node3173;
	wire [4-1:0] node3177;
	wire [4-1:0] node3178;
	wire [4-1:0] node3179;
	wire [4-1:0] node3182;
	wire [4-1:0] node3183;
	wire [4-1:0] node3186;
	wire [4-1:0] node3189;
	wire [4-1:0] node3190;
	wire [4-1:0] node3194;
	wire [4-1:0] node3195;
	wire [4-1:0] node3196;
	wire [4-1:0] node3197;
	wire [4-1:0] node3198;
	wire [4-1:0] node3200;
	wire [4-1:0] node3203;
	wire [4-1:0] node3204;
	wire [4-1:0] node3205;
	wire [4-1:0] node3206;
	wire [4-1:0] node3209;
	wire [4-1:0] node3213;
	wire [4-1:0] node3216;
	wire [4-1:0] node3217;
	wire [4-1:0] node3220;
	wire [4-1:0] node3221;
	wire [4-1:0] node3224;
	wire [4-1:0] node3227;
	wire [4-1:0] node3228;
	wire [4-1:0] node3229;
	wire [4-1:0] node3231;
	wire [4-1:0] node3233;
	wire [4-1:0] node3236;
	wire [4-1:0] node3237;
	wire [4-1:0] node3239;
	wire [4-1:0] node3240;
	wire [4-1:0] node3245;
	wire [4-1:0] node3246;
	wire [4-1:0] node3247;
	wire [4-1:0] node3248;
	wire [4-1:0] node3252;
	wire [4-1:0] node3254;
	wire [4-1:0] node3257;
	wire [4-1:0] node3259;
	wire [4-1:0] node3261;
	wire [4-1:0] node3264;
	wire [4-1:0] node3265;
	wire [4-1:0] node3266;
	wire [4-1:0] node3267;
	wire [4-1:0] node3268;
	wire [4-1:0] node3270;
	wire [4-1:0] node3273;
	wire [4-1:0] node3276;
	wire [4-1:0] node3278;
	wire [4-1:0] node3279;
	wire [4-1:0] node3283;
	wire [4-1:0] node3284;
	wire [4-1:0] node3285;
	wire [4-1:0] node3289;
	wire [4-1:0] node3290;
	wire [4-1:0] node3291;
	wire [4-1:0] node3292;
	wire [4-1:0] node3298;
	wire [4-1:0] node3299;
	wire [4-1:0] node3300;
	wire [4-1:0] node3302;
	wire [4-1:0] node3305;
	wire [4-1:0] node3306;
	wire [4-1:0] node3309;
	wire [4-1:0] node3312;
	wire [4-1:0] node3313;
	wire [4-1:0] node3314;
	wire [4-1:0] node3318;
	wire [4-1:0] node3319;
	wire [4-1:0] node3323;
	wire [4-1:0] node3324;
	wire [4-1:0] node3325;
	wire [4-1:0] node3326;
	wire [4-1:0] node3328;
	wire [4-1:0] node3329;
	wire [4-1:0] node3330;
	wire [4-1:0] node3331;
	wire [4-1:0] node3337;
	wire [4-1:0] node3338;
	wire [4-1:0] node3339;
	wire [4-1:0] node3342;
	wire [4-1:0] node3343;
	wire [4-1:0] node3344;
	wire [4-1:0] node3348;
	wire [4-1:0] node3349;
	wire [4-1:0] node3353;
	wire [4-1:0] node3355;
	wire [4-1:0] node3358;
	wire [4-1:0] node3359;
	wire [4-1:0] node3360;
	wire [4-1:0] node3361;
	wire [4-1:0] node3363;
	wire [4-1:0] node3366;
	wire [4-1:0] node3367;
	wire [4-1:0] node3368;
	wire [4-1:0] node3372;
	wire [4-1:0] node3374;
	wire [4-1:0] node3377;
	wire [4-1:0] node3378;
	wire [4-1:0] node3379;
	wire [4-1:0] node3381;
	wire [4-1:0] node3384;
	wire [4-1:0] node3385;
	wire [4-1:0] node3389;
	wire [4-1:0] node3390;
	wire [4-1:0] node3392;
	wire [4-1:0] node3396;
	wire [4-1:0] node3397;
	wire [4-1:0] node3398;
	wire [4-1:0] node3399;
	wire [4-1:0] node3402;
	wire [4-1:0] node3403;
	wire [4-1:0] node3407;
	wire [4-1:0] node3408;
	wire [4-1:0] node3409;
	wire [4-1:0] node3410;
	wire [4-1:0] node3414;
	wire [4-1:0] node3417;
	wire [4-1:0] node3418;
	wire [4-1:0] node3422;
	wire [4-1:0] node3423;
	wire [4-1:0] node3424;
	wire [4-1:0] node3428;
	wire [4-1:0] node3429;
	wire [4-1:0] node3432;
	wire [4-1:0] node3434;
	wire [4-1:0] node3438;
	wire [4-1:0] node3439;
	wire [4-1:0] node3440;
	wire [4-1:0] node3441;
	wire [4-1:0] node3442;
	wire [4-1:0] node3443;
	wire [4-1:0] node3444;
	wire [4-1:0] node3445;
	wire [4-1:0] node3447;
	wire [4-1:0] node3450;
	wire [4-1:0] node3452;
	wire [4-1:0] node3455;
	wire [4-1:0] node3456;
	wire [4-1:0] node3457;
	wire [4-1:0] node3459;
	wire [4-1:0] node3462;
	wire [4-1:0] node3465;
	wire [4-1:0] node3467;
	wire [4-1:0] node3468;
	wire [4-1:0] node3472;
	wire [4-1:0] node3473;
	wire [4-1:0] node3474;
	wire [4-1:0] node3476;
	wire [4-1:0] node3479;
	wire [4-1:0] node3480;
	wire [4-1:0] node3484;
	wire [4-1:0] node3485;
	wire [4-1:0] node3486;
	wire [4-1:0] node3487;
	wire [4-1:0] node3492;
	wire [4-1:0] node3495;
	wire [4-1:0] node3496;
	wire [4-1:0] node3497;
	wire [4-1:0] node3498;
	wire [4-1:0] node3500;
	wire [4-1:0] node3502;
	wire [4-1:0] node3505;
	wire [4-1:0] node3506;
	wire [4-1:0] node3510;
	wire [4-1:0] node3512;
	wire [4-1:0] node3515;
	wire [4-1:0] node3516;
	wire [4-1:0] node3517;
	wire [4-1:0] node3518;
	wire [4-1:0] node3520;
	wire [4-1:0] node3523;
	wire [4-1:0] node3524;
	wire [4-1:0] node3527;
	wire [4-1:0] node3530;
	wire [4-1:0] node3533;
	wire [4-1:0] node3534;
	wire [4-1:0] node3537;
	wire [4-1:0] node3538;
	wire [4-1:0] node3542;
	wire [4-1:0] node3543;
	wire [4-1:0] node3544;
	wire [4-1:0] node3545;
	wire [4-1:0] node3546;
	wire [4-1:0] node3547;
	wire [4-1:0] node3548;
	wire [4-1:0] node3549;
	wire [4-1:0] node3555;
	wire [4-1:0] node3556;
	wire [4-1:0] node3558;
	wire [4-1:0] node3562;
	wire [4-1:0] node3565;
	wire [4-1:0] node3566;
	wire [4-1:0] node3569;
	wire [4-1:0] node3571;
	wire [4-1:0] node3573;
	wire [4-1:0] node3576;
	wire [4-1:0] node3577;
	wire [4-1:0] node3579;
	wire [4-1:0] node3580;
	wire [4-1:0] node3581;
	wire [4-1:0] node3585;
	wire [4-1:0] node3587;
	wire [4-1:0] node3588;
	wire [4-1:0] node3593;
	wire [4-1:0] node3594;
	wire [4-1:0] node3595;
	wire [4-1:0] node3596;
	wire [4-1:0] node3597;
	wire [4-1:0] node3599;
	wire [4-1:0] node3601;
	wire [4-1:0] node3604;
	wire [4-1:0] node3605;
	wire [4-1:0] node3609;
	wire [4-1:0] node3610;
	wire [4-1:0] node3611;
	wire [4-1:0] node3612;
	wire [4-1:0] node3616;
	wire [4-1:0] node3619;
	wire [4-1:0] node3620;
	wire [4-1:0] node3621;
	wire [4-1:0] node3624;
	wire [4-1:0] node3626;
	wire [4-1:0] node3629;
	wire [4-1:0] node3630;
	wire [4-1:0] node3634;
	wire [4-1:0] node3635;
	wire [4-1:0] node3636;
	wire [4-1:0] node3637;
	wire [4-1:0] node3639;
	wire [4-1:0] node3641;
	wire [4-1:0] node3644;
	wire [4-1:0] node3645;
	wire [4-1:0] node3649;
	wire [4-1:0] node3650;
	wire [4-1:0] node3651;
	wire [4-1:0] node3652;
	wire [4-1:0] node3655;
	wire [4-1:0] node3658;
	wire [4-1:0] node3660;
	wire [4-1:0] node3663;
	wire [4-1:0] node3664;
	wire [4-1:0] node3668;
	wire [4-1:0] node3669;
	wire [4-1:0] node3670;
	wire [4-1:0] node3671;
	wire [4-1:0] node3673;
	wire [4-1:0] node3674;
	wire [4-1:0] node3678;
	wire [4-1:0] node3681;
	wire [4-1:0] node3683;
	wire [4-1:0] node3686;
	wire [4-1:0] node3687;
	wire [4-1:0] node3689;
	wire [4-1:0] node3690;
	wire [4-1:0] node3695;
	wire [4-1:0] node3696;
	wire [4-1:0] node3697;
	wire [4-1:0] node3698;
	wire [4-1:0] node3699;
	wire [4-1:0] node3700;
	wire [4-1:0] node3704;
	wire [4-1:0] node3706;
	wire [4-1:0] node3709;
	wire [4-1:0] node3710;
	wire [4-1:0] node3713;
	wire [4-1:0] node3714;
	wire [4-1:0] node3716;
	wire [4-1:0] node3720;
	wire [4-1:0] node3721;
	wire [4-1:0] node3722;
	wire [4-1:0] node3724;
	wire [4-1:0] node3725;
	wire [4-1:0] node3729;
	wire [4-1:0] node3730;
	wire [4-1:0] node3734;
	wire [4-1:0] node3735;
	wire [4-1:0] node3738;
	wire [4-1:0] node3741;
	wire [4-1:0] node3742;
	wire [4-1:0] node3743;
	wire [4-1:0] node3745;
	wire [4-1:0] node3748;
	wire [4-1:0] node3749;
	wire [4-1:0] node3750;
	wire [4-1:0] node3754;
	wire [4-1:0] node3755;
	wire [4-1:0] node3759;
	wire [4-1:0] node3762;
	wire [4-1:0] node3763;
	wire [4-1:0] node3764;
	wire [4-1:0] node3765;
	wire [4-1:0] node3766;
	wire [4-1:0] node3767;
	wire [4-1:0] node3768;
	wire [4-1:0] node3769;
	wire [4-1:0] node3773;
	wire [4-1:0] node3774;
	wire [4-1:0] node3777;
	wire [4-1:0] node3780;
	wire [4-1:0] node3781;
	wire [4-1:0] node3783;
	wire [4-1:0] node3786;
	wire [4-1:0] node3787;
	wire [4-1:0] node3788;
	wire [4-1:0] node3793;
	wire [4-1:0] node3794;
	wire [4-1:0] node3795;
	wire [4-1:0] node3796;
	wire [4-1:0] node3800;
	wire [4-1:0] node3803;
	wire [4-1:0] node3805;
	wire [4-1:0] node3807;
	wire [4-1:0] node3810;
	wire [4-1:0] node3811;
	wire [4-1:0] node3812;
	wire [4-1:0] node3813;
	wire [4-1:0] node3815;
	wire [4-1:0] node3819;
	wire [4-1:0] node3820;
	wire [4-1:0] node3821;
	wire [4-1:0] node3822;
	wire [4-1:0] node3826;
	wire [4-1:0] node3827;
	wire [4-1:0] node3831;
	wire [4-1:0] node3833;
	wire [4-1:0] node3836;
	wire [4-1:0] node3837;
	wire [4-1:0] node3838;
	wire [4-1:0] node3839;
	wire [4-1:0] node3843;
	wire [4-1:0] node3844;
	wire [4-1:0] node3848;
	wire [4-1:0] node3850;
	wire [4-1:0] node3851;
	wire [4-1:0] node3854;
	wire [4-1:0] node3856;
	wire [4-1:0] node3859;
	wire [4-1:0] node3860;
	wire [4-1:0] node3861;
	wire [4-1:0] node3862;
	wire [4-1:0] node3864;
	wire [4-1:0] node3866;
	wire [4-1:0] node3869;
	wire [4-1:0] node3870;
	wire [4-1:0] node3872;
	wire [4-1:0] node3875;
	wire [4-1:0] node3877;
	wire [4-1:0] node3880;
	wire [4-1:0] node3881;
	wire [4-1:0] node3882;
	wire [4-1:0] node3884;
	wire [4-1:0] node3887;
	wire [4-1:0] node3889;
	wire [4-1:0] node3892;
	wire [4-1:0] node3895;
	wire [4-1:0] node3896;
	wire [4-1:0] node3897;
	wire [4-1:0] node3899;
	wire [4-1:0] node3902;
	wire [4-1:0] node3903;
	wire [4-1:0] node3907;
	wire [4-1:0] node3908;
	wire [4-1:0] node3910;
	wire [4-1:0] node3913;
	wire [4-1:0] node3915;
	wire [4-1:0] node3916;
	wire [4-1:0] node3918;
	wire [4-1:0] node3922;
	wire [4-1:0] node3923;
	wire [4-1:0] node3924;
	wire [4-1:0] node3925;
	wire [4-1:0] node3926;
	wire [4-1:0] node3927;
	wire [4-1:0] node3928;
	wire [4-1:0] node3932;
	wire [4-1:0] node3933;
	wire [4-1:0] node3934;
	wire [4-1:0] node3938;
	wire [4-1:0] node3940;
	wire [4-1:0] node3943;
	wire [4-1:0] node3944;
	wire [4-1:0] node3945;
	wire [4-1:0] node3950;
	wire [4-1:0] node3951;
	wire [4-1:0] node3952;
	wire [4-1:0] node3953;
	wire [4-1:0] node3957;
	wire [4-1:0] node3959;
	wire [4-1:0] node3962;
	wire [4-1:0] node3963;
	wire [4-1:0] node3964;
	wire [4-1:0] node3967;
	wire [4-1:0] node3970;
	wire [4-1:0] node3971;
	wire [4-1:0] node3974;
	wire [4-1:0] node3975;
	wire [4-1:0] node3979;
	wire [4-1:0] node3980;
	wire [4-1:0] node3981;
	wire [4-1:0] node3982;
	wire [4-1:0] node3984;
	wire [4-1:0] node3985;
	wire [4-1:0] node3990;
	wire [4-1:0] node3991;
	wire [4-1:0] node3994;
	wire [4-1:0] node3995;
	wire [4-1:0] node4000;
	wire [4-1:0] node4001;
	wire [4-1:0] node4002;
	wire [4-1:0] node4003;
	wire [4-1:0] node4004;
	wire [4-1:0] node4006;
	wire [4-1:0] node4008;
	wire [4-1:0] node4010;
	wire [4-1:0] node4014;
	wire [4-1:0] node4015;
	wire [4-1:0] node4016;
	wire [4-1:0] node4017;
	wire [4-1:0] node4022;
	wire [4-1:0] node4024;
	wire [4-1:0] node4027;
	wire [4-1:0] node4028;
	wire [4-1:0] node4030;
	wire [4-1:0] node4032;
	wire [4-1:0] node4034;
	wire [4-1:0] node4038;
	wire [4-1:0] node4040;
	wire [4-1:0] node4041;
	wire [4-1:0] node4042;
	wire [4-1:0] node4043;
	wire [4-1:0] node4049;
	wire [4-1:0] node4050;
	wire [4-1:0] node4051;
	wire [4-1:0] node4052;
	wire [4-1:0] node4053;
	wire [4-1:0] node4055;
	wire [4-1:0] node4056;
	wire [4-1:0] node4057;
	wire [4-1:0] node4059;
	wire [4-1:0] node4060;
	wire [4-1:0] node4063;
	wire [4-1:0] node4065;
	wire [4-1:0] node4068;
	wire [4-1:0] node4069;
	wire [4-1:0] node4070;
	wire [4-1:0] node4074;
	wire [4-1:0] node4076;
	wire [4-1:0] node4077;
	wire [4-1:0] node4081;
	wire [4-1:0] node4083;
	wire [4-1:0] node4084;
	wire [4-1:0] node4086;
	wire [4-1:0] node4088;
	wire [4-1:0] node4092;
	wire [4-1:0] node4093;
	wire [4-1:0] node4094;
	wire [4-1:0] node4095;
	wire [4-1:0] node4096;
	wire [4-1:0] node4097;
	wire [4-1:0] node4100;
	wire [4-1:0] node4101;
	wire [4-1:0] node4105;
	wire [4-1:0] node4106;
	wire [4-1:0] node4109;
	wire [4-1:0] node4112;
	wire [4-1:0] node4113;
	wire [4-1:0] node4114;
	wire [4-1:0] node4117;
	wire [4-1:0] node4118;
	wire [4-1:0] node4121;
	wire [4-1:0] node4124;
	wire [4-1:0] node4125;
	wire [4-1:0] node4126;
	wire [4-1:0] node4130;
	wire [4-1:0] node4133;
	wire [4-1:0] node4134;
	wire [4-1:0] node4135;
	wire [4-1:0] node4136;
	wire [4-1:0] node4139;
	wire [4-1:0] node4140;
	wire [4-1:0] node4143;
	wire [4-1:0] node4144;
	wire [4-1:0] node4145;
	wire [4-1:0] node4150;
	wire [4-1:0] node4151;
	wire [4-1:0] node4153;
	wire [4-1:0] node4154;
	wire [4-1:0] node4157;
	wire [4-1:0] node4160;
	wire [4-1:0] node4163;
	wire [4-1:0] node4164;
	wire [4-1:0] node4167;
	wire [4-1:0] node4169;
	wire [4-1:0] node4170;
	wire [4-1:0] node4174;
	wire [4-1:0] node4175;
	wire [4-1:0] node4176;
	wire [4-1:0] node4177;
	wire [4-1:0] node4178;
	wire [4-1:0] node4179;
	wire [4-1:0] node4183;
	wire [4-1:0] node4186;
	wire [4-1:0] node4187;
	wire [4-1:0] node4188;
	wire [4-1:0] node4192;
	wire [4-1:0] node4195;
	wire [4-1:0] node4196;
	wire [4-1:0] node4197;
	wire [4-1:0] node4201;
	wire [4-1:0] node4202;
	wire [4-1:0] node4206;
	wire [4-1:0] node4207;
	wire [4-1:0] node4208;
	wire [4-1:0] node4209;
	wire [4-1:0] node4211;
	wire [4-1:0] node4214;
	wire [4-1:0] node4216;
	wire [4-1:0] node4219;
	wire [4-1:0] node4220;
	wire [4-1:0] node4222;
	wire [4-1:0] node4225;
	wire [4-1:0] node4226;
	wire [4-1:0] node4230;
	wire [4-1:0] node4231;
	wire [4-1:0] node4232;
	wire [4-1:0] node4236;
	wire [4-1:0] node4238;
	wire [4-1:0] node4239;
	wire [4-1:0] node4243;
	wire [4-1:0] node4245;
	wire [4-1:0] node4247;
	wire [4-1:0] node4248;
	wire [4-1:0] node4249;
	wire [4-1:0] node4251;
	wire [4-1:0] node4254;
	wire [4-1:0] node4255;
	wire [4-1:0] node4256;
	wire [4-1:0] node4258;
	wire [4-1:0] node4261;
	wire [4-1:0] node4264;
	wire [4-1:0] node4265;
	wire [4-1:0] node4267;
	wire [4-1:0] node4271;
	wire [4-1:0] node4273;
	wire [4-1:0] node4275;
	wire [4-1:0] node4277;
	wire [4-1:0] node4280;
	wire [4-1:0] node4281;
	wire [4-1:0] node4282;
	wire [4-1:0] node4283;
	wire [4-1:0] node4284;
	wire [4-1:0] node4285;
	wire [4-1:0] node4286;
	wire [4-1:0] node4288;
	wire [4-1:0] node4291;
	wire [4-1:0] node4292;
	wire [4-1:0] node4296;
	wire [4-1:0] node4297;
	wire [4-1:0] node4298;
	wire [4-1:0] node4300;
	wire [4-1:0] node4304;
	wire [4-1:0] node4306;
	wire [4-1:0] node4309;
	wire [4-1:0] node4310;
	wire [4-1:0] node4311;
	wire [4-1:0] node4312;
	wire [4-1:0] node4316;
	wire [4-1:0] node4317;
	wire [4-1:0] node4321;
	wire [4-1:0] node4322;
	wire [4-1:0] node4323;
	wire [4-1:0] node4326;
	wire [4-1:0] node4327;
	wire [4-1:0] node4331;
	wire [4-1:0] node4333;
	wire [4-1:0] node4335;
	wire [4-1:0] node4337;
	wire [4-1:0] node4340;
	wire [4-1:0] node4341;
	wire [4-1:0] node4342;
	wire [4-1:0] node4343;
	wire [4-1:0] node4344;
	wire [4-1:0] node4345;
	wire [4-1:0] node4346;
	wire [4-1:0] node4351;
	wire [4-1:0] node4354;
	wire [4-1:0] node4356;
	wire [4-1:0] node4359;
	wire [4-1:0] node4360;
	wire [4-1:0] node4361;
	wire [4-1:0] node4364;
	wire [4-1:0] node4365;
	wire [4-1:0] node4369;
	wire [4-1:0] node4371;
	wire [4-1:0] node4372;
	wire [4-1:0] node4375;
	wire [4-1:0] node4378;
	wire [4-1:0] node4379;
	wire [4-1:0] node4380;
	wire [4-1:0] node4381;
	wire [4-1:0] node4382;
	wire [4-1:0] node4385;
	wire [4-1:0] node4387;
	wire [4-1:0] node4390;
	wire [4-1:0] node4391;
	wire [4-1:0] node4395;
	wire [4-1:0] node4396;
	wire [4-1:0] node4399;
	wire [4-1:0] node4402;
	wire [4-1:0] node4403;
	wire [4-1:0] node4404;
	wire [4-1:0] node4407;
	wire [4-1:0] node4408;
	wire [4-1:0] node4409;
	wire [4-1:0] node4414;
	wire [4-1:0] node4415;
	wire [4-1:0] node4419;
	wire [4-1:0] node4420;
	wire [4-1:0] node4421;
	wire [4-1:0] node4422;
	wire [4-1:0] node4423;
	wire [4-1:0] node4425;
	wire [4-1:0] node4426;
	wire [4-1:0] node4429;
	wire [4-1:0] node4432;
	wire [4-1:0] node4433;
	wire [4-1:0] node4435;
	wire [4-1:0] node4437;
	wire [4-1:0] node4440;
	wire [4-1:0] node4443;
	wire [4-1:0] node4444;
	wire [4-1:0] node4445;
	wire [4-1:0] node4446;
	wire [4-1:0] node4447;
	wire [4-1:0] node4451;
	wire [4-1:0] node4454;
	wire [4-1:0] node4456;
	wire [4-1:0] node4457;
	wire [4-1:0] node4461;
	wire [4-1:0] node4462;
	wire [4-1:0] node4463;
	wire [4-1:0] node4464;
	wire [4-1:0] node4467;
	wire [4-1:0] node4470;
	wire [4-1:0] node4474;
	wire [4-1:0] node4475;
	wire [4-1:0] node4476;
	wire [4-1:0] node4477;
	wire [4-1:0] node4479;
	wire [4-1:0] node4483;
	wire [4-1:0] node4484;
	wire [4-1:0] node4485;
	wire [4-1:0] node4488;
	wire [4-1:0] node4491;
	wire [4-1:0] node4492;
	wire [4-1:0] node4496;
	wire [4-1:0] node4497;
	wire [4-1:0] node4498;
	wire [4-1:0] node4500;
	wire [4-1:0] node4504;
	wire [4-1:0] node4505;
	wire [4-1:0] node4506;
	wire [4-1:0] node4509;
	wire [4-1:0] node4513;
	wire [4-1:0] node4514;
	wire [4-1:0] node4515;
	wire [4-1:0] node4516;
	wire [4-1:0] node4517;
	wire [4-1:0] node4519;
	wire [4-1:0] node4521;
	wire [4-1:0] node4524;
	wire [4-1:0] node4527;
	wire [4-1:0] node4528;
	wire [4-1:0] node4530;
	wire [4-1:0] node4533;
	wire [4-1:0] node4536;
	wire [4-1:0] node4537;
	wire [4-1:0] node4538;
	wire [4-1:0] node4541;
	wire [4-1:0] node4542;
	wire [4-1:0] node4543;
	wire [4-1:0] node4547;
	wire [4-1:0] node4551;
	wire [4-1:0] node4552;
	wire [4-1:0] node4553;
	wire [4-1:0] node4555;
	wire [4-1:0] node4556;
	wire [4-1:0] node4560;
	wire [4-1:0] node4561;
	wire [4-1:0] node4564;
	wire [4-1:0] node4566;
	wire [4-1:0] node4569;
	wire [4-1:0] node4570;
	wire [4-1:0] node4571;
	wire [4-1:0] node4572;
	wire [4-1:0] node4577;
	wire [4-1:0] node4578;
	wire [4-1:0] node4579;
	wire [4-1:0] node4581;
	wire [4-1:0] node4586;
	wire [4-1:0] node4587;
	wire [4-1:0] node4588;
	wire [4-1:0] node4589;
	wire [4-1:0] node4590;
	wire [4-1:0] node4591;
	wire [4-1:0] node4592;
	wire [4-1:0] node4596;
	wire [4-1:0] node4597;
	wire [4-1:0] node4598;
	wire [4-1:0] node4601;
	wire [4-1:0] node4604;
	wire [4-1:0] node4605;
	wire [4-1:0] node4608;
	wire [4-1:0] node4611;
	wire [4-1:0] node4612;
	wire [4-1:0] node4613;
	wire [4-1:0] node4616;
	wire [4-1:0] node4618;
	wire [4-1:0] node4621;
	wire [4-1:0] node4622;
	wire [4-1:0] node4625;
	wire [4-1:0] node4628;
	wire [4-1:0] node4629;
	wire [4-1:0] node4630;
	wire [4-1:0] node4632;
	wire [4-1:0] node4635;
	wire [4-1:0] node4636;
	wire [4-1:0] node4637;
	wire [4-1:0] node4641;
	wire [4-1:0] node4642;
	wire [4-1:0] node4646;
	wire [4-1:0] node4647;
	wire [4-1:0] node4648;
	wire [4-1:0] node4651;
	wire [4-1:0] node4652;
	wire [4-1:0] node4655;
	wire [4-1:0] node4658;
	wire [4-1:0] node4659;
	wire [4-1:0] node4660;
	wire [4-1:0] node4662;
	wire [4-1:0] node4663;
	wire [4-1:0] node4668;
	wire [4-1:0] node4671;
	wire [4-1:0] node4672;
	wire [4-1:0] node4673;
	wire [4-1:0] node4674;
	wire [4-1:0] node4675;
	wire [4-1:0] node4678;
	wire [4-1:0] node4679;
	wire [4-1:0] node4680;
	wire [4-1:0] node4684;
	wire [4-1:0] node4687;
	wire [4-1:0] node4688;
	wire [4-1:0] node4689;
	wire [4-1:0] node4694;
	wire [4-1:0] node4695;
	wire [4-1:0] node4696;
	wire [4-1:0] node4697;
	wire [4-1:0] node4701;
	wire [4-1:0] node4702;
	wire [4-1:0] node4703;
	wire [4-1:0] node4708;
	wire [4-1:0] node4709;
	wire [4-1:0] node4710;
	wire [4-1:0] node4714;
	wire [4-1:0] node4715;
	wire [4-1:0] node4717;
	wire [4-1:0] node4718;
	wire [4-1:0] node4721;
	wire [4-1:0] node4725;
	wire [4-1:0] node4726;
	wire [4-1:0] node4727;
	wire [4-1:0] node4728;
	wire [4-1:0] node4730;
	wire [4-1:0] node4733;
	wire [4-1:0] node4735;
	wire [4-1:0] node4736;
	wire [4-1:0] node4740;
	wire [4-1:0] node4741;
	wire [4-1:0] node4745;
	wire [4-1:0] node4746;
	wire [4-1:0] node4747;
	wire [4-1:0] node4748;
	wire [4-1:0] node4753;
	wire [4-1:0] node4754;
	wire [4-1:0] node4756;
	wire [4-1:0] node4760;
	wire [4-1:0] node4761;
	wire [4-1:0] node4762;
	wire [4-1:0] node4763;
	wire [4-1:0] node4764;
	wire [4-1:0] node4766;
	wire [4-1:0] node4767;
	wire [4-1:0] node4770;
	wire [4-1:0] node4773;
	wire [4-1:0] node4774;
	wire [4-1:0] node4775;
	wire [4-1:0] node4780;
	wire [4-1:0] node4781;
	wire [4-1:0] node4782;
	wire [4-1:0] node4784;
	wire [4-1:0] node4788;
	wire [4-1:0] node4789;
	wire [4-1:0] node4791;
	wire [4-1:0] node4793;
	wire [4-1:0] node4796;
	wire [4-1:0] node4799;
	wire [4-1:0] node4800;
	wire [4-1:0] node4801;
	wire [4-1:0] node4802;
	wire [4-1:0] node4805;
	wire [4-1:0] node4806;
	wire [4-1:0] node4810;
	wire [4-1:0] node4812;
	wire [4-1:0] node4815;
	wire [4-1:0] node4816;
	wire [4-1:0] node4818;
	wire [4-1:0] node4820;
	wire [4-1:0] node4822;
	wire [4-1:0] node4823;
	wire [4-1:0] node4827;
	wire [4-1:0] node4829;
	wire [4-1:0] node4832;
	wire [4-1:0] node4833;
	wire [4-1:0] node4834;
	wire [4-1:0] node4835;
	wire [4-1:0] node4836;
	wire [4-1:0] node4839;
	wire [4-1:0] node4840;
	wire [4-1:0] node4845;
	wire [4-1:0] node4846;
	wire [4-1:0] node4847;
	wire [4-1:0] node4849;
	wire [4-1:0] node4853;
	wire [4-1:0] node4854;
	wire [4-1:0] node4855;
	wire [4-1:0] node4856;
	wire [4-1:0] node4860;
	wire [4-1:0] node4864;
	wire [4-1:0] node4865;
	wire [4-1:0] node4867;
	wire [4-1:0] node4868;
	wire [4-1:0] node4871;
	wire [4-1:0] node4874;
	wire [4-1:0] node4876;
	wire [4-1:0] node4879;
	wire [4-1:0] node4881;
	wire [4-1:0] node4882;
	wire [4-1:0] node4883;
	wire [4-1:0] node4885;
	wire [4-1:0] node4886;
	wire [4-1:0] node4887;
	wire [4-1:0] node4889;
	wire [4-1:0] node4890;
	wire [4-1:0] node4891;
	wire [4-1:0] node4895;
	wire [4-1:0] node4897;
	wire [4-1:0] node4900;
	wire [4-1:0] node4901;
	wire [4-1:0] node4903;
	wire [4-1:0] node4904;
	wire [4-1:0] node4908;
	wire [4-1:0] node4909;
	wire [4-1:0] node4913;
	wire [4-1:0] node4915;
	wire [4-1:0] node4916;
	wire [4-1:0] node4917;
	wire [4-1:0] node4920;
	wire [4-1:0] node4922;
	wire [4-1:0] node4924;
	wire [4-1:0] node4928;
	wire [4-1:0] node4929;
	wire [4-1:0] node4930;
	wire [4-1:0] node4931;
	wire [4-1:0] node4932;
	wire [4-1:0] node4934;
	wire [4-1:0] node4935;
	wire [4-1:0] node4936;
	wire [4-1:0] node4937;
	wire [4-1:0] node4941;
	wire [4-1:0] node4945;
	wire [4-1:0] node4946;
	wire [4-1:0] node4949;
	wire [4-1:0] node4951;
	wire [4-1:0] node4953;
	wire [4-1:0] node4956;
	wire [4-1:0] node4957;
	wire [4-1:0] node4958;
	wire [4-1:0] node4960;
	wire [4-1:0] node4964;
	wire [4-1:0] node4965;
	wire [4-1:0] node4968;
	wire [4-1:0] node4969;
	wire [4-1:0] node4972;
	wire [4-1:0] node4973;
	wire [4-1:0] node4975;
	wire [4-1:0] node4979;
	wire [4-1:0] node4980;
	wire [4-1:0] node4981;
	wire [4-1:0] node4982;
	wire [4-1:0] node4985;
	wire [4-1:0] node4988;
	wire [4-1:0] node4989;
	wire [4-1:0] node4991;
	wire [4-1:0] node4994;
	wire [4-1:0] node4995;
	wire [4-1:0] node4999;
	wire [4-1:0] node5000;
	wire [4-1:0] node5001;
	wire [4-1:0] node5003;
	wire [4-1:0] node5006;
	wire [4-1:0] node5007;
	wire [4-1:0] node5008;
	wire [4-1:0] node5012;
	wire [4-1:0] node5013;
	wire [4-1:0] node5018;
	wire [4-1:0] node5019;
	wire [4-1:0] node5020;
	wire [4-1:0] node5021;
	wire [4-1:0] node5022;
	wire [4-1:0] node5025;
	wire [4-1:0] node5026;
	wire [4-1:0] node5027;
	wire [4-1:0] node5031;
	wire [4-1:0] node5034;
	wire [4-1:0] node5036;
	wire [4-1:0] node5039;
	wire [4-1:0] node5040;
	wire [4-1:0] node5041;
	wire [4-1:0] node5044;
	wire [4-1:0] node5045;
	wire [4-1:0] node5046;
	wire [4-1:0] node5052;
	wire [4-1:0] node5053;
	wire [4-1:0] node5054;
	wire [4-1:0] node5055;
	wire [4-1:0] node5056;
	wire [4-1:0] node5061;
	wire [4-1:0] node5062;
	wire [4-1:0] node5064;
	wire [4-1:0] node5065;
	wire [4-1:0] node5069;
	wire [4-1:0] node5071;
	wire [4-1:0] node5074;
	wire [4-1:0] node5075;
	wire [4-1:0] node5076;
	wire [4-1:0] node5077;
	wire [4-1:0] node5080;
	wire [4-1:0] node5084;
	wire [4-1:0] node5085;
	wire [4-1:0] node5087;
	wire [4-1:0] node5091;
	wire [4-1:0] node5093;
	wire [4-1:0] node5095;
	wire [4-1:0] node5096;
	wire [4-1:0] node5097;
	wire [4-1:0] node5098;
	wire [4-1:0] node5099;
	wire [4-1:0] node5100;
	wire [4-1:0] node5104;
	wire [4-1:0] node5105;
	wire [4-1:0] node5110;
	wire [4-1:0] node5112;
	wire [4-1:0] node5114;
	wire [4-1:0] node5117;
	wire [4-1:0] node5119;
	wire [4-1:0] node5121;
	wire [4-1:0] node5124;
	wire [4-1:0] node5125;
	wire [4-1:0] node5126;
	wire [4-1:0] node5127;
	wire [4-1:0] node5128;
	wire [4-1:0] node5129;
	wire [4-1:0] node5130;
	wire [4-1:0] node5131;
	wire [4-1:0] node5132;
	wire [4-1:0] node5133;
	wire [4-1:0] node5134;
	wire [4-1:0] node5135;
	wire [4-1:0] node5138;
	wire [4-1:0] node5141;
	wire [4-1:0] node5142;
	wire [4-1:0] node5146;
	wire [4-1:0] node5147;
	wire [4-1:0] node5148;
	wire [4-1:0] node5150;
	wire [4-1:0] node5153;
	wire [4-1:0] node5154;
	wire [4-1:0] node5155;
	wire [4-1:0] node5158;
	wire [4-1:0] node5162;
	wire [4-1:0] node5164;
	wire [4-1:0] node5167;
	wire [4-1:0] node5168;
	wire [4-1:0] node5169;
	wire [4-1:0] node5172;
	wire [4-1:0] node5173;
	wire [4-1:0] node5177;
	wire [4-1:0] node5178;
	wire [4-1:0] node5181;
	wire [4-1:0] node5182;
	wire [4-1:0] node5186;
	wire [4-1:0] node5187;
	wire [4-1:0] node5188;
	wire [4-1:0] node5189;
	wire [4-1:0] node5190;
	wire [4-1:0] node5193;
	wire [4-1:0] node5194;
	wire [4-1:0] node5198;
	wire [4-1:0] node5201;
	wire [4-1:0] node5202;
	wire [4-1:0] node5204;
	wire [4-1:0] node5207;
	wire [4-1:0] node5208;
	wire [4-1:0] node5211;
	wire [4-1:0] node5212;
	wire [4-1:0] node5215;
	wire [4-1:0] node5218;
	wire [4-1:0] node5219;
	wire [4-1:0] node5220;
	wire [4-1:0] node5221;
	wire [4-1:0] node5224;
	wire [4-1:0] node5227;
	wire [4-1:0] node5229;
	wire [4-1:0] node5232;
	wire [4-1:0] node5233;
	wire [4-1:0] node5236;
	wire [4-1:0] node5238;
	wire [4-1:0] node5240;
	wire [4-1:0] node5243;
	wire [4-1:0] node5244;
	wire [4-1:0] node5245;
	wire [4-1:0] node5246;
	wire [4-1:0] node5247;
	wire [4-1:0] node5248;
	wire [4-1:0] node5249;
	wire [4-1:0] node5250;
	wire [4-1:0] node5256;
	wire [4-1:0] node5258;
	wire [4-1:0] node5259;
	wire [4-1:0] node5263;
	wire [4-1:0] node5264;
	wire [4-1:0] node5266;
	wire [4-1:0] node5269;
	wire [4-1:0] node5271;
	wire [4-1:0] node5274;
	wire [4-1:0] node5275;
	wire [4-1:0] node5276;
	wire [4-1:0] node5277;
	wire [4-1:0] node5280;
	wire [4-1:0] node5282;
	wire [4-1:0] node5285;
	wire [4-1:0] node5287;
	wire [4-1:0] node5288;
	wire [4-1:0] node5289;
	wire [4-1:0] node5294;
	wire [4-1:0] node5295;
	wire [4-1:0] node5296;
	wire [4-1:0] node5298;
	wire [4-1:0] node5301;
	wire [4-1:0] node5304;
	wire [4-1:0] node5307;
	wire [4-1:0] node5308;
	wire [4-1:0] node5309;
	wire [4-1:0] node5310;
	wire [4-1:0] node5311;
	wire [4-1:0] node5312;
	wire [4-1:0] node5316;
	wire [4-1:0] node5319;
	wire [4-1:0] node5320;
	wire [4-1:0] node5321;
	wire [4-1:0] node5326;
	wire [4-1:0] node5327;
	wire [4-1:0] node5328;
	wire [4-1:0] node5330;
	wire [4-1:0] node5331;
	wire [4-1:0] node5334;
	wire [4-1:0] node5337;
	wire [4-1:0] node5338;
	wire [4-1:0] node5342;
	wire [4-1:0] node5343;
	wire [4-1:0] node5345;
	wire [4-1:0] node5347;
	wire [4-1:0] node5351;
	wire [4-1:0] node5352;
	wire [4-1:0] node5353;
	wire [4-1:0] node5355;
	wire [4-1:0] node5358;
	wire [4-1:0] node5359;
	wire [4-1:0] node5360;
	wire [4-1:0] node5365;
	wire [4-1:0] node5366;
	wire [4-1:0] node5367;
	wire [4-1:0] node5370;
	wire [4-1:0] node5373;
	wire [4-1:0] node5374;
	wire [4-1:0] node5376;
	wire [4-1:0] node5377;
	wire [4-1:0] node5380;
	wire [4-1:0] node5383;
	wire [4-1:0] node5386;
	wire [4-1:0] node5388;
	wire [4-1:0] node5389;
	wire [4-1:0] node5390;
	wire [4-1:0] node5391;
	wire [4-1:0] node5392;
	wire [4-1:0] node5394;
	wire [4-1:0] node5395;
	wire [4-1:0] node5396;
	wire [4-1:0] node5400;
	wire [4-1:0] node5401;
	wire [4-1:0] node5405;
	wire [4-1:0] node5406;
	wire [4-1:0] node5411;
	wire [4-1:0] node5412;
	wire [4-1:0] node5413;
	wire [4-1:0] node5414;
	wire [4-1:0] node5417;
	wire [4-1:0] node5418;
	wire [4-1:0] node5422;
	wire [4-1:0] node5423;
	wire [4-1:0] node5425;
	wire [4-1:0] node5428;
	wire [4-1:0] node5431;
	wire [4-1:0] node5432;
	wire [4-1:0] node5434;
	wire [4-1:0] node5435;
	wire [4-1:0] node5438;
	wire [4-1:0] node5441;
	wire [4-1:0] node5443;
	wire [4-1:0] node5446;
	wire [4-1:0] node5447;
	wire [4-1:0] node5448;
	wire [4-1:0] node5449;
	wire [4-1:0] node5450;
	wire [4-1:0] node5453;
	wire [4-1:0] node5456;
	wire [4-1:0] node5457;
	wire [4-1:0] node5458;
	wire [4-1:0] node5460;
	wire [4-1:0] node5464;
	wire [4-1:0] node5466;
	wire [4-1:0] node5467;
	wire [4-1:0] node5471;
	wire [4-1:0] node5472;
	wire [4-1:0] node5473;
	wire [4-1:0] node5476;
	wire [4-1:0] node5477;
	wire [4-1:0] node5481;
	wire [4-1:0] node5482;
	wire [4-1:0] node5485;
	wire [4-1:0] node5488;
	wire [4-1:0] node5489;
	wire [4-1:0] node5490;
	wire [4-1:0] node5491;
	wire [4-1:0] node5493;
	wire [4-1:0] node5494;
	wire [4-1:0] node5498;
	wire [4-1:0] node5499;
	wire [4-1:0] node5503;
	wire [4-1:0] node5506;
	wire [4-1:0] node5507;
	wire [4-1:0] node5508;
	wire [4-1:0] node5509;
	wire [4-1:0] node5514;
	wire [4-1:0] node5516;
	wire [4-1:0] node5520;
	wire [4-1:0] node5521;
	wire [4-1:0] node5522;
	wire [4-1:0] node5523;
	wire [4-1:0] node5524;
	wire [4-1:0] node5525;
	wire [4-1:0] node5526;
	wire [4-1:0] node5527;
	wire [4-1:0] node5529;
	wire [4-1:0] node5531;
	wire [4-1:0] node5534;
	wire [4-1:0] node5535;
	wire [4-1:0] node5536;
	wire [4-1:0] node5539;
	wire [4-1:0] node5543;
	wire [4-1:0] node5544;
	wire [4-1:0] node5545;
	wire [4-1:0] node5548;
	wire [4-1:0] node5551;
	wire [4-1:0] node5552;
	wire [4-1:0] node5555;
	wire [4-1:0] node5558;
	wire [4-1:0] node5559;
	wire [4-1:0] node5560;
	wire [4-1:0] node5561;
	wire [4-1:0] node5562;
	wire [4-1:0] node5566;
	wire [4-1:0] node5569;
	wire [4-1:0] node5570;
	wire [4-1:0] node5571;
	wire [4-1:0] node5572;
	wire [4-1:0] node5577;
	wire [4-1:0] node5580;
	wire [4-1:0] node5581;
	wire [4-1:0] node5582;
	wire [4-1:0] node5583;
	wire [4-1:0] node5585;
	wire [4-1:0] node5587;
	wire [4-1:0] node5591;
	wire [4-1:0] node5593;
	wire [4-1:0] node5594;
	wire [4-1:0] node5596;
	wire [4-1:0] node5600;
	wire [4-1:0] node5601;
	wire [4-1:0] node5602;
	wire [4-1:0] node5606;
	wire [4-1:0] node5607;
	wire [4-1:0] node5610;
	wire [4-1:0] node5613;
	wire [4-1:0] node5614;
	wire [4-1:0] node5615;
	wire [4-1:0] node5616;
	wire [4-1:0] node5617;
	wire [4-1:0] node5618;
	wire [4-1:0] node5619;
	wire [4-1:0] node5624;
	wire [4-1:0] node5625;
	wire [4-1:0] node5629;
	wire [4-1:0] node5630;
	wire [4-1:0] node5631;
	wire [4-1:0] node5635;
	wire [4-1:0] node5637;
	wire [4-1:0] node5640;
	wire [4-1:0] node5641;
	wire [4-1:0] node5642;
	wire [4-1:0] node5644;
	wire [4-1:0] node5647;
	wire [4-1:0] node5649;
	wire [4-1:0] node5652;
	wire [4-1:0] node5653;
	wire [4-1:0] node5654;
	wire [4-1:0] node5658;
	wire [4-1:0] node5659;
	wire [4-1:0] node5661;
	wire [4-1:0] node5665;
	wire [4-1:0] node5666;
	wire [4-1:0] node5667;
	wire [4-1:0] node5668;
	wire [4-1:0] node5670;
	wire [4-1:0] node5671;
	wire [4-1:0] node5675;
	wire [4-1:0] node5677;
	wire [4-1:0] node5680;
	wire [4-1:0] node5681;
	wire [4-1:0] node5683;
	wire [4-1:0] node5686;
	wire [4-1:0] node5689;
	wire [4-1:0] node5690;
	wire [4-1:0] node5691;
	wire [4-1:0] node5694;
	wire [4-1:0] node5697;
	wire [4-1:0] node5700;
	wire [4-1:0] node5701;
	wire [4-1:0] node5702;
	wire [4-1:0] node5703;
	wire [4-1:0] node5704;
	wire [4-1:0] node5705;
	wire [4-1:0] node5706;
	wire [4-1:0] node5710;
	wire [4-1:0] node5713;
	wire [4-1:0] node5714;
	wire [4-1:0] node5716;
	wire [4-1:0] node5720;
	wire [4-1:0] node5721;
	wire [4-1:0] node5722;
	wire [4-1:0] node5723;
	wire [4-1:0] node5727;
	wire [4-1:0] node5729;
	wire [4-1:0] node5732;
	wire [4-1:0] node5733;
	wire [4-1:0] node5737;
	wire [4-1:0] node5738;
	wire [4-1:0] node5739;
	wire [4-1:0] node5740;
	wire [4-1:0] node5742;
	wire [4-1:0] node5743;
	wire [4-1:0] node5747;
	wire [4-1:0] node5748;
	wire [4-1:0] node5751;
	wire [4-1:0] node5754;
	wire [4-1:0] node5755;
	wire [4-1:0] node5758;
	wire [4-1:0] node5760;
	wire [4-1:0] node5762;
	wire [4-1:0] node5765;
	wire [4-1:0] node5766;
	wire [4-1:0] node5767;
	wire [4-1:0] node5770;
	wire [4-1:0] node5771;
	wire [4-1:0] node5775;
	wire [4-1:0] node5776;
	wire [4-1:0] node5778;
	wire [4-1:0] node5779;
	wire [4-1:0] node5783;
	wire [4-1:0] node5784;
	wire [4-1:0] node5787;
	wire [4-1:0] node5790;
	wire [4-1:0] node5791;
	wire [4-1:0] node5792;
	wire [4-1:0] node5793;
	wire [4-1:0] node5794;
	wire [4-1:0] node5795;
	wire [4-1:0] node5800;
	wire [4-1:0] node5801;
	wire [4-1:0] node5803;
	wire [4-1:0] node5804;
	wire [4-1:0] node5808;
	wire [4-1:0] node5811;
	wire [4-1:0] node5812;
	wire [4-1:0] node5813;
	wire [4-1:0] node5814;
	wire [4-1:0] node5815;
	wire [4-1:0] node5818;
	wire [4-1:0] node5822;
	wire [4-1:0] node5825;
	wire [4-1:0] node5826;
	wire [4-1:0] node5827;
	wire [4-1:0] node5829;
	wire [4-1:0] node5833;
	wire [4-1:0] node5835;
	wire [4-1:0] node5838;
	wire [4-1:0] node5839;
	wire [4-1:0] node5840;
	wire [4-1:0] node5842;
	wire [4-1:0] node5846;
	wire [4-1:0] node5847;
	wire [4-1:0] node5848;
	wire [4-1:0] node5850;
	wire [4-1:0] node5854;
	wire [4-1:0] node5855;
	wire [4-1:0] node5856;
	wire [4-1:0] node5861;
	wire [4-1:0] node5862;
	wire [4-1:0] node5863;
	wire [4-1:0] node5864;
	wire [4-1:0] node5865;
	wire [4-1:0] node5866;
	wire [4-1:0] node5867;
	wire [4-1:0] node5868;
	wire [4-1:0] node5873;
	wire [4-1:0] node5874;
	wire [4-1:0] node5875;
	wire [4-1:0] node5879;
	wire [4-1:0] node5883;
	wire [4-1:0] node5884;
	wire [4-1:0] node5885;
	wire [4-1:0] node5886;
	wire [4-1:0] node5888;
	wire [4-1:0] node5891;
	wire [4-1:0] node5894;
	wire [4-1:0] node5895;
	wire [4-1:0] node5898;
	wire [4-1:0] node5901;
	wire [4-1:0] node5902;
	wire [4-1:0] node5904;
	wire [4-1:0] node5907;
	wire [4-1:0] node5908;
	wire [4-1:0] node5911;
	wire [4-1:0] node5914;
	wire [4-1:0] node5915;
	wire [4-1:0] node5916;
	wire [4-1:0] node5917;
	wire [4-1:0] node5919;
	wire [4-1:0] node5922;
	wire [4-1:0] node5923;
	wire [4-1:0] node5924;
	wire [4-1:0] node5928;
	wire [4-1:0] node5929;
	wire [4-1:0] node5931;
	wire [4-1:0] node5935;
	wire [4-1:0] node5936;
	wire [4-1:0] node5937;
	wire [4-1:0] node5938;
	wire [4-1:0] node5943;
	wire [4-1:0] node5944;
	wire [4-1:0] node5945;
	wire [4-1:0] node5949;
	wire [4-1:0] node5952;
	wire [4-1:0] node5953;
	wire [4-1:0] node5954;
	wire [4-1:0] node5955;
	wire [4-1:0] node5956;
	wire [4-1:0] node5960;
	wire [4-1:0] node5963;
	wire [4-1:0] node5964;
	wire [4-1:0] node5968;
	wire [4-1:0] node5969;
	wire [4-1:0] node5971;
	wire [4-1:0] node5974;
	wire [4-1:0] node5975;
	wire [4-1:0] node5977;
	wire [4-1:0] node5980;
	wire [4-1:0] node5984;
	wire [4-1:0] node5985;
	wire [4-1:0] node5986;
	wire [4-1:0] node5987;
	wire [4-1:0] node5988;
	wire [4-1:0] node5989;
	wire [4-1:0] node5990;
	wire [4-1:0] node5991;
	wire [4-1:0] node5994;
	wire [4-1:0] node5996;
	wire [4-1:0] node5999;
	wire [4-1:0] node6000;
	wire [4-1:0] node6002;
	wire [4-1:0] node6005;
	wire [4-1:0] node6007;
	wire [4-1:0] node6010;
	wire [4-1:0] node6011;
	wire [4-1:0] node6013;
	wire [4-1:0] node6014;
	wire [4-1:0] node6017;
	wire [4-1:0] node6020;
	wire [4-1:0] node6021;
	wire [4-1:0] node6022;
	wire [4-1:0] node6026;
	wire [4-1:0] node6027;
	wire [4-1:0] node6031;
	wire [4-1:0] node6032;
	wire [4-1:0] node6033;
	wire [4-1:0] node6034;
	wire [4-1:0] node6037;
	wire [4-1:0] node6039;
	wire [4-1:0] node6042;
	wire [4-1:0] node6043;
	wire [4-1:0] node6046;
	wire [4-1:0] node6047;
	wire [4-1:0] node6051;
	wire [4-1:0] node6052;
	wire [4-1:0] node6053;
	wire [4-1:0] node6054;
	wire [4-1:0] node6058;
	wire [4-1:0] node6059;
	wire [4-1:0] node6064;
	wire [4-1:0] node6065;
	wire [4-1:0] node6066;
	wire [4-1:0] node6067;
	wire [4-1:0] node6069;
	wire [4-1:0] node6070;
	wire [4-1:0] node6073;
	wire [4-1:0] node6076;
	wire [4-1:0] node6078;
	wire [4-1:0] node6081;
	wire [4-1:0] node6082;
	wire [4-1:0] node6084;
	wire [4-1:0] node6085;
	wire [4-1:0] node6089;
	wire [4-1:0] node6091;
	wire [4-1:0] node6094;
	wire [4-1:0] node6095;
	wire [4-1:0] node6096;
	wire [4-1:0] node6097;
	wire [4-1:0] node6100;
	wire [4-1:0] node6101;
	wire [4-1:0] node6102;
	wire [4-1:0] node6106;
	wire [4-1:0] node6109;
	wire [4-1:0] node6110;
	wire [4-1:0] node6111;
	wire [4-1:0] node6115;
	wire [4-1:0] node6119;
	wire [4-1:0] node6120;
	wire [4-1:0] node6121;
	wire [4-1:0] node6122;
	wire [4-1:0] node6123;
	wire [4-1:0] node6124;
	wire [4-1:0] node6125;
	wire [4-1:0] node6127;
	wire [4-1:0] node6131;
	wire [4-1:0] node6134;
	wire [4-1:0] node6135;
	wire [4-1:0] node6137;
	wire [4-1:0] node6140;
	wire [4-1:0] node6142;
	wire [4-1:0] node6143;
	wire [4-1:0] node6146;
	wire [4-1:0] node6149;
	wire [4-1:0] node6150;
	wire [4-1:0] node6151;
	wire [4-1:0] node6152;
	wire [4-1:0] node6153;
	wire [4-1:0] node6157;
	wire [4-1:0] node6160;
	wire [4-1:0] node6161;
	wire [4-1:0] node6164;
	wire [4-1:0] node6167;
	wire [4-1:0] node6168;
	wire [4-1:0] node6170;
	wire [4-1:0] node6172;
	wire [4-1:0] node6175;
	wire [4-1:0] node6178;
	wire [4-1:0] node6179;
	wire [4-1:0] node6180;
	wire [4-1:0] node6181;
	wire [4-1:0] node6185;
	wire [4-1:0] node6187;
	wire [4-1:0] node6189;
	wire [4-1:0] node6192;
	wire [4-1:0] node6193;
	wire [4-1:0] node6194;
	wire [4-1:0] node6196;
	wire [4-1:0] node6199;
	wire [4-1:0] node6200;
	wire [4-1:0] node6202;
	wire [4-1:0] node6206;
	wire [4-1:0] node6207;
	wire [4-1:0] node6211;
	wire [4-1:0] node6212;
	wire [4-1:0] node6213;
	wire [4-1:0] node6214;
	wire [4-1:0] node6215;
	wire [4-1:0] node6217;
	wire [4-1:0] node6220;
	wire [4-1:0] node6221;
	wire [4-1:0] node6224;
	wire [4-1:0] node6227;
	wire [4-1:0] node6228;
	wire [4-1:0] node6229;
	wire [4-1:0] node6232;
	wire [4-1:0] node6235;
	wire [4-1:0] node6238;
	wire [4-1:0] node6239;
	wire [4-1:0] node6240;
	wire [4-1:0] node6243;
	wire [4-1:0] node6244;
	wire [4-1:0] node6248;
	wire [4-1:0] node6249;
	wire [4-1:0] node6252;
	wire [4-1:0] node6253;
	wire [4-1:0] node6257;
	wire [4-1:0] node6258;
	wire [4-1:0] node6259;
	wire [4-1:0] node6260;
	wire [4-1:0] node6261;
	wire [4-1:0] node6264;
	wire [4-1:0] node6266;
	wire [4-1:0] node6269;
	wire [4-1:0] node6270;
	wire [4-1:0] node6271;
	wire [4-1:0] node6276;
	wire [4-1:0] node6277;
	wire [4-1:0] node6280;
	wire [4-1:0] node6282;
	wire [4-1:0] node6284;
	wire [4-1:0] node6287;
	wire [4-1:0] node6288;
	wire [4-1:0] node6289;
	wire [4-1:0] node6291;
	wire [4-1:0] node6294;
	wire [4-1:0] node6295;
	wire [4-1:0] node6298;
	wire [4-1:0] node6302;
	wire [4-1:0] node6303;
	wire [4-1:0] node6304;
	wire [4-1:0] node6305;
	wire [4-1:0] node6306;
	wire [4-1:0] node6307;
	wire [4-1:0] node6308;
	wire [4-1:0] node6311;
	wire [4-1:0] node6314;
	wire [4-1:0] node6315;
	wire [4-1:0] node6316;
	wire [4-1:0] node6320;
	wire [4-1:0] node6323;
	wire [4-1:0] node6324;
	wire [4-1:0] node6325;
	wire [4-1:0] node6326;
	wire [4-1:0] node6330;
	wire [4-1:0] node6331;
	wire [4-1:0] node6334;
	wire [4-1:0] node6338;
	wire [4-1:0] node6339;
	wire [4-1:0] node6340;
	wire [4-1:0] node6341;
	wire [4-1:0] node6342;
	wire [4-1:0] node6346;
	wire [4-1:0] node6349;
	wire [4-1:0] node6350;
	wire [4-1:0] node6351;
	wire [4-1:0] node6355;
	wire [4-1:0] node6358;
	wire [4-1:0] node6359;
	wire [4-1:0] node6360;
	wire [4-1:0] node6361;
	wire [4-1:0] node6363;
	wire [4-1:0] node6365;
	wire [4-1:0] node6369;
	wire [4-1:0] node6371;
	wire [4-1:0] node6372;
	wire [4-1:0] node6376;
	wire [4-1:0] node6377;
	wire [4-1:0] node6380;
	wire [4-1:0] node6383;
	wire [4-1:0] node6384;
	wire [4-1:0] node6385;
	wire [4-1:0] node6386;
	wire [4-1:0] node6387;
	wire [4-1:0] node6388;
	wire [4-1:0] node6390;
	wire [4-1:0] node6393;
	wire [4-1:0] node6395;
	wire [4-1:0] node6399;
	wire [4-1:0] node6401;
	wire [4-1:0] node6403;
	wire [4-1:0] node6406;
	wire [4-1:0] node6407;
	wire [4-1:0] node6408;
	wire [4-1:0] node6409;
	wire [4-1:0] node6410;
	wire [4-1:0] node6416;
	wire [4-1:0] node6418;
	wire [4-1:0] node6419;
	wire [4-1:0] node6422;
	wire [4-1:0] node6425;
	wire [4-1:0] node6426;
	wire [4-1:0] node6427;
	wire [4-1:0] node6431;
	wire [4-1:0] node6432;
	wire [4-1:0] node6433;
	wire [4-1:0] node6438;
	wire [4-1:0] node6439;
	wire [4-1:0] node6440;
	wire [4-1:0] node6441;
	wire [4-1:0] node6442;
	wire [4-1:0] node6443;
	wire [4-1:0] node6444;
	wire [4-1:0] node6448;
	wire [4-1:0] node6449;
	wire [4-1:0] node6452;
	wire [4-1:0] node6455;
	wire [4-1:0] node6456;
	wire [4-1:0] node6458;
	wire [4-1:0] node6459;
	wire [4-1:0] node6463;
	wire [4-1:0] node6464;
	wire [4-1:0] node6466;
	wire [4-1:0] node6470;
	wire [4-1:0] node6471;
	wire [4-1:0] node6473;
	wire [4-1:0] node6474;
	wire [4-1:0] node6478;
	wire [4-1:0] node6479;
	wire [4-1:0] node6481;
	wire [4-1:0] node6484;
	wire [4-1:0] node6485;
	wire [4-1:0] node6486;
	wire [4-1:0] node6489;
	wire [4-1:0] node6493;
	wire [4-1:0] node6494;
	wire [4-1:0] node6495;
	wire [4-1:0] node6496;
	wire [4-1:0] node6497;
	wire [4-1:0] node6501;
	wire [4-1:0] node6502;
	wire [4-1:0] node6503;
	wire [4-1:0] node6507;
	wire [4-1:0] node6510;
	wire [4-1:0] node6511;
	wire [4-1:0] node6512;
	wire [4-1:0] node6517;
	wire [4-1:0] node6518;
	wire [4-1:0] node6520;
	wire [4-1:0] node6521;
	wire [4-1:0] node6522;
	wire [4-1:0] node6528;
	wire [4-1:0] node6529;
	wire [4-1:0] node6530;
	wire [4-1:0] node6531;
	wire [4-1:0] node6533;
	wire [4-1:0] node6536;
	wire [4-1:0] node6537;
	wire [4-1:0] node6540;
	wire [4-1:0] node6541;
	wire [4-1:0] node6544;
	wire [4-1:0] node6547;
	wire [4-1:0] node6548;
	wire [4-1:0] node6549;
	wire [4-1:0] node6550;
	wire [4-1:0] node6554;
	wire [4-1:0] node6558;
	wire [4-1:0] node6559;
	wire [4-1:0] node6561;
	wire [4-1:0] node6562;
	wire [4-1:0] node6567;
	wire [4-1:0] node6568;
	wire [4-1:0] node6569;
	wire [4-1:0] node6570;
	wire [4-1:0] node6571;
	wire [4-1:0] node6573;
	wire [4-1:0] node6574;
	wire [4-1:0] node6575;
	wire [4-1:0] node6576;
	wire [4-1:0] node6577;
	wire [4-1:0] node6578;
	wire [4-1:0] node6579;
	wire [4-1:0] node6586;
	wire [4-1:0] node6587;
	wire [4-1:0] node6589;
	wire [4-1:0] node6590;
	wire [4-1:0] node6592;
	wire [4-1:0] node6595;
	wire [4-1:0] node6596;
	wire [4-1:0] node6600;
	wire [4-1:0] node6601;
	wire [4-1:0] node6602;
	wire [4-1:0] node6607;
	wire [4-1:0] node6608;
	wire [4-1:0] node6609;
	wire [4-1:0] node6610;
	wire [4-1:0] node6614;
	wire [4-1:0] node6615;
	wire [4-1:0] node6618;
	wire [4-1:0] node6619;
	wire [4-1:0] node6623;
	wire [4-1:0] node6624;
	wire [4-1:0] node6625;
	wire [4-1:0] node6627;
	wire [4-1:0] node6630;
	wire [4-1:0] node6633;
	wire [4-1:0] node6635;
	wire [4-1:0] node6636;
	wire [4-1:0] node6640;
	wire [4-1:0] node6641;
	wire [4-1:0] node6642;
	wire [4-1:0] node6643;
	wire [4-1:0] node6644;
	wire [4-1:0] node6645;
	wire [4-1:0] node6648;
	wire [4-1:0] node6649;
	wire [4-1:0] node6653;
	wire [4-1:0] node6655;
	wire [4-1:0] node6656;
	wire [4-1:0] node6658;
	wire [4-1:0] node6662;
	wire [4-1:0] node6663;
	wire [4-1:0] node6664;
	wire [4-1:0] node6667;
	wire [4-1:0] node6668;
	wire [4-1:0] node6670;
	wire [4-1:0] node6671;
	wire [4-1:0] node6675;
	wire [4-1:0] node6677;
	wire [4-1:0] node6680;
	wire [4-1:0] node6683;
	wire [4-1:0] node6684;
	wire [4-1:0] node6685;
	wire [4-1:0] node6686;
	wire [4-1:0] node6687;
	wire [4-1:0] node6691;
	wire [4-1:0] node6692;
	wire [4-1:0] node6696;
	wire [4-1:0] node6698;
	wire [4-1:0] node6701;
	wire [4-1:0] node6702;
	wire [4-1:0] node6704;
	wire [4-1:0] node6705;
	wire [4-1:0] node6709;
	wire [4-1:0] node6710;
	wire [4-1:0] node6713;
	wire [4-1:0] node6716;
	wire [4-1:0] node6717;
	wire [4-1:0] node6718;
	wire [4-1:0] node6719;
	wire [4-1:0] node6720;
	wire [4-1:0] node6724;
	wire [4-1:0] node6725;
	wire [4-1:0] node6727;
	wire [4-1:0] node6730;
	wire [4-1:0] node6733;
	wire [4-1:0] node6734;
	wire [4-1:0] node6735;
	wire [4-1:0] node6736;
	wire [4-1:0] node6741;
	wire [4-1:0] node6742;
	wire [4-1:0] node6744;
	wire [4-1:0] node6746;
	wire [4-1:0] node6749;
	wire [4-1:0] node6751;
	wire [4-1:0] node6753;
	wire [4-1:0] node6755;
	wire [4-1:0] node6758;
	wire [4-1:0] node6759;
	wire [4-1:0] node6760;
	wire [4-1:0] node6761;
	wire [4-1:0] node6763;
	wire [4-1:0] node6764;
	wire [4-1:0] node6767;
	wire [4-1:0] node6769;
	wire [4-1:0] node6772;
	wire [4-1:0] node6774;
	wire [4-1:0] node6777;
	wire [4-1:0] node6778;
	wire [4-1:0] node6779;
	wire [4-1:0] node6783;
	wire [4-1:0] node6786;
	wire [4-1:0] node6787;
	wire [4-1:0] node6788;
	wire [4-1:0] node6790;
	wire [4-1:0] node6794;
	wire [4-1:0] node6795;
	wire [4-1:0] node6798;
	wire [4-1:0] node6799;
	wire [4-1:0] node6803;
	wire [4-1:0] node6805;
	wire [4-1:0] node6807;
	wire [4-1:0] node6808;
	wire [4-1:0] node6809;
	wire [4-1:0] node6810;
	wire [4-1:0] node6811;
	wire [4-1:0] node6812;
	wire [4-1:0] node6814;
	wire [4-1:0] node6819;
	wire [4-1:0] node6820;
	wire [4-1:0] node6822;
	wire [4-1:0] node6825;
	wire [4-1:0] node6827;
	wire [4-1:0] node6829;
	wire [4-1:0] node6832;
	wire [4-1:0] node6834;
	wire [4-1:0] node6835;
	wire [4-1:0] node6837;
	wire [4-1:0] node6840;
	wire [4-1:0] node6841;
	wire [4-1:0] node6844;
	wire [4-1:0] node6847;
	wire [4-1:0] node6848;
	wire [4-1:0] node6849;
	wire [4-1:0] node6850;
	wire [4-1:0] node6851;
	wire [4-1:0] node6855;
	wire [4-1:0] node6858;
	wire [4-1:0] node6861;
	wire [4-1:0] node6862;
	wire [4-1:0] node6863;
	wire [4-1:0] node6865;
	wire [4-1:0] node6868;
	wire [4-1:0] node6869;
	wire [4-1:0] node6873;
	wire [4-1:0] node6874;
	wire [4-1:0] node6878;
	wire [4-1:0] node6879;
	wire [4-1:0] node6880;
	wire [4-1:0] node6881;
	wire [4-1:0] node6882;
	wire [4-1:0] node6883;
	wire [4-1:0] node6884;
	wire [4-1:0] node6885;
	wire [4-1:0] node6887;
	wire [4-1:0] node6890;
	wire [4-1:0] node6892;
	wire [4-1:0] node6896;
	wire [4-1:0] node6897;
	wire [4-1:0] node6899;
	wire [4-1:0] node6902;
	wire [4-1:0] node6903;
	wire [4-1:0] node6904;
	wire [4-1:0] node6907;
	wire [4-1:0] node6910;
	wire [4-1:0] node6911;
	wire [4-1:0] node6914;
	wire [4-1:0] node6917;
	wire [4-1:0] node6918;
	wire [4-1:0] node6919;
	wire [4-1:0] node6920;
	wire [4-1:0] node6923;
	wire [4-1:0] node6925;
	wire [4-1:0] node6928;
	wire [4-1:0] node6929;
	wire [4-1:0] node6932;
	wire [4-1:0] node6933;
	wire [4-1:0] node6935;
	wire [4-1:0] node6937;
	wire [4-1:0] node6940;
	wire [4-1:0] node6942;
	wire [4-1:0] node6945;
	wire [4-1:0] node6946;
	wire [4-1:0] node6947;
	wire [4-1:0] node6948;
	wire [4-1:0] node6952;
	wire [4-1:0] node6955;
	wire [4-1:0] node6956;
	wire [4-1:0] node6957;
	wire [4-1:0] node6958;
	wire [4-1:0] node6961;
	wire [4-1:0] node6964;
	wire [4-1:0] node6967;
	wire [4-1:0] node6968;
	wire [4-1:0] node6969;
	wire [4-1:0] node6970;
	wire [4-1:0] node6976;
	wire [4-1:0] node6977;
	wire [4-1:0] node6978;
	wire [4-1:0] node6979;
	wire [4-1:0] node6980;
	wire [4-1:0] node6983;
	wire [4-1:0] node6984;
	wire [4-1:0] node6985;
	wire [4-1:0] node6990;
	wire [4-1:0] node6991;
	wire [4-1:0] node6992;
	wire [4-1:0] node6993;
	wire [4-1:0] node6998;
	wire [4-1:0] node7000;
	wire [4-1:0] node7001;
	wire [4-1:0] node7003;
	wire [4-1:0] node7006;
	wire [4-1:0] node7009;
	wire [4-1:0] node7010;
	wire [4-1:0] node7012;
	wire [4-1:0] node7015;
	wire [4-1:0] node7016;
	wire [4-1:0] node7019;
	wire [4-1:0] node7020;
	wire [4-1:0] node7023;
	wire [4-1:0] node7025;
	wire [4-1:0] node7028;
	wire [4-1:0] node7029;
	wire [4-1:0] node7030;
	wire [4-1:0] node7031;
	wire [4-1:0] node7033;
	wire [4-1:0] node7036;
	wire [4-1:0] node7037;
	wire [4-1:0] node7041;
	wire [4-1:0] node7042;
	wire [4-1:0] node7046;
	wire [4-1:0] node7047;
	wire [4-1:0] node7048;
	wire [4-1:0] node7051;
	wire [4-1:0] node7052;
	wire [4-1:0] node7056;
	wire [4-1:0] node7057;
	wire [4-1:0] node7060;
	wire [4-1:0] node7062;
	wire [4-1:0] node7063;
	wire [4-1:0] node7067;
	wire [4-1:0] node7068;
	wire [4-1:0] node7069;
	wire [4-1:0] node7070;
	wire [4-1:0] node7071;
	wire [4-1:0] node7072;
	wire [4-1:0] node7074;
	wire [4-1:0] node7078;
	wire [4-1:0] node7079;
	wire [4-1:0] node7081;
	wire [4-1:0] node7084;
	wire [4-1:0] node7086;
	wire [4-1:0] node7087;
	wire [4-1:0] node7091;
	wire [4-1:0] node7092;
	wire [4-1:0] node7093;
	wire [4-1:0] node7094;
	wire [4-1:0] node7098;
	wire [4-1:0] node7099;
	wire [4-1:0] node7103;
	wire [4-1:0] node7104;
	wire [4-1:0] node7105;
	wire [4-1:0] node7108;
	wire [4-1:0] node7110;
	wire [4-1:0] node7113;
	wire [4-1:0] node7114;
	wire [4-1:0] node7118;
	wire [4-1:0] node7119;
	wire [4-1:0] node7120;
	wire [4-1:0] node7121;
	wire [4-1:0] node7123;
	wire [4-1:0] node7125;
	wire [4-1:0] node7127;
	wire [4-1:0] node7131;
	wire [4-1:0] node7132;
	wire [4-1:0] node7134;
	wire [4-1:0] node7137;
	wire [4-1:0] node7140;
	wire [4-1:0] node7141;
	wire [4-1:0] node7143;
	wire [4-1:0] node7145;
	wire [4-1:0] node7148;
	wire [4-1:0] node7149;
	wire [4-1:0] node7151;
	wire [4-1:0] node7152;
	wire [4-1:0] node7155;
	wire [4-1:0] node7158;
	wire [4-1:0] node7160;
	wire [4-1:0] node7163;
	wire [4-1:0] node7164;
	wire [4-1:0] node7165;
	wire [4-1:0] node7166;
	wire [4-1:0] node7167;
	wire [4-1:0] node7169;
	wire [4-1:0] node7172;
	wire [4-1:0] node7174;
	wire [4-1:0] node7177;
	wire [4-1:0] node7179;
	wire [4-1:0] node7182;
	wire [4-1:0] node7183;
	wire [4-1:0] node7186;
	wire [4-1:0] node7188;
	wire [4-1:0] node7191;
	wire [4-1:0] node7192;
	wire [4-1:0] node7193;
	wire [4-1:0] node7195;
	wire [4-1:0] node7198;
	wire [4-1:0] node7201;
	wire [4-1:0] node7202;
	wire [4-1:0] node7203;
	wire [4-1:0] node7206;
	wire [4-1:0] node7207;
	wire [4-1:0] node7208;
	wire [4-1:0] node7213;
	wire [4-1:0] node7214;
	wire [4-1:0] node7215;
	wire [4-1:0] node7218;
	wire [4-1:0] node7221;
	wire [4-1:0] node7224;
	wire [4-1:0] node7225;
	wire [4-1:0] node7226;
	wire [4-1:0] node7227;
	wire [4-1:0] node7228;
	wire [4-1:0] node7229;
	wire [4-1:0] node7232;
	wire [4-1:0] node7234;
	wire [4-1:0] node7235;
	wire [4-1:0] node7238;
	wire [4-1:0] node7241;
	wire [4-1:0] node7242;
	wire [4-1:0] node7244;
	wire [4-1:0] node7246;
	wire [4-1:0] node7249;
	wire [4-1:0] node7250;
	wire [4-1:0] node7251;
	wire [4-1:0] node7255;
	wire [4-1:0] node7256;
	wire [4-1:0] node7259;
	wire [4-1:0] node7262;
	wire [4-1:0] node7263;
	wire [4-1:0] node7264;
	wire [4-1:0] node7265;
	wire [4-1:0] node7266;
	wire [4-1:0] node7269;
	wire [4-1:0] node7272;
	wire [4-1:0] node7273;
	wire [4-1:0] node7276;
	wire [4-1:0] node7279;
	wire [4-1:0] node7280;
	wire [4-1:0] node7282;
	wire [4-1:0] node7284;
	wire [4-1:0] node7288;
	wire [4-1:0] node7289;
	wire [4-1:0] node7290;
	wire [4-1:0] node7291;
	wire [4-1:0] node7294;
	wire [4-1:0] node7298;
	wire [4-1:0] node7300;
	wire [4-1:0] node7303;
	wire [4-1:0] node7304;
	wire [4-1:0] node7305;
	wire [4-1:0] node7306;
	wire [4-1:0] node7307;
	wire [4-1:0] node7308;
	wire [4-1:0] node7312;
	wire [4-1:0] node7315;
	wire [4-1:0] node7317;
	wire [4-1:0] node7319;
	wire [4-1:0] node7322;
	wire [4-1:0] node7323;
	wire [4-1:0] node7324;
	wire [4-1:0] node7327;
	wire [4-1:0] node7328;
	wire [4-1:0] node7332;
	wire [4-1:0] node7333;
	wire [4-1:0] node7334;
	wire [4-1:0] node7335;
	wire [4-1:0] node7339;
	wire [4-1:0] node7342;
	wire [4-1:0] node7343;
	wire [4-1:0] node7344;
	wire [4-1:0] node7349;
	wire [4-1:0] node7350;
	wire [4-1:0] node7351;
	wire [4-1:0] node7352;
	wire [4-1:0] node7353;
	wire [4-1:0] node7357;
	wire [4-1:0] node7358;
	wire [4-1:0] node7359;
	wire [4-1:0] node7361;
	wire [4-1:0] node7366;
	wire [4-1:0] node7367;
	wire [4-1:0] node7369;
	wire [4-1:0] node7372;
	wire [4-1:0] node7373;
	wire [4-1:0] node7374;
	wire [4-1:0] node7377;
	wire [4-1:0] node7381;
	wire [4-1:0] node7382;
	wire [4-1:0] node7383;
	wire [4-1:0] node7386;
	wire [4-1:0] node7387;
	wire [4-1:0] node7388;
	wire [4-1:0] node7392;
	wire [4-1:0] node7396;
	wire [4-1:0] node7397;
	wire [4-1:0] node7398;
	wire [4-1:0] node7399;
	wire [4-1:0] node7400;
	wire [4-1:0] node7401;
	wire [4-1:0] node7404;
	wire [4-1:0] node7405;
	wire [4-1:0] node7406;
	wire [4-1:0] node7410;
	wire [4-1:0] node7413;
	wire [4-1:0] node7414;
	wire [4-1:0] node7416;
	wire [4-1:0] node7419;
	wire [4-1:0] node7421;
	wire [4-1:0] node7422;
	wire [4-1:0] node7425;
	wire [4-1:0] node7428;
	wire [4-1:0] node7429;
	wire [4-1:0] node7430;
	wire [4-1:0] node7432;
	wire [4-1:0] node7433;
	wire [4-1:0] node7437;
	wire [4-1:0] node7438;
	wire [4-1:0] node7441;
	wire [4-1:0] node7444;
	wire [4-1:0] node7445;
	wire [4-1:0] node7447;
	wire [4-1:0] node7448;
	wire [4-1:0] node7452;
	wire [4-1:0] node7453;
	wire [4-1:0] node7456;
	wire [4-1:0] node7459;
	wire [4-1:0] node7460;
	wire [4-1:0] node7461;
	wire [4-1:0] node7463;
	wire [4-1:0] node7464;
	wire [4-1:0] node7468;
	wire [4-1:0] node7469;
	wire [4-1:0] node7472;
	wire [4-1:0] node7475;
	wire [4-1:0] node7476;
	wire [4-1:0] node7479;
	wire [4-1:0] node7480;
	wire [4-1:0] node7484;
	wire [4-1:0] node7485;
	wire [4-1:0] node7486;
	wire [4-1:0] node7487;
	wire [4-1:0] node7488;
	wire [4-1:0] node7491;
	wire [4-1:0] node7494;
	wire [4-1:0] node7496;
	wire [4-1:0] node7498;
	wire [4-1:0] node7499;
	wire [4-1:0] node7502;
	wire [4-1:0] node7505;
	wire [4-1:0] node7506;
	wire [4-1:0] node7507;
	wire [4-1:0] node7508;
	wire [4-1:0] node7509;
	wire [4-1:0] node7515;
	wire [4-1:0] node7516;
	wire [4-1:0] node7519;
	wire [4-1:0] node7520;
	wire [4-1:0] node7522;
	wire [4-1:0] node7523;
	wire [4-1:0] node7526;
	wire [4-1:0] node7530;
	wire [4-1:0] node7531;
	wire [4-1:0] node7532;
	wire [4-1:0] node7533;
	wire [4-1:0] node7535;
	wire [4-1:0] node7539;
	wire [4-1:0] node7543;
	wire [4-1:0] node7545;
	wire [4-1:0] node7546;
	wire [4-1:0] node7548;
	wire [4-1:0] node7549;
	wire [4-1:0] node7550;
	wire [4-1:0] node7551;
	wire [4-1:0] node7552;
	wire [4-1:0] node7553;
	wire [4-1:0] node7554;
	wire [4-1:0] node7558;
	wire [4-1:0] node7560;
	wire [4-1:0] node7563;
	wire [4-1:0] node7564;
	wire [4-1:0] node7568;
	wire [4-1:0] node7570;
	wire [4-1:0] node7571;
	wire [4-1:0] node7573;
	wire [4-1:0] node7577;
	wire [4-1:0] node7578;
	wire [4-1:0] node7579;
	wire [4-1:0] node7581;
	wire [4-1:0] node7582;
	wire [4-1:0] node7585;
	wire [4-1:0] node7588;
	wire [4-1:0] node7590;
	wire [4-1:0] node7592;
	wire [4-1:0] node7595;
	wire [4-1:0] node7596;
	wire [4-1:0] node7597;
	wire [4-1:0] node7598;
	wire [4-1:0] node7602;
	wire [4-1:0] node7605;
	wire [4-1:0] node7609;
	wire [4-1:0] node7610;
	wire [4-1:0] node7611;
	wire [4-1:0] node7612;
	wire [4-1:0] node7613;
	wire [4-1:0] node7614;
	wire [4-1:0] node7616;
	wire [4-1:0] node7619;
	wire [4-1:0] node7620;
	wire [4-1:0] node7623;
	wire [4-1:0] node7624;
	wire [4-1:0] node7625;
	wire [4-1:0] node7630;
	wire [4-1:0] node7631;
	wire [4-1:0] node7632;
	wire [4-1:0] node7634;
	wire [4-1:0] node7637;
	wire [4-1:0] node7640;
	wire [4-1:0] node7641;
	wire [4-1:0] node7643;
	wire [4-1:0] node7644;
	wire [4-1:0] node7649;
	wire [4-1:0] node7650;
	wire [4-1:0] node7651;
	wire [4-1:0] node7652;
	wire [4-1:0] node7653;
	wire [4-1:0] node7656;
	wire [4-1:0] node7660;
	wire [4-1:0] node7661;
	wire [4-1:0] node7662;
	wire [4-1:0] node7666;
	wire [4-1:0] node7668;
	wire [4-1:0] node7671;
	wire [4-1:0] node7672;
	wire [4-1:0] node7673;
	wire [4-1:0] node7674;
	wire [4-1:0] node7678;
	wire [4-1:0] node7681;
	wire [4-1:0] node7682;
	wire [4-1:0] node7683;
	wire [4-1:0] node7687;
	wire [4-1:0] node7688;
	wire [4-1:0] node7692;
	wire [4-1:0] node7693;
	wire [4-1:0] node7694;
	wire [4-1:0] node7695;
	wire [4-1:0] node7696;
	wire [4-1:0] node7697;
	wire [4-1:0] node7702;
	wire [4-1:0] node7703;
	wire [4-1:0] node7704;
	wire [4-1:0] node7705;
	wire [4-1:0] node7710;
	wire [4-1:0] node7713;
	wire [4-1:0] node7714;
	wire [4-1:0] node7716;
	wire [4-1:0] node7717;
	wire [4-1:0] node7721;
	wire [4-1:0] node7722;
	wire [4-1:0] node7723;
	wire [4-1:0] node7724;
	wire [4-1:0] node7728;
	wire [4-1:0] node7731;
	wire [4-1:0] node7734;
	wire [4-1:0] node7735;
	wire [4-1:0] node7736;
	wire [4-1:0] node7737;
	wire [4-1:0] node7738;
	wire [4-1:0] node7742;
	wire [4-1:0] node7743;
	wire [4-1:0] node7747;
	wire [4-1:0] node7748;
	wire [4-1:0] node7751;
	wire [4-1:0] node7752;
	wire [4-1:0] node7756;
	wire [4-1:0] node7757;
	wire [4-1:0] node7758;
	wire [4-1:0] node7759;
	wire [4-1:0] node7760;
	wire [4-1:0] node7762;
	wire [4-1:0] node7765;
	wire [4-1:0] node7771;
	wire [4-1:0] node7773;
	wire [4-1:0] node7774;
	wire [4-1:0] node7775;
	wire [4-1:0] node7776;
	wire [4-1:0] node7777;
	wire [4-1:0] node7779;
	wire [4-1:0] node7782;
	wire [4-1:0] node7785;
	wire [4-1:0] node7786;
	wire [4-1:0] node7787;
	wire [4-1:0] node7789;
	wire [4-1:0] node7792;
	wire [4-1:0] node7796;
	wire [4-1:0] node7797;
	wire [4-1:0] node7798;
	wire [4-1:0] node7799;
	wire [4-1:0] node7800;
	wire [4-1:0] node7804;
	wire [4-1:0] node7807;
	wire [4-1:0] node7809;
	wire [4-1:0] node7812;
	wire [4-1:0] node7813;
	wire [4-1:0] node7817;
	wire [4-1:0] node7819;
	wire [4-1:0] node7820;
	wire [4-1:0] node7822;
	wire [4-1:0] node7823;
	wire [4-1:0] node7827;
	wire [4-1:0] node7828;
	wire [4-1:0] node7832;
	wire [4-1:0] node7833;
	wire [4-1:0] node7834;
	wire [4-1:0] node7835;
	wire [4-1:0] node7836;
	wire [4-1:0] node7837;
	wire [4-1:0] node7838;
	wire [4-1:0] node7839;
	wire [4-1:0] node7840;
	wire [4-1:0] node7842;
	wire [4-1:0] node7845;
	wire [4-1:0] node7846;
	wire [4-1:0] node7847;
	wire [4-1:0] node7849;
	wire [4-1:0] node7852;
	wire [4-1:0] node7853;
	wire [4-1:0] node7857;
	wire [4-1:0] node7858;
	wire [4-1:0] node7860;
	wire [4-1:0] node7863;
	wire [4-1:0] node7866;
	wire [4-1:0] node7868;
	wire [4-1:0] node7870;
	wire [4-1:0] node7872;
	wire [4-1:0] node7873;
	wire [4-1:0] node7877;
	wire [4-1:0] node7878;
	wire [4-1:0] node7879;
	wire [4-1:0] node7880;
	wire [4-1:0] node7883;
	wire [4-1:0] node7886;
	wire [4-1:0] node7887;
	wire [4-1:0] node7888;
	wire [4-1:0] node7892;
	wire [4-1:0] node7893;
	wire [4-1:0] node7894;
	wire [4-1:0] node7897;
	wire [4-1:0] node7900;
	wire [4-1:0] node7902;
	wire [4-1:0] node7903;
	wire [4-1:0] node7907;
	wire [4-1:0] node7908;
	wire [4-1:0] node7909;
	wire [4-1:0] node7910;
	wire [4-1:0] node7914;
	wire [4-1:0] node7916;
	wire [4-1:0] node7917;
	wire [4-1:0] node7919;
	wire [4-1:0] node7922;
	wire [4-1:0] node7925;
	wire [4-1:0] node7926;
	wire [4-1:0] node7928;
	wire [4-1:0] node7929;
	wire [4-1:0] node7930;
	wire [4-1:0] node7933;
	wire [4-1:0] node7937;
	wire [4-1:0] node7938;
	wire [4-1:0] node7939;
	wire [4-1:0] node7943;
	wire [4-1:0] node7944;
	wire [4-1:0] node7949;
	wire [4-1:0] node7950;
	wire [4-1:0] node7951;
	wire [4-1:0] node7952;
	wire [4-1:0] node7953;
	wire [4-1:0] node7954;
	wire [4-1:0] node7955;
	wire [4-1:0] node7957;
	wire [4-1:0] node7959;
	wire [4-1:0] node7960;
	wire [4-1:0] node7964;
	wire [4-1:0] node7966;
	wire [4-1:0] node7969;
	wire [4-1:0] node7970;
	wire [4-1:0] node7972;
	wire [4-1:0] node7975;
	wire [4-1:0] node7976;
	wire [4-1:0] node7980;
	wire [4-1:0] node7981;
	wire [4-1:0] node7982;
	wire [4-1:0] node7983;
	wire [4-1:0] node7986;
	wire [4-1:0] node7990;
	wire [4-1:0] node7991;
	wire [4-1:0] node7994;
	wire [4-1:0] node7995;
	wire [4-1:0] node7998;
	wire [4-1:0] node8001;
	wire [4-1:0] node8002;
	wire [4-1:0] node8003;
	wire [4-1:0] node8004;
	wire [4-1:0] node8007;
	wire [4-1:0] node8011;
	wire [4-1:0] node8012;
	wire [4-1:0] node8013;
	wire [4-1:0] node8016;
	wire [4-1:0] node8019;
	wire [4-1:0] node8020;
	wire [4-1:0] node8021;
	wire [4-1:0] node8025;
	wire [4-1:0] node8028;
	wire [4-1:0] node8029;
	wire [4-1:0] node8030;
	wire [4-1:0] node8031;
	wire [4-1:0] node8034;
	wire [4-1:0] node8035;
	wire [4-1:0] node8036;
	wire [4-1:0] node8039;
	wire [4-1:0] node8043;
	wire [4-1:0] node8045;
	wire [4-1:0] node8046;
	wire [4-1:0] node8049;
	wire [4-1:0] node8052;
	wire [4-1:0] node8053;
	wire [4-1:0] node8054;
	wire [4-1:0] node8056;
	wire [4-1:0] node8059;
	wire [4-1:0] node8060;
	wire [4-1:0] node8061;
	wire [4-1:0] node8065;
	wire [4-1:0] node8067;
	wire [4-1:0] node8070;
	wire [4-1:0] node8071;
	wire [4-1:0] node8072;
	wire [4-1:0] node8073;
	wire [4-1:0] node8078;
	wire [4-1:0] node8079;
	wire [4-1:0] node8080;
	wire [4-1:0] node8084;
	wire [4-1:0] node8087;
	wire [4-1:0] node8088;
	wire [4-1:0] node8089;
	wire [4-1:0] node8090;
	wire [4-1:0] node8091;
	wire [4-1:0] node8093;
	wire [4-1:0] node8094;
	wire [4-1:0] node8097;
	wire [4-1:0] node8100;
	wire [4-1:0] node8101;
	wire [4-1:0] node8102;
	wire [4-1:0] node8107;
	wire [4-1:0] node8108;
	wire [4-1:0] node8109;
	wire [4-1:0] node8110;
	wire [4-1:0] node8111;
	wire [4-1:0] node8114;
	wire [4-1:0] node8118;
	wire [4-1:0] node8119;
	wire [4-1:0] node8123;
	wire [4-1:0] node8125;
	wire [4-1:0] node8126;
	wire [4-1:0] node8129;
	wire [4-1:0] node8132;
	wire [4-1:0] node8133;
	wire [4-1:0] node8134;
	wire [4-1:0] node8135;
	wire [4-1:0] node8139;
	wire [4-1:0] node8140;
	wire [4-1:0] node8143;
	wire [4-1:0] node8146;
	wire [4-1:0] node8147;
	wire [4-1:0] node8150;
	wire [4-1:0] node8151;
	wire [4-1:0] node8152;
	wire [4-1:0] node8156;
	wire [4-1:0] node8157;
	wire [4-1:0] node8158;
	wire [4-1:0] node8163;
	wire [4-1:0] node8164;
	wire [4-1:0] node8165;
	wire [4-1:0] node8166;
	wire [4-1:0] node8167;
	wire [4-1:0] node8168;
	wire [4-1:0] node8172;
	wire [4-1:0] node8173;
	wire [4-1:0] node8178;
	wire [4-1:0] node8179;
	wire [4-1:0] node8181;
	wire [4-1:0] node8183;
	wire [4-1:0] node8187;
	wire [4-1:0] node8188;
	wire [4-1:0] node8189;
	wire [4-1:0] node8192;
	wire [4-1:0] node8194;
	wire [4-1:0] node8197;
	wire [4-1:0] node8199;
	wire [4-1:0] node8200;
	wire [4-1:0] node8203;
	wire [4-1:0] node8207;
	wire [4-1:0] node8208;
	wire [4-1:0] node8209;
	wire [4-1:0] node8210;
	wire [4-1:0] node8211;
	wire [4-1:0] node8212;
	wire [4-1:0] node8213;
	wire [4-1:0] node8214;
	wire [4-1:0] node8215;
	wire [4-1:0] node8219;
	wire [4-1:0] node8220;
	wire [4-1:0] node8221;
	wire [4-1:0] node8224;
	wire [4-1:0] node8225;
	wire [4-1:0] node8229;
	wire [4-1:0] node8231;
	wire [4-1:0] node8232;
	wire [4-1:0] node8236;
	wire [4-1:0] node8237;
	wire [4-1:0] node8238;
	wire [4-1:0] node8239;
	wire [4-1:0] node8242;
	wire [4-1:0] node8245;
	wire [4-1:0] node8247;
	wire [4-1:0] node8249;
	wire [4-1:0] node8252;
	wire [4-1:0] node8253;
	wire [4-1:0] node8255;
	wire [4-1:0] node8257;
	wire [4-1:0] node8260;
	wire [4-1:0] node8263;
	wire [4-1:0] node8264;
	wire [4-1:0] node8265;
	wire [4-1:0] node8267;
	wire [4-1:0] node8271;
	wire [4-1:0] node8272;
	wire [4-1:0] node8273;
	wire [4-1:0] node8277;
	wire [4-1:0] node8279;
	wire [4-1:0] node8282;
	wire [4-1:0] node8283;
	wire [4-1:0] node8284;
	wire [4-1:0] node8285;
	wire [4-1:0] node8286;
	wire [4-1:0] node8287;
	wire [4-1:0] node8292;
	wire [4-1:0] node8293;
	wire [4-1:0] node8297;
	wire [4-1:0] node8298;
	wire [4-1:0] node8299;
	wire [4-1:0] node8300;
	wire [4-1:0] node8303;
	wire [4-1:0] node8305;
	wire [4-1:0] node8308;
	wire [4-1:0] node8309;
	wire [4-1:0] node8311;
	wire [4-1:0] node8312;
	wire [4-1:0] node8317;
	wire [4-1:0] node8318;
	wire [4-1:0] node8320;
	wire [4-1:0] node8321;
	wire [4-1:0] node8322;
	wire [4-1:0] node8328;
	wire [4-1:0] node8329;
	wire [4-1:0] node8330;
	wire [4-1:0] node8331;
	wire [4-1:0] node8332;
	wire [4-1:0] node8336;
	wire [4-1:0] node8337;
	wire [4-1:0] node8339;
	wire [4-1:0] node8343;
	wire [4-1:0] node8345;
	wire [4-1:0] node8346;
	wire [4-1:0] node8350;
	wire [4-1:0] node8351;
	wire [4-1:0] node8352;
	wire [4-1:0] node8353;
	wire [4-1:0] node8357;
	wire [4-1:0] node8359;
	wire [4-1:0] node8362;
	wire [4-1:0] node8364;
	wire [4-1:0] node8365;
	wire [4-1:0] node8367;
	wire [4-1:0] node8371;
	wire [4-1:0] node8372;
	wire [4-1:0] node8373;
	wire [4-1:0] node8374;
	wire [4-1:0] node8376;
	wire [4-1:0] node8377;
	wire [4-1:0] node8378;
	wire [4-1:0] node8381;
	wire [4-1:0] node8385;
	wire [4-1:0] node8386;
	wire [4-1:0] node8387;
	wire [4-1:0] node8388;
	wire [4-1:0] node8391;
	wire [4-1:0] node8392;
	wire [4-1:0] node8397;
	wire [4-1:0] node8398;
	wire [4-1:0] node8399;
	wire [4-1:0] node8402;
	wire [4-1:0] node8406;
	wire [4-1:0] node8407;
	wire [4-1:0] node8408;
	wire [4-1:0] node8409;
	wire [4-1:0] node8412;
	wire [4-1:0] node8414;
	wire [4-1:0] node8417;
	wire [4-1:0] node8419;
	wire [4-1:0] node8420;
	wire [4-1:0] node8423;
	wire [4-1:0] node8426;
	wire [4-1:0] node8427;
	wire [4-1:0] node8429;
	wire [4-1:0] node8430;
	wire [4-1:0] node8434;
	wire [4-1:0] node8435;
	wire [4-1:0] node8438;
	wire [4-1:0] node8441;
	wire [4-1:0] node8442;
	wire [4-1:0] node8443;
	wire [4-1:0] node8444;
	wire [4-1:0] node8445;
	wire [4-1:0] node8449;
	wire [4-1:0] node8450;
	wire [4-1:0] node8451;
	wire [4-1:0] node8455;
	wire [4-1:0] node8458;
	wire [4-1:0] node8459;
	wire [4-1:0] node8460;
	wire [4-1:0] node8463;
	wire [4-1:0] node8464;
	wire [4-1:0] node8468;
	wire [4-1:0] node8469;
	wire [4-1:0] node8471;
	wire [4-1:0] node8474;
	wire [4-1:0] node8476;
	wire [4-1:0] node8477;
	wire [4-1:0] node8480;
	wire [4-1:0] node8483;
	wire [4-1:0] node8484;
	wire [4-1:0] node8485;
	wire [4-1:0] node8486;
	wire [4-1:0] node8488;
	wire [4-1:0] node8492;
	wire [4-1:0] node8494;
	wire [4-1:0] node8497;
	wire [4-1:0] node8499;
	wire [4-1:0] node8502;
	wire [4-1:0] node8503;
	wire [4-1:0] node8504;
	wire [4-1:0] node8505;
	wire [4-1:0] node8507;
	wire [4-1:0] node8508;
	wire [4-1:0] node8509;
	wire [4-1:0] node8511;
	wire [4-1:0] node8516;
	wire [4-1:0] node8517;
	wire [4-1:0] node8518;
	wire [4-1:0] node8519;
	wire [4-1:0] node8520;
	wire [4-1:0] node8521;
	wire [4-1:0] node8525;
	wire [4-1:0] node8528;
	wire [4-1:0] node8530;
	wire [4-1:0] node8533;
	wire [4-1:0] node8534;
	wire [4-1:0] node8537;
	wire [4-1:0] node8540;
	wire [4-1:0] node8542;
	wire [4-1:0] node8544;
	wire [4-1:0] node8547;
	wire [4-1:0] node8548;
	wire [4-1:0] node8549;
	wire [4-1:0] node8550;
	wire [4-1:0] node8552;
	wire [4-1:0] node8553;
	wire [4-1:0] node8556;
	wire [4-1:0] node8558;
	wire [4-1:0] node8561;
	wire [4-1:0] node8562;
	wire [4-1:0] node8563;
	wire [4-1:0] node8567;
	wire [4-1:0] node8570;
	wire [4-1:0] node8571;
	wire [4-1:0] node8572;
	wire [4-1:0] node8576;
	wire [4-1:0] node8577;
	wire [4-1:0] node8578;
	wire [4-1:0] node8579;
	wire [4-1:0] node8584;
	wire [4-1:0] node8586;
	wire [4-1:0] node8587;
	wire [4-1:0] node8590;
	wire [4-1:0] node8593;
	wire [4-1:0] node8594;
	wire [4-1:0] node8595;
	wire [4-1:0] node8596;
	wire [4-1:0] node8597;
	wire [4-1:0] node8601;
	wire [4-1:0] node8603;
	wire [4-1:0] node8606;
	wire [4-1:0] node8607;
	wire [4-1:0] node8610;
	wire [4-1:0] node8612;
	wire [4-1:0] node8615;
	wire [4-1:0] node8616;
	wire [4-1:0] node8617;
	wire [4-1:0] node8618;
	wire [4-1:0] node8622;
	wire [4-1:0] node8625;
	wire [4-1:0] node8627;
	wire [4-1:0] node8631;
	wire [4-1:0] node8632;
	wire [4-1:0] node8633;
	wire [4-1:0] node8634;
	wire [4-1:0] node8635;
	wire [4-1:0] node8636;
	wire [4-1:0] node8637;
	wire [4-1:0] node8638;
	wire [4-1:0] node8640;
	wire [4-1:0] node8641;
	wire [4-1:0] node8645;
	wire [4-1:0] node8646;
	wire [4-1:0] node8650;
	wire [4-1:0] node8652;
	wire [4-1:0] node8653;
	wire [4-1:0] node8656;
	wire [4-1:0] node8658;
	wire [4-1:0] node8661;
	wire [4-1:0] node8662;
	wire [4-1:0] node8663;
	wire [4-1:0] node8664;
	wire [4-1:0] node8667;
	wire [4-1:0] node8671;
	wire [4-1:0] node8672;
	wire [4-1:0] node8673;
	wire [4-1:0] node8678;
	wire [4-1:0] node8679;
	wire [4-1:0] node8680;
	wire [4-1:0] node8682;
	wire [4-1:0] node8685;
	wire [4-1:0] node8686;
	wire [4-1:0] node8687;
	wire [4-1:0] node8689;
	wire [4-1:0] node8693;
	wire [4-1:0] node8696;
	wire [4-1:0] node8697;
	wire [4-1:0] node8698;
	wire [4-1:0] node8699;
	wire [4-1:0] node8700;
	wire [4-1:0] node8702;
	wire [4-1:0] node8705;
	wire [4-1:0] node8708;
	wire [4-1:0] node8710;
	wire [4-1:0] node8713;
	wire [4-1:0] node8714;
	wire [4-1:0] node8718;
	wire [4-1:0] node8719;
	wire [4-1:0] node8721;
	wire [4-1:0] node8722;
	wire [4-1:0] node8726;
	wire [4-1:0] node8728;
	wire [4-1:0] node8730;
	wire [4-1:0] node8733;
	wire [4-1:0] node8734;
	wire [4-1:0] node8735;
	wire [4-1:0] node8736;
	wire [4-1:0] node8737;
	wire [4-1:0] node8738;
	wire [4-1:0] node8742;
	wire [4-1:0] node8743;
	wire [4-1:0] node8745;
	wire [4-1:0] node8749;
	wire [4-1:0] node8750;
	wire [4-1:0] node8751;
	wire [4-1:0] node8752;
	wire [4-1:0] node8754;
	wire [4-1:0] node8758;
	wire [4-1:0] node8762;
	wire [4-1:0] node8763;
	wire [4-1:0] node8765;
	wire [4-1:0] node8768;
	wire [4-1:0] node8770;
	wire [4-1:0] node8772;
	wire [4-1:0] node8775;
	wire [4-1:0] node8776;
	wire [4-1:0] node8778;
	wire [4-1:0] node8779;
	wire [4-1:0] node8781;
	wire [4-1:0] node8784;
	wire [4-1:0] node8786;
	wire [4-1:0] node8790;
	wire [4-1:0] node8791;
	wire [4-1:0] node8792;
	wire [4-1:0] node8793;
	wire [4-1:0] node8794;
	wire [4-1:0] node8795;
	wire [4-1:0] node8796;
	wire [4-1:0] node8799;
	wire [4-1:0] node8802;
	wire [4-1:0] node8805;
	wire [4-1:0] node8806;
	wire [4-1:0] node8807;
	wire [4-1:0] node8808;
	wire [4-1:0] node8809;
	wire [4-1:0] node8814;
	wire [4-1:0] node8815;
	wire [4-1:0] node8819;
	wire [4-1:0] node8822;
	wire [4-1:0] node8823;
	wire [4-1:0] node8824;
	wire [4-1:0] node8825;
	wire [4-1:0] node8826;
	wire [4-1:0] node8831;
	wire [4-1:0] node8833;
	wire [4-1:0] node8836;
	wire [4-1:0] node8837;
	wire [4-1:0] node8839;
	wire [4-1:0] node8842;
	wire [4-1:0] node8843;
	wire [4-1:0] node8847;
	wire [4-1:0] node8848;
	wire [4-1:0] node8849;
	wire [4-1:0] node8851;
	wire [4-1:0] node8852;
	wire [4-1:0] node8853;
	wire [4-1:0] node8858;
	wire [4-1:0] node8859;
	wire [4-1:0] node8860;
	wire [4-1:0] node8863;
	wire [4-1:0] node8864;
	wire [4-1:0] node8869;
	wire [4-1:0] node8870;
	wire [4-1:0] node8871;
	wire [4-1:0] node8873;
	wire [4-1:0] node8877;
	wire [4-1:0] node8878;
	wire [4-1:0] node8879;
	wire [4-1:0] node8883;
	wire [4-1:0] node8884;
	wire [4-1:0] node8888;
	wire [4-1:0] node8889;
	wire [4-1:0] node8890;
	wire [4-1:0] node8891;
	wire [4-1:0] node8892;
	wire [4-1:0] node8893;
	wire [4-1:0] node8896;
	wire [4-1:0] node8898;
	wire [4-1:0] node8901;
	wire [4-1:0] node8902;
	wire [4-1:0] node8905;
	wire [4-1:0] node8908;
	wire [4-1:0] node8910;
	wire [4-1:0] node8913;
	wire [4-1:0] node8914;
	wire [4-1:0] node8915;
	wire [4-1:0] node8916;
	wire [4-1:0] node8921;
	wire [4-1:0] node8924;
	wire [4-1:0] node8925;
	wire [4-1:0] node8926;
	wire [4-1:0] node8927;
	wire [4-1:0] node8929;
	wire [4-1:0] node8931;
	wire [4-1:0] node8934;
	wire [4-1:0] node8937;
	wire [4-1:0] node8939;
	wire [4-1:0] node8940;
	wire [4-1:0] node8943;
	wire [4-1:0] node8946;
	wire [4-1:0] node8948;
	wire [4-1:0] node8949;
	wire [4-1:0] node8951;
	wire [4-1:0] node8954;
	wire [4-1:0] node8957;
	wire [4-1:0] node8958;
	wire [4-1:0] node8959;
	wire [4-1:0] node8960;
	wire [4-1:0] node8961;
	wire [4-1:0] node8962;
	wire [4-1:0] node8963;
	wire [4-1:0] node8964;
	wire [4-1:0] node8967;
	wire [4-1:0] node8969;
	wire [4-1:0] node8971;
	wire [4-1:0] node8975;
	wire [4-1:0] node8977;
	wire [4-1:0] node8980;
	wire [4-1:0] node8981;
	wire [4-1:0] node8982;
	wire [4-1:0] node8984;
	wire [4-1:0] node8985;
	wire [4-1:0] node8990;
	wire [4-1:0] node8991;
	wire [4-1:0] node8994;
	wire [4-1:0] node8996;
	wire [4-1:0] node8999;
	wire [4-1:0] node9000;
	wire [4-1:0] node9001;
	wire [4-1:0] node9002;
	wire [4-1:0] node9005;
	wire [4-1:0] node9006;
	wire [4-1:0] node9008;
	wire [4-1:0] node9010;
	wire [4-1:0] node9014;
	wire [4-1:0] node9016;
	wire [4-1:0] node9019;
	wire [4-1:0] node9020;
	wire [4-1:0] node9021;
	wire [4-1:0] node9024;
	wire [4-1:0] node9025;
	wire [4-1:0] node9029;
	wire [4-1:0] node9031;
	wire [4-1:0] node9032;
	wire [4-1:0] node9033;
	wire [4-1:0] node9038;
	wire [4-1:0] node9039;
	wire [4-1:0] node9040;
	wire [4-1:0] node9041;
	wire [4-1:0] node9042;
	wire [4-1:0] node9045;
	wire [4-1:0] node9046;
	wire [4-1:0] node9050;
	wire [4-1:0] node9051;
	wire [4-1:0] node9052;
	wire [4-1:0] node9056;
	wire [4-1:0] node9058;
	wire [4-1:0] node9060;
	wire [4-1:0] node9063;
	wire [4-1:0] node9064;
	wire [4-1:0] node9065;
	wire [4-1:0] node9069;
	wire [4-1:0] node9070;
	wire [4-1:0] node9071;
	wire [4-1:0] node9073;
	wire [4-1:0] node9077;
	wire [4-1:0] node9078;
	wire [4-1:0] node9080;
	wire [4-1:0] node9083;
	wire [4-1:0] node9086;
	wire [4-1:0] node9087;
	wire [4-1:0] node9088;
	wire [4-1:0] node9089;
	wire [4-1:0] node9090;
	wire [4-1:0] node9092;
	wire [4-1:0] node9095;
	wire [4-1:0] node9099;
	wire [4-1:0] node9102;
	wire [4-1:0] node9103;
	wire [4-1:0] node9104;
	wire [4-1:0] node9106;
	wire [4-1:0] node9111;
	wire [4-1:0] node9112;
	wire [4-1:0] node9113;
	wire [4-1:0] node9114;
	wire [4-1:0] node9115;
	wire [4-1:0] node9117;
	wire [4-1:0] node9118;
	wire [4-1:0] node9122;
	wire [4-1:0] node9123;
	wire [4-1:0] node9125;
	wire [4-1:0] node9128;
	wire [4-1:0] node9131;
	wire [4-1:0] node9132;
	wire [4-1:0] node9133;
	wire [4-1:0] node9134;
	wire [4-1:0] node9135;
	wire [4-1:0] node9141;
	wire [4-1:0] node9142;
	wire [4-1:0] node9144;
	wire [4-1:0] node9147;
	wire [4-1:0] node9148;
	wire [4-1:0] node9151;
	wire [4-1:0] node9152;
	wire [4-1:0] node9154;
	wire [4-1:0] node9158;
	wire [4-1:0] node9159;
	wire [4-1:0] node9160;
	wire [4-1:0] node9163;
	wire [4-1:0] node9164;
	wire [4-1:0] node9165;
	wire [4-1:0] node9168;
	wire [4-1:0] node9170;
	wire [4-1:0] node9173;
	wire [4-1:0] node9174;
	wire [4-1:0] node9177;
	wire [4-1:0] node9181;
	wire [4-1:0] node9182;
	wire [4-1:0] node9183;
	wire [4-1:0] node9184;
	wire [4-1:0] node9186;
	wire [4-1:0] node9188;
	wire [4-1:0] node9191;
	wire [4-1:0] node9192;
	wire [4-1:0] node9193;
	wire [4-1:0] node9197;
	wire [4-1:0] node9198;
	wire [4-1:0] node9202;
	wire [4-1:0] node9203;
	wire [4-1:0] node9206;
	wire [4-1:0] node9207;
	wire [4-1:0] node9208;
	wire [4-1:0] node9211;
	wire [4-1:0] node9212;
	wire [4-1:0] node9216;
	wire [4-1:0] node9218;
	wire [4-1:0] node9221;
	wire [4-1:0] node9222;
	wire [4-1:0] node9223;
	wire [4-1:0] node9224;
	wire [4-1:0] node9227;
	wire [4-1:0] node9229;
	wire [4-1:0] node9234;
	wire [4-1:0] node9235;
	wire [4-1:0] node9236;
	wire [4-1:0] node9237;
	wire [4-1:0] node9238;
	wire [4-1:0] node9240;
	wire [4-1:0] node9241;
	wire [4-1:0] node9243;
	wire [4-1:0] node9245;
	wire [4-1:0] node9247;
	wire [4-1:0] node9250;
	wire [4-1:0] node9251;
	wire [4-1:0] node9252;
	wire [4-1:0] node9254;
	wire [4-1:0] node9257;
	wire [4-1:0] node9258;
	wire [4-1:0] node9259;
	wire [4-1:0] node9262;
	wire [4-1:0] node9265;
	wire [4-1:0] node9267;
	wire [4-1:0] node9270;
	wire [4-1:0] node9272;
	wire [4-1:0] node9275;
	wire [4-1:0] node9276;
	wire [4-1:0] node9277;
	wire [4-1:0] node9278;
	wire [4-1:0] node9279;
	wire [4-1:0] node9280;
	wire [4-1:0] node9282;
	wire [4-1:0] node9284;
	wire [4-1:0] node9288;
	wire [4-1:0] node9289;
	wire [4-1:0] node9290;
	wire [4-1:0] node9294;
	wire [4-1:0] node9295;
	wire [4-1:0] node9299;
	wire [4-1:0] node9300;
	wire [4-1:0] node9301;
	wire [4-1:0] node9302;
	wire [4-1:0] node9306;
	wire [4-1:0] node9308;
	wire [4-1:0] node9309;
	wire [4-1:0] node9312;
	wire [4-1:0] node9315;
	wire [4-1:0] node9316;
	wire [4-1:0] node9319;
	wire [4-1:0] node9320;
	wire [4-1:0] node9324;
	wire [4-1:0] node9325;
	wire [4-1:0] node9327;
	wire [4-1:0] node9328;
	wire [4-1:0] node9329;
	wire [4-1:0] node9333;
	wire [4-1:0] node9336;
	wire [4-1:0] node9337;
	wire [4-1:0] node9338;
	wire [4-1:0] node9341;
	wire [4-1:0] node9344;
	wire [4-1:0] node9345;
	wire [4-1:0] node9349;
	wire [4-1:0] node9350;
	wire [4-1:0] node9351;
	wire [4-1:0] node9352;
	wire [4-1:0] node9353;
	wire [4-1:0] node9357;
	wire [4-1:0] node9358;
	wire [4-1:0] node9361;
	wire [4-1:0] node9362;
	wire [4-1:0] node9364;
	wire [4-1:0] node9365;
	wire [4-1:0] node9368;
	wire [4-1:0] node9372;
	wire [4-1:0] node9373;
	wire [4-1:0] node9374;
	wire [4-1:0] node9377;
	wire [4-1:0] node9379;
	wire [4-1:0] node9382;
	wire [4-1:0] node9384;
	wire [4-1:0] node9385;
	wire [4-1:0] node9389;
	wire [4-1:0] node9390;
	wire [4-1:0] node9391;
	wire [4-1:0] node9394;
	wire [4-1:0] node9396;
	wire [4-1:0] node9397;
	wire [4-1:0] node9398;
	wire [4-1:0] node9402;
	wire [4-1:0] node9405;
	wire [4-1:0] node9406;
	wire [4-1:0] node9408;
	wire [4-1:0] node9409;
	wire [4-1:0] node9413;
	wire [4-1:0] node9414;
	wire [4-1:0] node9416;
	wire [4-1:0] node9417;
	wire [4-1:0] node9418;
	wire [4-1:0] node9421;
	wire [4-1:0] node9425;
	wire [4-1:0] node9427;
	wire [4-1:0] node9430;
	wire [4-1:0] node9432;
	wire [4-1:0] node9434;
	wire [4-1:0] node9435;
	wire [4-1:0] node9437;
	wire [4-1:0] node9438;
	wire [4-1:0] node9439;
	wire [4-1:0] node9442;
	wire [4-1:0] node9444;
	wire [4-1:0] node9446;
	wire [4-1:0] node9450;
	wire [4-1:0] node9451;
	wire [4-1:0] node9452;
	wire [4-1:0] node9453;
	wire [4-1:0] node9455;
	wire [4-1:0] node9456;
	wire [4-1:0] node9461;
	wire [4-1:0] node9462;
	wire [4-1:0] node9464;
	wire [4-1:0] node9465;
	wire [4-1:0] node9469;
	wire [4-1:0] node9472;
	wire [4-1:0] node9473;
	wire [4-1:0] node9475;
	wire [4-1:0] node9477;
	wire [4-1:0] node9481;
	wire [4-1:0] node9482;
	wire [4-1:0] node9483;
	wire [4-1:0] node9484;
	wire [4-1:0] node9485;
	wire [4-1:0] node9486;
	wire [4-1:0] node9487;
	wire [4-1:0] node9488;
	wire [4-1:0] node9489;
	wire [4-1:0] node9491;
	wire [4-1:0] node9494;
	wire [4-1:0] node9499;
	wire [4-1:0] node9500;
	wire [4-1:0] node9502;
	wire [4-1:0] node9506;
	wire [4-1:0] node9507;
	wire [4-1:0] node9508;
	wire [4-1:0] node9510;
	wire [4-1:0] node9513;
	wire [4-1:0] node9514;
	wire [4-1:0] node9516;
	wire [4-1:0] node9519;
	wire [4-1:0] node9520;
	wire [4-1:0] node9523;
	wire [4-1:0] node9524;
	wire [4-1:0] node9528;
	wire [4-1:0] node9529;
	wire [4-1:0] node9530;
	wire [4-1:0] node9532;
	wire [4-1:0] node9535;
	wire [4-1:0] node9537;
	wire [4-1:0] node9538;
	wire [4-1:0] node9542;
	wire [4-1:0] node9544;
	wire [4-1:0] node9546;
	wire [4-1:0] node9549;
	wire [4-1:0] node9550;
	wire [4-1:0] node9551;
	wire [4-1:0] node9552;
	wire [4-1:0] node9553;
	wire [4-1:0] node9556;
	wire [4-1:0] node9558;
	wire [4-1:0] node9561;
	wire [4-1:0] node9562;
	wire [4-1:0] node9564;
	wire [4-1:0] node9567;
	wire [4-1:0] node9570;
	wire [4-1:0] node9571;
	wire [4-1:0] node9572;
	wire [4-1:0] node9575;
	wire [4-1:0] node9576;
	wire [4-1:0] node9578;
	wire [4-1:0] node9581;
	wire [4-1:0] node9582;
	wire [4-1:0] node9586;
	wire [4-1:0] node9587;
	wire [4-1:0] node9588;
	wire [4-1:0] node9592;
	wire [4-1:0] node9595;
	wire [4-1:0] node9596;
	wire [4-1:0] node9597;
	wire [4-1:0] node9598;
	wire [4-1:0] node9601;
	wire [4-1:0] node9602;
	wire [4-1:0] node9606;
	wire [4-1:0] node9607;
	wire [4-1:0] node9608;
	wire [4-1:0] node9612;
	wire [4-1:0] node9613;
	wire [4-1:0] node9617;
	wire [4-1:0] node9618;
	wire [4-1:0] node9620;
	wire [4-1:0] node9621;
	wire [4-1:0] node9625;
	wire [4-1:0] node9628;
	wire [4-1:0] node9629;
	wire [4-1:0] node9630;
	wire [4-1:0] node9631;
	wire [4-1:0] node9632;
	wire [4-1:0] node9633;
	wire [4-1:0] node9635;
	wire [4-1:0] node9638;
	wire [4-1:0] node9641;
	wire [4-1:0] node9642;
	wire [4-1:0] node9645;
	wire [4-1:0] node9646;
	wire [4-1:0] node9649;
	wire [4-1:0] node9652;
	wire [4-1:0] node9653;
	wire [4-1:0] node9654;
	wire [4-1:0] node9655;
	wire [4-1:0] node9659;
	wire [4-1:0] node9662;
	wire [4-1:0] node9663;
	wire [4-1:0] node9666;
	wire [4-1:0] node9667;
	wire [4-1:0] node9671;
	wire [4-1:0] node9672;
	wire [4-1:0] node9673;
	wire [4-1:0] node9674;
	wire [4-1:0] node9677;
	wire [4-1:0] node9680;
	wire [4-1:0] node9681;
	wire [4-1:0] node9682;
	wire [4-1:0] node9687;
	wire [4-1:0] node9688;
	wire [4-1:0] node9691;
	wire [4-1:0] node9693;
	wire [4-1:0] node9694;
	wire [4-1:0] node9695;
	wire [4-1:0] node9696;
	wire [4-1:0] node9702;
	wire [4-1:0] node9703;
	wire [4-1:0] node9704;
	wire [4-1:0] node9705;
	wire [4-1:0] node9707;
	wire [4-1:0] node9710;
	wire [4-1:0] node9712;
	wire [4-1:0] node9714;
	wire [4-1:0] node9717;
	wire [4-1:0] node9718;
	wire [4-1:0] node9719;
	wire [4-1:0] node9720;
	wire [4-1:0] node9724;
	wire [4-1:0] node9727;
	wire [4-1:0] node9728;
	wire [4-1:0] node9730;
	wire [4-1:0] node9733;
	wire [4-1:0] node9734;
	wire [4-1:0] node9738;
	wire [4-1:0] node9739;
	wire [4-1:0] node9740;
	wire [4-1:0] node9741;
	wire [4-1:0] node9745;
	wire [4-1:0] node9746;
	wire [4-1:0] node9749;
	wire [4-1:0] node9750;
	wire [4-1:0] node9752;
	wire [4-1:0] node9756;
	wire [4-1:0] node9757;
	wire [4-1:0] node9758;
	wire [4-1:0] node9762;
	wire [4-1:0] node9765;
	wire [4-1:0] node9766;
	wire [4-1:0] node9767;
	wire [4-1:0] node9768;
	wire [4-1:0] node9769;
	wire [4-1:0] node9770;
	wire [4-1:0] node9771;
	wire [4-1:0] node9772;
	wire [4-1:0] node9773;
	wire [4-1:0] node9778;
	wire [4-1:0] node9779;
	wire [4-1:0] node9782;
	wire [4-1:0] node9785;
	wire [4-1:0] node9786;
	wire [4-1:0] node9788;
	wire [4-1:0] node9790;
	wire [4-1:0] node9793;
	wire [4-1:0] node9794;
	wire [4-1:0] node9798;
	wire [4-1:0] node9799;
	wire [4-1:0] node9800;
	wire [4-1:0] node9801;
	wire [4-1:0] node9805;
	wire [4-1:0] node9808;
	wire [4-1:0] node9809;
	wire [4-1:0] node9811;
	wire [4-1:0] node9814;
	wire [4-1:0] node9815;
	wire [4-1:0] node9819;
	wire [4-1:0] node9820;
	wire [4-1:0] node9821;
	wire [4-1:0] node9822;
	wire [4-1:0] node9824;
	wire [4-1:0] node9827;
	wire [4-1:0] node9828;
	wire [4-1:0] node9832;
	wire [4-1:0] node9834;
	wire [4-1:0] node9836;
	wire [4-1:0] node9839;
	wire [4-1:0] node9840;
	wire [4-1:0] node9841;
	wire [4-1:0] node9844;
	wire [4-1:0] node9847;
	wire [4-1:0] node9849;
	wire [4-1:0] node9850;
	wire [4-1:0] node9853;
	wire [4-1:0] node9856;
	wire [4-1:0] node9857;
	wire [4-1:0] node9858;
	wire [4-1:0] node9859;
	wire [4-1:0] node9860;
	wire [4-1:0] node9862;
	wire [4-1:0] node9863;
	wire [4-1:0] node9865;
	wire [4-1:0] node9869;
	wire [4-1:0] node9872;
	wire [4-1:0] node9873;
	wire [4-1:0] node9874;
	wire [4-1:0] node9877;
	wire [4-1:0] node9880;
	wire [4-1:0] node9881;
	wire [4-1:0] node9883;
	wire [4-1:0] node9885;
	wire [4-1:0] node9889;
	wire [4-1:0] node9890;
	wire [4-1:0] node9891;
	wire [4-1:0] node9892;
	wire [4-1:0] node9893;
	wire [4-1:0] node9898;
	wire [4-1:0] node9901;
	wire [4-1:0] node9902;
	wire [4-1:0] node9903;
	wire [4-1:0] node9908;
	wire [4-1:0] node9909;
	wire [4-1:0] node9910;
	wire [4-1:0] node9911;
	wire [4-1:0] node9913;
	wire [4-1:0] node9915;
	wire [4-1:0] node9919;
	wire [4-1:0] node9920;
	wire [4-1:0] node9923;
	wire [4-1:0] node9924;
	wire [4-1:0] node9926;
	wire [4-1:0] node9929;
	wire [4-1:0] node9931;
	wire [4-1:0] node9934;
	wire [4-1:0] node9935;
	wire [4-1:0] node9936;
	wire [4-1:0] node9938;
	wire [4-1:0] node9941;
	wire [4-1:0] node9943;
	wire [4-1:0] node9947;
	wire [4-1:0] node9948;
	wire [4-1:0] node9949;
	wire [4-1:0] node9950;
	wire [4-1:0] node9951;
	wire [4-1:0] node9952;
	wire [4-1:0] node9953;
	wire [4-1:0] node9957;
	wire [4-1:0] node9960;
	wire [4-1:0] node9962;
	wire [4-1:0] node9963;
	wire [4-1:0] node9967;
	wire [4-1:0] node9968;
	wire [4-1:0] node9969;
	wire [4-1:0] node9970;
	wire [4-1:0] node9974;
	wire [4-1:0] node9975;
	wire [4-1:0] node9979;
	wire [4-1:0] node9980;
	wire [4-1:0] node9981;
	wire [4-1:0] node9986;
	wire [4-1:0] node9987;
	wire [4-1:0] node9988;
	wire [4-1:0] node9989;
	wire [4-1:0] node9992;
	wire [4-1:0] node9995;
	wire [4-1:0] node9997;
	wire [4-1:0] node10000;
	wire [4-1:0] node10001;
	wire [4-1:0] node10003;
	wire [4-1:0] node10005;
	wire [4-1:0] node10008;
	wire [4-1:0] node10010;
	wire [4-1:0] node10013;
	wire [4-1:0] node10014;
	wire [4-1:0] node10015;
	wire [4-1:0] node10016;
	wire [4-1:0] node10017;
	wire [4-1:0] node10018;
	wire [4-1:0] node10021;
	wire [4-1:0] node10024;
	wire [4-1:0] node10025;
	wire [4-1:0] node10028;
	wire [4-1:0] node10031;
	wire [4-1:0] node10032;
	wire [4-1:0] node10033;
	wire [4-1:0] node10038;
	wire [4-1:0] node10039;
	wire [4-1:0] node10040;
	wire [4-1:0] node10042;
	wire [4-1:0] node10045;
	wire [4-1:0] node10048;
	wire [4-1:0] node10050;
	wire [4-1:0] node10053;
	wire [4-1:0] node10055;
	wire [4-1:0] node10056;
	wire [4-1:0] node10057;
	wire [4-1:0] node10059;
	wire [4-1:0] node10063;
	wire [4-1:0] node10065;
	wire [4-1:0] node10068;
	wire [4-1:0] node10070;
	wire [4-1:0] node10071;
	wire [4-1:0] node10072;
	wire [4-1:0] node10074;
	wire [4-1:0] node10075;
	wire [4-1:0] node10076;
	wire [4-1:0] node10077;
	wire [4-1:0] node10079;
	wire [4-1:0] node10083;
	wire [4-1:0] node10084;
	wire [4-1:0] node10085;
	wire [4-1:0] node10086;
	wire [4-1:0] node10087;
	wire [4-1:0] node10092;
	wire [4-1:0] node10093;
	wire [4-1:0] node10096;
	wire [4-1:0] node10099;
	wire [4-1:0] node10103;
	wire [4-1:0] node10104;
	wire [4-1:0] node10105;
	wire [4-1:0] node10106;
	wire [4-1:0] node10107;
	wire [4-1:0] node10108;
	wire [4-1:0] node10109;
	wire [4-1:0] node10110;
	wire [4-1:0] node10113;
	wire [4-1:0] node10116;
	wire [4-1:0] node10117;
	wire [4-1:0] node10121;
	wire [4-1:0] node10122;
	wire [4-1:0] node10123;
	wire [4-1:0] node10126;
	wire [4-1:0] node10129;
	wire [4-1:0] node10130;
	wire [4-1:0] node10133;
	wire [4-1:0] node10136;
	wire [4-1:0] node10137;
	wire [4-1:0] node10138;
	wire [4-1:0] node10142;
	wire [4-1:0] node10145;
	wire [4-1:0] node10146;
	wire [4-1:0] node10147;
	wire [4-1:0] node10148;
	wire [4-1:0] node10152;
	wire [4-1:0] node10153;
	wire [4-1:0] node10157;
	wire [4-1:0] node10159;
	wire [4-1:0] node10162;
	wire [4-1:0] node10163;
	wire [4-1:0] node10164;
	wire [4-1:0] node10165;
	wire [4-1:0] node10167;
	wire [4-1:0] node10170;
	wire [4-1:0] node10173;
	wire [4-1:0] node10174;
	wire [4-1:0] node10176;
	wire [4-1:0] node10179;
	wire [4-1:0] node10180;
	wire [4-1:0] node10182;
	wire [4-1:0] node10185;
	wire [4-1:0] node10188;
	wire [4-1:0] node10189;
	wire [4-1:0] node10191;
	wire [4-1:0] node10194;
	wire [4-1:0] node10195;
	wire [4-1:0] node10196;
	wire [4-1:0] node10197;
	wire [4-1:0] node10202;
	wire [4-1:0] node10203;
	wire [4-1:0] node10204;
	wire [4-1:0] node10207;
	wire [4-1:0] node10209;
	wire [4-1:0] node10213;
	wire [4-1:0] node10214;
	wire [4-1:0] node10215;
	wire [4-1:0] node10216;
	wire [4-1:0] node10217;
	wire [4-1:0] node10222;
	wire [4-1:0] node10223;
	wire [4-1:0] node10224;
	wire [4-1:0] node10225;
	wire [4-1:0] node10229;
	wire [4-1:0] node10232;
	wire [4-1:0] node10233;
	wire [4-1:0] node10237;
	wire [4-1:0] node10238;
	wire [4-1:0] node10239;
	wire [4-1:0] node10241;
	wire [4-1:0] node10242;
	wire [4-1:0] node10245;
	wire [4-1:0] node10248;
	wire [4-1:0] node10249;
	wire [4-1:0] node10250;
	wire [4-1:0] node10251;
	wire [4-1:0] node10256;
	wire [4-1:0] node10259;
	wire [4-1:0] node10260;
	wire [4-1:0] node10261;
	wire [4-1:0] node10264;
	wire [4-1:0] node10265;
	wire [4-1:0] node10270;
	wire [4-1:0] node10272;
	wire [4-1:0] node10274;
	wire [4-1:0] node10275;
	wire [4-1:0] node10277;
	wire [4-1:0] node10278;
	wire [4-1:0] node10280;
	wire [4-1:0] node10281;
	wire [4-1:0] node10282;
	wire [4-1:0] node10287;
	wire [4-1:0] node10288;
	wire [4-1:0] node10289;

	assign outp = (inp[8]) ? node5124 : node1;
		assign node1 = (inp[9]) ? node2645 : node2;
			assign node2 = (inp[6]) ? node694 : node3;
				assign node3 = (inp[15]) ? node409 : node4;
					assign node4 = (inp[0]) ? 4'b1101 : node5;
						assign node5 = (inp[5]) ? node149 : node6;
							assign node6 = (inp[2]) ? 4'b1111 : node7;
								assign node7 = (inp[1]) ? node73 : node8;
									assign node8 = (inp[14]) ? node32 : node9;
										assign node9 = (inp[13]) ? node21 : node10;
											assign node10 = (inp[10]) ? node16 : node11;
												assign node11 = (inp[3]) ? 4'b1000 : node12;
													assign node12 = (inp[7]) ? 4'b1111 : 4'b0000;
												assign node16 = (inp[3]) ? node18 : 4'b0000;
													assign node18 = (inp[7]) ? 4'b0000 : 4'b0100;
											assign node21 = (inp[3]) ? node25 : node22;
												assign node22 = (inp[7]) ? 4'b1111 : 4'b1000;
												assign node25 = (inp[12]) ? node27 : 4'b1100;
													assign node27 = (inp[10]) ? node29 : 4'b0100;
														assign node29 = (inp[7]) ? 4'b1000 : 4'b1100;
										assign node32 = (inp[11]) ? node54 : node33;
											assign node33 = (inp[13]) ? node41 : node34;
												assign node34 = (inp[3]) ? 4'b1001 : node35;
													assign node35 = (inp[4]) ? node37 : 4'b1111;
														assign node37 = (inp[7]) ? 4'b1111 : 4'b1001;
												assign node41 = (inp[12]) ? node47 : node42;
													assign node42 = (inp[10]) ? node44 : 4'b0001;
														assign node44 = (inp[7]) ? 4'b1001 : 4'b1101;
													assign node47 = (inp[7]) ? node49 : 4'b0101;
														assign node49 = (inp[10]) ? 4'b0001 : node50;
															assign node50 = (inp[3]) ? 4'b0101 : 4'b0001;
											assign node54 = (inp[4]) ? node64 : node55;
												assign node55 = (inp[3]) ? 4'b1000 : node56;
													assign node56 = (inp[7]) ? 4'b1111 : node57;
														assign node57 = (inp[12]) ? node59 : 4'b0000;
															assign node59 = (inp[10]) ? 4'b1000 : 4'b1111;
												assign node64 = (inp[3]) ? node70 : node65;
													assign node65 = (inp[13]) ? 4'b1000 : node66;
														assign node66 = (inp[10]) ? 4'b0000 : 4'b1000;
													assign node70 = (inp[13]) ? 4'b1100 : 4'b0100;
									assign node73 = (inp[3]) ? node107 : node74;
										assign node74 = (inp[4]) ? node84 : node75;
											assign node75 = (inp[7]) ? 4'b1111 : node76;
												assign node76 = (inp[13]) ? 4'b1001 : node77;
													assign node77 = (inp[12]) ? 4'b1111 : node78;
														assign node78 = (inp[11]) ? 4'b0001 : 4'b0000;
											assign node84 = (inp[13]) ? node96 : node85;
												assign node85 = (inp[12]) ? node93 : node86;
													assign node86 = (inp[10]) ? 4'b0001 : node87;
														assign node87 = (inp[7]) ? node89 : 4'b0001;
															assign node89 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node93 = (inp[11]) ? 4'b0001 : 4'b1111;
												assign node96 = (inp[14]) ? node102 : node97;
													assign node97 = (inp[10]) ? 4'b1001 : node98;
														assign node98 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node102 = (inp[11]) ? 4'b1001 : node103;
														assign node103 = (inp[10]) ? 4'b1000 : 4'b0000;
										assign node107 = (inp[4]) ? node131 : node108;
											assign node108 = (inp[7]) ? node120 : node109;
												assign node109 = (inp[14]) ? node115 : node110;
													assign node110 = (inp[12]) ? node112 : 4'b0101;
														assign node112 = (inp[10]) ? 4'b0101 : 4'b1001;
													assign node115 = (inp[13]) ? node117 : 4'b1000;
														assign node117 = (inp[10]) ? 4'b1100 : 4'b0100;
												assign node120 = (inp[14]) ? node126 : node121;
													assign node121 = (inp[10]) ? node123 : 4'b1001;
														assign node123 = (inp[13]) ? 4'b1001 : 4'b0001;
													assign node126 = (inp[10]) ? 4'b1001 : node127;
														assign node127 = (inp[11]) ? 4'b0001 : 4'b0000;
											assign node131 = (inp[13]) ? node141 : node132;
												assign node132 = (inp[11]) ? node136 : node133;
													assign node133 = (inp[14]) ? 4'b0100 : 4'b0101;
													assign node136 = (inp[12]) ? node138 : 4'b0101;
														assign node138 = (inp[10]) ? 4'b0101 : 4'b1101;
												assign node141 = (inp[10]) ? node143 : 4'b0101;
													assign node143 = (inp[14]) ? node145 : 4'b1101;
														assign node145 = (inp[7]) ? 4'b1100 : 4'b1101;
							assign node149 = (inp[1]) ? node291 : node150;
								assign node150 = (inp[14]) ? node204 : node151;
									assign node151 = (inp[13]) ? node181 : node152;
										assign node152 = (inp[10]) ? node168 : node153;
											assign node153 = (inp[12]) ? node163 : node154;
												assign node154 = (inp[3]) ? node160 : node155;
													assign node155 = (inp[4]) ? 4'b0000 : node156;
														assign node156 = (inp[11]) ? 4'b1111 : 4'b0000;
													assign node160 = (inp[2]) ? 4'b0000 : 4'b0100;
												assign node163 = (inp[3]) ? 4'b1000 : node164;
													assign node164 = (inp[7]) ? 4'b1111 : 4'b1000;
											assign node168 = (inp[3]) ? node176 : node169;
												assign node169 = (inp[4]) ? 4'b0000 : node170;
													assign node170 = (inp[7]) ? node172 : 4'b0000;
														assign node172 = (inp[2]) ? 4'b1111 : 4'b0100;
												assign node176 = (inp[7]) ? node178 : 4'b0100;
													assign node178 = (inp[4]) ? 4'b0100 : 4'b0000;
										assign node181 = (inp[12]) ? node189 : node182;
											assign node182 = (inp[3]) ? node186 : node183;
												assign node183 = (inp[7]) ? 4'b1100 : 4'b1000;
												assign node186 = (inp[4]) ? 4'b1100 : 4'b1000;
											assign node189 = (inp[10]) ? node201 : node190;
												assign node190 = (inp[7]) ? node194 : node191;
													assign node191 = (inp[3]) ? 4'b0100 : 4'b0000;
													assign node194 = (inp[11]) ? 4'b1111 : node195;
														assign node195 = (inp[3]) ? node197 : 4'b0000;
															assign node197 = (inp[4]) ? 4'b0100 : 4'b0000;
												assign node201 = (inp[2]) ? 4'b1000 : 4'b1100;
									assign node204 = (inp[11]) ? node250 : node205;
										assign node205 = (inp[13]) ? node225 : node206;
											assign node206 = (inp[2]) ? node214 : node207;
												assign node207 = (inp[3]) ? node209 : 4'b1101;
													assign node209 = (inp[7]) ? 4'b1001 : node210;
														assign node210 = (inp[4]) ? 4'b1101 : 4'b1001;
												assign node214 = (inp[12]) ? node220 : node215;
													assign node215 = (inp[10]) ? node217 : 4'b1111;
														assign node217 = (inp[3]) ? 4'b0101 : 4'b0001;
													assign node220 = (inp[4]) ? node222 : 4'b1001;
														assign node222 = (inp[3]) ? 4'b1101 : 4'b1001;
											assign node225 = (inp[12]) ? node239 : node226;
												assign node226 = (inp[10]) ? node232 : node227;
													assign node227 = (inp[7]) ? node229 : 4'b0001;
														assign node229 = (inp[3]) ? 4'b0001 : 4'b0101;
													assign node232 = (inp[2]) ? 4'b1001 : node233;
														assign node233 = (inp[3]) ? 4'b1101 : node234;
															assign node234 = (inp[4]) ? 4'b1001 : 4'b1101;
												assign node239 = (inp[2]) ? node247 : node240;
													assign node240 = (inp[7]) ? node242 : 4'b0001;
														assign node242 = (inp[3]) ? node244 : 4'b0101;
															assign node244 = (inp[10]) ? 4'b0001 : 4'b0101;
													assign node247 = (inp[3]) ? 4'b0101 : 4'b1111;
										assign node250 = (inp[13]) ? node272 : node251;
											assign node251 = (inp[3]) ? node263 : node252;
												assign node252 = (inp[4]) ? node258 : node253;
													assign node253 = (inp[10]) ? 4'b1111 : node254;
														assign node254 = (inp[7]) ? 4'b1100 : 4'b0000;
													assign node258 = (inp[12]) ? node260 : 4'b0000;
														assign node260 = (inp[7]) ? 4'b0000 : 4'b1000;
												assign node263 = (inp[4]) ? 4'b0100 : node264;
													assign node264 = (inp[7]) ? 4'b0000 : node265;
														assign node265 = (inp[10]) ? 4'b0100 : node266;
															assign node266 = (inp[2]) ? 4'b0100 : 4'b1000;
											assign node272 = (inp[2]) ? node286 : node273;
												assign node273 = (inp[10]) ? node279 : node274;
													assign node274 = (inp[7]) ? 4'b0100 : node275;
														assign node275 = (inp[3]) ? 4'b1100 : 4'b1000;
													assign node279 = (inp[4]) ? 4'b1000 : node280;
														assign node280 = (inp[3]) ? 4'b1000 : node281;
															assign node281 = (inp[7]) ? 4'b1100 : 4'b1000;
												assign node286 = (inp[3]) ? node288 : 4'b1111;
													assign node288 = (inp[7]) ? 4'b0100 : 4'b1100;
								assign node291 = (inp[11]) ? node349 : node292;
									assign node292 = (inp[14]) ? node322 : node293;
										assign node293 = (inp[7]) ? node309 : node294;
											assign node294 = (inp[3]) ? node302 : node295;
												assign node295 = (inp[13]) ? 4'b1001 : node296;
													assign node296 = (inp[10]) ? 4'b0001 : node297;
														assign node297 = (inp[4]) ? 4'b0001 : 4'b1111;
												assign node302 = (inp[12]) ? node304 : 4'b0101;
													assign node304 = (inp[4]) ? 4'b1101 : node305;
														assign node305 = (inp[10]) ? 4'b1101 : 4'b1001;
											assign node309 = (inp[2]) ? node315 : node310;
												assign node310 = (inp[13]) ? node312 : 4'b0101;
													assign node312 = (inp[4]) ? 4'b0001 : 4'b0101;
												assign node315 = (inp[3]) ? 4'b0001 : node316;
													assign node316 = (inp[4]) ? node318 : 4'b1111;
														assign node318 = (inp[10]) ? 4'b0001 : 4'b1111;
										assign node322 = (inp[13]) ? node336 : node323;
											assign node323 = (inp[3]) ? node329 : node324;
												assign node324 = (inp[7]) ? node326 : 4'b0000;
													assign node326 = (inp[4]) ? 4'b0000 : 4'b0100;
												assign node329 = (inp[10]) ? node333 : node330;
													assign node330 = (inp[12]) ? 4'b1000 : 4'b0100;
													assign node333 = (inp[7]) ? 4'b0000 : 4'b0100;
											assign node336 = (inp[3]) ? node342 : node337;
												assign node337 = (inp[4]) ? 4'b1000 : node338;
													assign node338 = (inp[2]) ? 4'b1111 : 4'b1000;
												assign node342 = (inp[10]) ? 4'b1100 : node343;
													assign node343 = (inp[7]) ? 4'b0000 : node344;
														assign node344 = (inp[12]) ? 4'b0100 : 4'b1100;
									assign node349 = (inp[3]) ? node379 : node350;
										assign node350 = (inp[7]) ? node362 : node351;
											assign node351 = (inp[13]) ? node357 : node352;
												assign node352 = (inp[10]) ? 4'b0001 : node353;
													assign node353 = (inp[14]) ? 4'b0001 : 4'b1111;
												assign node357 = (inp[2]) ? node359 : 4'b1001;
													assign node359 = (inp[12]) ? 4'b0001 : 4'b1001;
											assign node362 = (inp[2]) ? node374 : node363;
												assign node363 = (inp[4]) ? node371 : node364;
													assign node364 = (inp[14]) ? node366 : 4'b1101;
														assign node366 = (inp[13]) ? 4'b0101 : node367;
															assign node367 = (inp[12]) ? 4'b1101 : 4'b0101;
													assign node371 = (inp[13]) ? 4'b1001 : 4'b1101;
												assign node374 = (inp[4]) ? node376 : 4'b1111;
													assign node376 = (inp[10]) ? 4'b0001 : 4'b1111;
										assign node379 = (inp[7]) ? node389 : node380;
											assign node380 = (inp[13]) ? node386 : node381;
												assign node381 = (inp[10]) ? 4'b0101 : node382;
													assign node382 = (inp[12]) ? 4'b1101 : 4'b0101;
												assign node386 = (inp[10]) ? 4'b1101 : 4'b0101;
											assign node389 = (inp[4]) ? node399 : node390;
												assign node390 = (inp[2]) ? node392 : 4'b0001;
													assign node392 = (inp[13]) ? node396 : node393;
														assign node393 = (inp[10]) ? 4'b0001 : 4'b1001;
														assign node396 = (inp[10]) ? 4'b1001 : 4'b0001;
												assign node399 = (inp[2]) ? node403 : node400;
													assign node400 = (inp[14]) ? 4'b1101 : 4'b1001;
													assign node403 = (inp[10]) ? 4'b0101 : node404;
														assign node404 = (inp[14]) ? 4'b0101 : 4'b1101;
					assign node409 = (inp[0]) ? 4'b1001 : node410;
						assign node410 = (inp[5]) ? node476 : node411;
							assign node411 = (inp[3]) ? node413 : 4'b1011;
								assign node413 = (inp[2]) ? 4'b1011 : node414;
									assign node414 = (inp[4]) ? node434 : node415;
										assign node415 = (inp[7]) ? 4'b1011 : node416;
											assign node416 = (inp[13]) ? node426 : node417;
												assign node417 = (inp[10]) ? node423 : node418;
													assign node418 = (inp[14]) ? 4'b1011 : node419;
														assign node419 = (inp[12]) ? 4'b1011 : 4'b0001;
													assign node423 = (inp[1]) ? 4'b0001 : 4'b0000;
												assign node426 = (inp[10]) ? node428 : 4'b0000;
													assign node428 = (inp[11]) ? node430 : 4'b1001;
														assign node430 = (inp[12]) ? 4'b1001 : 4'b1000;
										assign node434 = (inp[1]) ? node454 : node435;
											assign node435 = (inp[14]) ? node443 : node436;
												assign node436 = (inp[13]) ? node438 : 4'b0000;
													assign node438 = (inp[12]) ? node440 : 4'b1000;
														assign node440 = (inp[10]) ? 4'b1000 : 4'b0000;
												assign node443 = (inp[11]) ? node451 : node444;
													assign node444 = (inp[10]) ? node446 : 4'b0001;
														assign node446 = (inp[7]) ? node448 : 4'b1001;
															assign node448 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node451 = (inp[13]) ? 4'b1000 : 4'b0000;
											assign node454 = (inp[11]) ? node466 : node455;
												assign node455 = (inp[14]) ? node459 : node456;
													assign node456 = (inp[13]) ? 4'b1001 : 4'b0001;
													assign node459 = (inp[10]) ? 4'b1000 : node460;
														assign node460 = (inp[7]) ? node462 : 4'b0000;
															assign node462 = (inp[13]) ? 4'b0000 : 4'b1011;
												assign node466 = (inp[7]) ? node472 : node467;
													assign node467 = (inp[10]) ? node469 : 4'b1001;
														assign node469 = (inp[13]) ? 4'b1001 : 4'b0001;
													assign node472 = (inp[13]) ? 4'b1001 : 4'b1011;
							assign node476 = (inp[2]) ? node640 : node477;
								assign node477 = (inp[1]) ? node563 : node478;
									assign node478 = (inp[14]) ? node516 : node479;
										assign node479 = (inp[13]) ? node495 : node480;
											assign node480 = (inp[10]) ? node490 : node481;
												assign node481 = (inp[12]) ? node487 : node482;
													assign node482 = (inp[4]) ? 4'b0000 : node483;
														assign node483 = (inp[11]) ? 4'b0000 : 4'b0100;
													assign node487 = (inp[4]) ? 4'b1100 : 4'b1000;
												assign node490 = (inp[3]) ? node492 : 4'b0100;
													assign node492 = (inp[7]) ? 4'b0100 : 4'b0000;
											assign node495 = (inp[12]) ? node503 : node496;
												assign node496 = (inp[4]) ? 4'b1100 : node497;
													assign node497 = (inp[3]) ? node499 : 4'b1000;
														assign node499 = (inp[7]) ? 4'b1100 : 4'b1000;
												assign node503 = (inp[10]) ? node513 : node504;
													assign node504 = (inp[11]) ? node510 : node505;
														assign node505 = (inp[3]) ? 4'b0000 : node506;
															assign node506 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node510 = (inp[3]) ? 4'b0100 : 4'b0000;
													assign node513 = (inp[7]) ? 4'b1000 : 4'b1100;
										assign node516 = (inp[11]) ? node538 : node517;
											assign node517 = (inp[3]) ? node533 : node518;
												assign node518 = (inp[4]) ? node528 : node519;
													assign node519 = (inp[7]) ? node521 : 4'b1001;
														assign node521 = (inp[13]) ? node525 : node522;
															assign node522 = (inp[10]) ? 4'b0001 : 4'b1001;
															assign node525 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node528 = (inp[13]) ? 4'b0101 : node529;
														assign node529 = (inp[7]) ? 4'b1001 : 4'b1101;
												assign node533 = (inp[7]) ? 4'b1101 : node534;
													assign node534 = (inp[10]) ? 4'b1001 : 4'b0001;
											assign node538 = (inp[13]) ? node554 : node539;
												assign node539 = (inp[10]) ? node547 : node540;
													assign node540 = (inp[12]) ? node544 : node541;
														assign node541 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node544 = (inp[7]) ? 4'b1100 : 4'b1000;
													assign node547 = (inp[7]) ? node549 : 4'b0100;
														assign node549 = (inp[3]) ? node551 : 4'b0000;
															assign node551 = (inp[4]) ? 4'b0000 : 4'b0100;
												assign node554 = (inp[10]) ? node558 : node555;
													assign node555 = (inp[3]) ? 4'b1000 : 4'b0000;
													assign node558 = (inp[12]) ? node560 : 4'b1000;
														assign node560 = (inp[3]) ? 4'b1000 : 4'b1100;
									assign node563 = (inp[13]) ? node605 : node564;
										assign node564 = (inp[10]) ? node586 : node565;
											assign node565 = (inp[12]) ? node575 : node566;
												assign node566 = (inp[3]) ? 4'b0001 : node567;
													assign node567 = (inp[11]) ? 4'b0101 : node568;
														assign node568 = (inp[4]) ? 4'b0101 : node569;
															assign node569 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node575 = (inp[3]) ? 4'b1101 : node576;
													assign node576 = (inp[7]) ? node582 : node577;
														assign node577 = (inp[4]) ? node579 : 4'b1001;
															assign node579 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node582 = (inp[11]) ? 4'b1001 : 4'b1000;
											assign node586 = (inp[14]) ? node598 : node587;
												assign node587 = (inp[3]) ? node593 : node588;
													assign node588 = (inp[4]) ? 4'b0101 : node589;
														assign node589 = (inp[7]) ? 4'b0001 : 4'b0101;
													assign node593 = (inp[4]) ? 4'b0001 : node594;
														assign node594 = (inp[7]) ? 4'b0101 : 4'b0001;
												assign node598 = (inp[11]) ? 4'b0001 : node599;
													assign node599 = (inp[4]) ? node601 : 4'b0100;
														assign node601 = (inp[3]) ? 4'b0000 : 4'b0100;
										assign node605 = (inp[14]) ? node621 : node606;
											assign node606 = (inp[3]) ? node616 : node607;
												assign node607 = (inp[10]) ? node611 : node608;
													assign node608 = (inp[4]) ? 4'b0101 : 4'b1101;
													assign node611 = (inp[11]) ? 4'b1101 : node612;
														assign node612 = (inp[4]) ? 4'b1101 : 4'b1001;
												assign node616 = (inp[4]) ? 4'b1001 : node617;
													assign node617 = (inp[7]) ? 4'b1101 : 4'b1001;
											assign node621 = (inp[11]) ? node629 : node622;
												assign node622 = (inp[12]) ? 4'b1000 : node623;
													assign node623 = (inp[7]) ? 4'b1100 : node624;
														assign node624 = (inp[3]) ? 4'b1000 : 4'b1100;
												assign node629 = (inp[12]) ? node633 : node630;
													assign node630 = (inp[3]) ? 4'b1101 : 4'b1001;
													assign node633 = (inp[4]) ? 4'b1101 : node634;
														assign node634 = (inp[3]) ? 4'b0001 : node635;
															assign node635 = (inp[7]) ? 4'b0001 : 4'b0101;
								assign node640 = (inp[3]) ? node642 : 4'b1011;
									assign node642 = (inp[4]) ? node660 : node643;
										assign node643 = (inp[7]) ? 4'b1011 : node644;
											assign node644 = (inp[14]) ? node656 : node645;
												assign node645 = (inp[1]) ? node651 : node646;
													assign node646 = (inp[11]) ? node648 : 4'b0000;
														assign node648 = (inp[13]) ? 4'b1000 : 4'b0000;
													assign node651 = (inp[13]) ? 4'b1001 : node652;
														assign node652 = (inp[12]) ? 4'b1011 : 4'b0001;
												assign node656 = (inp[1]) ? 4'b0000 : 4'b0001;
										assign node660 = (inp[1]) ? node676 : node661;
											assign node661 = (inp[13]) ? node669 : node662;
												assign node662 = (inp[11]) ? 4'b0000 : node663;
													assign node663 = (inp[14]) ? node665 : 4'b0000;
														assign node665 = (inp[10]) ? 4'b1011 : 4'b1001;
												assign node669 = (inp[11]) ? 4'b1000 : node670;
													assign node670 = (inp[7]) ? node672 : 4'b1000;
														assign node672 = (inp[14]) ? 4'b0001 : 4'b0000;
											assign node676 = (inp[13]) ? node684 : node677;
												assign node677 = (inp[11]) ? node679 : 4'b0000;
													assign node679 = (inp[12]) ? node681 : 4'b0001;
														assign node681 = (inp[10]) ? 4'b0001 : 4'b1001;
												assign node684 = (inp[12]) ? node690 : node685;
													assign node685 = (inp[14]) ? node687 : 4'b1001;
														assign node687 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node690 = (inp[10]) ? 4'b1001 : 4'b0001;
				assign node694 = (inp[5]) ? node1558 : node695;
					assign node695 = (inp[0]) ? node1355 : node696;
						assign node696 = (inp[11]) ? node1034 : node697;
							assign node697 = (inp[2]) ? node873 : node698;
								assign node698 = (inp[10]) ? node774 : node699;
									assign node699 = (inp[1]) ? node741 : node700;
										assign node700 = (inp[12]) ? node722 : node701;
											assign node701 = (inp[15]) ? node713 : node702;
												assign node702 = (inp[3]) ? node708 : node703;
													assign node703 = (inp[14]) ? node705 : 4'b0000;
														assign node705 = (inp[4]) ? 4'b0100 : 4'b0000;
													assign node708 = (inp[4]) ? node710 : 4'b0000;
														assign node710 = (inp[14]) ? 4'b1000 : 4'b1001;
												assign node713 = (inp[4]) ? node717 : node714;
													assign node714 = (inp[3]) ? 4'b0100 : 4'b1100;
													assign node717 = (inp[7]) ? node719 : 4'b0000;
														assign node719 = (inp[13]) ? 4'b0000 : 4'b0100;
											assign node722 = (inp[14]) ? node734 : node723;
												assign node723 = (inp[3]) ? node731 : node724;
													assign node724 = (inp[4]) ? node726 : 4'b1100;
														assign node726 = (inp[7]) ? 4'b1000 : node727;
															assign node727 = (inp[13]) ? 4'b1100 : 4'b1000;
													assign node731 = (inp[15]) ? 4'b1000 : 4'b0001;
												assign node734 = (inp[3]) ? 4'b1100 : node735;
													assign node735 = (inp[13]) ? 4'b0101 : node736;
														assign node736 = (inp[7]) ? 4'b1000 : 4'b1001;
										assign node741 = (inp[15]) ? node759 : node742;
											assign node742 = (inp[3]) ? node752 : node743;
												assign node743 = (inp[12]) ? node749 : node744;
													assign node744 = (inp[7]) ? 4'b0000 : node745;
														assign node745 = (inp[4]) ? 4'b0100 : 4'b0000;
													assign node749 = (inp[4]) ? 4'b0100 : 4'b1100;
												assign node752 = (inp[4]) ? node754 : 4'b0000;
													assign node754 = (inp[7]) ? 4'b1001 : node755;
														assign node755 = (inp[13]) ? 4'b0100 : 4'b1000;
											assign node759 = (inp[14]) ? 4'b0000 : node760;
												assign node760 = (inp[7]) ? node762 : 4'b1101;
													assign node762 = (inp[3]) ? node768 : node763;
														assign node763 = (inp[13]) ? node765 : 4'b0101;
															assign node765 = (inp[4]) ? 4'b0000 : 4'b0001;
														assign node768 = (inp[4]) ? node770 : 4'b0100;
															assign node770 = (inp[13]) ? 4'b0000 : 4'b0100;
									assign node774 = (inp[1]) ? node818 : node775;
										assign node775 = (inp[12]) ? node797 : node776;
											assign node776 = (inp[14]) ? node794 : node777;
												assign node777 = (inp[3]) ? node787 : node778;
													assign node778 = (inp[7]) ? 4'b0100 : node779;
														assign node779 = (inp[15]) ? node783 : node780;
															assign node780 = (inp[4]) ? 4'b1100 : 4'b1000;
															assign node783 = (inp[13]) ? 4'b1000 : 4'b0100;
													assign node787 = (inp[4]) ? node791 : node788;
														assign node788 = (inp[7]) ? 4'b1100 : 4'b1000;
														assign node791 = (inp[13]) ? 4'b0001 : 4'b1000;
												assign node794 = (inp[3]) ? 4'b1100 : 4'b1000;
											assign node797 = (inp[13]) ? node811 : node798;
												assign node798 = (inp[14]) ? node806 : node799;
													assign node799 = (inp[7]) ? node801 : 4'b0100;
														assign node801 = (inp[15]) ? node803 : 4'b0000;
															assign node803 = (inp[4]) ? 4'b0100 : 4'b0000;
													assign node806 = (inp[15]) ? node808 : 4'b0000;
														assign node808 = (inp[4]) ? 4'b0000 : 4'b0100;
												assign node811 = (inp[4]) ? node815 : node812;
													assign node812 = (inp[3]) ? 4'b0100 : 4'b0101;
													assign node815 = (inp[3]) ? 4'b0001 : 4'b0000;
										assign node818 = (inp[13]) ? node854 : node819;
											assign node819 = (inp[7]) ? node835 : node820;
												assign node820 = (inp[3]) ? node830 : node821;
													assign node821 = (inp[4]) ? node827 : node822;
														assign node822 = (inp[15]) ? node824 : 4'b1000;
															assign node824 = (inp[14]) ? 4'b0100 : 4'b0101;
														assign node827 = (inp[12]) ? 4'b1100 : 4'b1000;
													assign node830 = (inp[4]) ? 4'b0101 : node831;
														assign node831 = (inp[15]) ? 4'b1100 : 4'b1000;
												assign node835 = (inp[3]) ? node849 : node836;
													assign node836 = (inp[14]) ? node842 : node837;
														assign node837 = (inp[12]) ? node839 : 4'b0101;
															assign node839 = (inp[4]) ? 4'b1000 : 4'b0101;
														assign node842 = (inp[4]) ? node846 : node843;
															assign node843 = (inp[15]) ? 4'b0000 : 4'b0100;
															assign node846 = (inp[15]) ? 4'b0100 : 4'b1000;
													assign node849 = (inp[4]) ? 4'b0000 : node850;
														assign node850 = (inp[12]) ? 4'b1000 : 4'b1100;
											assign node854 = (inp[4]) ? node864 : node855;
												assign node855 = (inp[15]) ? node861 : node856;
													assign node856 = (inp[14]) ? node858 : 4'b1000;
														assign node858 = (inp[3]) ? 4'b0001 : 4'b1000;
													assign node861 = (inp[3]) ? 4'b1100 : 4'b1000;
												assign node864 = (inp[3]) ? node866 : 4'b1100;
													assign node866 = (inp[15]) ? node870 : node867;
														assign node867 = (inp[12]) ? 4'b0101 : 4'b1101;
														assign node870 = (inp[12]) ? 4'b1000 : 4'b1001;
								assign node873 = (inp[3]) ? node955 : node874;
									assign node874 = (inp[15]) ? node912 : node875;
										assign node875 = (inp[10]) ? node895 : node876;
											assign node876 = (inp[7]) ? node886 : node877;
												assign node877 = (inp[13]) ? node881 : node878;
													assign node878 = (inp[12]) ? 4'b1000 : 4'b0001;
													assign node881 = (inp[14]) ? 4'b0001 : node882;
														assign node882 = (inp[1]) ? 4'b0001 : 4'b0000;
												assign node886 = (inp[4]) ? node888 : 4'b0100;
													assign node888 = (inp[13]) ? node892 : node889;
														assign node889 = (inp[1]) ? 4'b0001 : 4'b0000;
														assign node892 = (inp[12]) ? 4'b0000 : 4'b1000;
											assign node895 = (inp[7]) ? node901 : node896;
												assign node896 = (inp[13]) ? node898 : 4'b0001;
													assign node898 = (inp[12]) ? 4'b1001 : 4'b1000;
												assign node901 = (inp[14]) ? node903 : 4'b0101;
													assign node903 = (inp[4]) ? node909 : node904;
														assign node904 = (inp[13]) ? node906 : 4'b1101;
															assign node906 = (inp[12]) ? 4'b0101 : 4'b1101;
														assign node909 = (inp[12]) ? 4'b1101 : 4'b0001;
										assign node912 = (inp[7]) ? node938 : node913;
											assign node913 = (inp[12]) ? node919 : node914;
												assign node914 = (inp[13]) ? 4'b1100 : node915;
													assign node915 = (inp[1]) ? 4'b0101 : 4'b0100;
												assign node919 = (inp[10]) ? node927 : node920;
													assign node920 = (inp[13]) ? node922 : 4'b1101;
														assign node922 = (inp[14]) ? node924 : 4'b0101;
															assign node924 = (inp[4]) ? 4'b0101 : 4'b0100;
													assign node927 = (inp[4]) ? node933 : node928;
														assign node928 = (inp[1]) ? node930 : 4'b1001;
															assign node930 = (inp[14]) ? 4'b0100 : 4'b1101;
														assign node933 = (inp[1]) ? 4'b1101 : node934;
															assign node934 = (inp[14]) ? 4'b1101 : 4'b1100;
											assign node938 = (inp[12]) ? node946 : node939;
												assign node939 = (inp[4]) ? node943 : node940;
													assign node940 = (inp[13]) ? 4'b1000 : 4'b0000;
													assign node943 = (inp[10]) ? 4'b0100 : 4'b1100;
												assign node946 = (inp[1]) ? node950 : node947;
													assign node947 = (inp[14]) ? 4'b1001 : 4'b1000;
													assign node950 = (inp[13]) ? node952 : 4'b1000;
														assign node952 = (inp[4]) ? 4'b0101 : 4'b0001;
									assign node955 = (inp[15]) ? node995 : node956;
										assign node956 = (inp[4]) ? node978 : node957;
											assign node957 = (inp[7]) ? node963 : node958;
												assign node958 = (inp[10]) ? 4'b1000 : node959;
													assign node959 = (inp[12]) ? 4'b1000 : 4'b0000;
												assign node963 = (inp[12]) ? node965 : 4'b0000;
													assign node965 = (inp[10]) ? node969 : node966;
														assign node966 = (inp[1]) ? 4'b1000 : 4'b1001;
														assign node969 = (inp[13]) ? node975 : node970;
															assign node970 = (inp[1]) ? node972 : 4'b0000;
																assign node972 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node975 = (inp[14]) ? 4'b0000 : 4'b1000;
											assign node978 = (inp[13]) ? node986 : node979;
												assign node979 = (inp[10]) ? node981 : 4'b1000;
													assign node981 = (inp[12]) ? node983 : 4'b1000;
														assign node983 = (inp[7]) ? 4'b0000 : 4'b0100;
												assign node986 = (inp[7]) ? node992 : node987;
													assign node987 = (inp[12]) ? 4'b1100 : node988;
														assign node988 = (inp[1]) ? 4'b0100 : 4'b1100;
													assign node992 = (inp[12]) ? 4'b0100 : 4'b1100;
										assign node995 = (inp[14]) ? node1019 : node996;
											assign node996 = (inp[1]) ? node1006 : node997;
												assign node997 = (inp[13]) ? node1003 : node998;
													assign node998 = (inp[12]) ? node1000 : 4'b0000;
														assign node1000 = (inp[4]) ? 4'b0000 : 4'b0100;
													assign node1003 = (inp[4]) ? 4'b0000 : 4'b1000;
												assign node1006 = (inp[12]) ? node1010 : node1007;
													assign node1007 = (inp[7]) ? 4'b0001 : 4'b0000;
													assign node1010 = (inp[7]) ? node1012 : 4'b0001;
														assign node1012 = (inp[4]) ? node1014 : 4'b1101;
															assign node1014 = (inp[13]) ? 4'b0000 : node1015;
																assign node1015 = (inp[10]) ? 4'b0001 : 4'b1101;
											assign node1019 = (inp[1]) ? node1031 : node1020;
												assign node1020 = (inp[13]) ? node1022 : 4'b1101;
													assign node1022 = (inp[4]) ? node1028 : node1023;
														assign node1023 = (inp[7]) ? 4'b0101 : node1024;
															assign node1024 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node1028 = (inp[7]) ? 4'b0000 : 4'b1000;
												assign node1031 = (inp[13]) ? 4'b1000 : 4'b0000;
							assign node1034 = (inp[1]) ? node1196 : node1035;
								assign node1035 = (inp[13]) ? node1111 : node1036;
									assign node1036 = (inp[2]) ? node1078 : node1037;
										assign node1037 = (inp[12]) ? node1059 : node1038;
											assign node1038 = (inp[10]) ? node1050 : node1039;
												assign node1039 = (inp[7]) ? node1045 : node1040;
													assign node1040 = (inp[15]) ? 4'b0001 : node1041;
														assign node1041 = (inp[4]) ? 4'b0101 : 4'b0001;
													assign node1045 = (inp[15]) ? node1047 : 4'b0000;
														assign node1047 = (inp[14]) ? 4'b0100 : 4'b0101;
												assign node1050 = (inp[14]) ? node1056 : node1051;
													assign node1051 = (inp[3]) ? 4'b0000 : node1052;
														assign node1052 = (inp[7]) ? 4'b0000 : 4'b0100;
													assign node1056 = (inp[15]) ? 4'b1001 : 4'b0100;
											assign node1059 = (inp[10]) ? node1067 : node1060;
												assign node1060 = (inp[15]) ? node1064 : node1061;
													assign node1061 = (inp[7]) ? 4'b0000 : 4'b1001;
													assign node1064 = (inp[3]) ? 4'b1101 : 4'b1000;
												assign node1067 = (inp[14]) ? node1071 : node1068;
													assign node1068 = (inp[4]) ? 4'b0001 : 4'b0101;
													assign node1071 = (inp[15]) ? node1075 : node1072;
														assign node1072 = (inp[7]) ? 4'b1000 : 4'b0001;
														assign node1075 = (inp[4]) ? 4'b0101 : 4'b0000;
										assign node1078 = (inp[12]) ? node1098 : node1079;
											assign node1079 = (inp[15]) ? node1087 : node1080;
												assign node1080 = (inp[3]) ? node1082 : 4'b0000;
													assign node1082 = (inp[7]) ? 4'b0000 : node1083;
														assign node1083 = (inp[10]) ? 4'b1001 : 4'b0001;
												assign node1087 = (inp[3]) ? node1093 : node1088;
													assign node1088 = (inp[7]) ? node1090 : 4'b0100;
														assign node1090 = (inp[14]) ? 4'b0100 : 4'b0000;
													assign node1093 = (inp[4]) ? 4'b1001 : node1094;
														assign node1094 = (inp[7]) ? 4'b0100 : 4'b0000;
											assign node1098 = (inp[10]) ? node1106 : node1099;
												assign node1099 = (inp[14]) ? node1101 : 4'b1100;
													assign node1101 = (inp[7]) ? node1103 : 4'b1000;
														assign node1103 = (inp[3]) ? 4'b1100 : 4'b1000;
												assign node1106 = (inp[4]) ? node1108 : 4'b0100;
													assign node1108 = (inp[15]) ? 4'b0100 : 4'b0000;
									assign node1111 = (inp[12]) ? node1157 : node1112;
										assign node1112 = (inp[2]) ? node1138 : node1113;
											assign node1113 = (inp[10]) ? node1133 : node1114;
												assign node1114 = (inp[7]) ? node1128 : node1115;
													assign node1115 = (inp[14]) ? node1125 : node1116;
														assign node1116 = (inp[3]) ? node1120 : node1117;
															assign node1117 = (inp[15]) ? 4'b0001 : 4'b0101;
															assign node1120 = (inp[4]) ? node1122 : 4'b0101;
																assign node1122 = (inp[15]) ? 4'b1000 : 4'b1100;
														assign node1125 = (inp[3]) ? 4'b1000 : 4'b1100;
													assign node1128 = (inp[15]) ? node1130 : 4'b0001;
														assign node1130 = (inp[4]) ? 4'b0001 : 4'b0101;
												assign node1133 = (inp[4]) ? 4'b1100 : node1134;
													assign node1134 = (inp[14]) ? 4'b1001 : 4'b1101;
											assign node1138 = (inp[15]) ? node1146 : node1139;
												assign node1139 = (inp[3]) ? node1141 : 4'b1000;
													assign node1141 = (inp[4]) ? 4'b1101 : node1142;
														assign node1142 = (inp[7]) ? 4'b0001 : 4'b1001;
												assign node1146 = (inp[14]) ? node1152 : node1147;
													assign node1147 = (inp[4]) ? node1149 : 4'b1000;
														assign node1149 = (inp[7]) ? 4'b1001 : 4'b1100;
													assign node1152 = (inp[4]) ? 4'b1100 : node1153;
														assign node1153 = (inp[3]) ? 4'b1100 : 4'b1000;
										assign node1157 = (inp[10]) ? node1179 : node1158;
											assign node1158 = (inp[3]) ? node1166 : node1159;
												assign node1159 = (inp[4]) ? node1163 : node1160;
													assign node1160 = (inp[15]) ? 4'b0000 : 4'b0100;
													assign node1163 = (inp[15]) ? 4'b1001 : 4'b1101;
												assign node1166 = (inp[15]) ? node1176 : node1167;
													assign node1167 = (inp[14]) ? node1171 : node1168;
														assign node1168 = (inp[7]) ? 4'b1101 : 4'b1001;
														assign node1171 = (inp[4]) ? node1173 : 4'b1001;
															assign node1173 = (inp[2]) ? 4'b1001 : 4'b1000;
													assign node1176 = (inp[14]) ? 4'b1101 : 4'b1001;
											assign node1179 = (inp[4]) ? node1187 : node1180;
												assign node1180 = (inp[3]) ? node1184 : node1181;
													assign node1181 = (inp[14]) ? 4'b1100 : 4'b1000;
													assign node1184 = (inp[14]) ? 4'b0101 : 4'b0001;
												assign node1187 = (inp[15]) ? node1189 : 4'b0101;
													assign node1189 = (inp[14]) ? 4'b0001 : node1190;
														assign node1190 = (inp[7]) ? node1192 : 4'b0001;
															assign node1192 = (inp[3]) ? 4'b0000 : 4'b0001;
								assign node1196 = (inp[10]) ? node1280 : node1197;
									assign node1197 = (inp[7]) ? node1227 : node1198;
										assign node1198 = (inp[15]) ? node1206 : node1199;
											assign node1199 = (inp[4]) ? node1201 : 4'b0001;
												assign node1201 = (inp[13]) ? 4'b0101 : node1202;
													assign node1202 = (inp[2]) ? 4'b0001 : 4'b1001;
											assign node1206 = (inp[3]) ? node1216 : node1207;
												assign node1207 = (inp[14]) ? node1211 : node1208;
													assign node1208 = (inp[4]) ? 4'b0001 : 4'b0101;
													assign node1211 = (inp[2]) ? 4'b1101 : node1212;
														assign node1212 = (inp[12]) ? 4'b1001 : 4'b0001;
												assign node1216 = (inp[13]) ? node1218 : 4'b0001;
													assign node1218 = (inp[4]) ? node1222 : node1219;
														assign node1219 = (inp[14]) ? 4'b0001 : 4'b1001;
														assign node1222 = (inp[14]) ? node1224 : 4'b0001;
															assign node1224 = (inp[12]) ? 4'b1001 : 4'b0001;
										assign node1227 = (inp[3]) ? node1253 : node1228;
											assign node1228 = (inp[15]) ? node1238 : node1229;
												assign node1229 = (inp[2]) ? node1233 : node1230;
													assign node1230 = (inp[12]) ? 4'b1101 : 4'b0101;
													assign node1233 = (inp[12]) ? 4'b0101 : node1234;
														assign node1234 = (inp[14]) ? 4'b0001 : 4'b1001;
												assign node1238 = (inp[2]) ? node1244 : node1239;
													assign node1239 = (inp[12]) ? 4'b1001 : node1240;
														assign node1240 = (inp[13]) ? 4'b1001 : 4'b0001;
													assign node1244 = (inp[4]) ? node1250 : node1245;
														assign node1245 = (inp[12]) ? 4'b0001 : node1246;
															assign node1246 = (inp[13]) ? 4'b1001 : 4'b0001;
														assign node1250 = (inp[13]) ? 4'b0101 : 4'b1001;
											assign node1253 = (inp[2]) ? node1263 : node1254;
												assign node1254 = (inp[13]) ? 4'b0001 : node1255;
													assign node1255 = (inp[14]) ? 4'b0101 : node1256;
														assign node1256 = (inp[15]) ? node1258 : 4'b1001;
															assign node1258 = (inp[4]) ? 4'b0101 : 4'b0001;
												assign node1263 = (inp[12]) ? node1271 : node1264;
													assign node1264 = (inp[4]) ? 4'b0001 : node1265;
														assign node1265 = (inp[15]) ? node1267 : 4'b0001;
															assign node1267 = (inp[13]) ? 4'b1101 : 4'b0101;
													assign node1271 = (inp[13]) ? node1275 : node1272;
														assign node1272 = (inp[15]) ? 4'b1101 : 4'b1001;
														assign node1275 = (inp[14]) ? node1277 : 4'b0101;
															assign node1277 = (inp[4]) ? 4'b0001 : 4'b0101;
									assign node1280 = (inp[13]) ? node1328 : node1281;
										assign node1281 = (inp[2]) ? node1313 : node1282;
											assign node1282 = (inp[14]) ? node1294 : node1283;
												assign node1283 = (inp[15]) ? node1291 : node1284;
													assign node1284 = (inp[3]) ? node1288 : node1285;
														assign node1285 = (inp[4]) ? 4'b1001 : 4'b0101;
														assign node1288 = (inp[4]) ? 4'b0101 : 4'b1001;
													assign node1291 = (inp[3]) ? 4'b1101 : 4'b0101;
												assign node1294 = (inp[3]) ? node1304 : node1295;
													assign node1295 = (inp[4]) ? node1299 : node1296;
														assign node1296 = (inp[7]) ? 4'b0101 : 4'b1001;
														assign node1299 = (inp[7]) ? 4'b1001 : node1300;
															assign node1300 = (inp[15]) ? 4'b1001 : 4'b1101;
													assign node1304 = (inp[4]) ? node1308 : node1305;
														assign node1305 = (inp[7]) ? 4'b1001 : 4'b1101;
														assign node1308 = (inp[15]) ? 4'b0001 : node1309;
															assign node1309 = (inp[7]) ? 4'b0001 : 4'b0101;
											assign node1313 = (inp[15]) ? node1317 : node1314;
												assign node1314 = (inp[3]) ? 4'b1001 : 4'b0001;
												assign node1317 = (inp[7]) ? node1321 : node1318;
													assign node1318 = (inp[4]) ? 4'b1001 : 4'b0001;
													assign node1321 = (inp[3]) ? node1325 : node1322;
														assign node1322 = (inp[4]) ? 4'b0101 : 4'b0001;
														assign node1325 = (inp[4]) ? 4'b0001 : 4'b0101;
										assign node1328 = (inp[2]) ? node1340 : node1329;
											assign node1329 = (inp[14]) ? node1331 : 4'b1001;
												assign node1331 = (inp[7]) ? node1337 : node1332;
													assign node1332 = (inp[4]) ? 4'b1001 : node1333;
														assign node1333 = (inp[15]) ? 4'b1101 : 4'b1001;
													assign node1337 = (inp[12]) ? 4'b1001 : 4'b1101;
											assign node1340 = (inp[7]) ? node1350 : node1341;
												assign node1341 = (inp[15]) ? node1347 : node1342;
													assign node1342 = (inp[3]) ? node1344 : 4'b1001;
														assign node1344 = (inp[14]) ? 4'b1101 : 4'b1001;
													assign node1347 = (inp[3]) ? 4'b1001 : 4'b1101;
												assign node1350 = (inp[4]) ? 4'b1001 : node1351;
													assign node1351 = (inp[3]) ? 4'b1001 : 4'b1101;
						assign node1355 = (inp[15]) ? node1507 : node1356;
							assign node1356 = (inp[2]) ? 4'b1101 : node1357;
								assign node1357 = (inp[1]) ? node1433 : node1358;
									assign node1358 = (inp[11]) ? node1406 : node1359;
										assign node1359 = (inp[14]) ? node1381 : node1360;
											assign node1360 = (inp[4]) ? node1376 : node1361;
												assign node1361 = (inp[10]) ? node1363 : 4'b1101;
													assign node1363 = (inp[13]) ? node1369 : node1364;
														assign node1364 = (inp[12]) ? node1366 : 4'b0000;
															assign node1366 = (inp[3]) ? 4'b0000 : 4'b1101;
														assign node1369 = (inp[7]) ? node1373 : node1370;
															assign node1370 = (inp[3]) ? 4'b1100 : 4'b1000;
															assign node1373 = (inp[3]) ? 4'b1000 : 4'b1101;
												assign node1376 = (inp[12]) ? node1378 : 4'b0100;
													assign node1378 = (inp[10]) ? 4'b0000 : 4'b1000;
											assign node1381 = (inp[13]) ? node1391 : node1382;
												assign node1382 = (inp[3]) ? node1386 : node1383;
													assign node1383 = (inp[12]) ? 4'b1101 : 4'b0001;
													assign node1386 = (inp[7]) ? 4'b1001 : node1387;
														assign node1387 = (inp[4]) ? 4'b1101 : 4'b1001;
												assign node1391 = (inp[10]) ? node1397 : node1392;
													assign node1392 = (inp[3]) ? 4'b0101 : node1393;
														assign node1393 = (inp[12]) ? 4'b1101 : 4'b0001;
													assign node1397 = (inp[12]) ? 4'b0001 : node1398;
														assign node1398 = (inp[7]) ? node1400 : 4'b1001;
															assign node1400 = (inp[3]) ? node1402 : 4'b1101;
																assign node1402 = (inp[4]) ? 4'b1101 : 4'b1001;
										assign node1406 = (inp[13]) ? node1418 : node1407;
											assign node1407 = (inp[3]) ? node1413 : node1408;
												assign node1408 = (inp[10]) ? 4'b0000 : node1409;
													assign node1409 = (inp[7]) ? 4'b1101 : 4'b1000;
												assign node1413 = (inp[4]) ? 4'b0100 : node1414;
													assign node1414 = (inp[7]) ? 4'b0000 : 4'b0100;
											assign node1418 = (inp[3]) ? node1424 : node1419;
												assign node1419 = (inp[10]) ? node1421 : 4'b0000;
													assign node1421 = (inp[4]) ? 4'b1000 : 4'b1101;
												assign node1424 = (inp[4]) ? node1428 : node1425;
													assign node1425 = (inp[7]) ? 4'b1000 : 4'b1100;
													assign node1428 = (inp[10]) ? 4'b1100 : node1429;
														assign node1429 = (inp[7]) ? 4'b1100 : 4'b0100;
									assign node1433 = (inp[14]) ? node1465 : node1434;
										assign node1434 = (inp[13]) ? node1446 : node1435;
											assign node1435 = (inp[10]) ? 4'b0001 : node1436;
												assign node1436 = (inp[12]) ? node1442 : node1437;
													assign node1437 = (inp[7]) ? node1439 : 4'b0001;
														assign node1439 = (inp[3]) ? 4'b0001 : 4'b1101;
													assign node1442 = (inp[4]) ? 4'b1101 : 4'b1001;
											assign node1446 = (inp[3]) ? node1454 : node1447;
												assign node1447 = (inp[10]) ? 4'b1001 : node1448;
													assign node1448 = (inp[12]) ? node1450 : 4'b1001;
														assign node1450 = (inp[7]) ? 4'b1101 : 4'b0001;
												assign node1454 = (inp[4]) ? node1460 : node1455;
													assign node1455 = (inp[7]) ? 4'b1001 : node1456;
														assign node1456 = (inp[12]) ? 4'b0101 : 4'b1101;
													assign node1460 = (inp[10]) ? 4'b1101 : node1461;
														assign node1461 = (inp[12]) ? 4'b0101 : 4'b1101;
										assign node1465 = (inp[11]) ? node1489 : node1466;
											assign node1466 = (inp[3]) ? node1480 : node1467;
												assign node1467 = (inp[7]) ? node1475 : node1468;
													assign node1468 = (inp[12]) ? node1470 : 4'b1000;
														assign node1470 = (inp[13]) ? node1472 : 4'b0000;
															assign node1472 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node1475 = (inp[12]) ? 4'b1101 : node1476;
														assign node1476 = (inp[10]) ? 4'b1000 : 4'b1101;
												assign node1480 = (inp[4]) ? node1482 : 4'b1000;
													assign node1482 = (inp[13]) ? 4'b1100 : node1483;
														assign node1483 = (inp[10]) ? 4'b0100 : node1484;
															assign node1484 = (inp[12]) ? 4'b1100 : 4'b0100;
											assign node1489 = (inp[13]) ? node1497 : node1490;
												assign node1490 = (inp[7]) ? node1492 : 4'b0101;
													assign node1492 = (inp[12]) ? 4'b1001 : node1493;
														assign node1493 = (inp[10]) ? 4'b0001 : 4'b0101;
												assign node1497 = (inp[4]) ? 4'b1101 : node1498;
													assign node1498 = (inp[7]) ? node1502 : node1499;
														assign node1499 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node1502 = (inp[3]) ? 4'b1001 : 4'b1101;
							assign node1507 = (inp[2]) ? 4'b1001 : node1508;
								assign node1508 = (inp[3]) ? node1510 : 4'b1001;
									assign node1510 = (inp[4]) ? node1524 : node1511;
										assign node1511 = (inp[7]) ? 4'b1001 : node1512;
											assign node1512 = (inp[1]) ? node1518 : node1513;
												assign node1513 = (inp[13]) ? node1515 : 4'b0000;
													assign node1515 = (inp[11]) ? 4'b1000 : 4'b1001;
												assign node1518 = (inp[13]) ? 4'b1001 : node1519;
													assign node1519 = (inp[10]) ? 4'b0001 : 4'b1001;
										assign node1524 = (inp[13]) ? node1538 : node1525;
											assign node1525 = (inp[12]) ? node1533 : node1526;
												assign node1526 = (inp[10]) ? node1530 : node1527;
													assign node1527 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node1530 = (inp[11]) ? 4'b0000 : 4'b0001;
												assign node1533 = (inp[10]) ? node1535 : 4'b1001;
													assign node1535 = (inp[11]) ? 4'b0001 : 4'b0000;
											assign node1538 = (inp[1]) ? node1548 : node1539;
												assign node1539 = (inp[12]) ? node1541 : 4'b1000;
													assign node1541 = (inp[10]) ? node1543 : 4'b0000;
														assign node1543 = (inp[11]) ? 4'b1000 : node1544;
															assign node1544 = (inp[14]) ? 4'b0001 : 4'b1000;
												assign node1548 = (inp[10]) ? node1552 : node1549;
													assign node1549 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node1552 = (inp[14]) ? node1554 : 4'b1001;
														assign node1554 = (inp[11]) ? 4'b1001 : 4'b1000;
					assign node1558 = (inp[3]) ? node2120 : node1559;
						assign node1559 = (inp[4]) ? node1833 : node1560;
							assign node1560 = (inp[0]) ? node1726 : node1561;
								assign node1561 = (inp[11]) ? node1653 : node1562;
									assign node1562 = (inp[2]) ? node1620 : node1563;
										assign node1563 = (inp[14]) ? node1591 : node1564;
											assign node1564 = (inp[1]) ? node1582 : node1565;
												assign node1565 = (inp[13]) ? node1577 : node1566;
													assign node1566 = (inp[7]) ? node1574 : node1567;
														assign node1567 = (inp[12]) ? node1569 : 4'b0101;
															assign node1569 = (inp[10]) ? node1571 : 4'b1101;
																assign node1571 = (inp[15]) ? 4'b1101 : 4'b1001;
														assign node1574 = (inp[15]) ? 4'b1001 : 4'b0001;
													assign node1577 = (inp[10]) ? node1579 : 4'b0101;
														assign node1579 = (inp[7]) ? 4'b0101 : 4'b0000;
												assign node1582 = (inp[7]) ? node1586 : node1583;
													assign node1583 = (inp[15]) ? 4'b0100 : 4'b0001;
													assign node1586 = (inp[15]) ? 4'b1100 : node1587;
														assign node1587 = (inp[13]) ? 4'b1001 : 4'b1100;
											assign node1591 = (inp[1]) ? node1603 : node1592;
												assign node1592 = (inp[15]) ? node1596 : node1593;
													assign node1593 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node1596 = (inp[13]) ? 4'b0100 : node1597;
														assign node1597 = (inp[7]) ? 4'b1000 : node1598;
															assign node1598 = (inp[10]) ? 4'b1100 : 4'b1000;
												assign node1603 = (inp[12]) ? node1615 : node1604;
													assign node1604 = (inp[13]) ? node1610 : node1605;
														assign node1605 = (inp[7]) ? node1607 : 4'b1001;
															assign node1607 = (inp[10]) ? 4'b0101 : 4'b0001;
														assign node1610 = (inp[10]) ? node1612 : 4'b1101;
															assign node1612 = (inp[15]) ? 4'b1001 : 4'b1000;
													assign node1615 = (inp[13]) ? node1617 : 4'b0001;
														assign node1617 = (inp[10]) ? 4'b0000 : 4'b0001;
										assign node1620 = (inp[15]) ? node1636 : node1621;
											assign node1621 = (inp[13]) ? node1631 : node1622;
												assign node1622 = (inp[12]) ? node1628 : node1623;
													assign node1623 = (inp[10]) ? node1625 : 4'b0100;
														assign node1625 = (inp[14]) ? 4'b0001 : 4'b0000;
													assign node1628 = (inp[10]) ? 4'b0100 : 4'b1100;
												assign node1631 = (inp[14]) ? node1633 : 4'b0001;
													assign node1633 = (inp[10]) ? 4'b0000 : 4'b1000;
											assign node1636 = (inp[10]) ? node1644 : node1637;
												assign node1637 = (inp[13]) ? 4'b0100 : node1638;
													assign node1638 = (inp[1]) ? 4'b0100 : node1639;
														assign node1639 = (inp[7]) ? 4'b0000 : 4'b1000;
												assign node1644 = (inp[14]) ? node1650 : node1645;
													assign node1645 = (inp[12]) ? 4'b1100 : node1646;
														assign node1646 = (inp[1]) ? 4'b1000 : 4'b1100;
													assign node1650 = (inp[13]) ? 4'b0000 : 4'b1100;
									assign node1653 = (inp[1]) ? node1689 : node1654;
										assign node1654 = (inp[15]) ? node1672 : node1655;
											assign node1655 = (inp[2]) ? node1665 : node1656;
												assign node1656 = (inp[13]) ? node1658 : 4'b0001;
													assign node1658 = (inp[7]) ? node1662 : node1659;
														assign node1659 = (inp[10]) ? 4'b0000 : 4'b0101;
														assign node1662 = (inp[10]) ? 4'b0101 : 4'b0001;
												assign node1665 = (inp[14]) ? node1667 : 4'b0000;
													assign node1667 = (inp[12]) ? node1669 : 4'b1100;
														assign node1669 = (inp[13]) ? 4'b0100 : 4'b0101;
											assign node1672 = (inp[2]) ? node1678 : node1673;
												assign node1673 = (inp[12]) ? 4'b1100 : node1674;
													assign node1674 = (inp[7]) ? 4'b1100 : 4'b0001;
												assign node1678 = (inp[12]) ? node1682 : node1679;
													assign node1679 = (inp[10]) ? 4'b1101 : 4'b0101;
													assign node1682 = (inp[10]) ? node1684 : 4'b1001;
														assign node1684 = (inp[7]) ? node1686 : 4'b0101;
															assign node1686 = (inp[13]) ? 4'b0101 : 4'b0001;
										assign node1689 = (inp[13]) ? node1709 : node1690;
											assign node1690 = (inp[14]) ? node1702 : node1691;
												assign node1691 = (inp[2]) ? node1693 : 4'b0101;
													assign node1693 = (inp[12]) ? node1695 : 4'b0001;
														assign node1695 = (inp[10]) ? 4'b0001 : node1696;
															assign node1696 = (inp[15]) ? node1698 : 4'b0101;
																assign node1698 = (inp[7]) ? 4'b0001 : 4'b0101;
												assign node1702 = (inp[15]) ? node1706 : node1703;
													assign node1703 = (inp[2]) ? 4'b0001 : 4'b1001;
													assign node1706 = (inp[7]) ? 4'b1001 : 4'b1101;
											assign node1709 = (inp[10]) ? node1717 : node1710;
												assign node1710 = (inp[2]) ? node1712 : 4'b1001;
													assign node1712 = (inp[7]) ? node1714 : 4'b0101;
														assign node1714 = (inp[15]) ? 4'b0101 : 4'b1001;
												assign node1717 = (inp[15]) ? node1723 : node1718;
													assign node1718 = (inp[7]) ? node1720 : 4'b1101;
														assign node1720 = (inp[2]) ? 4'b1001 : 4'b1101;
													assign node1723 = (inp[7]) ? 4'b1101 : 4'b1001;
								assign node1726 = (inp[2]) ? node1810 : node1727;
									assign node1727 = (inp[1]) ? node1779 : node1728;
										assign node1728 = (inp[12]) ? node1754 : node1729;
											assign node1729 = (inp[10]) ? node1743 : node1730;
												assign node1730 = (inp[14]) ? node1738 : node1731;
													assign node1731 = (inp[15]) ? 4'b0100 : node1732;
														assign node1732 = (inp[11]) ? 4'b0001 : node1733;
															assign node1733 = (inp[7]) ? 4'b0100 : 4'b0000;
													assign node1738 = (inp[15]) ? node1740 : 4'b0000;
														assign node1740 = (inp[13]) ? 4'b0001 : 4'b1001;
												assign node1743 = (inp[14]) ? node1745 : 4'b1001;
													assign node1745 = (inp[7]) ? 4'b0100 : node1746;
														assign node1746 = (inp[15]) ? node1750 : node1747;
															assign node1747 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node1750 = (inp[11]) ? 4'b1100 : 4'b1101;
											assign node1754 = (inp[7]) ? node1772 : node1755;
												assign node1755 = (inp[10]) ? node1767 : node1756;
													assign node1756 = (inp[14]) ? node1762 : node1757;
														assign node1757 = (inp[13]) ? 4'b0100 : node1758;
															assign node1758 = (inp[11]) ? 4'b1100 : 4'b1000;
														assign node1762 = (inp[13]) ? 4'b1001 : node1763;
															assign node1763 = (inp[11]) ? 4'b1100 : 4'b1101;
													assign node1767 = (inp[13]) ? 4'b1100 : node1768;
														assign node1768 = (inp[15]) ? 4'b0100 : 4'b0000;
												assign node1772 = (inp[15]) ? node1774 : 4'b0100;
													assign node1774 = (inp[13]) ? node1776 : 4'b0000;
														assign node1776 = (inp[10]) ? 4'b1000 : 4'b0000;
										assign node1779 = (inp[10]) ? node1805 : node1780;
											assign node1780 = (inp[11]) ? node1794 : node1781;
												assign node1781 = (inp[14]) ? node1789 : node1782;
													assign node1782 = (inp[15]) ? node1786 : node1783;
														assign node1783 = (inp[13]) ? 4'b0000 : 4'b1101;
														assign node1786 = (inp[12]) ? 4'b1001 : 4'b1101;
													assign node1789 = (inp[15]) ? node1791 : 4'b0000;
														assign node1791 = (inp[13]) ? 4'b0100 : 4'b0000;
												assign node1794 = (inp[12]) ? node1798 : node1795;
													assign node1795 = (inp[15]) ? 4'b0101 : 4'b0001;
													assign node1798 = (inp[13]) ? node1802 : node1799;
														assign node1799 = (inp[15]) ? 4'b1001 : 4'b1101;
														assign node1802 = (inp[7]) ? 4'b0001 : 4'b0101;
											assign node1805 = (inp[11]) ? 4'b1001 : node1806;
												assign node1806 = (inp[15]) ? 4'b1001 : 4'b1000;
									assign node1810 = (inp[15]) ? 4'b1001 : node1811;
										assign node1811 = (inp[7]) ? 4'b1101 : node1812;
											assign node1812 = (inp[13]) ? node1824 : node1813;
												assign node1813 = (inp[10]) ? node1815 : 4'b1101;
													assign node1815 = (inp[1]) ? 4'b0001 : node1816;
														assign node1816 = (inp[12]) ? node1818 : 4'b0001;
															assign node1818 = (inp[11]) ? 4'b0000 : node1819;
																assign node1819 = (inp[14]) ? 4'b1101 : 4'b0000;
												assign node1824 = (inp[1]) ? 4'b1001 : node1825;
													assign node1825 = (inp[10]) ? 4'b1000 : node1826;
														assign node1826 = (inp[12]) ? 4'b0000 : 4'b1000;
							assign node1833 = (inp[2]) ? node2007 : node1834;
								assign node1834 = (inp[11]) ? node1938 : node1835;
									assign node1835 = (inp[0]) ? node1887 : node1836;
										assign node1836 = (inp[13]) ? node1866 : node1837;
											assign node1837 = (inp[10]) ? node1851 : node1838;
												assign node1838 = (inp[15]) ? node1844 : node1839;
													assign node1839 = (inp[1]) ? node1841 : 4'b0000;
														assign node1841 = (inp[14]) ? 4'b1000 : 4'b1001;
													assign node1844 = (inp[7]) ? node1846 : 4'b0101;
														assign node1846 = (inp[14]) ? 4'b1001 : node1847;
															assign node1847 = (inp[1]) ? 4'b0001 : 4'b1001;
												assign node1851 = (inp[7]) ? node1859 : node1852;
													assign node1852 = (inp[15]) ? node1854 : 4'b1100;
														assign node1854 = (inp[12]) ? 4'b0000 : node1855;
															assign node1855 = (inp[1]) ? 4'b0000 : 4'b0001;
													assign node1859 = (inp[15]) ? node1861 : 4'b0001;
														assign node1861 = (inp[1]) ? node1863 : 4'b0101;
															assign node1863 = (inp[12]) ? 4'b0101 : 4'b0000;
											assign node1866 = (inp[1]) ? node1876 : node1867;
												assign node1867 = (inp[10]) ? node1873 : node1868;
													assign node1868 = (inp[14]) ? 4'b0001 : node1869;
														assign node1869 = (inp[15]) ? 4'b1000 : 4'b0000;
													assign node1873 = (inp[12]) ? 4'b1000 : 4'b0100;
												assign node1876 = (inp[12]) ? node1878 : 4'b0000;
													assign node1878 = (inp[10]) ? node1884 : node1879;
														assign node1879 = (inp[7]) ? 4'b0001 : node1880;
															assign node1880 = (inp[14]) ? 4'b0100 : 4'b0101;
														assign node1884 = (inp[14]) ? 4'b0001 : 4'b0000;
										assign node1887 = (inp[13]) ? node1913 : node1888;
											assign node1888 = (inp[12]) ? node1894 : node1889;
												assign node1889 = (inp[15]) ? 4'b0101 : node1890;
													assign node1890 = (inp[7]) ? 4'b0000 : 4'b0100;
												assign node1894 = (inp[10]) ? node1904 : node1895;
													assign node1895 = (inp[7]) ? node1897 : 4'b0100;
														assign node1897 = (inp[15]) ? node1901 : node1898;
															assign node1898 = (inp[1]) ? 4'b0000 : 4'b1000;
															assign node1901 = (inp[1]) ? 4'b1001 : 4'b1000;
													assign node1904 = (inp[7]) ? 4'b0100 : node1905;
														assign node1905 = (inp[15]) ? 4'b0000 : node1906;
															assign node1906 = (inp[14]) ? 4'b1100 : node1907;
																assign node1907 = (inp[1]) ? 4'b0000 : 4'b0100;
											assign node1913 = (inp[10]) ? node1933 : node1914;
												assign node1914 = (inp[7]) ? node1924 : node1915;
													assign node1915 = (inp[1]) ? node1919 : node1916;
														assign node1916 = (inp[14]) ? 4'b0000 : 4'b1001;
														assign node1919 = (inp[14]) ? 4'b1001 : node1920;
															assign node1920 = (inp[12]) ? 4'b1000 : 4'b0000;
													assign node1924 = (inp[1]) ? 4'b0000 : node1925;
														assign node1925 = (inp[14]) ? node1929 : node1926;
															assign node1926 = (inp[12]) ? 4'b0100 : 4'b0000;
															assign node1929 = (inp[15]) ? 4'b0101 : 4'b0100;
												assign node1933 = (inp[15]) ? 4'b1000 : node1934;
													assign node1934 = (inp[12]) ? 4'b0001 : 4'b1001;
									assign node1938 = (inp[1]) ? node1982 : node1939;
										assign node1939 = (inp[15]) ? node1961 : node1940;
											assign node1940 = (inp[7]) ? node1952 : node1941;
												assign node1941 = (inp[0]) ? node1943 : 4'b1000;
													assign node1943 = (inp[13]) ? node1949 : node1944;
														assign node1944 = (inp[12]) ? 4'b0101 : node1945;
															assign node1945 = (inp[10]) ? 4'b0000 : 4'b0101;
														assign node1949 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node1952 = (inp[0]) ? 4'b1001 : node1953;
													assign node1953 = (inp[13]) ? node1957 : node1954;
														assign node1954 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node1957 = (inp[10]) ? 4'b1001 : 4'b0001;
											assign node1961 = (inp[0]) ? node1975 : node1962;
												assign node1962 = (inp[14]) ? node1970 : node1963;
													assign node1963 = (inp[7]) ? node1967 : node1964;
														assign node1964 = (inp[13]) ? 4'b1001 : 4'b1000;
														assign node1967 = (inp[10]) ? 4'b0101 : 4'b0000;
													assign node1970 = (inp[7]) ? node1972 : 4'b0101;
														assign node1972 = (inp[10]) ? 4'b0101 : 4'b0001;
												assign node1975 = (inp[13]) ? node1977 : 4'b0001;
													assign node1977 = (inp[7]) ? 4'b0001 : node1978;
														assign node1978 = (inp[14]) ? 4'b1001 : 4'b0001;
										assign node1982 = (inp[10]) ? node1996 : node1983;
											assign node1983 = (inp[15]) ? 4'b0001 : node1984;
												assign node1984 = (inp[12]) ? node1990 : node1985;
													assign node1985 = (inp[7]) ? 4'b0001 : node1986;
														assign node1986 = (inp[13]) ? 4'b0001 : 4'b0101;
													assign node1990 = (inp[0]) ? 4'b0101 : node1991;
														assign node1991 = (inp[13]) ? 4'b0001 : 4'b1001;
											assign node1996 = (inp[13]) ? 4'b1001 : node1997;
												assign node1997 = (inp[0]) ? node1999 : 4'b0101;
													assign node1999 = (inp[7]) ? node2003 : node2000;
														assign node2000 = (inp[15]) ? 4'b1001 : 4'b0001;
														assign node2003 = (inp[15]) ? 4'b0101 : 4'b1001;
								assign node2007 = (inp[15]) ? node2081 : node2008;
									assign node2008 = (inp[1]) ? node2048 : node2009;
										assign node2009 = (inp[0]) ? node2031 : node2010;
											assign node2010 = (inp[11]) ? node2020 : node2011;
												assign node2011 = (inp[12]) ? node2017 : node2012;
													assign node2012 = (inp[10]) ? 4'b0001 : node2013;
														assign node2013 = (inp[14]) ? 4'b0100 : 4'b0101;
													assign node2017 = (inp[14]) ? 4'b1100 : 4'b1101;
												assign node2020 = (inp[10]) ? node2028 : node2021;
													assign node2021 = (inp[13]) ? node2023 : 4'b0100;
														assign node2023 = (inp[12]) ? node2025 : 4'b0000;
															assign node2025 = (inp[7]) ? 4'b0001 : 4'b0101;
													assign node2028 = (inp[13]) ? 4'b0000 : 4'b0001;
											assign node2031 = (inp[10]) ? node2043 : node2032;
												assign node2032 = (inp[11]) ? node2038 : node2033;
													assign node2033 = (inp[7]) ? 4'b1101 : node2034;
														assign node2034 = (inp[13]) ? 4'b0001 : 4'b1000;
													assign node2038 = (inp[12]) ? node2040 : 4'b0000;
														assign node2040 = (inp[13]) ? 4'b0000 : 4'b1101;
												assign node2043 = (inp[13]) ? node2045 : 4'b0000;
													assign node2045 = (inp[7]) ? 4'b1000 : 4'b1001;
										assign node2048 = (inp[11]) ? node2064 : node2049;
											assign node2049 = (inp[14]) ? node2057 : node2050;
												assign node2050 = (inp[10]) ? node2052 : 4'b0100;
													assign node2052 = (inp[13]) ? node2054 : 4'b0001;
														assign node2054 = (inp[0]) ? 4'b1001 : 4'b0001;
												assign node2057 = (inp[0]) ? node2061 : node2058;
													assign node2058 = (inp[13]) ? 4'b0000 : 4'b0001;
													assign node2061 = (inp[12]) ? 4'b1000 : 4'b0000;
											assign node2064 = (inp[0]) ? node2070 : node2065;
												assign node2065 = (inp[10]) ? 4'b1001 : node2066;
													assign node2066 = (inp[12]) ? 4'b0101 : 4'b1101;
												assign node2070 = (inp[13]) ? node2076 : node2071;
													assign node2071 = (inp[10]) ? 4'b0001 : node2072;
														assign node2072 = (inp[14]) ? 4'b1001 : 4'b0001;
													assign node2076 = (inp[10]) ? 4'b1001 : node2077;
														assign node2077 = (inp[12]) ? 4'b0001 : 4'b1001;
									assign node2081 = (inp[0]) ? 4'b1001 : node2082;
										assign node2082 = (inp[1]) ? node2104 : node2083;
											assign node2083 = (inp[11]) ? node2099 : node2084;
												assign node2084 = (inp[12]) ? node2094 : node2085;
													assign node2085 = (inp[14]) ? 4'b0001 : node2086;
														assign node2086 = (inp[10]) ? 4'b1001 : node2087;
															assign node2087 = (inp[13]) ? node2089 : 4'b0001;
																assign node2089 = (inp[7]) ? 4'b1001 : 4'b0001;
													assign node2094 = (inp[13]) ? 4'b0000 : node2095;
														assign node2095 = (inp[10]) ? 4'b1001 : 4'b1100;
												assign node2099 = (inp[10]) ? 4'b1000 : node2100;
													assign node2100 = (inp[13]) ? 4'b1000 : 4'b0000;
											assign node2104 = (inp[11]) ? node2114 : node2105;
												assign node2105 = (inp[7]) ? node2109 : node2106;
													assign node2106 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node2109 = (inp[13]) ? node2111 : 4'b0001;
														assign node2111 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node2114 = (inp[13]) ? 4'b1001 : node2115;
													assign node2115 = (inp[10]) ? 4'b0101 : 4'b1001;
						assign node2120 = (inp[4]) ? node2440 : node2121;
							assign node2121 = (inp[1]) ? node2297 : node2122;
								assign node2122 = (inp[15]) ? node2202 : node2123;
									assign node2123 = (inp[11]) ? node2165 : node2124;
										assign node2124 = (inp[2]) ? node2154 : node2125;
											assign node2125 = (inp[0]) ? node2137 : node2126;
												assign node2126 = (inp[12]) ? node2130 : node2127;
													assign node2127 = (inp[13]) ? 4'b1001 : 4'b1000;
													assign node2130 = (inp[13]) ? 4'b0000 : node2131;
														assign node2131 = (inp[14]) ? node2133 : 4'b0001;
															assign node2133 = (inp[7]) ? 4'b0000 : 4'b0001;
												assign node2137 = (inp[12]) ? node2149 : node2138;
													assign node2138 = (inp[13]) ? node2144 : node2139;
														assign node2139 = (inp[7]) ? node2141 : 4'b0001;
															assign node2141 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node2144 = (inp[10]) ? node2146 : 4'b1001;
															assign node2146 = (inp[7]) ? 4'b1001 : 4'b1000;
													assign node2149 = (inp[10]) ? node2151 : 4'b1000;
														assign node2151 = (inp[13]) ? 4'b1000 : 4'b1001;
											assign node2154 = (inp[12]) ? node2162 : node2155;
												assign node2155 = (inp[10]) ? node2157 : 4'b0000;
													assign node2157 = (inp[7]) ? node2159 : 4'b0000;
														assign node2159 = (inp[0]) ? 4'b1000 : 4'b0000;
												assign node2162 = (inp[13]) ? 4'b0000 : 4'b1000;
										assign node2165 = (inp[2]) ? node2181 : node2166;
											assign node2166 = (inp[0]) ? node2170 : node2167;
												assign node2167 = (inp[10]) ? 4'b0000 : 4'b1000;
												assign node2170 = (inp[13]) ? node2176 : node2171;
													assign node2171 = (inp[14]) ? node2173 : 4'b0001;
														assign node2173 = (inp[10]) ? 4'b0001 : 4'b0000;
													assign node2176 = (inp[12]) ? node2178 : 4'b0000;
														assign node2178 = (inp[7]) ? 4'b0000 : 4'b1000;
											assign node2181 = (inp[12]) ? node2197 : node2182;
												assign node2182 = (inp[10]) ? node2190 : node2183;
													assign node2183 = (inp[7]) ? node2187 : node2184;
														assign node2184 = (inp[0]) ? 4'b0001 : 4'b1001;
														assign node2187 = (inp[0]) ? 4'b0001 : 4'b0000;
													assign node2190 = (inp[0]) ? node2192 : 4'b1000;
														assign node2192 = (inp[7]) ? node2194 : 4'b1001;
															assign node2194 = (inp[13]) ? 4'b1001 : 4'b0000;
												assign node2197 = (inp[10]) ? 4'b0001 : node2198;
													assign node2198 = (inp[0]) ? 4'b1000 : 4'b0001;
									assign node2202 = (inp[11]) ? node2246 : node2203;
										assign node2203 = (inp[0]) ? node2225 : node2204;
											assign node2204 = (inp[7]) ? node2218 : node2205;
												assign node2205 = (inp[10]) ? node2211 : node2206;
													assign node2206 = (inp[2]) ? 4'b0000 : node2207;
														assign node2207 = (inp[13]) ? 4'b0000 : 4'b0001;
													assign node2211 = (inp[14]) ? 4'b0001 : node2212;
														assign node2212 = (inp[12]) ? 4'b0001 : node2213;
															assign node2213 = (inp[13]) ? 4'b1001 : 4'b1000;
												assign node2218 = (inp[13]) ? node2220 : 4'b0000;
													assign node2220 = (inp[10]) ? 4'b0000 : node2221;
														assign node2221 = (inp[14]) ? 4'b0001 : 4'b0000;
											assign node2225 = (inp[2]) ? node2243 : node2226;
												assign node2226 = (inp[14]) ? node2238 : node2227;
													assign node2227 = (inp[13]) ? node2233 : node2228;
														assign node2228 = (inp[12]) ? node2230 : 4'b0001;
															assign node2230 = (inp[10]) ? 4'b1001 : 4'b1000;
														assign node2233 = (inp[7]) ? 4'b0001 : node2234;
															assign node2234 = (inp[10]) ? 4'b0000 : 4'b0001;
													assign node2238 = (inp[12]) ? 4'b1000 : node2239;
														assign node2239 = (inp[13]) ? 4'b1000 : 4'b0000;
												assign node2243 = (inp[7]) ? 4'b1001 : 4'b0001;
										assign node2246 = (inp[0]) ? node2280 : node2247;
											assign node2247 = (inp[7]) ? node2263 : node2248;
												assign node2248 = (inp[10]) ? node2250 : 4'b1000;
													assign node2250 = (inp[12]) ? node2260 : node2251;
														assign node2251 = (inp[14]) ? node2255 : node2252;
															assign node2252 = (inp[13]) ? 4'b0001 : 4'b1001;
															assign node2255 = (inp[13]) ? 4'b1001 : node2256;
																assign node2256 = (inp[2]) ? 4'b0001 : 4'b1001;
														assign node2260 = (inp[13]) ? 4'b1001 : 4'b1000;
												assign node2263 = (inp[10]) ? node2273 : node2264;
													assign node2264 = (inp[12]) ? node2270 : node2265;
														assign node2265 = (inp[13]) ? node2267 : 4'b1001;
															assign node2267 = (inp[2]) ? 4'b1001 : 4'b1000;
														assign node2270 = (inp[2]) ? 4'b0001 : 4'b0000;
													assign node2273 = (inp[13]) ? node2275 : 4'b1000;
														assign node2275 = (inp[12]) ? 4'b1000 : node2276;
															assign node2276 = (inp[2]) ? 4'b0000 : 4'b1000;
											assign node2280 = (inp[7]) ? node2290 : node2281;
												assign node2281 = (inp[12]) ? node2283 : 4'b0000;
													assign node2283 = (inp[13]) ? node2287 : node2284;
														assign node2284 = (inp[10]) ? 4'b0000 : 4'b1001;
														assign node2287 = (inp[10]) ? 4'b1000 : 4'b0000;
												assign node2290 = (inp[2]) ? 4'b1001 : node2291;
													assign node2291 = (inp[10]) ? 4'b0001 : node2292;
														assign node2292 = (inp[13]) ? 4'b1000 : 4'b0001;
								assign node2297 = (inp[11]) ? node2389 : node2298;
									assign node2298 = (inp[14]) ? node2342 : node2299;
										assign node2299 = (inp[0]) ? node2329 : node2300;
											assign node2300 = (inp[12]) ? node2318 : node2301;
												assign node2301 = (inp[13]) ? node2307 : node2302;
													assign node2302 = (inp[10]) ? node2304 : 4'b0000;
														assign node2304 = (inp[2]) ? 4'b1000 : 4'b0001;
													assign node2307 = (inp[7]) ? node2309 : 4'b0001;
														assign node2309 = (inp[10]) ? node2315 : node2310;
															assign node2310 = (inp[15]) ? node2312 : 4'b0001;
																assign node2312 = (inp[2]) ? 4'b0000 : 4'b0001;
															assign node2315 = (inp[15]) ? 4'b0001 : 4'b0000;
												assign node2318 = (inp[2]) ? node2322 : node2319;
													assign node2319 = (inp[7]) ? 4'b1001 : 4'b1000;
													assign node2322 = (inp[10]) ? node2324 : 4'b1000;
														assign node2324 = (inp[15]) ? node2326 : 4'b0000;
															assign node2326 = (inp[13]) ? 4'b0001 : 4'b0000;
											assign node2329 = (inp[15]) ? 4'b1001 : node2330;
												assign node2330 = (inp[2]) ? node2336 : node2331;
													assign node2331 = (inp[12]) ? 4'b0001 : node2332;
														assign node2332 = (inp[10]) ? 4'b0001 : 4'b1001;
													assign node2336 = (inp[13]) ? 4'b1000 : node2337;
														assign node2337 = (inp[7]) ? 4'b0001 : 4'b0000;
										assign node2342 = (inp[12]) ? node2358 : node2343;
											assign node2343 = (inp[15]) ? node2353 : node2344;
												assign node2344 = (inp[0]) ? 4'b0000 : node2345;
													assign node2345 = (inp[13]) ? node2349 : node2346;
														assign node2346 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node2349 = (inp[2]) ? 4'b0001 : 4'b0000;
												assign node2353 = (inp[10]) ? node2355 : 4'b1001;
													assign node2355 = (inp[7]) ? 4'b0001 : 4'b0000;
											assign node2358 = (inp[0]) ? node2368 : node2359;
												assign node2359 = (inp[15]) ? node2365 : node2360;
													assign node2360 = (inp[10]) ? node2362 : 4'b0001;
														assign node2362 = (inp[13]) ? 4'b1000 : 4'b1001;
													assign node2365 = (inp[2]) ? 4'b0000 : 4'b1000;
												assign node2368 = (inp[2]) ? node2380 : node2369;
													assign node2369 = (inp[10]) ? node2375 : node2370;
														assign node2370 = (inp[13]) ? 4'b0000 : node2371;
															assign node2371 = (inp[15]) ? 4'b0000 : 4'b0001;
														assign node2375 = (inp[15]) ? node2377 : 4'b0001;
															assign node2377 = (inp[7]) ? 4'b0001 : 4'b0000;
													assign node2380 = (inp[15]) ? 4'b1001 : node2381;
														assign node2381 = (inp[13]) ? 4'b0000 : node2382;
															assign node2382 = (inp[10]) ? 4'b0000 : node2383;
																assign node2383 = (inp[7]) ? 4'b1000 : 4'b0000;
									assign node2389 = (inp[13]) ? node2417 : node2390;
										assign node2390 = (inp[0]) ? node2402 : node2391;
											assign node2391 = (inp[12]) ? node2395 : node2392;
												assign node2392 = (inp[10]) ? 4'b1001 : 4'b0001;
												assign node2395 = (inp[10]) ? 4'b0001 : node2396;
													assign node2396 = (inp[15]) ? node2398 : 4'b1001;
														assign node2398 = (inp[14]) ? 4'b0001 : 4'b1001;
											assign node2402 = (inp[2]) ? node2408 : node2403;
												assign node2403 = (inp[10]) ? 4'b0001 : node2404;
													assign node2404 = (inp[7]) ? 4'b0001 : 4'b1001;
												assign node2408 = (inp[12]) ? node2414 : node2409;
													assign node2409 = (inp[14]) ? 4'b0001 : node2410;
														assign node2410 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node2414 = (inp[14]) ? 4'b1001 : 4'b0001;
										assign node2417 = (inp[10]) ? 4'b1001 : node2418;
											assign node2418 = (inp[0]) ? node2428 : node2419;
												assign node2419 = (inp[15]) ? 4'b0001 : node2420;
													assign node2420 = (inp[2]) ? 4'b0001 : node2421;
														assign node2421 = (inp[12]) ? 4'b1001 : node2422;
															assign node2422 = (inp[14]) ? 4'b0001 : 4'b1001;
												assign node2428 = (inp[15]) ? node2434 : node2429;
													assign node2429 = (inp[12]) ? 4'b0001 : node2430;
														assign node2430 = (inp[2]) ? 4'b0001 : 4'b1001;
													assign node2434 = (inp[2]) ? 4'b1001 : node2435;
														assign node2435 = (inp[7]) ? 4'b0001 : 4'b1001;
							assign node2440 = (inp[13]) ? node2596 : node2441;
								assign node2441 = (inp[1]) ? node2541 : node2442;
									assign node2442 = (inp[2]) ? node2498 : node2443;
										assign node2443 = (inp[7]) ? node2479 : node2444;
											assign node2444 = (inp[12]) ? node2462 : node2445;
												assign node2445 = (inp[11]) ? node2453 : node2446;
													assign node2446 = (inp[14]) ? node2448 : 4'b0001;
														assign node2448 = (inp[10]) ? 4'b0000 : node2449;
															assign node2449 = (inp[15]) ? 4'b0000 : 4'b0001;
													assign node2453 = (inp[10]) ? node2457 : node2454;
														assign node2454 = (inp[15]) ? 4'b1001 : 4'b0001;
														assign node2457 = (inp[15]) ? node2459 : 4'b0001;
															assign node2459 = (inp[14]) ? 4'b0001 : 4'b0000;
												assign node2462 = (inp[0]) ? node2468 : node2463;
													assign node2463 = (inp[15]) ? node2465 : 4'b1000;
														assign node2465 = (inp[14]) ? 4'b1000 : 4'b1001;
													assign node2468 = (inp[15]) ? node2474 : node2469;
														assign node2469 = (inp[10]) ? node2471 : 4'b1001;
															assign node2471 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node2474 = (inp[11]) ? 4'b0000 : node2475;
															assign node2475 = (inp[10]) ? 4'b0001 : 4'b0000;
											assign node2479 = (inp[12]) ? node2489 : node2480;
												assign node2480 = (inp[0]) ? node2482 : 4'b1000;
													assign node2482 = (inp[11]) ? 4'b1000 : node2483;
														assign node2483 = (inp[15]) ? node2485 : 4'b0001;
															assign node2485 = (inp[10]) ? 4'b0001 : 4'b0000;
												assign node2489 = (inp[10]) ? 4'b0000 : node2490;
													assign node2490 = (inp[14]) ? node2494 : node2491;
														assign node2491 = (inp[15]) ? 4'b0001 : 4'b1001;
														assign node2494 = (inp[11]) ? 4'b1000 : 4'b1001;
										assign node2498 = (inp[12]) ? node2518 : node2499;
											assign node2499 = (inp[11]) ? node2509 : node2500;
												assign node2500 = (inp[0]) ? node2506 : node2501;
													assign node2501 = (inp[15]) ? node2503 : 4'b1000;
														assign node2503 = (inp[10]) ? 4'b0000 : 4'b0001;
													assign node2506 = (inp[15]) ? 4'b1000 : 4'b0001;
												assign node2509 = (inp[15]) ? 4'b0001 : node2510;
													assign node2510 = (inp[14]) ? node2512 : 4'b0000;
														assign node2512 = (inp[0]) ? 4'b0001 : node2513;
															assign node2513 = (inp[10]) ? 4'b0000 : 4'b0001;
											assign node2518 = (inp[11]) ? node2526 : node2519;
												assign node2519 = (inp[0]) ? node2523 : node2520;
													assign node2520 = (inp[7]) ? 4'b0001 : 4'b1001;
													assign node2523 = (inp[14]) ? 4'b0001 : 4'b0000;
												assign node2526 = (inp[15]) ? node2536 : node2527;
													assign node2527 = (inp[10]) ? node2533 : node2528;
														assign node2528 = (inp[7]) ? node2530 : 4'b0001;
															assign node2530 = (inp[0]) ? 4'b0000 : 4'b0001;
														assign node2533 = (inp[14]) ? 4'b0000 : 4'b1000;
													assign node2536 = (inp[7]) ? 4'b1000 : node2537;
														assign node2537 = (inp[0]) ? 4'b1000 : 4'b0000;
									assign node2541 = (inp[11]) ? node2581 : node2542;
										assign node2542 = (inp[7]) ? node2562 : node2543;
											assign node2543 = (inp[2]) ? node2553 : node2544;
												assign node2544 = (inp[10]) ? 4'b0001 : node2545;
													assign node2545 = (inp[15]) ? node2547 : 4'b0001;
														assign node2547 = (inp[14]) ? node2549 : 4'b0000;
															assign node2549 = (inp[12]) ? 4'b1001 : 4'b0000;
												assign node2553 = (inp[0]) ? 4'b0001 : node2554;
													assign node2554 = (inp[12]) ? 4'b0000 : node2555;
														assign node2555 = (inp[15]) ? 4'b0001 : node2556;
															assign node2556 = (inp[14]) ? 4'b0000 : 4'b0001;
											assign node2562 = (inp[2]) ? node2568 : node2563;
												assign node2563 = (inp[0]) ? node2565 : 4'b0000;
													assign node2565 = (inp[12]) ? 4'b0001 : 4'b0000;
												assign node2568 = (inp[12]) ? node2578 : node2569;
													assign node2569 = (inp[0]) ? 4'b0000 : node2570;
														assign node2570 = (inp[15]) ? 4'b0001 : node2571;
															assign node2571 = (inp[10]) ? 4'b0000 : node2572;
																assign node2572 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node2578 = (inp[10]) ? 4'b0001 : 4'b1001;
										assign node2581 = (inp[10]) ? 4'b0001 : node2582;
											assign node2582 = (inp[14]) ? node2590 : node2583;
												assign node2583 = (inp[15]) ? 4'b1001 : node2584;
													assign node2584 = (inp[2]) ? 4'b0001 : node2585;
														assign node2585 = (inp[12]) ? 4'b1001 : 4'b0001;
												assign node2590 = (inp[15]) ? 4'b0001 : node2591;
													assign node2591 = (inp[12]) ? 4'b1001 : 4'b0001;
								assign node2596 = (inp[10]) ? node2636 : node2597;
									assign node2597 = (inp[11]) ? node2615 : node2598;
										assign node2598 = (inp[15]) ? node2610 : node2599;
											assign node2599 = (inp[0]) ? node2605 : node2600;
												assign node2600 = (inp[12]) ? node2602 : 4'b0000;
													assign node2602 = (inp[1]) ? 4'b0000 : 4'b0001;
												assign node2605 = (inp[14]) ? node2607 : 4'b0001;
													assign node2607 = (inp[2]) ? 4'b0001 : 4'b0000;
											assign node2610 = (inp[7]) ? node2612 : 4'b0000;
												assign node2612 = (inp[0]) ? 4'b0000 : 4'b0001;
										assign node2615 = (inp[1]) ? 4'b0001 : node2616;
											assign node2616 = (inp[14]) ? node2628 : node2617;
												assign node2617 = (inp[15]) ? node2623 : node2618;
													assign node2618 = (inp[12]) ? node2620 : 4'b0001;
														assign node2620 = (inp[7]) ? 4'b0001 : 4'b0000;
													assign node2623 = (inp[0]) ? node2625 : 4'b0000;
														assign node2625 = (inp[12]) ? 4'b0001 : 4'b0000;
												assign node2628 = (inp[7]) ? 4'b0000 : node2629;
													assign node2629 = (inp[2]) ? node2631 : 4'b0000;
														assign node2631 = (inp[15]) ? 4'b0001 : 4'b0000;
									assign node2636 = (inp[15]) ? node2638 : 4'b0000;
										assign node2638 = (inp[14]) ? 4'b0000 : node2639;
											assign node2639 = (inp[7]) ? node2641 : 4'b0000;
												assign node2641 = (inp[11]) ? 4'b0000 : 4'b0001;
			assign node2645 = (inp[15]) ? node4049 : node2646;
				assign node2646 = (inp[6]) ? node3022 : node2647;
					assign node2647 = (inp[0]) ? 4'b0101 : node2648;
						assign node2648 = (inp[5]) ? node2780 : node2649;
							assign node2649 = (inp[2]) ? 4'b0111 : node2650;
								assign node2650 = (inp[3]) ? node2706 : node2651;
									assign node2651 = (inp[4]) ? node2663 : node2652;
										assign node2652 = (inp[7]) ? 4'b0111 : node2653;
											assign node2653 = (inp[13]) ? node2655 : 4'b0111;
												assign node2655 = (inp[12]) ? 4'b0111 : node2656;
													assign node2656 = (inp[10]) ? 4'b0000 : node2657;
														assign node2657 = (inp[14]) ? 4'b0111 : 4'b0000;
										assign node2663 = (inp[7]) ? node2689 : node2664;
											assign node2664 = (inp[1]) ? node2678 : node2665;
												assign node2665 = (inp[11]) ? node2671 : node2666;
													assign node2666 = (inp[14]) ? node2668 : 4'b1000;
														assign node2668 = (inp[13]) ? 4'b1001 : 4'b0001;
													assign node2671 = (inp[12]) ? node2673 : 4'b1000;
														assign node2673 = (inp[13]) ? node2675 : 4'b0000;
															assign node2675 = (inp[10]) ? 4'b0000 : 4'b1000;
												assign node2678 = (inp[14]) ? node2684 : node2679;
													assign node2679 = (inp[10]) ? node2681 : 4'b1001;
														assign node2681 = (inp[13]) ? 4'b0001 : 4'b1001;
													assign node2684 = (inp[10]) ? node2686 : 4'b0000;
														assign node2686 = (inp[12]) ? 4'b1001 : 4'b1000;
											assign node2689 = (inp[13]) ? node2691 : 4'b0111;
												assign node2691 = (inp[10]) ? node2697 : node2692;
													assign node2692 = (inp[12]) ? 4'b0111 : node2693;
														assign node2693 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node2697 = (inp[11]) ? 4'b0001 : node2698;
														assign node2698 = (inp[12]) ? node2702 : node2699;
															assign node2699 = (inp[1]) ? 4'b0000 : 4'b0001;
															assign node2702 = (inp[1]) ? 4'b0001 : 4'b0000;
									assign node2706 = (inp[13]) ? node2740 : node2707;
										assign node2707 = (inp[1]) ? node2721 : node2708;
											assign node2708 = (inp[14]) ? node2716 : node2709;
												assign node2709 = (inp[11]) ? node2711 : 4'b1000;
													assign node2711 = (inp[10]) ? node2713 : 4'b0000;
														assign node2713 = (inp[4]) ? 4'b1100 : 4'b1000;
												assign node2716 = (inp[11]) ? node2718 : 4'b0001;
													assign node2718 = (inp[12]) ? 4'b0000 : 4'b1000;
											assign node2721 = (inp[14]) ? node2727 : node2722;
												assign node2722 = (inp[4]) ? node2724 : 4'b1001;
													assign node2724 = (inp[7]) ? 4'b1001 : 4'b1101;
												assign node2727 = (inp[11]) ? node2731 : node2728;
													assign node2728 = (inp[4]) ? 4'b1000 : 4'b0000;
													assign node2731 = (inp[4]) ? node2737 : node2732;
														assign node2732 = (inp[12]) ? node2734 : 4'b1001;
															assign node2734 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node2737 = (inp[7]) ? 4'b0001 : 4'b0101;
										assign node2740 = (inp[7]) ? node2752 : node2741;
											assign node2741 = (inp[1]) ? node2747 : node2742;
												assign node2742 = (inp[12]) ? node2744 : 4'b0100;
													assign node2744 = (inp[11]) ? 4'b1100 : 4'b1101;
												assign node2747 = (inp[14]) ? node2749 : 4'b0101;
													assign node2749 = (inp[11]) ? 4'b0101 : 4'b0100;
											assign node2752 = (inp[4]) ? node2766 : node2753;
												assign node2753 = (inp[12]) ? node2759 : node2754;
													assign node2754 = (inp[11]) ? 4'b0001 : node2755;
														assign node2755 = (inp[1]) ? 4'b0000 : 4'b0001;
													assign node2759 = (inp[10]) ? 4'b0000 : node2760;
														assign node2760 = (inp[1]) ? 4'b1000 : node2761;
															assign node2761 = (inp[14]) ? 4'b1001 : 4'b1000;
												assign node2766 = (inp[12]) ? node2772 : node2767;
													assign node2767 = (inp[14]) ? node2769 : 4'b0101;
														assign node2769 = (inp[11]) ? 4'b0101 : 4'b0100;
													assign node2772 = (inp[14]) ? node2774 : 4'b0100;
														assign node2774 = (inp[11]) ? 4'b0100 : node2775;
															assign node2775 = (inp[1]) ? 4'b0100 : 4'b1001;
							assign node2780 = (inp[1]) ? node2896 : node2781;
								assign node2781 = (inp[3]) ? node2845 : node2782;
									assign node2782 = (inp[2]) ? node2818 : node2783;
										assign node2783 = (inp[11]) ? node2807 : node2784;
											assign node2784 = (inp[14]) ? node2796 : node2785;
												assign node2785 = (inp[7]) ? node2791 : node2786;
													assign node2786 = (inp[4]) ? node2788 : 4'b1100;
														assign node2788 = (inp[12]) ? 4'b1000 : 4'b0000;
													assign node2791 = (inp[4]) ? 4'b1100 : node2792;
														assign node2792 = (inp[13]) ? 4'b1100 : 4'b0100;
												assign node2796 = (inp[4]) ? node2804 : node2797;
													assign node2797 = (inp[10]) ? node2801 : node2798;
														assign node2798 = (inp[13]) ? 4'b1101 : 4'b0101;
														assign node2801 = (inp[7]) ? 4'b0101 : 4'b0001;
													assign node2804 = (inp[7]) ? 4'b1101 : 4'b1001;
											assign node2807 = (inp[13]) ? node2813 : node2808;
												assign node2808 = (inp[4]) ? node2810 : 4'b1100;
													assign node2810 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node2813 = (inp[10]) ? 4'b0000 : node2814;
													assign node2814 = (inp[12]) ? 4'b1100 : 4'b0000;
										assign node2818 = (inp[4]) ? node2828 : node2819;
											assign node2819 = (inp[11]) ? node2821 : 4'b0111;
												assign node2821 = (inp[13]) ? node2823 : 4'b0111;
													assign node2823 = (inp[10]) ? node2825 : 4'b0111;
														assign node2825 = (inp[7]) ? 4'b0111 : 4'b0000;
											assign node2828 = (inp[7]) ? node2840 : node2829;
												assign node2829 = (inp[14]) ? node2837 : node2830;
													assign node2830 = (inp[11]) ? node2832 : 4'b0000;
														assign node2832 = (inp[13]) ? node2834 : 4'b1000;
															assign node2834 = (inp[12]) ? 4'b1000 : 4'b0000;
													assign node2837 = (inp[11]) ? 4'b1000 : 4'b1001;
												assign node2840 = (inp[10]) ? node2842 : 4'b0111;
													assign node2842 = (inp[13]) ? 4'b0000 : 4'b0111;
									assign node2845 = (inp[11]) ? node2869 : node2846;
										assign node2846 = (inp[14]) ? node2856 : node2847;
											assign node2847 = (inp[13]) ? node2849 : 4'b1000;
												assign node2849 = (inp[4]) ? 4'b0100 : node2850;
													assign node2850 = (inp[10]) ? 4'b0100 : node2851;
														assign node2851 = (inp[12]) ? 4'b1000 : 4'b0000;
											assign node2856 = (inp[7]) ? node2862 : node2857;
												assign node2857 = (inp[4]) ? 4'b0101 : node2858;
													assign node2858 = (inp[13]) ? 4'b1001 : 4'b0001;
												assign node2862 = (inp[13]) ? 4'b1001 : node2863;
													assign node2863 = (inp[10]) ? node2865 : 4'b0001;
														assign node2865 = (inp[12]) ? 4'b0001 : 4'b1001;
										assign node2869 = (inp[4]) ? node2883 : node2870;
											assign node2870 = (inp[10]) ? node2878 : node2871;
												assign node2871 = (inp[7]) ? 4'b0000 : node2872;
													assign node2872 = (inp[13]) ? 4'b1000 : node2873;
														assign node2873 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node2878 = (inp[7]) ? 4'b0000 : node2879;
													assign node2879 = (inp[13]) ? 4'b0100 : 4'b1000;
											assign node2883 = (inp[13]) ? node2891 : node2884;
												assign node2884 = (inp[7]) ? 4'b1000 : node2885;
													assign node2885 = (inp[2]) ? node2887 : 4'b1100;
														assign node2887 = (inp[10]) ? 4'b1100 : 4'b0100;
												assign node2891 = (inp[12]) ? node2893 : 4'b0100;
													assign node2893 = (inp[10]) ? 4'b0100 : 4'b1100;
								assign node2896 = (inp[13]) ? node2954 : node2897;
									assign node2897 = (inp[3]) ? node2923 : node2898;
										assign node2898 = (inp[2]) ? node2916 : node2899;
											assign node2899 = (inp[10]) ? node2907 : node2900;
												assign node2900 = (inp[12]) ? node2904 : node2901;
													assign node2901 = (inp[7]) ? 4'b1101 : 4'b1001;
													assign node2904 = (inp[4]) ? 4'b0001 : 4'b0101;
												assign node2907 = (inp[14]) ? node2913 : node2908;
													assign node2908 = (inp[7]) ? 4'b1101 : node2909;
														assign node2909 = (inp[4]) ? 4'b1001 : 4'b1101;
													assign node2913 = (inp[11]) ? 4'b1101 : 4'b1100;
											assign node2916 = (inp[4]) ? node2918 : 4'b0111;
												assign node2918 = (inp[7]) ? 4'b0111 : node2919;
													assign node2919 = (inp[14]) ? 4'b1000 : 4'b1001;
										assign node2923 = (inp[4]) ? node2935 : node2924;
											assign node2924 = (inp[12]) ? node2930 : node2925;
												assign node2925 = (inp[14]) ? node2927 : 4'b1001;
													assign node2927 = (inp[11]) ? 4'b1001 : 4'b1000;
												assign node2930 = (inp[10]) ? node2932 : 4'b0001;
													assign node2932 = (inp[11]) ? 4'b1001 : 4'b1000;
											assign node2935 = (inp[7]) ? node2945 : node2936;
												assign node2936 = (inp[14]) ? node2942 : node2937;
													assign node2937 = (inp[12]) ? node2939 : 4'b1101;
														assign node2939 = (inp[10]) ? 4'b1101 : 4'b0101;
													assign node2942 = (inp[11]) ? 4'b1101 : 4'b1100;
												assign node2945 = (inp[14]) ? node2951 : node2946;
													assign node2946 = (inp[10]) ? 4'b1001 : node2947;
														assign node2947 = (inp[11]) ? 4'b0001 : 4'b1001;
													assign node2951 = (inp[11]) ? 4'b1001 : 4'b1000;
									assign node2954 = (inp[14]) ? node2978 : node2955;
										assign node2955 = (inp[3]) ? node2967 : node2956;
											assign node2956 = (inp[12]) ? node2962 : node2957;
												assign node2957 = (inp[7]) ? node2959 : 4'b0001;
													assign node2959 = (inp[4]) ? 4'b0001 : 4'b0111;
												assign node2962 = (inp[2]) ? node2964 : 4'b1101;
													assign node2964 = (inp[4]) ? 4'b0001 : 4'b0111;
											assign node2967 = (inp[4]) ? node2973 : node2968;
												assign node2968 = (inp[7]) ? 4'b0001 : node2969;
													assign node2969 = (inp[10]) ? 4'b0101 : 4'b1001;
												assign node2973 = (inp[10]) ? 4'b0101 : node2974;
													assign node2974 = (inp[2]) ? 4'b1001 : 4'b0101;
										assign node2978 = (inp[11]) ? node2998 : node2979;
											assign node2979 = (inp[10]) ? node2989 : node2980;
												assign node2980 = (inp[3]) ? node2984 : node2981;
													assign node2981 = (inp[7]) ? 4'b0100 : 4'b0000;
													assign node2984 = (inp[4]) ? node2986 : 4'b1000;
														assign node2986 = (inp[7]) ? 4'b1000 : 4'b1100;
												assign node2989 = (inp[3]) ? node2993 : node2990;
													assign node2990 = (inp[7]) ? 4'b0100 : 4'b0000;
													assign node2993 = (inp[7]) ? node2995 : 4'b0100;
														assign node2995 = (inp[4]) ? 4'b0100 : 4'b0000;
											assign node2998 = (inp[12]) ? node3014 : node2999;
												assign node2999 = (inp[10]) ? node3011 : node3000;
													assign node3000 = (inp[2]) ? 4'b0001 : node3001;
														assign node3001 = (inp[7]) ? node3003 : 4'b0101;
															assign node3003 = (inp[4]) ? node3007 : node3004;
																assign node3004 = (inp[3]) ? 4'b0001 : 4'b0101;
																assign node3007 = (inp[3]) ? 4'b0101 : 4'b0001;
													assign node3011 = (inp[4]) ? 4'b0101 : 4'b0111;
												assign node3014 = (inp[4]) ? node3018 : node3015;
													assign node3015 = (inp[10]) ? 4'b0001 : 4'b1001;
													assign node3018 = (inp[10]) ? 4'b0001 : 4'b0111;
					assign node3022 = (inp[5]) ? node3438 : node3023;
						assign node3023 = (inp[0]) ? node3323 : node3024;
							assign node3024 = (inp[11]) ? node3194 : node3025;
								assign node3025 = (inp[10]) ? node3107 : node3026;
									assign node3026 = (inp[4]) ? node3070 : node3027;
										assign node3027 = (inp[7]) ? node3049 : node3028;
											assign node3028 = (inp[13]) ? node3038 : node3029;
												assign node3029 = (inp[12]) ? node3035 : node3030;
													assign node3030 = (inp[2]) ? node3032 : 4'b1100;
														assign node3032 = (inp[3]) ? 4'b1000 : 4'b1100;
													assign node3035 = (inp[2]) ? 4'b0100 : 4'b1100;
												assign node3038 = (inp[14]) ? 4'b1000 : node3039;
													assign node3039 = (inp[1]) ? 4'b1000 : node3040;
														assign node3040 = (inp[2]) ? node3042 : 4'b0000;
															assign node3042 = (inp[3]) ? 4'b0000 : node3043;
																assign node3043 = (inp[12]) ? 4'b1100 : 4'b0000;
											assign node3049 = (inp[2]) ? node3061 : node3050;
												assign node3050 = (inp[14]) ? node3054 : node3051;
													assign node3051 = (inp[3]) ? 4'b1100 : 4'b1101;
													assign node3054 = (inp[12]) ? node3056 : 4'b1100;
														assign node3056 = (inp[13]) ? node3058 : 4'b0100;
															assign node3058 = (inp[3]) ? 4'b0100 : 4'b1100;
												assign node3061 = (inp[3]) ? node3067 : node3062;
													assign node3062 = (inp[1]) ? node3064 : 4'b0101;
														assign node3064 = (inp[13]) ? 4'b0100 : 4'b1100;
													assign node3067 = (inp[12]) ? 4'b0001 : 4'b0000;
										assign node3070 = (inp[3]) ? node3088 : node3071;
											assign node3071 = (inp[2]) ? node3075 : node3072;
												assign node3072 = (inp[13]) ? 4'b1100 : 4'b1000;
												assign node3075 = (inp[7]) ? node3081 : node3076;
													assign node3076 = (inp[14]) ? 4'b1000 : node3077;
														assign node3077 = (inp[13]) ? 4'b1001 : 4'b0001;
													assign node3081 = (inp[12]) ? 4'b0101 : node3082;
														assign node3082 = (inp[14]) ? node3084 : 4'b1101;
															assign node3084 = (inp[1]) ? 4'b1100 : 4'b1101;
											assign node3088 = (inp[7]) ? node3098 : node3089;
												assign node3089 = (inp[1]) ? node3095 : node3090;
													assign node3090 = (inp[12]) ? node3092 : 4'b0100;
														assign node3092 = (inp[13]) ? 4'b1000 : 4'b0000;
													assign node3095 = (inp[13]) ? 4'b1100 : 4'b1001;
												assign node3098 = (inp[14]) ? 4'b1000 : node3099;
													assign node3099 = (inp[12]) ? 4'b0000 : node3100;
														assign node3100 = (inp[1]) ? node3102 : 4'b1000;
															assign node3102 = (inp[13]) ? 4'b1000 : 4'b0000;
									assign node3107 = (inp[1]) ? node3159 : node3108;
										assign node3108 = (inp[3]) ? node3138 : node3109;
											assign node3109 = (inp[14]) ? node3119 : node3110;
												assign node3110 = (inp[13]) ? node3116 : node3111;
													assign node3111 = (inp[4]) ? node3113 : 4'b1100;
														assign node3113 = (inp[7]) ? 4'b1100 : 4'b1000;
													assign node3116 = (inp[2]) ? 4'b0100 : 4'b0000;
												assign node3119 = (inp[4]) ? node3127 : node3120;
													assign node3120 = (inp[12]) ? node3124 : node3121;
														assign node3121 = (inp[13]) ? 4'b0001 : 4'b1101;
														assign node3124 = (inp[13]) ? 4'b1101 : 4'b0101;
													assign node3127 = (inp[2]) ? node3135 : node3128;
														assign node3128 = (inp[12]) ? node3132 : node3129;
															assign node3129 = (inp[7]) ? 4'b0000 : 4'b0100;
															assign node3132 = (inp[13]) ? 4'b1100 : 4'b1000;
														assign node3135 = (inp[13]) ? 4'b0001 : 4'b0101;
											assign node3138 = (inp[12]) ? node3150 : node3139;
												assign node3139 = (inp[2]) ? node3145 : node3140;
													assign node3140 = (inp[7]) ? node3142 : 4'b0000;
														assign node3142 = (inp[13]) ? 4'b0000 : 4'b0100;
													assign node3145 = (inp[7]) ? node3147 : 4'b0000;
														assign node3147 = (inp[13]) ? 4'b0000 : 4'b1001;
												assign node3150 = (inp[2]) ? node3154 : node3151;
													assign node3151 = (inp[7]) ? 4'b1100 : 4'b1000;
													assign node3154 = (inp[13]) ? 4'b1000 : node3155;
														assign node3155 = (inp[4]) ? 4'b1000 : 4'b0001;
										assign node3159 = (inp[4]) ? node3177 : node3160;
											assign node3160 = (inp[7]) ? node3168 : node3161;
												assign node3161 = (inp[2]) ? node3163 : 4'b0000;
													assign node3163 = (inp[14]) ? 4'b0000 : node3164;
														assign node3164 = (inp[3]) ? 4'b0000 : 4'b0001;
												assign node3168 = (inp[14]) ? node3170 : 4'b0000;
													assign node3170 = (inp[13]) ? node3172 : 4'b0100;
														assign node3172 = (inp[3]) ? 4'b0000 : node3173;
															assign node3173 = (inp[2]) ? 4'b0100 : 4'b0000;
											assign node3177 = (inp[13]) ? node3189 : node3178;
												assign node3178 = (inp[2]) ? node3182 : node3179;
													assign node3179 = (inp[3]) ? 4'b0001 : 4'b0000;
													assign node3182 = (inp[14]) ? node3186 : node3183;
														assign node3183 = (inp[12]) ? 4'b1101 : 4'b1001;
														assign node3186 = (inp[7]) ? 4'b1100 : 4'b1000;
												assign node3189 = (inp[3]) ? 4'b0100 : node3190;
													assign node3190 = (inp[7]) ? 4'b0001 : 4'b0000;
								assign node3194 = (inp[1]) ? node3264 : node3195;
									assign node3195 = (inp[3]) ? node3227 : node3196;
										assign node3196 = (inp[13]) ? node3216 : node3197;
											assign node3197 = (inp[4]) ? node3203 : node3198;
												assign node3198 = (inp[12]) ? node3200 : 4'b1100;
													assign node3200 = (inp[10]) ? 4'b1100 : 4'b0100;
												assign node3203 = (inp[2]) ? node3213 : node3204;
													assign node3204 = (inp[14]) ? 4'b0101 : node3205;
														assign node3205 = (inp[12]) ? node3209 : node3206;
															assign node3206 = (inp[7]) ? 4'b0001 : 4'b1001;
															assign node3209 = (inp[7]) ? 4'b1001 : 4'b0001;
													assign node3213 = (inp[12]) ? 4'b0100 : 4'b1100;
											assign node3216 = (inp[12]) ? node3220 : node3217;
												assign node3217 = (inp[2]) ? 4'b0000 : 4'b0001;
												assign node3220 = (inp[14]) ? node3224 : node3221;
													assign node3221 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node3224 = (inp[10]) ? 4'b0100 : 4'b1100;
										assign node3227 = (inp[2]) ? node3245 : node3228;
											assign node3228 = (inp[4]) ? node3236 : node3229;
												assign node3229 = (inp[13]) ? node3231 : 4'b0101;
													assign node3231 = (inp[12]) ? node3233 : 4'b0000;
														assign node3233 = (inp[10]) ? 4'b1001 : 4'b0001;
												assign node3236 = (inp[13]) ? 4'b0100 : node3237;
													assign node3237 = (inp[12]) ? node3239 : 4'b1000;
														assign node3239 = (inp[10]) ? 4'b0000 : node3240;
															assign node3240 = (inp[7]) ? 4'b0001 : 4'b1000;
											assign node3245 = (inp[4]) ? node3257 : node3246;
												assign node3246 = (inp[12]) ? node3252 : node3247;
													assign node3247 = (inp[7]) ? 4'b0000 : node3248;
														assign node3248 = (inp[10]) ? 4'b0001 : 4'b1001;
													assign node3252 = (inp[10]) ? node3254 : 4'b1000;
														assign node3254 = (inp[13]) ? 4'b1001 : 4'b1000;
												assign node3257 = (inp[13]) ? node3259 : 4'b0001;
													assign node3259 = (inp[12]) ? node3261 : 4'b1001;
														assign node3261 = (inp[10]) ? 4'b1101 : 4'b0101;
									assign node3264 = (inp[10]) ? node3298 : node3265;
										assign node3265 = (inp[4]) ? node3283 : node3266;
											assign node3266 = (inp[2]) ? node3276 : node3267;
												assign node3267 = (inp[13]) ? node3273 : node3268;
													assign node3268 = (inp[12]) ? node3270 : 4'b1101;
														assign node3270 = (inp[7]) ? 4'b0101 : 4'b1101;
													assign node3273 = (inp[7]) ? 4'b0101 : 4'b1001;
												assign node3276 = (inp[3]) ? node3278 : 4'b1101;
													assign node3278 = (inp[13]) ? 4'b1001 : node3279;
														assign node3279 = (inp[12]) ? 4'b0001 : 4'b1001;
											assign node3283 = (inp[2]) ? node3289 : node3284;
												assign node3284 = (inp[3]) ? 4'b0001 : node3285;
													assign node3285 = (inp[13]) ? 4'b1101 : 4'b1001;
												assign node3289 = (inp[3]) ? 4'b1001 : node3290;
													assign node3290 = (inp[13]) ? 4'b0001 : node3291;
														assign node3291 = (inp[7]) ? 4'b1101 : node3292;
															assign node3292 = (inp[12]) ? 4'b0001 : 4'b1001;
										assign node3298 = (inp[13]) ? node3312 : node3299;
											assign node3299 = (inp[7]) ? node3305 : node3300;
												assign node3300 = (inp[4]) ? node3302 : 4'b0001;
													assign node3302 = (inp[14]) ? 4'b1001 : 4'b0101;
												assign node3305 = (inp[2]) ? node3309 : node3306;
													assign node3306 = (inp[3]) ? 4'b0101 : 4'b1101;
													assign node3309 = (inp[3]) ? 4'b1001 : 4'b1101;
											assign node3312 = (inp[4]) ? node3318 : node3313;
												assign node3313 = (inp[3]) ? 4'b0001 : node3314;
													assign node3314 = (inp[7]) ? 4'b0101 : 4'b0001;
												assign node3318 = (inp[3]) ? 4'b0101 : node3319;
													assign node3319 = (inp[2]) ? 4'b0001 : 4'b0101;
							assign node3323 = (inp[2]) ? 4'b0101 : node3324;
								assign node3324 = (inp[3]) ? node3358 : node3325;
									assign node3325 = (inp[4]) ? node3337 : node3326;
										assign node3326 = (inp[13]) ? node3328 : 4'b0101;
											assign node3328 = (inp[1]) ? 4'b0101 : node3329;
												assign node3329 = (inp[7]) ? 4'b0101 : node3330;
													assign node3330 = (inp[11]) ? 4'b0000 : node3331;
														assign node3331 = (inp[12]) ? 4'b0101 : 4'b0001;
										assign node3337 = (inp[7]) ? node3353 : node3338;
											assign node3338 = (inp[13]) ? node3342 : node3339;
												assign node3339 = (inp[10]) ? 4'b1000 : 4'b0000;
												assign node3342 = (inp[12]) ? node3348 : node3343;
													assign node3343 = (inp[1]) ? 4'b0001 : node3344;
														assign node3344 = (inp[10]) ? 4'b0001 : 4'b1001;
													assign node3348 = (inp[10]) ? 4'b0000 : node3349;
														assign node3349 = (inp[11]) ? 4'b1001 : 4'b1000;
											assign node3353 = (inp[13]) ? node3355 : 4'b0101;
												assign node3355 = (inp[1]) ? 4'b0001 : 4'b0000;
									assign node3358 = (inp[13]) ? node3396 : node3359;
										assign node3359 = (inp[7]) ? node3377 : node3360;
											assign node3360 = (inp[4]) ? node3366 : node3361;
												assign node3361 = (inp[14]) ? node3363 : 4'b1000;
													assign node3363 = (inp[11]) ? 4'b1000 : 4'b0001;
												assign node3366 = (inp[12]) ? node3372 : node3367;
													assign node3367 = (inp[11]) ? 4'b1100 : node3368;
														assign node3368 = (inp[1]) ? 4'b1100 : 4'b1101;
													assign node3372 = (inp[11]) ? node3374 : 4'b0101;
														assign node3374 = (inp[1]) ? 4'b1101 : 4'b1100;
											assign node3377 = (inp[1]) ? node3389 : node3378;
												assign node3378 = (inp[11]) ? node3384 : node3379;
													assign node3379 = (inp[14]) ? node3381 : 4'b1000;
														assign node3381 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node3384 = (inp[10]) ? 4'b1000 : node3385;
														assign node3385 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node3389 = (inp[10]) ? 4'b1001 : node3390;
													assign node3390 = (inp[12]) ? node3392 : 4'b1001;
														assign node3392 = (inp[11]) ? 4'b0001 : 4'b0000;
										assign node3396 = (inp[10]) ? node3422 : node3397;
											assign node3397 = (inp[12]) ? node3407 : node3398;
												assign node3398 = (inp[14]) ? node3402 : node3399;
													assign node3399 = (inp[1]) ? 4'b0101 : 4'b0100;
													assign node3402 = (inp[4]) ? 4'b1001 : node3403;
														assign node3403 = (inp[7]) ? 4'b0001 : 4'b0101;
												assign node3407 = (inp[7]) ? node3417 : node3408;
													assign node3408 = (inp[4]) ? node3414 : node3409;
														assign node3409 = (inp[11]) ? 4'b1001 : node3410;
															assign node3410 = (inp[1]) ? 4'b1000 : 4'b1001;
														assign node3414 = (inp[1]) ? 4'b1101 : 4'b1100;
													assign node3417 = (inp[11]) ? 4'b1001 : node3418;
														assign node3418 = (inp[1]) ? 4'b1000 : 4'b1001;
											assign node3422 = (inp[1]) ? node3428 : node3423;
												assign node3423 = (inp[11]) ? 4'b0100 : node3424;
													assign node3424 = (inp[4]) ? 4'b0100 : 4'b0000;
												assign node3428 = (inp[11]) ? node3432 : node3429;
													assign node3429 = (inp[14]) ? 4'b0100 : 4'b0101;
													assign node3432 = (inp[7]) ? node3434 : 4'b0101;
														assign node3434 = (inp[4]) ? 4'b0101 : 4'b0001;
						assign node3438 = (inp[3]) ? node3762 : node3439;
							assign node3439 = (inp[4]) ? node3593 : node3440;
								assign node3440 = (inp[0]) ? node3542 : node3441;
									assign node3441 = (inp[13]) ? node3495 : node3442;
										assign node3442 = (inp[10]) ? node3472 : node3443;
											assign node3443 = (inp[14]) ? node3455 : node3444;
												assign node3444 = (inp[2]) ? node3450 : node3445;
													assign node3445 = (inp[11]) ? node3447 : 4'b1101;
														assign node3447 = (inp[1]) ? 4'b1101 : 4'b1100;
													assign node3450 = (inp[7]) ? node3452 : 4'b1101;
														assign node3452 = (inp[1]) ? 4'b1101 : 4'b0101;
												assign node3455 = (inp[7]) ? node3465 : node3456;
													assign node3456 = (inp[1]) ? node3462 : node3457;
														assign node3457 = (inp[2]) ? node3459 : 4'b1100;
															assign node3459 = (inp[12]) ? 4'b0101 : 4'b1101;
														assign node3462 = (inp[2]) ? 4'b1100 : 4'b0001;
													assign node3465 = (inp[1]) ? node3467 : 4'b1100;
														assign node3467 = (inp[2]) ? 4'b1100 : node3468;
															assign node3468 = (inp[12]) ? 4'b1101 : 4'b0101;
											assign node3472 = (inp[7]) ? node3484 : node3473;
												assign node3473 = (inp[2]) ? node3479 : node3474;
													assign node3474 = (inp[11]) ? node3476 : 4'b0001;
														assign node3476 = (inp[1]) ? 4'b0001 : 4'b1001;
													assign node3479 = (inp[1]) ? 4'b1001 : node3480;
														assign node3480 = (inp[12]) ? 4'b0001 : 4'b1000;
												assign node3484 = (inp[1]) ? node3492 : node3485;
													assign node3485 = (inp[14]) ? 4'b0100 : node3486;
														assign node3486 = (inp[11]) ? 4'b0101 : node3487;
															assign node3487 = (inp[2]) ? 4'b1100 : 4'b0101;
													assign node3492 = (inp[2]) ? 4'b0100 : 4'b0001;
										assign node3495 = (inp[1]) ? node3515 : node3496;
											assign node3496 = (inp[2]) ? node3510 : node3497;
												assign node3497 = (inp[11]) ? node3505 : node3498;
													assign node3498 = (inp[12]) ? node3500 : 4'b1001;
														assign node3500 = (inp[10]) ? node3502 : 4'b0001;
															assign node3502 = (inp[7]) ? 4'b0001 : 4'b0101;
													assign node3505 = (inp[7]) ? 4'b1001 : node3506;
														assign node3506 = (inp[10]) ? 4'b1101 : 4'b1001;
												assign node3510 = (inp[10]) ? node3512 : 4'b0000;
													assign node3512 = (inp[14]) ? 4'b1000 : 4'b1001;
											assign node3515 = (inp[14]) ? node3533 : node3516;
												assign node3516 = (inp[12]) ? node3530 : node3517;
													assign node3517 = (inp[2]) ? node3523 : node3518;
														assign node3518 = (inp[7]) ? node3520 : 4'b0101;
															assign node3520 = (inp[10]) ? 4'b0101 : 4'b0001;
														assign node3523 = (inp[11]) ? node3527 : node3524;
															assign node3524 = (inp[7]) ? 4'b0000 : 4'b1000;
															assign node3527 = (inp[7]) ? 4'b0001 : 4'b0101;
													assign node3530 = (inp[11]) ? 4'b0101 : 4'b1101;
												assign node3533 = (inp[2]) ? node3537 : node3534;
													assign node3534 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node3537 = (inp[11]) ? 4'b1001 : node3538;
														assign node3538 = (inp[10]) ? 4'b1001 : 4'b0001;
									assign node3542 = (inp[2]) ? node3576 : node3543;
										assign node3543 = (inp[13]) ? node3565 : node3544;
											assign node3544 = (inp[7]) ? node3562 : node3545;
												assign node3545 = (inp[12]) ? node3555 : node3546;
													assign node3546 = (inp[10]) ? 4'b0001 : node3547;
														assign node3547 = (inp[11]) ? 4'b1101 : node3548;
															assign node3548 = (inp[14]) ? 4'b1100 : node3549;
																assign node3549 = (inp[1]) ? 4'b1101 : 4'b1100;
													assign node3555 = (inp[10]) ? 4'b1100 : node3556;
														assign node3556 = (inp[11]) ? node3558 : 4'b0101;
															assign node3558 = (inp[1]) ? 4'b0101 : 4'b0100;
												assign node3562 = (inp[10]) ? 4'b1100 : 4'b0100;
											assign node3565 = (inp[10]) ? node3569 : node3566;
												assign node3566 = (inp[7]) ? 4'b0100 : 4'b1000;
												assign node3569 = (inp[11]) ? node3571 : 4'b0000;
													assign node3571 = (inp[12]) ? node3573 : 4'b0001;
														assign node3573 = (inp[1]) ? 4'b0001 : 4'b1001;
										assign node3576 = (inp[7]) ? 4'b0101 : node3577;
											assign node3577 = (inp[13]) ? node3579 : 4'b0101;
												assign node3579 = (inp[10]) ? node3585 : node3580;
													assign node3580 = (inp[12]) ? 4'b0101 : node3581;
														assign node3581 = (inp[1]) ? 4'b0001 : 4'b0101;
													assign node3585 = (inp[14]) ? node3587 : 4'b0000;
														assign node3587 = (inp[1]) ? 4'b0000 : node3588;
															assign node3588 = (inp[12]) ? 4'b0101 : 4'b0001;
								assign node3593 = (inp[1]) ? node3695 : node3594;
									assign node3594 = (inp[7]) ? node3634 : node3595;
										assign node3595 = (inp[11]) ? node3609 : node3596;
											assign node3596 = (inp[13]) ? node3604 : node3597;
												assign node3597 = (inp[0]) ? node3599 : 4'b1001;
													assign node3599 = (inp[12]) ? node3601 : 4'b1000;
														assign node3601 = (inp[14]) ? 4'b0000 : 4'b1000;
												assign node3604 = (inp[0]) ? 4'b1001 : node3605;
													assign node3605 = (inp[10]) ? 4'b0001 : 4'b1001;
											assign node3609 = (inp[13]) ? node3619 : node3610;
												assign node3610 = (inp[2]) ? node3616 : node3611;
													assign node3611 = (inp[10]) ? 4'b0100 : node3612;
														assign node3612 = (inp[14]) ? 4'b1000 : 4'b0000;
													assign node3616 = (inp[10]) ? 4'b1001 : 4'b1100;
												assign node3619 = (inp[14]) ? node3629 : node3620;
													assign node3620 = (inp[10]) ? node3624 : node3621;
														assign node3621 = (inp[0]) ? 4'b0000 : 4'b0001;
														assign node3624 = (inp[12]) ? node3626 : 4'b1000;
															assign node3626 = (inp[2]) ? 4'b0000 : 4'b1000;
													assign node3629 = (inp[2]) ? 4'b1000 : node3630;
														assign node3630 = (inp[12]) ? 4'b1001 : 4'b1000;
										assign node3634 = (inp[14]) ? node3668 : node3635;
											assign node3635 = (inp[10]) ? node3649 : node3636;
												assign node3636 = (inp[2]) ? node3644 : node3637;
													assign node3637 = (inp[12]) ? node3639 : 4'b0001;
														assign node3639 = (inp[0]) ? node3641 : 4'b0100;
															assign node3641 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node3644 = (inp[0]) ? 4'b0101 : node3645;
														assign node3645 = (inp[11]) ? 4'b1001 : 4'b0001;
												assign node3649 = (inp[2]) ? node3663 : node3650;
													assign node3650 = (inp[11]) ? node3658 : node3651;
														assign node3651 = (inp[12]) ? node3655 : node3652;
															assign node3652 = (inp[13]) ? 4'b0100 : 4'b0000;
															assign node3655 = (inp[0]) ? 4'b1000 : 4'b0000;
														assign node3658 = (inp[13]) ? node3660 : 4'b0001;
															assign node3660 = (inp[0]) ? 4'b0000 : 4'b0001;
													assign node3663 = (inp[13]) ? 4'b0000 : node3664;
														assign node3664 = (inp[0]) ? 4'b0101 : 4'b1100;
											assign node3668 = (inp[11]) ? node3686 : node3669;
												assign node3669 = (inp[12]) ? node3681 : node3670;
													assign node3670 = (inp[13]) ? node3678 : node3671;
														assign node3671 = (inp[2]) ? node3673 : 4'b1000;
															assign node3673 = (inp[0]) ? 4'b0101 : node3674;
																assign node3674 = (inp[10]) ? 4'b0100 : 4'b1000;
														assign node3678 = (inp[2]) ? 4'b1001 : 4'b0101;
													assign node3681 = (inp[13]) ? node3683 : 4'b0101;
														assign node3683 = (inp[2]) ? 4'b0101 : 4'b0000;
												assign node3686 = (inp[10]) ? 4'b1001 : node3687;
													assign node3687 = (inp[0]) ? node3689 : 4'b0100;
														assign node3689 = (inp[2]) ? 4'b0000 : node3690;
															assign node3690 = (inp[12]) ? 4'b0001 : 4'b1001;
									assign node3695 = (inp[11]) ? node3741 : node3696;
										assign node3696 = (inp[2]) ? node3720 : node3697;
											assign node3697 = (inp[13]) ? node3709 : node3698;
												assign node3698 = (inp[10]) ? node3704 : node3699;
													assign node3699 = (inp[0]) ? 4'b1000 : node3700;
														assign node3700 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node3704 = (inp[12]) ? node3706 : 4'b0000;
														assign node3706 = (inp[14]) ? 4'b0100 : 4'b0101;
												assign node3709 = (inp[0]) ? node3713 : node3710;
													assign node3710 = (inp[10]) ? 4'b1001 : 4'b1000;
													assign node3713 = (inp[14]) ? 4'b0001 : node3714;
														assign node3714 = (inp[7]) ? node3716 : 4'b0000;
															assign node3716 = (inp[12]) ? 4'b0000 : 4'b1000;
											assign node3720 = (inp[10]) ? node3734 : node3721;
												assign node3721 = (inp[12]) ? node3729 : node3722;
													assign node3722 = (inp[14]) ? node3724 : 4'b0001;
														assign node3724 = (inp[7]) ? 4'b0101 : node3725;
															assign node3725 = (inp[13]) ? 4'b0101 : 4'b0001;
													assign node3729 = (inp[0]) ? 4'b0101 : node3730;
														assign node3730 = (inp[7]) ? 4'b1001 : 4'b1101;
												assign node3734 = (inp[0]) ? node3738 : node3735;
													assign node3735 = (inp[12]) ? 4'b1001 : 4'b0001;
													assign node3738 = (inp[14]) ? 4'b1000 : 4'b1001;
										assign node3741 = (inp[12]) ? node3759 : node3742;
											assign node3742 = (inp[2]) ? node3748 : node3743;
												assign node3743 = (inp[10]) ? node3745 : 4'b1001;
													assign node3745 = (inp[14]) ? 4'b0101 : 4'b0001;
												assign node3748 = (inp[7]) ? node3754 : node3749;
													assign node3749 = (inp[13]) ? 4'b0001 : node3750;
														assign node3750 = (inp[0]) ? 4'b1001 : 4'b0001;
													assign node3754 = (inp[13]) ? 4'b0001 : node3755;
														assign node3755 = (inp[10]) ? 4'b0001 : 4'b0101;
											assign node3759 = (inp[0]) ? 4'b0101 : 4'b0001;
							assign node3762 = (inp[13]) ? node3922 : node3763;
								assign node3763 = (inp[11]) ? node3859 : node3764;
									assign node3764 = (inp[10]) ? node3810 : node3765;
										assign node3765 = (inp[2]) ? node3793 : node3766;
											assign node3766 = (inp[14]) ? node3780 : node3767;
												assign node3767 = (inp[12]) ? node3773 : node3768;
													assign node3768 = (inp[0]) ? 4'b0001 : node3769;
														assign node3769 = (inp[1]) ? 4'b1001 : 4'b0001;
													assign node3773 = (inp[0]) ? node3777 : node3774;
														assign node3774 = (inp[4]) ? 4'b0001 : 4'b1001;
														assign node3777 = (inp[7]) ? 4'b1000 : 4'b1001;
												assign node3780 = (inp[7]) ? node3786 : node3781;
													assign node3781 = (inp[1]) ? node3783 : 4'b0000;
														assign node3783 = (inp[0]) ? 4'b1001 : 4'b1000;
													assign node3786 = (inp[1]) ? 4'b0000 : node3787;
														assign node3787 = (inp[4]) ? 4'b1000 : node3788;
															assign node3788 = (inp[0]) ? 4'b0000 : 4'b1000;
											assign node3793 = (inp[4]) ? node3803 : node3794;
												assign node3794 = (inp[12]) ? node3800 : node3795;
													assign node3795 = (inp[14]) ? 4'b1001 : node3796;
														assign node3796 = (inp[1]) ? 4'b1001 : 4'b1000;
													assign node3800 = (inp[14]) ? 4'b0001 : 4'b0000;
												assign node3803 = (inp[12]) ? node3805 : 4'b1000;
													assign node3805 = (inp[0]) ? node3807 : 4'b1000;
														assign node3807 = (inp[1]) ? 4'b1000 : 4'b0000;
										assign node3810 = (inp[4]) ? node3836 : node3811;
											assign node3811 = (inp[2]) ? node3819 : node3812;
												assign node3812 = (inp[14]) ? 4'b1001 : node3813;
													assign node3813 = (inp[12]) ? node3815 : 4'b0001;
														assign node3815 = (inp[7]) ? 4'b0001 : 4'b0000;
												assign node3819 = (inp[14]) ? node3831 : node3820;
													assign node3820 = (inp[0]) ? node3826 : node3821;
														assign node3821 = (inp[12]) ? 4'b0000 : node3822;
															assign node3822 = (inp[7]) ? 4'b0000 : 4'b1000;
														assign node3826 = (inp[1]) ? 4'b1001 : node3827;
															assign node3827 = (inp[12]) ? 4'b1000 : 4'b0000;
													assign node3831 = (inp[12]) ? node3833 : 4'b0000;
														assign node3833 = (inp[1]) ? 4'b1000 : 4'b0000;
											assign node3836 = (inp[2]) ? node3848 : node3837;
												assign node3837 = (inp[12]) ? node3843 : node3838;
													assign node3838 = (inp[7]) ? 4'b1001 : node3839;
														assign node3839 = (inp[14]) ? 4'b0000 : 4'b1000;
													assign node3843 = (inp[7]) ? 4'b0000 : node3844;
														assign node3844 = (inp[1]) ? 4'b0001 : 4'b0000;
												assign node3848 = (inp[1]) ? node3850 : 4'b0001;
													assign node3850 = (inp[14]) ? node3854 : node3851;
														assign node3851 = (inp[7]) ? 4'b0000 : 4'b1000;
														assign node3854 = (inp[12]) ? node3856 : 4'b0001;
															assign node3856 = (inp[0]) ? 4'b0000 : 4'b0001;
									assign node3859 = (inp[1]) ? node3895 : node3860;
										assign node3860 = (inp[10]) ? node3880 : node3861;
											assign node3861 = (inp[4]) ? node3869 : node3862;
												assign node3862 = (inp[12]) ? node3864 : 4'b0000;
													assign node3864 = (inp[0]) ? node3866 : 4'b1000;
														assign node3866 = (inp[2]) ? 4'b0000 : 4'b1000;
												assign node3869 = (inp[2]) ? node3875 : node3870;
													assign node3870 = (inp[7]) ? node3872 : 4'b0001;
														assign node3872 = (inp[0]) ? 4'b0000 : 4'b0001;
													assign node3875 = (inp[14]) ? node3877 : 4'b0001;
														assign node3877 = (inp[12]) ? 4'b1000 : 4'b1001;
											assign node3880 = (inp[0]) ? node3892 : node3881;
												assign node3881 = (inp[4]) ? node3887 : node3882;
													assign node3882 = (inp[7]) ? node3884 : 4'b0001;
														assign node3884 = (inp[2]) ? 4'b1001 : 4'b0001;
													assign node3887 = (inp[14]) ? node3889 : 4'b0001;
														assign node3889 = (inp[7]) ? 4'b0000 : 4'b0001;
												assign node3892 = (inp[7]) ? 4'b1000 : 4'b0001;
										assign node3895 = (inp[12]) ? node3907 : node3896;
											assign node3896 = (inp[10]) ? node3902 : node3897;
												assign node3897 = (inp[7]) ? node3899 : 4'b1001;
													assign node3899 = (inp[2]) ? 4'b1001 : 4'b0001;
												assign node3902 = (inp[14]) ? 4'b0001 : node3903;
													assign node3903 = (inp[7]) ? 4'b1001 : 4'b0001;
											assign node3907 = (inp[10]) ? node3913 : node3908;
												assign node3908 = (inp[14]) ? node3910 : 4'b0001;
													assign node3910 = (inp[4]) ? 4'b1001 : 4'b0001;
												assign node3913 = (inp[7]) ? node3915 : 4'b0001;
													assign node3915 = (inp[4]) ? 4'b0001 : node3916;
														assign node3916 = (inp[0]) ? node3918 : 4'b1001;
															assign node3918 = (inp[2]) ? 4'b1001 : 4'b0001;
								assign node3922 = (inp[4]) ? node4000 : node3923;
									assign node3923 = (inp[1]) ? node3979 : node3924;
										assign node3924 = (inp[11]) ? node3950 : node3925;
											assign node3925 = (inp[10]) ? node3943 : node3926;
												assign node3926 = (inp[12]) ? node3932 : node3927;
													assign node3927 = (inp[7]) ? 4'b0000 : node3928;
														assign node3928 = (inp[14]) ? 4'b0001 : 4'b0000;
													assign node3932 = (inp[7]) ? node3938 : node3933;
														assign node3933 = (inp[2]) ? 4'b0001 : node3934;
															assign node3934 = (inp[0]) ? 4'b0001 : 4'b1000;
														assign node3938 = (inp[0]) ? node3940 : 4'b0001;
															assign node3940 = (inp[2]) ? 4'b1000 : 4'b0001;
												assign node3943 = (inp[0]) ? 4'b0000 : node3944;
													assign node3944 = (inp[12]) ? 4'b0000 : node3945;
														assign node3945 = (inp[7]) ? 4'b1001 : 4'b1000;
											assign node3950 = (inp[12]) ? node3962 : node3951;
												assign node3951 = (inp[2]) ? node3957 : node3952;
													assign node3952 = (inp[7]) ? 4'b1001 : node3953;
														assign node3953 = (inp[10]) ? 4'b1001 : 4'b0000;
													assign node3957 = (inp[7]) ? node3959 : 4'b1001;
														assign node3959 = (inp[10]) ? 4'b0001 : 4'b0000;
												assign node3962 = (inp[10]) ? node3970 : node3963;
													assign node3963 = (inp[7]) ? node3967 : node3964;
														assign node3964 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node3967 = (inp[2]) ? 4'b1000 : 4'b0001;
													assign node3970 = (inp[7]) ? node3974 : node3971;
														assign node3971 = (inp[14]) ? 4'b1001 : 4'b0001;
														assign node3974 = (inp[2]) ? 4'b0000 : node3975;
															assign node3975 = (inp[0]) ? 4'b1000 : 4'b1001;
										assign node3979 = (inp[11]) ? 4'b0001 : node3980;
											assign node3980 = (inp[10]) ? node3990 : node3981;
												assign node3981 = (inp[12]) ? 4'b1001 : node3982;
													assign node3982 = (inp[14]) ? node3984 : 4'b0001;
														assign node3984 = (inp[2]) ? 4'b0000 : node3985;
															assign node3985 = (inp[0]) ? 4'b0001 : 4'b0000;
												assign node3990 = (inp[0]) ? node3994 : node3991;
													assign node3991 = (inp[12]) ? 4'b0000 : 4'b1001;
													assign node3994 = (inp[7]) ? 4'b0000 : node3995;
														assign node3995 = (inp[2]) ? 4'b0001 : 4'b0000;
									assign node4000 = (inp[10]) ? node4038 : node4001;
										assign node4001 = (inp[1]) ? node4027 : node4002;
											assign node4002 = (inp[0]) ? node4014 : node4003;
												assign node4003 = (inp[11]) ? 4'b0000 : node4004;
													assign node4004 = (inp[14]) ? node4006 : 4'b0000;
														assign node4006 = (inp[12]) ? node4008 : 4'b0000;
															assign node4008 = (inp[2]) ? node4010 : 4'b0001;
																assign node4010 = (inp[7]) ? 4'b0000 : 4'b0001;
												assign node4014 = (inp[7]) ? node4022 : node4015;
													assign node4015 = (inp[11]) ? 4'b0000 : node4016;
														assign node4016 = (inp[14]) ? 4'b0001 : node4017;
															assign node4017 = (inp[2]) ? 4'b0001 : 4'b0000;
													assign node4022 = (inp[12]) ? node4024 : 4'b0001;
														assign node4024 = (inp[11]) ? 4'b0001 : 4'b0000;
											assign node4027 = (inp[11]) ? 4'b0001 : node4028;
												assign node4028 = (inp[14]) ? node4030 : 4'b0000;
													assign node4030 = (inp[0]) ? node4032 : 4'b0000;
														assign node4032 = (inp[2]) ? node4034 : 4'b0001;
															assign node4034 = (inp[12]) ? 4'b0000 : 4'b0001;
										assign node4038 = (inp[12]) ? node4040 : 4'b0000;
											assign node4040 = (inp[7]) ? 4'b0000 : node4041;
												assign node4041 = (inp[0]) ? 4'b0000 : node4042;
													assign node4042 = (inp[1]) ? 4'b0000 : node4043;
														assign node4043 = (inp[2]) ? 4'b0000 : 4'b0001;
				assign node4049 = (inp[0]) ? node4879 : node4050;
					assign node4050 = (inp[6]) ? node4280 : node4051;
						assign node4051 = (inp[2]) ? node4243 : node4052;
							assign node4052 = (inp[5]) ? node4092 : node4053;
								assign node4053 = (inp[3]) ? node4055 : 4'b0011;
									assign node4055 = (inp[7]) ? node4081 : node4056;
										assign node4056 = (inp[4]) ? node4068 : node4057;
											assign node4057 = (inp[13]) ? node4059 : 4'b0011;
												assign node4059 = (inp[12]) ? node4063 : node4060;
													assign node4060 = (inp[1]) ? 4'b0001 : 4'b0000;
													assign node4063 = (inp[10]) ? node4065 : 4'b0011;
														assign node4065 = (inp[14]) ? 4'b0000 : 4'b0001;
											assign node4068 = (inp[1]) ? node4074 : node4069;
												assign node4069 = (inp[11]) ? 4'b1000 : node4070;
													assign node4070 = (inp[13]) ? 4'b0000 : 4'b0001;
												assign node4074 = (inp[11]) ? node4076 : 4'b0000;
													assign node4076 = (inp[13]) ? 4'b0001 : node4077;
														assign node4077 = (inp[10]) ? 4'b1001 : 4'b0001;
										assign node4081 = (inp[13]) ? node4083 : 4'b0011;
											assign node4083 = (inp[14]) ? 4'b0011 : node4084;
												assign node4084 = (inp[4]) ? node4086 : 4'b0011;
													assign node4086 = (inp[1]) ? node4088 : 4'b0000;
														assign node4088 = (inp[11]) ? 4'b0001 : 4'b0011;
								assign node4092 = (inp[1]) ? node4174 : node4093;
									assign node4093 = (inp[14]) ? node4133 : node4094;
										assign node4094 = (inp[13]) ? node4112 : node4095;
											assign node4095 = (inp[11]) ? node4105 : node4096;
												assign node4096 = (inp[3]) ? node4100 : node4097;
													assign node4097 = (inp[7]) ? 4'b1000 : 4'b1100;
													assign node4100 = (inp[10]) ? 4'b1100 : node4101;
														assign node4101 = (inp[4]) ? 4'b0100 : 4'b1100;
												assign node4105 = (inp[3]) ? node4109 : node4106;
													assign node4106 = (inp[7]) ? 4'b1000 : 4'b1100;
													assign node4109 = (inp[7]) ? 4'b1100 : 4'b1000;
											assign node4112 = (inp[10]) ? node4124 : node4113;
												assign node4113 = (inp[12]) ? node4117 : node4114;
													assign node4114 = (inp[11]) ? 4'b0000 : 4'b0100;
													assign node4117 = (inp[4]) ? node4121 : node4118;
														assign node4118 = (inp[3]) ? 4'b1100 : 4'b1000;
														assign node4121 = (inp[3]) ? 4'b1000 : 4'b1100;
												assign node4124 = (inp[4]) ? node4130 : node4125;
													assign node4125 = (inp[12]) ? 4'b0100 : node4126;
														assign node4126 = (inp[11]) ? 4'b0000 : 4'b0100;
													assign node4130 = (inp[3]) ? 4'b0000 : 4'b0100;
										assign node4133 = (inp[11]) ? node4163 : node4134;
											assign node4134 = (inp[13]) ? node4150 : node4135;
												assign node4135 = (inp[12]) ? node4139 : node4136;
													assign node4136 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node4139 = (inp[4]) ? node4143 : node4140;
														assign node4140 = (inp[3]) ? 4'b0101 : 4'b0001;
														assign node4143 = (inp[10]) ? 4'b0101 : node4144;
															assign node4144 = (inp[7]) ? 4'b0001 : node4145;
																assign node4145 = (inp[3]) ? 4'b0001 : 4'b0101;
												assign node4150 = (inp[10]) ? node4160 : node4151;
													assign node4151 = (inp[4]) ? node4153 : 4'b1001;
														assign node4153 = (inp[3]) ? node4157 : node4154;
															assign node4154 = (inp[7]) ? 4'b1001 : 4'b1101;
															assign node4157 = (inp[7]) ? 4'b1101 : 4'b1001;
													assign node4160 = (inp[7]) ? 4'b1101 : 4'b0101;
											assign node4163 = (inp[13]) ? node4167 : node4164;
												assign node4164 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node4167 = (inp[3]) ? node4169 : 4'b0100;
													assign node4169 = (inp[10]) ? 4'b0000 : node4170;
														assign node4170 = (inp[12]) ? 4'b1100 : 4'b0000;
									assign node4174 = (inp[13]) ? node4206 : node4175;
										assign node4175 = (inp[11]) ? node4195 : node4176;
											assign node4176 = (inp[14]) ? node4186 : node4177;
												assign node4177 = (inp[12]) ? node4183 : node4178;
													assign node4178 = (inp[3]) ? 4'b1101 : node4179;
														assign node4179 = (inp[7]) ? 4'b1001 : 4'b1101;
													assign node4183 = (inp[10]) ? 4'b1001 : 4'b0101;
												assign node4186 = (inp[3]) ? node4192 : node4187;
													assign node4187 = (inp[10]) ? 4'b1000 : node4188;
														assign node4188 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node4192 = (inp[12]) ? 4'b0100 : 4'b1100;
											assign node4195 = (inp[3]) ? node4201 : node4196;
												assign node4196 = (inp[7]) ? 4'b1001 : node4197;
													assign node4197 = (inp[4]) ? 4'b1101 : 4'b1001;
												assign node4201 = (inp[7]) ? 4'b1101 : node4202;
													assign node4202 = (inp[4]) ? 4'b1001 : 4'b1101;
										assign node4206 = (inp[10]) ? node4230 : node4207;
											assign node4207 = (inp[12]) ? node4219 : node4208;
												assign node4208 = (inp[3]) ? node4214 : node4209;
													assign node4209 = (inp[11]) ? node4211 : 4'b0100;
														assign node4211 = (inp[7]) ? 4'b0001 : 4'b0101;
													assign node4214 = (inp[14]) ? node4216 : 4'b0001;
														assign node4216 = (inp[7]) ? 4'b0001 : 4'b0000;
												assign node4219 = (inp[3]) ? node4225 : node4220;
													assign node4220 = (inp[11]) ? node4222 : 4'b1000;
														assign node4222 = (inp[14]) ? 4'b1001 : 4'b1101;
													assign node4225 = (inp[11]) ? 4'b1101 : node4226;
														assign node4226 = (inp[14]) ? 4'b1100 : 4'b1101;
											assign node4230 = (inp[11]) ? node4236 : node4231;
												assign node4231 = (inp[14]) ? 4'b0000 : node4232;
													assign node4232 = (inp[3]) ? 4'b0001 : 4'b0101;
												assign node4236 = (inp[14]) ? node4238 : 4'b0001;
													assign node4238 = (inp[12]) ? 4'b0101 : node4239;
														assign node4239 = (inp[7]) ? 4'b0001 : 4'b0101;
							assign node4243 = (inp[3]) ? node4245 : 4'b0011;
								assign node4245 = (inp[5]) ? node4247 : 4'b0011;
									assign node4247 = (inp[7]) ? node4271 : node4248;
										assign node4248 = (inp[4]) ? node4254 : node4249;
											assign node4249 = (inp[13]) ? node4251 : 4'b0011;
												assign node4251 = (inp[1]) ? 4'b0001 : 4'b0000;
											assign node4254 = (inp[13]) ? node4264 : node4255;
												assign node4255 = (inp[12]) ? node4261 : node4256;
													assign node4256 = (inp[14]) ? node4258 : 4'b1001;
														assign node4258 = (inp[1]) ? 4'b1000 : 4'b1001;
													assign node4261 = (inp[10]) ? 4'b1001 : 4'b0001;
												assign node4264 = (inp[11]) ? 4'b0000 : node4265;
													assign node4265 = (inp[1]) ? node4267 : 4'b1001;
														assign node4267 = (inp[12]) ? 4'b1001 : 4'b0001;
										assign node4271 = (inp[4]) ? node4273 : 4'b0011;
											assign node4273 = (inp[13]) ? node4275 : 4'b0011;
												assign node4275 = (inp[10]) ? node4277 : 4'b0011;
													assign node4277 = (inp[14]) ? 4'b0000 : 4'b0001;
						assign node4280 = (inp[1]) ? node4586 : node4281;
							assign node4281 = (inp[5]) ? node4419 : node4282;
								assign node4282 = (inp[3]) ? node4340 : node4283;
									assign node4283 = (inp[4]) ? node4309 : node4284;
										assign node4284 = (inp[14]) ? node4296 : node4285;
											assign node4285 = (inp[13]) ? node4291 : node4286;
												assign node4286 = (inp[12]) ? node4288 : 4'b1000;
													assign node4288 = (inp[10]) ? 4'b1000 : 4'b0000;
												assign node4291 = (inp[7]) ? 4'b0000 : node4292;
													assign node4292 = (inp[11]) ? 4'b0100 : 4'b1000;
											assign node4296 = (inp[11]) ? node4304 : node4297;
												assign node4297 = (inp[13]) ? 4'b1001 : node4298;
													assign node4298 = (inp[10]) ? node4300 : 4'b0001;
														assign node4300 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node4304 = (inp[2]) ? node4306 : 4'b1000;
													assign node4306 = (inp[7]) ? 4'b0000 : 4'b1000;
										assign node4309 = (inp[13]) ? node4321 : node4310;
											assign node4310 = (inp[7]) ? node4316 : node4311;
												assign node4311 = (inp[11]) ? 4'b1100 : node4312;
													assign node4312 = (inp[12]) ? 4'b0100 : 4'b1100;
												assign node4316 = (inp[10]) ? 4'b1000 : node4317;
													assign node4317 = (inp[12]) ? 4'b0000 : 4'b1000;
											assign node4321 = (inp[2]) ? node4331 : node4322;
												assign node4322 = (inp[11]) ? node4326 : node4323;
													assign node4323 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node4326 = (inp[12]) ? 4'b1001 : node4327;
														assign node4327 = (inp[10]) ? 4'b0001 : 4'b1001;
												assign node4331 = (inp[12]) ? node4333 : 4'b0100;
													assign node4333 = (inp[10]) ? node4335 : 4'b1100;
														assign node4335 = (inp[14]) ? node4337 : 4'b0100;
															assign node4337 = (inp[11]) ? 4'b0100 : 4'b1001;
									assign node4340 = (inp[13]) ? node4378 : node4341;
										assign node4341 = (inp[2]) ? node4359 : node4342;
											assign node4342 = (inp[11]) ? node4354 : node4343;
												assign node4343 = (inp[4]) ? node4351 : node4344;
													assign node4344 = (inp[7]) ? 4'b1000 : node4345;
														assign node4345 = (inp[10]) ? 4'b0100 : node4346;
															assign node4346 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node4351 = (inp[12]) ? 4'b1100 : 4'b0100;
												assign node4354 = (inp[7]) ? node4356 : 4'b0101;
													assign node4356 = (inp[10]) ? 4'b0001 : 4'b1001;
											assign node4359 = (inp[14]) ? node4369 : node4360;
												assign node4360 = (inp[10]) ? node4364 : node4361;
													assign node4361 = (inp[12]) ? 4'b0100 : 4'b1100;
													assign node4364 = (inp[7]) ? 4'b1100 : node4365;
														assign node4365 = (inp[4]) ? 4'b0000 : 4'b1100;
												assign node4369 = (inp[11]) ? node4371 : 4'b0101;
													assign node4371 = (inp[12]) ? node4375 : node4372;
														assign node4372 = (inp[10]) ? 4'b0001 : 4'b1000;
														assign node4375 = (inp[10]) ? 4'b1100 : 4'b0100;
										assign node4378 = (inp[11]) ? node4402 : node4379;
											assign node4379 = (inp[12]) ? node4395 : node4380;
												assign node4380 = (inp[4]) ? node4390 : node4381;
													assign node4381 = (inp[2]) ? node4385 : node4382;
														assign node4382 = (inp[10]) ? 4'b0100 : 4'b1000;
														assign node4385 = (inp[10]) ? node4387 : 4'b1101;
															assign node4387 = (inp[7]) ? 4'b0101 : 4'b0001;
													assign node4390 = (inp[2]) ? 4'b0000 : node4391;
														assign node4391 = (inp[10]) ? 4'b1001 : 4'b0001;
												assign node4395 = (inp[14]) ? node4399 : node4396;
													assign node4396 = (inp[7]) ? 4'b1100 : 4'b0000;
													assign node4399 = (inp[2]) ? 4'b1101 : 4'b1100;
											assign node4402 = (inp[2]) ? node4414 : node4403;
												assign node4403 = (inp[12]) ? node4407 : node4404;
													assign node4404 = (inp[4]) ? 4'b0000 : 4'b0101;
													assign node4407 = (inp[10]) ? 4'b1101 : node4408;
														assign node4408 = (inp[4]) ? 4'b0101 : node4409;
															assign node4409 = (inp[7]) ? 4'b0001 : 4'b0101;
												assign node4414 = (inp[4]) ? 4'b0001 : node4415;
													assign node4415 = (inp[7]) ? 4'b0100 : 4'b0000;
								assign node4419 = (inp[3]) ? node4513 : node4420;
									assign node4420 = (inp[4]) ? node4474 : node4421;
										assign node4421 = (inp[13]) ? node4443 : node4422;
											assign node4422 = (inp[12]) ? node4432 : node4423;
												assign node4423 = (inp[10]) ? node4425 : 4'b1000;
													assign node4425 = (inp[7]) ? node4429 : node4426;
														assign node4426 = (inp[11]) ? 4'b1100 : 4'b0100;
														assign node4429 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node4432 = (inp[2]) ? node4440 : node4433;
													assign node4433 = (inp[14]) ? node4435 : 4'b0001;
														assign node4435 = (inp[10]) ? node4437 : 4'b0000;
															assign node4437 = (inp[7]) ? 4'b0000 : 4'b0100;
													assign node4440 = (inp[11]) ? 4'b0001 : 4'b0000;
											assign node4443 = (inp[10]) ? node4461 : node4444;
												assign node4444 = (inp[7]) ? node4454 : node4445;
													assign node4445 = (inp[2]) ? node4451 : node4446;
														assign node4446 = (inp[12]) ? 4'b1101 : node4447;
															assign node4447 = (inp[11]) ? 4'b0100 : 4'b0101;
														assign node4451 = (inp[12]) ? 4'b0101 : 4'b1101;
													assign node4454 = (inp[2]) ? node4456 : 4'b0100;
														assign node4456 = (inp[14]) ? 4'b1001 : node4457;
															assign node4457 = (inp[11]) ? 4'b0001 : 4'b0000;
												assign node4461 = (inp[11]) ? 4'b1001 : node4462;
													assign node4462 = (inp[2]) ? node4470 : node4463;
														assign node4463 = (inp[7]) ? node4467 : node4464;
															assign node4464 = (inp[12]) ? 4'b0001 : 4'b1001;
															assign node4467 = (inp[14]) ? 4'b1100 : 4'b1101;
														assign node4470 = (inp[12]) ? 4'b1100 : 4'b0100;
										assign node4474 = (inp[13]) ? node4496 : node4475;
											assign node4475 = (inp[2]) ? node4483 : node4476;
												assign node4476 = (inp[10]) ? 4'b0000 : node4477;
													assign node4477 = (inp[14]) ? node4479 : 4'b1001;
														assign node4479 = (inp[11]) ? 4'b1001 : 4'b0001;
												assign node4483 = (inp[12]) ? node4491 : node4484;
													assign node4484 = (inp[10]) ? node4488 : node4485;
														assign node4485 = (inp[7]) ? 4'b1100 : 4'b1000;
														assign node4488 = (inp[11]) ? 4'b1000 : 4'b0001;
													assign node4491 = (inp[14]) ? 4'b0000 : node4492;
														assign node4492 = (inp[7]) ? 4'b0100 : 4'b0001;
											assign node4496 = (inp[11]) ? node4504 : node4497;
												assign node4497 = (inp[2]) ? 4'b1001 : node4498;
													assign node4498 = (inp[14]) ? node4500 : 4'b0000;
														assign node4500 = (inp[7]) ? 4'b0001 : 4'b0000;
												assign node4504 = (inp[10]) ? 4'b0100 : node4505;
													assign node4505 = (inp[2]) ? node4509 : node4506;
														assign node4506 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node4509 = (inp[7]) ? 4'b0000 : 4'b0100;
									assign node4513 = (inp[14]) ? node4551 : node4514;
										assign node4514 = (inp[4]) ? node4536 : node4515;
											assign node4515 = (inp[12]) ? node4527 : node4516;
												assign node4516 = (inp[10]) ? node4524 : node4517;
													assign node4517 = (inp[7]) ? node4519 : 4'b0000;
														assign node4519 = (inp[13]) ? node4521 : 4'b0001;
															assign node4521 = (inp[2]) ? 4'b0001 : 4'b0000;
													assign node4524 = (inp[7]) ? 4'b0000 : 4'b0001;
												assign node4527 = (inp[10]) ? node4533 : node4528;
													assign node4528 = (inp[2]) ? node4530 : 4'b0000;
														assign node4530 = (inp[11]) ? 4'b1001 : 4'b0001;
													assign node4533 = (inp[7]) ? 4'b0000 : 4'b1000;
											assign node4536 = (inp[13]) ? 4'b0000 : node4537;
												assign node4537 = (inp[12]) ? node4541 : node4538;
													assign node4538 = (inp[11]) ? 4'b1000 : 4'b0000;
													assign node4541 = (inp[10]) ? node4547 : node4542;
														assign node4542 = (inp[7]) ? 4'b0000 : node4543;
															assign node4543 = (inp[2]) ? 4'b1000 : 4'b0000;
														assign node4547 = (inp[11]) ? 4'b0000 : 4'b0001;
										assign node4551 = (inp[4]) ? node4569 : node4552;
											assign node4552 = (inp[2]) ? node4560 : node4553;
												assign node4553 = (inp[10]) ? node4555 : 4'b1001;
													assign node4555 = (inp[11]) ? 4'b0000 : node4556;
														assign node4556 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node4560 = (inp[12]) ? node4564 : node4561;
													assign node4561 = (inp[10]) ? 4'b1001 : 4'b1000;
													assign node4564 = (inp[7]) ? node4566 : 4'b1001;
														assign node4566 = (inp[13]) ? 4'b1001 : 4'b0001;
											assign node4569 = (inp[2]) ? node4577 : node4570;
												assign node4570 = (inp[13]) ? 4'b0000 : node4571;
													assign node4571 = (inp[12]) ? 4'b1000 : node4572;
														assign node4572 = (inp[10]) ? 4'b1000 : 4'b0001;
												assign node4577 = (inp[12]) ? 4'b0001 : node4578;
													assign node4578 = (inp[11]) ? 4'b0000 : node4579;
														assign node4579 = (inp[13]) ? node4581 : 4'b0001;
															assign node4581 = (inp[7]) ? 4'b0001 : 4'b0000;
							assign node4586 = (inp[11]) ? node4760 : node4587;
								assign node4587 = (inp[5]) ? node4671 : node4588;
									assign node4588 = (inp[14]) ? node4628 : node4589;
										assign node4589 = (inp[3]) ? node4611 : node4590;
											assign node4590 = (inp[13]) ? node4596 : node4591;
												assign node4591 = (inp[7]) ? 4'b1001 : node4592;
													assign node4592 = (inp[12]) ? 4'b0101 : 4'b1001;
												assign node4596 = (inp[2]) ? node4604 : node4597;
													assign node4597 = (inp[10]) ? node4601 : node4598;
														assign node4598 = (inp[7]) ? 4'b1001 : 4'b1000;
														assign node4601 = (inp[7]) ? 4'b0001 : 4'b0101;
													assign node4604 = (inp[4]) ? node4608 : node4605;
														assign node4605 = (inp[10]) ? 4'b0001 : 4'b0101;
														assign node4608 = (inp[12]) ? 4'b1101 : 4'b0101;
											assign node4611 = (inp[2]) ? node4621 : node4612;
												assign node4612 = (inp[10]) ? node4616 : node4613;
													assign node4613 = (inp[13]) ? 4'b1100 : 4'b1000;
													assign node4616 = (inp[4]) ? node4618 : 4'b0100;
														assign node4618 = (inp[7]) ? 4'b0100 : 4'b0000;
												assign node4621 = (inp[12]) ? node4625 : node4622;
													assign node4622 = (inp[13]) ? 4'b1000 : 4'b1101;
													assign node4625 = (inp[10]) ? 4'b0101 : 4'b1101;
										assign node4628 = (inp[13]) ? node4646 : node4629;
											assign node4629 = (inp[3]) ? node4635 : node4630;
												assign node4630 = (inp[4]) ? node4632 : 4'b1000;
													assign node4632 = (inp[7]) ? 4'b1000 : 4'b1100;
												assign node4635 = (inp[12]) ? node4641 : node4636;
													assign node4636 = (inp[7]) ? 4'b1100 : node4637;
														assign node4637 = (inp[10]) ? 4'b0100 : 4'b1000;
													assign node4641 = (inp[2]) ? 4'b0100 : node4642;
														assign node4642 = (inp[10]) ? 4'b0100 : 4'b1000;
											assign node4646 = (inp[12]) ? node4658 : node4647;
												assign node4647 = (inp[7]) ? node4651 : node4648;
													assign node4648 = (inp[4]) ? 4'b0001 : 4'b0000;
													assign node4651 = (inp[4]) ? node4655 : node4652;
														assign node4652 = (inp[3]) ? 4'b0100 : 4'b0000;
														assign node4655 = (inp[3]) ? 4'b0000 : 4'b0100;
												assign node4658 = (inp[10]) ? node4668 : node4659;
													assign node4659 = (inp[2]) ? 4'b1000 : node4660;
														assign node4660 = (inp[3]) ? node4662 : 4'b1000;
															assign node4662 = (inp[7]) ? 4'b1100 : node4663;
																assign node4663 = (inp[4]) ? 4'b0001 : 4'b1100;
													assign node4668 = (inp[7]) ? 4'b0000 : 4'b0100;
									assign node4671 = (inp[3]) ? node4725 : node4672;
										assign node4672 = (inp[4]) ? node4694 : node4673;
											assign node4673 = (inp[14]) ? node4687 : node4674;
												assign node4674 = (inp[7]) ? node4678 : node4675;
													assign node4675 = (inp[13]) ? 4'b1100 : 4'b0100;
													assign node4678 = (inp[13]) ? node4684 : node4679;
														assign node4679 = (inp[2]) ? 4'b1000 : node4680;
															assign node4680 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node4684 = (inp[12]) ? 4'b0100 : 4'b1100;
												assign node4687 = (inp[2]) ? 4'b1100 : node4688;
													assign node4688 = (inp[12]) ? 4'b0101 : node4689;
														assign node4689 = (inp[13]) ? 4'b0001 : 4'b1101;
											assign node4694 = (inp[2]) ? node4708 : node4695;
												assign node4695 = (inp[10]) ? node4701 : node4696;
													assign node4696 = (inp[12]) ? 4'b1001 : node4697;
														assign node4697 = (inp[14]) ? 4'b1000 : 4'b1001;
													assign node4701 = (inp[13]) ? 4'b1001 : node4702;
														assign node4702 = (inp[7]) ? 4'b0101 : node4703;
															assign node4703 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node4708 = (inp[14]) ? node4714 : node4709;
													assign node4709 = (inp[10]) ? 4'b0001 : node4710;
														assign node4710 = (inp[12]) ? 4'b0100 : 4'b0000;
													assign node4714 = (inp[7]) ? 4'b0001 : node4715;
														assign node4715 = (inp[10]) ? node4717 : 4'b0001;
															assign node4717 = (inp[13]) ? node4721 : node4718;
																assign node4718 = (inp[12]) ? 4'b0001 : 4'b1001;
																assign node4721 = (inp[12]) ? 4'b1001 : 4'b0001;
										assign node4725 = (inp[4]) ? node4745 : node4726;
											assign node4726 = (inp[10]) ? node4740 : node4727;
												assign node4727 = (inp[13]) ? node4733 : node4728;
													assign node4728 = (inp[12]) ? node4730 : 4'b1000;
														assign node4730 = (inp[7]) ? 4'b1001 : 4'b0001;
													assign node4733 = (inp[14]) ? node4735 : 4'b0000;
														assign node4735 = (inp[7]) ? 4'b0000 : node4736;
															assign node4736 = (inp[2]) ? 4'b0001 : 4'b0000;
												assign node4740 = (inp[2]) ? 4'b1001 : node4741;
													assign node4741 = (inp[14]) ? 4'b0001 : 4'b0000;
											assign node4745 = (inp[14]) ? node4753 : node4746;
												assign node4746 = (inp[12]) ? 4'b0000 : node4747;
													assign node4747 = (inp[7]) ? 4'b0000 : node4748;
														assign node4748 = (inp[10]) ? 4'b0001 : 4'b1000;
												assign node4753 = (inp[10]) ? 4'b0000 : node4754;
													assign node4754 = (inp[12]) ? node4756 : 4'b0001;
														assign node4756 = (inp[13]) ? 4'b0000 : 4'b0001;
								assign node4760 = (inp[5]) ? node4832 : node4761;
									assign node4761 = (inp[10]) ? node4799 : node4762;
										assign node4762 = (inp[3]) ? node4780 : node4763;
											assign node4763 = (inp[4]) ? node4773 : node4764;
												assign node4764 = (inp[7]) ? node4766 : 4'b0001;
													assign node4766 = (inp[13]) ? node4770 : node4767;
														assign node4767 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node4770 = (inp[12]) ? 4'b1001 : 4'b0001;
												assign node4773 = (inp[7]) ? 4'b1001 : node4774;
													assign node4774 = (inp[13]) ? 4'b1001 : node4775;
														assign node4775 = (inp[12]) ? 4'b0101 : 4'b1101;
											assign node4780 = (inp[12]) ? node4788 : node4781;
												assign node4781 = (inp[2]) ? 4'b1001 : node4782;
													assign node4782 = (inp[7]) ? node4784 : 4'b1101;
														assign node4784 = (inp[4]) ? 4'b1101 : 4'b1001;
												assign node4788 = (inp[7]) ? node4796 : node4789;
													assign node4789 = (inp[14]) ? node4791 : 4'b1001;
														assign node4791 = (inp[4]) ? node4793 : 4'b1101;
															assign node4793 = (inp[13]) ? 4'b1001 : 4'b1101;
													assign node4796 = (inp[4]) ? 4'b1101 : 4'b0101;
										assign node4799 = (inp[13]) ? node4815 : node4800;
											assign node4800 = (inp[7]) ? node4810 : node4801;
												assign node4801 = (inp[4]) ? node4805 : node4802;
													assign node4802 = (inp[2]) ? 4'b1101 : 4'b0101;
													assign node4805 = (inp[3]) ? 4'b0001 : node4806;
														assign node4806 = (inp[2]) ? 4'b1101 : 4'b0001;
												assign node4810 = (inp[3]) ? node4812 : 4'b1001;
													assign node4812 = (inp[2]) ? 4'b1101 : 4'b0101;
											assign node4815 = (inp[4]) ? node4827 : node4816;
												assign node4816 = (inp[2]) ? node4818 : 4'b0101;
													assign node4818 = (inp[14]) ? node4820 : 4'b0001;
														assign node4820 = (inp[12]) ? node4822 : 4'b0001;
															assign node4822 = (inp[3]) ? 4'b0101 : node4823;
																assign node4823 = (inp[7]) ? 4'b0001 : 4'b0101;
												assign node4827 = (inp[2]) ? node4829 : 4'b0001;
													assign node4829 = (inp[7]) ? 4'b0001 : 4'b0101;
									assign node4832 = (inp[3]) ? node4864 : node4833;
										assign node4833 = (inp[13]) ? node4845 : node4834;
											assign node4834 = (inp[2]) ? 4'b1001 : node4835;
												assign node4835 = (inp[10]) ? node4839 : node4836;
													assign node4836 = (inp[7]) ? 4'b0001 : 4'b0101;
													assign node4839 = (inp[7]) ? 4'b0101 : node4840;
														assign node4840 = (inp[4]) ? 4'b1001 : 4'b1101;
											assign node4845 = (inp[4]) ? node4853 : node4846;
												assign node4846 = (inp[7]) ? 4'b0101 : node4847;
													assign node4847 = (inp[12]) ? node4849 : 4'b0001;
														assign node4849 = (inp[10]) ? 4'b0001 : 4'b1101;
												assign node4853 = (inp[2]) ? 4'b0001 : node4854;
													assign node4854 = (inp[12]) ? node4860 : node4855;
														assign node4855 = (inp[10]) ? 4'b0001 : node4856;
															assign node4856 = (inp[7]) ? 4'b0001 : 4'b0101;
														assign node4860 = (inp[7]) ? 4'b0001 : 4'b1001;
										assign node4864 = (inp[4]) ? node4874 : node4865;
											assign node4865 = (inp[7]) ? node4867 : 4'b0001;
												assign node4867 = (inp[13]) ? node4871 : node4868;
													assign node4868 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node4871 = (inp[10]) ? 4'b0001 : 4'b1001;
											assign node4874 = (inp[10]) ? node4876 : 4'b0001;
												assign node4876 = (inp[13]) ? 4'b0000 : 4'b0001;
					assign node4879 = (inp[6]) ? node4881 : 4'b0001;
						assign node4881 = (inp[2]) ? node5091 : node4882;
							assign node4882 = (inp[5]) ? node4928 : node4883;
								assign node4883 = (inp[3]) ? node4885 : 4'b0001;
									assign node4885 = (inp[7]) ? node4913 : node4886;
										assign node4886 = (inp[4]) ? node4900 : node4887;
											assign node4887 = (inp[13]) ? node4889 : 4'b0001;
												assign node4889 = (inp[14]) ? node4895 : node4890;
													assign node4890 = (inp[1]) ? 4'b0001 : node4891;
														assign node4891 = (inp[12]) ? 4'b0001 : 4'b0000;
													assign node4895 = (inp[1]) ? node4897 : 4'b0000;
														assign node4897 = (inp[11]) ? 4'b0001 : 4'b0000;
											assign node4900 = (inp[1]) ? node4908 : node4901;
												assign node4901 = (inp[13]) ? node4903 : 4'b1000;
													assign node4903 = (inp[10]) ? 4'b0000 : node4904;
														assign node4904 = (inp[12]) ? 4'b1000 : 4'b0000;
												assign node4908 = (inp[10]) ? 4'b0001 : node4909;
													assign node4909 = (inp[12]) ? 4'b0000 : 4'b1001;
										assign node4913 = (inp[13]) ? node4915 : 4'b0001;
											assign node4915 = (inp[1]) ? 4'b0001 : node4916;
												assign node4916 = (inp[12]) ? node4920 : node4917;
													assign node4917 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node4920 = (inp[14]) ? node4922 : 4'b0001;
														assign node4922 = (inp[10]) ? node4924 : 4'b0001;
															assign node4924 = (inp[11]) ? 4'b0000 : 4'b0001;
								assign node4928 = (inp[1]) ? node5018 : node4929;
									assign node4929 = (inp[3]) ? node4979 : node4930;
										assign node4930 = (inp[14]) ? node4956 : node4931;
											assign node4931 = (inp[10]) ? node4945 : node4932;
												assign node4932 = (inp[4]) ? node4934 : 4'b1000;
													assign node4934 = (inp[12]) ? 4'b1000 : node4935;
														assign node4935 = (inp[11]) ? node4941 : node4936;
															assign node4936 = (inp[7]) ? 4'b1000 : node4937;
																assign node4937 = (inp[13]) ? 4'b1000 : 4'b1100;
															assign node4941 = (inp[13]) ? 4'b0100 : 4'b1100;
												assign node4945 = (inp[13]) ? node4949 : node4946;
													assign node4946 = (inp[11]) ? 4'b1100 : 4'b1000;
													assign node4949 = (inp[7]) ? node4951 : 4'b0100;
														assign node4951 = (inp[12]) ? node4953 : 4'b0000;
															assign node4953 = (inp[4]) ? 4'b0100 : 4'b0000;
											assign node4956 = (inp[11]) ? node4964 : node4957;
												assign node4957 = (inp[12]) ? 4'b1001 : node4958;
													assign node4958 = (inp[7]) ? node4960 : 4'b0101;
														assign node4960 = (inp[13]) ? 4'b0001 : 4'b1001;
												assign node4964 = (inp[7]) ? node4968 : node4965;
													assign node4965 = (inp[4]) ? 4'b1001 : 4'b1000;
													assign node4968 = (inp[12]) ? node4972 : node4969;
														assign node4969 = (inp[13]) ? 4'b0100 : 4'b1000;
														assign node4972 = (inp[4]) ? 4'b1000 : node4973;
															assign node4973 = (inp[13]) ? node4975 : 4'b0000;
																assign node4975 = (inp[10]) ? 4'b0000 : 4'b1000;
										assign node4979 = (inp[13]) ? node4999 : node4980;
											assign node4980 = (inp[10]) ? node4988 : node4981;
												assign node4981 = (inp[4]) ? node4985 : node4982;
													assign node4982 = (inp[14]) ? 4'b0001 : 4'b1001;
													assign node4985 = (inp[7]) ? 4'b1001 : 4'b1000;
												assign node4988 = (inp[11]) ? node4994 : node4989;
													assign node4989 = (inp[12]) ? node4991 : 4'b0000;
														assign node4991 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node4994 = (inp[4]) ? 4'b0001 : node4995;
														assign node4995 = (inp[14]) ? 4'b0001 : 4'b1001;
											assign node4999 = (inp[11]) ? 4'b0000 : node5000;
												assign node5000 = (inp[14]) ? node5006 : node5001;
													assign node5001 = (inp[7]) ? node5003 : 4'b0001;
														assign node5003 = (inp[4]) ? 4'b0000 : 4'b0001;
													assign node5006 = (inp[4]) ? node5012 : node5007;
														assign node5007 = (inp[12]) ? 4'b1000 : node5008;
															assign node5008 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node5012 = (inp[7]) ? 4'b0000 : node5013;
															assign node5013 = (inp[12]) ? 4'b0000 : 4'b0001;
									assign node5018 = (inp[11]) ? node5052 : node5019;
										assign node5019 = (inp[4]) ? node5039 : node5020;
											assign node5020 = (inp[14]) ? node5034 : node5021;
												assign node5021 = (inp[3]) ? node5025 : node5022;
													assign node5022 = (inp[7]) ? 4'b0001 : 4'b0101;
													assign node5025 = (inp[13]) ? node5031 : node5026;
														assign node5026 = (inp[7]) ? 4'b1000 : node5027;
															assign node5027 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node5031 = (inp[10]) ? 4'b1001 : 4'b0001;
												assign node5034 = (inp[7]) ? node5036 : 4'b1000;
													assign node5036 = (inp[12]) ? 4'b1000 : 4'b0000;
											assign node5039 = (inp[10]) ? 4'b0000 : node5040;
												assign node5040 = (inp[3]) ? node5044 : node5041;
													assign node5041 = (inp[7]) ? 4'b0100 : 4'b1000;
													assign node5044 = (inp[13]) ? 4'b0001 : node5045;
														assign node5045 = (inp[14]) ? 4'b0000 : node5046;
															assign node5046 = (inp[7]) ? 4'b0001 : 4'b0000;
										assign node5052 = (inp[3]) ? node5074 : node5053;
											assign node5053 = (inp[13]) ? node5061 : node5054;
												assign node5054 = (inp[12]) ? 4'b0001 : node5055;
													assign node5055 = (inp[14]) ? 4'b1001 : node5056;
														assign node5056 = (inp[7]) ? 4'b1001 : 4'b0001;
												assign node5061 = (inp[12]) ? node5069 : node5062;
													assign node5062 = (inp[7]) ? node5064 : 4'b0101;
														assign node5064 = (inp[10]) ? 4'b0001 : node5065;
															assign node5065 = (inp[4]) ? 4'b0101 : 4'b0001;
													assign node5069 = (inp[10]) ? node5071 : 4'b1001;
														assign node5071 = (inp[4]) ? 4'b0001 : 4'b0101;
											assign node5074 = (inp[7]) ? node5084 : node5075;
												assign node5075 = (inp[14]) ? 4'b0001 : node5076;
													assign node5076 = (inp[13]) ? node5080 : node5077;
														assign node5077 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node5080 = (inp[4]) ? 4'b0000 : 4'b0001;
												assign node5084 = (inp[10]) ? 4'b0001 : node5085;
													assign node5085 = (inp[13]) ? node5087 : 4'b1001;
														assign node5087 = (inp[4]) ? 4'b0001 : 4'b1001;
							assign node5091 = (inp[3]) ? node5093 : 4'b0001;
								assign node5093 = (inp[5]) ? node5095 : 4'b0001;
									assign node5095 = (inp[7]) ? node5117 : node5096;
										assign node5096 = (inp[1]) ? node5110 : node5097;
											assign node5097 = (inp[11]) ? 4'b0000 : node5098;
												assign node5098 = (inp[13]) ? node5104 : node5099;
													assign node5099 = (inp[12]) ? 4'b0001 : node5100;
														assign node5100 = (inp[14]) ? 4'b0000 : 4'b1000;
													assign node5104 = (inp[12]) ? 4'b0000 : node5105;
														assign node5105 = (inp[14]) ? 4'b0000 : 4'b0001;
											assign node5110 = (inp[4]) ? node5112 : 4'b0001;
												assign node5112 = (inp[11]) ? node5114 : 4'b0000;
													assign node5114 = (inp[13]) ? 4'b0000 : 4'b0001;
										assign node5117 = (inp[4]) ? node5119 : 4'b0001;
											assign node5119 = (inp[10]) ? node5121 : 4'b0001;
												assign node5121 = (inp[13]) ? 4'b0000 : 4'b0001;
		assign node5124 = (inp[9]) ? node7832 : node5125;
			assign node5125 = (inp[15]) ? node6567 : node5126;
				assign node5126 = (inp[6]) ? node5520 : node5127;
					assign node5127 = (inp[0]) ? 4'b1100 : node5128;
						assign node5128 = (inp[2]) ? node5386 : node5129;
							assign node5129 = (inp[1]) ? node5243 : node5130;
								assign node5130 = (inp[14]) ? node5186 : node5131;
									assign node5131 = (inp[13]) ? node5167 : node5132;
										assign node5132 = (inp[10]) ? node5146 : node5133;
											assign node5133 = (inp[3]) ? node5141 : node5134;
												assign node5134 = (inp[4]) ? node5138 : node5135;
													assign node5135 = (inp[5]) ? 4'b1101 : 4'b1110;
													assign node5138 = (inp[7]) ? 4'b1101 : 4'b1001;
												assign node5141 = (inp[7]) ? 4'b1001 : node5142;
													assign node5142 = (inp[4]) ? 4'b1101 : 4'b1001;
											assign node5146 = (inp[12]) ? node5162 : node5147;
												assign node5147 = (inp[11]) ? node5153 : node5148;
													assign node5148 = (inp[5]) ? node5150 : 4'b1110;
														assign node5150 = (inp[4]) ? 4'b0101 : 4'b0001;
													assign node5153 = (inp[4]) ? 4'b0001 : node5154;
														assign node5154 = (inp[7]) ? node5158 : node5155;
															assign node5155 = (inp[3]) ? 4'b0101 : 4'b0001;
															assign node5158 = (inp[3]) ? 4'b0001 : 4'b0101;
												assign node5162 = (inp[5]) ? node5164 : 4'b1001;
													assign node5164 = (inp[4]) ? 4'b1101 : 4'b1001;
										assign node5167 = (inp[3]) ? node5177 : node5168;
											assign node5168 = (inp[4]) ? node5172 : node5169;
												assign node5169 = (inp[7]) ? 4'b1110 : 4'b0001;
												assign node5172 = (inp[12]) ? 4'b0001 : node5173;
													assign node5173 = (inp[10]) ? 4'b1001 : 4'b0001;
											assign node5177 = (inp[4]) ? node5181 : node5178;
												assign node5178 = (inp[7]) ? 4'b0001 : 4'b0101;
												assign node5181 = (inp[12]) ? 4'b0101 : node5182;
													assign node5182 = (inp[10]) ? 4'b1101 : 4'b0101;
									assign node5186 = (inp[11]) ? node5218 : node5187;
										assign node5187 = (inp[13]) ? node5201 : node5188;
											assign node5188 = (inp[10]) ? node5198 : node5189;
												assign node5189 = (inp[5]) ? node5193 : node5190;
													assign node5190 = (inp[7]) ? 4'b1110 : 4'b1100;
													assign node5193 = (inp[4]) ? 4'b1000 : node5194;
														assign node5194 = (inp[3]) ? 4'b1000 : 4'b1100;
												assign node5198 = (inp[12]) ? 4'b1000 : 4'b0000;
											assign node5201 = (inp[10]) ? node5207 : node5202;
												assign node5202 = (inp[3]) ? node5204 : 4'b0000;
													assign node5204 = (inp[4]) ? 4'b0100 : 4'b0000;
												assign node5207 = (inp[12]) ? node5211 : node5208;
													assign node5208 = (inp[7]) ? 4'b1000 : 4'b1100;
													assign node5211 = (inp[3]) ? node5215 : node5212;
														assign node5212 = (inp[4]) ? 4'b0000 : 4'b1110;
														assign node5215 = (inp[4]) ? 4'b0100 : 4'b0000;
										assign node5218 = (inp[13]) ? node5232 : node5219;
											assign node5219 = (inp[3]) ? node5227 : node5220;
												assign node5220 = (inp[7]) ? node5224 : node5221;
													assign node5221 = (inp[4]) ? 4'b1001 : 4'b1101;
													assign node5224 = (inp[5]) ? 4'b1101 : 4'b1110;
												assign node5227 = (inp[12]) ? node5229 : 4'b0101;
													assign node5229 = (inp[4]) ? 4'b1101 : 4'b1001;
											assign node5232 = (inp[12]) ? node5236 : node5233;
												assign node5233 = (inp[5]) ? 4'b1001 : 4'b0001;
												assign node5236 = (inp[3]) ? node5238 : 4'b0001;
													assign node5238 = (inp[7]) ? node5240 : 4'b0101;
														assign node5240 = (inp[4]) ? 4'b0101 : 4'b0001;
								assign node5243 = (inp[14]) ? node5307 : node5244;
									assign node5244 = (inp[3]) ? node5274 : node5245;
										assign node5245 = (inp[4]) ? node5263 : node5246;
											assign node5246 = (inp[7]) ? node5256 : node5247;
												assign node5247 = (inp[10]) ? 4'b0000 : node5248;
													assign node5248 = (inp[11]) ? 4'b1000 : node5249;
														assign node5249 = (inp[5]) ? 4'b0000 : node5250;
															assign node5250 = (inp[12]) ? 4'b1110 : 4'b0000;
												assign node5256 = (inp[5]) ? node5258 : 4'b1110;
													assign node5258 = (inp[12]) ? 4'b0100 : node5259;
														assign node5259 = (inp[11]) ? 4'b0100 : 4'b1100;
											assign node5263 = (inp[13]) ? node5269 : node5264;
												assign node5264 = (inp[12]) ? node5266 : 4'b0000;
													assign node5266 = (inp[10]) ? 4'b0000 : 4'b1000;
												assign node5269 = (inp[12]) ? node5271 : 4'b1000;
													assign node5271 = (inp[10]) ? 4'b1000 : 4'b0000;
										assign node5274 = (inp[4]) ? node5294 : node5275;
											assign node5275 = (inp[7]) ? node5285 : node5276;
												assign node5276 = (inp[12]) ? node5280 : node5277;
													assign node5277 = (inp[13]) ? 4'b1100 : 4'b0100;
													assign node5280 = (inp[10]) ? node5282 : 4'b1000;
														assign node5282 = (inp[5]) ? 4'b0100 : 4'b1100;
												assign node5285 = (inp[11]) ? node5287 : 4'b1000;
													assign node5287 = (inp[10]) ? 4'b1000 : node5288;
														assign node5288 = (inp[5]) ? 4'b0000 : node5289;
															assign node5289 = (inp[12]) ? 4'b1000 : 4'b0000;
											assign node5294 = (inp[10]) ? node5304 : node5295;
												assign node5295 = (inp[13]) ? node5301 : node5296;
													assign node5296 = (inp[12]) ? node5298 : 4'b0100;
														assign node5298 = (inp[7]) ? 4'b1000 : 4'b1100;
													assign node5301 = (inp[12]) ? 4'b0100 : 4'b1100;
												assign node5304 = (inp[13]) ? 4'b1100 : 4'b0100;
									assign node5307 = (inp[11]) ? node5351 : node5308;
										assign node5308 = (inp[13]) ? node5326 : node5309;
											assign node5309 = (inp[3]) ? node5319 : node5310;
												assign node5310 = (inp[5]) ? node5316 : node5311;
													assign node5311 = (inp[7]) ? 4'b1110 : node5312;
														assign node5312 = (inp[10]) ? 4'b1001 : 4'b1110;
													assign node5316 = (inp[12]) ? 4'b1101 : 4'b0101;
												assign node5319 = (inp[7]) ? 4'b1001 : node5320;
													assign node5320 = (inp[10]) ? 4'b0101 : node5321;
														assign node5321 = (inp[4]) ? 4'b1101 : 4'b1001;
											assign node5326 = (inp[10]) ? node5342 : node5327;
												assign node5327 = (inp[12]) ? node5337 : node5328;
													assign node5328 = (inp[7]) ? node5330 : 4'b0101;
														assign node5330 = (inp[3]) ? node5334 : node5331;
															assign node5331 = (inp[4]) ? 4'b0001 : 4'b0101;
															assign node5334 = (inp[4]) ? 4'b0101 : 4'b0001;
													assign node5337 = (inp[4]) ? 4'b0001 : node5338;
														assign node5338 = (inp[7]) ? 4'b0101 : 4'b0001;
												assign node5342 = (inp[12]) ? 4'b0001 : node5343;
													assign node5343 = (inp[3]) ? node5345 : 4'b1001;
														assign node5345 = (inp[7]) ? node5347 : 4'b1101;
															assign node5347 = (inp[5]) ? 4'b1101 : 4'b1001;
										assign node5351 = (inp[12]) ? node5365 : node5352;
											assign node5352 = (inp[13]) ? node5358 : node5353;
												assign node5353 = (inp[5]) ? node5355 : 4'b0000;
													assign node5355 = (inp[4]) ? 4'b0000 : 4'b0100;
												assign node5358 = (inp[3]) ? 4'b1100 : node5359;
													assign node5359 = (inp[10]) ? 4'b1000 : node5360;
														assign node5360 = (inp[4]) ? 4'b1000 : 4'b1100;
											assign node5365 = (inp[5]) ? node5373 : node5366;
												assign node5366 = (inp[7]) ? node5370 : node5367;
													assign node5367 = (inp[3]) ? 4'b1100 : 4'b1000;
													assign node5370 = (inp[10]) ? 4'b1110 : 4'b1000;
												assign node5373 = (inp[4]) ? node5383 : node5374;
													assign node5374 = (inp[3]) ? node5376 : 4'b1100;
														assign node5376 = (inp[10]) ? node5380 : node5377;
															assign node5377 = (inp[13]) ? 4'b0000 : 4'b1000;
															assign node5380 = (inp[13]) ? 4'b1100 : 4'b0100;
													assign node5383 = (inp[3]) ? 4'b0100 : 4'b0000;
							assign node5386 = (inp[5]) ? node5388 : 4'b1110;
								assign node5388 = (inp[3]) ? node5446 : node5389;
									assign node5389 = (inp[4]) ? node5411 : node5390;
										assign node5390 = (inp[7]) ? 4'b1110 : node5391;
											assign node5391 = (inp[13]) ? node5405 : node5392;
												assign node5392 = (inp[1]) ? node5394 : 4'b1110;
													assign node5394 = (inp[11]) ? node5400 : node5395;
														assign node5395 = (inp[12]) ? 4'b1110 : node5396;
															assign node5396 = (inp[10]) ? 4'b0001 : 4'b1110;
														assign node5400 = (inp[10]) ? 4'b0000 : node5401;
															assign node5401 = (inp[12]) ? 4'b1110 : 4'b0000;
												assign node5405 = (inp[14]) ? 4'b0001 : node5406;
													assign node5406 = (inp[1]) ? 4'b1000 : 4'b0001;
										assign node5411 = (inp[1]) ? node5431 : node5412;
											assign node5412 = (inp[13]) ? node5422 : node5413;
												assign node5413 = (inp[7]) ? node5417 : node5414;
													assign node5414 = (inp[14]) ? 4'b0001 : 4'b1001;
													assign node5417 = (inp[12]) ? 4'b1110 : node5418;
														assign node5418 = (inp[10]) ? 4'b0001 : 4'b1110;
												assign node5422 = (inp[10]) ? node5428 : node5423;
													assign node5423 = (inp[14]) ? node5425 : 4'b0001;
														assign node5425 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node5428 = (inp[12]) ? 4'b0001 : 4'b1001;
											assign node5431 = (inp[11]) ? node5441 : node5432;
												assign node5432 = (inp[7]) ? node5434 : 4'b1001;
													assign node5434 = (inp[12]) ? node5438 : node5435;
														assign node5435 = (inp[13]) ? 4'b1000 : 4'b0000;
														assign node5438 = (inp[13]) ? 4'b0001 : 4'b1110;
												assign node5441 = (inp[13]) ? node5443 : 4'b0000;
													assign node5443 = (inp[12]) ? 4'b0000 : 4'b1000;
									assign node5446 = (inp[4]) ? node5488 : node5447;
										assign node5447 = (inp[7]) ? node5471 : node5448;
											assign node5448 = (inp[13]) ? node5456 : node5449;
												assign node5449 = (inp[14]) ? node5453 : node5450;
													assign node5450 = (inp[11]) ? 4'b0101 : 4'b0100;
													assign node5453 = (inp[11]) ? 4'b1001 : 4'b1000;
												assign node5456 = (inp[12]) ? node5464 : node5457;
													assign node5457 = (inp[11]) ? 4'b1100 : node5458;
														assign node5458 = (inp[10]) ? node5460 : 4'b0101;
															assign node5460 = (inp[14]) ? 4'b1100 : 4'b1101;
													assign node5464 = (inp[1]) ? node5466 : 4'b0101;
														assign node5466 = (inp[11]) ? 4'b1100 : node5467;
															assign node5467 = (inp[14]) ? 4'b0101 : 4'b0100;
											assign node5471 = (inp[1]) ? node5481 : node5472;
												assign node5472 = (inp[13]) ? node5476 : node5473;
													assign node5473 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node5476 = (inp[12]) ? 4'b0001 : node5477;
														assign node5477 = (inp[10]) ? 4'b1001 : 4'b0001;
												assign node5481 = (inp[11]) ? node5485 : node5482;
													assign node5482 = (inp[14]) ? 4'b1001 : 4'b1000;
													assign node5485 = (inp[13]) ? 4'b1000 : 4'b0000;
										assign node5488 = (inp[1]) ? node5506 : node5489;
											assign node5489 = (inp[13]) ? node5503 : node5490;
												assign node5490 = (inp[12]) ? node5498 : node5491;
													assign node5491 = (inp[10]) ? node5493 : 4'b1101;
														assign node5493 = (inp[7]) ? 4'b0101 : node5494;
															assign node5494 = (inp[11]) ? 4'b0101 : 4'b0100;
													assign node5498 = (inp[7]) ? 4'b1001 : node5499;
														assign node5499 = (inp[10]) ? 4'b1101 : 4'b1100;
												assign node5503 = (inp[14]) ? 4'b0100 : 4'b0101;
											assign node5506 = (inp[13]) ? node5514 : node5507;
												assign node5507 = (inp[11]) ? 4'b0100 : node5508;
													assign node5508 = (inp[14]) ? 4'b1101 : node5509;
														assign node5509 = (inp[10]) ? 4'b0100 : 4'b1100;
												assign node5514 = (inp[12]) ? node5516 : 4'b1100;
													assign node5516 = (inp[10]) ? 4'b1100 : 4'b0100;
					assign node5520 = (inp[5]) ? node5984 : node5521;
						assign node5521 = (inp[0]) ? node5861 : node5522;
							assign node5522 = (inp[11]) ? node5700 : node5523;
								assign node5523 = (inp[13]) ? node5613 : node5524;
									assign node5524 = (inp[4]) ? node5558 : node5525;
										assign node5525 = (inp[12]) ? node5543 : node5526;
											assign node5526 = (inp[7]) ? node5534 : node5527;
												assign node5527 = (inp[1]) ? node5529 : 4'b0001;
													assign node5529 = (inp[3]) ? node5531 : 4'b1101;
														assign node5531 = (inp[10]) ? 4'b1001 : 4'b0001;
												assign node5534 = (inp[3]) ? 4'b0000 : node5535;
													assign node5535 = (inp[1]) ? node5539 : node5536;
														assign node5536 = (inp[14]) ? 4'b1100 : 4'b1101;
														assign node5539 = (inp[10]) ? 4'b0101 : 4'b0100;
											assign node5543 = (inp[3]) ? node5551 : node5544;
												assign node5544 = (inp[14]) ? node5548 : node5545;
													assign node5545 = (inp[1]) ? 4'b1100 : 4'b1101;
													assign node5548 = (inp[1]) ? 4'b1101 : 4'b1100;
												assign node5551 = (inp[10]) ? node5555 : node5552;
													assign node5552 = (inp[2]) ? 4'b1000 : 4'b1101;
													assign node5555 = (inp[7]) ? 4'b0101 : 4'b0001;
										assign node5558 = (inp[10]) ? node5580 : node5559;
											assign node5559 = (inp[3]) ? node5569 : node5560;
												assign node5560 = (inp[7]) ? node5566 : node5561;
													assign node5561 = (inp[1]) ? 4'b1001 : node5562;
														assign node5562 = (inp[14]) ? 4'b1000 : 4'b1001;
													assign node5566 = (inp[2]) ? 4'b1101 : 4'b1001;
												assign node5569 = (inp[1]) ? node5577 : node5570;
													assign node5570 = (inp[14]) ? 4'b1001 : node5571;
														assign node5571 = (inp[2]) ? 4'b1001 : node5572;
															assign node5572 = (inp[12]) ? 4'b1000 : 4'b0000;
													assign node5577 = (inp[14]) ? 4'b0000 : 4'b0001;
											assign node5580 = (inp[7]) ? node5600 : node5581;
												assign node5581 = (inp[14]) ? node5591 : node5582;
													assign node5582 = (inp[12]) ? 4'b0101 : node5583;
														assign node5583 = (inp[1]) ? node5585 : 4'b1000;
															assign node5585 = (inp[3]) ? node5587 : 4'b1101;
																assign node5587 = (inp[2]) ? 4'b1101 : 4'b0101;
													assign node5591 = (inp[3]) ? node5593 : 4'b1000;
														assign node5593 = (inp[2]) ? 4'b0101 : node5594;
															assign node5594 = (inp[1]) ? node5596 : 4'b0001;
																assign node5596 = (inp[12]) ? 4'b1000 : 4'b0100;
												assign node5600 = (inp[3]) ? node5606 : node5601;
													assign node5601 = (inp[12]) ? 4'b1100 : node5602;
														assign node5602 = (inp[1]) ? 4'b0000 : 4'b0001;
													assign node5606 = (inp[1]) ? node5610 : node5607;
														assign node5607 = (inp[12]) ? 4'b1000 : 4'b1001;
														assign node5610 = (inp[14]) ? 4'b0001 : 4'b1001;
									assign node5613 = (inp[4]) ? node5665 : node5614;
										assign node5614 = (inp[7]) ? node5640 : node5615;
											assign node5615 = (inp[10]) ? node5629 : node5616;
												assign node5616 = (inp[3]) ? node5624 : node5617;
													assign node5617 = (inp[14]) ? 4'b0001 : node5618;
														assign node5618 = (inp[12]) ? 4'b0001 : node5619;
															assign node5619 = (inp[1]) ? 4'b1000 : 4'b1001;
													assign node5624 = (inp[12]) ? 4'b1001 : node5625;
														assign node5625 = (inp[1]) ? 4'b0001 : 4'b1001;
												assign node5629 = (inp[1]) ? node5635 : node5630;
													assign node5630 = (inp[3]) ? 4'b0000 : node5631;
														assign node5631 = (inp[12]) ? 4'b0000 : 4'b0001;
													assign node5635 = (inp[2]) ? node5637 : 4'b0000;
														assign node5637 = (inp[14]) ? 4'b1001 : 4'b1000;
											assign node5640 = (inp[2]) ? node5652 : node5641;
												assign node5641 = (inp[10]) ? node5647 : node5642;
													assign node5642 = (inp[1]) ? node5644 : 4'b1101;
														assign node5644 = (inp[12]) ? 4'b0101 : 4'b0001;
													assign node5647 = (inp[1]) ? node5649 : 4'b0001;
														assign node5649 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node5652 = (inp[3]) ? node5658 : node5653;
													assign node5653 = (inp[10]) ? 4'b0101 : node5654;
														assign node5654 = (inp[12]) ? 4'b0100 : 4'b1100;
													assign node5658 = (inp[10]) ? 4'b0001 : node5659;
														assign node5659 = (inp[1]) ? node5661 : 4'b0000;
															assign node5661 = (inp[14]) ? 4'b0001 : 4'b0000;
										assign node5665 = (inp[7]) ? node5689 : node5666;
											assign node5666 = (inp[2]) ? node5680 : node5667;
												assign node5667 = (inp[3]) ? node5675 : node5668;
													assign node5668 = (inp[10]) ? node5670 : 4'b1101;
														assign node5670 = (inp[12]) ? 4'b0101 : node5671;
															assign node5671 = (inp[14]) ? 4'b0101 : 4'b1101;
													assign node5675 = (inp[10]) ? node5677 : 4'b0101;
														assign node5677 = (inp[14]) ? 4'b1101 : 4'b0101;
												assign node5680 = (inp[12]) ? node5686 : node5681;
													assign node5681 = (inp[1]) ? node5683 : 4'b1001;
														assign node5683 = (inp[10]) ? 4'b1101 : 4'b0101;
													assign node5686 = (inp[1]) ? 4'b0001 : 4'b0000;
											assign node5689 = (inp[10]) ? node5697 : node5690;
												assign node5690 = (inp[3]) ? node5694 : node5691;
													assign node5691 = (inp[1]) ? 4'b0101 : 4'b1001;
													assign node5694 = (inp[12]) ? 4'b1001 : 4'b1000;
												assign node5697 = (inp[12]) ? 4'b0101 : 4'b1001;
								assign node5700 = (inp[1]) ? node5790 : node5701;
									assign node5701 = (inp[13]) ? node5737 : node5702;
										assign node5702 = (inp[4]) ? node5720 : node5703;
											assign node5703 = (inp[2]) ? node5713 : node5704;
												assign node5704 = (inp[7]) ? node5710 : node5705;
													assign node5705 = (inp[3]) ? 4'b1100 : node5706;
														assign node5706 = (inp[14]) ? 4'b0000 : 4'b1000;
													assign node5710 = (inp[3]) ? 4'b1100 : 4'b1101;
												assign node5713 = (inp[3]) ? 4'b1001 : node5714;
													assign node5714 = (inp[10]) ? node5716 : 4'b1101;
														assign node5716 = (inp[12]) ? 4'b1101 : 4'b0101;
											assign node5720 = (inp[10]) ? node5732 : node5721;
												assign node5721 = (inp[12]) ? node5727 : node5722;
													assign node5722 = (inp[3]) ? 4'b0100 : node5723;
														assign node5723 = (inp[7]) ? 4'b0000 : 4'b1001;
													assign node5727 = (inp[3]) ? node5729 : 4'b1000;
														assign node5729 = (inp[14]) ? 4'b1000 : 4'b1001;
												assign node5732 = (inp[12]) ? 4'b1101 : node5733;
													assign node5733 = (inp[7]) ? 4'b1000 : 4'b1100;
										assign node5737 = (inp[4]) ? node5765 : node5738;
											assign node5738 = (inp[2]) ? node5754 : node5739;
												assign node5739 = (inp[12]) ? node5747 : node5740;
													assign node5740 = (inp[10]) ? node5742 : 4'b0000;
														assign node5742 = (inp[7]) ? 4'b1000 : node5743;
															assign node5743 = (inp[3]) ? 4'b0001 : 4'b1000;
													assign node5747 = (inp[3]) ? node5751 : node5748;
														assign node5748 = (inp[7]) ? 4'b0101 : 4'b0000;
														assign node5751 = (inp[7]) ? 4'b1100 : 4'b1000;
												assign node5754 = (inp[3]) ? node5758 : node5755;
													assign node5755 = (inp[7]) ? 4'b0101 : 4'b0001;
													assign node5758 = (inp[14]) ? node5760 : 4'b0000;
														assign node5760 = (inp[7]) ? node5762 : 4'b1000;
															assign node5762 = (inp[12]) ? 4'b0001 : 4'b0000;
											assign node5765 = (inp[12]) ? node5775 : node5766;
												assign node5766 = (inp[3]) ? node5770 : node5767;
													assign node5767 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node5770 = (inp[2]) ? 4'b0100 : node5771;
														assign node5771 = (inp[14]) ? 4'b1001 : 4'b0101;
												assign node5775 = (inp[10]) ? node5783 : node5776;
													assign node5776 = (inp[7]) ? node5778 : 4'b1100;
														assign node5778 = (inp[2]) ? 4'b1000 : node5779;
															assign node5779 = (inp[3]) ? 4'b0001 : 4'b1000;
													assign node5783 = (inp[2]) ? node5787 : node5784;
														assign node5784 = (inp[3]) ? 4'b0101 : 4'b0100;
														assign node5787 = (inp[7]) ? 4'b0001 : 4'b0100;
									assign node5790 = (inp[10]) ? node5838 : node5791;
										assign node5791 = (inp[7]) ? node5811 : node5792;
											assign node5792 = (inp[4]) ? node5800 : node5793;
												assign node5793 = (inp[12]) ? 4'b0000 : node5794;
													assign node5794 = (inp[3]) ? 4'b0000 : node5795;
														assign node5795 = (inp[13]) ? 4'b1000 : 4'b0000;
												assign node5800 = (inp[3]) ? node5808 : node5801;
													assign node5801 = (inp[2]) ? node5803 : 4'b0100;
														assign node5803 = (inp[13]) ? 4'b0000 : node5804;
															assign node5804 = (inp[12]) ? 4'b1000 : 4'b0000;
													assign node5808 = (inp[2]) ? 4'b0100 : 4'b0000;
											assign node5811 = (inp[12]) ? node5825 : node5812;
												assign node5812 = (inp[14]) ? node5822 : node5813;
													assign node5813 = (inp[2]) ? 4'b0100 : node5814;
														assign node5814 = (inp[13]) ? node5818 : node5815;
															assign node5815 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node5818 = (inp[4]) ? 4'b0100 : 4'b0000;
													assign node5822 = (inp[3]) ? 4'b0000 : 4'b0100;
												assign node5825 = (inp[14]) ? node5833 : node5826;
													assign node5826 = (inp[2]) ? 4'b0000 : node5827;
														assign node5827 = (inp[13]) ? node5829 : 4'b0000;
															assign node5829 = (inp[4]) ? 4'b0100 : 4'b0000;
													assign node5833 = (inp[4]) ? node5835 : 4'b0100;
														assign node5835 = (inp[3]) ? 4'b1000 : 4'b0000;
										assign node5838 = (inp[4]) ? node5846 : node5839;
											assign node5839 = (inp[3]) ? 4'b1000 : node5840;
												assign node5840 = (inp[7]) ? node5842 : 4'b1000;
													assign node5842 = (inp[13]) ? 4'b1100 : 4'b0100;
											assign node5846 = (inp[7]) ? node5854 : node5847;
												assign node5847 = (inp[3]) ? 4'b1100 : node5848;
													assign node5848 = (inp[2]) ? node5850 : 4'b1100;
														assign node5850 = (inp[13]) ? 4'b1000 : 4'b0000;
												assign node5854 = (inp[13]) ? 4'b1000 : node5855;
													assign node5855 = (inp[2]) ? 4'b0000 : node5856;
														assign node5856 = (inp[3]) ? 4'b0000 : 4'b1000;
							assign node5861 = (inp[2]) ? 4'b1100 : node5862;
								assign node5862 = (inp[4]) ? node5914 : node5863;
									assign node5863 = (inp[3]) ? node5883 : node5864;
										assign node5864 = (inp[7]) ? 4'b1100 : node5865;
											assign node5865 = (inp[13]) ? node5873 : node5866;
												assign node5866 = (inp[14]) ? 4'b1100 : node5867;
													assign node5867 = (inp[12]) ? 4'b1100 : node5868;
														assign node5868 = (inp[10]) ? 4'b0001 : 4'b0000;
												assign node5873 = (inp[1]) ? node5879 : node5874;
													assign node5874 = (inp[11]) ? 4'b0001 : node5875;
														assign node5875 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node5879 = (inp[10]) ? 4'b1000 : 4'b0000;
										assign node5883 = (inp[7]) ? node5901 : node5884;
											assign node5884 = (inp[13]) ? node5894 : node5885;
												assign node5885 = (inp[10]) ? node5891 : node5886;
													assign node5886 = (inp[12]) ? node5888 : 4'b1001;
														assign node5888 = (inp[1]) ? 4'b1001 : 4'b1000;
													assign node5891 = (inp[12]) ? 4'b1001 : 4'b0100;
												assign node5894 = (inp[11]) ? node5898 : node5895;
													assign node5895 = (inp[14]) ? 4'b0101 : 4'b0100;
													assign node5898 = (inp[12]) ? 4'b0100 : 4'b1100;
											assign node5901 = (inp[1]) ? node5907 : node5902;
												assign node5902 = (inp[11]) ? node5904 : 4'b1000;
													assign node5904 = (inp[13]) ? 4'b0001 : 4'b1001;
												assign node5907 = (inp[14]) ? node5911 : node5908;
													assign node5908 = (inp[13]) ? 4'b1000 : 4'b0000;
													assign node5911 = (inp[11]) ? 4'b1000 : 4'b1001;
									assign node5914 = (inp[3]) ? node5952 : node5915;
										assign node5915 = (inp[13]) ? node5935 : node5916;
											assign node5916 = (inp[7]) ? node5922 : node5917;
												assign node5917 = (inp[12]) ? node5919 : 4'b1001;
													assign node5919 = (inp[14]) ? 4'b1000 : 4'b1001;
												assign node5922 = (inp[10]) ? node5928 : node5923;
													assign node5923 = (inp[14]) ? 4'b1100 : node5924;
														assign node5924 = (inp[1]) ? 4'b0000 : 4'b1100;
													assign node5928 = (inp[12]) ? 4'b1100 : node5929;
														assign node5929 = (inp[1]) ? node5931 : 4'b0001;
															assign node5931 = (inp[14]) ? 4'b0001 : 4'b0000;
											assign node5935 = (inp[12]) ? node5943 : node5936;
												assign node5936 = (inp[1]) ? 4'b1000 : node5937;
													assign node5937 = (inp[11]) ? 4'b0001 : node5938;
														assign node5938 = (inp[10]) ? 4'b1000 : 4'b0000;
												assign node5943 = (inp[1]) ? node5949 : node5944;
													assign node5944 = (inp[11]) ? 4'b0001 : node5945;
														assign node5945 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node5949 = (inp[11]) ? 4'b0000 : 4'b0001;
										assign node5952 = (inp[13]) ? node5968 : node5953;
											assign node5953 = (inp[1]) ? node5963 : node5954;
												assign node5954 = (inp[7]) ? node5960 : node5955;
													assign node5955 = (inp[10]) ? 4'b0100 : node5956;
														assign node5956 = (inp[11]) ? 4'b1101 : 4'b1100;
													assign node5960 = (inp[11]) ? 4'b1001 : 4'b1000;
												assign node5963 = (inp[12]) ? 4'b1100 : node5964;
													assign node5964 = (inp[11]) ? 4'b0100 : 4'b0101;
											assign node5968 = (inp[12]) ? node5974 : node5969;
												assign node5969 = (inp[14]) ? node5971 : 4'b1100;
													assign node5971 = (inp[10]) ? 4'b1100 : 4'b0101;
												assign node5974 = (inp[1]) ? node5980 : node5975;
													assign node5975 = (inp[10]) ? node5977 : 4'b0101;
														assign node5977 = (inp[11]) ? 4'b0101 : 4'b0100;
													assign node5980 = (inp[11]) ? 4'b0100 : 4'b0101;
						assign node5984 = (inp[3]) ? node6302 : node5985;
							assign node5985 = (inp[4]) ? node6119 : node5986;
								assign node5986 = (inp[7]) ? node6064 : node5987;
									assign node5987 = (inp[11]) ? node6031 : node5988;
										assign node5988 = (inp[13]) ? node6010 : node5989;
											assign node5989 = (inp[10]) ? node5999 : node5990;
												assign node5990 = (inp[14]) ? node5994 : node5991;
													assign node5991 = (inp[12]) ? 4'b1100 : 4'b1000;
													assign node5994 = (inp[12]) ? node5996 : 4'b1100;
														assign node5996 = (inp[2]) ? 4'b1100 : 4'b1101;
												assign node5999 = (inp[0]) ? node6005 : node6000;
													assign node6000 = (inp[12]) ? node6002 : 4'b1000;
														assign node6002 = (inp[2]) ? 4'b1000 : 4'b0000;
													assign node6005 = (inp[12]) ? node6007 : 4'b0001;
														assign node6007 = (inp[14]) ? 4'b1100 : 4'b0001;
											assign node6010 = (inp[0]) ? node6020 : node6011;
												assign node6011 = (inp[2]) ? node6013 : 4'b0100;
													assign node6013 = (inp[1]) ? node6017 : node6014;
														assign node6014 = (inp[10]) ? 4'b0101 : 4'b0001;
														assign node6017 = (inp[14]) ? 4'b1100 : 4'b1101;
												assign node6020 = (inp[2]) ? node6026 : node6021;
													assign node6021 = (inp[12]) ? 4'b1001 : node6022;
														assign node6022 = (inp[14]) ? 4'b0001 : 4'b1001;
													assign node6026 = (inp[14]) ? 4'b0000 : node6027;
														assign node6027 = (inp[12]) ? 4'b0000 : 4'b1000;
										assign node6031 = (inp[1]) ? node6051 : node6032;
											assign node6032 = (inp[2]) ? node6042 : node6033;
												assign node6033 = (inp[0]) ? node6037 : node6034;
													assign node6034 = (inp[13]) ? 4'b0001 : 4'b0000;
													assign node6037 = (inp[12]) ? node6039 : 4'b1000;
														assign node6039 = (inp[10]) ? 4'b0000 : 4'b1000;
												assign node6042 = (inp[13]) ? node6046 : node6043;
													assign node6043 = (inp[10]) ? 4'b1001 : 4'b1100;
													assign node6046 = (inp[10]) ? 4'b0101 : node6047;
														assign node6047 = (inp[0]) ? 4'b0001 : 4'b1001;
											assign node6051 = (inp[13]) ? 4'b1000 : node6052;
												assign node6052 = (inp[2]) ? node6058 : node6053;
													assign node6053 = (inp[12]) ? 4'b1000 : node6054;
														assign node6054 = (inp[14]) ? 4'b1000 : 4'b0000;
													assign node6058 = (inp[14]) ? 4'b0000 : node6059;
														assign node6059 = (inp[10]) ? 4'b0000 : 4'b1000;
									assign node6064 = (inp[2]) ? node6094 : node6065;
										assign node6065 = (inp[10]) ? node6081 : node6066;
											assign node6066 = (inp[13]) ? node6076 : node6067;
												assign node6067 = (inp[1]) ? node6069 : 4'b1101;
													assign node6069 = (inp[0]) ? node6073 : node6070;
														assign node6070 = (inp[11]) ? 4'b0100 : 4'b0101;
														assign node6073 = (inp[14]) ? 4'b1101 : 4'b1100;
												assign node6076 = (inp[0]) ? node6078 : 4'b1000;
													assign node6078 = (inp[12]) ? 4'b0101 : 4'b0001;
											assign node6081 = (inp[13]) ? node6089 : node6082;
												assign node6082 = (inp[0]) ? node6084 : 4'b0000;
													assign node6084 = (inp[1]) ? 4'b0100 : node6085;
														assign node6085 = (inp[14]) ? 4'b0100 : 4'b0101;
												assign node6089 = (inp[1]) ? node6091 : 4'b0100;
													assign node6091 = (inp[12]) ? 4'b0100 : 4'b1100;
										assign node6094 = (inp[0]) ? 4'b1100 : node6095;
											assign node6095 = (inp[13]) ? node6109 : node6096;
												assign node6096 = (inp[11]) ? node6100 : node6097;
													assign node6097 = (inp[1]) ? 4'b0101 : 4'b1101;
													assign node6100 = (inp[1]) ? node6106 : node6101;
														assign node6101 = (inp[14]) ? 4'b1100 : node6102;
															assign node6102 = (inp[12]) ? 4'b1100 : 4'b0100;
														assign node6106 = (inp[12]) ? 4'b0100 : 4'b0000;
												assign node6109 = (inp[10]) ? node6115 : node6110;
													assign node6110 = (inp[1]) ? 4'b1001 : node6111;
														assign node6111 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node6115 = (inp[11]) ? 4'b1000 : 4'b0000;
								assign node6119 = (inp[2]) ? node6211 : node6120;
									assign node6120 = (inp[11]) ? node6178 : node6121;
										assign node6121 = (inp[10]) ? node6149 : node6122;
											assign node6122 = (inp[7]) ? node6134 : node6123;
												assign node6123 = (inp[14]) ? node6131 : node6124;
													assign node6124 = (inp[12]) ? 4'b1000 : node6125;
														assign node6125 = (inp[0]) ? node6127 : 4'b1001;
															assign node6127 = (inp[13]) ? 4'b1000 : 4'b1001;
													assign node6131 = (inp[0]) ? 4'b1000 : 4'b0000;
												assign node6134 = (inp[14]) ? node6140 : node6135;
													assign node6135 = (inp[13]) ? node6137 : 4'b0001;
														assign node6137 = (inp[1]) ? 4'b1001 : 4'b0001;
													assign node6140 = (inp[13]) ? node6142 : 4'b1001;
														assign node6142 = (inp[0]) ? node6146 : node6143;
															assign node6143 = (inp[1]) ? 4'b1001 : 4'b0001;
															assign node6146 = (inp[1]) ? 4'b0101 : 4'b1001;
											assign node6149 = (inp[0]) ? node6167 : node6150;
												assign node6150 = (inp[14]) ? node6160 : node6151;
													assign node6151 = (inp[7]) ? node6157 : node6152;
														assign node6152 = (inp[13]) ? 4'b1000 : node6153;
															assign node6153 = (inp[1]) ? 4'b0001 : 4'b0101;
														assign node6157 = (inp[1]) ? 4'b1000 : 4'b1001;
													assign node6160 = (inp[13]) ? node6164 : node6161;
														assign node6161 = (inp[1]) ? 4'b0001 : 4'b0000;
														assign node6164 = (inp[1]) ? 4'b0000 : 4'b0001;
												assign node6167 = (inp[1]) ? node6175 : node6168;
													assign node6168 = (inp[12]) ? node6170 : 4'b0001;
														assign node6170 = (inp[13]) ? node6172 : 4'b0101;
															assign node6172 = (inp[7]) ? 4'b0101 : 4'b1001;
													assign node6175 = (inp[12]) ? 4'b0001 : 4'b1001;
										assign node6178 = (inp[10]) ? node6192 : node6179;
											assign node6179 = (inp[0]) ? node6185 : node6180;
												assign node6180 = (inp[13]) ? 4'b0000 : node6181;
													assign node6181 = (inp[12]) ? 4'b0001 : 4'b0000;
												assign node6185 = (inp[7]) ? node6187 : 4'b0100;
													assign node6187 = (inp[12]) ? node6189 : 4'b0000;
														assign node6189 = (inp[1]) ? 4'b0100 : 4'b1000;
											assign node6192 = (inp[1]) ? node6206 : node6193;
												assign node6193 = (inp[0]) ? node6199 : node6194;
													assign node6194 = (inp[12]) ? node6196 : 4'b1001;
														assign node6196 = (inp[13]) ? 4'b1001 : 4'b0001;
													assign node6199 = (inp[13]) ? 4'b0001 : node6200;
														assign node6200 = (inp[12]) ? node6202 : 4'b1100;
															assign node6202 = (inp[7]) ? 4'b0000 : 4'b0100;
												assign node6206 = (inp[7]) ? 4'b1000 : node6207;
													assign node6207 = (inp[0]) ? 4'b0000 : 4'b1000;
									assign node6211 = (inp[1]) ? node6257 : node6212;
										assign node6212 = (inp[11]) ? node6238 : node6213;
											assign node6213 = (inp[12]) ? node6227 : node6214;
												assign node6214 = (inp[7]) ? node6220 : node6215;
													assign node6215 = (inp[0]) ? node6217 : 4'b0100;
														assign node6217 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node6220 = (inp[10]) ? node6224 : node6221;
														assign node6221 = (inp[0]) ? 4'b1100 : 4'b1001;
														assign node6224 = (inp[0]) ? 4'b0000 : 4'b0100;
												assign node6227 = (inp[13]) ? node6235 : node6228;
													assign node6228 = (inp[0]) ? node6232 : node6229;
														assign node6229 = (inp[10]) ? 4'b0101 : 4'b1001;
														assign node6232 = (inp[7]) ? 4'b1100 : 4'b1000;
													assign node6235 = (inp[0]) ? 4'b0000 : 4'b1000;
											assign node6238 = (inp[10]) ? node6248 : node6239;
												assign node6239 = (inp[13]) ? node6243 : node6240;
													assign node6240 = (inp[0]) ? 4'b1100 : 4'b0101;
													assign node6243 = (inp[0]) ? 4'b0001 : node6244;
														assign node6244 = (inp[14]) ? 4'b0100 : 4'b0000;
												assign node6248 = (inp[0]) ? node6252 : node6249;
													assign node6249 = (inp[13]) ? 4'b0001 : 4'b0000;
													assign node6252 = (inp[7]) ? 4'b0001 : node6253;
														assign node6253 = (inp[13]) ? 4'b1001 : 4'b0001;
										assign node6257 = (inp[11]) ? node6287 : node6258;
											assign node6258 = (inp[10]) ? node6276 : node6259;
												assign node6259 = (inp[0]) ? node6269 : node6260;
													assign node6260 = (inp[7]) ? node6264 : node6261;
														assign node6261 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node6264 = (inp[14]) ? node6266 : 4'b0101;
															assign node6266 = (inp[13]) ? 4'b0000 : 4'b0100;
													assign node6269 = (inp[12]) ? 4'b1100 : node6270;
														assign node6270 = (inp[14]) ? 4'b1100 : node6271;
															assign node6271 = (inp[13]) ? 4'b1000 : 4'b0000;
												assign node6276 = (inp[0]) ? node6280 : node6277;
													assign node6277 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node6280 = (inp[14]) ? node6282 : 4'b0000;
														assign node6282 = (inp[13]) ? node6284 : 4'b0001;
															assign node6284 = (inp[12]) ? 4'b0001 : 4'b1001;
											assign node6287 = (inp[13]) ? 4'b1000 : node6288;
												assign node6288 = (inp[7]) ? node6294 : node6289;
													assign node6289 = (inp[0]) ? node6291 : 4'b1000;
														assign node6291 = (inp[14]) ? 4'b1000 : 4'b0000;
													assign node6294 = (inp[10]) ? node6298 : node6295;
														assign node6295 = (inp[12]) ? 4'b0100 : 4'b1100;
														assign node6298 = (inp[0]) ? 4'b0000 : 4'b1000;
							assign node6302 = (inp[4]) ? node6438 : node6303;
								assign node6303 = (inp[1]) ? node6383 : node6304;
									assign node6304 = (inp[10]) ? node6338 : node6305;
										assign node6305 = (inp[11]) ? node6323 : node6306;
											assign node6306 = (inp[2]) ? node6314 : node6307;
												assign node6307 = (inp[14]) ? node6311 : node6308;
													assign node6308 = (inp[12]) ? 4'b1000 : 4'b0000;
													assign node6311 = (inp[13]) ? 4'b1000 : 4'b1001;
												assign node6314 = (inp[7]) ? node6320 : node6315;
													assign node6315 = (inp[0]) ? 4'b1001 : node6316;
														assign node6316 = (inp[13]) ? 4'b0000 : 4'b0001;
													assign node6320 = (inp[14]) ? 4'b0000 : 4'b1000;
											assign node6323 = (inp[0]) ? 4'b1001 : node6324;
												assign node6324 = (inp[12]) ? node6330 : node6325;
													assign node6325 = (inp[2]) ? 4'b1000 : node6326;
														assign node6326 = (inp[13]) ? 4'b1001 : 4'b1000;
													assign node6330 = (inp[7]) ? node6334 : node6331;
														assign node6331 = (inp[13]) ? 4'b0001 : 4'b0000;
														assign node6334 = (inp[13]) ? 4'b1000 : 4'b0001;
										assign node6338 = (inp[2]) ? node6358 : node6339;
											assign node6339 = (inp[0]) ? node6349 : node6340;
												assign node6340 = (inp[12]) ? node6346 : node6341;
													assign node6341 = (inp[7]) ? 4'b0001 : node6342;
														assign node6342 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node6346 = (inp[11]) ? 4'b1001 : 4'b0000;
												assign node6349 = (inp[12]) ? node6355 : node6350;
													assign node6350 = (inp[11]) ? 4'b0000 : node6351;
														assign node6351 = (inp[7]) ? 4'b1000 : 4'b0000;
													assign node6355 = (inp[11]) ? 4'b0000 : 4'b0001;
											assign node6358 = (inp[14]) ? node6376 : node6359;
												assign node6359 = (inp[11]) ? node6369 : node6360;
													assign node6360 = (inp[0]) ? 4'b0001 : node6361;
														assign node6361 = (inp[13]) ? node6363 : 4'b1001;
															assign node6363 = (inp[7]) ? node6365 : 4'b1001;
																assign node6365 = (inp[12]) ? 4'b0000 : 4'b0001;
													assign node6369 = (inp[12]) ? node6371 : 4'b1000;
														assign node6371 = (inp[13]) ? 4'b0001 : node6372;
															assign node6372 = (inp[7]) ? 4'b1000 : 4'b0001;
												assign node6376 = (inp[13]) ? node6380 : node6377;
													assign node6377 = (inp[11]) ? 4'b0001 : 4'b1001;
													assign node6380 = (inp[12]) ? 4'b0001 : 4'b0000;
									assign node6383 = (inp[11]) ? node6425 : node6384;
										assign node6384 = (inp[2]) ? node6406 : node6385;
											assign node6385 = (inp[10]) ? node6399 : node6386;
												assign node6386 = (inp[14]) ? 4'b0000 : node6387;
													assign node6387 = (inp[12]) ? node6393 : node6388;
														assign node6388 = (inp[13]) ? node6390 : 4'b0000;
															assign node6390 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node6393 = (inp[0]) ? node6395 : 4'b0001;
															assign node6395 = (inp[13]) ? 4'b0000 : 4'b0001;
												assign node6399 = (inp[0]) ? node6401 : 4'b1001;
													assign node6401 = (inp[7]) ? node6403 : 4'b0000;
														assign node6403 = (inp[12]) ? 4'b0000 : 4'b1000;
											assign node6406 = (inp[10]) ? node6416 : node6407;
												assign node6407 = (inp[0]) ? 4'b1001 : node6408;
													assign node6408 = (inp[13]) ? 4'b0000 : node6409;
														assign node6409 = (inp[14]) ? 4'b0001 : node6410;
															assign node6410 = (inp[7]) ? 4'b1000 : 4'b1001;
												assign node6416 = (inp[13]) ? node6418 : 4'b0001;
													assign node6418 = (inp[0]) ? node6422 : node6419;
														assign node6419 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node6422 = (inp[14]) ? 4'b0000 : 4'b1001;
										assign node6425 = (inp[13]) ? node6431 : node6426;
											assign node6426 = (inp[14]) ? 4'b0000 : node6427;
												assign node6427 = (inp[0]) ? 4'b1000 : 4'b0000;
											assign node6431 = (inp[10]) ? 4'b1000 : node6432;
												assign node6432 = (inp[0]) ? 4'b0000 : node6433;
													assign node6433 = (inp[7]) ? 4'b1000 : 4'b0000;
								assign node6438 = (inp[13]) ? node6528 : node6439;
									assign node6439 = (inp[10]) ? node6493 : node6440;
										assign node6440 = (inp[14]) ? node6470 : node6441;
											assign node6441 = (inp[11]) ? node6455 : node6442;
												assign node6442 = (inp[1]) ? node6448 : node6443;
													assign node6443 = (inp[12]) ? 4'b1000 : node6444;
														assign node6444 = (inp[2]) ? 4'b1000 : 4'b0000;
													assign node6448 = (inp[0]) ? node6452 : node6449;
														assign node6449 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node6452 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node6455 = (inp[1]) ? node6463 : node6456;
													assign node6456 = (inp[12]) ? node6458 : 4'b1001;
														assign node6458 = (inp[0]) ? 4'b0001 : node6459;
															assign node6459 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node6463 = (inp[12]) ? 4'b1000 : node6464;
														assign node6464 = (inp[2]) ? node6466 : 4'b0000;
															assign node6466 = (inp[7]) ? 4'b0000 : 4'b1000;
											assign node6470 = (inp[7]) ? node6478 : node6471;
												assign node6471 = (inp[2]) ? node6473 : 4'b0000;
													assign node6473 = (inp[1]) ? 4'b0001 : node6474;
														assign node6474 = (inp[11]) ? 4'b0001 : 4'b0000;
												assign node6478 = (inp[12]) ? node6484 : node6479;
													assign node6479 = (inp[11]) ? node6481 : 4'b0001;
														assign node6481 = (inp[2]) ? 4'b0000 : 4'b1001;
													assign node6484 = (inp[0]) ? 4'b0000 : node6485;
														assign node6485 = (inp[11]) ? node6489 : node6486;
															assign node6486 = (inp[2]) ? 4'b1000 : 4'b1001;
															assign node6489 = (inp[1]) ? 4'b0000 : 4'b1000;
										assign node6493 = (inp[14]) ? node6517 : node6494;
											assign node6494 = (inp[11]) ? node6510 : node6495;
												assign node6495 = (inp[1]) ? node6501 : node6496;
													assign node6496 = (inp[0]) ? 4'b0001 : node6497;
														assign node6497 = (inp[12]) ? 4'b1000 : 4'b0001;
													assign node6501 = (inp[2]) ? node6507 : node6502;
														assign node6502 = (inp[12]) ? 4'b1000 : node6503;
															assign node6503 = (inp[0]) ? 4'b1000 : 4'b0000;
														assign node6507 = (inp[7]) ? 4'b0000 : 4'b0001;
												assign node6510 = (inp[2]) ? 4'b0000 : node6511;
													assign node6511 = (inp[1]) ? 4'b0000 : node6512;
														assign node6512 = (inp[0]) ? 4'b0000 : 4'b0001;
											assign node6517 = (inp[1]) ? 4'b0000 : node6518;
												assign node6518 = (inp[11]) ? node6520 : 4'b0000;
													assign node6520 = (inp[12]) ? 4'b0000 : node6521;
														assign node6521 = (inp[7]) ? 4'b1000 : node6522;
															assign node6522 = (inp[0]) ? 4'b0000 : 4'b1000;
									assign node6528 = (inp[1]) ? node6558 : node6529;
										assign node6529 = (inp[10]) ? node6547 : node6530;
											assign node6530 = (inp[0]) ? node6536 : node6531;
												assign node6531 = (inp[14]) ? node6533 : 4'b0000;
													assign node6533 = (inp[11]) ? 4'b0000 : 4'b0001;
												assign node6536 = (inp[2]) ? node6540 : node6537;
													assign node6537 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node6540 = (inp[12]) ? node6544 : node6541;
														assign node6541 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node6544 = (inp[7]) ? 4'b0000 : 4'b0001;
											assign node6547 = (inp[11]) ? 4'b0000 : node6548;
												assign node6548 = (inp[7]) ? node6554 : node6549;
													assign node6549 = (inp[14]) ? 4'b0000 : node6550;
														assign node6550 = (inp[2]) ? 4'b0000 : 4'b0001;
													assign node6554 = (inp[14]) ? 4'b0001 : 4'b0000;
										assign node6558 = (inp[14]) ? 4'b0000 : node6559;
											assign node6559 = (inp[7]) ? node6561 : 4'b0000;
												assign node6561 = (inp[2]) ? 4'b0000 : node6562;
													assign node6562 = (inp[11]) ? 4'b0000 : 4'b0001;
				assign node6567 = (inp[0]) ? node7543 : node6568;
					assign node6568 = (inp[6]) ? node6878 : node6569;
						assign node6569 = (inp[2]) ? node6803 : node6570;
							assign node6570 = (inp[5]) ? node6640 : node6571;
								assign node6571 = (inp[3]) ? node6573 : 4'b1010;
									assign node6573 = (inp[13]) ? node6607 : node6574;
										assign node6574 = (inp[4]) ? node6586 : node6575;
											assign node6575 = (inp[14]) ? 4'b1010 : node6576;
												assign node6576 = (inp[7]) ? 4'b1010 : node6577;
													assign node6577 = (inp[1]) ? 4'b0000 : node6578;
														assign node6578 = (inp[12]) ? 4'b1010 : node6579;
															assign node6579 = (inp[11]) ? 4'b0001 : 4'b1010;
											assign node6586 = (inp[7]) ? node6600 : node6587;
												assign node6587 = (inp[1]) ? node6589 : 4'b1001;
													assign node6589 = (inp[14]) ? node6595 : node6590;
														assign node6590 = (inp[12]) ? node6592 : 4'b0000;
															assign node6592 = (inp[10]) ? 4'b0000 : 4'b1000;
														assign node6595 = (inp[12]) ? 4'b0000 : node6596;
															assign node6596 = (inp[10]) ? 4'b0001 : 4'b1001;
												assign node6600 = (inp[12]) ? 4'b1010 : node6601;
													assign node6601 = (inp[14]) ? 4'b1010 : node6602;
														assign node6602 = (inp[10]) ? 4'b0001 : 4'b0000;
										assign node6607 = (inp[10]) ? node6623 : node6608;
											assign node6608 = (inp[1]) ? node6614 : node6609;
												assign node6609 = (inp[11]) ? 4'b0001 : node6610;
													assign node6610 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node6614 = (inp[12]) ? node6618 : node6615;
													assign node6615 = (inp[7]) ? 4'b1010 : 4'b1000;
													assign node6618 = (inp[11]) ? 4'b0000 : node6619;
														assign node6619 = (inp[14]) ? 4'b0001 : 4'b0000;
											assign node6623 = (inp[1]) ? node6633 : node6624;
												assign node6624 = (inp[12]) ? node6630 : node6625;
													assign node6625 = (inp[14]) ? node6627 : 4'b1001;
														assign node6627 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node6630 = (inp[11]) ? 4'b0001 : 4'b0000;
												assign node6633 = (inp[14]) ? node6635 : 4'b1000;
													assign node6635 = (inp[11]) ? 4'b1000 : node6636;
														assign node6636 = (inp[12]) ? 4'b0001 : 4'b1001;
								assign node6640 = (inp[1]) ? node6716 : node6641;
									assign node6641 = (inp[11]) ? node6683 : node6642;
										assign node6642 = (inp[14]) ? node6662 : node6643;
											assign node6643 = (inp[7]) ? node6653 : node6644;
												assign node6644 = (inp[3]) ? node6648 : node6645;
													assign node6645 = (inp[12]) ? 4'b0101 : 4'b1101;
													assign node6648 = (inp[12]) ? 4'b0001 : node6649;
														assign node6649 = (inp[13]) ? 4'b1001 : 4'b0001;
												assign node6653 = (inp[3]) ? node6655 : 4'b0001;
													assign node6655 = (inp[13]) ? 4'b0101 : node6656;
														assign node6656 = (inp[10]) ? node6658 : 4'b1101;
															assign node6658 = (inp[12]) ? 4'b1101 : 4'b0101;
											assign node6662 = (inp[13]) ? node6680 : node6663;
												assign node6663 = (inp[12]) ? node6667 : node6664;
													assign node6664 = (inp[10]) ? 4'b0100 : 4'b1100;
													assign node6667 = (inp[10]) ? node6675 : node6668;
														assign node6668 = (inp[3]) ? node6670 : 4'b1000;
															assign node6670 = (inp[7]) ? 4'b1100 : node6671;
																assign node6671 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node6675 = (inp[3]) ? node6677 : 4'b1100;
															assign node6677 = (inp[4]) ? 4'b1000 : 4'b1100;
												assign node6680 = (inp[12]) ? 4'b0100 : 4'b0000;
										assign node6683 = (inp[13]) ? node6701 : node6684;
											assign node6684 = (inp[12]) ? node6696 : node6685;
												assign node6685 = (inp[10]) ? node6691 : node6686;
													assign node6686 = (inp[14]) ? 4'b1101 : node6687;
														assign node6687 = (inp[4]) ? 4'b1001 : 4'b1101;
													assign node6691 = (inp[3]) ? 4'b0001 : node6692;
														assign node6692 = (inp[7]) ? 4'b0001 : 4'b0101;
												assign node6696 = (inp[3]) ? node6698 : 4'b1001;
													assign node6698 = (inp[7]) ? 4'b1101 : 4'b1001;
											assign node6701 = (inp[10]) ? node6709 : node6702;
												assign node6702 = (inp[7]) ? node6704 : 4'b0001;
													assign node6704 = (inp[3]) ? 4'b0101 : node6705;
														assign node6705 = (inp[4]) ? 4'b0101 : 4'b0001;
												assign node6709 = (inp[12]) ? node6713 : node6710;
													assign node6710 = (inp[3]) ? 4'b1001 : 4'b1101;
													assign node6713 = (inp[14]) ? 4'b0101 : 4'b0001;
									assign node6716 = (inp[14]) ? node6758 : node6717;
										assign node6717 = (inp[13]) ? node6733 : node6718;
											assign node6718 = (inp[10]) ? node6724 : node6719;
												assign node6719 = (inp[12]) ? 4'b1100 : node6720;
													assign node6720 = (inp[3]) ? 4'b0000 : 4'b0100;
												assign node6724 = (inp[4]) ? node6730 : node6725;
													assign node6725 = (inp[12]) ? node6727 : 4'b0100;
														assign node6727 = (inp[11]) ? 4'b0000 : 4'b0100;
													assign node6730 = (inp[3]) ? 4'b0000 : 4'b0100;
											assign node6733 = (inp[12]) ? node6741 : node6734;
												assign node6734 = (inp[10]) ? 4'b1100 : node6735;
													assign node6735 = (inp[3]) ? 4'b1000 : node6736;
														assign node6736 = (inp[4]) ? 4'b1100 : 4'b1000;
												assign node6741 = (inp[10]) ? node6749 : node6742;
													assign node6742 = (inp[3]) ? node6744 : 4'b0100;
														assign node6744 = (inp[7]) ? node6746 : 4'b0000;
															assign node6746 = (inp[4]) ? 4'b0000 : 4'b0100;
													assign node6749 = (inp[11]) ? node6751 : 4'b1000;
														assign node6751 = (inp[7]) ? node6753 : 4'b1100;
															assign node6753 = (inp[4]) ? node6755 : 4'b1000;
																assign node6755 = (inp[3]) ? 4'b1000 : 4'b1100;
										assign node6758 = (inp[11]) ? node6786 : node6759;
											assign node6759 = (inp[13]) ? node6777 : node6760;
												assign node6760 = (inp[12]) ? node6772 : node6761;
													assign node6761 = (inp[10]) ? node6763 : 4'b1001;
														assign node6763 = (inp[3]) ? node6767 : node6764;
															assign node6764 = (inp[4]) ? 4'b0101 : 4'b0001;
															assign node6767 = (inp[7]) ? node6769 : 4'b0001;
																assign node6769 = (inp[4]) ? 4'b0001 : 4'b0101;
													assign node6772 = (inp[3]) ? node6774 : 4'b1001;
														assign node6774 = (inp[7]) ? 4'b1101 : 4'b1001;
												assign node6777 = (inp[3]) ? node6783 : node6778;
													assign node6778 = (inp[7]) ? 4'b0001 : node6779;
														assign node6779 = (inp[10]) ? 4'b1101 : 4'b0101;
													assign node6783 = (inp[4]) ? 4'b0001 : 4'b1001;
											assign node6786 = (inp[13]) ? node6794 : node6787;
												assign node6787 = (inp[10]) ? 4'b0100 : node6788;
													assign node6788 = (inp[12]) ? node6790 : 4'b0100;
														assign node6790 = (inp[7]) ? 4'b1000 : 4'b1100;
												assign node6794 = (inp[10]) ? node6798 : node6795;
													assign node6795 = (inp[7]) ? 4'b0100 : 4'b0000;
													assign node6798 = (inp[12]) ? 4'b1100 : node6799;
														assign node6799 = (inp[3]) ? 4'b1000 : 4'b1100;
							assign node6803 = (inp[3]) ? node6805 : 4'b1010;
								assign node6805 = (inp[5]) ? node6807 : 4'b1010;
									assign node6807 = (inp[13]) ? node6847 : node6808;
										assign node6808 = (inp[7]) ? node6832 : node6809;
											assign node6809 = (inp[10]) ? node6819 : node6810;
												assign node6810 = (inp[4]) ? 4'b1000 : node6811;
													assign node6811 = (inp[14]) ? 4'b1010 : node6812;
														assign node6812 = (inp[1]) ? node6814 : 4'b1010;
															assign node6814 = (inp[12]) ? 4'b1010 : 4'b0000;
												assign node6819 = (inp[12]) ? node6825 : node6820;
													assign node6820 = (inp[1]) ? node6822 : 4'b0001;
														assign node6822 = (inp[14]) ? 4'b0001 : 4'b0000;
													assign node6825 = (inp[4]) ? node6827 : 4'b1010;
														assign node6827 = (inp[1]) ? node6829 : 4'b1001;
															assign node6829 = (inp[11]) ? 4'b0000 : 4'b1001;
											assign node6832 = (inp[4]) ? node6834 : 4'b1010;
												assign node6834 = (inp[1]) ? node6840 : node6835;
													assign node6835 = (inp[10]) ? node6837 : 4'b1010;
														assign node6837 = (inp[12]) ? 4'b1010 : 4'b0000;
													assign node6840 = (inp[12]) ? node6844 : node6841;
														assign node6841 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node6844 = (inp[10]) ? 4'b0000 : 4'b1010;
										assign node6847 = (inp[1]) ? node6861 : node6848;
											assign node6848 = (inp[10]) ? node6858 : node6849;
												assign node6849 = (inp[12]) ? node6855 : node6850;
													assign node6850 = (inp[11]) ? 4'b0001 : node6851;
														assign node6851 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node6855 = (inp[4]) ? 4'b0001 : 4'b1010;
												assign node6858 = (inp[12]) ? 4'b0001 : 4'b1001;
											assign node6861 = (inp[11]) ? node6873 : node6862;
												assign node6862 = (inp[14]) ? node6868 : node6863;
													assign node6863 = (inp[12]) ? node6865 : 4'b1000;
														assign node6865 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node6868 = (inp[4]) ? 4'b0001 : node6869;
														assign node6869 = (inp[7]) ? 4'b1010 : 4'b0001;
												assign node6873 = (inp[10]) ? 4'b1000 : node6874;
													assign node6874 = (inp[12]) ? 4'b0000 : 4'b1000;
						assign node6878 = (inp[5]) ? node7224 : node6879;
							assign node6879 = (inp[1]) ? node7067 : node6880;
								assign node6880 = (inp[13]) ? node6976 : node6881;
									assign node6881 = (inp[14]) ? node6917 : node6882;
										assign node6882 = (inp[3]) ? node6896 : node6883;
											assign node6883 = (inp[7]) ? 4'b1001 : node6884;
												assign node6884 = (inp[4]) ? node6890 : node6885;
													assign node6885 = (inp[10]) ? node6887 : 4'b1001;
														assign node6887 = (inp[11]) ? 4'b0101 : 4'b1001;
													assign node6890 = (inp[10]) ? node6892 : 4'b1101;
														assign node6892 = (inp[12]) ? 4'b1101 : 4'b0101;
											assign node6896 = (inp[11]) ? node6902 : node6897;
												assign node6897 = (inp[10]) ? node6899 : 4'b1101;
													assign node6899 = (inp[4]) ? 4'b1101 : 4'b0101;
												assign node6902 = (inp[7]) ? node6910 : node6903;
													assign node6903 = (inp[12]) ? node6907 : node6904;
														assign node6904 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node6907 = (inp[10]) ? 4'b0000 : 4'b1000;
													assign node6910 = (inp[2]) ? node6914 : node6911;
														assign node6911 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node6914 = (inp[10]) ? 4'b0101 : 4'b1101;
										assign node6917 = (inp[12]) ? node6945 : node6918;
											assign node6918 = (inp[3]) ? node6928 : node6919;
												assign node6919 = (inp[10]) ? node6923 : node6920;
													assign node6920 = (inp[11]) ? 4'b0000 : 4'b1000;
													assign node6923 = (inp[7]) ? node6925 : 4'b0100;
														assign node6925 = (inp[4]) ? 4'b0100 : 4'b0000;
												assign node6928 = (inp[11]) ? node6932 : node6929;
													assign node6929 = (inp[10]) ? 4'b0001 : 4'b1001;
													assign node6932 = (inp[2]) ? node6940 : node6933;
														assign node6933 = (inp[10]) ? node6935 : 4'b0000;
															assign node6935 = (inp[4]) ? node6937 : 4'b1000;
																assign node6937 = (inp[7]) ? 4'b1100 : 4'b1000;
														assign node6940 = (inp[7]) ? node6942 : 4'b0000;
															assign node6942 = (inp[4]) ? 4'b0001 : 4'b0101;
											assign node6945 = (inp[3]) ? node6955 : node6946;
												assign node6946 = (inp[11]) ? node6952 : node6947;
													assign node6947 = (inp[10]) ? 4'b1000 : node6948;
														assign node6948 = (inp[2]) ? 4'b1100 : 4'b1000;
													assign node6952 = (inp[7]) ? 4'b1001 : 4'b0000;
												assign node6955 = (inp[10]) ? node6967 : node6956;
													assign node6956 = (inp[2]) ? node6964 : node6957;
														assign node6957 = (inp[11]) ? node6961 : node6958;
															assign node6958 = (inp[4]) ? 4'b1101 : 4'b1001;
															assign node6961 = (inp[7]) ? 4'b1100 : 4'b1000;
														assign node6964 = (inp[11]) ? 4'b1101 : 4'b1100;
													assign node6967 = (inp[4]) ? 4'b0000 : node6968;
														assign node6968 = (inp[2]) ? 4'b1101 : node6969;
															assign node6969 = (inp[11]) ? 4'b0000 : node6970;
																assign node6970 = (inp[7]) ? 4'b0001 : 4'b0101;
									assign node6976 = (inp[2]) ? node7028 : node6977;
										assign node6977 = (inp[14]) ? node7009 : node6978;
											assign node6978 = (inp[4]) ? node6990 : node6979;
												assign node6979 = (inp[7]) ? node6983 : node6980;
													assign node6980 = (inp[11]) ? 4'b1100 : 4'b0101;
													assign node6983 = (inp[11]) ? 4'b0001 : node6984;
														assign node6984 = (inp[10]) ? 4'b1001 : node6985;
															assign node6985 = (inp[12]) ? 4'b1001 : 4'b0001;
												assign node6990 = (inp[10]) ? node6998 : node6991;
													assign node6991 = (inp[11]) ? 4'b0000 : node6992;
														assign node6992 = (inp[12]) ? 4'b0000 : node6993;
															assign node6993 = (inp[3]) ? 4'b1000 : 4'b1001;
													assign node6998 = (inp[7]) ? node7000 : 4'b0001;
														assign node7000 = (inp[3]) ? node7006 : node7001;
															assign node7001 = (inp[11]) ? node7003 : 4'b0001;
																assign node7003 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node7006 = (inp[11]) ? 4'b0001 : 4'b0000;
											assign node7009 = (inp[3]) ? node7015 : node7010;
												assign node7010 = (inp[7]) ? node7012 : 4'b1000;
													assign node7012 = (inp[4]) ? 4'b0101 : 4'b0000;
												assign node7015 = (inp[4]) ? node7019 : node7016;
													assign node7016 = (inp[11]) ? 4'b1100 : 4'b0101;
													assign node7019 = (inp[11]) ? node7023 : node7020;
														assign node7020 = (inp[10]) ? 4'b1001 : 4'b1101;
														assign node7023 = (inp[12]) ? node7025 : 4'b0001;
															assign node7025 = (inp[7]) ? 4'b1100 : 4'b0001;
										assign node7028 = (inp[3]) ? node7046 : node7029;
											assign node7029 = (inp[11]) ? node7041 : node7030;
												assign node7030 = (inp[14]) ? node7036 : node7031;
													assign node7031 = (inp[10]) ? node7033 : 4'b0001;
														assign node7033 = (inp[12]) ? 4'b0101 : 4'b1101;
													assign node7036 = (inp[10]) ? 4'b1100 : node7037;
														assign node7037 = (inp[7]) ? 4'b0000 : 4'b0100;
												assign node7041 = (inp[12]) ? 4'b0101 : node7042;
													assign node7042 = (inp[14]) ? 4'b1101 : 4'b0101;
											assign node7046 = (inp[4]) ? node7056 : node7047;
												assign node7047 = (inp[10]) ? node7051 : node7048;
													assign node7048 = (inp[7]) ? 4'b0101 : 4'b0001;
													assign node7051 = (inp[12]) ? 4'b0100 : node7052;
														assign node7052 = (inp[11]) ? 4'b1101 : 4'b1100;
												assign node7056 = (inp[11]) ? node7060 : node7057;
													assign node7057 = (inp[10]) ? 4'b0001 : 4'b0000;
													assign node7060 = (inp[12]) ? node7062 : 4'b1000;
														assign node7062 = (inp[7]) ? 4'b0001 : node7063;
															assign node7063 = (inp[10]) ? 4'b0000 : 4'b1000;
								assign node7067 = (inp[11]) ? node7163 : node7068;
									assign node7068 = (inp[14]) ? node7118 : node7069;
										assign node7069 = (inp[2]) ? node7091 : node7070;
											assign node7070 = (inp[4]) ? node7078 : node7071;
												assign node7071 = (inp[7]) ? 4'b1000 : node7072;
													assign node7072 = (inp[3]) ? node7074 : 4'b0100;
														assign node7074 = (inp[12]) ? 4'b0101 : 4'b1101;
												assign node7078 = (inp[13]) ? node7084 : node7079;
													assign node7079 = (inp[7]) ? node7081 : 4'b0001;
														assign node7081 = (inp[3]) ? 4'b0101 : 4'b0100;
													assign node7084 = (inp[3]) ? node7086 : 4'b0001;
														assign node7086 = (inp[12]) ? 4'b0001 : node7087;
															assign node7087 = (inp[7]) ? 4'b0001 : 4'b1001;
											assign node7091 = (inp[3]) ? node7103 : node7092;
												assign node7092 = (inp[13]) ? node7098 : node7093;
													assign node7093 = (inp[4]) ? 4'b0100 : node7094;
														assign node7094 = (inp[12]) ? 4'b1000 : 4'b0000;
													assign node7098 = (inp[4]) ? 4'b1100 : node7099;
														assign node7099 = (inp[12]) ? 4'b0100 : 4'b1100;
												assign node7103 = (inp[7]) ? node7113 : node7104;
													assign node7104 = (inp[4]) ? node7108 : node7105;
														assign node7105 = (inp[13]) ? 4'b1000 : 4'b0000;
														assign node7108 = (inp[10]) ? node7110 : 4'b1000;
															assign node7110 = (inp[13]) ? 4'b0001 : 4'b1001;
													assign node7113 = (inp[12]) ? 4'b1100 : node7114;
														assign node7114 = (inp[10]) ? 4'b0100 : 4'b0001;
										assign node7118 = (inp[7]) ? node7140 : node7119;
											assign node7119 = (inp[4]) ? node7131 : node7120;
												assign node7120 = (inp[12]) ? 4'b1101 : node7121;
													assign node7121 = (inp[10]) ? node7123 : 4'b0101;
														assign node7123 = (inp[2]) ? node7125 : 4'b1101;
															assign node7125 = (inp[13]) ? node7127 : 4'b0001;
																assign node7127 = (inp[3]) ? 4'b1001 : 4'b1101;
												assign node7131 = (inp[10]) ? node7137 : node7132;
													assign node7132 = (inp[13]) ? node7134 : 4'b1101;
														assign node7134 = (inp[2]) ? 4'b1001 : 4'b1000;
													assign node7137 = (inp[12]) ? 4'b0001 : 4'b1001;
											assign node7140 = (inp[13]) ? node7148 : node7141;
												assign node7141 = (inp[12]) ? node7143 : 4'b0101;
													assign node7143 = (inp[10]) ? node7145 : 4'b1001;
														assign node7145 = (inp[4]) ? 4'b0101 : 4'b1101;
												assign node7148 = (inp[10]) ? node7158 : node7149;
													assign node7149 = (inp[4]) ? node7151 : 4'b0001;
														assign node7151 = (inp[12]) ? node7155 : node7152;
															assign node7152 = (inp[3]) ? 4'b0001 : 4'b0101;
															assign node7155 = (inp[3]) ? 4'b1101 : 4'b0101;
													assign node7158 = (inp[4]) ? node7160 : 4'b1001;
														assign node7160 = (inp[12]) ? 4'b0000 : 4'b1000;
									assign node7163 = (inp[4]) ? node7191 : node7164;
										assign node7164 = (inp[7]) ? node7182 : node7165;
											assign node7165 = (inp[12]) ? node7177 : node7166;
												assign node7166 = (inp[13]) ? node7172 : node7167;
													assign node7167 = (inp[3]) ? node7169 : 4'b0100;
														assign node7169 = (inp[2]) ? 4'b0000 : 4'b1100;
													assign node7172 = (inp[3]) ? node7174 : 4'b1100;
														assign node7174 = (inp[14]) ? 4'b1100 : 4'b0100;
												assign node7177 = (inp[2]) ? node7179 : 4'b0100;
													assign node7179 = (inp[3]) ? 4'b0000 : 4'b0100;
											assign node7182 = (inp[10]) ? node7186 : node7183;
												assign node7183 = (inp[14]) ? 4'b0100 : 4'b1000;
												assign node7186 = (inp[2]) ? node7188 : 4'b1000;
													assign node7188 = (inp[13]) ? 4'b1000 : 4'b0000;
										assign node7191 = (inp[7]) ? node7201 : node7192;
											assign node7192 = (inp[12]) ? node7198 : node7193;
												assign node7193 = (inp[2]) ? node7195 : 4'b0000;
													assign node7195 = (inp[13]) ? 4'b0000 : 4'b0100;
												assign node7198 = (inp[3]) ? 4'b0000 : 4'b1000;
											assign node7201 = (inp[3]) ? node7213 : node7202;
												assign node7202 = (inp[2]) ? node7206 : node7203;
													assign node7203 = (inp[13]) ? 4'b0000 : 4'b0100;
													assign node7206 = (inp[14]) ? 4'b1100 : node7207;
														assign node7207 = (inp[13]) ? 4'b0100 : node7208;
															assign node7208 = (inp[12]) ? 4'b1000 : 4'b0100;
												assign node7213 = (inp[13]) ? node7221 : node7214;
													assign node7214 = (inp[12]) ? node7218 : node7215;
														assign node7215 = (inp[2]) ? 4'b0000 : 4'b1100;
														assign node7218 = (inp[2]) ? 4'b1100 : 4'b0100;
													assign node7221 = (inp[10]) ? 4'b1000 : 4'b0000;
							assign node7224 = (inp[3]) ? node7396 : node7225;
								assign node7225 = (inp[11]) ? node7303 : node7226;
									assign node7226 = (inp[4]) ? node7262 : node7227;
										assign node7227 = (inp[10]) ? node7241 : node7228;
											assign node7228 = (inp[13]) ? node7232 : node7229;
												assign node7229 = (inp[1]) ? 4'b0001 : 4'b1001;
												assign node7232 = (inp[12]) ? node7234 : 4'b0101;
													assign node7234 = (inp[7]) ? node7238 : node7235;
														assign node7235 = (inp[2]) ? 4'b1101 : 4'b0101;
														assign node7238 = (inp[14]) ? 4'b1100 : 4'b1101;
											assign node7241 = (inp[13]) ? node7249 : node7242;
												assign node7242 = (inp[7]) ? node7244 : 4'b1101;
													assign node7244 = (inp[2]) ? node7246 : 4'b1001;
														assign node7246 = (inp[1]) ? 4'b1001 : 4'b0001;
												assign node7249 = (inp[2]) ? node7255 : node7250;
													assign node7250 = (inp[12]) ? 4'b1000 : node7251;
														assign node7251 = (inp[1]) ? 4'b1000 : 4'b0000;
													assign node7255 = (inp[14]) ? node7259 : node7256;
														assign node7256 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node7259 = (inp[12]) ? 4'b0000 : 4'b0001;
										assign node7262 = (inp[10]) ? node7288 : node7263;
											assign node7263 = (inp[2]) ? node7279 : node7264;
												assign node7264 = (inp[7]) ? node7272 : node7265;
													assign node7265 = (inp[13]) ? node7269 : node7266;
														assign node7266 = (inp[12]) ? 4'b1000 : 4'b1100;
														assign node7269 = (inp[14]) ? 4'b0101 : 4'b0100;
													assign node7272 = (inp[14]) ? node7276 : node7273;
														assign node7273 = (inp[1]) ? 4'b0000 : 4'b1000;
														assign node7276 = (inp[12]) ? 4'b1001 : 4'b1000;
												assign node7279 = (inp[12]) ? 4'b0000 : node7280;
													assign node7280 = (inp[14]) ? node7282 : 4'b0001;
														assign node7282 = (inp[1]) ? node7284 : 4'b0001;
															assign node7284 = (inp[13]) ? 4'b1000 : 4'b0000;
											assign node7288 = (inp[2]) ? node7298 : node7289;
												assign node7289 = (inp[1]) ? 4'b0001 : node7290;
													assign node7290 = (inp[7]) ? node7294 : node7291;
														assign node7291 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node7294 = (inp[13]) ? 4'b1001 : 4'b1000;
												assign node7298 = (inp[7]) ? node7300 : 4'b1000;
													assign node7300 = (inp[13]) ? 4'b0000 : 4'b1000;
									assign node7303 = (inp[1]) ? node7349 : node7304;
										assign node7304 = (inp[2]) ? node7322 : node7305;
											assign node7305 = (inp[13]) ? node7315 : node7306;
												assign node7306 = (inp[4]) ? node7312 : node7307;
													assign node7307 = (inp[12]) ? 4'b1001 : node7308;
														assign node7308 = (inp[10]) ? 4'b1101 : 4'b0001;
													assign node7312 = (inp[12]) ? 4'b0001 : 4'b0100;
												assign node7315 = (inp[7]) ? node7317 : 4'b0000;
													assign node7317 = (inp[14]) ? node7319 : 4'b0000;
														assign node7319 = (inp[4]) ? 4'b1001 : 4'b1101;
											assign node7322 = (inp[7]) ? node7332 : node7323;
												assign node7323 = (inp[4]) ? node7327 : node7324;
													assign node7324 = (inp[13]) ? 4'b0001 : 4'b0100;
													assign node7327 = (inp[13]) ? 4'b0000 : node7328;
														assign node7328 = (inp[12]) ? 4'b1001 : 4'b0001;
												assign node7332 = (inp[13]) ? node7342 : node7333;
													assign node7333 = (inp[4]) ? node7339 : node7334;
														assign node7334 = (inp[14]) ? 4'b0000 : node7335;
															assign node7335 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node7339 = (inp[12]) ? 4'b1100 : 4'b1001;
													assign node7342 = (inp[4]) ? 4'b0000 : node7343;
														assign node7343 = (inp[12]) ? 4'b1000 : node7344;
															assign node7344 = (inp[10]) ? 4'b1100 : 4'b0100;
										assign node7349 = (inp[13]) ? node7381 : node7350;
											assign node7350 = (inp[7]) ? node7366 : node7351;
												assign node7351 = (inp[4]) ? node7357 : node7352;
													assign node7352 = (inp[2]) ? 4'b0100 : node7353;
														assign node7353 = (inp[10]) ? 4'b0100 : 4'b1100;
													assign node7357 = (inp[14]) ? 4'b1000 : node7358;
														assign node7358 = (inp[10]) ? 4'b0100 : node7359;
															assign node7359 = (inp[12]) ? node7361 : 4'b0000;
																assign node7361 = (inp[2]) ? 4'b0000 : 4'b1100;
												assign node7366 = (inp[12]) ? node7372 : node7367;
													assign node7367 = (inp[4]) ? node7369 : 4'b1000;
														assign node7369 = (inp[10]) ? 4'b0000 : 4'b1000;
													assign node7372 = (inp[14]) ? 4'b0000 : node7373;
														assign node7373 = (inp[2]) ? node7377 : node7374;
															assign node7374 = (inp[10]) ? 4'b0000 : 4'b1000;
															assign node7377 = (inp[10]) ? 4'b1000 : 4'b0000;
											assign node7381 = (inp[10]) ? 4'b1000 : node7382;
												assign node7382 = (inp[7]) ? node7386 : node7383;
													assign node7383 = (inp[4]) ? 4'b0000 : 4'b1000;
													assign node7386 = (inp[14]) ? node7392 : node7387;
														assign node7387 = (inp[12]) ? 4'b1000 : node7388;
															assign node7388 = (inp[2]) ? 4'b0100 : 4'b1000;
														assign node7392 = (inp[4]) ? 4'b0100 : 4'b1100;
								assign node7396 = (inp[4]) ? node7484 : node7397;
									assign node7397 = (inp[1]) ? node7459 : node7398;
										assign node7398 = (inp[11]) ? node7428 : node7399;
											assign node7399 = (inp[10]) ? node7413 : node7400;
												assign node7400 = (inp[13]) ? node7404 : node7401;
													assign node7401 = (inp[12]) ? 4'b1000 : 4'b0000;
													assign node7404 = (inp[7]) ? node7410 : node7405;
														assign node7405 = (inp[12]) ? 4'b1001 : node7406;
															assign node7406 = (inp[2]) ? 4'b0001 : 4'b1000;
														assign node7410 = (inp[12]) ? 4'b0000 : 4'b0001;
												assign node7413 = (inp[7]) ? node7419 : node7414;
													assign node7414 = (inp[13]) ? node7416 : 4'b0000;
														assign node7416 = (inp[2]) ? 4'b0000 : 4'b0001;
													assign node7419 = (inp[2]) ? node7421 : 4'b1001;
														assign node7421 = (inp[14]) ? node7425 : node7422;
															assign node7422 = (inp[13]) ? 4'b0000 : 4'b0001;
															assign node7425 = (inp[12]) ? 4'b0001 : 4'b0000;
											assign node7428 = (inp[12]) ? node7444 : node7429;
												assign node7429 = (inp[13]) ? node7437 : node7430;
													assign node7430 = (inp[2]) ? node7432 : 4'b1000;
														assign node7432 = (inp[10]) ? 4'b1001 : node7433;
															assign node7433 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node7437 = (inp[2]) ? node7441 : node7438;
														assign node7438 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node7441 = (inp[7]) ? 4'b1000 : 4'b0001;
												assign node7444 = (inp[10]) ? node7452 : node7445;
													assign node7445 = (inp[2]) ? node7447 : 4'b0001;
														assign node7447 = (inp[13]) ? 4'b0000 : node7448;
															assign node7448 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node7452 = (inp[2]) ? node7456 : node7453;
														assign node7453 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node7456 = (inp[7]) ? 4'b1001 : 4'b0001;
										assign node7459 = (inp[11]) ? node7475 : node7460;
											assign node7460 = (inp[10]) ? node7468 : node7461;
												assign node7461 = (inp[12]) ? node7463 : 4'b1000;
													assign node7463 = (inp[2]) ? 4'b0001 : node7464;
														assign node7464 = (inp[13]) ? 4'b1000 : 4'b1001;
												assign node7468 = (inp[14]) ? node7472 : node7469;
													assign node7469 = (inp[12]) ? 4'b1000 : 4'b0000;
													assign node7472 = (inp[2]) ? 4'b0001 : 4'b0000;
											assign node7475 = (inp[10]) ? node7479 : node7476;
												assign node7476 = (inp[13]) ? 4'b0000 : 4'b1000;
												assign node7479 = (inp[7]) ? 4'b1000 : node7480;
													assign node7480 = (inp[14]) ? 4'b1000 : 4'b0000;
									assign node7484 = (inp[1]) ? node7530 : node7485;
										assign node7485 = (inp[13]) ? node7505 : node7486;
											assign node7486 = (inp[10]) ? node7494 : node7487;
												assign node7487 = (inp[12]) ? node7491 : node7488;
													assign node7488 = (inp[2]) ? 4'b0001 : 4'b1001;
													assign node7491 = (inp[2]) ? 4'b1000 : 4'b0000;
												assign node7494 = (inp[7]) ? node7496 : 4'b0001;
													assign node7496 = (inp[12]) ? node7498 : 4'b0000;
														assign node7498 = (inp[11]) ? node7502 : node7499;
															assign node7499 = (inp[2]) ? 4'b0000 : 4'b0001;
															assign node7502 = (inp[2]) ? 4'b0001 : 4'b0000;
											assign node7505 = (inp[12]) ? node7515 : node7506;
												assign node7506 = (inp[11]) ? 4'b0000 : node7507;
													assign node7507 = (inp[14]) ? 4'b0000 : node7508;
														assign node7508 = (inp[10]) ? 4'b0000 : node7509;
															assign node7509 = (inp[2]) ? 4'b0000 : 4'b0001;
												assign node7515 = (inp[7]) ? node7519 : node7516;
													assign node7516 = (inp[2]) ? 4'b0001 : 4'b0000;
													assign node7519 = (inp[11]) ? 4'b0000 : node7520;
														assign node7520 = (inp[14]) ? node7522 : 4'b0000;
															assign node7522 = (inp[2]) ? node7526 : node7523;
																assign node7523 = (inp[10]) ? 4'b0001 : 4'b0000;
																assign node7526 = (inp[10]) ? 4'b0000 : 4'b0001;
										assign node7530 = (inp[11]) ? 4'b0000 : node7531;
											assign node7531 = (inp[2]) ? node7539 : node7532;
												assign node7532 = (inp[13]) ? 4'b0000 : node7533;
													assign node7533 = (inp[10]) ? node7535 : 4'b1000;
														assign node7535 = (inp[14]) ? 4'b0001 : 4'b0000;
												assign node7539 = (inp[10]) ? 4'b0000 : 4'b0001;
					assign node7543 = (inp[6]) ? node7545 : 4'b1000;
						assign node7545 = (inp[5]) ? node7609 : node7546;
							assign node7546 = (inp[3]) ? node7548 : 4'b1000;
								assign node7548 = (inp[2]) ? 4'b1000 : node7549;
									assign node7549 = (inp[1]) ? node7577 : node7550;
										assign node7550 = (inp[7]) ? node7568 : node7551;
											assign node7551 = (inp[11]) ? node7563 : node7552;
												assign node7552 = (inp[14]) ? node7558 : node7553;
													assign node7553 = (inp[13]) ? 4'b0001 : node7554;
														assign node7554 = (inp[10]) ? 4'b0001 : 4'b1000;
													assign node7558 = (inp[12]) ? node7560 : 4'b0000;
														assign node7560 = (inp[13]) ? 4'b0000 : 4'b1000;
												assign node7563 = (inp[12]) ? 4'b1001 : node7564;
													assign node7564 = (inp[10]) ? 4'b1001 : 4'b0001;
											assign node7568 = (inp[4]) ? node7570 : 4'b1000;
												assign node7570 = (inp[11]) ? 4'b0001 : node7571;
													assign node7571 = (inp[14]) ? node7573 : 4'b1001;
														assign node7573 = (inp[13]) ? 4'b0000 : 4'b1000;
										assign node7577 = (inp[14]) ? node7595 : node7578;
											assign node7578 = (inp[11]) ? node7588 : node7579;
												assign node7579 = (inp[12]) ? node7581 : 4'b1000;
													assign node7581 = (inp[7]) ? node7585 : node7582;
														assign node7582 = (inp[4]) ? 4'b1000 : 4'b0000;
														assign node7585 = (inp[10]) ? 4'b0000 : 4'b1000;
												assign node7588 = (inp[7]) ? node7590 : 4'b0000;
													assign node7590 = (inp[13]) ? node7592 : 4'b1000;
														assign node7592 = (inp[10]) ? 4'b1000 : 4'b0000;
											assign node7595 = (inp[11]) ? node7605 : node7596;
												assign node7596 = (inp[4]) ? node7602 : node7597;
													assign node7597 = (inp[12]) ? 4'b1000 : node7598;
														assign node7598 = (inp[13]) ? 4'b1001 : 4'b1000;
													assign node7602 = (inp[7]) ? 4'b0001 : 4'b1001;
												assign node7605 = (inp[13]) ? 4'b1000 : 4'b0000;
							assign node7609 = (inp[2]) ? node7771 : node7610;
								assign node7610 = (inp[3]) ? node7692 : node7611;
									assign node7611 = (inp[7]) ? node7649 : node7612;
										assign node7612 = (inp[4]) ? node7630 : node7613;
											assign node7613 = (inp[1]) ? node7619 : node7614;
												assign node7614 = (inp[13]) ? node7616 : 4'b1001;
													assign node7616 = (inp[12]) ? 4'b0101 : 4'b1101;
												assign node7619 = (inp[14]) ? node7623 : node7620;
													assign node7620 = (inp[13]) ? 4'b1100 : 4'b0100;
													assign node7623 = (inp[11]) ? 4'b0100 : node7624;
														assign node7624 = (inp[13]) ? 4'b0101 : node7625;
															assign node7625 = (inp[10]) ? 4'b0101 : 4'b1001;
											assign node7630 = (inp[11]) ? node7640 : node7631;
												assign node7631 = (inp[12]) ? node7637 : node7632;
													assign node7632 = (inp[10]) ? node7634 : 4'b0001;
														assign node7634 = (inp[1]) ? 4'b1001 : 4'b0001;
													assign node7637 = (inp[10]) ? 4'b0001 : 4'b1100;
												assign node7640 = (inp[1]) ? 4'b1000 : node7641;
													assign node7641 = (inp[14]) ? node7643 : 4'b0000;
														assign node7643 = (inp[12]) ? 4'b0000 : node7644;
															assign node7644 = (inp[13]) ? 4'b0000 : 4'b1000;
										assign node7649 = (inp[12]) ? node7671 : node7650;
											assign node7650 = (inp[10]) ? node7660 : node7651;
												assign node7651 = (inp[11]) ? 4'b0000 : node7652;
													assign node7652 = (inp[13]) ? node7656 : node7653;
														assign node7653 = (inp[4]) ? 4'b1001 : 4'b1000;
														assign node7656 = (inp[14]) ? 4'b0100 : 4'b1000;
												assign node7660 = (inp[13]) ? node7666 : node7661;
													assign node7661 = (inp[4]) ? 4'b0101 : node7662;
														assign node7662 = (inp[1]) ? 4'b0000 : 4'b0001;
													assign node7666 = (inp[4]) ? node7668 : 4'b1001;
														assign node7668 = (inp[1]) ? 4'b1001 : 4'b1000;
											assign node7671 = (inp[13]) ? node7681 : node7672;
												assign node7672 = (inp[1]) ? node7678 : node7673;
													assign node7673 = (inp[11]) ? 4'b1001 : node7674;
														assign node7674 = (inp[14]) ? 4'b1000 : 4'b1001;
													assign node7678 = (inp[10]) ? 4'b0000 : 4'b1000;
												assign node7681 = (inp[4]) ? node7687 : node7682;
													assign node7682 = (inp[1]) ? 4'b0001 : node7683;
														assign node7683 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node7687 = (inp[1]) ? 4'b1000 : node7688;
														assign node7688 = (inp[11]) ? 4'b0000 : 4'b0001;
									assign node7692 = (inp[1]) ? node7734 : node7693;
										assign node7693 = (inp[13]) ? node7713 : node7694;
											assign node7694 = (inp[4]) ? node7702 : node7695;
												assign node7695 = (inp[10]) ? 4'b1001 : node7696;
													assign node7696 = (inp[12]) ? 4'b1001 : node7697;
														assign node7697 = (inp[11]) ? 4'b0001 : 4'b0000;
												assign node7702 = (inp[10]) ? node7710 : node7703;
													assign node7703 = (inp[7]) ? 4'b1000 : node7704;
														assign node7704 = (inp[11]) ? 4'b1000 : node7705;
															assign node7705 = (inp[12]) ? 4'b1001 : 4'b0001;
													assign node7710 = (inp[11]) ? 4'b0001 : 4'b0000;
											assign node7713 = (inp[7]) ? node7721 : node7714;
												assign node7714 = (inp[11]) ? node7716 : 4'b0000;
													assign node7716 = (inp[12]) ? 4'b0000 : node7717;
														assign node7717 = (inp[4]) ? 4'b0000 : 4'b0001;
												assign node7721 = (inp[4]) ? node7731 : node7722;
													assign node7722 = (inp[12]) ? node7728 : node7723;
														assign node7723 = (inp[10]) ? 4'b0000 : node7724;
															assign node7724 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node7728 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node7731 = (inp[14]) ? 4'b0000 : 4'b0001;
										assign node7734 = (inp[4]) ? node7756 : node7735;
											assign node7735 = (inp[13]) ? node7747 : node7736;
												assign node7736 = (inp[11]) ? node7742 : node7737;
													assign node7737 = (inp[7]) ? 4'b0001 : node7738;
														assign node7738 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node7742 = (inp[7]) ? 4'b0000 : node7743;
														assign node7743 = (inp[10]) ? 4'b0000 : 4'b1000;
												assign node7747 = (inp[7]) ? node7751 : node7748;
													assign node7748 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node7751 = (inp[14]) ? 4'b1000 : node7752;
														assign node7752 = (inp[10]) ? 4'b1000 : 4'b1001;
											assign node7756 = (inp[13]) ? 4'b0000 : node7757;
												assign node7757 = (inp[12]) ? 4'b0000 : node7758;
													assign node7758 = (inp[11]) ? 4'b1000 : node7759;
														assign node7759 = (inp[7]) ? node7765 : node7760;
															assign node7760 = (inp[14]) ? node7762 : 4'b0001;
																assign node7762 = (inp[10]) ? 4'b0001 : 4'b0000;
															assign node7765 = (inp[10]) ? 4'b0000 : 4'b1000;
								assign node7771 = (inp[3]) ? node7773 : 4'b1000;
									assign node7773 = (inp[7]) ? node7817 : node7774;
										assign node7774 = (inp[1]) ? node7796 : node7775;
											assign node7775 = (inp[11]) ? node7785 : node7776;
												assign node7776 = (inp[4]) ? node7782 : node7777;
													assign node7777 = (inp[14]) ? node7779 : 4'b1001;
														assign node7779 = (inp[13]) ? 4'b0000 : 4'b1000;
													assign node7782 = (inp[13]) ? 4'b0000 : 4'b0001;
												assign node7785 = (inp[4]) ? 4'b1001 : node7786;
													assign node7786 = (inp[14]) ? node7792 : node7787;
														assign node7787 = (inp[13]) ? node7789 : 4'b0001;
															assign node7789 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node7792 = (inp[13]) ? 4'b0001 : 4'b1000;
											assign node7796 = (inp[11]) ? node7812 : node7797;
												assign node7797 = (inp[14]) ? node7807 : node7798;
													assign node7798 = (inp[12]) ? node7804 : node7799;
														assign node7799 = (inp[10]) ? 4'b1000 : node7800;
															assign node7800 = (inp[4]) ? 4'b0001 : 4'b0000;
														assign node7804 = (inp[13]) ? 4'b0000 : 4'b1000;
													assign node7807 = (inp[13]) ? node7809 : 4'b1001;
														assign node7809 = (inp[10]) ? 4'b0001 : 4'b0000;
												assign node7812 = (inp[4]) ? 4'b0000 : node7813;
													assign node7813 = (inp[13]) ? 4'b1000 : 4'b0000;
										assign node7817 = (inp[4]) ? node7819 : 4'b1000;
											assign node7819 = (inp[13]) ? node7827 : node7820;
												assign node7820 = (inp[10]) ? node7822 : 4'b1000;
													assign node7822 = (inp[12]) ? 4'b1000 : node7823;
														assign node7823 = (inp[1]) ? 4'b0000 : 4'b0001;
												assign node7827 = (inp[10]) ? 4'b0000 : node7828;
													assign node7828 = (inp[14]) ? 4'b0001 : 4'b0000;
			assign node7832 = (inp[15]) ? node9234 : node7833;
				assign node7833 = (inp[6]) ? node8207 : node7834;
					assign node7834 = (inp[0]) ? 4'b0100 : node7835;
						assign node7835 = (inp[5]) ? node7949 : node7836;
							assign node7836 = (inp[2]) ? 4'b0110 : node7837;
								assign node7837 = (inp[3]) ? node7877 : node7838;
									assign node7838 = (inp[7]) ? node7866 : node7839;
										assign node7839 = (inp[4]) ? node7845 : node7840;
											assign node7840 = (inp[13]) ? node7842 : 4'b0110;
												assign node7842 = (inp[10]) ? 4'b0000 : 4'b0110;
											assign node7845 = (inp[1]) ? node7857 : node7846;
												assign node7846 = (inp[11]) ? node7852 : node7847;
													assign node7847 = (inp[14]) ? node7849 : 4'b1001;
														assign node7849 = (inp[13]) ? 4'b1000 : 4'b0000;
													assign node7852 = (inp[13]) ? 4'b1001 : node7853;
														assign node7853 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node7857 = (inp[14]) ? node7863 : node7858;
													assign node7858 = (inp[10]) ? node7860 : 4'b0000;
														assign node7860 = (inp[13]) ? 4'b0000 : 4'b1000;
													assign node7863 = (inp[11]) ? 4'b0000 : 4'b0001;
										assign node7866 = (inp[13]) ? node7868 : 4'b0110;
											assign node7868 = (inp[4]) ? node7870 : 4'b0110;
												assign node7870 = (inp[1]) ? node7872 : 4'b0110;
													assign node7872 = (inp[11]) ? 4'b0000 : node7873;
														assign node7873 = (inp[14]) ? 4'b0001 : 4'b0000;
									assign node7877 = (inp[1]) ? node7907 : node7878;
										assign node7878 = (inp[10]) ? node7886 : node7879;
											assign node7879 = (inp[13]) ? node7883 : node7880;
												assign node7880 = (inp[11]) ? 4'b0001 : 4'b0000;
												assign node7883 = (inp[14]) ? 4'b1000 : 4'b1001;
											assign node7886 = (inp[7]) ? node7892 : node7887;
												assign node7887 = (inp[4]) ? 4'b0101 : node7888;
													assign node7888 = (inp[12]) ? 4'b0001 : 4'b0101;
												assign node7892 = (inp[14]) ? node7900 : node7893;
													assign node7893 = (inp[13]) ? node7897 : node7894;
														assign node7894 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node7897 = (inp[11]) ? 4'b0101 : 4'b0001;
													assign node7900 = (inp[11]) ? node7902 : 4'b0000;
														assign node7902 = (inp[12]) ? 4'b1001 : node7903;
															assign node7903 = (inp[13]) ? 4'b0001 : 4'b1001;
										assign node7907 = (inp[4]) ? node7925 : node7908;
											assign node7908 = (inp[10]) ? node7914 : node7909;
												assign node7909 = (inp[13]) ? 4'b1000 : node7910;
													assign node7910 = (inp[7]) ? 4'b0000 : 4'b1000;
												assign node7914 = (inp[7]) ? node7916 : 4'b0100;
													assign node7916 = (inp[11]) ? node7922 : node7917;
														assign node7917 = (inp[13]) ? node7919 : 4'b0001;
															assign node7919 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node7922 = (inp[13]) ? 4'b0000 : 4'b1000;
											assign node7925 = (inp[11]) ? node7937 : node7926;
												assign node7926 = (inp[14]) ? node7928 : 4'b0100;
													assign node7928 = (inp[7]) ? 4'b0101 : node7929;
														assign node7929 = (inp[10]) ? node7933 : node7930;
															assign node7930 = (inp[13]) ? 4'b1101 : 4'b0101;
															assign node7933 = (inp[13]) ? 4'b0101 : 4'b1101;
												assign node7937 = (inp[7]) ? node7943 : node7938;
													assign node7938 = (inp[10]) ? 4'b1100 : node7939;
														assign node7939 = (inp[13]) ? 4'b1100 : 4'b0100;
													assign node7943 = (inp[13]) ? 4'b0100 : node7944;
														assign node7944 = (inp[10]) ? 4'b1000 : 4'b0000;
							assign node7949 = (inp[1]) ? node8087 : node7950;
								assign node7950 = (inp[11]) ? node8028 : node7951;
									assign node7951 = (inp[14]) ? node8001 : node7952;
										assign node7952 = (inp[2]) ? node7980 : node7953;
											assign node7953 = (inp[12]) ? node7969 : node7954;
												assign node7954 = (inp[13]) ? node7964 : node7955;
													assign node7955 = (inp[10]) ? node7957 : 4'b0101;
														assign node7957 = (inp[4]) ? node7959 : 4'b1001;
															assign node7959 = (inp[3]) ? 4'b1101 : node7960;
																assign node7960 = (inp[7]) ? 4'b1101 : 4'b1001;
													assign node7964 = (inp[10]) ? node7966 : 4'b1001;
														assign node7966 = (inp[3]) ? 4'b0101 : 4'b0001;
												assign node7969 = (inp[13]) ? node7975 : node7970;
													assign node7970 = (inp[3]) ? node7972 : 4'b0101;
														assign node7972 = (inp[10]) ? 4'b0101 : 4'b0001;
													assign node7975 = (inp[10]) ? 4'b1101 : node7976;
														assign node7976 = (inp[4]) ? 4'b1101 : 4'b1001;
											assign node7980 = (inp[3]) ? node7990 : node7981;
												assign node7981 = (inp[7]) ? 4'b0110 : node7982;
													assign node7982 = (inp[4]) ? node7986 : node7983;
														assign node7983 = (inp[13]) ? 4'b0001 : 4'b0110;
														assign node7986 = (inp[13]) ? 4'b1001 : 4'b0001;
												assign node7990 = (inp[13]) ? node7994 : node7991;
													assign node7991 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node7994 = (inp[10]) ? node7998 : node7995;
														assign node7995 = (inp[7]) ? 4'b1001 : 4'b1101;
														assign node7998 = (inp[12]) ? 4'b1101 : 4'b0101;
										assign node8001 = (inp[3]) ? node8011 : node8002;
											assign node8002 = (inp[2]) ? 4'b0110 : node8003;
												assign node8003 = (inp[4]) ? node8007 : node8004;
													assign node8004 = (inp[13]) ? 4'b1100 : 4'b0100;
													assign node8007 = (inp[10]) ? 4'b0000 : 4'b1000;
											assign node8011 = (inp[4]) ? node8019 : node8012;
												assign node8012 = (inp[10]) ? node8016 : node8013;
													assign node8013 = (inp[13]) ? 4'b1000 : 4'b0000;
													assign node8016 = (inp[7]) ? 4'b0000 : 4'b0100;
												assign node8019 = (inp[7]) ? node8025 : node8020;
													assign node8020 = (inp[12]) ? 4'b0100 : node8021;
														assign node8021 = (inp[2]) ? 4'b1100 : 4'b0100;
													assign node8025 = (inp[13]) ? 4'b0100 : 4'b0000;
									assign node8028 = (inp[3]) ? node8052 : node8029;
										assign node8029 = (inp[2]) ? node8043 : node8030;
											assign node8030 = (inp[7]) ? node8034 : node8031;
												assign node8031 = (inp[4]) ? 4'b1001 : 4'b1101;
												assign node8034 = (inp[12]) ? 4'b1101 : node8035;
													assign node8035 = (inp[10]) ? node8039 : node8036;
														assign node8036 = (inp[14]) ? 4'b1101 : 4'b0101;
														assign node8039 = (inp[13]) ? 4'b0001 : 4'b1101;
											assign node8043 = (inp[4]) ? node8045 : 4'b0110;
												assign node8045 = (inp[7]) ? node8049 : node8046;
													assign node8046 = (inp[13]) ? 4'b1001 : 4'b0001;
													assign node8049 = (inp[13]) ? 4'b0001 : 4'b0110;
										assign node8052 = (inp[4]) ? node8070 : node8053;
											assign node8053 = (inp[2]) ? node8059 : node8054;
												assign node8054 = (inp[13]) ? node8056 : 4'b0001;
													assign node8056 = (inp[14]) ? 4'b0001 : 4'b1001;
												assign node8059 = (inp[14]) ? node8065 : node8060;
													assign node8060 = (inp[13]) ? 4'b1001 : node8061;
														assign node8061 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node8065 = (inp[13]) ? node8067 : 4'b1001;
														assign node8067 = (inp[10]) ? 4'b0001 : 4'b1001;
											assign node8070 = (inp[7]) ? node8078 : node8071;
												assign node8071 = (inp[2]) ? 4'b1101 : node8072;
													assign node8072 = (inp[10]) ? 4'b0101 : node8073;
														assign node8073 = (inp[13]) ? 4'b1101 : 4'b0101;
												assign node8078 = (inp[13]) ? node8084 : node8079;
													assign node8079 = (inp[12]) ? 4'b0001 : node8080;
														assign node8080 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node8084 = (inp[12]) ? 4'b1001 : 4'b0101;
								assign node8087 = (inp[11]) ? node8163 : node8088;
									assign node8088 = (inp[14]) ? node8132 : node8089;
										assign node8089 = (inp[13]) ? node8107 : node8090;
											assign node8090 = (inp[3]) ? node8100 : node8091;
												assign node8091 = (inp[4]) ? node8093 : 4'b0110;
													assign node8093 = (inp[7]) ? node8097 : node8094;
														assign node8094 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node8097 = (inp[2]) ? 4'b0110 : 4'b1100;
												assign node8100 = (inp[4]) ? 4'b1100 : node8101;
													assign node8101 = (inp[10]) ? 4'b1000 : node8102;
														assign node8102 = (inp[12]) ? 4'b0000 : 4'b1000;
											assign node8107 = (inp[10]) ? node8123 : node8108;
												assign node8108 = (inp[12]) ? node8118 : node8109;
													assign node8109 = (inp[4]) ? 4'b0000 : node8110;
														assign node8110 = (inp[7]) ? node8114 : node8111;
															assign node8111 = (inp[3]) ? 4'b0100 : 4'b0000;
															assign node8114 = (inp[3]) ? 4'b0000 : 4'b0100;
													assign node8118 = (inp[3]) ? 4'b1000 : node8119;
														assign node8119 = (inp[7]) ? 4'b1100 : 4'b1000;
												assign node8123 = (inp[7]) ? node8125 : 4'b0000;
													assign node8125 = (inp[4]) ? node8129 : node8126;
														assign node8126 = (inp[3]) ? 4'b0000 : 4'b0100;
														assign node8129 = (inp[3]) ? 4'b0100 : 4'b0000;
										assign node8132 = (inp[3]) ? node8146 : node8133;
											assign node8133 = (inp[7]) ? node8139 : node8134;
												assign node8134 = (inp[12]) ? 4'b0001 : node8135;
													assign node8135 = (inp[13]) ? 4'b0001 : 4'b1001;
												assign node8139 = (inp[2]) ? node8143 : node8140;
													assign node8140 = (inp[13]) ? 4'b1101 : 4'b0101;
													assign node8143 = (inp[10]) ? 4'b0001 : 4'b0110;
											assign node8146 = (inp[10]) ? node8150 : node8147;
												assign node8147 = (inp[13]) ? 4'b1001 : 4'b0001;
												assign node8150 = (inp[12]) ? node8156 : node8151;
													assign node8151 = (inp[13]) ? 4'b0101 : node8152;
														assign node8152 = (inp[7]) ? 4'b1001 : 4'b1101;
													assign node8156 = (inp[13]) ? 4'b1001 : node8157;
														assign node8157 = (inp[7]) ? 4'b0001 : node8158;
															assign node8158 = (inp[4]) ? 4'b0101 : 4'b0001;
									assign node8163 = (inp[3]) ? node8187 : node8164;
										assign node8164 = (inp[7]) ? node8178 : node8165;
											assign node8165 = (inp[13]) ? 4'b0000 : node8166;
												assign node8166 = (inp[4]) ? node8172 : node8167;
													assign node8167 = (inp[2]) ? 4'b0110 : node8168;
														assign node8168 = (inp[12]) ? 4'b0100 : 4'b1100;
													assign node8172 = (inp[14]) ? 4'b1000 : node8173;
														assign node8173 = (inp[10]) ? 4'b1000 : 4'b0000;
											assign node8178 = (inp[2]) ? 4'b0110 : node8179;
												assign node8179 = (inp[14]) ? node8181 : 4'b1100;
													assign node8181 = (inp[12]) ? node8183 : 4'b0000;
														assign node8183 = (inp[13]) ? 4'b1100 : 4'b0100;
										assign node8187 = (inp[13]) ? node8197 : node8188;
											assign node8188 = (inp[10]) ? node8192 : node8189;
												assign node8189 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node8192 = (inp[4]) ? node8194 : 4'b1000;
													assign node8194 = (inp[7]) ? 4'b1000 : 4'b1100;
											assign node8197 = (inp[7]) ? node8199 : 4'b0100;
												assign node8199 = (inp[12]) ? node8203 : node8200;
													assign node8200 = (inp[4]) ? 4'b0100 : 4'b0000;
													assign node8203 = (inp[10]) ? 4'b0000 : 4'b1000;
					assign node8207 = (inp[5]) ? node8631 : node8208;
						assign node8208 = (inp[0]) ? node8502 : node8209;
							assign node8209 = (inp[11]) ? node8371 : node8210;
								assign node8210 = (inp[4]) ? node8282 : node8211;
									assign node8211 = (inp[3]) ? node8263 : node8212;
										assign node8212 = (inp[2]) ? node8236 : node8213;
											assign node8213 = (inp[13]) ? node8219 : node8214;
												assign node8214 = (inp[14]) ? 4'b0101 : node8215;
													assign node8215 = (inp[1]) ? 4'b0100 : 4'b0101;
												assign node8219 = (inp[7]) ? node8229 : node8220;
													assign node8220 = (inp[1]) ? node8224 : node8221;
														assign node8221 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node8224 = (inp[12]) ? 4'b1001 : node8225;
															assign node8225 = (inp[10]) ? 4'b0001 : 4'b1001;
													assign node8229 = (inp[14]) ? node8231 : 4'b0100;
														assign node8231 = (inp[12]) ? 4'b1101 : node8232;
															assign node8232 = (inp[10]) ? 4'b0001 : 4'b1101;
											assign node8236 = (inp[12]) ? node8252 : node8237;
												assign node8237 = (inp[14]) ? node8245 : node8238;
													assign node8238 = (inp[1]) ? node8242 : node8239;
														assign node8239 = (inp[10]) ? 4'b1101 : 4'b0101;
														assign node8242 = (inp[13]) ? 4'b0100 : 4'b1100;
													assign node8245 = (inp[1]) ? node8247 : 4'b0100;
														assign node8247 = (inp[10]) ? node8249 : 4'b0101;
															assign node8249 = (inp[7]) ? 4'b0101 : 4'b0001;
												assign node8252 = (inp[14]) ? node8260 : node8253;
													assign node8253 = (inp[1]) ? node8255 : 4'b1101;
														assign node8255 = (inp[10]) ? node8257 : 4'b0100;
															assign node8257 = (inp[13]) ? 4'b0100 : 4'b1100;
													assign node8260 = (inp[1]) ? 4'b1101 : 4'b1100;
										assign node8263 = (inp[2]) ? node8271 : node8264;
											assign node8264 = (inp[14]) ? 4'b1101 : node8265;
												assign node8265 = (inp[12]) ? node8267 : 4'b0001;
													assign node8267 = (inp[10]) ? 4'b1101 : 4'b0101;
											assign node8271 = (inp[10]) ? node8277 : node8272;
												assign node8272 = (inp[1]) ? 4'b0001 : node8273;
													assign node8273 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node8277 = (inp[12]) ? node8279 : 4'b0001;
													assign node8279 = (inp[13]) ? 4'b1001 : 4'b1000;
									assign node8282 = (inp[10]) ? node8328 : node8283;
										assign node8283 = (inp[13]) ? node8297 : node8284;
											assign node8284 = (inp[12]) ? node8292 : node8285;
												assign node8285 = (inp[1]) ? 4'b1001 : node8286;
													assign node8286 = (inp[3]) ? 4'b0001 : node8287;
														assign node8287 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node8292 = (inp[3]) ? 4'b0001 : node8293;
													assign node8293 = (inp[14]) ? 4'b0001 : 4'b0100;
											assign node8297 = (inp[7]) ? node8317 : node8298;
												assign node8298 = (inp[2]) ? node8308 : node8299;
													assign node8299 = (inp[3]) ? node8303 : node8300;
														assign node8300 = (inp[1]) ? 4'b1101 : 4'b0101;
														assign node8303 = (inp[14]) ? node8305 : 4'b0100;
															assign node8305 = (inp[12]) ? 4'b0100 : 4'b1001;
													assign node8308 = (inp[3]) ? 4'b0101 : node8309;
														assign node8309 = (inp[1]) ? node8311 : 4'b1001;
															assign node8311 = (inp[14]) ? 4'b1001 : node8312;
																assign node8312 = (inp[12]) ? 4'b1000 : 4'b0000;
												assign node8317 = (inp[12]) ? 4'b0001 : node8318;
													assign node8318 = (inp[3]) ? node8320 : 4'b1100;
														assign node8320 = (inp[2]) ? 4'b0001 : node8321;
															assign node8321 = (inp[1]) ? 4'b0000 : node8322;
																assign node8322 = (inp[14]) ? 4'b1001 : 4'b0000;
										assign node8328 = (inp[12]) ? node8350 : node8329;
											assign node8329 = (inp[1]) ? node8343 : node8330;
												assign node8330 = (inp[3]) ? node8336 : node8331;
													assign node8331 = (inp[2]) ? 4'b0001 : node8332;
														assign node8332 = (inp[13]) ? 4'b1101 : 4'b1001;
													assign node8336 = (inp[14]) ? 4'b1001 : node8337;
														assign node8337 = (inp[13]) ? node8339 : 4'b0000;
															assign node8339 = (inp[7]) ? 4'b1000 : 4'b1100;
												assign node8343 = (inp[7]) ? node8345 : 4'b0101;
													assign node8345 = (inp[13]) ? 4'b0100 : node8346;
														assign node8346 = (inp[3]) ? 4'b1000 : 4'b1101;
											assign node8350 = (inp[1]) ? node8362 : node8351;
												assign node8351 = (inp[3]) ? node8357 : node8352;
													assign node8352 = (inp[7]) ? 4'b0100 : node8353;
														assign node8353 = (inp[14]) ? 4'b1000 : 4'b1001;
													assign node8357 = (inp[13]) ? node8359 : 4'b1001;
														assign node8359 = (inp[2]) ? 4'b1101 : 4'b1000;
												assign node8362 = (inp[7]) ? node8364 : 4'b1000;
													assign node8364 = (inp[2]) ? 4'b1001 : node8365;
														assign node8365 = (inp[3]) ? node8367 : 4'b1001;
															assign node8367 = (inp[13]) ? 4'b1000 : 4'b0000;
								assign node8371 = (inp[1]) ? node8441 : node8372;
									assign node8372 = (inp[13]) ? node8406 : node8373;
										assign node8373 = (inp[4]) ? node8385 : node8374;
											assign node8374 = (inp[3]) ? node8376 : 4'b0101;
												assign node8376 = (inp[2]) ? 4'b0001 : node8377;
													assign node8377 = (inp[12]) ? node8381 : node8378;
														assign node8378 = (inp[7]) ? 4'b0100 : 4'b1100;
														assign node8381 = (inp[10]) ? 4'b1100 : 4'b0100;
											assign node8385 = (inp[10]) ? node8397 : node8386;
												assign node8386 = (inp[12]) ? 4'b0000 : node8387;
													assign node8387 = (inp[3]) ? node8391 : node8388;
														assign node8388 = (inp[7]) ? 4'b0101 : 4'b1000;
														assign node8391 = (inp[2]) ? 4'b1000 : node8392;
															assign node8392 = (inp[7]) ? 4'b1000 : 4'b1001;
												assign node8397 = (inp[12]) ? 4'b0001 : node8398;
													assign node8398 = (inp[3]) ? node8402 : node8399;
														assign node8399 = (inp[2]) ? 4'b1001 : 4'b0100;
														assign node8402 = (inp[2]) ? 4'b0100 : 4'b0001;
										assign node8406 = (inp[2]) ? node8426 : node8407;
											assign node8407 = (inp[3]) ? node8417 : node8408;
												assign node8408 = (inp[7]) ? node8412 : node8409;
													assign node8409 = (inp[4]) ? 4'b0100 : 4'b0000;
													assign node8412 = (inp[4]) ? node8414 : 4'b1101;
														assign node8414 = (inp[14]) ? 4'b0100 : 4'b1000;
												assign node8417 = (inp[4]) ? node8419 : 4'b1100;
													assign node8419 = (inp[7]) ? node8423 : node8420;
														assign node8420 = (inp[10]) ? 4'b1101 : 4'b1001;
														assign node8423 = (inp[10]) ? 4'b1001 : 4'b0001;
											assign node8426 = (inp[3]) ? node8434 : node8427;
												assign node8427 = (inp[12]) ? node8429 : 4'b1001;
													assign node8429 = (inp[7]) ? 4'b1101 : node8430;
														assign node8430 = (inp[4]) ? 4'b1001 : 4'b1101;
												assign node8434 = (inp[7]) ? node8438 : node8435;
													assign node8435 = (inp[4]) ? 4'b1100 : 4'b1000;
													assign node8438 = (inp[4]) ? 4'b1000 : 4'b1001;
									assign node8441 = (inp[13]) ? node8483 : node8442;
										assign node8442 = (inp[3]) ? node8458 : node8443;
											assign node8443 = (inp[12]) ? node8449 : node8444;
												assign node8444 = (inp[7]) ? 4'b1100 : node8445;
													assign node8445 = (inp[4]) ? 4'b1000 : 4'b1100;
												assign node8449 = (inp[7]) ? node8455 : node8450;
													assign node8450 = (inp[14]) ? 4'b1100 : node8451;
														assign node8451 = (inp[4]) ? 4'b1000 : 4'b0000;
													assign node8455 = (inp[10]) ? 4'b0000 : 4'b0100;
											assign node8458 = (inp[10]) ? node8468 : node8459;
												assign node8459 = (inp[4]) ? node8463 : node8460;
													assign node8460 = (inp[2]) ? 4'b1000 : 4'b1100;
													assign node8463 = (inp[2]) ? 4'b1000 : node8464;
														assign node8464 = (inp[7]) ? 4'b1000 : 4'b0000;
												assign node8468 = (inp[7]) ? node8474 : node8469;
													assign node8469 = (inp[4]) ? node8471 : 4'b0000;
														assign node8471 = (inp[2]) ? 4'b0100 : 4'b1000;
													assign node8474 = (inp[12]) ? node8476 : 4'b1000;
														assign node8476 = (inp[2]) ? node8480 : node8477;
															assign node8477 = (inp[4]) ? 4'b1000 : 4'b0100;
															assign node8480 = (inp[4]) ? 4'b0000 : 4'b1000;
										assign node8483 = (inp[10]) ? node8497 : node8484;
											assign node8484 = (inp[12]) ? node8492 : node8485;
												assign node8485 = (inp[14]) ? 4'b0000 : node8486;
													assign node8486 = (inp[4]) ? node8488 : 4'b1000;
														assign node8488 = (inp[7]) ? 4'b1000 : 4'b1100;
												assign node8492 = (inp[3]) ? node8494 : 4'b1100;
													assign node8494 = (inp[2]) ? 4'b1100 : 4'b0100;
											assign node8497 = (inp[4]) ? node8499 : 4'b0000;
												assign node8499 = (inp[3]) ? 4'b0100 : 4'b0000;
							assign node8502 = (inp[2]) ? 4'b0100 : node8503;
								assign node8503 = (inp[3]) ? node8547 : node8504;
									assign node8504 = (inp[4]) ? node8516 : node8505;
										assign node8505 = (inp[13]) ? node8507 : 4'b0100;
											assign node8507 = (inp[11]) ? 4'b0100 : node8508;
												assign node8508 = (inp[7]) ? 4'b0100 : node8509;
													assign node8509 = (inp[14]) ? node8511 : 4'b0100;
														assign node8511 = (inp[10]) ? 4'b0001 : 4'b0100;
										assign node8516 = (inp[7]) ? node8540 : node8517;
											assign node8517 = (inp[1]) ? node8533 : node8518;
												assign node8518 = (inp[12]) ? node8528 : node8519;
													assign node8519 = (inp[14]) ? node8525 : node8520;
														assign node8520 = (inp[10]) ? 4'b0001 : node8521;
															assign node8521 = (inp[13]) ? 4'b1001 : 4'b0001;
														assign node8525 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node8528 = (inp[14]) ? node8530 : 4'b0001;
														assign node8530 = (inp[11]) ? 4'b0001 : 4'b0000;
												assign node8533 = (inp[11]) ? node8537 : node8534;
													assign node8534 = (inp[14]) ? 4'b0001 : 4'b0000;
													assign node8537 = (inp[12]) ? 4'b1000 : 4'b0000;
											assign node8540 = (inp[1]) ? node8542 : 4'b0100;
												assign node8542 = (inp[10]) ? node8544 : 4'b0100;
													assign node8544 = (inp[14]) ? 4'b0100 : 4'b0000;
									assign node8547 = (inp[7]) ? node8593 : node8548;
										assign node8548 = (inp[4]) ? node8570 : node8549;
											assign node8549 = (inp[13]) ? node8561 : node8550;
												assign node8550 = (inp[12]) ? node8552 : 4'b1001;
													assign node8552 = (inp[1]) ? node8556 : node8553;
														assign node8553 = (inp[10]) ? 4'b0000 : 4'b0001;
														assign node8556 = (inp[11]) ? node8558 : 4'b0001;
															assign node8558 = (inp[10]) ? 4'b1000 : 4'b0000;
												assign node8561 = (inp[1]) ? node8567 : node8562;
													assign node8562 = (inp[11]) ? 4'b1001 : node8563;
														assign node8563 = (inp[10]) ? 4'b0100 : 4'b1000;
													assign node8567 = (inp[14]) ? 4'b0101 : 4'b0100;
											assign node8570 = (inp[14]) ? node8576 : node8571;
												assign node8571 = (inp[1]) ? 4'b0100 : node8572;
													assign node8572 = (inp[12]) ? 4'b0101 : 4'b1101;
												assign node8576 = (inp[11]) ? node8584 : node8577;
													assign node8577 = (inp[1]) ? 4'b1101 : node8578;
														assign node8578 = (inp[13]) ? 4'b1100 : node8579;
															assign node8579 = (inp[12]) ? 4'b0100 : 4'b1100;
													assign node8584 = (inp[1]) ? node8586 : 4'b0101;
														assign node8586 = (inp[13]) ? node8590 : node8587;
															assign node8587 = (inp[10]) ? 4'b1100 : 4'b0100;
															assign node8590 = (inp[12]) ? 4'b1100 : 4'b0100;
										assign node8593 = (inp[1]) ? node8615 : node8594;
											assign node8594 = (inp[10]) ? node8606 : node8595;
												assign node8595 = (inp[13]) ? node8601 : node8596;
													assign node8596 = (inp[11]) ? 4'b0001 : node8597;
														assign node8597 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node8601 = (inp[12]) ? node8603 : 4'b1001;
														assign node8603 = (inp[14]) ? 4'b1000 : 4'b1001;
												assign node8606 = (inp[13]) ? node8610 : node8607;
													assign node8607 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node8610 = (inp[14]) ? node8612 : 4'b0101;
														assign node8612 = (inp[11]) ? 4'b0101 : 4'b0100;
											assign node8615 = (inp[11]) ? node8625 : node8616;
												assign node8616 = (inp[14]) ? node8622 : node8617;
													assign node8617 = (inp[13]) ? 4'b0100 : node8618;
														assign node8618 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node8622 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node8625 = (inp[13]) ? node8627 : 4'b1000;
													assign node8627 = (inp[4]) ? 4'b1000 : 4'b0000;
						assign node8631 = (inp[3]) ? node8957 : node8632;
							assign node8632 = (inp[4]) ? node8790 : node8633;
								assign node8633 = (inp[2]) ? node8733 : node8634;
									assign node8634 = (inp[0]) ? node8678 : node8635;
										assign node8635 = (inp[1]) ? node8661 : node8636;
											assign node8636 = (inp[13]) ? node8650 : node8637;
												assign node8637 = (inp[7]) ? node8645 : node8638;
													assign node8638 = (inp[10]) ? node8640 : 4'b0101;
														assign node8640 = (inp[14]) ? 4'b1000 : node8641;
															assign node8641 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node8645 = (inp[12]) ? 4'b0101 : node8646;
														assign node8646 = (inp[14]) ? 4'b0101 : 4'b1100;
												assign node8650 = (inp[12]) ? node8652 : 4'b1000;
													assign node8652 = (inp[11]) ? node8656 : node8653;
														assign node8653 = (inp[14]) ? 4'b0000 : 4'b0100;
														assign node8656 = (inp[10]) ? node8658 : 4'b1000;
															assign node8658 = (inp[7]) ? 4'b1000 : 4'b1100;
											assign node8661 = (inp[12]) ? node8671 : node8662;
												assign node8662 = (inp[10]) ? 4'b0100 : node8663;
													assign node8663 = (inp[7]) ? node8667 : node8664;
														assign node8664 = (inp[13]) ? 4'b0100 : 4'b0000;
														assign node8667 = (inp[14]) ? 4'b0100 : 4'b0000;
												assign node8671 = (inp[10]) ? 4'b0000 : node8672;
													assign node8672 = (inp[7]) ? 4'b1100 : node8673;
														assign node8673 = (inp[11]) ? 4'b0100 : 4'b1000;
										assign node8678 = (inp[7]) ? node8696 : node8679;
											assign node8679 = (inp[11]) ? node8685 : node8680;
												assign node8680 = (inp[12]) ? node8682 : 4'b0001;
													assign node8682 = (inp[13]) ? 4'b1001 : 4'b0101;
												assign node8685 = (inp[13]) ? node8693 : node8686;
													assign node8686 = (inp[14]) ? 4'b0101 : node8687;
														assign node8687 = (inp[1]) ? node8689 : 4'b0000;
															assign node8689 = (inp[12]) ? 4'b0100 : 4'b1100;
													assign node8693 = (inp[1]) ? 4'b1000 : 4'b0000;
											assign node8696 = (inp[1]) ? node8718 : node8697;
												assign node8697 = (inp[14]) ? node8713 : node8698;
													assign node8698 = (inp[11]) ? node8708 : node8699;
														assign node8699 = (inp[12]) ? node8705 : node8700;
															assign node8700 = (inp[10]) ? node8702 : 4'b1101;
																assign node8702 = (inp[13]) ? 4'b0101 : 4'b1101;
															assign node8705 = (inp[13]) ? 4'b1101 : 4'b0101;
														assign node8708 = (inp[12]) ? node8710 : 4'b0000;
															assign node8710 = (inp[13]) ? 4'b1101 : 4'b0101;
													assign node8713 = (inp[13]) ? 4'b1100 : node8714;
														assign node8714 = (inp[11]) ? 4'b0101 : 4'b0100;
												assign node8718 = (inp[14]) ? node8726 : node8719;
													assign node8719 = (inp[13]) ? node8721 : 4'b1100;
														assign node8721 = (inp[10]) ? 4'b0100 : node8722;
															assign node8722 = (inp[12]) ? 4'b1100 : 4'b0100;
													assign node8726 = (inp[11]) ? node8728 : 4'b1101;
														assign node8728 = (inp[10]) ? node8730 : 4'b1100;
															assign node8730 = (inp[13]) ? 4'b0000 : 4'b1100;
									assign node8733 = (inp[0]) ? node8775 : node8734;
										assign node8734 = (inp[11]) ? node8762 : node8735;
											assign node8735 = (inp[13]) ? node8749 : node8736;
												assign node8736 = (inp[10]) ? node8742 : node8737;
													assign node8737 = (inp[12]) ? 4'b0101 : node8738;
														assign node8738 = (inp[1]) ? 4'b1101 : 4'b0101;
													assign node8742 = (inp[14]) ? 4'b1101 : node8743;
														assign node8743 = (inp[12]) ? node8745 : 4'b1001;
															assign node8745 = (inp[1]) ? 4'b0001 : 4'b0000;
												assign node8749 = (inp[10]) ? 4'b1001 : node8750;
													assign node8750 = (inp[7]) ? node8758 : node8751;
														assign node8751 = (inp[1]) ? 4'b0001 : node8752;
															assign node8752 = (inp[12]) ? node8754 : 4'b0000;
																assign node8754 = (inp[14]) ? 4'b1001 : 4'b1000;
														assign node8758 = (inp[1]) ? 4'b0000 : 4'b0101;
											assign node8762 = (inp[13]) ? node8768 : node8763;
												assign node8763 = (inp[1]) ? node8765 : 4'b0100;
													assign node8765 = (inp[10]) ? 4'b0100 : 4'b1100;
												assign node8768 = (inp[1]) ? node8770 : 4'b1001;
													assign node8770 = (inp[12]) ? node8772 : 4'b0000;
														assign node8772 = (inp[10]) ? 4'b0100 : 4'b0000;
										assign node8775 = (inp[7]) ? 4'b0100 : node8776;
											assign node8776 = (inp[13]) ? node8778 : 4'b0100;
												assign node8778 = (inp[10]) ? node8784 : node8779;
													assign node8779 = (inp[1]) ? node8781 : 4'b0100;
														assign node8781 = (inp[12]) ? 4'b0100 : 4'b0000;
													assign node8784 = (inp[1]) ? node8786 : 4'b0001;
														assign node8786 = (inp[14]) ? 4'b0100 : 4'b0000;
								assign node8790 = (inp[2]) ? node8888 : node8791;
									assign node8791 = (inp[11]) ? node8847 : node8792;
										assign node8792 = (inp[10]) ? node8822 : node8793;
											assign node8793 = (inp[13]) ? node8805 : node8794;
												assign node8794 = (inp[0]) ? node8802 : node8795;
													assign node8795 = (inp[7]) ? node8799 : node8796;
														assign node8796 = (inp[12]) ? 4'b1001 : 4'b1000;
														assign node8799 = (inp[14]) ? 4'b1100 : 4'b0100;
													assign node8802 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node8805 = (inp[14]) ? node8819 : node8806;
													assign node8806 = (inp[7]) ? node8814 : node8807;
														assign node8807 = (inp[0]) ? 4'b0101 : node8808;
															assign node8808 = (inp[1]) ? 4'b0001 : node8809;
																assign node8809 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node8814 = (inp[0]) ? 4'b1001 : node8815;
															assign node8815 = (inp[12]) ? 4'b1001 : 4'b0101;
													assign node8819 = (inp[0]) ? 4'b0000 : 4'b0001;
											assign node8822 = (inp[1]) ? node8836 : node8823;
												assign node8823 = (inp[0]) ? node8831 : node8824;
													assign node8824 = (inp[7]) ? 4'b1000 : node8825;
														assign node8825 = (inp[12]) ? 4'b1001 : node8826;
															assign node8826 = (inp[14]) ? 4'b1000 : 4'b1001;
													assign node8831 = (inp[13]) ? node8833 : 4'b1001;
														assign node8833 = (inp[12]) ? 4'b1000 : 4'b1001;
												assign node8836 = (inp[12]) ? node8842 : node8837;
													assign node8837 = (inp[0]) ? node8839 : 4'b1001;
														assign node8839 = (inp[7]) ? 4'b0001 : 4'b0101;
													assign node8842 = (inp[7]) ? 4'b1001 : node8843;
														assign node8843 = (inp[14]) ? 4'b1000 : 4'b1001;
										assign node8847 = (inp[1]) ? node8869 : node8848;
											assign node8848 = (inp[13]) ? node8858 : node8849;
												assign node8849 = (inp[0]) ? node8851 : 4'b1001;
													assign node8851 = (inp[14]) ? 4'b0000 : node8852;
														assign node8852 = (inp[12]) ? 4'b1000 : node8853;
															assign node8853 = (inp[10]) ? 4'b0100 : 4'b1000;
												assign node8858 = (inp[14]) ? 4'b1001 : node8859;
													assign node8859 = (inp[12]) ? node8863 : node8860;
														assign node8860 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node8863 = (inp[10]) ? 4'b0001 : node8864;
															assign node8864 = (inp[7]) ? 4'b0101 : 4'b0100;
											assign node8869 = (inp[10]) ? node8877 : node8870;
												assign node8870 = (inp[13]) ? 4'b1000 : node8871;
													assign node8871 = (inp[12]) ? node8873 : 4'b1000;
														assign node8873 = (inp[0]) ? 4'b1000 : 4'b0000;
												assign node8877 = (inp[7]) ? node8883 : node8878;
													assign node8878 = (inp[13]) ? 4'b0000 : node8879;
														assign node8879 = (inp[0]) ? 4'b0100 : 4'b0000;
													assign node8883 = (inp[0]) ? 4'b0000 : node8884;
														assign node8884 = (inp[13]) ? 4'b0000 : 4'b1000;
									assign node8888 = (inp[7]) ? node8924 : node8889;
										assign node8889 = (inp[14]) ? node8913 : node8890;
											assign node8890 = (inp[0]) ? node8908 : node8891;
												assign node8891 = (inp[10]) ? node8901 : node8892;
													assign node8892 = (inp[12]) ? node8896 : node8893;
														assign node8893 = (inp[1]) ? 4'b0000 : 4'b1000;
														assign node8896 = (inp[13]) ? node8898 : 4'b0100;
															assign node8898 = (inp[11]) ? 4'b0100 : 4'b1000;
													assign node8901 = (inp[1]) ? node8905 : node8902;
														assign node8902 = (inp[11]) ? 4'b1000 : 4'b0000;
														assign node8905 = (inp[12]) ? 4'b1000 : 4'b0000;
												assign node8908 = (inp[1]) ? node8910 : 4'b0001;
													assign node8910 = (inp[13]) ? 4'b0000 : 4'b1000;
											assign node8913 = (inp[1]) ? node8921 : node8914;
												assign node8914 = (inp[11]) ? 4'b0001 : node8915;
													assign node8915 = (inp[0]) ? 4'b1000 : node8916;
														assign node8916 = (inp[13]) ? 4'b0000 : 4'b1000;
												assign node8921 = (inp[0]) ? 4'b0001 : 4'b1001;
										assign node8924 = (inp[0]) ? node8946 : node8925;
											assign node8925 = (inp[13]) ? node8937 : node8926;
												assign node8926 = (inp[11]) ? node8934 : node8927;
													assign node8927 = (inp[12]) ? node8929 : 4'b0101;
														assign node8929 = (inp[14]) ? node8931 : 4'b1001;
															assign node8931 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node8934 = (inp[10]) ? 4'b0000 : 4'b0100;
												assign node8937 = (inp[12]) ? node8939 : 4'b1000;
													assign node8939 = (inp[1]) ? node8943 : node8940;
														assign node8940 = (inp[11]) ? 4'b1000 : 4'b0000;
														assign node8943 = (inp[11]) ? 4'b0000 : 4'b1000;
											assign node8946 = (inp[13]) ? node8948 : 4'b0100;
												assign node8948 = (inp[11]) ? node8954 : node8949;
													assign node8949 = (inp[1]) ? node8951 : 4'b0100;
														assign node8951 = (inp[14]) ? 4'b0100 : 4'b0000;
													assign node8954 = (inp[1]) ? 4'b0000 : 4'b0001;
							assign node8957 = (inp[11]) ? node9111 : node8958;
								assign node8958 = (inp[4]) ? node9038 : node8959;
									assign node8959 = (inp[2]) ? node8999 : node8960;
										assign node8960 = (inp[10]) ? node8980 : node8961;
											assign node8961 = (inp[1]) ? node8975 : node8962;
												assign node8962 = (inp[14]) ? 4'b0001 : node8963;
													assign node8963 = (inp[13]) ? node8967 : node8964;
														assign node8964 = (inp[7]) ? 4'b1000 : 4'b0000;
														assign node8967 = (inp[0]) ? node8969 : 4'b0001;
															assign node8969 = (inp[7]) ? node8971 : 4'b0001;
																assign node8971 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node8975 = (inp[7]) ? node8977 : 4'b1000;
													assign node8977 = (inp[0]) ? 4'b1000 : 4'b1001;
											assign node8980 = (inp[14]) ? node8990 : node8981;
												assign node8981 = (inp[7]) ? 4'b0000 : node8982;
													assign node8982 = (inp[0]) ? node8984 : 4'b0001;
														assign node8984 = (inp[12]) ? 4'b0000 : node8985;
															assign node8985 = (inp[1]) ? 4'b0000 : 4'b1000;
												assign node8990 = (inp[13]) ? node8994 : node8991;
													assign node8991 = (inp[0]) ? 4'b0000 : 4'b1000;
													assign node8994 = (inp[1]) ? node8996 : 4'b0000;
														assign node8996 = (inp[0]) ? 4'b1001 : 4'b0001;
										assign node8999 = (inp[1]) ? node9019 : node9000;
											assign node9000 = (inp[12]) ? node9014 : node9001;
												assign node9001 = (inp[7]) ? node9005 : node9002;
													assign node9002 = (inp[14]) ? 4'b1000 : 4'b1001;
													assign node9005 = (inp[0]) ? 4'b1001 : node9006;
														assign node9006 = (inp[14]) ? node9008 : 4'b0000;
															assign node9008 = (inp[10]) ? node9010 : 4'b0001;
																assign node9010 = (inp[13]) ? 4'b1000 : 4'b0001;
												assign node9014 = (inp[10]) ? node9016 : 4'b0000;
													assign node9016 = (inp[14]) ? 4'b1000 : 4'b0001;
											assign node9019 = (inp[13]) ? node9029 : node9020;
												assign node9020 = (inp[0]) ? node9024 : node9021;
													assign node9021 = (inp[7]) ? 4'b1001 : 4'b0001;
													assign node9024 = (inp[14]) ? 4'b0001 : node9025;
														assign node9025 = (inp[10]) ? 4'b0001 : 4'b1000;
												assign node9029 = (inp[12]) ? node9031 : 4'b0001;
													assign node9031 = (inp[0]) ? 4'b1001 : node9032;
														assign node9032 = (inp[14]) ? 4'b1000 : node9033;
															assign node9033 = (inp[7]) ? 4'b1001 : 4'b1000;
									assign node9038 = (inp[13]) ? node9086 : node9039;
										assign node9039 = (inp[7]) ? node9063 : node9040;
											assign node9040 = (inp[12]) ? node9050 : node9041;
												assign node9041 = (inp[0]) ? node9045 : node9042;
													assign node9042 = (inp[1]) ? 4'b1000 : 4'b0000;
													assign node9045 = (inp[2]) ? 4'b1000 : node9046;
														assign node9046 = (inp[14]) ? 4'b1000 : 4'b0000;
												assign node9050 = (inp[10]) ? node9056 : node9051;
													assign node9051 = (inp[1]) ? 4'b1000 : node9052;
														assign node9052 = (inp[0]) ? 4'b0001 : 4'b0000;
													assign node9056 = (inp[2]) ? node9058 : 4'b0001;
														assign node9058 = (inp[0]) ? node9060 : 4'b0000;
															assign node9060 = (inp[14]) ? 4'b0001 : 4'b0000;
											assign node9063 = (inp[2]) ? node9069 : node9064;
												assign node9064 = (inp[0]) ? 4'b1000 : node9065;
													assign node9065 = (inp[14]) ? 4'b0001 : 4'b0000;
												assign node9069 = (inp[10]) ? node9077 : node9070;
													assign node9070 = (inp[14]) ? 4'b1001 : node9071;
														assign node9071 = (inp[1]) ? node9073 : 4'b1001;
															assign node9073 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node9077 = (inp[1]) ? node9083 : node9078;
														assign node9078 = (inp[0]) ? node9080 : 4'b1001;
															assign node9080 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node9083 = (inp[0]) ? 4'b0000 : 4'b1000;
										assign node9086 = (inp[10]) ? node9102 : node9087;
											assign node9087 = (inp[0]) ? node9099 : node9088;
												assign node9088 = (inp[7]) ? 4'b0001 : node9089;
													assign node9089 = (inp[1]) ? node9095 : node9090;
														assign node9090 = (inp[2]) ? node9092 : 4'b0001;
															assign node9092 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node9095 = (inp[12]) ? 4'b0001 : 4'b0000;
												assign node9099 = (inp[1]) ? 4'b0001 : 4'b0000;
											assign node9102 = (inp[1]) ? 4'b0000 : node9103;
												assign node9103 = (inp[2]) ? 4'b0000 : node9104;
													assign node9104 = (inp[12]) ? node9106 : 4'b0001;
														assign node9106 = (inp[14]) ? 4'b0001 : 4'b0000;
								assign node9111 = (inp[1]) ? node9181 : node9112;
									assign node9112 = (inp[4]) ? node9158 : node9113;
										assign node9113 = (inp[7]) ? node9131 : node9114;
											assign node9114 = (inp[2]) ? node9122 : node9115;
												assign node9115 = (inp[10]) ? node9117 : 4'b0001;
													assign node9117 = (inp[0]) ? 4'b1000 : node9118;
														assign node9118 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node9122 = (inp[0]) ? node9128 : node9123;
													assign node9123 = (inp[10]) ? node9125 : 4'b0000;
														assign node9125 = (inp[14]) ? 4'b1000 : 4'b0000;
													assign node9128 = (inp[13]) ? 4'b0000 : 4'b0001;
											assign node9131 = (inp[13]) ? node9141 : node9132;
												assign node9132 = (inp[0]) ? 4'b0001 : node9133;
													assign node9133 = (inp[10]) ? 4'b1000 : node9134;
														assign node9134 = (inp[12]) ? 4'b1001 : node9135;
															assign node9135 = (inp[2]) ? 4'b1001 : 4'b0001;
												assign node9141 = (inp[0]) ? node9147 : node9142;
													assign node9142 = (inp[2]) ? node9144 : 4'b1000;
														assign node9144 = (inp[10]) ? 4'b0000 : 4'b0001;
													assign node9147 = (inp[10]) ? node9151 : node9148;
														assign node9148 = (inp[2]) ? 4'b1001 : 4'b1000;
														assign node9151 = (inp[14]) ? 4'b1001 : node9152;
															assign node9152 = (inp[12]) ? node9154 : 4'b0000;
																assign node9154 = (inp[2]) ? 4'b1001 : 4'b0001;
										assign node9158 = (inp[13]) ? 4'b0000 : node9159;
											assign node9159 = (inp[0]) ? node9163 : node9160;
												assign node9160 = (inp[10]) ? 4'b0000 : 4'b1000;
												assign node9163 = (inp[2]) ? node9173 : node9164;
													assign node9164 = (inp[10]) ? node9168 : node9165;
														assign node9165 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node9168 = (inp[7]) ? node9170 : 4'b0001;
															assign node9170 = (inp[12]) ? 4'b0001 : 4'b0000;
													assign node9173 = (inp[12]) ? node9177 : node9174;
														assign node9174 = (inp[7]) ? 4'b0001 : 4'b1001;
														assign node9177 = (inp[14]) ? 4'b0000 : 4'b1000;
									assign node9181 = (inp[10]) ? node9221 : node9182;
										assign node9182 = (inp[2]) ? node9202 : node9183;
											assign node9183 = (inp[7]) ? node9191 : node9184;
												assign node9184 = (inp[13]) ? node9186 : 4'b0000;
													assign node9186 = (inp[0]) ? node9188 : 4'b0000;
														assign node9188 = (inp[12]) ? 4'b1000 : 4'b0000;
												assign node9191 = (inp[13]) ? node9197 : node9192;
													assign node9192 = (inp[4]) ? 4'b1000 : node9193;
														assign node9193 = (inp[14]) ? 4'b1000 : 4'b0000;
													assign node9197 = (inp[4]) ? 4'b0000 : node9198;
														assign node9198 = (inp[14]) ? 4'b1000 : 4'b0000;
											assign node9202 = (inp[0]) ? node9206 : node9203;
												assign node9203 = (inp[13]) ? 4'b0000 : 4'b1000;
												assign node9206 = (inp[4]) ? node9216 : node9207;
													assign node9207 = (inp[13]) ? node9211 : node9208;
														assign node9208 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node9211 = (inp[12]) ? 4'b1000 : node9212;
															assign node9212 = (inp[7]) ? 4'b0000 : 4'b1000;
													assign node9216 = (inp[12]) ? node9218 : 4'b0000;
														assign node9218 = (inp[7]) ? 4'b1000 : 4'b0000;
										assign node9221 = (inp[4]) ? 4'b0000 : node9222;
											assign node9222 = (inp[13]) ? 4'b0000 : node9223;
												assign node9223 = (inp[0]) ? node9227 : node9224;
													assign node9224 = (inp[14]) ? 4'b0000 : 4'b1000;
													assign node9227 = (inp[2]) ? node9229 : 4'b0000;
														assign node9229 = (inp[7]) ? 4'b1000 : 4'b0000;
				assign node9234 = (inp[0]) ? node10068 : node9235;
					assign node9235 = (inp[6]) ? node9481 : node9236;
						assign node9236 = (inp[2]) ? node9430 : node9237;
							assign node9237 = (inp[5]) ? node9275 : node9238;
								assign node9238 = (inp[3]) ? node9240 : 4'b0010;
									assign node9240 = (inp[4]) ? node9250 : node9241;
										assign node9241 = (inp[13]) ? node9243 : 4'b0010;
											assign node9243 = (inp[11]) ? node9245 : 4'b0010;
												assign node9245 = (inp[10]) ? node9247 : 4'b0010;
													assign node9247 = (inp[1]) ? 4'b0000 : 4'b0010;
										assign node9250 = (inp[7]) ? node9270 : node9251;
											assign node9251 = (inp[1]) ? node9257 : node9252;
												assign node9252 = (inp[11]) ? node9254 : 4'b1001;
													assign node9254 = (inp[14]) ? 4'b1001 : 4'b0001;
												assign node9257 = (inp[14]) ? node9265 : node9258;
													assign node9258 = (inp[13]) ? node9262 : node9259;
														assign node9259 = (inp[11]) ? 4'b0000 : 4'b1000;
														assign node9262 = (inp[12]) ? 4'b1000 : 4'b0000;
													assign node9265 = (inp[11]) ? node9267 : 4'b1001;
														assign node9267 = (inp[13]) ? 4'b0000 : 4'b1000;
											assign node9270 = (inp[13]) ? node9272 : 4'b0010;
												assign node9272 = (inp[1]) ? 4'b0000 : 4'b0010;
								assign node9275 = (inp[1]) ? node9349 : node9276;
									assign node9276 = (inp[11]) ? node9324 : node9277;
										assign node9277 = (inp[14]) ? node9299 : node9278;
											assign node9278 = (inp[4]) ? node9288 : node9279;
												assign node9279 = (inp[7]) ? 4'b0001 : node9280;
													assign node9280 = (inp[10]) ? node9282 : 4'b1101;
														assign node9282 = (inp[3]) ? node9284 : 4'b0101;
															assign node9284 = (inp[12]) ? 4'b0101 : 4'b1101;
												assign node9288 = (inp[3]) ? node9294 : node9289;
													assign node9289 = (inp[10]) ? 4'b0101 : node9290;
														assign node9290 = (inp[13]) ? 4'b1001 : 4'b0001;
													assign node9294 = (inp[12]) ? 4'b1001 : node9295;
														assign node9295 = (inp[13]) ? 4'b0001 : 4'b1001;
											assign node9299 = (inp[3]) ? node9315 : node9300;
												assign node9300 = (inp[7]) ? node9306 : node9301;
													assign node9301 = (inp[10]) ? 4'b0100 : node9302;
														assign node9302 = (inp[4]) ? 4'b0100 : 4'b0000;
													assign node9306 = (inp[10]) ? node9308 : 4'b1000;
														assign node9308 = (inp[13]) ? node9312 : node9309;
															assign node9309 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node9312 = (inp[4]) ? 4'b0100 : 4'b0000;
												assign node9315 = (inp[13]) ? node9319 : node9316;
													assign node9316 = (inp[7]) ? 4'b0100 : 4'b1100;
													assign node9319 = (inp[7]) ? 4'b1100 : node9320;
														assign node9320 = (inp[4]) ? 4'b1000 : 4'b0000;
										assign node9324 = (inp[3]) ? node9336 : node9325;
											assign node9325 = (inp[7]) ? node9327 : 4'b1001;
												assign node9327 = (inp[13]) ? node9333 : node9328;
													assign node9328 = (inp[12]) ? 4'b0001 : node9329;
														assign node9329 = (inp[4]) ? 4'b0001 : 4'b1001;
													assign node9333 = (inp[4]) ? 4'b1001 : 4'b0001;
											assign node9336 = (inp[7]) ? node9344 : node9337;
												assign node9337 = (inp[10]) ? node9341 : node9338;
													assign node9338 = (inp[13]) ? 4'b1001 : 4'b0001;
													assign node9341 = (inp[12]) ? 4'b0101 : 4'b0001;
												assign node9344 = (inp[13]) ? 4'b1101 : node9345;
													assign node9345 = (inp[12]) ? 4'b0101 : 4'b1101;
									assign node9349 = (inp[11]) ? node9389 : node9350;
										assign node9350 = (inp[14]) ? node9372 : node9351;
											assign node9351 = (inp[4]) ? node9357 : node9352;
												assign node9352 = (inp[10]) ? 4'b0100 : node9353;
													assign node9353 = (inp[7]) ? 4'b0000 : 4'b0100;
												assign node9357 = (inp[3]) ? node9361 : node9358;
													assign node9358 = (inp[12]) ? 4'b1100 : 4'b0100;
													assign node9361 = (inp[7]) ? 4'b1100 : node9362;
														assign node9362 = (inp[12]) ? node9364 : 4'b1000;
															assign node9364 = (inp[13]) ? node9368 : node9365;
																assign node9365 = (inp[10]) ? 4'b1000 : 4'b0000;
																assign node9368 = (inp[10]) ? 4'b0000 : 4'b1000;
											assign node9372 = (inp[13]) ? node9382 : node9373;
												assign node9373 = (inp[12]) ? node9377 : node9374;
													assign node9374 = (inp[10]) ? 4'b1101 : 4'b0101;
													assign node9377 = (inp[4]) ? node9379 : 4'b0001;
														assign node9379 = (inp[10]) ? 4'b0101 : 4'b0001;
												assign node9382 = (inp[10]) ? node9384 : 4'b1101;
													assign node9384 = (inp[4]) ? 4'b0001 : node9385;
														assign node9385 = (inp[12]) ? 4'b1101 : 4'b0101;
										assign node9389 = (inp[13]) ? node9405 : node9390;
											assign node9390 = (inp[3]) ? node9394 : node9391;
												assign node9391 = (inp[7]) ? 4'b1000 : 4'b0000;
												assign node9394 = (inp[14]) ? node9396 : 4'b1100;
													assign node9396 = (inp[7]) ? node9402 : node9397;
														assign node9397 = (inp[10]) ? 4'b1000 : node9398;
															assign node9398 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node9402 = (inp[12]) ? 4'b0100 : 4'b1100;
											assign node9405 = (inp[12]) ? node9413 : node9406;
												assign node9406 = (inp[3]) ? node9408 : 4'b0100;
													assign node9408 = (inp[4]) ? 4'b0000 : node9409;
														assign node9409 = (inp[7]) ? 4'b0100 : 4'b0000;
												assign node9413 = (inp[10]) ? node9425 : node9414;
													assign node9414 = (inp[4]) ? node9416 : 4'b1100;
														assign node9416 = (inp[14]) ? 4'b1000 : node9417;
															assign node9417 = (inp[3]) ? node9421 : node9418;
																assign node9418 = (inp[7]) ? 4'b1000 : 4'b1100;
																assign node9421 = (inp[7]) ? 4'b1100 : 4'b1000;
													assign node9425 = (inp[14]) ? node9427 : 4'b0000;
														assign node9427 = (inp[3]) ? 4'b0100 : 4'b0000;
							assign node9430 = (inp[5]) ? node9432 : 4'b0010;
								assign node9432 = (inp[3]) ? node9434 : 4'b0010;
									assign node9434 = (inp[4]) ? node9450 : node9435;
										assign node9435 = (inp[13]) ? node9437 : 4'b0010;
											assign node9437 = (inp[7]) ? 4'b0010 : node9438;
												assign node9438 = (inp[14]) ? node9442 : node9439;
													assign node9439 = (inp[1]) ? 4'b0000 : 4'b0001;
													assign node9442 = (inp[10]) ? node9444 : 4'b0010;
														assign node9444 = (inp[11]) ? node9446 : 4'b0010;
															assign node9446 = (inp[1]) ? 4'b0000 : 4'b0010;
										assign node9450 = (inp[7]) ? node9472 : node9451;
											assign node9451 = (inp[13]) ? node9461 : node9452;
												assign node9452 = (inp[10]) ? 4'b1000 : node9453;
													assign node9453 = (inp[1]) ? node9455 : 4'b0001;
														assign node9455 = (inp[14]) ? 4'b0001 : node9456;
															assign node9456 = (inp[11]) ? 4'b0000 : 4'b1000;
												assign node9461 = (inp[11]) ? node9469 : node9462;
													assign node9462 = (inp[12]) ? node9464 : 4'b1001;
														assign node9464 = (inp[10]) ? 4'b1001 : node9465;
															assign node9465 = (inp[1]) ? 4'b1001 : 4'b1000;
													assign node9469 = (inp[10]) ? 4'b0000 : 4'b1001;
											assign node9472 = (inp[12]) ? 4'b0010 : node9473;
												assign node9473 = (inp[10]) ? node9475 : 4'b0010;
													assign node9475 = (inp[13]) ? node9477 : 4'b0010;
														assign node9477 = (inp[11]) ? 4'b0001 : 4'b0000;
						assign node9481 = (inp[5]) ? node9765 : node9482;
							assign node9482 = (inp[1]) ? node9628 : node9483;
								assign node9483 = (inp[3]) ? node9549 : node9484;
									assign node9484 = (inp[14]) ? node9506 : node9485;
										assign node9485 = (inp[7]) ? node9499 : node9486;
											assign node9486 = (inp[2]) ? 4'b0101 : node9487;
												assign node9487 = (inp[13]) ? 4'b1001 : node9488;
													assign node9488 = (inp[4]) ? node9494 : node9489;
														assign node9489 = (inp[10]) ? node9491 : 4'b0001;
															assign node9491 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node9494 = (inp[10]) ? 4'b1101 : 4'b0101;
											assign node9499 = (inp[13]) ? 4'b1001 : node9500;
												assign node9500 = (inp[10]) ? node9502 : 4'b0001;
													assign node9502 = (inp[12]) ? 4'b0001 : 4'b1001;
										assign node9506 = (inp[11]) ? node9528 : node9507;
											assign node9507 = (inp[2]) ? node9513 : node9508;
												assign node9508 = (inp[7]) ? node9510 : 4'b1001;
													assign node9510 = (inp[13]) ? 4'b1000 : 4'b0000;
												assign node9513 = (inp[13]) ? node9519 : node9514;
													assign node9514 = (inp[10]) ? node9516 : 4'b0000;
														assign node9516 = (inp[7]) ? 4'b1000 : 4'b0000;
													assign node9519 = (inp[10]) ? node9523 : node9520;
														assign node9520 = (inp[7]) ? 4'b1000 : 4'b1100;
														assign node9523 = (inp[4]) ? 4'b0100 : node9524;
															assign node9524 = (inp[7]) ? 4'b0000 : 4'b0100;
											assign node9528 = (inp[2]) ? node9542 : node9529;
												assign node9529 = (inp[7]) ? node9535 : node9530;
													assign node9530 = (inp[13]) ? node9532 : 4'b0000;
														assign node9532 = (inp[4]) ? 4'b1000 : 4'b1001;
													assign node9535 = (inp[4]) ? node9537 : 4'b1001;
														assign node9537 = (inp[13]) ? 4'b1001 : node9538;
															assign node9538 = (inp[10]) ? 4'b1001 : 4'b0001;
												assign node9542 = (inp[13]) ? node9544 : 4'b0001;
													assign node9544 = (inp[12]) ? node9546 : 4'b0101;
														assign node9546 = (inp[4]) ? 4'b1101 : 4'b1001;
									assign node9549 = (inp[10]) ? node9595 : node9550;
										assign node9550 = (inp[11]) ? node9570 : node9551;
											assign node9551 = (inp[2]) ? node9561 : node9552;
												assign node9552 = (inp[13]) ? node9556 : node9553;
													assign node9553 = (inp[4]) ? 4'b0101 : 4'b0001;
													assign node9556 = (inp[4]) ? node9558 : 4'b0101;
														assign node9558 = (inp[7]) ? 4'b0101 : 4'b0001;
												assign node9561 = (inp[14]) ? node9567 : node9562;
													assign node9562 = (inp[13]) ? node9564 : 4'b0101;
														assign node9564 = (inp[12]) ? 4'b1101 : 4'b0001;
													assign node9567 = (inp[13]) ? 4'b1100 : 4'b0100;
											assign node9570 = (inp[2]) ? node9586 : node9571;
												assign node9571 = (inp[12]) ? node9575 : node9572;
													assign node9572 = (inp[4]) ? 4'b0001 : 4'b1000;
													assign node9575 = (inp[4]) ? node9581 : node9576;
														assign node9576 = (inp[13]) ? node9578 : 4'b0000;
															assign node9578 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node9581 = (inp[14]) ? 4'b0100 : node9582;
															assign node9582 = (inp[13]) ? 4'b0000 : 4'b0100;
												assign node9586 = (inp[13]) ? node9592 : node9587;
													assign node9587 = (inp[7]) ? 4'b0101 : node9588;
														assign node9588 = (inp[12]) ? 4'b0001 : 4'b0101;
													assign node9592 = (inp[14]) ? 4'b0000 : 4'b1000;
										assign node9595 = (inp[11]) ? node9617 : node9596;
											assign node9596 = (inp[2]) ? node9606 : node9597;
												assign node9597 = (inp[4]) ? node9601 : node9598;
													assign node9598 = (inp[7]) ? 4'b1001 : 4'b1101;
													assign node9601 = (inp[7]) ? 4'b1101 : node9602;
														assign node9602 = (inp[13]) ? 4'b1001 : 4'b1101;
												assign node9606 = (inp[4]) ? node9612 : node9607;
													assign node9607 = (inp[14]) ? 4'b1100 : node9608;
														assign node9608 = (inp[13]) ? 4'b0101 : 4'b1101;
													assign node9612 = (inp[13]) ? 4'b0000 : node9613;
														assign node9613 = (inp[12]) ? 4'b0001 : 4'b1001;
											assign node9617 = (inp[2]) ? node9625 : node9618;
												assign node9618 = (inp[12]) ? node9620 : 4'b0000;
													assign node9620 = (inp[7]) ? 4'b1000 : node9621;
														assign node9621 = (inp[14]) ? 4'b1100 : 4'b1000;
												assign node9625 = (inp[4]) ? 4'b1101 : 4'b0101;
								assign node9628 = (inp[11]) ? node9702 : node9629;
									assign node9629 = (inp[14]) ? node9671 : node9630;
										assign node9630 = (inp[2]) ? node9652 : node9631;
											assign node9631 = (inp[3]) ? node9641 : node9632;
												assign node9632 = (inp[7]) ? node9638 : node9633;
													assign node9633 = (inp[4]) ? node9635 : 4'b0100;
														assign node9635 = (inp[13]) ? 4'b0001 : 4'b0100;
													assign node9638 = (inp[4]) ? 4'b0100 : 4'b1000;
												assign node9641 = (inp[7]) ? node9645 : node9642;
													assign node9642 = (inp[13]) ? 4'b1101 : 4'b0101;
													assign node9645 = (inp[4]) ? node9649 : node9646;
														assign node9646 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node9649 = (inp[12]) ? 4'b0101 : 4'b0001;
											assign node9652 = (inp[13]) ? node9662 : node9653;
												assign node9653 = (inp[3]) ? node9659 : node9654;
													assign node9654 = (inp[10]) ? 4'b1000 : node9655;
														assign node9655 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node9659 = (inp[7]) ? 4'b1100 : 4'b1000;
												assign node9662 = (inp[10]) ? node9666 : node9663;
													assign node9663 = (inp[12]) ? 4'b1100 : 4'b0100;
													assign node9666 = (inp[7]) ? 4'b0000 : node9667;
														assign node9667 = (inp[3]) ? 4'b0000 : 4'b0100;
										assign node9671 = (inp[4]) ? node9687 : node9672;
											assign node9672 = (inp[3]) ? node9680 : node9673;
												assign node9673 = (inp[13]) ? node9677 : node9674;
													assign node9674 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node9677 = (inp[7]) ? 4'b0001 : 4'b0101;
												assign node9680 = (inp[10]) ? 4'b0101 : node9681;
													assign node9681 = (inp[12]) ? 4'b0101 : node9682;
														assign node9682 = (inp[13]) ? 4'b1101 : 4'b1001;
											assign node9687 = (inp[2]) ? node9691 : node9688;
												assign node9688 = (inp[3]) ? 4'b0000 : 4'b0001;
												assign node9691 = (inp[12]) ? node9693 : 4'b0001;
													assign node9693 = (inp[13]) ? 4'b1101 : node9694;
														assign node9694 = (inp[10]) ? 4'b0101 : node9695;
															assign node9695 = (inp[7]) ? 4'b0001 : node9696;
																assign node9696 = (inp[3]) ? 4'b0001 : 4'b0101;
									assign node9702 = (inp[10]) ? node9738 : node9703;
										assign node9703 = (inp[2]) ? node9717 : node9704;
											assign node9704 = (inp[4]) ? node9710 : node9705;
												assign node9705 = (inp[13]) ? node9707 : 4'b1000;
													assign node9707 = (inp[7]) ? 4'b1000 : 4'b1100;
												assign node9710 = (inp[13]) ? node9712 : 4'b0000;
													assign node9712 = (inp[3]) ? node9714 : 4'b1000;
														assign node9714 = (inp[12]) ? 4'b0000 : 4'b1000;
											assign node9717 = (inp[12]) ? node9727 : node9718;
												assign node9718 = (inp[13]) ? node9724 : node9719;
													assign node9719 = (inp[3]) ? 4'b1100 : node9720;
														assign node9720 = (inp[7]) ? 4'b1000 : 4'b1100;
													assign node9724 = (inp[3]) ? 4'b0000 : 4'b0100;
												assign node9727 = (inp[13]) ? node9733 : node9728;
													assign node9728 = (inp[3]) ? node9730 : 4'b0000;
														assign node9730 = (inp[4]) ? 4'b0000 : 4'b0100;
													assign node9733 = (inp[7]) ? 4'b1000 : node9734;
														assign node9734 = (inp[3]) ? 4'b1000 : 4'b1100;
										assign node9738 = (inp[13]) ? node9756 : node9739;
											assign node9739 = (inp[2]) ? node9745 : node9740;
												assign node9740 = (inp[7]) ? 4'b0100 : node9741;
													assign node9741 = (inp[4]) ? 4'b0000 : 4'b1000;
												assign node9745 = (inp[12]) ? node9749 : node9746;
													assign node9746 = (inp[4]) ? 4'b0000 : 4'b1100;
													assign node9749 = (inp[3]) ? 4'b1100 : node9750;
														assign node9750 = (inp[4]) ? node9752 : 4'b1000;
															assign node9752 = (inp[7]) ? 4'b1000 : 4'b1100;
											assign node9756 = (inp[4]) ? node9762 : node9757;
												assign node9757 = (inp[3]) ? 4'b0100 : node9758;
													assign node9758 = (inp[12]) ? 4'b0100 : 4'b0000;
												assign node9762 = (inp[3]) ? 4'b0000 : 4'b0100;
							assign node9765 = (inp[11]) ? node9947 : node9766;
								assign node9766 = (inp[3]) ? node9856 : node9767;
									assign node9767 = (inp[4]) ? node9819 : node9768;
										assign node9768 = (inp[2]) ? node9798 : node9769;
											assign node9769 = (inp[13]) ? node9785 : node9770;
												assign node9770 = (inp[7]) ? node9778 : node9771;
													assign node9771 = (inp[10]) ? 4'b0100 : node9772;
														assign node9772 = (inp[1]) ? 4'b1001 : node9773;
															assign node9773 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node9778 = (inp[10]) ? node9782 : node9779;
														assign node9779 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node9782 = (inp[1]) ? 4'b0001 : 4'b1001;
												assign node9785 = (inp[1]) ? node9793 : node9786;
													assign node9786 = (inp[14]) ? node9788 : 4'b1000;
														assign node9788 = (inp[7]) ? node9790 : 4'b1101;
															assign node9790 = (inp[10]) ? 4'b1101 : 4'b1001;
													assign node9793 = (inp[10]) ? 4'b0000 : node9794;
														assign node9794 = (inp[14]) ? 4'b0100 : 4'b0101;
											assign node9798 = (inp[10]) ? node9808 : node9799;
												assign node9799 = (inp[13]) ? node9805 : node9800;
													assign node9800 = (inp[12]) ? 4'b0001 : node9801;
														assign node9801 = (inp[14]) ? 4'b1001 : 4'b0001;
													assign node9805 = (inp[7]) ? 4'b0001 : 4'b0101;
												assign node9808 = (inp[12]) ? node9814 : node9809;
													assign node9809 = (inp[7]) ? node9811 : 4'b0000;
														assign node9811 = (inp[13]) ? 4'b0101 : 4'b0001;
													assign node9814 = (inp[7]) ? 4'b1001 : node9815;
														assign node9815 = (inp[13]) ? 4'b1101 : 4'b1001;
										assign node9819 = (inp[13]) ? node9839 : node9820;
											assign node9820 = (inp[12]) ? node9832 : node9821;
												assign node9821 = (inp[2]) ? node9827 : node9822;
													assign node9822 = (inp[1]) ? node9824 : 4'b1000;
														assign node9824 = (inp[14]) ? 4'b0100 : 4'b1000;
													assign node9827 = (inp[7]) ? 4'b1101 : node9828;
														assign node9828 = (inp[14]) ? 4'b1000 : 4'b1001;
												assign node9832 = (inp[2]) ? node9834 : 4'b1000;
													assign node9834 = (inp[1]) ? node9836 : 4'b0000;
														assign node9836 = (inp[10]) ? 4'b0000 : 4'b0101;
											assign node9839 = (inp[2]) ? node9847 : node9840;
												assign node9840 = (inp[12]) ? node9844 : node9841;
													assign node9841 = (inp[1]) ? 4'b1001 : 4'b0001;
													assign node9844 = (inp[1]) ? 4'b0001 : 4'b0100;
												assign node9847 = (inp[7]) ? node9849 : 4'b1000;
													assign node9849 = (inp[1]) ? node9853 : node9850;
														assign node9850 = (inp[14]) ? 4'b1001 : 4'b1000;
														assign node9853 = (inp[12]) ? 4'b1001 : 4'b0001;
									assign node9856 = (inp[2]) ? node9908 : node9857;
										assign node9857 = (inp[10]) ? node9889 : node9858;
											assign node9858 = (inp[7]) ? node9872 : node9859;
												assign node9859 = (inp[1]) ? node9869 : node9860;
													assign node9860 = (inp[14]) ? node9862 : 4'b0001;
														assign node9862 = (inp[13]) ? 4'b0000 : node9863;
															assign node9863 = (inp[12]) ? node9865 : 4'b0001;
																assign node9865 = (inp[4]) ? 4'b1000 : 4'b0001;
													assign node9869 = (inp[13]) ? 4'b0001 : 4'b0000;
												assign node9872 = (inp[1]) ? node9880 : node9873;
													assign node9873 = (inp[4]) ? node9877 : node9874;
														assign node9874 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node9877 = (inp[12]) ? 4'b1000 : 4'b0000;
													assign node9880 = (inp[4]) ? 4'b0001 : node9881;
														assign node9881 = (inp[13]) ? node9883 : 4'b0001;
															assign node9883 = (inp[12]) ? node9885 : 4'b1000;
																assign node9885 = (inp[14]) ? 4'b0001 : 4'b0000;
											assign node9889 = (inp[1]) ? node9901 : node9890;
												assign node9890 = (inp[4]) ? node9898 : node9891;
													assign node9891 = (inp[14]) ? 4'b0001 : node9892;
														assign node9892 = (inp[12]) ? 4'b0000 : node9893;
															assign node9893 = (inp[7]) ? 4'b0001 : 4'b0000;
													assign node9898 = (inp[13]) ? 4'b0000 : 4'b1000;
												assign node9901 = (inp[12]) ? 4'b0000 : node9902;
													assign node9902 = (inp[14]) ? 4'b1000 : node9903;
														assign node9903 = (inp[13]) ? 4'b1001 : 4'b1000;
										assign node9908 = (inp[14]) ? node9934 : node9909;
											assign node9909 = (inp[12]) ? node9919 : node9910;
												assign node9910 = (inp[10]) ? 4'b0001 : node9911;
													assign node9911 = (inp[4]) ? node9913 : 4'b0001;
														assign node9913 = (inp[1]) ? node9915 : 4'b1000;
															assign node9915 = (inp[13]) ? 4'b0000 : 4'b0001;
												assign node9919 = (inp[7]) ? node9923 : node9920;
													assign node9920 = (inp[4]) ? 4'b0000 : 4'b1000;
													assign node9923 = (inp[13]) ? node9929 : node9924;
														assign node9924 = (inp[10]) ? node9926 : 4'b1000;
															assign node9926 = (inp[4]) ? 4'b0001 : 4'b0000;
														assign node9929 = (inp[4]) ? node9931 : 4'b1001;
															assign node9931 = (inp[10]) ? 4'b0000 : 4'b0001;
											assign node9934 = (inp[4]) ? 4'b0000 : node9935;
												assign node9935 = (inp[7]) ? node9941 : node9936;
													assign node9936 = (inp[13]) ? node9938 : 4'b1000;
														assign node9938 = (inp[10]) ? 4'b1000 : 4'b0001;
													assign node9941 = (inp[1]) ? node9943 : 4'b0000;
														assign node9943 = (inp[10]) ? 4'b0001 : 4'b1000;
								assign node9947 = (inp[1]) ? node10013 : node9948;
									assign node9948 = (inp[3]) ? node9986 : node9949;
										assign node9949 = (inp[2]) ? node9967 : node9950;
											assign node9950 = (inp[13]) ? node9960 : node9951;
												assign node9951 = (inp[4]) ? node9957 : node9952;
													assign node9952 = (inp[12]) ? 4'b0001 : node9953;
														assign node9953 = (inp[10]) ? 4'b0001 : 4'b1001;
													assign node9957 = (inp[14]) ? 4'b1000 : 4'b0001;
												assign node9960 = (inp[12]) ? node9962 : 4'b0101;
													assign node9962 = (inp[14]) ? 4'b1000 : node9963;
														assign node9963 = (inp[7]) ? 4'b1001 : 4'b0001;
											assign node9967 = (inp[4]) ? node9979 : node9968;
												assign node9968 = (inp[12]) ? node9974 : node9969;
													assign node9969 = (inp[10]) ? 4'b0100 : node9970;
														assign node9970 = (inp[13]) ? 4'b1100 : 4'b1000;
													assign node9974 = (inp[10]) ? 4'b1000 : node9975;
														assign node9975 = (inp[7]) ? 4'b0000 : 4'b0100;
												assign node9979 = (inp[10]) ? 4'b1001 : node9980;
													assign node9980 = (inp[12]) ? 4'b0001 : node9981;
														assign node9981 = (inp[14]) ? 4'b0101 : 4'b0001;
										assign node9986 = (inp[7]) ? node10000 : node9987;
											assign node9987 = (inp[12]) ? node9995 : node9988;
												assign node9988 = (inp[2]) ? node9992 : node9989;
													assign node9989 = (inp[10]) ? 4'b0000 : 4'b0001;
													assign node9992 = (inp[13]) ? 4'b0000 : 4'b1000;
												assign node9995 = (inp[2]) ? node9997 : 4'b1000;
													assign node9997 = (inp[4]) ? 4'b0000 : 4'b1000;
											assign node10000 = (inp[10]) ? node10008 : node10001;
												assign node10001 = (inp[12]) ? node10003 : 4'b0000;
													assign node10003 = (inp[13]) ? node10005 : 4'b1001;
														assign node10005 = (inp[2]) ? 4'b0001 : 4'b0000;
												assign node10008 = (inp[12]) ? node10010 : 4'b0001;
													assign node10010 = (inp[4]) ? 4'b0000 : 4'b0001;
									assign node10013 = (inp[4]) ? node10053 : node10014;
										assign node10014 = (inp[10]) ? node10038 : node10015;
											assign node10015 = (inp[14]) ? node10031 : node10016;
												assign node10016 = (inp[12]) ? node10024 : node10017;
													assign node10017 = (inp[2]) ? node10021 : node10018;
														assign node10018 = (inp[13]) ? 4'b0000 : 4'b0100;
														assign node10021 = (inp[3]) ? 4'b1000 : 4'b1100;
													assign node10024 = (inp[2]) ? node10028 : node10025;
														assign node10025 = (inp[3]) ? 4'b1000 : 4'b0000;
														assign node10028 = (inp[3]) ? 4'b0000 : 4'b1000;
												assign node10031 = (inp[13]) ? 4'b1000 : node10032;
													assign node10032 = (inp[12]) ? 4'b1000 : node10033;
														assign node10033 = (inp[2]) ? 4'b1000 : 4'b0000;
											assign node10038 = (inp[13]) ? node10048 : node10039;
												assign node10039 = (inp[12]) ? node10045 : node10040;
													assign node10040 = (inp[7]) ? node10042 : 4'b1100;
														assign node10042 = (inp[3]) ? 4'b1000 : 4'b0000;
													assign node10045 = (inp[3]) ? 4'b0000 : 4'b1000;
												assign node10048 = (inp[2]) ? node10050 : 4'b0000;
													assign node10050 = (inp[3]) ? 4'b0000 : 4'b0100;
										assign node10053 = (inp[12]) ? node10055 : 4'b0000;
											assign node10055 = (inp[3]) ? node10063 : node10056;
												assign node10056 = (inp[7]) ? 4'b1000 : node10057;
													assign node10057 = (inp[13]) ? node10059 : 4'b0100;
														assign node10059 = (inp[14]) ? 4'b1000 : 4'b0000;
												assign node10063 = (inp[2]) ? node10065 : 4'b0000;
													assign node10065 = (inp[10]) ? 4'b0000 : 4'b1000;
					assign node10068 = (inp[6]) ? node10070 : 4'b0000;
						assign node10070 = (inp[2]) ? node10270 : node10071;
							assign node10071 = (inp[5]) ? node10103 : node10072;
								assign node10072 = (inp[3]) ? node10074 : 4'b0000;
									assign node10074 = (inp[7]) ? 4'b0000 : node10075;
										assign node10075 = (inp[4]) ? node10083 : node10076;
											assign node10076 = (inp[12]) ? 4'b0000 : node10077;
												assign node10077 = (inp[13]) ? node10079 : 4'b0000;
													assign node10079 = (inp[10]) ? 4'b0001 : 4'b0000;
											assign node10083 = (inp[11]) ? node10099 : node10084;
												assign node10084 = (inp[1]) ? node10092 : node10085;
													assign node10085 = (inp[14]) ? 4'b1000 : node10086;
														assign node10086 = (inp[13]) ? 4'b0001 : node10087;
															assign node10087 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node10092 = (inp[14]) ? node10096 : node10093;
														assign node10093 = (inp[13]) ? 4'b0000 : 4'b1000;
														assign node10096 = (inp[13]) ? 4'b1001 : 4'b0001;
												assign node10099 = (inp[12]) ? 4'b1000 : 4'b1001;
								assign node10103 = (inp[11]) ? node10213 : node10104;
									assign node10104 = (inp[3]) ? node10162 : node10105;
										assign node10105 = (inp[12]) ? node10145 : node10106;
											assign node10106 = (inp[10]) ? node10136 : node10107;
												assign node10107 = (inp[4]) ? node10121 : node10108;
													assign node10108 = (inp[7]) ? node10116 : node10109;
														assign node10109 = (inp[13]) ? node10113 : node10110;
															assign node10110 = (inp[14]) ? 4'b0000 : 4'b1000;
															assign node10113 = (inp[1]) ? 4'b1001 : 4'b1000;
														assign node10116 = (inp[13]) ? 4'b0000 : node10117;
															assign node10117 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node10121 = (inp[1]) ? node10129 : node10122;
														assign node10122 = (inp[13]) ? node10126 : node10123;
															assign node10123 = (inp[7]) ? 4'b0001 : 4'b0101;
															assign node10126 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node10129 = (inp[7]) ? node10133 : node10130;
															assign node10130 = (inp[13]) ? 4'b1001 : 4'b1100;
															assign node10133 = (inp[13]) ? 4'b0100 : 4'b1000;
												assign node10136 = (inp[4]) ? node10142 : node10137;
													assign node10137 = (inp[14]) ? 4'b1001 : node10138;
														assign node10138 = (inp[1]) ? 4'b0100 : 4'b0101;
													assign node10142 = (inp[1]) ? 4'b0001 : 4'b1001;
											assign node10145 = (inp[13]) ? node10157 : node10146;
												assign node10146 = (inp[4]) ? node10152 : node10147;
													assign node10147 = (inp[14]) ? 4'b0001 : node10148;
														assign node10148 = (inp[1]) ? 4'b0000 : 4'b0001;
													assign node10152 = (inp[10]) ? 4'b0101 : node10153;
														assign node10153 = (inp[14]) ? 4'b0100 : 4'b0101;
												assign node10157 = (inp[4]) ? node10159 : 4'b1001;
													assign node10159 = (inp[10]) ? 4'b1001 : 4'b0001;
										assign node10162 = (inp[13]) ? node10188 : node10163;
											assign node10163 = (inp[4]) ? node10173 : node10164;
												assign node10164 = (inp[1]) ? node10170 : node10165;
													assign node10165 = (inp[10]) ? node10167 : 4'b0001;
														assign node10167 = (inp[14]) ? 4'b0001 : 4'b0000;
													assign node10170 = (inp[10]) ? 4'b1001 : 4'b0001;
												assign node10173 = (inp[1]) ? node10179 : node10174;
													assign node10174 = (inp[10]) ? node10176 : 4'b1000;
														assign node10176 = (inp[14]) ? 4'b0001 : 4'b1001;
													assign node10179 = (inp[14]) ? node10185 : node10180;
														assign node10180 = (inp[10]) ? node10182 : 4'b0000;
															assign node10182 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node10185 = (inp[10]) ? 4'b0000 : 4'b0001;
											assign node10188 = (inp[7]) ? node10194 : node10189;
												assign node10189 = (inp[14]) ? node10191 : 4'b0000;
													assign node10191 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node10194 = (inp[1]) ? node10202 : node10195;
													assign node10195 = (inp[4]) ? 4'b0001 : node10196;
														assign node10196 = (inp[12]) ? 4'b0001 : node10197;
															assign node10197 = (inp[14]) ? 4'b1001 : 4'b1000;
													assign node10202 = (inp[10]) ? 4'b0000 : node10203;
														assign node10203 = (inp[4]) ? node10207 : node10204;
															assign node10204 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node10207 = (inp[14]) ? node10209 : 4'b0000;
																assign node10209 = (inp[12]) ? 4'b0000 : 4'b0001;
									assign node10213 = (inp[1]) ? node10237 : node10214;
										assign node10214 = (inp[3]) ? node10222 : node10215;
											assign node10215 = (inp[7]) ? 4'b0001 : node10216;
												assign node10216 = (inp[4]) ? 4'b0000 : node10217;
													assign node10217 = (inp[12]) ? 4'b1001 : 4'b0101;
											assign node10222 = (inp[4]) ? node10232 : node10223;
												assign node10223 = (inp[10]) ? node10229 : node10224;
													assign node10224 = (inp[13]) ? 4'b0001 : node10225;
														assign node10225 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node10229 = (inp[7]) ? 4'b1001 : 4'b1000;
												assign node10232 = (inp[13]) ? 4'b0000 : node10233;
													assign node10233 = (inp[14]) ? 4'b0000 : 4'b1000;
										assign node10237 = (inp[10]) ? node10259 : node10238;
											assign node10238 = (inp[13]) ? node10248 : node10239;
												assign node10239 = (inp[3]) ? node10241 : 4'b0000;
													assign node10241 = (inp[14]) ? node10245 : node10242;
														assign node10242 = (inp[7]) ? 4'b1000 : 4'b0000;
														assign node10245 = (inp[7]) ? 4'b0000 : 4'b1000;
												assign node10248 = (inp[3]) ? node10256 : node10249;
													assign node10249 = (inp[12]) ? 4'b1000 : node10250;
														assign node10250 = (inp[7]) ? 4'b0100 : node10251;
															assign node10251 = (inp[14]) ? 4'b0100 : 4'b1000;
													assign node10256 = (inp[7]) ? 4'b1000 : 4'b0000;
											assign node10259 = (inp[4]) ? 4'b0000 : node10260;
												assign node10260 = (inp[13]) ? node10264 : node10261;
													assign node10261 = (inp[14]) ? 4'b0000 : 4'b1000;
													assign node10264 = (inp[7]) ? 4'b0000 : node10265;
														assign node10265 = (inp[12]) ? 4'b0000 : 4'b0100;
							assign node10270 = (inp[4]) ? node10272 : 4'b0000;
								assign node10272 = (inp[3]) ? node10274 : 4'b0000;
									assign node10274 = (inp[7]) ? 4'b0000 : node10275;
										assign node10275 = (inp[5]) ? node10277 : 4'b0000;
											assign node10277 = (inp[1]) ? node10287 : node10278;
												assign node10278 = (inp[10]) ? node10280 : 4'b0001;
													assign node10280 = (inp[12]) ? 4'b0001 : node10281;
														assign node10281 = (inp[13]) ? 4'b0000 : node10282;
															assign node10282 = (inp[11]) ? 4'b0000 : 4'b1001;
												assign node10287 = (inp[13]) ? 4'b0000 : node10288;
													assign node10288 = (inp[12]) ? 4'b1000 : node10289;
														assign node10289 = (inp[11]) ? 4'b1000 : 4'b0001;

endmodule