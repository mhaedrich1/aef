module dtc_split5_bm75 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node7;
	wire [3-1:0] node8;
	wire [3-1:0] node9;
	wire [3-1:0] node12;
	wire [3-1:0] node15;
	wire [3-1:0] node16;
	wire [3-1:0] node20;
	wire [3-1:0] node21;
	wire [3-1:0] node22;
	wire [3-1:0] node25;
	wire [3-1:0] node28;
	wire [3-1:0] node29;
	wire [3-1:0] node32;
	wire [3-1:0] node35;
	wire [3-1:0] node36;
	wire [3-1:0] node37;
	wire [3-1:0] node38;
	wire [3-1:0] node41;
	wire [3-1:0] node44;
	wire [3-1:0] node45;
	wire [3-1:0] node48;
	wire [3-1:0] node51;
	wire [3-1:0] node52;
	wire [3-1:0] node54;
	wire [3-1:0] node57;
	wire [3-1:0] node59;
	wire [3-1:0] node62;
	wire [3-1:0] node63;
	wire [3-1:0] node64;
	wire [3-1:0] node66;
	wire [3-1:0] node67;
	wire [3-1:0] node72;
	wire [3-1:0] node73;
	wire [3-1:0] node74;
	wire [3-1:0] node75;
	wire [3-1:0] node79;
	wire [3-1:0] node81;
	wire [3-1:0] node84;
	wire [3-1:0] node86;
	wire [3-1:0] node87;
	wire [3-1:0] node91;
	wire [3-1:0] node92;
	wire [3-1:0] node93;
	wire [3-1:0] node95;
	wire [3-1:0] node96;
	wire [3-1:0] node97;
	wire [3-1:0] node102;
	wire [3-1:0] node103;
	wire [3-1:0] node104;
	wire [3-1:0] node105;
	wire [3-1:0] node110;
	wire [3-1:0] node111;
	wire [3-1:0] node112;
	wire [3-1:0] node116;
	wire [3-1:0] node117;
	wire [3-1:0] node121;
	wire [3-1:0] node122;
	wire [3-1:0] node123;
	wire [3-1:0] node125;
	wire [3-1:0] node127;
	wire [3-1:0] node132;
	wire [3-1:0] node133;
	wire [3-1:0] node134;
	wire [3-1:0] node135;
	wire [3-1:0] node136;
	wire [3-1:0] node137;
	wire [3-1:0] node138;
	wire [3-1:0] node141;
	wire [3-1:0] node145;
	wire [3-1:0] node146;
	wire [3-1:0] node147;
	wire [3-1:0] node151;
	wire [3-1:0] node152;
	wire [3-1:0] node155;
	wire [3-1:0] node158;
	wire [3-1:0] node159;
	wire [3-1:0] node160;
	wire [3-1:0] node162;
	wire [3-1:0] node165;
	wire [3-1:0] node167;
	wire [3-1:0] node170;
	wire [3-1:0] node171;
	wire [3-1:0] node172;
	wire [3-1:0] node175;
	wire [3-1:0] node178;
	wire [3-1:0] node180;
	wire [3-1:0] node183;
	wire [3-1:0] node184;
	wire [3-1:0] node185;
	wire [3-1:0] node186;
	wire [3-1:0] node188;
	wire [3-1:0] node191;
	wire [3-1:0] node192;
	wire [3-1:0] node195;
	wire [3-1:0] node198;
	wire [3-1:0] node199;
	wire [3-1:0] node200;
	wire [3-1:0] node203;
	wire [3-1:0] node206;
	wire [3-1:0] node207;
	wire [3-1:0] node210;
	wire [3-1:0] node213;
	wire [3-1:0] node214;
	wire [3-1:0] node215;
	wire [3-1:0] node218;
	wire [3-1:0] node219;
	wire [3-1:0] node222;
	wire [3-1:0] node225;
	wire [3-1:0] node226;
	wire [3-1:0] node227;
	wire [3-1:0] node231;
	wire [3-1:0] node232;
	wire [3-1:0] node236;
	wire [3-1:0] node237;
	wire [3-1:0] node238;
	wire [3-1:0] node239;
	wire [3-1:0] node240;
	wire [3-1:0] node241;
	wire [3-1:0] node244;
	wire [3-1:0] node247;
	wire [3-1:0] node249;
	wire [3-1:0] node252;
	wire [3-1:0] node253;
	wire [3-1:0] node254;
	wire [3-1:0] node257;
	wire [3-1:0] node260;
	wire [3-1:0] node261;
	wire [3-1:0] node264;
	wire [3-1:0] node267;
	wire [3-1:0] node268;
	wire [3-1:0] node269;
	wire [3-1:0] node270;
	wire [3-1:0] node273;
	wire [3-1:0] node276;
	wire [3-1:0] node278;
	wire [3-1:0] node281;
	wire [3-1:0] node282;
	wire [3-1:0] node283;
	wire [3-1:0] node286;
	wire [3-1:0] node289;
	wire [3-1:0] node290;
	wire [3-1:0] node293;
	wire [3-1:0] node296;
	wire [3-1:0] node297;
	wire [3-1:0] node299;
	wire [3-1:0] node300;
	wire [3-1:0] node301;
	wire [3-1:0] node304;
	wire [3-1:0] node308;
	wire [3-1:0] node309;
	wire [3-1:0] node310;
	wire [3-1:0] node311;
	wire [3-1:0] node314;
	wire [3-1:0] node318;
	wire [3-1:0] node319;
	wire [3-1:0] node320;
	wire [3-1:0] node323;
	wire [3-1:0] node326;
	wire [3-1:0] node328;
	wire [3-1:0] node331;
	wire [3-1:0] node332;
	wire [3-1:0] node333;
	wire [3-1:0] node334;
	wire [3-1:0] node335;
	wire [3-1:0] node336;
	wire [3-1:0] node337;
	wire [3-1:0] node338;
	wire [3-1:0] node342;
	wire [3-1:0] node344;
	wire [3-1:0] node347;
	wire [3-1:0] node348;
	wire [3-1:0] node350;
	wire [3-1:0] node353;
	wire [3-1:0] node354;
	wire [3-1:0] node357;
	wire [3-1:0] node360;
	wire [3-1:0] node361;
	wire [3-1:0] node362;
	wire [3-1:0] node363;
	wire [3-1:0] node367;
	wire [3-1:0] node368;
	wire [3-1:0] node371;
	wire [3-1:0] node374;
	wire [3-1:0] node375;
	wire [3-1:0] node376;
	wire [3-1:0] node379;
	wire [3-1:0] node382;
	wire [3-1:0] node383;
	wire [3-1:0] node386;
	wire [3-1:0] node389;
	wire [3-1:0] node390;
	wire [3-1:0] node391;
	wire [3-1:0] node392;
	wire [3-1:0] node394;
	wire [3-1:0] node397;
	wire [3-1:0] node399;
	wire [3-1:0] node402;
	wire [3-1:0] node403;
	wire [3-1:0] node404;
	wire [3-1:0] node408;
	wire [3-1:0] node409;
	wire [3-1:0] node412;
	wire [3-1:0] node415;
	wire [3-1:0] node416;
	wire [3-1:0] node417;
	wire [3-1:0] node418;
	wire [3-1:0] node421;
	wire [3-1:0] node424;
	wire [3-1:0] node426;
	wire [3-1:0] node429;
	wire [3-1:0] node430;
	wire [3-1:0] node431;
	wire [3-1:0] node434;
	wire [3-1:0] node437;
	wire [3-1:0] node438;
	wire [3-1:0] node441;
	wire [3-1:0] node444;
	wire [3-1:0] node445;
	wire [3-1:0] node446;
	wire [3-1:0] node447;
	wire [3-1:0] node448;
	wire [3-1:0] node449;
	wire [3-1:0] node452;
	wire [3-1:0] node455;
	wire [3-1:0] node456;
	wire [3-1:0] node460;
	wire [3-1:0] node461;
	wire [3-1:0] node462;
	wire [3-1:0] node465;
	wire [3-1:0] node468;
	wire [3-1:0] node469;
	wire [3-1:0] node472;
	wire [3-1:0] node475;
	wire [3-1:0] node476;
	wire [3-1:0] node477;
	wire [3-1:0] node480;
	wire [3-1:0] node481;
	wire [3-1:0] node485;
	wire [3-1:0] node486;
	wire [3-1:0] node487;
	wire [3-1:0] node490;
	wire [3-1:0] node493;
	wire [3-1:0] node496;
	wire [3-1:0] node497;
	wire [3-1:0] node498;
	wire [3-1:0] node499;
	wire [3-1:0] node500;
	wire [3-1:0] node504;
	wire [3-1:0] node505;
	wire [3-1:0] node508;
	wire [3-1:0] node512;
	wire [3-1:0] node513;
	wire [3-1:0] node514;
	wire [3-1:0] node515;
	wire [3-1:0] node519;
	wire [3-1:0] node520;
	wire [3-1:0] node523;
	wire [3-1:0] node526;
	wire [3-1:0] node527;
	wire [3-1:0] node528;
	wire [3-1:0] node531;
	wire [3-1:0] node534;
	wire [3-1:0] node535;
	wire [3-1:0] node538;
	wire [3-1:0] node541;
	wire [3-1:0] node542;
	wire [3-1:0] node543;
	wire [3-1:0] node544;
	wire [3-1:0] node545;
	wire [3-1:0] node546;
	wire [3-1:0] node549;
	wire [3-1:0] node551;
	wire [3-1:0] node554;
	wire [3-1:0] node555;
	wire [3-1:0] node556;
	wire [3-1:0] node559;
	wire [3-1:0] node562;
	wire [3-1:0] node565;
	wire [3-1:0] node566;
	wire [3-1:0] node567;
	wire [3-1:0] node568;
	wire [3-1:0] node571;
	wire [3-1:0] node574;
	wire [3-1:0] node575;
	wire [3-1:0] node579;
	wire [3-1:0] node581;
	wire [3-1:0] node582;
	wire [3-1:0] node585;
	wire [3-1:0] node588;
	wire [3-1:0] node589;
	wire [3-1:0] node590;
	wire [3-1:0] node591;
	wire [3-1:0] node592;
	wire [3-1:0] node595;
	wire [3-1:0] node599;
	wire [3-1:0] node600;
	wire [3-1:0] node603;
	wire [3-1:0] node605;
	wire [3-1:0] node608;
	wire [3-1:0] node609;
	wire [3-1:0] node610;
	wire [3-1:0] node612;
	wire [3-1:0] node615;
	wire [3-1:0] node616;
	wire [3-1:0] node619;
	wire [3-1:0] node622;
	wire [3-1:0] node623;
	wire [3-1:0] node624;
	wire [3-1:0] node627;
	wire [3-1:0] node630;
	wire [3-1:0] node632;
	wire [3-1:0] node635;
	wire [3-1:0] node636;
	wire [3-1:0] node637;
	wire [3-1:0] node638;
	wire [3-1:0] node639;
	wire [3-1:0] node640;
	wire [3-1:0] node644;
	wire [3-1:0] node645;
	wire [3-1:0] node648;
	wire [3-1:0] node651;
	wire [3-1:0] node652;
	wire [3-1:0] node653;
	wire [3-1:0] node657;
	wire [3-1:0] node659;
	wire [3-1:0] node662;
	wire [3-1:0] node663;
	wire [3-1:0] node664;
	wire [3-1:0] node665;
	wire [3-1:0] node668;
	wire [3-1:0] node671;
	wire [3-1:0] node672;
	wire [3-1:0] node676;
	wire [3-1:0] node677;
	wire [3-1:0] node678;
	wire [3-1:0] node681;
	wire [3-1:0] node684;
	wire [3-1:0] node685;
	wire [3-1:0] node689;
	wire [3-1:0] node690;
	wire [3-1:0] node691;
	wire [3-1:0] node692;
	wire [3-1:0] node693;
	wire [3-1:0] node696;
	wire [3-1:0] node699;
	wire [3-1:0] node700;
	wire [3-1:0] node703;
	wire [3-1:0] node706;
	wire [3-1:0] node707;
	wire [3-1:0] node708;
	wire [3-1:0] node711;
	wire [3-1:0] node714;
	wire [3-1:0] node715;
	wire [3-1:0] node718;
	wire [3-1:0] node721;
	wire [3-1:0] node722;
	wire [3-1:0] node723;
	wire [3-1:0] node725;
	wire [3-1:0] node728;
	wire [3-1:0] node730;
	wire [3-1:0] node733;
	wire [3-1:0] node734;
	wire [3-1:0] node735;
	wire [3-1:0] node739;
	wire [3-1:0] node741;
	wire [3-1:0] node744;
	wire [3-1:0] node745;
	wire [3-1:0] node746;
	wire [3-1:0] node747;
	wire [3-1:0] node748;
	wire [3-1:0] node749;
	wire [3-1:0] node750;
	wire [3-1:0] node751;
	wire [3-1:0] node752;
	wire [3-1:0] node755;
	wire [3-1:0] node759;
	wire [3-1:0] node760;
	wire [3-1:0] node761;
	wire [3-1:0] node764;
	wire [3-1:0] node767;
	wire [3-1:0] node768;
	wire [3-1:0] node771;
	wire [3-1:0] node774;
	wire [3-1:0] node775;
	wire [3-1:0] node776;
	wire [3-1:0] node777;
	wire [3-1:0] node781;
	wire [3-1:0] node783;
	wire [3-1:0] node786;
	wire [3-1:0] node787;
	wire [3-1:0] node789;
	wire [3-1:0] node792;
	wire [3-1:0] node793;
	wire [3-1:0] node796;
	wire [3-1:0] node799;
	wire [3-1:0] node800;
	wire [3-1:0] node801;
	wire [3-1:0] node802;
	wire [3-1:0] node804;
	wire [3-1:0] node807;
	wire [3-1:0] node809;
	wire [3-1:0] node812;
	wire [3-1:0] node813;
	wire [3-1:0] node814;
	wire [3-1:0] node817;
	wire [3-1:0] node820;
	wire [3-1:0] node821;
	wire [3-1:0] node825;
	wire [3-1:0] node826;
	wire [3-1:0] node827;
	wire [3-1:0] node829;
	wire [3-1:0] node832;
	wire [3-1:0] node834;
	wire [3-1:0] node837;
	wire [3-1:0] node838;
	wire [3-1:0] node839;
	wire [3-1:0] node843;
	wire [3-1:0] node844;
	wire [3-1:0] node847;
	wire [3-1:0] node850;
	wire [3-1:0] node851;
	wire [3-1:0] node852;
	wire [3-1:0] node853;
	wire [3-1:0] node855;
	wire [3-1:0] node856;
	wire [3-1:0] node859;
	wire [3-1:0] node862;
	wire [3-1:0] node863;
	wire [3-1:0] node865;
	wire [3-1:0] node868;
	wire [3-1:0] node869;
	wire [3-1:0] node872;
	wire [3-1:0] node875;
	wire [3-1:0] node876;
	wire [3-1:0] node877;
	wire [3-1:0] node878;
	wire [3-1:0] node881;
	wire [3-1:0] node884;
	wire [3-1:0] node885;
	wire [3-1:0] node888;
	wire [3-1:0] node891;
	wire [3-1:0] node892;
	wire [3-1:0] node893;
	wire [3-1:0] node896;
	wire [3-1:0] node899;
	wire [3-1:0] node900;
	wire [3-1:0] node903;
	wire [3-1:0] node906;
	wire [3-1:0] node907;
	wire [3-1:0] node908;
	wire [3-1:0] node909;
	wire [3-1:0] node911;
	wire [3-1:0] node914;
	wire [3-1:0] node916;
	wire [3-1:0] node919;
	wire [3-1:0] node920;
	wire [3-1:0] node922;
	wire [3-1:0] node925;
	wire [3-1:0] node926;
	wire [3-1:0] node930;
	wire [3-1:0] node931;
	wire [3-1:0] node932;
	wire [3-1:0] node933;
	wire [3-1:0] node936;
	wire [3-1:0] node939;
	wire [3-1:0] node940;
	wire [3-1:0] node943;
	wire [3-1:0] node946;
	wire [3-1:0] node947;
	wire [3-1:0] node949;
	wire [3-1:0] node952;
	wire [3-1:0] node953;
	wire [3-1:0] node956;
	wire [3-1:0] node959;
	wire [3-1:0] node960;
	wire [3-1:0] node961;
	wire [3-1:0] node962;
	wire [3-1:0] node964;
	wire [3-1:0] node965;
	wire [3-1:0] node968;
	wire [3-1:0] node970;
	wire [3-1:0] node974;
	wire [3-1:0] node975;
	wire [3-1:0] node976;
	wire [3-1:0] node977;
	wire [3-1:0] node980;
	wire [3-1:0] node981;
	wire [3-1:0] node985;
	wire [3-1:0] node986;
	wire [3-1:0] node987;
	wire [3-1:0] node990;
	wire [3-1:0] node993;
	wire [3-1:0] node995;
	wire [3-1:0] node998;
	wire [3-1:0] node999;
	wire [3-1:0] node1001;
	wire [3-1:0] node1003;
	wire [3-1:0] node1006;
	wire [3-1:0] node1008;
	wire [3-1:0] node1010;
	wire [3-1:0] node1013;
	wire [3-1:0] node1014;
	wire [3-1:0] node1015;
	wire [3-1:0] node1016;
	wire [3-1:0] node1017;
	wire [3-1:0] node1018;
	wire [3-1:0] node1022;
	wire [3-1:0] node1023;
	wire [3-1:0] node1027;
	wire [3-1:0] node1028;
	wire [3-1:0] node1029;
	wire [3-1:0] node1032;
	wire [3-1:0] node1035;
	wire [3-1:0] node1036;
	wire [3-1:0] node1040;
	wire [3-1:0] node1042;
	wire [3-1:0] node1043;
	wire [3-1:0] node1045;
	wire [3-1:0] node1048;
	wire [3-1:0] node1049;
	wire [3-1:0] node1052;
	wire [3-1:0] node1055;
	wire [3-1:0] node1056;
	wire [3-1:0] node1057;
	wire [3-1:0] node1058;
	wire [3-1:0] node1060;
	wire [3-1:0] node1063;
	wire [3-1:0] node1064;
	wire [3-1:0] node1067;
	wire [3-1:0] node1070;
	wire [3-1:0] node1071;
	wire [3-1:0] node1072;
	wire [3-1:0] node1075;
	wire [3-1:0] node1078;
	wire [3-1:0] node1079;
	wire [3-1:0] node1082;
	wire [3-1:0] node1085;
	wire [3-1:0] node1086;
	wire [3-1:0] node1087;
	wire [3-1:0] node1088;
	wire [3-1:0] node1091;
	wire [3-1:0] node1094;
	wire [3-1:0] node1095;
	wire [3-1:0] node1099;
	wire [3-1:0] node1100;
	wire [3-1:0] node1102;
	wire [3-1:0] node1105;
	wire [3-1:0] node1106;
	wire [3-1:0] node1109;
	wire [3-1:0] node1112;
	wire [3-1:0] node1113;
	wire [3-1:0] node1114;
	wire [3-1:0] node1115;
	wire [3-1:0] node1117;
	wire [3-1:0] node1119;
	wire [3-1:0] node1120;
	wire [3-1:0] node1121;
	wire [3-1:0] node1124;
	wire [3-1:0] node1127;
	wire [3-1:0] node1128;
	wire [3-1:0] node1132;
	wire [3-1:0] node1133;
	wire [3-1:0] node1134;
	wire [3-1:0] node1135;
	wire [3-1:0] node1136;
	wire [3-1:0] node1139;
	wire [3-1:0] node1142;
	wire [3-1:0] node1143;
	wire [3-1:0] node1147;
	wire [3-1:0] node1148;
	wire [3-1:0] node1150;
	wire [3-1:0] node1154;
	wire [3-1:0] node1155;
	wire [3-1:0] node1156;
	wire [3-1:0] node1157;
	wire [3-1:0] node1160;
	wire [3-1:0] node1163;
	wire [3-1:0] node1165;
	wire [3-1:0] node1168;
	wire [3-1:0] node1170;
	wire [3-1:0] node1172;
	wire [3-1:0] node1175;
	wire [3-1:0] node1176;
	wire [3-1:0] node1177;
	wire [3-1:0] node1178;
	wire [3-1:0] node1179;
	wire [3-1:0] node1180;
	wire [3-1:0] node1183;
	wire [3-1:0] node1186;
	wire [3-1:0] node1187;
	wire [3-1:0] node1191;
	wire [3-1:0] node1192;
	wire [3-1:0] node1193;
	wire [3-1:0] node1197;
	wire [3-1:0] node1198;
	wire [3-1:0] node1202;
	wire [3-1:0] node1203;
	wire [3-1:0] node1204;
	wire [3-1:0] node1205;
	wire [3-1:0] node1208;
	wire [3-1:0] node1211;
	wire [3-1:0] node1212;
	wire [3-1:0] node1216;
	wire [3-1:0] node1218;
	wire [3-1:0] node1221;
	wire [3-1:0] node1222;
	wire [3-1:0] node1223;
	wire [3-1:0] node1224;
	wire [3-1:0] node1225;
	wire [3-1:0] node1228;
	wire [3-1:0] node1231;
	wire [3-1:0] node1233;
	wire [3-1:0] node1236;
	wire [3-1:0] node1237;
	wire [3-1:0] node1238;
	wire [3-1:0] node1241;
	wire [3-1:0] node1244;
	wire [3-1:0] node1245;
	wire [3-1:0] node1248;
	wire [3-1:0] node1251;
	wire [3-1:0] node1252;
	wire [3-1:0] node1253;
	wire [3-1:0] node1254;
	wire [3-1:0] node1257;
	wire [3-1:0] node1260;
	wire [3-1:0] node1261;
	wire [3-1:0] node1265;
	wire [3-1:0] node1266;
	wire [3-1:0] node1268;
	wire [3-1:0] node1271;
	wire [3-1:0] node1272;
	wire [3-1:0] node1275;
	wire [3-1:0] node1278;
	wire [3-1:0] node1279;
	wire [3-1:0] node1281;
	wire [3-1:0] node1283;
	wire [3-1:0] node1284;
	wire [3-1:0] node1285;
	wire [3-1:0] node1287;
	wire [3-1:0] node1292;
	wire [3-1:0] node1293;
	wire [3-1:0] node1295;
	wire [3-1:0] node1296;
	wire [3-1:0] node1298;
	wire [3-1:0] node1299;
	wire [3-1:0] node1304;
	wire [3-1:0] node1305;
	wire [3-1:0] node1306;
	wire [3-1:0] node1307;
	wire [3-1:0] node1308;
	wire [3-1:0] node1312;
	wire [3-1:0] node1313;
	wire [3-1:0] node1317;
	wire [3-1:0] node1319;
	wire [3-1:0] node1320;
	wire [3-1:0] node1324;
	wire [3-1:0] node1326;
	wire [3-1:0] node1328;

	assign outp = (inp[3]) ? node744 : node1;
		assign node1 = (inp[9]) ? node331 : node2;
			assign node2 = (inp[4]) ? node132 : node3;
				assign node3 = (inp[0]) ? node91 : node4;
					assign node4 = (inp[6]) ? node62 : node5;
						assign node5 = (inp[10]) ? node35 : node6;
							assign node6 = (inp[5]) ? node20 : node7;
								assign node7 = (inp[1]) ? node15 : node8;
									assign node8 = (inp[7]) ? node12 : node9;
										assign node9 = (inp[11]) ? 3'b011 : 3'b011;
										assign node12 = (inp[11]) ? 3'b011 : 3'b111;
									assign node15 = (inp[7]) ? 3'b111 : node16;
										assign node16 = (inp[2]) ? 3'b111 : 3'b011;
								assign node20 = (inp[7]) ? node28 : node21;
									assign node21 = (inp[2]) ? node25 : node22;
										assign node22 = (inp[11]) ? 3'b001 : 3'b101;
										assign node25 = (inp[8]) ? 3'b011 : 3'b101;
									assign node28 = (inp[2]) ? node32 : node29;
										assign node29 = (inp[11]) ? 3'b101 : 3'b011;
										assign node32 = (inp[11]) ? 3'b011 : 3'b011;
							assign node35 = (inp[2]) ? node51 : node36;
								assign node36 = (inp[7]) ? node44 : node37;
									assign node37 = (inp[1]) ? node41 : node38;
										assign node38 = (inp[8]) ? 3'b001 : 3'b000;
										assign node41 = (inp[5]) ? 3'b001 : 3'b101;
									assign node44 = (inp[1]) ? node48 : node45;
										assign node45 = (inp[5]) ? 3'b001 : 3'b101;
										assign node48 = (inp[5]) ? 3'b101 : 3'b011;
								assign node51 = (inp[1]) ? node57 : node52;
									assign node52 = (inp[11]) ? node54 : 3'b101;
										assign node54 = (inp[8]) ? 3'b001 : 3'b001;
									assign node57 = (inp[7]) ? node59 : 3'b101;
										assign node59 = (inp[11]) ? 3'b101 : 3'b111;
						assign node62 = (inp[5]) ? node72 : node63;
							assign node63 = (inp[7]) ? 3'b111 : node64;
								assign node64 = (inp[11]) ? node66 : 3'b111;
									assign node66 = (inp[8]) ? 3'b111 : node67;
										assign node67 = (inp[10]) ? 3'b011 : 3'b111;
							assign node72 = (inp[1]) ? node84 : node73;
								assign node73 = (inp[10]) ? node79 : node74;
									assign node74 = (inp[7]) ? 3'b111 : node75;
										assign node75 = (inp[11]) ? 3'b011 : 3'b111;
									assign node79 = (inp[11]) ? node81 : 3'b011;
										assign node81 = (inp[7]) ? 3'b011 : 3'b101;
								assign node84 = (inp[10]) ? node86 : 3'b111;
									assign node86 = (inp[7]) ? 3'b111 : node87;
										assign node87 = (inp[8]) ? 3'b011 : 3'b001;
					assign node91 = (inp[6]) ? node121 : node92;
						assign node92 = (inp[10]) ? node102 : node93;
							assign node93 = (inp[5]) ? node95 : 3'b111;
								assign node95 = (inp[1]) ? 3'b111 : node96;
									assign node96 = (inp[7]) ? 3'b111 : node97;
										assign node97 = (inp[2]) ? 3'b111 : 3'b011;
							assign node102 = (inp[5]) ? node110 : node103;
								assign node103 = (inp[1]) ? 3'b111 : node104;
									assign node104 = (inp[8]) ? 3'b111 : node105;
										assign node105 = (inp[11]) ? 3'b011 : 3'b011;
								assign node110 = (inp[2]) ? node116 : node111;
									assign node111 = (inp[7]) ? 3'b011 : node112;
										assign node112 = (inp[8]) ? 3'b011 : 3'b101;
									assign node116 = (inp[8]) ? 3'b111 : node117;
										assign node117 = (inp[1]) ? 3'b011 : 3'b001;
						assign node121 = (inp[7]) ? 3'b111 : node122;
							assign node122 = (inp[8]) ? 3'b111 : node123;
								assign node123 = (inp[10]) ? node125 : 3'b111;
									assign node125 = (inp[11]) ? node127 : 3'b111;
										assign node127 = (inp[2]) ? 3'b111 : 3'b011;
				assign node132 = (inp[6]) ? node236 : node133;
					assign node133 = (inp[7]) ? node183 : node134;
						assign node134 = (inp[0]) ? node158 : node135;
							assign node135 = (inp[10]) ? node145 : node136;
								assign node136 = (inp[5]) ? 3'b110 : node137;
									assign node137 = (inp[1]) ? node141 : node138;
										assign node138 = (inp[11]) ? 3'b110 : 3'b001;
										assign node141 = (inp[8]) ? 3'b101 : 3'b001;
								assign node145 = (inp[5]) ? node151 : node146;
									assign node146 = (inp[1]) ? 3'b110 : node147;
										assign node147 = (inp[11]) ? 3'b010 : 3'b110;
									assign node151 = (inp[2]) ? node155 : node152;
										assign node152 = (inp[1]) ? 3'b010 : 3'b000;
										assign node155 = (inp[1]) ? 3'b010 : 3'b010;
							assign node158 = (inp[5]) ? node170 : node159;
								assign node159 = (inp[1]) ? node165 : node160;
									assign node160 = (inp[10]) ? node162 : 3'b101;
										assign node162 = (inp[8]) ? 3'b001 : 3'b000;
									assign node165 = (inp[10]) ? node167 : 3'b011;
										assign node167 = (inp[2]) ? 3'b001 : 3'b101;
								assign node170 = (inp[10]) ? node178 : node171;
									assign node171 = (inp[8]) ? node175 : node172;
										assign node172 = (inp[11]) ? 3'b001 : 3'b101;
										assign node175 = (inp[11]) ? 3'b101 : 3'b001;
									assign node178 = (inp[1]) ? node180 : 3'b110;
										assign node180 = (inp[11]) ? 3'b110 : 3'b001;
						assign node183 = (inp[10]) ? node213 : node184;
							assign node184 = (inp[5]) ? node198 : node185;
								assign node185 = (inp[0]) ? node191 : node186;
									assign node186 = (inp[8]) ? node188 : 3'b101;
										assign node188 = (inp[11]) ? 3'b001 : 3'b011;
									assign node191 = (inp[8]) ? node195 : node192;
										assign node192 = (inp[11]) ? 3'b011 : 3'b011;
										assign node195 = (inp[1]) ? 3'b111 : 3'b011;
								assign node198 = (inp[1]) ? node206 : node199;
									assign node199 = (inp[8]) ? node203 : node200;
										assign node200 = (inp[11]) ? 3'b001 : 3'b101;
										assign node203 = (inp[0]) ? 3'b011 : 3'b110;
									assign node206 = (inp[0]) ? node210 : node207;
										assign node207 = (inp[11]) ? 3'b001 : 3'b101;
										assign node210 = (inp[11]) ? 3'b101 : 3'b011;
							assign node213 = (inp[0]) ? node225 : node214;
								assign node214 = (inp[8]) ? node218 : node215;
									assign node215 = (inp[2]) ? 3'b110 : 3'b010;
									assign node218 = (inp[5]) ? node222 : node219;
										assign node219 = (inp[2]) ? 3'b001 : 3'b001;
										assign node222 = (inp[2]) ? 3'b000 : 3'b110;
								assign node225 = (inp[5]) ? node231 : node226;
									assign node226 = (inp[11]) ? 3'b101 : node227;
										assign node227 = (inp[1]) ? 3'b011 : 3'b101;
									assign node231 = (inp[11]) ? 3'b001 : node232;
										assign node232 = (inp[1]) ? 3'b101 : 3'b001;
					assign node236 = (inp[0]) ? node296 : node237;
						assign node237 = (inp[10]) ? node267 : node238;
							assign node238 = (inp[5]) ? node252 : node239;
								assign node239 = (inp[1]) ? node247 : node240;
									assign node240 = (inp[11]) ? node244 : node241;
										assign node241 = (inp[8]) ? 3'b011 : 3'b011;
										assign node244 = (inp[7]) ? 3'b011 : 3'b101;
									assign node247 = (inp[11]) ? node249 : 3'b111;
										assign node249 = (inp[8]) ? 3'b011 : 3'b111;
								assign node252 = (inp[1]) ? node260 : node253;
									assign node253 = (inp[2]) ? node257 : node254;
										assign node254 = (inp[8]) ? 3'b101 : 3'b001;
										assign node257 = (inp[8]) ? 3'b101 : 3'b101;
									assign node260 = (inp[7]) ? node264 : node261;
										assign node261 = (inp[11]) ? 3'b001 : 3'b101;
										assign node264 = (inp[2]) ? 3'b011 : 3'b011;
							assign node267 = (inp[2]) ? node281 : node268;
								assign node268 = (inp[8]) ? node276 : node269;
									assign node269 = (inp[5]) ? node273 : node270;
										assign node270 = (inp[11]) ? 3'b001 : 3'b011;
										assign node273 = (inp[11]) ? 3'b110 : 3'b001;
									assign node276 = (inp[7]) ? node278 : 3'b001;
										assign node278 = (inp[5]) ? 3'b001 : 3'b101;
								assign node281 = (inp[1]) ? node289 : node282;
									assign node282 = (inp[5]) ? node286 : node283;
										assign node283 = (inp[11]) ? 3'b001 : 3'b101;
										assign node286 = (inp[7]) ? 3'b101 : 3'b110;
									assign node289 = (inp[5]) ? node293 : node290;
										assign node290 = (inp[7]) ? 3'b011 : 3'b101;
										assign node293 = (inp[7]) ? 3'b101 : 3'b001;
						assign node296 = (inp[5]) ? node308 : node297;
							assign node297 = (inp[10]) ? node299 : 3'b111;
								assign node299 = (inp[7]) ? 3'b111 : node300;
									assign node300 = (inp[1]) ? node304 : node301;
										assign node301 = (inp[11]) ? 3'b101 : 3'b011;
										assign node304 = (inp[8]) ? 3'b111 : 3'b011;
							assign node308 = (inp[10]) ? node318 : node309;
								assign node309 = (inp[1]) ? 3'b111 : node310;
									assign node310 = (inp[7]) ? node314 : node311;
										assign node311 = (inp[11]) ? 3'b001 : 3'b011;
										assign node314 = (inp[11]) ? 3'b011 : 3'b111;
								assign node318 = (inp[7]) ? node326 : node319;
									assign node319 = (inp[8]) ? node323 : node320;
										assign node320 = (inp[1]) ? 3'b101 : 3'b001;
										assign node323 = (inp[1]) ? 3'b011 : 3'b101;
									assign node326 = (inp[8]) ? node328 : 3'b011;
										assign node328 = (inp[11]) ? 3'b101 : 3'b011;
			assign node331 = (inp[4]) ? node541 : node332;
				assign node332 = (inp[0]) ? node444 : node333;
					assign node333 = (inp[6]) ? node389 : node334;
						assign node334 = (inp[10]) ? node360 : node335;
							assign node335 = (inp[5]) ? node347 : node336;
								assign node336 = (inp[7]) ? node342 : node337;
									assign node337 = (inp[8]) ? 3'b001 : node338;
										assign node338 = (inp[1]) ? 3'b001 : 3'b110;
									assign node342 = (inp[11]) ? node344 : 3'b101;
										assign node344 = (inp[1]) ? 3'b101 : 3'b001;
								assign node347 = (inp[1]) ? node353 : node348;
									assign node348 = (inp[8]) ? node350 : 3'b110;
										assign node350 = (inp[7]) ? 3'b001 : 3'b110;
									assign node353 = (inp[7]) ? node357 : node354;
										assign node354 = (inp[11]) ? 3'b110 : 3'b001;
										assign node357 = (inp[8]) ? 3'b001 : 3'b001;
							assign node360 = (inp[11]) ? node374 : node361;
								assign node361 = (inp[8]) ? node367 : node362;
									assign node362 = (inp[7]) ? 3'b110 : node363;
										assign node363 = (inp[2]) ? 3'b010 : 3'b110;
									assign node367 = (inp[5]) ? node371 : node368;
										assign node368 = (inp[7]) ? 3'b001 : 3'b000;
										assign node371 = (inp[1]) ? 3'b000 : 3'b110;
								assign node374 = (inp[5]) ? node382 : node375;
									assign node375 = (inp[7]) ? node379 : node376;
										assign node376 = (inp[1]) ? 3'b110 : 3'b010;
										assign node379 = (inp[1]) ? 3'b001 : 3'b110;
									assign node382 = (inp[2]) ? node386 : node383;
										assign node383 = (inp[1]) ? 3'b010 : 3'b100;
										assign node386 = (inp[1]) ? 3'b110 : 3'b010;
						assign node389 = (inp[10]) ? node415 : node390;
							assign node390 = (inp[7]) ? node402 : node391;
								assign node391 = (inp[2]) ? node397 : node392;
									assign node392 = (inp[5]) ? node394 : 3'b011;
										assign node394 = (inp[1]) ? 3'b101 : 3'b001;
									assign node397 = (inp[5]) ? node399 : 3'b101;
										assign node399 = (inp[1]) ? 3'b101 : 3'b001;
								assign node402 = (inp[5]) ? node408 : node403;
									assign node403 = (inp[1]) ? 3'b111 : node404;
										assign node404 = (inp[2]) ? 3'b011 : 3'b011;
									assign node408 = (inp[1]) ? node412 : node409;
										assign node409 = (inp[11]) ? 3'b101 : 3'b001;
										assign node412 = (inp[8]) ? 3'b011 : 3'b001;
							assign node415 = (inp[5]) ? node429 : node416;
								assign node416 = (inp[1]) ? node424 : node417;
									assign node417 = (inp[7]) ? node421 : node418;
										assign node418 = (inp[11]) ? 3'b001 : 3'b001;
										assign node421 = (inp[2]) ? 3'b011 : 3'b101;
									assign node424 = (inp[8]) ? node426 : 3'b101;
										assign node426 = (inp[7]) ? 3'b011 : 3'b101;
								assign node429 = (inp[7]) ? node437 : node430;
									assign node430 = (inp[1]) ? node434 : node431;
										assign node431 = (inp[8]) ? 3'b110 : 3'b010;
										assign node434 = (inp[8]) ? 3'b001 : 3'b001;
									assign node437 = (inp[1]) ? node441 : node438;
										assign node438 = (inp[8]) ? 3'b001 : 3'b001;
										assign node441 = (inp[11]) ? 3'b001 : 3'b101;
					assign node444 = (inp[6]) ? node496 : node445;
						assign node445 = (inp[10]) ? node475 : node446;
							assign node446 = (inp[5]) ? node460 : node447;
								assign node447 = (inp[1]) ? node455 : node448;
									assign node448 = (inp[7]) ? node452 : node449;
										assign node449 = (inp[11]) ? 3'b001 : 3'b101;
										assign node452 = (inp[11]) ? 3'b101 : 3'b011;
									assign node455 = (inp[11]) ? 3'b011 : node456;
										assign node456 = (inp[7]) ? 3'b111 : 3'b011;
								assign node460 = (inp[8]) ? node468 : node461;
									assign node461 = (inp[11]) ? node465 : node462;
										assign node462 = (inp[1]) ? 3'b011 : 3'b001;
										assign node465 = (inp[2]) ? 3'b101 : 3'b001;
									assign node468 = (inp[7]) ? node472 : node469;
										assign node469 = (inp[1]) ? 3'b101 : 3'b001;
										assign node472 = (inp[1]) ? 3'b011 : 3'b101;
							assign node475 = (inp[5]) ? node485 : node476;
								assign node476 = (inp[7]) ? node480 : node477;
									assign node477 = (inp[11]) ? 3'b001 : 3'b101;
									assign node480 = (inp[8]) ? 3'b101 : node481;
										assign node481 = (inp[11]) ? 3'b101 : 3'b001;
								assign node485 = (inp[1]) ? node493 : node486;
									assign node486 = (inp[7]) ? node490 : node487;
										assign node487 = (inp[2]) ? 3'b000 : 3'b110;
										assign node490 = (inp[8]) ? 3'b001 : 3'b000;
									assign node493 = (inp[7]) ? 3'b101 : 3'b001;
						assign node496 = (inp[10]) ? node512 : node497;
							assign node497 = (inp[7]) ? 3'b111 : node498;
								assign node498 = (inp[5]) ? node504 : node499;
									assign node499 = (inp[8]) ? 3'b111 : node500;
										assign node500 = (inp[1]) ? 3'b111 : 3'b011;
									assign node504 = (inp[2]) ? node508 : node505;
										assign node505 = (inp[8]) ? 3'b011 : 3'b011;
										assign node508 = (inp[1]) ? 3'b111 : 3'b001;
							assign node512 = (inp[5]) ? node526 : node513;
								assign node513 = (inp[11]) ? node519 : node514;
									assign node514 = (inp[7]) ? 3'b111 : node515;
										assign node515 = (inp[2]) ? 3'b111 : 3'b011;
									assign node519 = (inp[8]) ? node523 : node520;
										assign node520 = (inp[1]) ? 3'b011 : 3'b001;
										assign node523 = (inp[1]) ? 3'b111 : 3'b011;
								assign node526 = (inp[1]) ? node534 : node527;
									assign node527 = (inp[7]) ? node531 : node528;
										assign node528 = (inp[11]) ? 3'b001 : 3'b101;
										assign node531 = (inp[11]) ? 3'b101 : 3'b011;
									assign node534 = (inp[7]) ? node538 : node535;
										assign node535 = (inp[2]) ? 3'b011 : 3'b101;
										assign node538 = (inp[11]) ? 3'b011 : 3'b011;
				assign node541 = (inp[6]) ? node635 : node542;
					assign node542 = (inp[0]) ? node588 : node543;
						assign node543 = (inp[5]) ? node565 : node544;
							assign node544 = (inp[10]) ? node554 : node545;
								assign node545 = (inp[11]) ? node549 : node546;
									assign node546 = (inp[1]) ? 3'b110 : 3'b010;
									assign node549 = (inp[8]) ? node551 : 3'b010;
										assign node551 = (inp[2]) ? 3'b010 : 3'b010;
								assign node554 = (inp[7]) ? node562 : node555;
									assign node555 = (inp[2]) ? node559 : node556;
										assign node556 = (inp[11]) ? 3'b000 : 3'b100;
										assign node559 = (inp[11]) ? 3'b100 : 3'b000;
									assign node562 = (inp[1]) ? 3'b010 : 3'b100;
							assign node565 = (inp[10]) ? node579 : node566;
								assign node566 = (inp[7]) ? node574 : node567;
									assign node567 = (inp[1]) ? node571 : node568;
										assign node568 = (inp[8]) ? 3'b100 : 3'b000;
										assign node571 = (inp[8]) ? 3'b100 : 3'b100;
									assign node574 = (inp[1]) ? 3'b010 : node575;
										assign node575 = (inp[11]) ? 3'b100 : 3'b010;
								assign node579 = (inp[1]) ? node581 : 3'b000;
									assign node581 = (inp[7]) ? node585 : node582;
										assign node582 = (inp[8]) ? 3'b000 : 3'b000;
										assign node585 = (inp[11]) ? 3'b100 : 3'b100;
						assign node588 = (inp[10]) ? node608 : node589;
							assign node589 = (inp[1]) ? node599 : node590;
								assign node590 = (inp[8]) ? 3'b110 : node591;
									assign node591 = (inp[7]) ? node595 : node592;
										assign node592 = (inp[5]) ? 3'b000 : 3'b110;
										assign node595 = (inp[2]) ? 3'b001 : 3'b010;
								assign node599 = (inp[11]) ? node603 : node600;
									assign node600 = (inp[2]) ? 3'b101 : 3'b001;
									assign node603 = (inp[2]) ? node605 : 3'b110;
										assign node605 = (inp[8]) ? 3'b001 : 3'b001;
							assign node608 = (inp[5]) ? node622 : node609;
								assign node609 = (inp[1]) ? node615 : node610;
									assign node610 = (inp[2]) ? node612 : 3'b010;
										assign node612 = (inp[7]) ? 3'b110 : 3'b010;
									assign node615 = (inp[7]) ? node619 : node616;
										assign node616 = (inp[11]) ? 3'b010 : 3'b110;
										assign node619 = (inp[2]) ? 3'b001 : 3'b110;
								assign node622 = (inp[7]) ? node630 : node623;
									assign node623 = (inp[2]) ? node627 : node624;
										assign node624 = (inp[1]) ? 3'b100 : 3'b000;
										assign node627 = (inp[8]) ? 3'b010 : 3'b100;
									assign node630 = (inp[8]) ? node632 : 3'b010;
										assign node632 = (inp[1]) ? 3'b110 : 3'b010;
					assign node635 = (inp[0]) ? node689 : node636;
						assign node636 = (inp[5]) ? node662 : node637;
							assign node637 = (inp[10]) ? node651 : node638;
								assign node638 = (inp[7]) ? node644 : node639;
									assign node639 = (inp[1]) ? 3'b001 : node640;
										assign node640 = (inp[2]) ? 3'b001 : 3'b110;
									assign node644 = (inp[1]) ? node648 : node645;
										assign node645 = (inp[11]) ? 3'b000 : 3'b001;
										assign node648 = (inp[11]) ? 3'b001 : 3'b101;
								assign node651 = (inp[7]) ? node657 : node652;
									assign node652 = (inp[1]) ? 3'b110 : node653;
										assign node653 = (inp[8]) ? 3'b010 : 3'b010;
									assign node657 = (inp[1]) ? node659 : 3'b110;
										assign node659 = (inp[11]) ? 3'b000 : 3'b001;
							assign node662 = (inp[10]) ? node676 : node663;
								assign node663 = (inp[1]) ? node671 : node664;
									assign node664 = (inp[8]) ? node668 : node665;
										assign node665 = (inp[7]) ? 3'b010 : 3'b010;
										assign node668 = (inp[2]) ? 3'b110 : 3'b010;
									assign node671 = (inp[2]) ? 3'b001 : node672;
										assign node672 = (inp[11]) ? 3'b110 : 3'b001;
								assign node676 = (inp[7]) ? node684 : node677;
									assign node677 = (inp[8]) ? node681 : node678;
										assign node678 = (inp[2]) ? 3'b100 : 3'b000;
										assign node681 = (inp[11]) ? 3'b100 : 3'b010;
									assign node684 = (inp[1]) ? 3'b010 : node685;
										assign node685 = (inp[8]) ? 3'b010 : 3'b100;
						assign node689 = (inp[10]) ? node721 : node690;
							assign node690 = (inp[5]) ? node706 : node691;
								assign node691 = (inp[7]) ? node699 : node692;
									assign node692 = (inp[1]) ? node696 : node693;
										assign node693 = (inp[11]) ? 3'b001 : 3'b101;
										assign node696 = (inp[11]) ? 3'b101 : 3'b011;
									assign node699 = (inp[2]) ? node703 : node700;
										assign node700 = (inp[11]) ? 3'b101 : 3'b111;
										assign node703 = (inp[1]) ? 3'b011 : 3'b011;
								assign node706 = (inp[2]) ? node714 : node707;
									assign node707 = (inp[7]) ? node711 : node708;
										assign node708 = (inp[1]) ? 3'b001 : 3'b110;
										assign node711 = (inp[1]) ? 3'b001 : 3'b001;
									assign node714 = (inp[7]) ? node718 : node715;
										assign node715 = (inp[1]) ? 3'b001 : 3'b001;
										assign node718 = (inp[11]) ? 3'b101 : 3'b101;
							assign node721 = (inp[5]) ? node733 : node722;
								assign node722 = (inp[7]) ? node728 : node723;
									assign node723 = (inp[11]) ? node725 : 3'b001;
										assign node725 = (inp[8]) ? 3'b001 : 3'b110;
									assign node728 = (inp[11]) ? node730 : 3'b101;
										assign node730 = (inp[8]) ? 3'b101 : 3'b001;
								assign node733 = (inp[11]) ? node739 : node734;
									assign node734 = (inp[7]) ? 3'b001 : node735;
										assign node735 = (inp[1]) ? 3'b001 : 3'b110;
									assign node739 = (inp[2]) ? node741 : 3'b110;
										assign node741 = (inp[8]) ? 3'b110 : 3'b000;
		assign node744 = (inp[4]) ? node1112 : node745;
			assign node745 = (inp[9]) ? node959 : node746;
				assign node746 = (inp[6]) ? node850 : node747;
					assign node747 = (inp[0]) ? node799 : node748;
						assign node748 = (inp[5]) ? node774 : node749;
							assign node749 = (inp[7]) ? node759 : node750;
								assign node750 = (inp[10]) ? 3'b100 : node751;
									assign node751 = (inp[1]) ? node755 : node752;
										assign node752 = (inp[2]) ? 3'b010 : 3'b100;
										assign node755 = (inp[11]) ? 3'b010 : 3'b110;
								assign node759 = (inp[10]) ? node767 : node760;
									assign node760 = (inp[1]) ? node764 : node761;
										assign node761 = (inp[8]) ? 3'b110 : 3'b010;
										assign node764 = (inp[8]) ? 3'b000 : 3'b110;
									assign node767 = (inp[1]) ? node771 : node768;
										assign node768 = (inp[11]) ? 3'b100 : 3'b010;
										assign node771 = (inp[2]) ? 3'b010 : 3'b010;
							assign node774 = (inp[10]) ? node786 : node775;
								assign node775 = (inp[7]) ? node781 : node776;
									assign node776 = (inp[11]) ? 3'b000 : node777;
										assign node777 = (inp[8]) ? 3'b100 : 3'b000;
									assign node781 = (inp[11]) ? node783 : 3'b010;
										assign node783 = (inp[1]) ? 3'b010 : 3'b100;
								assign node786 = (inp[7]) ? node792 : node787;
									assign node787 = (inp[2]) ? node789 : 3'b000;
										assign node789 = (inp[1]) ? 3'b000 : 3'b000;
									assign node792 = (inp[1]) ? node796 : node793;
										assign node793 = (inp[8]) ? 3'b000 : 3'b000;
										assign node796 = (inp[8]) ? 3'b000 : 3'b100;
						assign node799 = (inp[7]) ? node825 : node800;
							assign node800 = (inp[10]) ? node812 : node801;
								assign node801 = (inp[5]) ? node807 : node802;
									assign node802 = (inp[1]) ? node804 : 3'b110;
										assign node804 = (inp[11]) ? 3'b000 : 3'b001;
									assign node807 = (inp[11]) ? node809 : 3'b110;
										assign node809 = (inp[2]) ? 3'b010 : 3'b110;
								assign node812 = (inp[5]) ? node820 : node813;
									assign node813 = (inp[11]) ? node817 : node814;
										assign node814 = (inp[1]) ? 3'b110 : 3'b010;
										assign node817 = (inp[2]) ? 3'b010 : 3'b010;
									assign node820 = (inp[11]) ? 3'b100 : node821;
										assign node821 = (inp[1]) ? 3'b010 : 3'b100;
							assign node825 = (inp[10]) ? node837 : node826;
								assign node826 = (inp[5]) ? node832 : node827;
									assign node827 = (inp[1]) ? node829 : 3'b001;
										assign node829 = (inp[2]) ? 3'b101 : 3'b001;
									assign node832 = (inp[1]) ? node834 : 3'b110;
										assign node834 = (inp[11]) ? 3'b000 : 3'b001;
								assign node837 = (inp[5]) ? node843 : node838;
									assign node838 = (inp[11]) ? 3'b110 : node839;
										assign node839 = (inp[1]) ? 3'b001 : 3'b110;
									assign node843 = (inp[11]) ? node847 : node844;
										assign node844 = (inp[1]) ? 3'b110 : 3'b010;
										assign node847 = (inp[1]) ? 3'b010 : 3'b100;
					assign node850 = (inp[0]) ? node906 : node851;
						assign node851 = (inp[5]) ? node875 : node852;
							assign node852 = (inp[10]) ? node862 : node853;
								assign node853 = (inp[7]) ? node855 : 3'b001;
									assign node855 = (inp[1]) ? node859 : node856;
										assign node856 = (inp[2]) ? 3'b001 : 3'b000;
										assign node859 = (inp[2]) ? 3'b101 : 3'b001;
								assign node862 = (inp[11]) ? node868 : node863;
									assign node863 = (inp[1]) ? node865 : 3'b110;
										assign node865 = (inp[7]) ? 3'b001 : 3'b110;
									assign node868 = (inp[1]) ? node872 : node869;
										assign node869 = (inp[7]) ? 3'b110 : 3'b100;
										assign node872 = (inp[8]) ? 3'b110 : 3'b010;
							assign node875 = (inp[8]) ? node891 : node876;
								assign node876 = (inp[7]) ? node884 : node877;
									assign node877 = (inp[10]) ? node881 : node878;
										assign node878 = (inp[1]) ? 3'b010 : 3'b010;
										assign node881 = (inp[11]) ? 3'b100 : 3'b010;
									assign node884 = (inp[10]) ? node888 : node885;
										assign node885 = (inp[2]) ? 3'b110 : 3'b010;
										assign node888 = (inp[2]) ? 3'b010 : 3'b110;
								assign node891 = (inp[10]) ? node899 : node892;
									assign node892 = (inp[11]) ? node896 : node893;
										assign node893 = (inp[1]) ? 3'b001 : 3'b110;
										assign node896 = (inp[7]) ? 3'b110 : 3'b110;
									assign node899 = (inp[7]) ? node903 : node900;
										assign node900 = (inp[2]) ? 3'b010 : 3'b100;
										assign node903 = (inp[2]) ? 3'b110 : 3'b010;
						assign node906 = (inp[7]) ? node930 : node907;
							assign node907 = (inp[10]) ? node919 : node908;
								assign node908 = (inp[1]) ? node914 : node909;
									assign node909 = (inp[5]) ? node911 : 3'b101;
										assign node911 = (inp[11]) ? 3'b000 : 3'b001;
									assign node914 = (inp[5]) ? node916 : 3'b011;
										assign node916 = (inp[2]) ? 3'b101 : 3'b001;
								assign node919 = (inp[5]) ? node925 : node920;
									assign node920 = (inp[1]) ? node922 : 3'b110;
										assign node922 = (inp[8]) ? 3'b101 : 3'b001;
									assign node925 = (inp[1]) ? 3'b110 : node926;
										assign node926 = (inp[8]) ? 3'b110 : 3'b010;
							assign node930 = (inp[10]) ? node946 : node931;
								assign node931 = (inp[5]) ? node939 : node932;
									assign node932 = (inp[11]) ? node936 : node933;
										assign node933 = (inp[1]) ? 3'b111 : 3'b011;
										assign node936 = (inp[1]) ? 3'b011 : 3'b001;
									assign node939 = (inp[1]) ? node943 : node940;
										assign node940 = (inp[11]) ? 3'b001 : 3'b101;
										assign node943 = (inp[2]) ? 3'b001 : 3'b101;
								assign node946 = (inp[8]) ? node952 : node947;
									assign node947 = (inp[1]) ? node949 : 3'b001;
										assign node949 = (inp[5]) ? 3'b001 : 3'b101;
									assign node952 = (inp[5]) ? node956 : node953;
										assign node953 = (inp[1]) ? 3'b001 : 3'b001;
										assign node956 = (inp[1]) ? 3'b001 : 3'b001;
				assign node959 = (inp[0]) ? node1013 : node960;
					assign node960 = (inp[6]) ? node974 : node961;
						assign node961 = (inp[11]) ? 3'b000 : node962;
							assign node962 = (inp[7]) ? node964 : 3'b000;
								assign node964 = (inp[10]) ? node968 : node965;
									assign node965 = (inp[1]) ? 3'b100 : 3'b000;
									assign node968 = (inp[8]) ? node970 : 3'b000;
										assign node970 = (inp[5]) ? 3'b000 : 3'b000;
						assign node974 = (inp[5]) ? node998 : node975;
							assign node975 = (inp[1]) ? node985 : node976;
								assign node976 = (inp[7]) ? node980 : node977;
									assign node977 = (inp[10]) ? 3'b000 : 3'b100;
									assign node980 = (inp[10]) ? 3'b100 : node981;
										assign node981 = (inp[2]) ? 3'b010 : 3'b100;
								assign node985 = (inp[8]) ? node993 : node986;
									assign node986 = (inp[11]) ? node990 : node987;
										assign node987 = (inp[10]) ? 3'b100 : 3'b110;
										assign node990 = (inp[10]) ? 3'b000 : 3'b100;
									assign node993 = (inp[10]) ? node995 : 3'b010;
										assign node995 = (inp[11]) ? 3'b000 : 3'b010;
							assign node998 = (inp[10]) ? node1006 : node999;
								assign node999 = (inp[11]) ? node1001 : 3'b100;
									assign node1001 = (inp[7]) ? node1003 : 3'b000;
										assign node1003 = (inp[8]) ? 3'b000 : 3'b100;
								assign node1006 = (inp[7]) ? node1008 : 3'b000;
									assign node1008 = (inp[1]) ? node1010 : 3'b000;
										assign node1010 = (inp[11]) ? 3'b000 : 3'b100;
					assign node1013 = (inp[6]) ? node1055 : node1014;
						assign node1014 = (inp[5]) ? node1040 : node1015;
							assign node1015 = (inp[7]) ? node1027 : node1016;
								assign node1016 = (inp[2]) ? node1022 : node1017;
									assign node1017 = (inp[10]) ? 3'b000 : node1018;
										assign node1018 = (inp[1]) ? 3'b100 : 3'b000;
									assign node1022 = (inp[11]) ? 3'b100 : node1023;
										assign node1023 = (inp[8]) ? 3'b010 : 3'b100;
								assign node1027 = (inp[10]) ? node1035 : node1028;
									assign node1028 = (inp[8]) ? node1032 : node1029;
										assign node1029 = (inp[1]) ? 3'b010 : 3'b100;
										assign node1032 = (inp[1]) ? 3'b010 : 3'b010;
									assign node1035 = (inp[11]) ? 3'b100 : node1036;
										assign node1036 = (inp[1]) ? 3'b010 : 3'b100;
							assign node1040 = (inp[1]) ? node1042 : 3'b000;
								assign node1042 = (inp[7]) ? node1048 : node1043;
									assign node1043 = (inp[8]) ? node1045 : 3'b000;
										assign node1045 = (inp[11]) ? 3'b000 : 3'b100;
									assign node1048 = (inp[10]) ? node1052 : node1049;
										assign node1049 = (inp[8]) ? 3'b010 : 3'b100;
										assign node1052 = (inp[8]) ? 3'b100 : 3'b000;
						assign node1055 = (inp[5]) ? node1085 : node1056;
							assign node1056 = (inp[7]) ? node1070 : node1057;
								assign node1057 = (inp[8]) ? node1063 : node1058;
									assign node1058 = (inp[11]) ? node1060 : 3'b010;
										assign node1060 = (inp[10]) ? 3'b100 : 3'b010;
									assign node1063 = (inp[10]) ? node1067 : node1064;
										assign node1064 = (inp[11]) ? 3'b110 : 3'b110;
										assign node1067 = (inp[11]) ? 3'b010 : 3'b010;
								assign node1070 = (inp[10]) ? node1078 : node1071;
									assign node1071 = (inp[8]) ? node1075 : node1072;
										assign node1072 = (inp[1]) ? 3'b001 : 3'b110;
										assign node1075 = (inp[1]) ? 3'b001 : 3'b001;
									assign node1078 = (inp[8]) ? node1082 : node1079;
										assign node1079 = (inp[2]) ? 3'b110 : 3'b010;
										assign node1082 = (inp[11]) ? 3'b110 : 3'b110;
							assign node1085 = (inp[7]) ? node1099 : node1086;
								assign node1086 = (inp[10]) ? node1094 : node1087;
									assign node1087 = (inp[1]) ? node1091 : node1088;
										assign node1088 = (inp[8]) ? 3'b010 : 3'b100;
										assign node1091 = (inp[11]) ? 3'b010 : 3'b010;
									assign node1094 = (inp[8]) ? 3'b100 : node1095;
										assign node1095 = (inp[11]) ? 3'b000 : 3'b100;
								assign node1099 = (inp[10]) ? node1105 : node1100;
									assign node1100 = (inp[11]) ? node1102 : 3'b110;
										assign node1102 = (inp[1]) ? 3'b110 : 3'b010;
									assign node1105 = (inp[1]) ? node1109 : node1106;
										assign node1106 = (inp[11]) ? 3'b100 : 3'b010;
										assign node1109 = (inp[8]) ? 3'b010 : 3'b010;
			assign node1112 = (inp[9]) ? node1278 : node1113;
				assign node1113 = (inp[6]) ? node1175 : node1114;
					assign node1114 = (inp[0]) ? node1132 : node1115;
						assign node1115 = (inp[7]) ? node1117 : 3'b000;
							assign node1117 = (inp[2]) ? node1119 : 3'b000;
								assign node1119 = (inp[10]) ? node1127 : node1120;
									assign node1120 = (inp[8]) ? node1124 : node1121;
										assign node1121 = (inp[5]) ? 3'b000 : 3'b100;
										assign node1124 = (inp[1]) ? 3'b100 : 3'b000;
									assign node1127 = (inp[11]) ? 3'b000 : node1128;
										assign node1128 = (inp[1]) ? 3'b000 : 3'b000;
						assign node1132 = (inp[10]) ? node1154 : node1133;
							assign node1133 = (inp[5]) ? node1147 : node1134;
								assign node1134 = (inp[7]) ? node1142 : node1135;
									assign node1135 = (inp[1]) ? node1139 : node1136;
										assign node1136 = (inp[2]) ? 3'b100 : 3'b000;
										assign node1139 = (inp[2]) ? 3'b010 : 3'b100;
									assign node1142 = (inp[11]) ? 3'b010 : node1143;
										assign node1143 = (inp[1]) ? 3'b110 : 3'b010;
								assign node1147 = (inp[1]) ? 3'b100 : node1148;
									assign node1148 = (inp[2]) ? node1150 : 3'b000;
										assign node1150 = (inp[8]) ? 3'b100 : 3'b000;
							assign node1154 = (inp[5]) ? node1168 : node1155;
								assign node1155 = (inp[2]) ? node1163 : node1156;
									assign node1156 = (inp[1]) ? node1160 : node1157;
										assign node1157 = (inp[11]) ? 3'b000 : 3'b000;
										assign node1160 = (inp[7]) ? 3'b010 : 3'b000;
									assign node1163 = (inp[11]) ? node1165 : 3'b100;
										assign node1165 = (inp[7]) ? 3'b100 : 3'b000;
								assign node1168 = (inp[1]) ? node1170 : 3'b000;
									assign node1170 = (inp[7]) ? node1172 : 3'b000;
										assign node1172 = (inp[8]) ? 3'b100 : 3'b000;
					assign node1175 = (inp[0]) ? node1221 : node1176;
						assign node1176 = (inp[5]) ? node1202 : node1177;
							assign node1177 = (inp[1]) ? node1191 : node1178;
								assign node1178 = (inp[8]) ? node1186 : node1179;
									assign node1179 = (inp[11]) ? node1183 : node1180;
										assign node1180 = (inp[10]) ? 3'b100 : 3'b000;
										assign node1183 = (inp[7]) ? 3'b100 : 3'b000;
									assign node1186 = (inp[11]) ? 3'b100 : node1187;
										assign node1187 = (inp[7]) ? 3'b100 : 3'b000;
								assign node1191 = (inp[7]) ? node1197 : node1192;
									assign node1192 = (inp[10]) ? 3'b100 : node1193;
										assign node1193 = (inp[8]) ? 3'b010 : 3'b000;
									assign node1197 = (inp[10]) ? 3'b010 : node1198;
										assign node1198 = (inp[8]) ? 3'b010 : 3'b010;
							assign node1202 = (inp[10]) ? node1216 : node1203;
								assign node1203 = (inp[11]) ? node1211 : node1204;
									assign node1204 = (inp[7]) ? node1208 : node1205;
										assign node1205 = (inp[8]) ? 3'b100 : 3'b000;
										assign node1208 = (inp[8]) ? 3'b010 : 3'b000;
									assign node1211 = (inp[8]) ? 3'b100 : node1212;
										assign node1212 = (inp[2]) ? 3'b100 : 3'b000;
								assign node1216 = (inp[7]) ? node1218 : 3'b000;
									assign node1218 = (inp[2]) ? 3'b100 : 3'b000;
						assign node1221 = (inp[1]) ? node1251 : node1222;
							assign node1222 = (inp[10]) ? node1236 : node1223;
								assign node1223 = (inp[2]) ? node1231 : node1224;
									assign node1224 = (inp[5]) ? node1228 : node1225;
										assign node1225 = (inp[8]) ? 3'b001 : 3'b110;
										assign node1228 = (inp[7]) ? 3'b110 : 3'b100;
									assign node1231 = (inp[11]) ? node1233 : 3'b110;
										assign node1233 = (inp[7]) ? 3'b110 : 3'b010;
								assign node1236 = (inp[5]) ? node1244 : node1237;
									assign node1237 = (inp[7]) ? node1241 : node1238;
										assign node1238 = (inp[2]) ? 3'b010 : 3'b100;
										assign node1241 = (inp[11]) ? 3'b010 : 3'b110;
									assign node1244 = (inp[11]) ? node1248 : node1245;
										assign node1245 = (inp[7]) ? 3'b010 : 3'b100;
										assign node1248 = (inp[7]) ? 3'b100 : 3'b000;
							assign node1251 = (inp[5]) ? node1265 : node1252;
								assign node1252 = (inp[10]) ? node1260 : node1253;
									assign node1253 = (inp[7]) ? node1257 : node1254;
										assign node1254 = (inp[11]) ? 3'b110 : 3'b001;
										assign node1257 = (inp[8]) ? 3'b001 : 3'b001;
									assign node1260 = (inp[11]) ? 3'b010 : node1261;
										assign node1261 = (inp[7]) ? 3'b000 : 3'b110;
								assign node1265 = (inp[2]) ? node1271 : node1266;
									assign node1266 = (inp[7]) ? node1268 : 3'b010;
										assign node1268 = (inp[10]) ? 3'b010 : 3'b110;
									assign node1271 = (inp[11]) ? node1275 : node1272;
										assign node1272 = (inp[7]) ? 3'b000 : 3'b110;
										assign node1275 = (inp[10]) ? 3'b100 : 3'b110;
				assign node1278 = (inp[0]) ? node1292 : node1279;
					assign node1279 = (inp[1]) ? node1281 : 3'b000;
						assign node1281 = (inp[6]) ? node1283 : 3'b000;
							assign node1283 = (inp[10]) ? 3'b000 : node1284;
								assign node1284 = (inp[5]) ? 3'b000 : node1285;
									assign node1285 = (inp[7]) ? node1287 : 3'b000;
										assign node1287 = (inp[2]) ? 3'b100 : 3'b000;
					assign node1292 = (inp[6]) ? node1304 : node1293;
						assign node1293 = (inp[1]) ? node1295 : 3'b000;
							assign node1295 = (inp[11]) ? 3'b000 : node1296;
								assign node1296 = (inp[7]) ? node1298 : 3'b000;
									assign node1298 = (inp[10]) ? 3'b000 : node1299;
										assign node1299 = (inp[2]) ? 3'b100 : 3'b000;
						assign node1304 = (inp[10]) ? node1324 : node1305;
							assign node1305 = (inp[5]) ? node1317 : node1306;
								assign node1306 = (inp[7]) ? node1312 : node1307;
									assign node1307 = (inp[11]) ? 3'b100 : node1308;
										assign node1308 = (inp[1]) ? 3'b000 : 3'b100;
									assign node1312 = (inp[2]) ? 3'b010 : node1313;
										assign node1313 = (inp[1]) ? 3'b010 : 3'b100;
								assign node1317 = (inp[7]) ? node1319 : 3'b000;
									assign node1319 = (inp[8]) ? 3'b100 : node1320;
										assign node1320 = (inp[1]) ? 3'b000 : 3'b000;
							assign node1324 = (inp[1]) ? node1326 : 3'b000;
								assign node1326 = (inp[7]) ? node1328 : 3'b000;
									assign node1328 = (inp[5]) ? 3'b000 : 3'b100;

endmodule