module dtc_split125_bm62 (
	input  wire [16-1:0] inp,
	output wire [4-1:0] outp
);

	wire [4-1:0] node1;
	wire [4-1:0] node2;
	wire [4-1:0] node3;
	wire [4-1:0] node4;
	wire [4-1:0] node5;
	wire [4-1:0] node6;
	wire [4-1:0] node7;
	wire [4-1:0] node8;
	wire [4-1:0] node9;
	wire [4-1:0] node10;
	wire [4-1:0] node11;
	wire [4-1:0] node13;
	wire [4-1:0] node15;
	wire [4-1:0] node18;
	wire [4-1:0] node19;
	wire [4-1:0] node23;
	wire [4-1:0] node24;
	wire [4-1:0] node25;
	wire [4-1:0] node26;
	wire [4-1:0] node31;
	wire [4-1:0] node33;
	wire [4-1:0] node36;
	wire [4-1:0] node37;
	wire [4-1:0] node38;
	wire [4-1:0] node40;
	wire [4-1:0] node43;
	wire [4-1:0] node44;
	wire [4-1:0] node46;
	wire [4-1:0] node49;
	wire [4-1:0] node50;
	wire [4-1:0] node53;
	wire [4-1:0] node56;
	wire [4-1:0] node57;
	wire [4-1:0] node59;
	wire [4-1:0] node62;
	wire [4-1:0] node64;
	wire [4-1:0] node67;
	wire [4-1:0] node68;
	wire [4-1:0] node69;
	wire [4-1:0] node71;
	wire [4-1:0] node72;
	wire [4-1:0] node73;
	wire [4-1:0] node78;
	wire [4-1:0] node79;
	wire [4-1:0] node81;
	wire [4-1:0] node83;
	wire [4-1:0] node86;
	wire [4-1:0] node88;
	wire [4-1:0] node91;
	wire [4-1:0] node92;
	wire [4-1:0] node94;
	wire [4-1:0] node95;
	wire [4-1:0] node99;
	wire [4-1:0] node100;
	wire [4-1:0] node101;
	wire [4-1:0] node104;
	wire [4-1:0] node107;
	wire [4-1:0] node110;
	wire [4-1:0] node111;
	wire [4-1:0] node112;
	wire [4-1:0] node113;
	wire [4-1:0] node115;
	wire [4-1:0] node117;
	wire [4-1:0] node120;
	wire [4-1:0] node121;
	wire [4-1:0] node122;
	wire [4-1:0] node126;
	wire [4-1:0] node127;
	wire [4-1:0] node131;
	wire [4-1:0] node132;
	wire [4-1:0] node133;
	wire [4-1:0] node136;
	wire [4-1:0] node138;
	wire [4-1:0] node141;
	wire [4-1:0] node142;
	wire [4-1:0] node143;
	wire [4-1:0] node146;
	wire [4-1:0] node148;
	wire [4-1:0] node152;
	wire [4-1:0] node153;
	wire [4-1:0] node154;
	wire [4-1:0] node155;
	wire [4-1:0] node158;
	wire [4-1:0] node159;
	wire [4-1:0] node160;
	wire [4-1:0] node164;
	wire [4-1:0] node167;
	wire [4-1:0] node168;
	wire [4-1:0] node169;
	wire [4-1:0] node170;
	wire [4-1:0] node173;
	wire [4-1:0] node176;
	wire [4-1:0] node178;
	wire [4-1:0] node182;
	wire [4-1:0] node183;
	wire [4-1:0] node186;
	wire [4-1:0] node187;
	wire [4-1:0] node188;
	wire [4-1:0] node189;
	wire [4-1:0] node193;
	wire [4-1:0] node196;
	wire [4-1:0] node197;
	wire [4-1:0] node199;
	wire [4-1:0] node202;
	wire [4-1:0] node205;
	wire [4-1:0] node206;
	wire [4-1:0] node207;
	wire [4-1:0] node208;
	wire [4-1:0] node209;
	wire [4-1:0] node210;
	wire [4-1:0] node211;
	wire [4-1:0] node214;
	wire [4-1:0] node215;
	wire [4-1:0] node218;
	wire [4-1:0] node222;
	wire [4-1:0] node223;
	wire [4-1:0] node224;
	wire [4-1:0] node227;
	wire [4-1:0] node230;
	wire [4-1:0] node233;
	wire [4-1:0] node234;
	wire [4-1:0] node235;
	wire [4-1:0] node239;
	wire [4-1:0] node240;
	wire [4-1:0] node243;
	wire [4-1:0] node244;
	wire [4-1:0] node245;
	wire [4-1:0] node250;
	wire [4-1:0] node251;
	wire [4-1:0] node252;
	wire [4-1:0] node253;
	wire [4-1:0] node256;
	wire [4-1:0] node257;
	wire [4-1:0] node261;
	wire [4-1:0] node262;
	wire [4-1:0] node263;
	wire [4-1:0] node264;
	wire [4-1:0] node268;
	wire [4-1:0] node271;
	wire [4-1:0] node274;
	wire [4-1:0] node275;
	wire [4-1:0] node276;
	wire [4-1:0] node278;
	wire [4-1:0] node281;
	wire [4-1:0] node282;
	wire [4-1:0] node285;
	wire [4-1:0] node286;
	wire [4-1:0] node290;
	wire [4-1:0] node291;
	wire [4-1:0] node292;
	wire [4-1:0] node296;
	wire [4-1:0] node297;
	wire [4-1:0] node301;
	wire [4-1:0] node302;
	wire [4-1:0] node303;
	wire [4-1:0] node304;
	wire [4-1:0] node305;
	wire [4-1:0] node307;
	wire [4-1:0] node310;
	wire [4-1:0] node311;
	wire [4-1:0] node312;
	wire [4-1:0] node317;
	wire [4-1:0] node318;
	wire [4-1:0] node319;
	wire [4-1:0] node320;
	wire [4-1:0] node323;
	wire [4-1:0] node326;
	wire [4-1:0] node329;
	wire [4-1:0] node330;
	wire [4-1:0] node334;
	wire [4-1:0] node335;
	wire [4-1:0] node337;
	wire [4-1:0] node339;
	wire [4-1:0] node342;
	wire [4-1:0] node343;
	wire [4-1:0] node344;
	wire [4-1:0] node348;
	wire [4-1:0] node349;
	wire [4-1:0] node353;
	wire [4-1:0] node354;
	wire [4-1:0] node355;
	wire [4-1:0] node357;
	wire [4-1:0] node358;
	wire [4-1:0] node360;
	wire [4-1:0] node364;
	wire [4-1:0] node365;
	wire [4-1:0] node369;
	wire [4-1:0] node370;
	wire [4-1:0] node371;
	wire [4-1:0] node374;
	wire [4-1:0] node375;
	wire [4-1:0] node379;
	wire [4-1:0] node380;
	wire [4-1:0] node383;
	wire [4-1:0] node385;
	wire [4-1:0] node388;
	wire [4-1:0] node389;
	wire [4-1:0] node390;
	wire [4-1:0] node391;
	wire [4-1:0] node392;
	wire [4-1:0] node393;
	wire [4-1:0] node395;
	wire [4-1:0] node397;
	wire [4-1:0] node400;
	wire [4-1:0] node401;
	wire [4-1:0] node403;
	wire [4-1:0] node404;
	wire [4-1:0] node408;
	wire [4-1:0] node411;
	wire [4-1:0] node412;
	wire [4-1:0] node413;
	wire [4-1:0] node414;
	wire [4-1:0] node417;
	wire [4-1:0] node421;
	wire [4-1:0] node422;
	wire [4-1:0] node424;
	wire [4-1:0] node428;
	wire [4-1:0] node429;
	wire [4-1:0] node430;
	wire [4-1:0] node431;
	wire [4-1:0] node432;
	wire [4-1:0] node437;
	wire [4-1:0] node438;
	wire [4-1:0] node440;
	wire [4-1:0] node443;
	wire [4-1:0] node446;
	wire [4-1:0] node448;
	wire [4-1:0] node449;
	wire [4-1:0] node451;
	wire [4-1:0] node454;
	wire [4-1:0] node455;
	wire [4-1:0] node458;
	wire [4-1:0] node459;
	wire [4-1:0] node463;
	wire [4-1:0] node464;
	wire [4-1:0] node465;
	wire [4-1:0] node466;
	wire [4-1:0] node469;
	wire [4-1:0] node470;
	wire [4-1:0] node471;
	wire [4-1:0] node474;
	wire [4-1:0] node477;
	wire [4-1:0] node478;
	wire [4-1:0] node482;
	wire [4-1:0] node483;
	wire [4-1:0] node484;
	wire [4-1:0] node486;
	wire [4-1:0] node490;
	wire [4-1:0] node492;
	wire [4-1:0] node494;
	wire [4-1:0] node497;
	wire [4-1:0] node498;
	wire [4-1:0] node499;
	wire [4-1:0] node500;
	wire [4-1:0] node502;
	wire [4-1:0] node504;
	wire [4-1:0] node507;
	wire [4-1:0] node510;
	wire [4-1:0] node511;
	wire [4-1:0] node513;
	wire [4-1:0] node514;
	wire [4-1:0] node518;
	wire [4-1:0] node519;
	wire [4-1:0] node521;
	wire [4-1:0] node524;
	wire [4-1:0] node527;
	wire [4-1:0] node528;
	wire [4-1:0] node529;
	wire [4-1:0] node533;
	wire [4-1:0] node534;
	wire [4-1:0] node535;
	wire [4-1:0] node540;
	wire [4-1:0] node541;
	wire [4-1:0] node542;
	wire [4-1:0] node543;
	wire [4-1:0] node544;
	wire [4-1:0] node545;
	wire [4-1:0] node546;
	wire [4-1:0] node549;
	wire [4-1:0] node552;
	wire [4-1:0] node555;
	wire [4-1:0] node556;
	wire [4-1:0] node558;
	wire [4-1:0] node561;
	wire [4-1:0] node562;
	wire [4-1:0] node565;
	wire [4-1:0] node568;
	wire [4-1:0] node569;
	wire [4-1:0] node570;
	wire [4-1:0] node572;
	wire [4-1:0] node575;
	wire [4-1:0] node577;
	wire [4-1:0] node579;
	wire [4-1:0] node582;
	wire [4-1:0] node583;
	wire [4-1:0] node584;
	wire [4-1:0] node586;
	wire [4-1:0] node589;
	wire [4-1:0] node592;
	wire [4-1:0] node593;
	wire [4-1:0] node597;
	wire [4-1:0] node598;
	wire [4-1:0] node599;
	wire [4-1:0] node600;
	wire [4-1:0] node601;
	wire [4-1:0] node605;
	wire [4-1:0] node608;
	wire [4-1:0] node609;
	wire [4-1:0] node610;
	wire [4-1:0] node613;
	wire [4-1:0] node614;
	wire [4-1:0] node618;
	wire [4-1:0] node619;
	wire [4-1:0] node622;
	wire [4-1:0] node623;
	wire [4-1:0] node627;
	wire [4-1:0] node628;
	wire [4-1:0] node629;
	wire [4-1:0] node633;
	wire [4-1:0] node635;
	wire [4-1:0] node638;
	wire [4-1:0] node639;
	wire [4-1:0] node640;
	wire [4-1:0] node641;
	wire [4-1:0] node642;
	wire [4-1:0] node644;
	wire [4-1:0] node647;
	wire [4-1:0] node648;
	wire [4-1:0] node652;
	wire [4-1:0] node653;
	wire [4-1:0] node654;
	wire [4-1:0] node656;
	wire [4-1:0] node660;
	wire [4-1:0] node663;
	wire [4-1:0] node664;
	wire [4-1:0] node665;
	wire [4-1:0] node666;
	wire [4-1:0] node667;
	wire [4-1:0] node672;
	wire [4-1:0] node674;
	wire [4-1:0] node677;
	wire [4-1:0] node679;
	wire [4-1:0] node682;
	wire [4-1:0] node683;
	wire [4-1:0] node684;
	wire [4-1:0] node685;
	wire [4-1:0] node686;
	wire [4-1:0] node687;
	wire [4-1:0] node691;
	wire [4-1:0] node694;
	wire [4-1:0] node696;
	wire [4-1:0] node697;
	wire [4-1:0] node701;
	wire [4-1:0] node702;
	wire [4-1:0] node705;
	wire [4-1:0] node706;
	wire [4-1:0] node709;
	wire [4-1:0] node710;
	wire [4-1:0] node713;
	wire [4-1:0] node716;
	wire [4-1:0] node717;
	wire [4-1:0] node720;
	wire [4-1:0] node721;
	wire [4-1:0] node722;
	wire [4-1:0] node723;
	wire [4-1:0] node727;
	wire [4-1:0] node728;
	wire [4-1:0] node731;
	wire [4-1:0] node734;
	wire [4-1:0] node737;
	wire [4-1:0] node738;
	wire [4-1:0] node739;
	wire [4-1:0] node740;
	wire [4-1:0] node741;
	wire [4-1:0] node742;
	wire [4-1:0] node743;
	wire [4-1:0] node744;
	wire [4-1:0] node747;
	wire [4-1:0] node749;
	wire [4-1:0] node750;
	wire [4-1:0] node754;
	wire [4-1:0] node755;
	wire [4-1:0] node758;
	wire [4-1:0] node760;
	wire [4-1:0] node763;
	wire [4-1:0] node764;
	wire [4-1:0] node766;
	wire [4-1:0] node768;
	wire [4-1:0] node771;
	wire [4-1:0] node774;
	wire [4-1:0] node775;
	wire [4-1:0] node776;
	wire [4-1:0] node778;
	wire [4-1:0] node779;
	wire [4-1:0] node780;
	wire [4-1:0] node783;
	wire [4-1:0] node787;
	wire [4-1:0] node788;
	wire [4-1:0] node790;
	wire [4-1:0] node793;
	wire [4-1:0] node795;
	wire [4-1:0] node796;
	wire [4-1:0] node800;
	wire [4-1:0] node801;
	wire [4-1:0] node802;
	wire [4-1:0] node804;
	wire [4-1:0] node805;
	wire [4-1:0] node809;
	wire [4-1:0] node810;
	wire [4-1:0] node811;
	wire [4-1:0] node816;
	wire [4-1:0] node817;
	wire [4-1:0] node818;
	wire [4-1:0] node822;
	wire [4-1:0] node823;
	wire [4-1:0] node824;
	wire [4-1:0] node828;
	wire [4-1:0] node830;
	wire [4-1:0] node833;
	wire [4-1:0] node834;
	wire [4-1:0] node835;
	wire [4-1:0] node836;
	wire [4-1:0] node837;
	wire [4-1:0] node838;
	wire [4-1:0] node839;
	wire [4-1:0] node845;
	wire [4-1:0] node846;
	wire [4-1:0] node847;
	wire [4-1:0] node850;
	wire [4-1:0] node853;
	wire [4-1:0] node855;
	wire [4-1:0] node858;
	wire [4-1:0] node859;
	wire [4-1:0] node860;
	wire [4-1:0] node861;
	wire [4-1:0] node865;
	wire [4-1:0] node867;
	wire [4-1:0] node869;
	wire [4-1:0] node872;
	wire [4-1:0] node874;
	wire [4-1:0] node875;
	wire [4-1:0] node877;
	wire [4-1:0] node881;
	wire [4-1:0] node882;
	wire [4-1:0] node883;
	wire [4-1:0] node885;
	wire [4-1:0] node886;
	wire [4-1:0] node890;
	wire [4-1:0] node891;
	wire [4-1:0] node892;
	wire [4-1:0] node895;
	wire [4-1:0] node899;
	wire [4-1:0] node900;
	wire [4-1:0] node901;
	wire [4-1:0] node902;
	wire [4-1:0] node907;
	wire [4-1:0] node908;
	wire [4-1:0] node909;
	wire [4-1:0] node910;
	wire [4-1:0] node916;
	wire [4-1:0] node917;
	wire [4-1:0] node918;
	wire [4-1:0] node919;
	wire [4-1:0] node920;
	wire [4-1:0] node921;
	wire [4-1:0] node923;
	wire [4-1:0] node926;
	wire [4-1:0] node929;
	wire [4-1:0] node930;
	wire [4-1:0] node932;
	wire [4-1:0] node935;
	wire [4-1:0] node938;
	wire [4-1:0] node939;
	wire [4-1:0] node940;
	wire [4-1:0] node944;
	wire [4-1:0] node945;
	wire [4-1:0] node946;
	wire [4-1:0] node951;
	wire [4-1:0] node952;
	wire [4-1:0] node953;
	wire [4-1:0] node954;
	wire [4-1:0] node957;
	wire [4-1:0] node960;
	wire [4-1:0] node962;
	wire [4-1:0] node963;
	wire [4-1:0] node965;
	wire [4-1:0] node969;
	wire [4-1:0] node970;
	wire [4-1:0] node971;
	wire [4-1:0] node973;
	wire [4-1:0] node976;
	wire [4-1:0] node977;
	wire [4-1:0] node979;
	wire [4-1:0] node983;
	wire [4-1:0] node984;
	wire [4-1:0] node986;
	wire [4-1:0] node987;
	wire [4-1:0] node991;
	wire [4-1:0] node993;
	wire [4-1:0] node996;
	wire [4-1:0] node997;
	wire [4-1:0] node998;
	wire [4-1:0] node999;
	wire [4-1:0] node1001;
	wire [4-1:0] node1004;
	wire [4-1:0] node1006;
	wire [4-1:0] node1009;
	wire [4-1:0] node1010;
	wire [4-1:0] node1012;
	wire [4-1:0] node1015;
	wire [4-1:0] node1016;
	wire [4-1:0] node1017;
	wire [4-1:0] node1018;
	wire [4-1:0] node1024;
	wire [4-1:0] node1025;
	wire [4-1:0] node1026;
	wire [4-1:0] node1027;
	wire [4-1:0] node1029;
	wire [4-1:0] node1032;
	wire [4-1:0] node1033;
	wire [4-1:0] node1036;
	wire [4-1:0] node1039;
	wire [4-1:0] node1041;
	wire [4-1:0] node1044;
	wire [4-1:0] node1045;
	wire [4-1:0] node1047;
	wire [4-1:0] node1049;
	wire [4-1:0] node1052;
	wire [4-1:0] node1053;
	wire [4-1:0] node1055;
	wire [4-1:0] node1056;
	wire [4-1:0] node1060;
	wire [4-1:0] node1063;
	wire [4-1:0] node1064;
	wire [4-1:0] node1065;
	wire [4-1:0] node1066;
	wire [4-1:0] node1067;
	wire [4-1:0] node1068;
	wire [4-1:0] node1069;
	wire [4-1:0] node1071;
	wire [4-1:0] node1072;
	wire [4-1:0] node1077;
	wire [4-1:0] node1078;
	wire [4-1:0] node1081;
	wire [4-1:0] node1082;
	wire [4-1:0] node1084;
	wire [4-1:0] node1088;
	wire [4-1:0] node1089;
	wire [4-1:0] node1090;
	wire [4-1:0] node1091;
	wire [4-1:0] node1095;
	wire [4-1:0] node1097;
	wire [4-1:0] node1099;
	wire [4-1:0] node1102;
	wire [4-1:0] node1104;
	wire [4-1:0] node1105;
	wire [4-1:0] node1108;
	wire [4-1:0] node1111;
	wire [4-1:0] node1112;
	wire [4-1:0] node1113;
	wire [4-1:0] node1114;
	wire [4-1:0] node1115;
	wire [4-1:0] node1117;
	wire [4-1:0] node1122;
	wire [4-1:0] node1123;
	wire [4-1:0] node1126;
	wire [4-1:0] node1129;
	wire [4-1:0] node1130;
	wire [4-1:0] node1131;
	wire [4-1:0] node1132;
	wire [4-1:0] node1135;
	wire [4-1:0] node1139;
	wire [4-1:0] node1140;
	wire [4-1:0] node1141;
	wire [4-1:0] node1142;
	wire [4-1:0] node1146;
	wire [4-1:0] node1149;
	wire [4-1:0] node1151;
	wire [4-1:0] node1154;
	wire [4-1:0] node1155;
	wire [4-1:0] node1156;
	wire [4-1:0] node1157;
	wire [4-1:0] node1158;
	wire [4-1:0] node1160;
	wire [4-1:0] node1162;
	wire [4-1:0] node1166;
	wire [4-1:0] node1167;
	wire [4-1:0] node1171;
	wire [4-1:0] node1172;
	wire [4-1:0] node1173;
	wire [4-1:0] node1176;
	wire [4-1:0] node1179;
	wire [4-1:0] node1180;
	wire [4-1:0] node1182;
	wire [4-1:0] node1185;
	wire [4-1:0] node1186;
	wire [4-1:0] node1190;
	wire [4-1:0] node1191;
	wire [4-1:0] node1192;
	wire [4-1:0] node1193;
	wire [4-1:0] node1197;
	wire [4-1:0] node1200;
	wire [4-1:0] node1201;
	wire [4-1:0] node1202;
	wire [4-1:0] node1203;
	wire [4-1:0] node1204;
	wire [4-1:0] node1209;
	wire [4-1:0] node1211;
	wire [4-1:0] node1213;
	wire [4-1:0] node1216;
	wire [4-1:0] node1217;
	wire [4-1:0] node1218;
	wire [4-1:0] node1220;
	wire [4-1:0] node1224;
	wire [4-1:0] node1225;
	wire [4-1:0] node1228;
	wire [4-1:0] node1231;
	wire [4-1:0] node1232;
	wire [4-1:0] node1233;
	wire [4-1:0] node1234;
	wire [4-1:0] node1235;
	wire [4-1:0] node1236;
	wire [4-1:0] node1239;
	wire [4-1:0] node1242;
	wire [4-1:0] node1243;
	wire [4-1:0] node1244;
	wire [4-1:0] node1246;
	wire [4-1:0] node1249;
	wire [4-1:0] node1253;
	wire [4-1:0] node1254;
	wire [4-1:0] node1255;
	wire [4-1:0] node1258;
	wire [4-1:0] node1260;
	wire [4-1:0] node1261;
	wire [4-1:0] node1264;
	wire [4-1:0] node1267;
	wire [4-1:0] node1268;
	wire [4-1:0] node1270;
	wire [4-1:0] node1273;
	wire [4-1:0] node1276;
	wire [4-1:0] node1277;
	wire [4-1:0] node1278;
	wire [4-1:0] node1279;
	wire [4-1:0] node1280;
	wire [4-1:0] node1283;
	wire [4-1:0] node1286;
	wire [4-1:0] node1287;
	wire [4-1:0] node1290;
	wire [4-1:0] node1292;
	wire [4-1:0] node1295;
	wire [4-1:0] node1296;
	wire [4-1:0] node1297;
	wire [4-1:0] node1298;
	wire [4-1:0] node1302;
	wire [4-1:0] node1306;
	wire [4-1:0] node1307;
	wire [4-1:0] node1308;
	wire [4-1:0] node1310;
	wire [4-1:0] node1314;
	wire [4-1:0] node1316;
	wire [4-1:0] node1317;
	wire [4-1:0] node1320;
	wire [4-1:0] node1323;
	wire [4-1:0] node1324;
	wire [4-1:0] node1325;
	wire [4-1:0] node1326;
	wire [4-1:0] node1328;
	wire [4-1:0] node1329;
	wire [4-1:0] node1330;
	wire [4-1:0] node1334;
	wire [4-1:0] node1337;
	wire [4-1:0] node1338;
	wire [4-1:0] node1341;
	wire [4-1:0] node1344;
	wire [4-1:0] node1345;
	wire [4-1:0] node1346;
	wire [4-1:0] node1347;
	wire [4-1:0] node1348;
	wire [4-1:0] node1353;
	wire [4-1:0] node1354;
	wire [4-1:0] node1355;
	wire [4-1:0] node1360;
	wire [4-1:0] node1361;
	wire [4-1:0] node1364;
	wire [4-1:0] node1365;
	wire [4-1:0] node1368;
	wire [4-1:0] node1371;
	wire [4-1:0] node1372;
	wire [4-1:0] node1373;
	wire [4-1:0] node1374;
	wire [4-1:0] node1376;
	wire [4-1:0] node1379;
	wire [4-1:0] node1380;
	wire [4-1:0] node1384;
	wire [4-1:0] node1385;
	wire [4-1:0] node1389;
	wire [4-1:0] node1390;
	wire [4-1:0] node1393;
	wire [4-1:0] node1394;
	wire [4-1:0] node1395;
	wire [4-1:0] node1398;
	wire [4-1:0] node1401;
	wire [4-1:0] node1403;
	wire [4-1:0] node1404;
	wire [4-1:0] node1408;
	wire [4-1:0] node1409;
	wire [4-1:0] node1410;
	wire [4-1:0] node1411;
	wire [4-1:0] node1412;
	wire [4-1:0] node1413;
	wire [4-1:0] node1414;
	wire [4-1:0] node1415;
	wire [4-1:0] node1417;
	wire [4-1:0] node1418;
	wire [4-1:0] node1419;
	wire [4-1:0] node1422;
	wire [4-1:0] node1426;
	wire [4-1:0] node1427;
	wire [4-1:0] node1429;
	wire [4-1:0] node1432;
	wire [4-1:0] node1435;
	wire [4-1:0] node1436;
	wire [4-1:0] node1438;
	wire [4-1:0] node1440;
	wire [4-1:0] node1443;
	wire [4-1:0] node1445;
	wire [4-1:0] node1446;
	wire [4-1:0] node1450;
	wire [4-1:0] node1451;
	wire [4-1:0] node1452;
	wire [4-1:0] node1453;
	wire [4-1:0] node1454;
	wire [4-1:0] node1458;
	wire [4-1:0] node1461;
	wire [4-1:0] node1463;
	wire [4-1:0] node1465;
	wire [4-1:0] node1468;
	wire [4-1:0] node1469;
	wire [4-1:0] node1470;
	wire [4-1:0] node1473;
	wire [4-1:0] node1474;
	wire [4-1:0] node1478;
	wire [4-1:0] node1481;
	wire [4-1:0] node1482;
	wire [4-1:0] node1483;
	wire [4-1:0] node1485;
	wire [4-1:0] node1486;
	wire [4-1:0] node1489;
	wire [4-1:0] node1490;
	wire [4-1:0] node1493;
	wire [4-1:0] node1496;
	wire [4-1:0] node1497;
	wire [4-1:0] node1498;
	wire [4-1:0] node1501;
	wire [4-1:0] node1503;
	wire [4-1:0] node1506;
	wire [4-1:0] node1508;
	wire [4-1:0] node1509;
	wire [4-1:0] node1511;
	wire [4-1:0] node1515;
	wire [4-1:0] node1516;
	wire [4-1:0] node1517;
	wire [4-1:0] node1518;
	wire [4-1:0] node1519;
	wire [4-1:0] node1523;
	wire [4-1:0] node1524;
	wire [4-1:0] node1525;
	wire [4-1:0] node1530;
	wire [4-1:0] node1531;
	wire [4-1:0] node1534;
	wire [4-1:0] node1535;
	wire [4-1:0] node1536;
	wire [4-1:0] node1540;
	wire [4-1:0] node1543;
	wire [4-1:0] node1544;
	wire [4-1:0] node1547;
	wire [4-1:0] node1548;
	wire [4-1:0] node1549;
	wire [4-1:0] node1551;
	wire [4-1:0] node1554;
	wire [4-1:0] node1556;
	wire [4-1:0] node1559;
	wire [4-1:0] node1561;
	wire [4-1:0] node1564;
	wire [4-1:0] node1565;
	wire [4-1:0] node1566;
	wire [4-1:0] node1567;
	wire [4-1:0] node1568;
	wire [4-1:0] node1570;
	wire [4-1:0] node1571;
	wire [4-1:0] node1575;
	wire [4-1:0] node1577;
	wire [4-1:0] node1578;
	wire [4-1:0] node1581;
	wire [4-1:0] node1582;
	wire [4-1:0] node1586;
	wire [4-1:0] node1587;
	wire [4-1:0] node1588;
	wire [4-1:0] node1589;
	wire [4-1:0] node1593;
	wire [4-1:0] node1595;
	wire [4-1:0] node1598;
	wire [4-1:0] node1599;
	wire [4-1:0] node1600;
	wire [4-1:0] node1602;
	wire [4-1:0] node1606;
	wire [4-1:0] node1608;
	wire [4-1:0] node1611;
	wire [4-1:0] node1612;
	wire [4-1:0] node1613;
	wire [4-1:0] node1614;
	wire [4-1:0] node1617;
	wire [4-1:0] node1618;
	wire [4-1:0] node1622;
	wire [4-1:0] node1623;
	wire [4-1:0] node1626;
	wire [4-1:0] node1627;
	wire [4-1:0] node1631;
	wire [4-1:0] node1632;
	wire [4-1:0] node1633;
	wire [4-1:0] node1634;
	wire [4-1:0] node1638;
	wire [4-1:0] node1641;
	wire [4-1:0] node1642;
	wire [4-1:0] node1644;
	wire [4-1:0] node1647;
	wire [4-1:0] node1649;
	wire [4-1:0] node1651;
	wire [4-1:0] node1654;
	wire [4-1:0] node1655;
	wire [4-1:0] node1656;
	wire [4-1:0] node1657;
	wire [4-1:0] node1658;
	wire [4-1:0] node1661;
	wire [4-1:0] node1664;
	wire [4-1:0] node1666;
	wire [4-1:0] node1667;
	wire [4-1:0] node1669;
	wire [4-1:0] node1673;
	wire [4-1:0] node1674;
	wire [4-1:0] node1675;
	wire [4-1:0] node1678;
	wire [4-1:0] node1679;
	wire [4-1:0] node1680;
	wire [4-1:0] node1683;
	wire [4-1:0] node1687;
	wire [4-1:0] node1688;
	wire [4-1:0] node1689;
	wire [4-1:0] node1692;
	wire [4-1:0] node1694;
	wire [4-1:0] node1697;
	wire [4-1:0] node1698;
	wire [4-1:0] node1699;
	wire [4-1:0] node1704;
	wire [4-1:0] node1705;
	wire [4-1:0] node1706;
	wire [4-1:0] node1707;
	wire [4-1:0] node1708;
	wire [4-1:0] node1711;
	wire [4-1:0] node1715;
	wire [4-1:0] node1716;
	wire [4-1:0] node1718;
	wire [4-1:0] node1721;
	wire [4-1:0] node1723;
	wire [4-1:0] node1726;
	wire [4-1:0] node1727;
	wire [4-1:0] node1728;
	wire [4-1:0] node1730;
	wire [4-1:0] node1733;
	wire [4-1:0] node1734;
	wire [4-1:0] node1735;
	wire [4-1:0] node1738;
	wire [4-1:0] node1742;
	wire [4-1:0] node1743;
	wire [4-1:0] node1744;
	wire [4-1:0] node1747;
	wire [4-1:0] node1750;
	wire [4-1:0] node1753;
	wire [4-1:0] node1754;
	wire [4-1:0] node1755;
	wire [4-1:0] node1756;
	wire [4-1:0] node1757;
	wire [4-1:0] node1758;
	wire [4-1:0] node1761;
	wire [4-1:0] node1763;
	wire [4-1:0] node1766;
	wire [4-1:0] node1767;
	wire [4-1:0] node1768;
	wire [4-1:0] node1769;
	wire [4-1:0] node1771;
	wire [4-1:0] node1774;
	wire [4-1:0] node1777;
	wire [4-1:0] node1778;
	wire [4-1:0] node1780;
	wire [4-1:0] node1784;
	wire [4-1:0] node1786;
	wire [4-1:0] node1787;
	wire [4-1:0] node1791;
	wire [4-1:0] node1792;
	wire [4-1:0] node1793;
	wire [4-1:0] node1794;
	wire [4-1:0] node1796;
	wire [4-1:0] node1799;
	wire [4-1:0] node1800;
	wire [4-1:0] node1801;
	wire [4-1:0] node1806;
	wire [4-1:0] node1807;
	wire [4-1:0] node1808;
	wire [4-1:0] node1810;
	wire [4-1:0] node1815;
	wire [4-1:0] node1816;
	wire [4-1:0] node1817;
	wire [4-1:0] node1818;
	wire [4-1:0] node1821;
	wire [4-1:0] node1825;
	wire [4-1:0] node1827;
	wire [4-1:0] node1828;
	wire [4-1:0] node1830;
	wire [4-1:0] node1833;
	wire [4-1:0] node1836;
	wire [4-1:0] node1837;
	wire [4-1:0] node1838;
	wire [4-1:0] node1839;
	wire [4-1:0] node1840;
	wire [4-1:0] node1842;
	wire [4-1:0] node1845;
	wire [4-1:0] node1846;
	wire [4-1:0] node1850;
	wire [4-1:0] node1851;
	wire [4-1:0] node1852;
	wire [4-1:0] node1853;
	wire [4-1:0] node1858;
	wire [4-1:0] node1859;
	wire [4-1:0] node1861;
	wire [4-1:0] node1864;
	wire [4-1:0] node1866;
	wire [4-1:0] node1869;
	wire [4-1:0] node1870;
	wire [4-1:0] node1871;
	wire [4-1:0] node1873;
	wire [4-1:0] node1875;
	wire [4-1:0] node1878;
	wire [4-1:0] node1881;
	wire [4-1:0] node1883;
	wire [4-1:0] node1885;
	wire [4-1:0] node1888;
	wire [4-1:0] node1889;
	wire [4-1:0] node1890;
	wire [4-1:0] node1892;
	wire [4-1:0] node1894;
	wire [4-1:0] node1897;
	wire [4-1:0] node1898;
	wire [4-1:0] node1899;
	wire [4-1:0] node1900;
	wire [4-1:0] node1903;
	wire [4-1:0] node1908;
	wire [4-1:0] node1909;
	wire [4-1:0] node1910;
	wire [4-1:0] node1912;
	wire [4-1:0] node1913;
	wire [4-1:0] node1917;
	wire [4-1:0] node1918;
	wire [4-1:0] node1922;
	wire [4-1:0] node1924;
	wire [4-1:0] node1927;
	wire [4-1:0] node1928;
	wire [4-1:0] node1929;
	wire [4-1:0] node1930;
	wire [4-1:0] node1931;
	wire [4-1:0] node1933;
	wire [4-1:0] node1936;
	wire [4-1:0] node1937;
	wire [4-1:0] node1940;
	wire [4-1:0] node1941;
	wire [4-1:0] node1944;
	wire [4-1:0] node1946;
	wire [4-1:0] node1949;
	wire [4-1:0] node1950;
	wire [4-1:0] node1951;
	wire [4-1:0] node1954;
	wire [4-1:0] node1955;
	wire [4-1:0] node1957;
	wire [4-1:0] node1961;
	wire [4-1:0] node1963;
	wire [4-1:0] node1964;
	wire [4-1:0] node1968;
	wire [4-1:0] node1969;
	wire [4-1:0] node1970;
	wire [4-1:0] node1972;
	wire [4-1:0] node1974;
	wire [4-1:0] node1977;
	wire [4-1:0] node1978;
	wire [4-1:0] node1982;
	wire [4-1:0] node1983;
	wire [4-1:0] node1984;
	wire [4-1:0] node1988;
	wire [4-1:0] node1989;
	wire [4-1:0] node1990;
	wire [4-1:0] node1991;
	wire [4-1:0] node1996;
	wire [4-1:0] node1998;
	wire [4-1:0] node2001;
	wire [4-1:0] node2002;
	wire [4-1:0] node2003;
	wire [4-1:0] node2004;
	wire [4-1:0] node2005;
	wire [4-1:0] node2007;
	wire [4-1:0] node2010;
	wire [4-1:0] node2013;
	wire [4-1:0] node2014;
	wire [4-1:0] node2017;
	wire [4-1:0] node2019;
	wire [4-1:0] node2022;
	wire [4-1:0] node2023;
	wire [4-1:0] node2024;
	wire [4-1:0] node2025;
	wire [4-1:0] node2027;
	wire [4-1:0] node2030;
	wire [4-1:0] node2031;
	wire [4-1:0] node2034;
	wire [4-1:0] node2037;
	wire [4-1:0] node2039;
	wire [4-1:0] node2040;
	wire [4-1:0] node2044;
	wire [4-1:0] node2045;
	wire [4-1:0] node2047;
	wire [4-1:0] node2050;
	wire [4-1:0] node2052;
	wire [4-1:0] node2054;
	wire [4-1:0] node2057;
	wire [4-1:0] node2058;
	wire [4-1:0] node2059;
	wire [4-1:0] node2060;
	wire [4-1:0] node2064;
	wire [4-1:0] node2065;
	wire [4-1:0] node2068;
	wire [4-1:0] node2070;
	wire [4-1:0] node2073;
	wire [4-1:0] node2074;
	wire [4-1:0] node2076;
	wire [4-1:0] node2077;
	wire [4-1:0] node2080;
	wire [4-1:0] node2083;
	wire [4-1:0] node2084;
	wire [4-1:0] node2087;
	wire [4-1:0] node2090;
	wire [4-1:0] node2091;
	wire [4-1:0] node2092;
	wire [4-1:0] node2093;
	wire [4-1:0] node2094;
	wire [4-1:0] node2095;
	wire [4-1:0] node2096;
	wire [4-1:0] node2097;
	wire [4-1:0] node2099;
	wire [4-1:0] node2102;
	wire [4-1:0] node2103;
	wire [4-1:0] node2104;
	wire [4-1:0] node2109;
	wire [4-1:0] node2110;
	wire [4-1:0] node2112;
	wire [4-1:0] node2115;
	wire [4-1:0] node2118;
	wire [4-1:0] node2119;
	wire [4-1:0] node2121;
	wire [4-1:0] node2124;
	wire [4-1:0] node2125;
	wire [4-1:0] node2126;
	wire [4-1:0] node2127;
	wire [4-1:0] node2131;
	wire [4-1:0] node2134;
	wire [4-1:0] node2136;
	wire [4-1:0] node2139;
	wire [4-1:0] node2140;
	wire [4-1:0] node2141;
	wire [4-1:0] node2142;
	wire [4-1:0] node2143;
	wire [4-1:0] node2144;
	wire [4-1:0] node2149;
	wire [4-1:0] node2152;
	wire [4-1:0] node2153;
	wire [4-1:0] node2157;
	wire [4-1:0] node2159;
	wire [4-1:0] node2161;
	wire [4-1:0] node2162;
	wire [4-1:0] node2165;
	wire [4-1:0] node2168;
	wire [4-1:0] node2169;
	wire [4-1:0] node2170;
	wire [4-1:0] node2171;
	wire [4-1:0] node2172;
	wire [4-1:0] node2174;
	wire [4-1:0] node2178;
	wire [4-1:0] node2179;
	wire [4-1:0] node2181;
	wire [4-1:0] node2182;
	wire [4-1:0] node2185;
	wire [4-1:0] node2188;
	wire [4-1:0] node2189;
	wire [4-1:0] node2191;
	wire [4-1:0] node2194;
	wire [4-1:0] node2195;
	wire [4-1:0] node2199;
	wire [4-1:0] node2200;
	wire [4-1:0] node2201;
	wire [4-1:0] node2203;
	wire [4-1:0] node2206;
	wire [4-1:0] node2209;
	wire [4-1:0] node2210;
	wire [4-1:0] node2211;
	wire [4-1:0] node2215;
	wire [4-1:0] node2218;
	wire [4-1:0] node2219;
	wire [4-1:0] node2220;
	wire [4-1:0] node2222;
	wire [4-1:0] node2223;
	wire [4-1:0] node2226;
	wire [4-1:0] node2229;
	wire [4-1:0] node2230;
	wire [4-1:0] node2231;
	wire [4-1:0] node2235;
	wire [4-1:0] node2236;
	wire [4-1:0] node2240;
	wire [4-1:0] node2241;
	wire [4-1:0] node2242;
	wire [4-1:0] node2245;
	wire [4-1:0] node2247;
	wire [4-1:0] node2251;
	wire [4-1:0] node2252;
	wire [4-1:0] node2253;
	wire [4-1:0] node2254;
	wire [4-1:0] node2255;
	wire [4-1:0] node2256;
	wire [4-1:0] node2257;
	wire [4-1:0] node2261;
	wire [4-1:0] node2262;
	wire [4-1:0] node2264;
	wire [4-1:0] node2268;
	wire [4-1:0] node2271;
	wire [4-1:0] node2272;
	wire [4-1:0] node2273;
	wire [4-1:0] node2274;
	wire [4-1:0] node2275;
	wire [4-1:0] node2280;
	wire [4-1:0] node2281;
	wire [4-1:0] node2284;
	wire [4-1:0] node2285;
	wire [4-1:0] node2289;
	wire [4-1:0] node2290;
	wire [4-1:0] node2291;
	wire [4-1:0] node2295;
	wire [4-1:0] node2296;
	wire [4-1:0] node2300;
	wire [4-1:0] node2301;
	wire [4-1:0] node2302;
	wire [4-1:0] node2303;
	wire [4-1:0] node2306;
	wire [4-1:0] node2307;
	wire [4-1:0] node2310;
	wire [4-1:0] node2313;
	wire [4-1:0] node2315;
	wire [4-1:0] node2316;
	wire [4-1:0] node2319;
	wire [4-1:0] node2322;
	wire [4-1:0] node2323;
	wire [4-1:0] node2324;
	wire [4-1:0] node2326;
	wire [4-1:0] node2327;
	wire [4-1:0] node2330;
	wire [4-1:0] node2333;
	wire [4-1:0] node2334;
	wire [4-1:0] node2337;
	wire [4-1:0] node2340;
	wire [4-1:0] node2341;
	wire [4-1:0] node2345;
	wire [4-1:0] node2346;
	wire [4-1:0] node2347;
	wire [4-1:0] node2348;
	wire [4-1:0] node2349;
	wire [4-1:0] node2351;
	wire [4-1:0] node2352;
	wire [4-1:0] node2355;
	wire [4-1:0] node2358;
	wire [4-1:0] node2359;
	wire [4-1:0] node2363;
	wire [4-1:0] node2364;
	wire [4-1:0] node2365;
	wire [4-1:0] node2366;
	wire [4-1:0] node2369;
	wire [4-1:0] node2372;
	wire [4-1:0] node2375;
	wire [4-1:0] node2376;
	wire [4-1:0] node2379;
	wire [4-1:0] node2382;
	wire [4-1:0] node2383;
	wire [4-1:0] node2384;
	wire [4-1:0] node2385;
	wire [4-1:0] node2388;
	wire [4-1:0] node2391;
	wire [4-1:0] node2392;
	wire [4-1:0] node2395;
	wire [4-1:0] node2398;
	wire [4-1:0] node2399;
	wire [4-1:0] node2400;
	wire [4-1:0] node2404;
	wire [4-1:0] node2405;
	wire [4-1:0] node2406;
	wire [4-1:0] node2409;
	wire [4-1:0] node2412;
	wire [4-1:0] node2415;
	wire [4-1:0] node2416;
	wire [4-1:0] node2417;
	wire [4-1:0] node2418;
	wire [4-1:0] node2421;
	wire [4-1:0] node2424;
	wire [4-1:0] node2425;
	wire [4-1:0] node2426;
	wire [4-1:0] node2428;
	wire [4-1:0] node2432;
	wire [4-1:0] node2433;
	wire [4-1:0] node2435;
	wire [4-1:0] node2438;
	wire [4-1:0] node2441;
	wire [4-1:0] node2442;
	wire [4-1:0] node2444;
	wire [4-1:0] node2446;
	wire [4-1:0] node2449;
	wire [4-1:0] node2450;
	wire [4-1:0] node2453;
	wire [4-1:0] node2455;
	wire [4-1:0] node2458;
	wire [4-1:0] node2459;
	wire [4-1:0] node2460;
	wire [4-1:0] node2461;
	wire [4-1:0] node2462;
	wire [4-1:0] node2463;
	wire [4-1:0] node2465;
	wire [4-1:0] node2468;
	wire [4-1:0] node2469;
	wire [4-1:0] node2470;
	wire [4-1:0] node2471;
	wire [4-1:0] node2474;
	wire [4-1:0] node2477;
	wire [4-1:0] node2478;
	wire [4-1:0] node2481;
	wire [4-1:0] node2484;
	wire [4-1:0] node2485;
	wire [4-1:0] node2486;
	wire [4-1:0] node2491;
	wire [4-1:0] node2492;
	wire [4-1:0] node2493;
	wire [4-1:0] node2495;
	wire [4-1:0] node2497;
	wire [4-1:0] node2500;
	wire [4-1:0] node2502;
	wire [4-1:0] node2504;
	wire [4-1:0] node2507;
	wire [4-1:0] node2508;
	wire [4-1:0] node2509;
	wire [4-1:0] node2512;
	wire [4-1:0] node2515;
	wire [4-1:0] node2518;
	wire [4-1:0] node2519;
	wire [4-1:0] node2520;
	wire [4-1:0] node2521;
	wire [4-1:0] node2523;
	wire [4-1:0] node2526;
	wire [4-1:0] node2527;
	wire [4-1:0] node2530;
	wire [4-1:0] node2533;
	wire [4-1:0] node2535;
	wire [4-1:0] node2536;
	wire [4-1:0] node2537;
	wire [4-1:0] node2540;
	wire [4-1:0] node2543;
	wire [4-1:0] node2545;
	wire [4-1:0] node2548;
	wire [4-1:0] node2549;
	wire [4-1:0] node2550;
	wire [4-1:0] node2551;
	wire [4-1:0] node2555;
	wire [4-1:0] node2556;
	wire [4-1:0] node2559;
	wire [4-1:0] node2562;
	wire [4-1:0] node2563;
	wire [4-1:0] node2564;
	wire [4-1:0] node2565;
	wire [4-1:0] node2570;
	wire [4-1:0] node2571;
	wire [4-1:0] node2572;
	wire [4-1:0] node2577;
	wire [4-1:0] node2578;
	wire [4-1:0] node2579;
	wire [4-1:0] node2580;
	wire [4-1:0] node2581;
	wire [4-1:0] node2583;
	wire [4-1:0] node2586;
	wire [4-1:0] node2587;
	wire [4-1:0] node2589;
	wire [4-1:0] node2593;
	wire [4-1:0] node2594;
	wire [4-1:0] node2596;
	wire [4-1:0] node2597;
	wire [4-1:0] node2601;
	wire [4-1:0] node2602;
	wire [4-1:0] node2606;
	wire [4-1:0] node2607;
	wire [4-1:0] node2608;
	wire [4-1:0] node2609;
	wire [4-1:0] node2610;
	wire [4-1:0] node2613;
	wire [4-1:0] node2616;
	wire [4-1:0] node2620;
	wire [4-1:0] node2622;
	wire [4-1:0] node2623;
	wire [4-1:0] node2626;
	wire [4-1:0] node2629;
	wire [4-1:0] node2630;
	wire [4-1:0] node2631;
	wire [4-1:0] node2633;
	wire [4-1:0] node2634;
	wire [4-1:0] node2637;
	wire [4-1:0] node2639;
	wire [4-1:0] node2642;
	wire [4-1:0] node2643;
	wire [4-1:0] node2646;
	wire [4-1:0] node2649;
	wire [4-1:0] node2650;
	wire [4-1:0] node2651;
	wire [4-1:0] node2655;
	wire [4-1:0] node2656;
	wire [4-1:0] node2659;
	wire [4-1:0] node2660;
	wire [4-1:0] node2663;
	wire [4-1:0] node2664;
	wire [4-1:0] node2668;
	wire [4-1:0] node2669;
	wire [4-1:0] node2670;
	wire [4-1:0] node2671;
	wire [4-1:0] node2672;
	wire [4-1:0] node2673;
	wire [4-1:0] node2674;
	wire [4-1:0] node2675;
	wire [4-1:0] node2680;
	wire [4-1:0] node2681;
	wire [4-1:0] node2682;
	wire [4-1:0] node2686;
	wire [4-1:0] node2689;
	wire [4-1:0] node2691;
	wire [4-1:0] node2694;
	wire [4-1:0] node2695;
	wire [4-1:0] node2697;
	wire [4-1:0] node2698;
	wire [4-1:0] node2701;
	wire [4-1:0] node2704;
	wire [4-1:0] node2707;
	wire [4-1:0] node2708;
	wire [4-1:0] node2709;
	wire [4-1:0] node2710;
	wire [4-1:0] node2713;
	wire [4-1:0] node2716;
	wire [4-1:0] node2719;
	wire [4-1:0] node2720;
	wire [4-1:0] node2721;
	wire [4-1:0] node2724;
	wire [4-1:0] node2725;
	wire [4-1:0] node2727;
	wire [4-1:0] node2731;
	wire [4-1:0] node2733;
	wire [4-1:0] node2736;
	wire [4-1:0] node2737;
	wire [4-1:0] node2738;
	wire [4-1:0] node2739;
	wire [4-1:0] node2740;
	wire [4-1:0] node2742;
	wire [4-1:0] node2745;
	wire [4-1:0] node2747;
	wire [4-1:0] node2750;
	wire [4-1:0] node2752;
	wire [4-1:0] node2753;
	wire [4-1:0] node2757;
	wire [4-1:0] node2758;
	wire [4-1:0] node2760;
	wire [4-1:0] node2763;
	wire [4-1:0] node2764;
	wire [4-1:0] node2765;
	wire [4-1:0] node2768;
	wire [4-1:0] node2769;
	wire [4-1:0] node2773;
	wire [4-1:0] node2776;
	wire [4-1:0] node2777;
	wire [4-1:0] node2778;
	wire [4-1:0] node2779;
	wire [4-1:0] node2782;
	wire [4-1:0] node2783;
	wire [4-1:0] node2784;
	wire [4-1:0] node2788;
	wire [4-1:0] node2791;
	wire [4-1:0] node2793;
	wire [4-1:0] node2795;
	wire [4-1:0] node2796;
	wire [4-1:0] node2800;
	wire [4-1:0] node2801;
	wire [4-1:0] node2802;
	wire [4-1:0] node2803;
	wire [4-1:0] node2804;
	wire [4-1:0] node2810;
	wire [4-1:0] node2811;
	wire [4-1:0] node2812;
	wire [4-1:0] node2813;
	wire [4-1:0] node2817;
	wire [4-1:0] node2820;
	wire [4-1:0] node2823;
	wire [4-1:0] node2824;
	wire [4-1:0] node2825;
	wire [4-1:0] node2826;
	wire [4-1:0] node2827;
	wire [4-1:0] node2828;
	wire [4-1:0] node2829;
	wire [4-1:0] node2830;
	wire [4-1:0] node2831;
	wire [4-1:0] node2833;
	wire [4-1:0] node2836;
	wire [4-1:0] node2839;
	wire [4-1:0] node2840;
	wire [4-1:0] node2841;
	wire [4-1:0] node2843;
	wire [4-1:0] node2844;
	wire [4-1:0] node2849;
	wire [4-1:0] node2851;
	wire [4-1:0] node2854;
	wire [4-1:0] node2855;
	wire [4-1:0] node2856;
	wire [4-1:0] node2857;
	wire [4-1:0] node2859;
	wire [4-1:0] node2863;
	wire [4-1:0] node2864;
	wire [4-1:0] node2865;
	wire [4-1:0] node2870;
	wire [4-1:0] node2871;
	wire [4-1:0] node2872;
	wire [4-1:0] node2873;
	wire [4-1:0] node2876;
	wire [4-1:0] node2879;
	wire [4-1:0] node2882;
	wire [4-1:0] node2883;
	wire [4-1:0] node2884;
	wire [4-1:0] node2888;
	wire [4-1:0] node2889;
	wire [4-1:0] node2893;
	wire [4-1:0] node2894;
	wire [4-1:0] node2895;
	wire [4-1:0] node2896;
	wire [4-1:0] node2897;
	wire [4-1:0] node2899;
	wire [4-1:0] node2902;
	wire [4-1:0] node2903;
	wire [4-1:0] node2904;
	wire [4-1:0] node2907;
	wire [4-1:0] node2910;
	wire [4-1:0] node2913;
	wire [4-1:0] node2914;
	wire [4-1:0] node2917;
	wire [4-1:0] node2919;
	wire [4-1:0] node2922;
	wire [4-1:0] node2923;
	wire [4-1:0] node2925;
	wire [4-1:0] node2926;
	wire [4-1:0] node2927;
	wire [4-1:0] node2932;
	wire [4-1:0] node2933;
	wire [4-1:0] node2934;
	wire [4-1:0] node2937;
	wire [4-1:0] node2940;
	wire [4-1:0] node2943;
	wire [4-1:0] node2944;
	wire [4-1:0] node2945;
	wire [4-1:0] node2946;
	wire [4-1:0] node2948;
	wire [4-1:0] node2951;
	wire [4-1:0] node2952;
	wire [4-1:0] node2956;
	wire [4-1:0] node2957;
	wire [4-1:0] node2958;
	wire [4-1:0] node2960;
	wire [4-1:0] node2964;
	wire [4-1:0] node2967;
	wire [4-1:0] node2968;
	wire [4-1:0] node2969;
	wire [4-1:0] node2972;
	wire [4-1:0] node2974;
	wire [4-1:0] node2976;
	wire [4-1:0] node2979;
	wire [4-1:0] node2980;
	wire [4-1:0] node2983;
	wire [4-1:0] node2984;
	wire [4-1:0] node2988;
	wire [4-1:0] node2989;
	wire [4-1:0] node2990;
	wire [4-1:0] node2991;
	wire [4-1:0] node2992;
	wire [4-1:0] node2993;
	wire [4-1:0] node2994;
	wire [4-1:0] node2996;
	wire [4-1:0] node3000;
	wire [4-1:0] node3001;
	wire [4-1:0] node3004;
	wire [4-1:0] node3007;
	wire [4-1:0] node3008;
	wire [4-1:0] node3012;
	wire [4-1:0] node3013;
	wire [4-1:0] node3014;
	wire [4-1:0] node3017;
	wire [4-1:0] node3020;
	wire [4-1:0] node3021;
	wire [4-1:0] node3023;
	wire [4-1:0] node3025;
	wire [4-1:0] node3028;
	wire [4-1:0] node3031;
	wire [4-1:0] node3032;
	wire [4-1:0] node3033;
	wire [4-1:0] node3036;
	wire [4-1:0] node3037;
	wire [4-1:0] node3038;
	wire [4-1:0] node3040;
	wire [4-1:0] node3043;
	wire [4-1:0] node3045;
	wire [4-1:0] node3049;
	wire [4-1:0] node3050;
	wire [4-1:0] node3051;
	wire [4-1:0] node3052;
	wire [4-1:0] node3053;
	wire [4-1:0] node3056;
	wire [4-1:0] node3059;
	wire [4-1:0] node3060;
	wire [4-1:0] node3064;
	wire [4-1:0] node3067;
	wire [4-1:0] node3068;
	wire [4-1:0] node3069;
	wire [4-1:0] node3073;
	wire [4-1:0] node3076;
	wire [4-1:0] node3077;
	wire [4-1:0] node3078;
	wire [4-1:0] node3079;
	wire [4-1:0] node3080;
	wire [4-1:0] node3083;
	wire [4-1:0] node3086;
	wire [4-1:0] node3088;
	wire [4-1:0] node3091;
	wire [4-1:0] node3092;
	wire [4-1:0] node3093;
	wire [4-1:0] node3095;
	wire [4-1:0] node3097;
	wire [4-1:0] node3101;
	wire [4-1:0] node3102;
	wire [4-1:0] node3104;
	wire [4-1:0] node3105;
	wire [4-1:0] node3110;
	wire [4-1:0] node3111;
	wire [4-1:0] node3112;
	wire [4-1:0] node3113;
	wire [4-1:0] node3115;
	wire [4-1:0] node3117;
	wire [4-1:0] node3120;
	wire [4-1:0] node3123;
	wire [4-1:0] node3125;
	wire [4-1:0] node3126;
	wire [4-1:0] node3130;
	wire [4-1:0] node3131;
	wire [4-1:0] node3132;
	wire [4-1:0] node3133;
	wire [4-1:0] node3137;
	wire [4-1:0] node3138;
	wire [4-1:0] node3142;
	wire [4-1:0] node3143;
	wire [4-1:0] node3146;
	wire [4-1:0] node3147;
	wire [4-1:0] node3148;
	wire [4-1:0] node3152;
	wire [4-1:0] node3155;
	wire [4-1:0] node3156;
	wire [4-1:0] node3157;
	wire [4-1:0] node3158;
	wire [4-1:0] node3159;
	wire [4-1:0] node3160;
	wire [4-1:0] node3162;
	wire [4-1:0] node3163;
	wire [4-1:0] node3165;
	wire [4-1:0] node3168;
	wire [4-1:0] node3169;
	wire [4-1:0] node3173;
	wire [4-1:0] node3174;
	wire [4-1:0] node3176;
	wire [4-1:0] node3178;
	wire [4-1:0] node3181;
	wire [4-1:0] node3184;
	wire [4-1:0] node3185;
	wire [4-1:0] node3186;
	wire [4-1:0] node3187;
	wire [4-1:0] node3190;
	wire [4-1:0] node3194;
	wire [4-1:0] node3195;
	wire [4-1:0] node3197;
	wire [4-1:0] node3200;
	wire [4-1:0] node3201;
	wire [4-1:0] node3204;
	wire [4-1:0] node3207;
	wire [4-1:0] node3208;
	wire [4-1:0] node3209;
	wire [4-1:0] node3210;
	wire [4-1:0] node3211;
	wire [4-1:0] node3212;
	wire [4-1:0] node3215;
	wire [4-1:0] node3218;
	wire [4-1:0] node3221;
	wire [4-1:0] node3222;
	wire [4-1:0] node3223;
	wire [4-1:0] node3228;
	wire [4-1:0] node3229;
	wire [4-1:0] node3232;
	wire [4-1:0] node3235;
	wire [4-1:0] node3236;
	wire [4-1:0] node3237;
	wire [4-1:0] node3239;
	wire [4-1:0] node3242;
	wire [4-1:0] node3245;
	wire [4-1:0] node3246;
	wire [4-1:0] node3248;
	wire [4-1:0] node3251;
	wire [4-1:0] node3252;
	wire [4-1:0] node3256;
	wire [4-1:0] node3257;
	wire [4-1:0] node3258;
	wire [4-1:0] node3259;
	wire [4-1:0] node3260;
	wire [4-1:0] node3261;
	wire [4-1:0] node3265;
	wire [4-1:0] node3266;
	wire [4-1:0] node3269;
	wire [4-1:0] node3271;
	wire [4-1:0] node3274;
	wire [4-1:0] node3275;
	wire [4-1:0] node3278;
	wire [4-1:0] node3279;
	wire [4-1:0] node3280;
	wire [4-1:0] node3283;
	wire [4-1:0] node3286;
	wire [4-1:0] node3287;
	wire [4-1:0] node3290;
	wire [4-1:0] node3293;
	wire [4-1:0] node3294;
	wire [4-1:0] node3295;
	wire [4-1:0] node3297;
	wire [4-1:0] node3301;
	wire [4-1:0] node3302;
	wire [4-1:0] node3303;
	wire [4-1:0] node3304;
	wire [4-1:0] node3309;
	wire [4-1:0] node3310;
	wire [4-1:0] node3312;
	wire [4-1:0] node3316;
	wire [4-1:0] node3317;
	wire [4-1:0] node3318;
	wire [4-1:0] node3319;
	wire [4-1:0] node3323;
	wire [4-1:0] node3324;
	wire [4-1:0] node3327;
	wire [4-1:0] node3328;
	wire [4-1:0] node3330;
	wire [4-1:0] node3333;
	wire [4-1:0] node3335;
	wire [4-1:0] node3338;
	wire [4-1:0] node3339;
	wire [4-1:0] node3341;
	wire [4-1:0] node3343;
	wire [4-1:0] node3346;
	wire [4-1:0] node3347;
	wire [4-1:0] node3348;
	wire [4-1:0] node3350;
	wire [4-1:0] node3353;
	wire [4-1:0] node3354;
	wire [4-1:0] node3358;
	wire [4-1:0] node3359;
	wire [4-1:0] node3361;
	wire [4-1:0] node3364;
	wire [4-1:0] node3367;
	wire [4-1:0] node3368;
	wire [4-1:0] node3369;
	wire [4-1:0] node3370;
	wire [4-1:0] node3371;
	wire [4-1:0] node3372;
	wire [4-1:0] node3373;
	wire [4-1:0] node3376;
	wire [4-1:0] node3380;
	wire [4-1:0] node3381;
	wire [4-1:0] node3384;
	wire [4-1:0] node3387;
	wire [4-1:0] node3388;
	wire [4-1:0] node3389;
	wire [4-1:0] node3390;
	wire [4-1:0] node3394;
	wire [4-1:0] node3395;
	wire [4-1:0] node3398;
	wire [4-1:0] node3401;
	wire [4-1:0] node3404;
	wire [4-1:0] node3405;
	wire [4-1:0] node3407;
	wire [4-1:0] node3408;
	wire [4-1:0] node3409;
	wire [4-1:0] node3412;
	wire [4-1:0] node3415;
	wire [4-1:0] node3417;
	wire [4-1:0] node3420;
	wire [4-1:0] node3421;
	wire [4-1:0] node3422;
	wire [4-1:0] node3424;
	wire [4-1:0] node3428;
	wire [4-1:0] node3429;
	wire [4-1:0] node3432;
	wire [4-1:0] node3435;
	wire [4-1:0] node3436;
	wire [4-1:0] node3437;
	wire [4-1:0] node3438;
	wire [4-1:0] node3439;
	wire [4-1:0] node3440;
	wire [4-1:0] node3442;
	wire [4-1:0] node3445;
	wire [4-1:0] node3449;
	wire [4-1:0] node3451;
	wire [4-1:0] node3452;
	wire [4-1:0] node3455;
	wire [4-1:0] node3458;
	wire [4-1:0] node3459;
	wire [4-1:0] node3460;
	wire [4-1:0] node3463;
	wire [4-1:0] node3465;
	wire [4-1:0] node3468;
	wire [4-1:0] node3469;
	wire [4-1:0] node3472;
	wire [4-1:0] node3475;
	wire [4-1:0] node3476;
	wire [4-1:0] node3477;
	wire [4-1:0] node3479;
	wire [4-1:0] node3480;
	wire [4-1:0] node3483;
	wire [4-1:0] node3484;
	wire [4-1:0] node3488;
	wire [4-1:0] node3489;
	wire [4-1:0] node3492;
	wire [4-1:0] node3493;
	wire [4-1:0] node3495;
	wire [4-1:0] node3499;
	wire [4-1:0] node3500;
	wire [4-1:0] node3501;
	wire [4-1:0] node3503;
	wire [4-1:0] node3506;
	wire [4-1:0] node3509;
	wire [4-1:0] node3511;
	wire [4-1:0] node3512;
	wire [4-1:0] node3515;
	wire [4-1:0] node3518;
	wire [4-1:0] node3519;
	wire [4-1:0] node3520;
	wire [4-1:0] node3521;
	wire [4-1:0] node3522;
	wire [4-1:0] node3523;
	wire [4-1:0] node3524;
	wire [4-1:0] node3525;
	wire [4-1:0] node3528;
	wire [4-1:0] node3530;
	wire [4-1:0] node3533;
	wire [4-1:0] node3534;
	wire [4-1:0] node3535;
	wire [4-1:0] node3537;
	wire [4-1:0] node3541;
	wire [4-1:0] node3542;
	wire [4-1:0] node3546;
	wire [4-1:0] node3547;
	wire [4-1:0] node3548;
	wire [4-1:0] node3549;
	wire [4-1:0] node3552;
	wire [4-1:0] node3553;
	wire [4-1:0] node3557;
	wire [4-1:0] node3559;
	wire [4-1:0] node3562;
	wire [4-1:0] node3563;
	wire [4-1:0] node3567;
	wire [4-1:0] node3568;
	wire [4-1:0] node3569;
	wire [4-1:0] node3571;
	wire [4-1:0] node3572;
	wire [4-1:0] node3574;
	wire [4-1:0] node3578;
	wire [4-1:0] node3579;
	wire [4-1:0] node3581;
	wire [4-1:0] node3582;
	wire [4-1:0] node3586;
	wire [4-1:0] node3587;
	wire [4-1:0] node3590;
	wire [4-1:0] node3591;
	wire [4-1:0] node3595;
	wire [4-1:0] node3596;
	wire [4-1:0] node3597;
	wire [4-1:0] node3601;
	wire [4-1:0] node3602;
	wire [4-1:0] node3604;
	wire [4-1:0] node3607;
	wire [4-1:0] node3610;
	wire [4-1:0] node3611;
	wire [4-1:0] node3612;
	wire [4-1:0] node3613;
	wire [4-1:0] node3615;
	wire [4-1:0] node3618;
	wire [4-1:0] node3619;
	wire [4-1:0] node3622;
	wire [4-1:0] node3625;
	wire [4-1:0] node3626;
	wire [4-1:0] node3627;
	wire [4-1:0] node3628;
	wire [4-1:0] node3629;
	wire [4-1:0] node3635;
	wire [4-1:0] node3637;
	wire [4-1:0] node3640;
	wire [4-1:0] node3641;
	wire [4-1:0] node3642;
	wire [4-1:0] node3644;
	wire [4-1:0] node3645;
	wire [4-1:0] node3648;
	wire [4-1:0] node3649;
	wire [4-1:0] node3652;
	wire [4-1:0] node3655;
	wire [4-1:0] node3656;
	wire [4-1:0] node3658;
	wire [4-1:0] node3659;
	wire [4-1:0] node3663;
	wire [4-1:0] node3664;
	wire [4-1:0] node3665;
	wire [4-1:0] node3669;
	wire [4-1:0] node3670;
	wire [4-1:0] node3674;
	wire [4-1:0] node3675;
	wire [4-1:0] node3676;
	wire [4-1:0] node3677;
	wire [4-1:0] node3680;
	wire [4-1:0] node3683;
	wire [4-1:0] node3684;
	wire [4-1:0] node3687;
	wire [4-1:0] node3690;
	wire [4-1:0] node3691;
	wire [4-1:0] node3692;
	wire [4-1:0] node3694;
	wire [4-1:0] node3697;
	wire [4-1:0] node3699;
	wire [4-1:0] node3702;
	wire [4-1:0] node3705;
	wire [4-1:0] node3706;
	wire [4-1:0] node3707;
	wire [4-1:0] node3708;
	wire [4-1:0] node3709;
	wire [4-1:0] node3711;
	wire [4-1:0] node3712;
	wire [4-1:0] node3715;
	wire [4-1:0] node3716;
	wire [4-1:0] node3720;
	wire [4-1:0] node3721;
	wire [4-1:0] node3722;
	wire [4-1:0] node3724;
	wire [4-1:0] node3728;
	wire [4-1:0] node3729;
	wire [4-1:0] node3731;
	wire [4-1:0] node3734;
	wire [4-1:0] node3737;
	wire [4-1:0] node3738;
	wire [4-1:0] node3739;
	wire [4-1:0] node3740;
	wire [4-1:0] node3743;
	wire [4-1:0] node3747;
	wire [4-1:0] node3749;
	wire [4-1:0] node3752;
	wire [4-1:0] node3753;
	wire [4-1:0] node3754;
	wire [4-1:0] node3755;
	wire [4-1:0] node3756;
	wire [4-1:0] node3758;
	wire [4-1:0] node3761;
	wire [4-1:0] node3764;
	wire [4-1:0] node3766;
	wire [4-1:0] node3769;
	wire [4-1:0] node3770;
	wire [4-1:0] node3771;
	wire [4-1:0] node3774;
	wire [4-1:0] node3777;
	wire [4-1:0] node3779;
	wire [4-1:0] node3782;
	wire [4-1:0] node3783;
	wire [4-1:0] node3784;
	wire [4-1:0] node3786;
	wire [4-1:0] node3789;
	wire [4-1:0] node3791;
	wire [4-1:0] node3792;
	wire [4-1:0] node3796;
	wire [4-1:0] node3797;
	wire [4-1:0] node3801;
	wire [4-1:0] node3802;
	wire [4-1:0] node3803;
	wire [4-1:0] node3804;
	wire [4-1:0] node3805;
	wire [4-1:0] node3808;
	wire [4-1:0] node3809;
	wire [4-1:0] node3813;
	wire [4-1:0] node3814;
	wire [4-1:0] node3815;
	wire [4-1:0] node3819;
	wire [4-1:0] node3822;
	wire [4-1:0] node3823;
	wire [4-1:0] node3824;
	wire [4-1:0] node3825;
	wire [4-1:0] node3828;
	wire [4-1:0] node3831;
	wire [4-1:0] node3833;
	wire [4-1:0] node3836;
	wire [4-1:0] node3837;
	wire [4-1:0] node3839;
	wire [4-1:0] node3841;
	wire [4-1:0] node3844;
	wire [4-1:0] node3846;
	wire [4-1:0] node3847;
	wire [4-1:0] node3851;
	wire [4-1:0] node3852;
	wire [4-1:0] node3853;
	wire [4-1:0] node3854;
	wire [4-1:0] node3858;
	wire [4-1:0] node3859;
	wire [4-1:0] node3860;
	wire [4-1:0] node3864;
	wire [4-1:0] node3866;
	wire [4-1:0] node3868;
	wire [4-1:0] node3871;
	wire [4-1:0] node3872;
	wire [4-1:0] node3873;
	wire [4-1:0] node3875;
	wire [4-1:0] node3878;
	wire [4-1:0] node3880;
	wire [4-1:0] node3881;
	wire [4-1:0] node3884;
	wire [4-1:0] node3887;
	wire [4-1:0] node3888;
	wire [4-1:0] node3889;
	wire [4-1:0] node3893;
	wire [4-1:0] node3895;
	wire [4-1:0] node3898;
	wire [4-1:0] node3899;
	wire [4-1:0] node3900;
	wire [4-1:0] node3901;
	wire [4-1:0] node3902;
	wire [4-1:0] node3903;
	wire [4-1:0] node3904;
	wire [4-1:0] node3905;
	wire [4-1:0] node3908;
	wire [4-1:0] node3911;
	wire [4-1:0] node3912;
	wire [4-1:0] node3914;
	wire [4-1:0] node3917;
	wire [4-1:0] node3920;
	wire [4-1:0] node3921;
	wire [4-1:0] node3924;
	wire [4-1:0] node3927;
	wire [4-1:0] node3928;
	wire [4-1:0] node3929;
	wire [4-1:0] node3931;
	wire [4-1:0] node3934;
	wire [4-1:0] node3935;
	wire [4-1:0] node3939;
	wire [4-1:0] node3940;
	wire [4-1:0] node3941;
	wire [4-1:0] node3945;
	wire [4-1:0] node3948;
	wire [4-1:0] node3949;
	wire [4-1:0] node3950;
	wire [4-1:0] node3952;
	wire [4-1:0] node3953;
	wire [4-1:0] node3954;
	wire [4-1:0] node3959;
	wire [4-1:0] node3961;
	wire [4-1:0] node3964;
	wire [4-1:0] node3965;
	wire [4-1:0] node3966;
	wire [4-1:0] node3969;
	wire [4-1:0] node3971;
	wire [4-1:0] node3972;
	wire [4-1:0] node3976;
	wire [4-1:0] node3977;
	wire [4-1:0] node3981;
	wire [4-1:0] node3982;
	wire [4-1:0] node3983;
	wire [4-1:0] node3984;
	wire [4-1:0] node3985;
	wire [4-1:0] node3986;
	wire [4-1:0] node3989;
	wire [4-1:0] node3990;
	wire [4-1:0] node3994;
	wire [4-1:0] node3997;
	wire [4-1:0] node3998;
	wire [4-1:0] node3999;
	wire [4-1:0] node4000;
	wire [4-1:0] node4004;
	wire [4-1:0] node4005;
	wire [4-1:0] node4010;
	wire [4-1:0] node4011;
	wire [4-1:0] node4013;
	wire [4-1:0] node4016;
	wire [4-1:0] node4018;
	wire [4-1:0] node4020;
	wire [4-1:0] node4023;
	wire [4-1:0] node4024;
	wire [4-1:0] node4025;
	wire [4-1:0] node4026;
	wire [4-1:0] node4028;
	wire [4-1:0] node4031;
	wire [4-1:0] node4034;
	wire [4-1:0] node4035;
	wire [4-1:0] node4037;
	wire [4-1:0] node4040;
	wire [4-1:0] node4041;
	wire [4-1:0] node4044;
	wire [4-1:0] node4046;
	wire [4-1:0] node4049;
	wire [4-1:0] node4050;
	wire [4-1:0] node4051;
	wire [4-1:0] node4053;
	wire [4-1:0] node4056;
	wire [4-1:0] node4057;
	wire [4-1:0] node4061;
	wire [4-1:0] node4062;
	wire [4-1:0] node4065;
	wire [4-1:0] node4066;
	wire [4-1:0] node4070;
	wire [4-1:0] node4071;
	wire [4-1:0] node4072;
	wire [4-1:0] node4073;
	wire [4-1:0] node4074;
	wire [4-1:0] node4075;
	wire [4-1:0] node4078;
	wire [4-1:0] node4079;
	wire [4-1:0] node4083;
	wire [4-1:0] node4084;
	wire [4-1:0] node4085;
	wire [4-1:0] node4086;
	wire [4-1:0] node4089;
	wire [4-1:0] node4092;
	wire [4-1:0] node4094;
	wire [4-1:0] node4097;
	wire [4-1:0] node4098;
	wire [4-1:0] node4100;
	wire [4-1:0] node4103;
	wire [4-1:0] node4106;
	wire [4-1:0] node4107;
	wire [4-1:0] node4108;
	wire [4-1:0] node4111;
	wire [4-1:0] node4114;
	wire [4-1:0] node4116;
	wire [4-1:0] node4119;
	wire [4-1:0] node4120;
	wire [4-1:0] node4121;
	wire [4-1:0] node4122;
	wire [4-1:0] node4126;
	wire [4-1:0] node4127;
	wire [4-1:0] node4128;
	wire [4-1:0] node4129;
	wire [4-1:0] node4134;
	wire [4-1:0] node4135;
	wire [4-1:0] node4139;
	wire [4-1:0] node4140;
	wire [4-1:0] node4142;
	wire [4-1:0] node4145;
	wire [4-1:0] node4146;
	wire [4-1:0] node4147;
	wire [4-1:0] node4148;
	wire [4-1:0] node4154;
	wire [4-1:0] node4155;
	wire [4-1:0] node4156;
	wire [4-1:0] node4157;
	wire [4-1:0] node4158;
	wire [4-1:0] node4161;
	wire [4-1:0] node4163;
	wire [4-1:0] node4166;
	wire [4-1:0] node4167;
	wire [4-1:0] node4168;
	wire [4-1:0] node4171;
	wire [4-1:0] node4172;
	wire [4-1:0] node4177;
	wire [4-1:0] node4178;
	wire [4-1:0] node4179;
	wire [4-1:0] node4180;
	wire [4-1:0] node4183;
	wire [4-1:0] node4186;
	wire [4-1:0] node4187;
	wire [4-1:0] node4190;
	wire [4-1:0] node4193;
	wire [4-1:0] node4195;
	wire [4-1:0] node4198;
	wire [4-1:0] node4199;
	wire [4-1:0] node4200;
	wire [4-1:0] node4201;
	wire [4-1:0] node4202;
	wire [4-1:0] node4204;
	wire [4-1:0] node4207;
	wire [4-1:0] node4209;
	wire [4-1:0] node4212;
	wire [4-1:0] node4213;
	wire [4-1:0] node4217;
	wire [4-1:0] node4218;
	wire [4-1:0] node4221;
	wire [4-1:0] node4224;
	wire [4-1:0] node4225;
	wire [4-1:0] node4226;
	wire [4-1:0] node4227;
	wire [4-1:0] node4231;
	wire [4-1:0] node4232;
	wire [4-1:0] node4235;
	wire [4-1:0] node4238;
	wire [4-1:0] node4239;
	wire [4-1:0] node4240;
	wire [4-1:0] node4242;
	wire [4-1:0] node4245;
	wire [4-1:0] node4247;
	wire [4-1:0] node4250;
	wire [4-1:0] node4252;
	wire [4-1:0] node4255;
	wire [4-1:0] node4256;
	wire [4-1:0] node4257;
	wire [4-1:0] node4258;
	wire [4-1:0] node4259;
	wire [4-1:0] node4260;
	wire [4-1:0] node4261;
	wire [4-1:0] node4262;
	wire [4-1:0] node4263;
	wire [4-1:0] node4266;
	wire [4-1:0] node4268;
	wire [4-1:0] node4271;
	wire [4-1:0] node4272;
	wire [4-1:0] node4273;
	wire [4-1:0] node4275;
	wire [4-1:0] node4278;
	wire [4-1:0] node4281;
	wire [4-1:0] node4284;
	wire [4-1:0] node4285;
	wire [4-1:0] node4286;
	wire [4-1:0] node4287;
	wire [4-1:0] node4291;
	wire [4-1:0] node4292;
	wire [4-1:0] node4295;
	wire [4-1:0] node4298;
	wire [4-1:0] node4299;
	wire [4-1:0] node4301;
	wire [4-1:0] node4302;
	wire [4-1:0] node4306;
	wire [4-1:0] node4309;
	wire [4-1:0] node4310;
	wire [4-1:0] node4311;
	wire [4-1:0] node4313;
	wire [4-1:0] node4316;
	wire [4-1:0] node4317;
	wire [4-1:0] node4318;
	wire [4-1:0] node4321;
	wire [4-1:0] node4325;
	wire [4-1:0] node4326;
	wire [4-1:0] node4327;
	wire [4-1:0] node4328;
	wire [4-1:0] node4330;
	wire [4-1:0] node4334;
	wire [4-1:0] node4335;
	wire [4-1:0] node4336;
	wire [4-1:0] node4341;
	wire [4-1:0] node4343;
	wire [4-1:0] node4344;
	wire [4-1:0] node4345;
	wire [4-1:0] node4350;
	wire [4-1:0] node4351;
	wire [4-1:0] node4352;
	wire [4-1:0] node4353;
	wire [4-1:0] node4354;
	wire [4-1:0] node4357;
	wire [4-1:0] node4359;
	wire [4-1:0] node4362;
	wire [4-1:0] node4363;
	wire [4-1:0] node4365;
	wire [4-1:0] node4369;
	wire [4-1:0] node4370;
	wire [4-1:0] node4372;
	wire [4-1:0] node4375;
	wire [4-1:0] node4376;
	wire [4-1:0] node4378;
	wire [4-1:0] node4379;
	wire [4-1:0] node4382;
	wire [4-1:0] node4385;
	wire [4-1:0] node4386;
	wire [4-1:0] node4389;
	wire [4-1:0] node4392;
	wire [4-1:0] node4393;
	wire [4-1:0] node4394;
	wire [4-1:0] node4396;
	wire [4-1:0] node4397;
	wire [4-1:0] node4398;
	wire [4-1:0] node4401;
	wire [4-1:0] node4405;
	wire [4-1:0] node4406;
	wire [4-1:0] node4407;
	wire [4-1:0] node4411;
	wire [4-1:0] node4412;
	wire [4-1:0] node4413;
	wire [4-1:0] node4418;
	wire [4-1:0] node4419;
	wire [4-1:0] node4420;
	wire [4-1:0] node4421;
	wire [4-1:0] node4425;
	wire [4-1:0] node4427;
	wire [4-1:0] node4430;
	wire [4-1:0] node4431;
	wire [4-1:0] node4434;
	wire [4-1:0] node4437;
	wire [4-1:0] node4438;
	wire [4-1:0] node4439;
	wire [4-1:0] node4440;
	wire [4-1:0] node4441;
	wire [4-1:0] node4442;
	wire [4-1:0] node4445;
	wire [4-1:0] node4446;
	wire [4-1:0] node4450;
	wire [4-1:0] node4452;
	wire [4-1:0] node4453;
	wire [4-1:0] node4457;
	wire [4-1:0] node4458;
	wire [4-1:0] node4459;
	wire [4-1:0] node4460;
	wire [4-1:0] node4462;
	wire [4-1:0] node4465;
	wire [4-1:0] node4468;
	wire [4-1:0] node4469;
	wire [4-1:0] node4470;
	wire [4-1:0] node4473;
	wire [4-1:0] node4476;
	wire [4-1:0] node4478;
	wire [4-1:0] node4481;
	wire [4-1:0] node4482;
	wire [4-1:0] node4485;
	wire [4-1:0] node4487;
	wire [4-1:0] node4490;
	wire [4-1:0] node4491;
	wire [4-1:0] node4492;
	wire [4-1:0] node4494;
	wire [4-1:0] node4495;
	wire [4-1:0] node4496;
	wire [4-1:0] node4501;
	wire [4-1:0] node4502;
	wire [4-1:0] node4503;
	wire [4-1:0] node4507;
	wire [4-1:0] node4508;
	wire [4-1:0] node4511;
	wire [4-1:0] node4512;
	wire [4-1:0] node4516;
	wire [4-1:0] node4517;
	wire [4-1:0] node4519;
	wire [4-1:0] node4522;
	wire [4-1:0] node4523;
	wire [4-1:0] node4524;
	wire [4-1:0] node4526;
	wire [4-1:0] node4529;
	wire [4-1:0] node4532;
	wire [4-1:0] node4533;
	wire [4-1:0] node4537;
	wire [4-1:0] node4538;
	wire [4-1:0] node4539;
	wire [4-1:0] node4540;
	wire [4-1:0] node4541;
	wire [4-1:0] node4542;
	wire [4-1:0] node4543;
	wire [4-1:0] node4547;
	wire [4-1:0] node4549;
	wire [4-1:0] node4552;
	wire [4-1:0] node4555;
	wire [4-1:0] node4556;
	wire [4-1:0] node4558;
	wire [4-1:0] node4561;
	wire [4-1:0] node4563;
	wire [4-1:0] node4566;
	wire [4-1:0] node4567;
	wire [4-1:0] node4568;
	wire [4-1:0] node4570;
	wire [4-1:0] node4572;
	wire [4-1:0] node4575;
	wire [4-1:0] node4578;
	wire [4-1:0] node4579;
	wire [4-1:0] node4582;
	wire [4-1:0] node4583;
	wire [4-1:0] node4587;
	wire [4-1:0] node4588;
	wire [4-1:0] node4589;
	wire [4-1:0] node4590;
	wire [4-1:0] node4593;
	wire [4-1:0] node4594;
	wire [4-1:0] node4598;
	wire [4-1:0] node4599;
	wire [4-1:0] node4600;
	wire [4-1:0] node4602;
	wire [4-1:0] node4606;
	wire [4-1:0] node4608;
	wire [4-1:0] node4611;
	wire [4-1:0] node4612;
	wire [4-1:0] node4613;
	wire [4-1:0] node4614;
	wire [4-1:0] node4618;
	wire [4-1:0] node4619;
	wire [4-1:0] node4623;
	wire [4-1:0] node4624;
	wire [4-1:0] node4626;
	wire [4-1:0] node4629;
	wire [4-1:0] node4630;
	wire [4-1:0] node4632;
	wire [4-1:0] node4636;
	wire [4-1:0] node4637;
	wire [4-1:0] node4638;
	wire [4-1:0] node4639;
	wire [4-1:0] node4640;
	wire [4-1:0] node4641;
	wire [4-1:0] node4642;
	wire [4-1:0] node4643;
	wire [4-1:0] node4648;
	wire [4-1:0] node4651;
	wire [4-1:0] node4652;
	wire [4-1:0] node4653;
	wire [4-1:0] node4654;
	wire [4-1:0] node4658;
	wire [4-1:0] node4661;
	wire [4-1:0] node4662;
	wire [4-1:0] node4663;
	wire [4-1:0] node4667;
	wire [4-1:0] node4670;
	wire [4-1:0] node4671;
	wire [4-1:0] node4672;
	wire [4-1:0] node4673;
	wire [4-1:0] node4675;
	wire [4-1:0] node4678;
	wire [4-1:0] node4680;
	wire [4-1:0] node4682;
	wire [4-1:0] node4685;
	wire [4-1:0] node4687;
	wire [4-1:0] node4688;
	wire [4-1:0] node4691;
	wire [4-1:0] node4692;
	wire [4-1:0] node4696;
	wire [4-1:0] node4697;
	wire [4-1:0] node4698;
	wire [4-1:0] node4702;
	wire [4-1:0] node4703;
	wire [4-1:0] node4704;
	wire [4-1:0] node4706;
	wire [4-1:0] node4709;
	wire [4-1:0] node4712;
	wire [4-1:0] node4713;
	wire [4-1:0] node4716;
	wire [4-1:0] node4719;
	wire [4-1:0] node4720;
	wire [4-1:0] node4721;
	wire [4-1:0] node4722;
	wire [4-1:0] node4723;
	wire [4-1:0] node4724;
	wire [4-1:0] node4726;
	wire [4-1:0] node4730;
	wire [4-1:0] node4731;
	wire [4-1:0] node4734;
	wire [4-1:0] node4737;
	wire [4-1:0] node4738;
	wire [4-1:0] node4740;
	wire [4-1:0] node4741;
	wire [4-1:0] node4745;
	wire [4-1:0] node4748;
	wire [4-1:0] node4749;
	wire [4-1:0] node4750;
	wire [4-1:0] node4754;
	wire [4-1:0] node4755;
	wire [4-1:0] node4756;
	wire [4-1:0] node4757;
	wire [4-1:0] node4762;
	wire [4-1:0] node4765;
	wire [4-1:0] node4766;
	wire [4-1:0] node4767;
	wire [4-1:0] node4768;
	wire [4-1:0] node4770;
	wire [4-1:0] node4773;
	wire [4-1:0] node4774;
	wire [4-1:0] node4778;
	wire [4-1:0] node4779;
	wire [4-1:0] node4780;
	wire [4-1:0] node4781;
	wire [4-1:0] node4785;
	wire [4-1:0] node4788;
	wire [4-1:0] node4791;
	wire [4-1:0] node4792;
	wire [4-1:0] node4793;
	wire [4-1:0] node4794;
	wire [4-1:0] node4798;
	wire [4-1:0] node4799;
	wire [4-1:0] node4801;
	wire [4-1:0] node4805;
	wire [4-1:0] node4806;
	wire [4-1:0] node4808;
	wire [4-1:0] node4811;
	wire [4-1:0] node4813;
	wire [4-1:0] node4816;
	wire [4-1:0] node4817;
	wire [4-1:0] node4818;
	wire [4-1:0] node4819;
	wire [4-1:0] node4820;
	wire [4-1:0] node4821;
	wire [4-1:0] node4822;
	wire [4-1:0] node4823;
	wire [4-1:0] node4826;
	wire [4-1:0] node4829;
	wire [4-1:0] node4832;
	wire [4-1:0] node4833;
	wire [4-1:0] node4835;
	wire [4-1:0] node4839;
	wire [4-1:0] node4840;
	wire [4-1:0] node4841;
	wire [4-1:0] node4844;
	wire [4-1:0] node4848;
	wire [4-1:0] node4849;
	wire [4-1:0] node4850;
	wire [4-1:0] node4852;
	wire [4-1:0] node4854;
	wire [4-1:0] node4857;
	wire [4-1:0] node4860;
	wire [4-1:0] node4861;
	wire [4-1:0] node4862;
	wire [4-1:0] node4865;
	wire [4-1:0] node4867;
	wire [4-1:0] node4870;
	wire [4-1:0] node4873;
	wire [4-1:0] node4874;
	wire [4-1:0] node4875;
	wire [4-1:0] node4876;
	wire [4-1:0] node4879;
	wire [4-1:0] node4881;
	wire [4-1:0] node4883;
	wire [4-1:0] node4886;
	wire [4-1:0] node4887;
	wire [4-1:0] node4890;
	wire [4-1:0] node4893;
	wire [4-1:0] node4894;
	wire [4-1:0] node4895;
	wire [4-1:0] node4896;
	wire [4-1:0] node4900;
	wire [4-1:0] node4901;
	wire [4-1:0] node4902;
	wire [4-1:0] node4905;
	wire [4-1:0] node4908;
	wire [4-1:0] node4909;
	wire [4-1:0] node4913;
	wire [4-1:0] node4915;
	wire [4-1:0] node4916;
	wire [4-1:0] node4919;
	wire [4-1:0] node4921;
	wire [4-1:0] node4924;
	wire [4-1:0] node4925;
	wire [4-1:0] node4926;
	wire [4-1:0] node4927;
	wire [4-1:0] node4928;
	wire [4-1:0] node4930;
	wire [4-1:0] node4933;
	wire [4-1:0] node4935;
	wire [4-1:0] node4938;
	wire [4-1:0] node4941;
	wire [4-1:0] node4942;
	wire [4-1:0] node4943;
	wire [4-1:0] node4945;
	wire [4-1:0] node4948;
	wire [4-1:0] node4951;
	wire [4-1:0] node4952;
	wire [4-1:0] node4953;
	wire [4-1:0] node4954;
	wire [4-1:0] node4958;
	wire [4-1:0] node4959;
	wire [4-1:0] node4964;
	wire [4-1:0] node4965;
	wire [4-1:0] node4966;
	wire [4-1:0] node4967;
	wire [4-1:0] node4969;
	wire [4-1:0] node4970;
	wire [4-1:0] node4975;
	wire [4-1:0] node4976;
	wire [4-1:0] node4977;
	wire [4-1:0] node4981;
	wire [4-1:0] node4983;
	wire [4-1:0] node4986;
	wire [4-1:0] node4987;
	wire [4-1:0] node4988;
	wire [4-1:0] node4991;
	wire [4-1:0] node4992;
	wire [4-1:0] node4995;
	wire [4-1:0] node4996;
	wire [4-1:0] node5000;
	wire [4-1:0] node5001;
	wire [4-1:0] node5005;
	wire [4-1:0] node5006;
	wire [4-1:0] node5007;
	wire [4-1:0] node5008;
	wire [4-1:0] node5009;
	wire [4-1:0] node5010;
	wire [4-1:0] node5011;
	wire [4-1:0] node5012;
	wire [4-1:0] node5014;
	wire [4-1:0] node5017;
	wire [4-1:0] node5018;
	wire [4-1:0] node5020;
	wire [4-1:0] node5024;
	wire [4-1:0] node5025;
	wire [4-1:0] node5026;
	wire [4-1:0] node5030;
	wire [4-1:0] node5033;
	wire [4-1:0] node5034;
	wire [4-1:0] node5035;
	wire [4-1:0] node5039;
	wire [4-1:0] node5040;
	wire [4-1:0] node5043;
	wire [4-1:0] node5046;
	wire [4-1:0] node5047;
	wire [4-1:0] node5048;
	wire [4-1:0] node5050;
	wire [4-1:0] node5054;
	wire [4-1:0] node5055;
	wire [4-1:0] node5056;
	wire [4-1:0] node5057;
	wire [4-1:0] node5061;
	wire [4-1:0] node5063;
	wire [4-1:0] node5064;
	wire [4-1:0] node5068;
	wire [4-1:0] node5069;
	wire [4-1:0] node5071;
	wire [4-1:0] node5075;
	wire [4-1:0] node5076;
	wire [4-1:0] node5077;
	wire [4-1:0] node5078;
	wire [4-1:0] node5079;
	wire [4-1:0] node5082;
	wire [4-1:0] node5083;
	wire [4-1:0] node5087;
	wire [4-1:0] node5088;
	wire [4-1:0] node5090;
	wire [4-1:0] node5093;
	wire [4-1:0] node5095;
	wire [4-1:0] node5096;
	wire [4-1:0] node5099;
	wire [4-1:0] node5102;
	wire [4-1:0] node5103;
	wire [4-1:0] node5104;
	wire [4-1:0] node5105;
	wire [4-1:0] node5109;
	wire [4-1:0] node5111;
	wire [4-1:0] node5114;
	wire [4-1:0] node5115;
	wire [4-1:0] node5116;
	wire [4-1:0] node5120;
	wire [4-1:0] node5122;
	wire [4-1:0] node5125;
	wire [4-1:0] node5126;
	wire [4-1:0] node5127;
	wire [4-1:0] node5128;
	wire [4-1:0] node5130;
	wire [4-1:0] node5133;
	wire [4-1:0] node5136;
	wire [4-1:0] node5137;
	wire [4-1:0] node5138;
	wire [4-1:0] node5140;
	wire [4-1:0] node5144;
	wire [4-1:0] node5145;
	wire [4-1:0] node5148;
	wire [4-1:0] node5149;
	wire [4-1:0] node5152;
	wire [4-1:0] node5155;
	wire [4-1:0] node5156;
	wire [4-1:0] node5158;
	wire [4-1:0] node5159;
	wire [4-1:0] node5160;
	wire [4-1:0] node5165;
	wire [4-1:0] node5166;
	wire [4-1:0] node5167;
	wire [4-1:0] node5168;
	wire [4-1:0] node5172;
	wire [4-1:0] node5173;
	wire [4-1:0] node5177;
	wire [4-1:0] node5179;
	wire [4-1:0] node5180;
	wire [4-1:0] node5184;
	wire [4-1:0] node5185;
	wire [4-1:0] node5186;
	wire [4-1:0] node5187;
	wire [4-1:0] node5188;
	wire [4-1:0] node5189;
	wire [4-1:0] node5191;
	wire [4-1:0] node5193;
	wire [4-1:0] node5196;
	wire [4-1:0] node5197;
	wire [4-1:0] node5201;
	wire [4-1:0] node5202;
	wire [4-1:0] node5203;
	wire [4-1:0] node5204;
	wire [4-1:0] node5209;
	wire [4-1:0] node5212;
	wire [4-1:0] node5213;
	wire [4-1:0] node5216;
	wire [4-1:0] node5217;
	wire [4-1:0] node5219;
	wire [4-1:0] node5221;
	wire [4-1:0] node5224;
	wire [4-1:0] node5225;
	wire [4-1:0] node5227;
	wire [4-1:0] node5231;
	wire [4-1:0] node5232;
	wire [4-1:0] node5233;
	wire [4-1:0] node5234;
	wire [4-1:0] node5235;
	wire [4-1:0] node5236;
	wire [4-1:0] node5241;
	wire [4-1:0] node5243;
	wire [4-1:0] node5246;
	wire [4-1:0] node5247;
	wire [4-1:0] node5248;
	wire [4-1:0] node5249;
	wire [4-1:0] node5253;
	wire [4-1:0] node5255;
	wire [4-1:0] node5258;
	wire [4-1:0] node5259;
	wire [4-1:0] node5263;
	wire [4-1:0] node5264;
	wire [4-1:0] node5267;
	wire [4-1:0] node5268;
	wire [4-1:0] node5269;
	wire [4-1:0] node5270;
	wire [4-1:0] node5275;
	wire [4-1:0] node5277;
	wire [4-1:0] node5278;
	wire [4-1:0] node5282;
	wire [4-1:0] node5283;
	wire [4-1:0] node5284;
	wire [4-1:0] node5285;
	wire [4-1:0] node5286;
	wire [4-1:0] node5289;
	wire [4-1:0] node5291;
	wire [4-1:0] node5293;
	wire [4-1:0] node5296;
	wire [4-1:0] node5297;
	wire [4-1:0] node5298;
	wire [4-1:0] node5301;
	wire [4-1:0] node5304;
	wire [4-1:0] node5305;
	wire [4-1:0] node5308;
	wire [4-1:0] node5309;
	wire [4-1:0] node5313;
	wire [4-1:0] node5314;
	wire [4-1:0] node5315;
	wire [4-1:0] node5318;
	wire [4-1:0] node5319;
	wire [4-1:0] node5322;
	wire [4-1:0] node5324;
	wire [4-1:0] node5327;
	wire [4-1:0] node5328;
	wire [4-1:0] node5330;
	wire [4-1:0] node5333;
	wire [4-1:0] node5336;
	wire [4-1:0] node5337;
	wire [4-1:0] node5338;
	wire [4-1:0] node5339;
	wire [4-1:0] node5341;
	wire [4-1:0] node5344;
	wire [4-1:0] node5346;
	wire [4-1:0] node5349;
	wire [4-1:0] node5350;
	wire [4-1:0] node5351;
	wire [4-1:0] node5354;
	wire [4-1:0] node5358;
	wire [4-1:0] node5359;
	wire [4-1:0] node5360;
	wire [4-1:0] node5361;
	wire [4-1:0] node5365;
	wire [4-1:0] node5366;
	wire [4-1:0] node5370;
	wire [4-1:0] node5371;
	wire [4-1:0] node5372;
	wire [4-1:0] node5377;
	wire [4-1:0] node5378;
	wire [4-1:0] node5379;
	wire [4-1:0] node5380;
	wire [4-1:0] node5381;
	wire [4-1:0] node5382;
	wire [4-1:0] node5383;
	wire [4-1:0] node5387;
	wire [4-1:0] node5388;
	wire [4-1:0] node5389;
	wire [4-1:0] node5394;
	wire [4-1:0] node5395;
	wire [4-1:0] node5396;
	wire [4-1:0] node5398;
	wire [4-1:0] node5401;
	wire [4-1:0] node5404;
	wire [4-1:0] node5405;
	wire [4-1:0] node5406;
	wire [4-1:0] node5408;
	wire [4-1:0] node5411;
	wire [4-1:0] node5414;
	wire [4-1:0] node5416;
	wire [4-1:0] node5419;
	wire [4-1:0] node5420;
	wire [4-1:0] node5421;
	wire [4-1:0] node5422;
	wire [4-1:0] node5424;
	wire [4-1:0] node5425;
	wire [4-1:0] node5429;
	wire [4-1:0] node5430;
	wire [4-1:0] node5431;
	wire [4-1:0] node5435;
	wire [4-1:0] node5438;
	wire [4-1:0] node5439;
	wire [4-1:0] node5441;
	wire [4-1:0] node5444;
	wire [4-1:0] node5447;
	wire [4-1:0] node5449;
	wire [4-1:0] node5450;
	wire [4-1:0] node5451;
	wire [4-1:0] node5455;
	wire [4-1:0] node5458;
	wire [4-1:0] node5459;
	wire [4-1:0] node5460;
	wire [4-1:0] node5461;
	wire [4-1:0] node5462;
	wire [4-1:0] node5463;
	wire [4-1:0] node5468;
	wire [4-1:0] node5470;
	wire [4-1:0] node5472;
	wire [4-1:0] node5473;
	wire [4-1:0] node5477;
	wire [4-1:0] node5478;
	wire [4-1:0] node5479;
	wire [4-1:0] node5480;
	wire [4-1:0] node5484;
	wire [4-1:0] node5486;
	wire [4-1:0] node5489;
	wire [4-1:0] node5491;
	wire [4-1:0] node5492;
	wire [4-1:0] node5493;
	wire [4-1:0] node5496;
	wire [4-1:0] node5500;
	wire [4-1:0] node5501;
	wire [4-1:0] node5502;
	wire [4-1:0] node5503;
	wire [4-1:0] node5504;
	wire [4-1:0] node5508;
	wire [4-1:0] node5509;
	wire [4-1:0] node5512;
	wire [4-1:0] node5515;
	wire [4-1:0] node5516;
	wire [4-1:0] node5520;
	wire [4-1:0] node5521;
	wire [4-1:0] node5523;
	wire [4-1:0] node5524;
	wire [4-1:0] node5525;
	wire [4-1:0] node5530;
	wire [4-1:0] node5531;
	wire [4-1:0] node5534;
	wire [4-1:0] node5535;
	wire [4-1:0] node5539;
	wire [4-1:0] node5540;
	wire [4-1:0] node5541;
	wire [4-1:0] node5542;
	wire [4-1:0] node5543;
	wire [4-1:0] node5544;
	wire [4-1:0] node5545;
	wire [4-1:0] node5548;
	wire [4-1:0] node5551;
	wire [4-1:0] node5554;
	wire [4-1:0] node5555;
	wire [4-1:0] node5557;
	wire [4-1:0] node5558;
	wire [4-1:0] node5563;
	wire [4-1:0] node5564;
	wire [4-1:0] node5565;
	wire [4-1:0] node5567;
	wire [4-1:0] node5571;
	wire [4-1:0] node5572;
	wire [4-1:0] node5575;
	wire [4-1:0] node5576;
	wire [4-1:0] node5577;
	wire [4-1:0] node5581;
	wire [4-1:0] node5584;
	wire [4-1:0] node5585;
	wire [4-1:0] node5586;
	wire [4-1:0] node5587;
	wire [4-1:0] node5589;
	wire [4-1:0] node5592;
	wire [4-1:0] node5594;
	wire [4-1:0] node5597;
	wire [4-1:0] node5598;
	wire [4-1:0] node5600;
	wire [4-1:0] node5604;
	wire [4-1:0] node5605;
	wire [4-1:0] node5607;
	wire [4-1:0] node5608;
	wire [4-1:0] node5612;
	wire [4-1:0] node5613;
	wire [4-1:0] node5616;
	wire [4-1:0] node5618;
	wire [4-1:0] node5621;
	wire [4-1:0] node5622;
	wire [4-1:0] node5623;
	wire [4-1:0] node5624;
	wire [4-1:0] node5626;
	wire [4-1:0] node5627;
	wire [4-1:0] node5628;
	wire [4-1:0] node5633;
	wire [4-1:0] node5635;
	wire [4-1:0] node5638;
	wire [4-1:0] node5639;
	wire [4-1:0] node5640;
	wire [4-1:0] node5642;
	wire [4-1:0] node5644;
	wire [4-1:0] node5647;
	wire [4-1:0] node5648;
	wire [4-1:0] node5649;
	wire [4-1:0] node5652;
	wire [4-1:0] node5656;
	wire [4-1:0] node5657;
	wire [4-1:0] node5658;
	wire [4-1:0] node5662;
	wire [4-1:0] node5663;
	wire [4-1:0] node5665;
	wire [4-1:0] node5668;
	wire [4-1:0] node5671;
	wire [4-1:0] node5672;
	wire [4-1:0] node5673;
	wire [4-1:0] node5674;
	wire [4-1:0] node5676;
	wire [4-1:0] node5680;
	wire [4-1:0] node5681;
	wire [4-1:0] node5684;
	wire [4-1:0] node5687;
	wire [4-1:0] node5688;
	wire [4-1:0] node5689;
	wire [4-1:0] node5690;
	wire [4-1:0] node5693;
	wire [4-1:0] node5694;
	wire [4-1:0] node5698;
	wire [4-1:0] node5699;
	wire [4-1:0] node5703;
	wire [4-1:0] node5705;
	wire [4-1:0] node5708;
	wire [4-1:0] node5709;
	wire [4-1:0] node5710;
	wire [4-1:0] node5711;
	wire [4-1:0] node5712;
	wire [4-1:0] node5713;
	wire [4-1:0] node5714;
	wire [4-1:0] node5715;
	wire [4-1:0] node5716;
	wire [4-1:0] node5717;
	wire [4-1:0] node5719;
	wire [4-1:0] node5722;
	wire [4-1:0] node5724;
	wire [4-1:0] node5727;
	wire [4-1:0] node5728;
	wire [4-1:0] node5730;
	wire [4-1:0] node5732;
	wire [4-1:0] node5735;
	wire [4-1:0] node5736;
	wire [4-1:0] node5740;
	wire [4-1:0] node5741;
	wire [4-1:0] node5742;
	wire [4-1:0] node5744;
	wire [4-1:0] node5746;
	wire [4-1:0] node5749;
	wire [4-1:0] node5750;
	wire [4-1:0] node5752;
	wire [4-1:0] node5756;
	wire [4-1:0] node5757;
	wire [4-1:0] node5758;
	wire [4-1:0] node5759;
	wire [4-1:0] node5763;
	wire [4-1:0] node5764;
	wire [4-1:0] node5768;
	wire [4-1:0] node5769;
	wire [4-1:0] node5772;
	wire [4-1:0] node5775;
	wire [4-1:0] node5776;
	wire [4-1:0] node5777;
	wire [4-1:0] node5778;
	wire [4-1:0] node5779;
	wire [4-1:0] node5780;
	wire [4-1:0] node5783;
	wire [4-1:0] node5785;
	wire [4-1:0] node5788;
	wire [4-1:0] node5791;
	wire [4-1:0] node5792;
	wire [4-1:0] node5795;
	wire [4-1:0] node5797;
	wire [4-1:0] node5798;
	wire [4-1:0] node5802;
	wire [4-1:0] node5803;
	wire [4-1:0] node5804;
	wire [4-1:0] node5805;
	wire [4-1:0] node5809;
	wire [4-1:0] node5810;
	wire [4-1:0] node5812;
	wire [4-1:0] node5815;
	wire [4-1:0] node5818;
	wire [4-1:0] node5820;
	wire [4-1:0] node5822;
	wire [4-1:0] node5825;
	wire [4-1:0] node5826;
	wire [4-1:0] node5827;
	wire [4-1:0] node5828;
	wire [4-1:0] node5829;
	wire [4-1:0] node5831;
	wire [4-1:0] node5836;
	wire [4-1:0] node5837;
	wire [4-1:0] node5840;
	wire [4-1:0] node5842;
	wire [4-1:0] node5845;
	wire [4-1:0] node5846;
	wire [4-1:0] node5848;
	wire [4-1:0] node5849;
	wire [4-1:0] node5853;
	wire [4-1:0] node5854;
	wire [4-1:0] node5857;
	wire [4-1:0] node5858;
	wire [4-1:0] node5862;
	wire [4-1:0] node5863;
	wire [4-1:0] node5864;
	wire [4-1:0] node5865;
	wire [4-1:0] node5866;
	wire [4-1:0] node5868;
	wire [4-1:0] node5870;
	wire [4-1:0] node5873;
	wire [4-1:0] node5875;
	wire [4-1:0] node5878;
	wire [4-1:0] node5879;
	wire [4-1:0] node5880;
	wire [4-1:0] node5882;
	wire [4-1:0] node5885;
	wire [4-1:0] node5887;
	wire [4-1:0] node5890;
	wire [4-1:0] node5892;
	wire [4-1:0] node5895;
	wire [4-1:0] node5896;
	wire [4-1:0] node5897;
	wire [4-1:0] node5900;
	wire [4-1:0] node5901;
	wire [4-1:0] node5904;
	wire [4-1:0] node5905;
	wire [4-1:0] node5907;
	wire [4-1:0] node5911;
	wire [4-1:0] node5912;
	wire [4-1:0] node5914;
	wire [4-1:0] node5915;
	wire [4-1:0] node5916;
	wire [4-1:0] node5920;
	wire [4-1:0] node5923;
	wire [4-1:0] node5924;
	wire [4-1:0] node5927;
	wire [4-1:0] node5930;
	wire [4-1:0] node5931;
	wire [4-1:0] node5932;
	wire [4-1:0] node5933;
	wire [4-1:0] node5934;
	wire [4-1:0] node5938;
	wire [4-1:0] node5939;
	wire [4-1:0] node5942;
	wire [4-1:0] node5943;
	wire [4-1:0] node5944;
	wire [4-1:0] node5948;
	wire [4-1:0] node5951;
	wire [4-1:0] node5952;
	wire [4-1:0] node5953;
	wire [4-1:0] node5957;
	wire [4-1:0] node5958;
	wire [4-1:0] node5960;
	wire [4-1:0] node5964;
	wire [4-1:0] node5965;
	wire [4-1:0] node5966;
	wire [4-1:0] node5968;
	wire [4-1:0] node5970;
	wire [4-1:0] node5972;
	wire [4-1:0] node5975;
	wire [4-1:0] node5976;
	wire [4-1:0] node5977;
	wire [4-1:0] node5980;
	wire [4-1:0] node5981;
	wire [4-1:0] node5985;
	wire [4-1:0] node5987;
	wire [4-1:0] node5990;
	wire [4-1:0] node5991;
	wire [4-1:0] node5992;
	wire [4-1:0] node5993;
	wire [4-1:0] node5995;
	wire [4-1:0] node5998;
	wire [4-1:0] node6001;
	wire [4-1:0] node6003;
	wire [4-1:0] node6006;
	wire [4-1:0] node6007;
	wire [4-1:0] node6008;
	wire [4-1:0] node6011;
	wire [4-1:0] node6014;
	wire [4-1:0] node6015;
	wire [4-1:0] node6016;
	wire [4-1:0] node6021;
	wire [4-1:0] node6022;
	wire [4-1:0] node6023;
	wire [4-1:0] node6024;
	wire [4-1:0] node6025;
	wire [4-1:0] node6026;
	wire [4-1:0] node6027;
	wire [4-1:0] node6031;
	wire [4-1:0] node6032;
	wire [4-1:0] node6034;
	wire [4-1:0] node6037;
	wire [4-1:0] node6038;
	wire [4-1:0] node6042;
	wire [4-1:0] node6044;
	wire [4-1:0] node6046;
	wire [4-1:0] node6048;
	wire [4-1:0] node6051;
	wire [4-1:0] node6052;
	wire [4-1:0] node6053;
	wire [4-1:0] node6054;
	wire [4-1:0] node6055;
	wire [4-1:0] node6056;
	wire [4-1:0] node6061;
	wire [4-1:0] node6062;
	wire [4-1:0] node6063;
	wire [4-1:0] node6067;
	wire [4-1:0] node6070;
	wire [4-1:0] node6072;
	wire [4-1:0] node6073;
	wire [4-1:0] node6074;
	wire [4-1:0] node6078;
	wire [4-1:0] node6081;
	wire [4-1:0] node6082;
	wire [4-1:0] node6083;
	wire [4-1:0] node6087;
	wire [4-1:0] node6088;
	wire [4-1:0] node6089;
	wire [4-1:0] node6091;
	wire [4-1:0] node6095;
	wire [4-1:0] node6096;
	wire [4-1:0] node6097;
	wire [4-1:0] node6102;
	wire [4-1:0] node6103;
	wire [4-1:0] node6104;
	wire [4-1:0] node6105;
	wire [4-1:0] node6107;
	wire [4-1:0] node6110;
	wire [4-1:0] node6111;
	wire [4-1:0] node6112;
	wire [4-1:0] node6114;
	wire [4-1:0] node6119;
	wire [4-1:0] node6120;
	wire [4-1:0] node6122;
	wire [4-1:0] node6125;
	wire [4-1:0] node6126;
	wire [4-1:0] node6129;
	wire [4-1:0] node6130;
	wire [4-1:0] node6132;
	wire [4-1:0] node6136;
	wire [4-1:0] node6137;
	wire [4-1:0] node6138;
	wire [4-1:0] node6139;
	wire [4-1:0] node6141;
	wire [4-1:0] node6145;
	wire [4-1:0] node6146;
	wire [4-1:0] node6149;
	wire [4-1:0] node6152;
	wire [4-1:0] node6153;
	wire [4-1:0] node6154;
	wire [4-1:0] node6156;
	wire [4-1:0] node6160;
	wire [4-1:0] node6162;
	wire [4-1:0] node6163;
	wire [4-1:0] node6164;
	wire [4-1:0] node6167;
	wire [4-1:0] node6171;
	wire [4-1:0] node6172;
	wire [4-1:0] node6173;
	wire [4-1:0] node6174;
	wire [4-1:0] node6175;
	wire [4-1:0] node6176;
	wire [4-1:0] node6177;
	wire [4-1:0] node6178;
	wire [4-1:0] node6182;
	wire [4-1:0] node6184;
	wire [4-1:0] node6188;
	wire [4-1:0] node6189;
	wire [4-1:0] node6190;
	wire [4-1:0] node6191;
	wire [4-1:0] node6196;
	wire [4-1:0] node6199;
	wire [4-1:0] node6200;
	wire [4-1:0] node6201;
	wire [4-1:0] node6203;
	wire [4-1:0] node6206;
	wire [4-1:0] node6208;
	wire [4-1:0] node6209;
	wire [4-1:0] node6213;
	wire [4-1:0] node6215;
	wire [4-1:0] node6216;
	wire [4-1:0] node6219;
	wire [4-1:0] node6221;
	wire [4-1:0] node6224;
	wire [4-1:0] node6225;
	wire [4-1:0] node6226;
	wire [4-1:0] node6228;
	wire [4-1:0] node6231;
	wire [4-1:0] node6232;
	wire [4-1:0] node6234;
	wire [4-1:0] node6237;
	wire [4-1:0] node6239;
	wire [4-1:0] node6241;
	wire [4-1:0] node6244;
	wire [4-1:0] node6245;
	wire [4-1:0] node6246;
	wire [4-1:0] node6248;
	wire [4-1:0] node6252;
	wire [4-1:0] node6253;
	wire [4-1:0] node6257;
	wire [4-1:0] node6258;
	wire [4-1:0] node6259;
	wire [4-1:0] node6260;
	wire [4-1:0] node6261;
	wire [4-1:0] node6263;
	wire [4-1:0] node6264;
	wire [4-1:0] node6269;
	wire [4-1:0] node6270;
	wire [4-1:0] node6271;
	wire [4-1:0] node6276;
	wire [4-1:0] node6277;
	wire [4-1:0] node6278;
	wire [4-1:0] node6279;
	wire [4-1:0] node6280;
	wire [4-1:0] node6285;
	wire [4-1:0] node6286;
	wire [4-1:0] node6290;
	wire [4-1:0] node6292;
	wire [4-1:0] node6293;
	wire [4-1:0] node6296;
	wire [4-1:0] node6299;
	wire [4-1:0] node6300;
	wire [4-1:0] node6302;
	wire [4-1:0] node6303;
	wire [4-1:0] node6304;
	wire [4-1:0] node6308;
	wire [4-1:0] node6311;
	wire [4-1:0] node6312;
	wire [4-1:0] node6313;
	wire [4-1:0] node6314;
	wire [4-1:0] node6316;
	wire [4-1:0] node6320;
	wire [4-1:0] node6322;
	wire [4-1:0] node6323;
	wire [4-1:0] node6327;
	wire [4-1:0] node6328;
	wire [4-1:0] node6331;
	wire [4-1:0] node6332;
	wire [4-1:0] node6335;
	wire [4-1:0] node6338;
	wire [4-1:0] node6339;
	wire [4-1:0] node6340;
	wire [4-1:0] node6341;
	wire [4-1:0] node6342;
	wire [4-1:0] node6343;
	wire [4-1:0] node6344;
	wire [4-1:0] node6345;
	wire [4-1:0] node6349;
	wire [4-1:0] node6350;
	wire [4-1:0] node6351;
	wire [4-1:0] node6353;
	wire [4-1:0] node6357;
	wire [4-1:0] node6359;
	wire [4-1:0] node6362;
	wire [4-1:0] node6363;
	wire [4-1:0] node6364;
	wire [4-1:0] node6366;
	wire [4-1:0] node6367;
	wire [4-1:0] node6371;
	wire [4-1:0] node6372;
	wire [4-1:0] node6375;
	wire [4-1:0] node6378;
	wire [4-1:0] node6379;
	wire [4-1:0] node6380;
	wire [4-1:0] node6382;
	wire [4-1:0] node6385;
	wire [4-1:0] node6386;
	wire [4-1:0] node6389;
	wire [4-1:0] node6393;
	wire [4-1:0] node6394;
	wire [4-1:0] node6395;
	wire [4-1:0] node6396;
	wire [4-1:0] node6399;
	wire [4-1:0] node6402;
	wire [4-1:0] node6403;
	wire [4-1:0] node6404;
	wire [4-1:0] node6408;
	wire [4-1:0] node6410;
	wire [4-1:0] node6412;
	wire [4-1:0] node6415;
	wire [4-1:0] node6416;
	wire [4-1:0] node6417;
	wire [4-1:0] node6420;
	wire [4-1:0] node6421;
	wire [4-1:0] node6424;
	wire [4-1:0] node6426;
	wire [4-1:0] node6429;
	wire [4-1:0] node6430;
	wire [4-1:0] node6432;
	wire [4-1:0] node6434;
	wire [4-1:0] node6438;
	wire [4-1:0] node6439;
	wire [4-1:0] node6440;
	wire [4-1:0] node6441;
	wire [4-1:0] node6442;
	wire [4-1:0] node6444;
	wire [4-1:0] node6445;
	wire [4-1:0] node6449;
	wire [4-1:0] node6450;
	wire [4-1:0] node6451;
	wire [4-1:0] node6455;
	wire [4-1:0] node6458;
	wire [4-1:0] node6460;
	wire [4-1:0] node6461;
	wire [4-1:0] node6465;
	wire [4-1:0] node6466;
	wire [4-1:0] node6467;
	wire [4-1:0] node6469;
	wire [4-1:0] node6472;
	wire [4-1:0] node6474;
	wire [4-1:0] node6477;
	wire [4-1:0] node6478;
	wire [4-1:0] node6480;
	wire [4-1:0] node6483;
	wire [4-1:0] node6485;
	wire [4-1:0] node6488;
	wire [4-1:0] node6489;
	wire [4-1:0] node6490;
	wire [4-1:0] node6491;
	wire [4-1:0] node6493;
	wire [4-1:0] node6496;
	wire [4-1:0] node6498;
	wire [4-1:0] node6500;
	wire [4-1:0] node6503;
	wire [4-1:0] node6504;
	wire [4-1:0] node6505;
	wire [4-1:0] node6507;
	wire [4-1:0] node6510;
	wire [4-1:0] node6512;
	wire [4-1:0] node6515;
	wire [4-1:0] node6518;
	wire [4-1:0] node6519;
	wire [4-1:0] node6520;
	wire [4-1:0] node6523;
	wire [4-1:0] node6524;
	wire [4-1:0] node6525;
	wire [4-1:0] node6530;
	wire [4-1:0] node6531;
	wire [4-1:0] node6533;
	wire [4-1:0] node6534;
	wire [4-1:0] node6538;
	wire [4-1:0] node6539;
	wire [4-1:0] node6543;
	wire [4-1:0] node6544;
	wire [4-1:0] node6545;
	wire [4-1:0] node6546;
	wire [4-1:0] node6547;
	wire [4-1:0] node6549;
	wire [4-1:0] node6552;
	wire [4-1:0] node6553;
	wire [4-1:0] node6557;
	wire [4-1:0] node6558;
	wire [4-1:0] node6559;
	wire [4-1:0] node6560;
	wire [4-1:0] node6564;
	wire [4-1:0] node6566;
	wire [4-1:0] node6569;
	wire [4-1:0] node6570;
	wire [4-1:0] node6571;
	wire [4-1:0] node6575;
	wire [4-1:0] node6576;
	wire [4-1:0] node6577;
	wire [4-1:0] node6581;
	wire [4-1:0] node6584;
	wire [4-1:0] node6585;
	wire [4-1:0] node6586;
	wire [4-1:0] node6587;
	wire [4-1:0] node6588;
	wire [4-1:0] node6592;
	wire [4-1:0] node6594;
	wire [4-1:0] node6597;
	wire [4-1:0] node6598;
	wire [4-1:0] node6601;
	wire [4-1:0] node6603;
	wire [4-1:0] node6606;
	wire [4-1:0] node6607;
	wire [4-1:0] node6609;
	wire [4-1:0] node6610;
	wire [4-1:0] node6611;
	wire [4-1:0] node6615;
	wire [4-1:0] node6618;
	wire [4-1:0] node6620;
	wire [4-1:0] node6623;
	wire [4-1:0] node6624;
	wire [4-1:0] node6625;
	wire [4-1:0] node6626;
	wire [4-1:0] node6627;
	wire [4-1:0] node6630;
	wire [4-1:0] node6633;
	wire [4-1:0] node6635;
	wire [4-1:0] node6638;
	wire [4-1:0] node6639;
	wire [4-1:0] node6640;
	wire [4-1:0] node6641;
	wire [4-1:0] node6645;
	wire [4-1:0] node6646;
	wire [4-1:0] node6650;
	wire [4-1:0] node6651;
	wire [4-1:0] node6655;
	wire [4-1:0] node6656;
	wire [4-1:0] node6657;
	wire [4-1:0] node6658;
	wire [4-1:0] node6659;
	wire [4-1:0] node6663;
	wire [4-1:0] node6664;
	wire [4-1:0] node6665;
	wire [4-1:0] node6669;
	wire [4-1:0] node6671;
	wire [4-1:0] node6674;
	wire [4-1:0] node6677;
	wire [4-1:0] node6678;
	wire [4-1:0] node6679;
	wire [4-1:0] node6680;
	wire [4-1:0] node6681;
	wire [4-1:0] node6686;
	wire [4-1:0] node6689;
	wire [4-1:0] node6690;
	wire [4-1:0] node6691;
	wire [4-1:0] node6692;
	wire [4-1:0] node6695;
	wire [4-1:0] node6698;
	wire [4-1:0] node6702;
	wire [4-1:0] node6703;
	wire [4-1:0] node6704;
	wire [4-1:0] node6705;
	wire [4-1:0] node6706;
	wire [4-1:0] node6707;
	wire [4-1:0] node6708;
	wire [4-1:0] node6710;
	wire [4-1:0] node6714;
	wire [4-1:0] node6715;
	wire [4-1:0] node6717;
	wire [4-1:0] node6719;
	wire [4-1:0] node6723;
	wire [4-1:0] node6724;
	wire [4-1:0] node6725;
	wire [4-1:0] node6728;
	wire [4-1:0] node6729;
	wire [4-1:0] node6732;
	wire [4-1:0] node6735;
	wire [4-1:0] node6736;
	wire [4-1:0] node6739;
	wire [4-1:0] node6742;
	wire [4-1:0] node6743;
	wire [4-1:0] node6744;
	wire [4-1:0] node6746;
	wire [4-1:0] node6748;
	wire [4-1:0] node6751;
	wire [4-1:0] node6752;
	wire [4-1:0] node6754;
	wire [4-1:0] node6757;
	wire [4-1:0] node6758;
	wire [4-1:0] node6759;
	wire [4-1:0] node6762;
	wire [4-1:0] node6765;
	wire [4-1:0] node6766;
	wire [4-1:0] node6769;
	wire [4-1:0] node6772;
	wire [4-1:0] node6773;
	wire [4-1:0] node6775;
	wire [4-1:0] node6778;
	wire [4-1:0] node6780;
	wire [4-1:0] node6781;
	wire [4-1:0] node6782;
	wire [4-1:0] node6786;
	wire [4-1:0] node6789;
	wire [4-1:0] node6790;
	wire [4-1:0] node6791;
	wire [4-1:0] node6792;
	wire [4-1:0] node6793;
	wire [4-1:0] node6796;
	wire [4-1:0] node6798;
	wire [4-1:0] node6799;
	wire [4-1:0] node6803;
	wire [4-1:0] node6804;
	wire [4-1:0] node6806;
	wire [4-1:0] node6810;
	wire [4-1:0] node6811;
	wire [4-1:0] node6812;
	wire [4-1:0] node6814;
	wire [4-1:0] node6815;
	wire [4-1:0] node6819;
	wire [4-1:0] node6820;
	wire [4-1:0] node6824;
	wire [4-1:0] node6825;
	wire [4-1:0] node6828;
	wire [4-1:0] node6830;
	wire [4-1:0] node6831;
	wire [4-1:0] node6835;
	wire [4-1:0] node6836;
	wire [4-1:0] node6837;
	wire [4-1:0] node6838;
	wire [4-1:0] node6840;
	wire [4-1:0] node6842;
	wire [4-1:0] node6845;
	wire [4-1:0] node6846;
	wire [4-1:0] node6850;
	wire [4-1:0] node6851;
	wire [4-1:0] node6852;
	wire [4-1:0] node6855;
	wire [4-1:0] node6857;
	wire [4-1:0] node6860;
	wire [4-1:0] node6863;
	wire [4-1:0] node6864;
	wire [4-1:0] node6866;
	wire [4-1:0] node6869;
	wire [4-1:0] node6870;
	wire [4-1:0] node6872;
	wire [4-1:0] node6873;
	wire [4-1:0] node6876;
	wire [4-1:0] node6880;
	wire [4-1:0] node6881;
	wire [4-1:0] node6882;
	wire [4-1:0] node6883;
	wire [4-1:0] node6884;
	wire [4-1:0] node6886;
	wire [4-1:0] node6887;
	wire [4-1:0] node6891;
	wire [4-1:0] node6892;
	wire [4-1:0] node6893;
	wire [4-1:0] node6894;
	wire [4-1:0] node6899;
	wire [4-1:0] node6902;
	wire [4-1:0] node6903;
	wire [4-1:0] node6904;
	wire [4-1:0] node6905;
	wire [4-1:0] node6909;
	wire [4-1:0] node6912;
	wire [4-1:0] node6913;
	wire [4-1:0] node6916;
	wire [4-1:0] node6919;
	wire [4-1:0] node6920;
	wire [4-1:0] node6921;
	wire [4-1:0] node6922;
	wire [4-1:0] node6925;
	wire [4-1:0] node6926;
	wire [4-1:0] node6927;
	wire [4-1:0] node6932;
	wire [4-1:0] node6933;
	wire [4-1:0] node6934;
	wire [4-1:0] node6938;
	wire [4-1:0] node6941;
	wire [4-1:0] node6942;
	wire [4-1:0] node6943;
	wire [4-1:0] node6945;
	wire [4-1:0] node6948;
	wire [4-1:0] node6951;
	wire [4-1:0] node6953;
	wire [4-1:0] node6956;
	wire [4-1:0] node6957;
	wire [4-1:0] node6958;
	wire [4-1:0] node6959;
	wire [4-1:0] node6960;
	wire [4-1:0] node6961;
	wire [4-1:0] node6964;
	wire [4-1:0] node6966;
	wire [4-1:0] node6969;
	wire [4-1:0] node6972;
	wire [4-1:0] node6974;
	wire [4-1:0] node6975;
	wire [4-1:0] node6976;
	wire [4-1:0] node6980;
	wire [4-1:0] node6981;
	wire [4-1:0] node6984;
	wire [4-1:0] node6987;
	wire [4-1:0] node6988;
	wire [4-1:0] node6990;
	wire [4-1:0] node6992;
	wire [4-1:0] node6993;
	wire [4-1:0] node6997;
	wire [4-1:0] node7000;
	wire [4-1:0] node7001;
	wire [4-1:0] node7002;
	wire [4-1:0] node7003;
	wire [4-1:0] node7005;
	wire [4-1:0] node7008;
	wire [4-1:0] node7011;
	wire [4-1:0] node7012;
	wire [4-1:0] node7013;
	wire [4-1:0] node7015;
	wire [4-1:0] node7020;
	wire [4-1:0] node7021;
	wire [4-1:0] node7022;
	wire [4-1:0] node7024;
	wire [4-1:0] node7028;
	wire [4-1:0] node7029;
	wire [4-1:0] node7031;
	wire [4-1:0] node7035;
	wire [4-1:0] node7036;
	wire [4-1:0] node7037;
	wire [4-1:0] node7038;
	wire [4-1:0] node7039;
	wire [4-1:0] node7040;
	wire [4-1:0] node7041;
	wire [4-1:0] node7042;
	wire [4-1:0] node7043;
	wire [4-1:0] node7044;
	wire [4-1:0] node7048;
	wire [4-1:0] node7049;
	wire [4-1:0] node7051;
	wire [4-1:0] node7054;
	wire [4-1:0] node7056;
	wire [4-1:0] node7059;
	wire [4-1:0] node7060;
	wire [4-1:0] node7061;
	wire [4-1:0] node7066;
	wire [4-1:0] node7067;
	wire [4-1:0] node7068;
	wire [4-1:0] node7070;
	wire [4-1:0] node7071;
	wire [4-1:0] node7075;
	wire [4-1:0] node7076;
	wire [4-1:0] node7078;
	wire [4-1:0] node7081;
	wire [4-1:0] node7083;
	wire [4-1:0] node7086;
	wire [4-1:0] node7089;
	wire [4-1:0] node7090;
	wire [4-1:0] node7091;
	wire [4-1:0] node7093;
	wire [4-1:0] node7095;
	wire [4-1:0] node7098;
	wire [4-1:0] node7099;
	wire [4-1:0] node7101;
	wire [4-1:0] node7102;
	wire [4-1:0] node7106;
	wire [4-1:0] node7107;
	wire [4-1:0] node7111;
	wire [4-1:0] node7112;
	wire [4-1:0] node7115;
	wire [4-1:0] node7116;
	wire [4-1:0] node7119;
	wire [4-1:0] node7121;
	wire [4-1:0] node7123;
	wire [4-1:0] node7126;
	wire [4-1:0] node7127;
	wire [4-1:0] node7128;
	wire [4-1:0] node7129;
	wire [4-1:0] node7130;
	wire [4-1:0] node7134;
	wire [4-1:0] node7136;
	wire [4-1:0] node7139;
	wire [4-1:0] node7140;
	wire [4-1:0] node7143;
	wire [4-1:0] node7144;
	wire [4-1:0] node7146;
	wire [4-1:0] node7147;
	wire [4-1:0] node7151;
	wire [4-1:0] node7153;
	wire [4-1:0] node7156;
	wire [4-1:0] node7157;
	wire [4-1:0] node7158;
	wire [4-1:0] node7159;
	wire [4-1:0] node7161;
	wire [4-1:0] node7164;
	wire [4-1:0] node7166;
	wire [4-1:0] node7169;
	wire [4-1:0] node7170;
	wire [4-1:0] node7171;
	wire [4-1:0] node7173;
	wire [4-1:0] node7176;
	wire [4-1:0] node7180;
	wire [4-1:0] node7181;
	wire [4-1:0] node7182;
	wire [4-1:0] node7184;
	wire [4-1:0] node7186;
	wire [4-1:0] node7189;
	wire [4-1:0] node7190;
	wire [4-1:0] node7194;
	wire [4-1:0] node7195;
	wire [4-1:0] node7197;
	wire [4-1:0] node7198;
	wire [4-1:0] node7203;
	wire [4-1:0] node7204;
	wire [4-1:0] node7205;
	wire [4-1:0] node7206;
	wire [4-1:0] node7207;
	wire [4-1:0] node7210;
	wire [4-1:0] node7212;
	wire [4-1:0] node7214;
	wire [4-1:0] node7216;
	wire [4-1:0] node7219;
	wire [4-1:0] node7220;
	wire [4-1:0] node7221;
	wire [4-1:0] node7223;
	wire [4-1:0] node7226;
	wire [4-1:0] node7227;
	wire [4-1:0] node7228;
	wire [4-1:0] node7233;
	wire [4-1:0] node7234;
	wire [4-1:0] node7235;
	wire [4-1:0] node7236;
	wire [4-1:0] node7241;
	wire [4-1:0] node7244;
	wire [4-1:0] node7245;
	wire [4-1:0] node7246;
	wire [4-1:0] node7247;
	wire [4-1:0] node7250;
	wire [4-1:0] node7253;
	wire [4-1:0] node7254;
	wire [4-1:0] node7258;
	wire [4-1:0] node7259;
	wire [4-1:0] node7261;
	wire [4-1:0] node7262;
	wire [4-1:0] node7263;
	wire [4-1:0] node7268;
	wire [4-1:0] node7269;
	wire [4-1:0] node7270;
	wire [4-1:0] node7271;
	wire [4-1:0] node7276;
	wire [4-1:0] node7278;
	wire [4-1:0] node7281;
	wire [4-1:0] node7282;
	wire [4-1:0] node7283;
	wire [4-1:0] node7284;
	wire [4-1:0] node7285;
	wire [4-1:0] node7288;
	wire [4-1:0] node7290;
	wire [4-1:0] node7293;
	wire [4-1:0] node7294;
	wire [4-1:0] node7295;
	wire [4-1:0] node7297;
	wire [4-1:0] node7301;
	wire [4-1:0] node7302;
	wire [4-1:0] node7305;
	wire [4-1:0] node7307;
	wire [4-1:0] node7310;
	wire [4-1:0] node7311;
	wire [4-1:0] node7314;
	wire [4-1:0] node7315;
	wire [4-1:0] node7316;
	wire [4-1:0] node7319;
	wire [4-1:0] node7322;
	wire [4-1:0] node7324;
	wire [4-1:0] node7327;
	wire [4-1:0] node7328;
	wire [4-1:0] node7329;
	wire [4-1:0] node7330;
	wire [4-1:0] node7333;
	wire [4-1:0] node7335;
	wire [4-1:0] node7338;
	wire [4-1:0] node7341;
	wire [4-1:0] node7342;
	wire [4-1:0] node7344;
	wire [4-1:0] node7348;
	wire [4-1:0] node7349;
	wire [4-1:0] node7350;
	wire [4-1:0] node7351;
	wire [4-1:0] node7352;
	wire [4-1:0] node7353;
	wire [4-1:0] node7354;
	wire [4-1:0] node7355;
	wire [4-1:0] node7357;
	wire [4-1:0] node7360;
	wire [4-1:0] node7361;
	wire [4-1:0] node7364;
	wire [4-1:0] node7367;
	wire [4-1:0] node7370;
	wire [4-1:0] node7372;
	wire [4-1:0] node7375;
	wire [4-1:0] node7376;
	wire [4-1:0] node7377;
	wire [4-1:0] node7380;
	wire [4-1:0] node7383;
	wire [4-1:0] node7386;
	wire [4-1:0] node7387;
	wire [4-1:0] node7388;
	wire [4-1:0] node7389;
	wire [4-1:0] node7392;
	wire [4-1:0] node7394;
	wire [4-1:0] node7395;
	wire [4-1:0] node7399;
	wire [4-1:0] node7401;
	wire [4-1:0] node7402;
	wire [4-1:0] node7406;
	wire [4-1:0] node7407;
	wire [4-1:0] node7409;
	wire [4-1:0] node7411;
	wire [4-1:0] node7414;
	wire [4-1:0] node7416;
	wire [4-1:0] node7417;
	wire [4-1:0] node7421;
	wire [4-1:0] node7422;
	wire [4-1:0] node7423;
	wire [4-1:0] node7424;
	wire [4-1:0] node7425;
	wire [4-1:0] node7428;
	wire [4-1:0] node7431;
	wire [4-1:0] node7432;
	wire [4-1:0] node7436;
	wire [4-1:0] node7437;
	wire [4-1:0] node7438;
	wire [4-1:0] node7440;
	wire [4-1:0] node7441;
	wire [4-1:0] node7445;
	wire [4-1:0] node7447;
	wire [4-1:0] node7450;
	wire [4-1:0] node7453;
	wire [4-1:0] node7454;
	wire [4-1:0] node7455;
	wire [4-1:0] node7457;
	wire [4-1:0] node7459;
	wire [4-1:0] node7462;
	wire [4-1:0] node7464;
	wire [4-1:0] node7466;
	wire [4-1:0] node7469;
	wire [4-1:0] node7470;
	wire [4-1:0] node7471;
	wire [4-1:0] node7472;
	wire [4-1:0] node7477;
	wire [4-1:0] node7478;
	wire [4-1:0] node7481;
	wire [4-1:0] node7482;
	wire [4-1:0] node7486;
	wire [4-1:0] node7487;
	wire [4-1:0] node7488;
	wire [4-1:0] node7489;
	wire [4-1:0] node7490;
	wire [4-1:0] node7491;
	wire [4-1:0] node7495;
	wire [4-1:0] node7496;
	wire [4-1:0] node7499;
	wire [4-1:0] node7500;
	wire [4-1:0] node7504;
	wire [4-1:0] node7505;
	wire [4-1:0] node7507;
	wire [4-1:0] node7509;
	wire [4-1:0] node7510;
	wire [4-1:0] node7514;
	wire [4-1:0] node7515;
	wire [4-1:0] node7519;
	wire [4-1:0] node7520;
	wire [4-1:0] node7521;
	wire [4-1:0] node7522;
	wire [4-1:0] node7524;
	wire [4-1:0] node7527;
	wire [4-1:0] node7528;
	wire [4-1:0] node7531;
	wire [4-1:0] node7532;
	wire [4-1:0] node7535;
	wire [4-1:0] node7538;
	wire [4-1:0] node7539;
	wire [4-1:0] node7540;
	wire [4-1:0] node7543;
	wire [4-1:0] node7546;
	wire [4-1:0] node7548;
	wire [4-1:0] node7551;
	wire [4-1:0] node7552;
	wire [4-1:0] node7553;
	wire [4-1:0] node7556;
	wire [4-1:0] node7557;
	wire [4-1:0] node7561;
	wire [4-1:0] node7562;
	wire [4-1:0] node7564;
	wire [4-1:0] node7567;
	wire [4-1:0] node7570;
	wire [4-1:0] node7571;
	wire [4-1:0] node7572;
	wire [4-1:0] node7573;
	wire [4-1:0] node7576;
	wire [4-1:0] node7578;
	wire [4-1:0] node7579;
	wire [4-1:0] node7580;
	wire [4-1:0] node7585;
	wire [4-1:0] node7586;
	wire [4-1:0] node7589;
	wire [4-1:0] node7591;
	wire [4-1:0] node7592;
	wire [4-1:0] node7596;
	wire [4-1:0] node7597;
	wire [4-1:0] node7598;
	wire [4-1:0] node7599;
	wire [4-1:0] node7600;
	wire [4-1:0] node7604;
	wire [4-1:0] node7607;
	wire [4-1:0] node7608;
	wire [4-1:0] node7609;
	wire [4-1:0] node7610;
	wire [4-1:0] node7614;
	wire [4-1:0] node7617;
	wire [4-1:0] node7618;
	wire [4-1:0] node7622;
	wire [4-1:0] node7623;
	wire [4-1:0] node7624;
	wire [4-1:0] node7627;
	wire [4-1:0] node7630;
	wire [4-1:0] node7632;
	wire [4-1:0] node7635;
	wire [4-1:0] node7636;
	wire [4-1:0] node7637;
	wire [4-1:0] node7638;
	wire [4-1:0] node7639;
	wire [4-1:0] node7640;
	wire [4-1:0] node7641;
	wire [4-1:0] node7642;
	wire [4-1:0] node7643;
	wire [4-1:0] node7646;
	wire [4-1:0] node7649;
	wire [4-1:0] node7650;
	wire [4-1:0] node7654;
	wire [4-1:0] node7655;
	wire [4-1:0] node7656;
	wire [4-1:0] node7657;
	wire [4-1:0] node7660;
	wire [4-1:0] node7664;
	wire [4-1:0] node7665;
	wire [4-1:0] node7669;
	wire [4-1:0] node7670;
	wire [4-1:0] node7672;
	wire [4-1:0] node7673;
	wire [4-1:0] node7675;
	wire [4-1:0] node7679;
	wire [4-1:0] node7680;
	wire [4-1:0] node7681;
	wire [4-1:0] node7683;
	wire [4-1:0] node7686;
	wire [4-1:0] node7689;
	wire [4-1:0] node7691;
	wire [4-1:0] node7693;
	wire [4-1:0] node7696;
	wire [4-1:0] node7697;
	wire [4-1:0] node7698;
	wire [4-1:0] node7699;
	wire [4-1:0] node7700;
	wire [4-1:0] node7701;
	wire [4-1:0] node7704;
	wire [4-1:0] node7709;
	wire [4-1:0] node7711;
	wire [4-1:0] node7713;
	wire [4-1:0] node7716;
	wire [4-1:0] node7717;
	wire [4-1:0] node7718;
	wire [4-1:0] node7719;
	wire [4-1:0] node7720;
	wire [4-1:0] node7724;
	wire [4-1:0] node7726;
	wire [4-1:0] node7729;
	wire [4-1:0] node7731;
	wire [4-1:0] node7734;
	wire [4-1:0] node7735;
	wire [4-1:0] node7738;
	wire [4-1:0] node7739;
	wire [4-1:0] node7743;
	wire [4-1:0] node7744;
	wire [4-1:0] node7745;
	wire [4-1:0] node7746;
	wire [4-1:0] node7747;
	wire [4-1:0] node7748;
	wire [4-1:0] node7752;
	wire [4-1:0] node7753;
	wire [4-1:0] node7756;
	wire [4-1:0] node7758;
	wire [4-1:0] node7761;
	wire [4-1:0] node7762;
	wire [4-1:0] node7763;
	wire [4-1:0] node7767;
	wire [4-1:0] node7768;
	wire [4-1:0] node7769;
	wire [4-1:0] node7773;
	wire [4-1:0] node7774;
	wire [4-1:0] node7778;
	wire [4-1:0] node7779;
	wire [4-1:0] node7780;
	wire [4-1:0] node7781;
	wire [4-1:0] node7785;
	wire [4-1:0] node7786;
	wire [4-1:0] node7789;
	wire [4-1:0] node7792;
	wire [4-1:0] node7793;
	wire [4-1:0] node7795;
	wire [4-1:0] node7798;
	wire [4-1:0] node7799;
	wire [4-1:0] node7803;
	wire [4-1:0] node7804;
	wire [4-1:0] node7805;
	wire [4-1:0] node7806;
	wire [4-1:0] node7807;
	wire [4-1:0] node7811;
	wire [4-1:0] node7813;
	wire [4-1:0] node7816;
	wire [4-1:0] node7817;
	wire [4-1:0] node7820;
	wire [4-1:0] node7823;
	wire [4-1:0] node7824;
	wire [4-1:0] node7825;
	wire [4-1:0] node7826;
	wire [4-1:0] node7827;
	wire [4-1:0] node7831;
	wire [4-1:0] node7835;
	wire [4-1:0] node7837;
	wire [4-1:0] node7839;
	wire [4-1:0] node7840;
	wire [4-1:0] node7844;
	wire [4-1:0] node7845;
	wire [4-1:0] node7846;
	wire [4-1:0] node7847;
	wire [4-1:0] node7848;
	wire [4-1:0] node7849;
	wire [4-1:0] node7851;
	wire [4-1:0] node7852;
	wire [4-1:0] node7858;
	wire [4-1:0] node7859;
	wire [4-1:0] node7860;
	wire [4-1:0] node7862;
	wire [4-1:0] node7865;
	wire [4-1:0] node7867;
	wire [4-1:0] node7868;
	wire [4-1:0] node7872;
	wire [4-1:0] node7873;
	wire [4-1:0] node7874;
	wire [4-1:0] node7877;
	wire [4-1:0] node7879;
	wire [4-1:0] node7882;
	wire [4-1:0] node7884;
	wire [4-1:0] node7887;
	wire [4-1:0] node7888;
	wire [4-1:0] node7889;
	wire [4-1:0] node7890;
	wire [4-1:0] node7891;
	wire [4-1:0] node7892;
	wire [4-1:0] node7896;
	wire [4-1:0] node7898;
	wire [4-1:0] node7901;
	wire [4-1:0] node7903;
	wire [4-1:0] node7906;
	wire [4-1:0] node7907;
	wire [4-1:0] node7908;
	wire [4-1:0] node7911;
	wire [4-1:0] node7914;
	wire [4-1:0] node7916;
	wire [4-1:0] node7919;
	wire [4-1:0] node7920;
	wire [4-1:0] node7921;
	wire [4-1:0] node7924;
	wire [4-1:0] node7926;
	wire [4-1:0] node7927;
	wire [4-1:0] node7930;
	wire [4-1:0] node7933;
	wire [4-1:0] node7934;
	wire [4-1:0] node7935;
	wire [4-1:0] node7939;
	wire [4-1:0] node7941;
	wire [4-1:0] node7944;
	wire [4-1:0] node7945;
	wire [4-1:0] node7946;
	wire [4-1:0] node7947;
	wire [4-1:0] node7948;
	wire [4-1:0] node7949;
	wire [4-1:0] node7952;
	wire [4-1:0] node7953;
	wire [4-1:0] node7958;
	wire [4-1:0] node7959;
	wire [4-1:0] node7962;
	wire [4-1:0] node7963;
	wire [4-1:0] node7964;
	wire [4-1:0] node7969;
	wire [4-1:0] node7970;
	wire [4-1:0] node7971;
	wire [4-1:0] node7972;
	wire [4-1:0] node7975;
	wire [4-1:0] node7976;
	wire [4-1:0] node7980;
	wire [4-1:0] node7983;
	wire [4-1:0] node7984;
	wire [4-1:0] node7985;
	wire [4-1:0] node7988;
	wire [4-1:0] node7991;
	wire [4-1:0] node7993;
	wire [4-1:0] node7994;
	wire [4-1:0] node7998;
	wire [4-1:0] node7999;
	wire [4-1:0] node8000;
	wire [4-1:0] node8001;
	wire [4-1:0] node8004;
	wire [4-1:0] node8005;
	wire [4-1:0] node8008;
	wire [4-1:0] node8009;
	wire [4-1:0] node8012;
	wire [4-1:0] node8015;
	wire [4-1:0] node8017;
	wire [4-1:0] node8018;
	wire [4-1:0] node8019;
	wire [4-1:0] node8023;
	wire [4-1:0] node8026;
	wire [4-1:0] node8027;
	wire [4-1:0] node8030;
	wire [4-1:0] node8031;
	wire [4-1:0] node8035;
	wire [4-1:0] node8036;
	wire [4-1:0] node8037;
	wire [4-1:0] node8038;
	wire [4-1:0] node8039;
	wire [4-1:0] node8040;
	wire [4-1:0] node8041;
	wire [4-1:0] node8042;
	wire [4-1:0] node8046;
	wire [4-1:0] node8048;
	wire [4-1:0] node8051;
	wire [4-1:0] node8052;
	wire [4-1:0] node8054;
	wire [4-1:0] node8055;
	wire [4-1:0] node8060;
	wire [4-1:0] node8061;
	wire [4-1:0] node8062;
	wire [4-1:0] node8063;
	wire [4-1:0] node8067;
	wire [4-1:0] node8069;
	wire [4-1:0] node8072;
	wire [4-1:0] node8073;
	wire [4-1:0] node8077;
	wire [4-1:0] node8078;
	wire [4-1:0] node8079;
	wire [4-1:0] node8080;
	wire [4-1:0] node8081;
	wire [4-1:0] node8086;
	wire [4-1:0] node8087;
	wire [4-1:0] node8089;
	wire [4-1:0] node8091;
	wire [4-1:0] node8094;
	wire [4-1:0] node8097;
	wire [4-1:0] node8098;
	wire [4-1:0] node8099;
	wire [4-1:0] node8101;
	wire [4-1:0] node8105;
	wire [4-1:0] node8106;
	wire [4-1:0] node8108;
	wire [4-1:0] node8111;
	wire [4-1:0] node8113;
	wire [4-1:0] node8116;
	wire [4-1:0] node8117;
	wire [4-1:0] node8118;
	wire [4-1:0] node8119;
	wire [4-1:0] node8120;
	wire [4-1:0] node8122;
	wire [4-1:0] node8125;
	wire [4-1:0] node8126;
	wire [4-1:0] node8130;
	wire [4-1:0] node8131;
	wire [4-1:0] node8132;
	wire [4-1:0] node8136;
	wire [4-1:0] node8137;
	wire [4-1:0] node8140;
	wire [4-1:0] node8143;
	wire [4-1:0] node8144;
	wire [4-1:0] node8145;
	wire [4-1:0] node8149;
	wire [4-1:0] node8150;
	wire [4-1:0] node8152;
	wire [4-1:0] node8155;
	wire [4-1:0] node8158;
	wire [4-1:0] node8159;
	wire [4-1:0] node8160;
	wire [4-1:0] node8162;
	wire [4-1:0] node8165;
	wire [4-1:0] node8166;
	wire [4-1:0] node8170;
	wire [4-1:0] node8171;
	wire [4-1:0] node8173;
	wire [4-1:0] node8174;
	wire [4-1:0] node8176;
	wire [4-1:0] node8180;
	wire [4-1:0] node8182;
	wire [4-1:0] node8184;
	wire [4-1:0] node8187;
	wire [4-1:0] node8188;
	wire [4-1:0] node8189;
	wire [4-1:0] node8190;
	wire [4-1:0] node8191;
	wire [4-1:0] node8192;
	wire [4-1:0] node8193;
	wire [4-1:0] node8197;
	wire [4-1:0] node8200;
	wire [4-1:0] node8203;
	wire [4-1:0] node8204;
	wire [4-1:0] node8205;
	wire [4-1:0] node8207;
	wire [4-1:0] node8209;
	wire [4-1:0] node8213;
	wire [4-1:0] node8214;
	wire [4-1:0] node8217;
	wire [4-1:0] node8219;
	wire [4-1:0] node8222;
	wire [4-1:0] node8223;
	wire [4-1:0] node8224;
	wire [4-1:0] node8226;
	wire [4-1:0] node8228;
	wire [4-1:0] node8231;
	wire [4-1:0] node8232;
	wire [4-1:0] node8234;
	wire [4-1:0] node8237;
	wire [4-1:0] node8238;
	wire [4-1:0] node8242;
	wire [4-1:0] node8243;
	wire [4-1:0] node8244;
	wire [4-1:0] node8247;
	wire [4-1:0] node8248;
	wire [4-1:0] node8249;
	wire [4-1:0] node8254;
	wire [4-1:0] node8256;
	wire [4-1:0] node8259;
	wire [4-1:0] node8260;
	wire [4-1:0] node8261;
	wire [4-1:0] node8262;
	wire [4-1:0] node8263;
	wire [4-1:0] node8266;
	wire [4-1:0] node8269;
	wire [4-1:0] node8271;
	wire [4-1:0] node8272;
	wire [4-1:0] node8274;
	wire [4-1:0] node8277;
	wire [4-1:0] node8278;
	wire [4-1:0] node8282;
	wire [4-1:0] node8283;
	wire [4-1:0] node8284;
	wire [4-1:0] node8289;
	wire [4-1:0] node8290;
	wire [4-1:0] node8291;
	wire [4-1:0] node8294;
	wire [4-1:0] node8296;
	wire [4-1:0] node8299;
	wire [4-1:0] node8300;
	wire [4-1:0] node8301;
	wire [4-1:0] node8302;
	wire [4-1:0] node8306;
	wire [4-1:0] node8310;
	wire [4-1:0] node8311;
	wire [4-1:0] node8312;
	wire [4-1:0] node8313;
	wire [4-1:0] node8314;
	wire [4-1:0] node8315;
	wire [4-1:0] node8316;
	wire [4-1:0] node8317;
	wire [4-1:0] node8318;
	wire [4-1:0] node8319;
	wire [4-1:0] node8320;
	wire [4-1:0] node8322;
	wire [4-1:0] node8326;
	wire [4-1:0] node8329;
	wire [4-1:0] node8330;
	wire [4-1:0] node8333;
	wire [4-1:0] node8334;
	wire [4-1:0] node8338;
	wire [4-1:0] node8339;
	wire [4-1:0] node8340;
	wire [4-1:0] node8344;
	wire [4-1:0] node8347;
	wire [4-1:0] node8348;
	wire [4-1:0] node8349;
	wire [4-1:0] node8350;
	wire [4-1:0] node8351;
	wire [4-1:0] node8356;
	wire [4-1:0] node8357;
	wire [4-1:0] node8359;
	wire [4-1:0] node8362;
	wire [4-1:0] node8365;
	wire [4-1:0] node8366;
	wire [4-1:0] node8368;
	wire [4-1:0] node8369;
	wire [4-1:0] node8370;
	wire [4-1:0] node8375;
	wire [4-1:0] node8376;
	wire [4-1:0] node8377;
	wire [4-1:0] node8380;
	wire [4-1:0] node8383;
	wire [4-1:0] node8386;
	wire [4-1:0] node8387;
	wire [4-1:0] node8388;
	wire [4-1:0] node8389;
	wire [4-1:0] node8390;
	wire [4-1:0] node8391;
	wire [4-1:0] node8394;
	wire [4-1:0] node8397;
	wire [4-1:0] node8399;
	wire [4-1:0] node8402;
	wire [4-1:0] node8404;
	wire [4-1:0] node8407;
	wire [4-1:0] node8408;
	wire [4-1:0] node8409;
	wire [4-1:0] node8411;
	wire [4-1:0] node8414;
	wire [4-1:0] node8417;
	wire [4-1:0] node8418;
	wire [4-1:0] node8419;
	wire [4-1:0] node8423;
	wire [4-1:0] node8425;
	wire [4-1:0] node8428;
	wire [4-1:0] node8429;
	wire [4-1:0] node8430;
	wire [4-1:0] node8431;
	wire [4-1:0] node8433;
	wire [4-1:0] node8435;
	wire [4-1:0] node8438;
	wire [4-1:0] node8441;
	wire [4-1:0] node8442;
	wire [4-1:0] node8445;
	wire [4-1:0] node8446;
	wire [4-1:0] node8449;
	wire [4-1:0] node8452;
	wire [4-1:0] node8453;
	wire [4-1:0] node8454;
	wire [4-1:0] node8457;
	wire [4-1:0] node8458;
	wire [4-1:0] node8459;
	wire [4-1:0] node8464;
	wire [4-1:0] node8467;
	wire [4-1:0] node8468;
	wire [4-1:0] node8469;
	wire [4-1:0] node8470;
	wire [4-1:0] node8471;
	wire [4-1:0] node8472;
	wire [4-1:0] node8473;
	wire [4-1:0] node8477;
	wire [4-1:0] node8480;
	wire [4-1:0] node8481;
	wire [4-1:0] node8482;
	wire [4-1:0] node8484;
	wire [4-1:0] node8487;
	wire [4-1:0] node8488;
	wire [4-1:0] node8492;
	wire [4-1:0] node8493;
	wire [4-1:0] node8496;
	wire [4-1:0] node8498;
	wire [4-1:0] node8501;
	wire [4-1:0] node8502;
	wire [4-1:0] node8503;
	wire [4-1:0] node8504;
	wire [4-1:0] node8505;
	wire [4-1:0] node8509;
	wire [4-1:0] node8511;
	wire [4-1:0] node8514;
	wire [4-1:0] node8515;
	wire [4-1:0] node8517;
	wire [4-1:0] node8520;
	wire [4-1:0] node8522;
	wire [4-1:0] node8525;
	wire [4-1:0] node8526;
	wire [4-1:0] node8530;
	wire [4-1:0] node8531;
	wire [4-1:0] node8532;
	wire [4-1:0] node8533;
	wire [4-1:0] node8535;
	wire [4-1:0] node8538;
	wire [4-1:0] node8540;
	wire [4-1:0] node8543;
	wire [4-1:0] node8545;
	wire [4-1:0] node8547;
	wire [4-1:0] node8549;
	wire [4-1:0] node8552;
	wire [4-1:0] node8553;
	wire [4-1:0] node8556;
	wire [4-1:0] node8557;
	wire [4-1:0] node8559;
	wire [4-1:0] node8563;
	wire [4-1:0] node8564;
	wire [4-1:0] node8565;
	wire [4-1:0] node8566;
	wire [4-1:0] node8567;
	wire [4-1:0] node8568;
	wire [4-1:0] node8573;
	wire [4-1:0] node8574;
	wire [4-1:0] node8575;
	wire [4-1:0] node8580;
	wire [4-1:0] node8581;
	wire [4-1:0] node8582;
	wire [4-1:0] node8584;
	wire [4-1:0] node8587;
	wire [4-1:0] node8590;
	wire [4-1:0] node8591;
	wire [4-1:0] node8594;
	wire [4-1:0] node8595;
	wire [4-1:0] node8599;
	wire [4-1:0] node8600;
	wire [4-1:0] node8601;
	wire [4-1:0] node8603;
	wire [4-1:0] node8606;
	wire [4-1:0] node8607;
	wire [4-1:0] node8608;
	wire [4-1:0] node8609;
	wire [4-1:0] node8614;
	wire [4-1:0] node8615;
	wire [4-1:0] node8616;
	wire [4-1:0] node8620;
	wire [4-1:0] node8621;
	wire [4-1:0] node8625;
	wire [4-1:0] node8626;
	wire [4-1:0] node8628;
	wire [4-1:0] node8630;
	wire [4-1:0] node8632;
	wire [4-1:0] node8635;
	wire [4-1:0] node8637;
	wire [4-1:0] node8638;
	wire [4-1:0] node8640;
	wire [4-1:0] node8643;
	wire [4-1:0] node8646;
	wire [4-1:0] node8647;
	wire [4-1:0] node8648;
	wire [4-1:0] node8649;
	wire [4-1:0] node8650;
	wire [4-1:0] node8651;
	wire [4-1:0] node8652;
	wire [4-1:0] node8653;
	wire [4-1:0] node8654;
	wire [4-1:0] node8657;
	wire [4-1:0] node8661;
	wire [4-1:0] node8662;
	wire [4-1:0] node8666;
	wire [4-1:0] node8667;
	wire [4-1:0] node8668;
	wire [4-1:0] node8672;
	wire [4-1:0] node8675;
	wire [4-1:0] node8676;
	wire [4-1:0] node8677;
	wire [4-1:0] node8678;
	wire [4-1:0] node8682;
	wire [4-1:0] node8683;
	wire [4-1:0] node8684;
	wire [4-1:0] node8688;
	wire [4-1:0] node8691;
	wire [4-1:0] node8692;
	wire [4-1:0] node8694;
	wire [4-1:0] node8697;
	wire [4-1:0] node8698;
	wire [4-1:0] node8702;
	wire [4-1:0] node8703;
	wire [4-1:0] node8704;
	wire [4-1:0] node8705;
	wire [4-1:0] node8706;
	wire [4-1:0] node8710;
	wire [4-1:0] node8712;
	wire [4-1:0] node8715;
	wire [4-1:0] node8718;
	wire [4-1:0] node8719;
	wire [4-1:0] node8720;
	wire [4-1:0] node8721;
	wire [4-1:0] node8722;
	wire [4-1:0] node8726;
	wire [4-1:0] node8729;
	wire [4-1:0] node8732;
	wire [4-1:0] node8733;
	wire [4-1:0] node8736;
	wire [4-1:0] node8739;
	wire [4-1:0] node8740;
	wire [4-1:0] node8741;
	wire [4-1:0] node8742;
	wire [4-1:0] node8744;
	wire [4-1:0] node8747;
	wire [4-1:0] node8748;
	wire [4-1:0] node8749;
	wire [4-1:0] node8753;
	wire [4-1:0] node8755;
	wire [4-1:0] node8756;
	wire [4-1:0] node8760;
	wire [4-1:0] node8761;
	wire [4-1:0] node8763;
	wire [4-1:0] node8764;
	wire [4-1:0] node8768;
	wire [4-1:0] node8770;
	wire [4-1:0] node8771;
	wire [4-1:0] node8775;
	wire [4-1:0] node8776;
	wire [4-1:0] node8777;
	wire [4-1:0] node8779;
	wire [4-1:0] node8782;
	wire [4-1:0] node8785;
	wire [4-1:0] node8786;
	wire [4-1:0] node8787;
	wire [4-1:0] node8791;
	wire [4-1:0] node8793;
	wire [4-1:0] node8796;
	wire [4-1:0] node8797;
	wire [4-1:0] node8798;
	wire [4-1:0] node8799;
	wire [4-1:0] node8800;
	wire [4-1:0] node8801;
	wire [4-1:0] node8803;
	wire [4-1:0] node8806;
	wire [4-1:0] node8808;
	wire [4-1:0] node8811;
	wire [4-1:0] node8813;
	wire [4-1:0] node8814;
	wire [4-1:0] node8815;
	wire [4-1:0] node8820;
	wire [4-1:0] node8821;
	wire [4-1:0] node8822;
	wire [4-1:0] node8825;
	wire [4-1:0] node8827;
	wire [4-1:0] node8828;
	wire [4-1:0] node8833;
	wire [4-1:0] node8834;
	wire [4-1:0] node8835;
	wire [4-1:0] node8838;
	wire [4-1:0] node8840;
	wire [4-1:0] node8841;
	wire [4-1:0] node8842;
	wire [4-1:0] node8846;
	wire [4-1:0] node8849;
	wire [4-1:0] node8850;
	wire [4-1:0] node8851;
	wire [4-1:0] node8852;
	wire [4-1:0] node8857;
	wire [4-1:0] node8858;
	wire [4-1:0] node8862;
	wire [4-1:0] node8863;
	wire [4-1:0] node8864;
	wire [4-1:0] node8865;
	wire [4-1:0] node8866;
	wire [4-1:0] node8868;
	wire [4-1:0] node8871;
	wire [4-1:0] node8875;
	wire [4-1:0] node8876;
	wire [4-1:0] node8877;
	wire [4-1:0] node8879;
	wire [4-1:0] node8881;
	wire [4-1:0] node8884;
	wire [4-1:0] node8886;
	wire [4-1:0] node8889;
	wire [4-1:0] node8890;
	wire [4-1:0] node8894;
	wire [4-1:0] node8895;
	wire [4-1:0] node8897;
	wire [4-1:0] node8898;
	wire [4-1:0] node8902;
	wire [4-1:0] node8903;
	wire [4-1:0] node8904;
	wire [4-1:0] node8905;
	wire [4-1:0] node8909;
	wire [4-1:0] node8912;
	wire [4-1:0] node8913;
	wire [4-1:0] node8914;
	wire [4-1:0] node8918;
	wire [4-1:0] node8920;
	wire [4-1:0] node8923;
	wire [4-1:0] node8924;
	wire [4-1:0] node8925;
	wire [4-1:0] node8926;
	wire [4-1:0] node8927;
	wire [4-1:0] node8928;
	wire [4-1:0] node8929;
	wire [4-1:0] node8932;
	wire [4-1:0] node8933;
	wire [4-1:0] node8936;
	wire [4-1:0] node8937;
	wire [4-1:0] node8940;
	wire [4-1:0] node8943;
	wire [4-1:0] node8944;
	wire [4-1:0] node8945;
	wire [4-1:0] node8946;
	wire [4-1:0] node8951;
	wire [4-1:0] node8953;
	wire [4-1:0] node8954;
	wire [4-1:0] node8955;
	wire [4-1:0] node8960;
	wire [4-1:0] node8961;
	wire [4-1:0] node8962;
	wire [4-1:0] node8963;
	wire [4-1:0] node8966;
	wire [4-1:0] node8969;
	wire [4-1:0] node8970;
	wire [4-1:0] node8971;
	wire [4-1:0] node8975;
	wire [4-1:0] node8976;
	wire [4-1:0] node8977;
	wire [4-1:0] node8982;
	wire [4-1:0] node8983;
	wire [4-1:0] node8984;
	wire [4-1:0] node8986;
	wire [4-1:0] node8989;
	wire [4-1:0] node8992;
	wire [4-1:0] node8994;
	wire [4-1:0] node8996;
	wire [4-1:0] node8998;
	wire [4-1:0] node9001;
	wire [4-1:0] node9002;
	wire [4-1:0] node9003;
	wire [4-1:0] node9004;
	wire [4-1:0] node9005;
	wire [4-1:0] node9007;
	wire [4-1:0] node9009;
	wire [4-1:0] node9012;
	wire [4-1:0] node9014;
	wire [4-1:0] node9015;
	wire [4-1:0] node9019;
	wire [4-1:0] node9020;
	wire [4-1:0] node9022;
	wire [4-1:0] node9023;
	wire [4-1:0] node9027;
	wire [4-1:0] node9030;
	wire [4-1:0] node9031;
	wire [4-1:0] node9032;
	wire [4-1:0] node9033;
	wire [4-1:0] node9037;
	wire [4-1:0] node9038;
	wire [4-1:0] node9041;
	wire [4-1:0] node9044;
	wire [4-1:0] node9046;
	wire [4-1:0] node9047;
	wire [4-1:0] node9050;
	wire [4-1:0] node9053;
	wire [4-1:0] node9054;
	wire [4-1:0] node9055;
	wire [4-1:0] node9057;
	wire [4-1:0] node9058;
	wire [4-1:0] node9062;
	wire [4-1:0] node9063;
	wire [4-1:0] node9066;
	wire [4-1:0] node9068;
	wire [4-1:0] node9069;
	wire [4-1:0] node9073;
	wire [4-1:0] node9074;
	wire [4-1:0] node9075;
	wire [4-1:0] node9076;
	wire [4-1:0] node9079;
	wire [4-1:0] node9082;
	wire [4-1:0] node9084;
	wire [4-1:0] node9087;
	wire [4-1:0] node9088;
	wire [4-1:0] node9091;
	wire [4-1:0] node9092;
	wire [4-1:0] node9094;
	wire [4-1:0] node9098;
	wire [4-1:0] node9099;
	wire [4-1:0] node9100;
	wire [4-1:0] node9101;
	wire [4-1:0] node9102;
	wire [4-1:0] node9103;
	wire [4-1:0] node9106;
	wire [4-1:0] node9109;
	wire [4-1:0] node9110;
	wire [4-1:0] node9113;
	wire [4-1:0] node9114;
	wire [4-1:0] node9118;
	wire [4-1:0] node9119;
	wire [4-1:0] node9120;
	wire [4-1:0] node9122;
	wire [4-1:0] node9126;
	wire [4-1:0] node9127;
	wire [4-1:0] node9129;
	wire [4-1:0] node9131;
	wire [4-1:0] node9134;
	wire [4-1:0] node9136;
	wire [4-1:0] node9137;
	wire [4-1:0] node9140;
	wire [4-1:0] node9143;
	wire [4-1:0] node9144;
	wire [4-1:0] node9145;
	wire [4-1:0] node9146;
	wire [4-1:0] node9147;
	wire [4-1:0] node9151;
	wire [4-1:0] node9153;
	wire [4-1:0] node9156;
	wire [4-1:0] node9157;
	wire [4-1:0] node9160;
	wire [4-1:0] node9161;
	wire [4-1:0] node9165;
	wire [4-1:0] node9166;
	wire [4-1:0] node9167;
	wire [4-1:0] node9169;
	wire [4-1:0] node9172;
	wire [4-1:0] node9175;
	wire [4-1:0] node9176;
	wire [4-1:0] node9178;
	wire [4-1:0] node9181;
	wire [4-1:0] node9183;
	wire [4-1:0] node9186;
	wire [4-1:0] node9187;
	wire [4-1:0] node9188;
	wire [4-1:0] node9189;
	wire [4-1:0] node9190;
	wire [4-1:0] node9191;
	wire [4-1:0] node9194;
	wire [4-1:0] node9196;
	wire [4-1:0] node9199;
	wire [4-1:0] node9200;
	wire [4-1:0] node9202;
	wire [4-1:0] node9206;
	wire [4-1:0] node9207;
	wire [4-1:0] node9209;
	wire [4-1:0] node9210;
	wire [4-1:0] node9214;
	wire [4-1:0] node9215;
	wire [4-1:0] node9218;
	wire [4-1:0] node9219;
	wire [4-1:0] node9223;
	wire [4-1:0] node9224;
	wire [4-1:0] node9225;
	wire [4-1:0] node9229;
	wire [4-1:0] node9231;
	wire [4-1:0] node9232;
	wire [4-1:0] node9236;
	wire [4-1:0] node9237;
	wire [4-1:0] node9238;
	wire [4-1:0] node9239;
	wire [4-1:0] node9242;
	wire [4-1:0] node9244;
	wire [4-1:0] node9245;
	wire [4-1:0] node9249;
	wire [4-1:0] node9250;
	wire [4-1:0] node9252;
	wire [4-1:0] node9254;
	wire [4-1:0] node9258;
	wire [4-1:0] node9259;
	wire [4-1:0] node9260;
	wire [4-1:0] node9261;
	wire [4-1:0] node9266;
	wire [4-1:0] node9267;
	wire [4-1:0] node9269;
	wire [4-1:0] node9272;
	wire [4-1:0] node9273;
	wire [4-1:0] node9277;
	wire [4-1:0] node9278;
	wire [4-1:0] node9279;
	wire [4-1:0] node9280;
	wire [4-1:0] node9281;
	wire [4-1:0] node9282;
	wire [4-1:0] node9284;
	wire [4-1:0] node9287;
	wire [4-1:0] node9288;
	wire [4-1:0] node9290;
	wire [4-1:0] node9294;
	wire [4-1:0] node9295;
	wire [4-1:0] node9296;
	wire [4-1:0] node9297;
	wire [4-1:0] node9301;
	wire [4-1:0] node9302;
	wire [4-1:0] node9306;
	wire [4-1:0] node9307;
	wire [4-1:0] node9308;
	wire [4-1:0] node9309;
	wire [4-1:0] node9315;
	wire [4-1:0] node9316;
	wire [4-1:0] node9317;
	wire [4-1:0] node9318;
	wire [4-1:0] node9319;
	wire [4-1:0] node9321;
	wire [4-1:0] node9325;
	wire [4-1:0] node9326;
	wire [4-1:0] node9327;
	wire [4-1:0] node9330;
	wire [4-1:0] node9333;
	wire [4-1:0] node9336;
	wire [4-1:0] node9337;
	wire [4-1:0] node9338;
	wire [4-1:0] node9342;
	wire [4-1:0] node9343;
	wire [4-1:0] node9347;
	wire [4-1:0] node9348;
	wire [4-1:0] node9350;
	wire [4-1:0] node9353;
	wire [4-1:0] node9354;
	wire [4-1:0] node9358;
	wire [4-1:0] node9359;
	wire [4-1:0] node9360;
	wire [4-1:0] node9361;
	wire [4-1:0] node9363;
	wire [4-1:0] node9366;
	wire [4-1:0] node9367;
	wire [4-1:0] node9369;
	wire [4-1:0] node9372;
	wire [4-1:0] node9374;
	wire [4-1:0] node9377;
	wire [4-1:0] node9378;
	wire [4-1:0] node9380;
	wire [4-1:0] node9381;
	wire [4-1:0] node9383;
	wire [4-1:0] node9387;
	wire [4-1:0] node9388;
	wire [4-1:0] node9389;
	wire [4-1:0] node9393;
	wire [4-1:0] node9395;
	wire [4-1:0] node9396;
	wire [4-1:0] node9400;
	wire [4-1:0] node9401;
	wire [4-1:0] node9402;
	wire [4-1:0] node9403;
	wire [4-1:0] node9406;
	wire [4-1:0] node9410;
	wire [4-1:0] node9411;
	wire [4-1:0] node9412;
	wire [4-1:0] node9414;
	wire [4-1:0] node9418;
	wire [4-1:0] node9419;
	wire [4-1:0] node9423;
	wire [4-1:0] node9424;
	wire [4-1:0] node9425;
	wire [4-1:0] node9426;
	wire [4-1:0] node9427;
	wire [4-1:0] node9429;
	wire [4-1:0] node9431;
	wire [4-1:0] node9434;
	wire [4-1:0] node9435;
	wire [4-1:0] node9437;
	wire [4-1:0] node9441;
	wire [4-1:0] node9442;
	wire [4-1:0] node9443;
	wire [4-1:0] node9445;
	wire [4-1:0] node9449;
	wire [4-1:0] node9451;
	wire [4-1:0] node9452;
	wire [4-1:0] node9453;
	wire [4-1:0] node9456;
	wire [4-1:0] node9460;
	wire [4-1:0] node9461;
	wire [4-1:0] node9462;
	wire [4-1:0] node9463;
	wire [4-1:0] node9466;
	wire [4-1:0] node9467;
	wire [4-1:0] node9471;
	wire [4-1:0] node9472;
	wire [4-1:0] node9476;
	wire [4-1:0] node9477;
	wire [4-1:0] node9479;
	wire [4-1:0] node9481;
	wire [4-1:0] node9484;
	wire [4-1:0] node9486;
	wire [4-1:0] node9489;
	wire [4-1:0] node9490;
	wire [4-1:0] node9491;
	wire [4-1:0] node9492;
	wire [4-1:0] node9493;
	wire [4-1:0] node9494;
	wire [4-1:0] node9497;
	wire [4-1:0] node9500;
	wire [4-1:0] node9501;
	wire [4-1:0] node9505;
	wire [4-1:0] node9506;
	wire [4-1:0] node9507;
	wire [4-1:0] node9508;
	wire [4-1:0] node9511;
	wire [4-1:0] node9516;
	wire [4-1:0] node9517;
	wire [4-1:0] node9518;
	wire [4-1:0] node9520;
	wire [4-1:0] node9523;
	wire [4-1:0] node9524;
	wire [4-1:0] node9527;
	wire [4-1:0] node9530;
	wire [4-1:0] node9531;
	wire [4-1:0] node9532;
	wire [4-1:0] node9536;
	wire [4-1:0] node9539;
	wire [4-1:0] node9540;
	wire [4-1:0] node9542;
	wire [4-1:0] node9543;
	wire [4-1:0] node9546;
	wire [4-1:0] node9547;
	wire [4-1:0] node9551;
	wire [4-1:0] node9552;
	wire [4-1:0] node9553;
	wire [4-1:0] node9556;
	wire [4-1:0] node9558;
	wire [4-1:0] node9559;
	wire [4-1:0] node9563;
	wire [4-1:0] node9564;
	wire [4-1:0] node9565;
	wire [4-1:0] node9569;
	wire [4-1:0] node9572;
	wire [4-1:0] node9573;
	wire [4-1:0] node9574;
	wire [4-1:0] node9575;
	wire [4-1:0] node9576;
	wire [4-1:0] node9577;
	wire [4-1:0] node9578;
	wire [4-1:0] node9579;
	wire [4-1:0] node9581;
	wire [4-1:0] node9583;
	wire [4-1:0] node9586;
	wire [4-1:0] node9587;
	wire [4-1:0] node9589;
	wire [4-1:0] node9592;
	wire [4-1:0] node9594;
	wire [4-1:0] node9597;
	wire [4-1:0] node9598;
	wire [4-1:0] node9599;
	wire [4-1:0] node9603;
	wire [4-1:0] node9604;
	wire [4-1:0] node9606;
	wire [4-1:0] node9610;
	wire [4-1:0] node9611;
	wire [4-1:0] node9612;
	wire [4-1:0] node9613;
	wire [4-1:0] node9614;
	wire [4-1:0] node9618;
	wire [4-1:0] node9619;
	wire [4-1:0] node9621;
	wire [4-1:0] node9625;
	wire [4-1:0] node9626;
	wire [4-1:0] node9627;
	wire [4-1:0] node9630;
	wire [4-1:0] node9632;
	wire [4-1:0] node9635;
	wire [4-1:0] node9637;
	wire [4-1:0] node9638;
	wire [4-1:0] node9642;
	wire [4-1:0] node9643;
	wire [4-1:0] node9644;
	wire [4-1:0] node9645;
	wire [4-1:0] node9649;
	wire [4-1:0] node9651;
	wire [4-1:0] node9653;
	wire [4-1:0] node9656;
	wire [4-1:0] node9657;
	wire [4-1:0] node9660;
	wire [4-1:0] node9663;
	wire [4-1:0] node9664;
	wire [4-1:0] node9665;
	wire [4-1:0] node9666;
	wire [4-1:0] node9667;
	wire [4-1:0] node9668;
	wire [4-1:0] node9672;
	wire [4-1:0] node9673;
	wire [4-1:0] node9676;
	wire [4-1:0] node9677;
	wire [4-1:0] node9681;
	wire [4-1:0] node9682;
	wire [4-1:0] node9685;
	wire [4-1:0] node9687;
	wire [4-1:0] node9689;
	wire [4-1:0] node9692;
	wire [4-1:0] node9693;
	wire [4-1:0] node9694;
	wire [4-1:0] node9695;
	wire [4-1:0] node9696;
	wire [4-1:0] node9700;
	wire [4-1:0] node9702;
	wire [4-1:0] node9705;
	wire [4-1:0] node9706;
	wire [4-1:0] node9710;
	wire [4-1:0] node9711;
	wire [4-1:0] node9713;
	wire [4-1:0] node9714;
	wire [4-1:0] node9718;
	wire [4-1:0] node9721;
	wire [4-1:0] node9722;
	wire [4-1:0] node9723;
	wire [4-1:0] node9724;
	wire [4-1:0] node9725;
	wire [4-1:0] node9726;
	wire [4-1:0] node9731;
	wire [4-1:0] node9734;
	wire [4-1:0] node9735;
	wire [4-1:0] node9736;
	wire [4-1:0] node9739;
	wire [4-1:0] node9741;
	wire [4-1:0] node9744;
	wire [4-1:0] node9745;
	wire [4-1:0] node9747;
	wire [4-1:0] node9750;
	wire [4-1:0] node9751;
	wire [4-1:0] node9754;
	wire [4-1:0] node9757;
	wire [4-1:0] node9758;
	wire [4-1:0] node9759;
	wire [4-1:0] node9760;
	wire [4-1:0] node9764;
	wire [4-1:0] node9767;
	wire [4-1:0] node9768;
	wire [4-1:0] node9770;
	wire [4-1:0] node9773;
	wire [4-1:0] node9775;
	wire [4-1:0] node9778;
	wire [4-1:0] node9779;
	wire [4-1:0] node9780;
	wire [4-1:0] node9781;
	wire [4-1:0] node9782;
	wire [4-1:0] node9783;
	wire [4-1:0] node9784;
	wire [4-1:0] node9785;
	wire [4-1:0] node9790;
	wire [4-1:0] node9792;
	wire [4-1:0] node9793;
	wire [4-1:0] node9797;
	wire [4-1:0] node9798;
	wire [4-1:0] node9800;
	wire [4-1:0] node9804;
	wire [4-1:0] node9805;
	wire [4-1:0] node9806;
	wire [4-1:0] node9809;
	wire [4-1:0] node9810;
	wire [4-1:0] node9814;
	wire [4-1:0] node9815;
	wire [4-1:0] node9816;
	wire [4-1:0] node9820;
	wire [4-1:0] node9821;
	wire [4-1:0] node9825;
	wire [4-1:0] node9826;
	wire [4-1:0] node9827;
	wire [4-1:0] node9828;
	wire [4-1:0] node9831;
	wire [4-1:0] node9834;
	wire [4-1:0] node9835;
	wire [4-1:0] node9837;
	wire [4-1:0] node9840;
	wire [4-1:0] node9843;
	wire [4-1:0] node9844;
	wire [4-1:0] node9846;
	wire [4-1:0] node9850;
	wire [4-1:0] node9851;
	wire [4-1:0] node9852;
	wire [4-1:0] node9853;
	wire [4-1:0] node9855;
	wire [4-1:0] node9857;
	wire [4-1:0] node9860;
	wire [4-1:0] node9862;
	wire [4-1:0] node9865;
	wire [4-1:0] node9866;
	wire [4-1:0] node9867;
	wire [4-1:0] node9868;
	wire [4-1:0] node9871;
	wire [4-1:0] node9873;
	wire [4-1:0] node9876;
	wire [4-1:0] node9879;
	wire [4-1:0] node9880;
	wire [4-1:0] node9882;
	wire [4-1:0] node9885;
	wire [4-1:0] node9888;
	wire [4-1:0] node9889;
	wire [4-1:0] node9890;
	wire [4-1:0] node9891;
	wire [4-1:0] node9892;
	wire [4-1:0] node9896;
	wire [4-1:0] node9899;
	wire [4-1:0] node9901;
	wire [4-1:0] node9904;
	wire [4-1:0] node9905;
	wire [4-1:0] node9906;
	wire [4-1:0] node9908;
	wire [4-1:0] node9911;
	wire [4-1:0] node9912;
	wire [4-1:0] node9916;
	wire [4-1:0] node9917;
	wire [4-1:0] node9920;
	wire [4-1:0] node9923;
	wire [4-1:0] node9924;
	wire [4-1:0] node9925;
	wire [4-1:0] node9926;
	wire [4-1:0] node9927;
	wire [4-1:0] node9928;
	wire [4-1:0] node9930;
	wire [4-1:0] node9932;
	wire [4-1:0] node9933;
	wire [4-1:0] node9936;
	wire [4-1:0] node9939;
	wire [4-1:0] node9940;
	wire [4-1:0] node9943;
	wire [4-1:0] node9945;
	wire [4-1:0] node9948;
	wire [4-1:0] node9949;
	wire [4-1:0] node9950;
	wire [4-1:0] node9952;
	wire [4-1:0] node9955;
	wire [4-1:0] node9958;
	wire [4-1:0] node9959;
	wire [4-1:0] node9963;
	wire [4-1:0] node9964;
	wire [4-1:0] node9965;
	wire [4-1:0] node9966;
	wire [4-1:0] node9967;
	wire [4-1:0] node9971;
	wire [4-1:0] node9973;
	wire [4-1:0] node9975;
	wire [4-1:0] node9978;
	wire [4-1:0] node9979;
	wire [4-1:0] node9981;
	wire [4-1:0] node9985;
	wire [4-1:0] node9987;
	wire [4-1:0] node9988;
	wire [4-1:0] node9991;
	wire [4-1:0] node9994;
	wire [4-1:0] node9995;
	wire [4-1:0] node9996;
	wire [4-1:0] node9997;
	wire [4-1:0] node9998;
	wire [4-1:0] node10000;
	wire [4-1:0] node10003;
	wire [4-1:0] node10005;
	wire [4-1:0] node10008;
	wire [4-1:0] node10009;
	wire [4-1:0] node10010;
	wire [4-1:0] node10015;
	wire [4-1:0] node10016;
	wire [4-1:0] node10017;
	wire [4-1:0] node10021;
	wire [4-1:0] node10022;
	wire [4-1:0] node10023;
	wire [4-1:0] node10027;
	wire [4-1:0] node10028;
	wire [4-1:0] node10032;
	wire [4-1:0] node10033;
	wire [4-1:0] node10034;
	wire [4-1:0] node10035;
	wire [4-1:0] node10037;
	wire [4-1:0] node10041;
	wire [4-1:0] node10042;
	wire [4-1:0] node10044;
	wire [4-1:0] node10046;
	wire [4-1:0] node10050;
	wire [4-1:0] node10051;
	wire [4-1:0] node10052;
	wire [4-1:0] node10056;
	wire [4-1:0] node10057;
	wire [4-1:0] node10060;
	wire [4-1:0] node10063;
	wire [4-1:0] node10064;
	wire [4-1:0] node10065;
	wire [4-1:0] node10066;
	wire [4-1:0] node10068;
	wire [4-1:0] node10069;
	wire [4-1:0] node10072;
	wire [4-1:0] node10073;
	wire [4-1:0] node10077;
	wire [4-1:0] node10078;
	wire [4-1:0] node10080;
	wire [4-1:0] node10081;
	wire [4-1:0] node10084;
	wire [4-1:0] node10087;
	wire [4-1:0] node10088;
	wire [4-1:0] node10090;
	wire [4-1:0] node10093;
	wire [4-1:0] node10094;
	wire [4-1:0] node10098;
	wire [4-1:0] node10099;
	wire [4-1:0] node10100;
	wire [4-1:0] node10101;
	wire [4-1:0] node10103;
	wire [4-1:0] node10106;
	wire [4-1:0] node10108;
	wire [4-1:0] node10109;
	wire [4-1:0] node10113;
	wire [4-1:0] node10114;
	wire [4-1:0] node10115;
	wire [4-1:0] node10116;
	wire [4-1:0] node10122;
	wire [4-1:0] node10123;
	wire [4-1:0] node10124;
	wire [4-1:0] node10127;
	wire [4-1:0] node10130;
	wire [4-1:0] node10131;
	wire [4-1:0] node10133;
	wire [4-1:0] node10135;
	wire [4-1:0] node10139;
	wire [4-1:0] node10140;
	wire [4-1:0] node10141;
	wire [4-1:0] node10142;
	wire [4-1:0] node10143;
	wire [4-1:0] node10144;
	wire [4-1:0] node10148;
	wire [4-1:0] node10151;
	wire [4-1:0] node10152;
	wire [4-1:0] node10155;
	wire [4-1:0] node10158;
	wire [4-1:0] node10159;
	wire [4-1:0] node10160;
	wire [4-1:0] node10162;
	wire [4-1:0] node10164;
	wire [4-1:0] node10167;
	wire [4-1:0] node10170;
	wire [4-1:0] node10172;
	wire [4-1:0] node10173;
	wire [4-1:0] node10175;
	wire [4-1:0] node10179;
	wire [4-1:0] node10180;
	wire [4-1:0] node10181;
	wire [4-1:0] node10182;
	wire [4-1:0] node10183;
	wire [4-1:0] node10184;
	wire [4-1:0] node10188;
	wire [4-1:0] node10191;
	wire [4-1:0] node10194;
	wire [4-1:0] node10195;
	wire [4-1:0] node10196;
	wire [4-1:0] node10200;
	wire [4-1:0] node10201;
	wire [4-1:0] node10205;
	wire [4-1:0] node10207;
	wire [4-1:0] node10208;
	wire [4-1:0] node10210;
	wire [4-1:0] node10214;
	wire [4-1:0] node10215;
	wire [4-1:0] node10216;
	wire [4-1:0] node10217;
	wire [4-1:0] node10218;
	wire [4-1:0] node10219;
	wire [4-1:0] node10220;
	wire [4-1:0] node10221;
	wire [4-1:0] node10222;
	wire [4-1:0] node10225;
	wire [4-1:0] node10226;
	wire [4-1:0] node10230;
	wire [4-1:0] node10231;
	wire [4-1:0] node10233;
	wire [4-1:0] node10236;
	wire [4-1:0] node10239;
	wire [4-1:0] node10240;
	wire [4-1:0] node10243;
	wire [4-1:0] node10245;
	wire [4-1:0] node10248;
	wire [4-1:0] node10249;
	wire [4-1:0] node10250;
	wire [4-1:0] node10251;
	wire [4-1:0] node10253;
	wire [4-1:0] node10258;
	wire [4-1:0] node10259;
	wire [4-1:0] node10262;
	wire [4-1:0] node10265;
	wire [4-1:0] node10266;
	wire [4-1:0] node10267;
	wire [4-1:0] node10268;
	wire [4-1:0] node10269;
	wire [4-1:0] node10271;
	wire [4-1:0] node10275;
	wire [4-1:0] node10277;
	wire [4-1:0] node10279;
	wire [4-1:0] node10282;
	wire [4-1:0] node10283;
	wire [4-1:0] node10284;
	wire [4-1:0] node10287;
	wire [4-1:0] node10288;
	wire [4-1:0] node10292;
	wire [4-1:0] node10293;
	wire [4-1:0] node10295;
	wire [4-1:0] node10299;
	wire [4-1:0] node10300;
	wire [4-1:0] node10301;
	wire [4-1:0] node10303;
	wire [4-1:0] node10306;
	wire [4-1:0] node10307;
	wire [4-1:0] node10310;
	wire [4-1:0] node10313;
	wire [4-1:0] node10314;
	wire [4-1:0] node10316;
	wire [4-1:0] node10318;
	wire [4-1:0] node10321;
	wire [4-1:0] node10322;
	wire [4-1:0] node10325;
	wire [4-1:0] node10328;
	wire [4-1:0] node10329;
	wire [4-1:0] node10330;
	wire [4-1:0] node10331;
	wire [4-1:0] node10332;
	wire [4-1:0] node10335;
	wire [4-1:0] node10336;
	wire [4-1:0] node10340;
	wire [4-1:0] node10341;
	wire [4-1:0] node10343;
	wire [4-1:0] node10347;
	wire [4-1:0] node10348;
	wire [4-1:0] node10350;
	wire [4-1:0] node10353;
	wire [4-1:0] node10354;
	wire [4-1:0] node10356;
	wire [4-1:0] node10360;
	wire [4-1:0] node10361;
	wire [4-1:0] node10362;
	wire [4-1:0] node10363;
	wire [4-1:0] node10367;
	wire [4-1:0] node10368;
	wire [4-1:0] node10371;
	wire [4-1:0] node10372;
	wire [4-1:0] node10374;
	wire [4-1:0] node10378;
	wire [4-1:0] node10379;
	wire [4-1:0] node10380;
	wire [4-1:0] node10381;
	wire [4-1:0] node10386;
	wire [4-1:0] node10387;
	wire [4-1:0] node10388;
	wire [4-1:0] node10389;
	wire [4-1:0] node10392;
	wire [4-1:0] node10395;
	wire [4-1:0] node10396;
	wire [4-1:0] node10400;
	wire [4-1:0] node10402;
	wire [4-1:0] node10403;
	wire [4-1:0] node10407;
	wire [4-1:0] node10408;
	wire [4-1:0] node10409;
	wire [4-1:0] node10410;
	wire [4-1:0] node10411;
	wire [4-1:0] node10413;
	wire [4-1:0] node10414;
	wire [4-1:0] node10417;
	wire [4-1:0] node10419;
	wire [4-1:0] node10422;
	wire [4-1:0] node10423;
	wire [4-1:0] node10426;
	wire [4-1:0] node10429;
	wire [4-1:0] node10430;
	wire [4-1:0] node10431;
	wire [4-1:0] node10435;
	wire [4-1:0] node10436;
	wire [4-1:0] node10439;
	wire [4-1:0] node10440;
	wire [4-1:0] node10444;
	wire [4-1:0] node10445;
	wire [4-1:0] node10446;
	wire [4-1:0] node10447;
	wire [4-1:0] node10448;
	wire [4-1:0] node10451;
	wire [4-1:0] node10452;
	wire [4-1:0] node10456;
	wire [4-1:0] node10457;
	wire [4-1:0] node10462;
	wire [4-1:0] node10463;
	wire [4-1:0] node10465;
	wire [4-1:0] node10468;
	wire [4-1:0] node10469;
	wire [4-1:0] node10470;
	wire [4-1:0] node10472;
	wire [4-1:0] node10476;
	wire [4-1:0] node10478;
	wire [4-1:0] node10480;
	wire [4-1:0] node10483;
	wire [4-1:0] node10484;
	wire [4-1:0] node10485;
	wire [4-1:0] node10486;
	wire [4-1:0] node10487;
	wire [4-1:0] node10490;
	wire [4-1:0] node10492;
	wire [4-1:0] node10493;
	wire [4-1:0] node10497;
	wire [4-1:0] node10498;
	wire [4-1:0] node10499;
	wire [4-1:0] node10501;
	wire [4-1:0] node10504;
	wire [4-1:0] node10507;
	wire [4-1:0] node10508;
	wire [4-1:0] node10510;
	wire [4-1:0] node10513;
	wire [4-1:0] node10515;
	wire [4-1:0] node10518;
	wire [4-1:0] node10519;
	wire [4-1:0] node10520;
	wire [4-1:0] node10522;
	wire [4-1:0] node10523;
	wire [4-1:0] node10527;
	wire [4-1:0] node10530;
	wire [4-1:0] node10531;
	wire [4-1:0] node10533;
	wire [4-1:0] node10536;
	wire [4-1:0] node10537;
	wire [4-1:0] node10538;
	wire [4-1:0] node10542;
	wire [4-1:0] node10544;
	wire [4-1:0] node10547;
	wire [4-1:0] node10548;
	wire [4-1:0] node10549;
	wire [4-1:0] node10550;
	wire [4-1:0] node10554;
	wire [4-1:0] node10555;
	wire [4-1:0] node10556;
	wire [4-1:0] node10560;
	wire [4-1:0] node10563;
	wire [4-1:0] node10564;
	wire [4-1:0] node10565;
	wire [4-1:0] node10567;
	wire [4-1:0] node10569;
	wire [4-1:0] node10572;
	wire [4-1:0] node10574;
	wire [4-1:0] node10577;
	wire [4-1:0] node10578;
	wire [4-1:0] node10580;
	wire [4-1:0] node10583;
	wire [4-1:0] node10586;
	wire [4-1:0] node10587;
	wire [4-1:0] node10588;
	wire [4-1:0] node10589;
	wire [4-1:0] node10590;
	wire [4-1:0] node10591;
	wire [4-1:0] node10592;
	wire [4-1:0] node10595;
	wire [4-1:0] node10596;
	wire [4-1:0] node10599;
	wire [4-1:0] node10602;
	wire [4-1:0] node10603;
	wire [4-1:0] node10604;
	wire [4-1:0] node10607;
	wire [4-1:0] node10610;
	wire [4-1:0] node10612;
	wire [4-1:0] node10615;
	wire [4-1:0] node10616;
	wire [4-1:0] node10618;
	wire [4-1:0] node10619;
	wire [4-1:0] node10621;
	wire [4-1:0] node10624;
	wire [4-1:0] node10627;
	wire [4-1:0] node10629;
	wire [4-1:0] node10632;
	wire [4-1:0] node10633;
	wire [4-1:0] node10634;
	wire [4-1:0] node10635;
	wire [4-1:0] node10639;
	wire [4-1:0] node10640;
	wire [4-1:0] node10644;
	wire [4-1:0] node10645;
	wire [4-1:0] node10646;
	wire [4-1:0] node10650;
	wire [4-1:0] node10653;
	wire [4-1:0] node10654;
	wire [4-1:0] node10655;
	wire [4-1:0] node10656;
	wire [4-1:0] node10657;
	wire [4-1:0] node10658;
	wire [4-1:0] node10660;
	wire [4-1:0] node10664;
	wire [4-1:0] node10666;
	wire [4-1:0] node10669;
	wire [4-1:0] node10670;
	wire [4-1:0] node10673;
	wire [4-1:0] node10675;
	wire [4-1:0] node10676;
	wire [4-1:0] node10680;
	wire [4-1:0] node10681;
	wire [4-1:0] node10682;
	wire [4-1:0] node10684;
	wire [4-1:0] node10687;
	wire [4-1:0] node10690;
	wire [4-1:0] node10691;
	wire [4-1:0] node10692;
	wire [4-1:0] node10696;
	wire [4-1:0] node10699;
	wire [4-1:0] node10700;
	wire [4-1:0] node10701;
	wire [4-1:0] node10704;
	wire [4-1:0] node10706;
	wire [4-1:0] node10709;
	wire [4-1:0] node10710;
	wire [4-1:0] node10712;
	wire [4-1:0] node10715;
	wire [4-1:0] node10718;
	wire [4-1:0] node10719;
	wire [4-1:0] node10720;
	wire [4-1:0] node10721;
	wire [4-1:0] node10722;
	wire [4-1:0] node10723;
	wire [4-1:0] node10724;
	wire [4-1:0] node10725;
	wire [4-1:0] node10729;
	wire [4-1:0] node10730;
	wire [4-1:0] node10734;
	wire [4-1:0] node10736;
	wire [4-1:0] node10737;
	wire [4-1:0] node10741;
	wire [4-1:0] node10744;
	wire [4-1:0] node10745;
	wire [4-1:0] node10746;
	wire [4-1:0] node10748;
	wire [4-1:0] node10749;
	wire [4-1:0] node10752;
	wire [4-1:0] node10755;
	wire [4-1:0] node10757;
	wire [4-1:0] node10760;
	wire [4-1:0] node10761;
	wire [4-1:0] node10762;
	wire [4-1:0] node10765;
	wire [4-1:0] node10767;
	wire [4-1:0] node10771;
	wire [4-1:0] node10772;
	wire [4-1:0] node10773;
	wire [4-1:0] node10776;
	wire [4-1:0] node10777;
	wire [4-1:0] node10780;
	wire [4-1:0] node10783;
	wire [4-1:0] node10784;
	wire [4-1:0] node10787;
	wire [4-1:0] node10788;
	wire [4-1:0] node10792;
	wire [4-1:0] node10793;
	wire [4-1:0] node10794;
	wire [4-1:0] node10795;
	wire [4-1:0] node10796;
	wire [4-1:0] node10798;
	wire [4-1:0] node10799;
	wire [4-1:0] node10802;
	wire [4-1:0] node10805;
	wire [4-1:0] node10806;
	wire [4-1:0] node10807;
	wire [4-1:0] node10811;
	wire [4-1:0] node10812;
	wire [4-1:0] node10816;
	wire [4-1:0] node10817;
	wire [4-1:0] node10818;
	wire [4-1:0] node10819;
	wire [4-1:0] node10824;
	wire [4-1:0] node10827;
	wire [4-1:0] node10828;
	wire [4-1:0] node10829;
	wire [4-1:0] node10831;
	wire [4-1:0] node10834;
	wire [4-1:0] node10835;
	wire [4-1:0] node10836;
	wire [4-1:0] node10841;
	wire [4-1:0] node10843;
	wire [4-1:0] node10844;
	wire [4-1:0] node10846;
	wire [4-1:0] node10849;
	wire [4-1:0] node10852;
	wire [4-1:0] node10853;
	wire [4-1:0] node10854;
	wire [4-1:0] node10856;
	wire [4-1:0] node10858;
	wire [4-1:0] node10861;
	wire [4-1:0] node10862;
	wire [4-1:0] node10863;
	wire [4-1:0] node10867;
	wire [4-1:0] node10870;
	wire [4-1:0] node10871;
	wire [4-1:0] node10872;
	wire [4-1:0] node10874;
	wire [4-1:0] node10876;
	wire [4-1:0] node10879;
	wire [4-1:0] node10881;

	assign outp = (inp[14]) ? node5708 : node1;
		assign node1 = (inp[7]) ? node2823 : node2;
			assign node2 = (inp[5]) ? node1408 : node3;
				assign node3 = (inp[0]) ? node737 : node4;
					assign node4 = (inp[15]) ? node388 : node5;
						assign node5 = (inp[3]) ? node205 : node6;
							assign node6 = (inp[2]) ? node110 : node7;
								assign node7 = (inp[8]) ? node67 : node8;
									assign node8 = (inp[1]) ? node36 : node9;
										assign node9 = (inp[9]) ? node23 : node10;
											assign node10 = (inp[6]) ? node18 : node11;
												assign node11 = (inp[10]) ? node13 : 4'b1111;
													assign node13 = (inp[4]) ? node15 : 4'b0011;
														assign node15 = (inp[12]) ? 4'b0111 : 4'b0011;
												assign node18 = (inp[11]) ? 4'b1111 : node19;
													assign node19 = (inp[12]) ? 4'b0011 : 4'b0111;
											assign node23 = (inp[6]) ? node31 : node24;
												assign node24 = (inp[11]) ? 4'b0111 : node25;
													assign node25 = (inp[4]) ? 4'b1111 : node26;
														assign node26 = (inp[12]) ? 4'b1111 : 4'b1011;
												assign node31 = (inp[11]) ? node33 : 4'b0111;
													assign node33 = (inp[12]) ? 4'b1011 : 4'b1111;
										assign node36 = (inp[10]) ? node56 : node37;
											assign node37 = (inp[6]) ? node43 : node38;
												assign node38 = (inp[9]) ? node40 : 4'b0011;
													assign node40 = (inp[4]) ? 4'b0111 : 4'b0011;
												assign node43 = (inp[12]) ? node49 : node44;
													assign node44 = (inp[13]) ? node46 : 4'b0011;
														assign node46 = (inp[11]) ? 4'b0111 : 4'b1111;
													assign node49 = (inp[4]) ? node53 : node50;
														assign node50 = (inp[11]) ? 4'b1011 : 4'b1111;
														assign node53 = (inp[9]) ? 4'b1011 : 4'b0011;
											assign node56 = (inp[9]) ? node62 : node57;
												assign node57 = (inp[13]) ? node59 : 4'b1011;
													assign node59 = (inp[11]) ? 4'b1011 : 4'b0111;
												assign node62 = (inp[6]) ? node64 : 4'b1011;
													assign node64 = (inp[13]) ? 4'b1011 : 4'b0011;
									assign node67 = (inp[9]) ? node91 : node68;
										assign node68 = (inp[4]) ? node78 : node69;
											assign node69 = (inp[11]) ? node71 : 4'b1110;
												assign node71 = (inp[1]) ? 4'b1010 : node72;
													assign node72 = (inp[12]) ? 4'b1010 : node73;
														assign node73 = (inp[10]) ? 4'b1010 : 4'b1110;
											assign node78 = (inp[10]) ? node86 : node79;
												assign node79 = (inp[6]) ? node81 : 4'b1010;
													assign node81 = (inp[11]) ? node83 : 4'b0010;
														assign node83 = (inp[13]) ? 4'b0010 : 4'b1010;
												assign node86 = (inp[12]) ? node88 : 4'b1010;
													assign node88 = (inp[6]) ? 4'b1110 : 4'b0110;
										assign node91 = (inp[11]) ? node99 : node92;
											assign node92 = (inp[4]) ? node94 : 4'b1110;
												assign node94 = (inp[12]) ? 4'b0110 : node95;
													assign node95 = (inp[13]) ? 4'b1110 : 4'b0110;
											assign node99 = (inp[6]) ? node107 : node100;
												assign node100 = (inp[1]) ? node104 : node101;
													assign node101 = (inp[13]) ? 4'b0010 : 4'b0110;
													assign node104 = (inp[10]) ? 4'b0010 : 4'b1010;
												assign node107 = (inp[12]) ? 4'b1010 : 4'b1110;
								assign node110 = (inp[8]) ? node152 : node111;
									assign node111 = (inp[13]) ? node131 : node112;
										assign node112 = (inp[12]) ? node120 : node113;
											assign node113 = (inp[11]) ? node115 : 4'b0110;
												assign node115 = (inp[4]) ? node117 : 4'b0010;
													assign node117 = (inp[9]) ? 4'b0110 : 4'b0010;
											assign node120 = (inp[10]) ? node126 : node121;
												assign node121 = (inp[11]) ? 4'b1110 : node122;
													assign node122 = (inp[1]) ? 4'b0010 : 4'b1010;
												assign node126 = (inp[11]) ? 4'b0010 : node127;
													assign node127 = (inp[6]) ? 4'b0010 : 4'b1010;
										assign node131 = (inp[11]) ? node141 : node132;
											assign node132 = (inp[10]) ? node136 : node133;
												assign node133 = (inp[1]) ? 4'b1010 : 4'b0110;
												assign node136 = (inp[1]) ? node138 : 4'b1110;
													assign node138 = (inp[6]) ? 4'b1110 : 4'b0110;
											assign node141 = (inp[10]) ? 4'b0010 : node142;
												assign node142 = (inp[6]) ? node146 : node143;
													assign node143 = (inp[1]) ? 4'b1110 : 4'b0110;
													assign node146 = (inp[9]) ? node148 : 4'b0110;
														assign node148 = (inp[12]) ? 4'b0010 : 4'b0110;
									assign node152 = (inp[9]) ? node182 : node153;
										assign node153 = (inp[12]) ? node167 : node154;
											assign node154 = (inp[4]) ? node158 : node155;
												assign node155 = (inp[11]) ? 4'b1011 : 4'b0111;
												assign node158 = (inp[6]) ? node164 : node159;
													assign node159 = (inp[1]) ? 4'b0011 : node160;
														assign node160 = (inp[13]) ? 4'b0011 : 4'b1011;
													assign node164 = (inp[10]) ? 4'b0111 : 4'b0011;
											assign node167 = (inp[4]) ? 4'b1111 : node168;
												assign node168 = (inp[13]) ? node176 : node169;
													assign node169 = (inp[1]) ? node173 : node170;
														assign node170 = (inp[11]) ? 4'b0111 : 4'b1111;
														assign node173 = (inp[10]) ? 4'b0011 : 4'b1011;
													assign node176 = (inp[6]) ? node178 : 4'b1011;
														assign node178 = (inp[11]) ? 4'b0011 : 4'b1011;
										assign node182 = (inp[12]) ? node186 : node183;
											assign node183 = (inp[4]) ? 4'b0111 : 4'b0011;
											assign node186 = (inp[6]) ? node196 : node187;
												assign node187 = (inp[10]) ? node193 : node188;
													assign node188 = (inp[1]) ? 4'b1111 : node189;
														assign node189 = (inp[4]) ? 4'b1111 : 4'b0011;
													assign node193 = (inp[4]) ? 4'b0011 : 4'b0111;
												assign node196 = (inp[13]) ? node202 : node197;
													assign node197 = (inp[1]) ? node199 : 4'b0011;
														assign node199 = (inp[11]) ? 4'b0011 : 4'b1011;
													assign node202 = (inp[4]) ? 4'b0011 : 4'b0111;
							assign node205 = (inp[9]) ? node301 : node206;
								assign node206 = (inp[4]) ? node250 : node207;
									assign node207 = (inp[11]) ? node233 : node208;
										assign node208 = (inp[10]) ? node222 : node209;
											assign node209 = (inp[6]) ? 4'b0111 : node210;
												assign node210 = (inp[1]) ? node214 : node211;
													assign node211 = (inp[13]) ? 4'b1110 : 4'b1111;
													assign node214 = (inp[13]) ? node218 : node215;
														assign node215 = (inp[12]) ? 4'b0111 : 4'b1110;
														assign node218 = (inp[8]) ? 4'b0110 : 4'b0111;
											assign node222 = (inp[13]) ? node230 : node223;
												assign node223 = (inp[12]) ? node227 : node224;
													assign node224 = (inp[6]) ? 4'b0110 : 4'b0111;
													assign node227 = (inp[2]) ? 4'b1010 : 4'b0011;
												assign node230 = (inp[8]) ? 4'b1011 : 4'b1010;
										assign node233 = (inp[6]) ? node239 : node234;
											assign node234 = (inp[1]) ? 4'b1010 : node235;
												assign node235 = (inp[8]) ? 4'b0110 : 4'b0111;
											assign node239 = (inp[8]) ? node243 : node240;
												assign node240 = (inp[2]) ? 4'b1010 : 4'b1011;
												assign node243 = (inp[1]) ? 4'b0010 : node244;
													assign node244 = (inp[10]) ? 4'b1010 : node245;
														assign node245 = (inp[13]) ? 4'b1110 : 4'b1010;
									assign node250 = (inp[6]) ? node274 : node251;
										assign node251 = (inp[11]) ? node261 : node252;
											assign node252 = (inp[8]) ? node256 : node253;
												assign node253 = (inp[2]) ? 4'b1010 : 4'b1011;
												assign node256 = (inp[2]) ? 4'b0011 : node257;
													assign node257 = (inp[12]) ? 4'b1010 : 4'b0010;
											assign node261 = (inp[10]) ? node271 : node262;
												assign node262 = (inp[1]) ? node268 : node263;
													assign node263 = (inp[13]) ? 4'b0010 : node264;
														assign node264 = (inp[8]) ? 4'b0011 : 4'b0010;
													assign node268 = (inp[13]) ? 4'b1100 : 4'b0010;
												assign node271 = (inp[2]) ? 4'b1101 : 4'b0011;
										assign node274 = (inp[11]) ? node290 : node275;
											assign node275 = (inp[13]) ? node281 : node276;
												assign node276 = (inp[2]) ? node278 : 4'b0010;
													assign node278 = (inp[8]) ? 4'b0011 : 4'b0010;
												assign node281 = (inp[12]) ? node285 : node282;
													assign node282 = (inp[1]) ? 4'b1010 : 4'b0010;
													assign node285 = (inp[8]) ? 4'b1101 : node286;
														assign node286 = (inp[2]) ? 4'b0010 : 4'b0101;
											assign node290 = (inp[2]) ? node296 : node291;
												assign node291 = (inp[8]) ? 4'b1100 : node292;
													assign node292 = (inp[13]) ? 4'b0101 : 4'b1101;
												assign node296 = (inp[8]) ? 4'b0101 : node297;
													assign node297 = (inp[13]) ? 4'b0010 : 4'b1010;
								assign node301 = (inp[4]) ? node353 : node302;
									assign node302 = (inp[12]) ? node334 : node303;
										assign node303 = (inp[10]) ? node317 : node304;
											assign node304 = (inp[13]) ? node310 : node305;
												assign node305 = (inp[1]) ? node307 : 4'b0011;
													assign node307 = (inp[2]) ? 4'b1010 : 4'b1011;
												assign node310 = (inp[6]) ? 4'b0010 : node311;
													assign node311 = (inp[11]) ? 4'b1010 : node312;
														assign node312 = (inp[1]) ? 4'b0010 : 4'b1010;
											assign node317 = (inp[13]) ? node329 : node318;
												assign node318 = (inp[1]) ? node326 : node319;
													assign node319 = (inp[8]) ? node323 : node320;
														assign node320 = (inp[6]) ? 4'b0000 : 4'b0010;
														assign node323 = (inp[2]) ? 4'b0011 : 4'b0010;
													assign node326 = (inp[6]) ? 4'b1101 : 4'b1011;
												assign node329 = (inp[8]) ? 4'b1101 : node330;
													assign node330 = (inp[11]) ? 4'b1100 : 4'b0010;
										assign node334 = (inp[11]) ? node342 : node335;
											assign node335 = (inp[10]) ? node337 : 4'b0011;
												assign node337 = (inp[6]) ? node339 : 4'b1100;
													assign node339 = (inp[1]) ? 4'b1101 : 4'b0101;
											assign node342 = (inp[10]) ? node348 : node343;
												assign node343 = (inp[6]) ? 4'b1100 : node344;
													assign node344 = (inp[8]) ? 4'b1100 : 4'b0010;
												assign node348 = (inp[1]) ? 4'b1100 : node349;
													assign node349 = (inp[6]) ? 4'b0101 : 4'b1101;
									assign node353 = (inp[12]) ? node369 : node354;
										assign node354 = (inp[10]) ? node364 : node355;
											assign node355 = (inp[11]) ? node357 : 4'b0100;
												assign node357 = (inp[8]) ? 4'b1101 : node358;
													assign node358 = (inp[2]) ? node360 : 4'b1101;
														assign node360 = (inp[6]) ? 4'b1100 : 4'b0100;
											assign node364 = (inp[1]) ? 4'b1000 : node365;
												assign node365 = (inp[2]) ? 4'b0100 : 4'b1100;
										assign node369 = (inp[2]) ? node379 : node370;
											assign node370 = (inp[8]) ? node374 : node371;
												assign node371 = (inp[10]) ? 4'b0001 : 4'b0101;
												assign node374 = (inp[11]) ? 4'b0000 : node375;
													assign node375 = (inp[1]) ? 4'b0100 : 4'b1100;
											assign node379 = (inp[8]) ? node383 : node380;
												assign node380 = (inp[13]) ? 4'b0000 : 4'b1000;
												assign node383 = (inp[11]) ? node385 : 4'b1001;
													assign node385 = (inp[1]) ? 4'b0001 : 4'b1001;
						assign node388 = (inp[3]) ? node540 : node389;
							assign node389 = (inp[2]) ? node463 : node390;
								assign node390 = (inp[8]) ? node428 : node391;
									assign node391 = (inp[12]) ? node411 : node392;
										assign node392 = (inp[6]) ? node400 : node393;
											assign node393 = (inp[1]) ? node395 : 4'b0001;
												assign node395 = (inp[10]) ? node397 : 4'b0101;
													assign node397 = (inp[13]) ? 4'b0101 : 4'b1101;
											assign node400 = (inp[10]) ? node408 : node401;
												assign node401 = (inp[1]) ? node403 : 4'b1101;
													assign node403 = (inp[11]) ? 4'b1001 : node404;
														assign node404 = (inp[4]) ? 4'b0101 : 4'b1001;
												assign node408 = (inp[9]) ? 4'b0101 : 4'b0001;
										assign node411 = (inp[13]) ? node421 : node412;
											assign node412 = (inp[4]) ? 4'b1001 : node413;
												assign node413 = (inp[10]) ? node417 : node414;
													assign node414 = (inp[11]) ? 4'b0101 : 4'b0001;
													assign node417 = (inp[11]) ? 4'b0001 : 4'b0101;
											assign node421 = (inp[6]) ? 4'b0101 : node422;
												assign node422 = (inp[10]) ? node424 : 4'b1101;
													assign node424 = (inp[11]) ? 4'b0001 : 4'b1001;
									assign node428 = (inp[13]) ? node446 : node429;
										assign node429 = (inp[9]) ? node437 : node430;
											assign node430 = (inp[11]) ? 4'b1100 : node431;
												assign node431 = (inp[4]) ? 4'b0000 : node432;
													assign node432 = (inp[12]) ? 4'b1100 : 4'b0100;
											assign node437 = (inp[4]) ? node443 : node438;
												assign node438 = (inp[1]) ? node440 : 4'b0000;
													assign node440 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node443 = (inp[1]) ? 4'b1100 : 4'b1000;
										assign node446 = (inp[1]) ? node448 : 4'b1100;
											assign node448 = (inp[10]) ? node454 : node449;
												assign node449 = (inp[6]) ? node451 : 4'b0100;
													assign node451 = (inp[11]) ? 4'b0100 : 4'b1100;
												assign node454 = (inp[9]) ? node458 : node455;
													assign node455 = (inp[4]) ? 4'b0100 : 4'b0000;
													assign node458 = (inp[6]) ? 4'b0100 : node459;
														assign node459 = (inp[4]) ? 4'b0100 : 4'b1100;
								assign node463 = (inp[8]) ? node497 : node464;
									assign node464 = (inp[9]) ? node482 : node465;
										assign node465 = (inp[10]) ? node469 : node466;
											assign node466 = (inp[4]) ? 4'b0000 : 4'b0100;
											assign node469 = (inp[13]) ? node477 : node470;
												assign node470 = (inp[12]) ? node474 : node471;
													assign node471 = (inp[4]) ? 4'b1000 : 4'b0100;
													assign node474 = (inp[4]) ? 4'b0100 : 4'b1000;
												assign node477 = (inp[1]) ? 4'b1100 : node478;
													assign node478 = (inp[11]) ? 4'b1000 : 4'b0000;
										assign node482 = (inp[13]) ? node490 : node483;
											assign node483 = (inp[1]) ? 4'b0000 : node484;
												assign node484 = (inp[6]) ? node486 : 4'b1000;
													assign node486 = (inp[11]) ? 4'b1000 : 4'b0000;
											assign node490 = (inp[11]) ? node492 : 4'b1100;
												assign node492 = (inp[10]) ? node494 : 4'b1000;
													assign node494 = (inp[4]) ? 4'b0000 : 4'b0100;
									assign node497 = (inp[12]) ? node527 : node498;
										assign node498 = (inp[13]) ? node510 : node499;
											assign node499 = (inp[4]) ? node507 : node500;
												assign node500 = (inp[9]) ? node502 : 4'b1001;
													assign node502 = (inp[1]) ? node504 : 4'b0001;
														assign node504 = (inp[6]) ? 4'b1001 : 4'b0001;
												assign node507 = (inp[9]) ? 4'b1101 : 4'b1001;
											assign node510 = (inp[9]) ? node518 : node511;
												assign node511 = (inp[1]) ? node513 : 4'b1001;
													assign node513 = (inp[4]) ? 4'b0101 : node514;
														assign node514 = (inp[10]) ? 4'b0001 : 4'b0101;
												assign node518 = (inp[10]) ? node524 : node519;
													assign node519 = (inp[4]) ? node521 : 4'b1001;
														assign node521 = (inp[6]) ? 4'b1101 : 4'b0101;
													assign node524 = (inp[4]) ? 4'b1001 : 4'b1101;
										assign node527 = (inp[13]) ? node533 : node528;
											assign node528 = (inp[9]) ? 4'b0101 : node529;
												assign node529 = (inp[1]) ? 4'b0101 : 4'b1101;
											assign node533 = (inp[10]) ? 4'b0101 : node534;
												assign node534 = (inp[1]) ? 4'b0001 : node535;
													assign node535 = (inp[9]) ? 4'b0001 : 4'b1001;
							assign node540 = (inp[9]) ? node638 : node541;
								assign node541 = (inp[4]) ? node597 : node542;
									assign node542 = (inp[10]) ? node568 : node543;
										assign node543 = (inp[11]) ? node555 : node544;
											assign node544 = (inp[1]) ? node552 : node545;
												assign node545 = (inp[8]) ? node549 : node546;
													assign node546 = (inp[2]) ? 4'b1100 : 4'b1101;
													assign node549 = (inp[13]) ? 4'b0101 : 4'b1101;
												assign node552 = (inp[12]) ? 4'b0100 : 4'b1100;
											assign node555 = (inp[12]) ? node561 : node556;
												assign node556 = (inp[2]) ? node558 : 4'b0100;
													assign node558 = (inp[8]) ? 4'b0101 : 4'b0100;
												assign node561 = (inp[8]) ? node565 : node562;
													assign node562 = (inp[13]) ? 4'b0101 : 4'b0100;
													assign node565 = (inp[2]) ? 4'b0001 : 4'b1000;
										assign node568 = (inp[12]) ? node582 : node569;
											assign node569 = (inp[2]) ? node575 : node570;
												assign node570 = (inp[8]) ? node572 : 4'b0101;
													assign node572 = (inp[11]) ? 4'b0100 : 4'b1100;
												assign node575 = (inp[8]) ? node577 : 4'b0000;
													assign node577 = (inp[11]) ? node579 : 4'b1001;
														assign node579 = (inp[6]) ? 4'b0001 : 4'b1001;
											assign node582 = (inp[13]) ? node592 : node583;
												assign node583 = (inp[1]) ? node589 : node584;
													assign node584 = (inp[8]) ? node586 : 4'b1000;
														assign node586 = (inp[6]) ? 4'b0001 : 4'b1001;
													assign node589 = (inp[6]) ? 4'b1001 : 4'b0001;
												assign node592 = (inp[8]) ? 4'b1000 : node593;
													assign node593 = (inp[11]) ? 4'b0001 : 4'b1000;
									assign node597 = (inp[10]) ? node627 : node598;
										assign node598 = (inp[12]) ? node608 : node599;
											assign node599 = (inp[2]) ? node605 : node600;
												assign node600 = (inp[1]) ? 4'b0000 : node601;
													assign node601 = (inp[13]) ? 4'b0000 : 4'b1000;
												assign node605 = (inp[8]) ? 4'b1001 : 4'b0000;
											assign node608 = (inp[6]) ? node618 : node609;
												assign node609 = (inp[11]) ? node613 : node610;
													assign node610 = (inp[13]) ? 4'b1000 : 4'b1001;
													assign node613 = (inp[8]) ? 4'b0000 : node614;
														assign node614 = (inp[2]) ? 4'b0000 : 4'b0001;
												assign node618 = (inp[11]) ? node622 : node619;
													assign node619 = (inp[8]) ? 4'b0000 : 4'b0001;
													assign node622 = (inp[1]) ? 4'b0111 : node623;
														assign node623 = (inp[8]) ? 4'b1110 : 4'b1111;
										assign node627 = (inp[12]) ? node633 : node628;
											assign node628 = (inp[11]) ? 4'b1110 : node629;
												assign node629 = (inp[13]) ? 4'b0001 : 4'b0000;
											assign node633 = (inp[1]) ? node635 : 4'b1110;
												assign node635 = (inp[6]) ? 4'b1111 : 4'b0111;
								assign node638 = (inp[4]) ? node682 : node639;
									assign node639 = (inp[12]) ? node663 : node640;
										assign node640 = (inp[10]) ? node652 : node641;
											assign node641 = (inp[13]) ? node647 : node642;
												assign node642 = (inp[11]) ? node644 : 4'b1000;
													assign node644 = (inp[1]) ? 4'b1000 : 4'b0000;
												assign node647 = (inp[8]) ? 4'b1000 : node648;
													assign node648 = (inp[2]) ? 4'b0000 : 4'b0001;
											assign node652 = (inp[8]) ? node660 : node653;
												assign node653 = (inp[11]) ? 4'b1110 : node654;
													assign node654 = (inp[2]) ? node656 : 4'b1001;
														assign node656 = (inp[6]) ? 4'b0000 : 4'b0000;
												assign node660 = (inp[11]) ? 4'b0111 : 4'b1111;
										assign node663 = (inp[2]) ? node677 : node664;
											assign node664 = (inp[1]) ? node672 : node665;
												assign node665 = (inp[10]) ? 4'b0111 : node666;
													assign node666 = (inp[6]) ? 4'b0001 : node667;
														assign node667 = (inp[11]) ? 4'b0001 : 4'b1001;
												assign node672 = (inp[6]) ? node674 : 4'b1000;
													assign node674 = (inp[13]) ? 4'b1111 : 4'b1110;
											assign node677 = (inp[8]) ? node679 : 4'b1110;
												assign node679 = (inp[1]) ? 4'b1111 : 4'b0111;
									assign node682 = (inp[12]) ? node716 : node683;
										assign node683 = (inp[10]) ? node701 : node684;
											assign node684 = (inp[11]) ? node694 : node685;
												assign node685 = (inp[8]) ? node691 : node686;
													assign node686 = (inp[1]) ? 4'b0111 : node687;
														assign node687 = (inp[6]) ? 4'b0110 : 4'b1110;
													assign node691 = (inp[6]) ? 4'b1111 : 4'b0111;
												assign node694 = (inp[1]) ? node696 : 4'b0111;
													assign node696 = (inp[2]) ? 4'b0111 : node697;
														assign node697 = (inp[13]) ? 4'b1111 : 4'b0111;
											assign node701 = (inp[6]) ? node705 : node702;
												assign node702 = (inp[1]) ? 4'b0111 : 4'b0110;
												assign node705 = (inp[11]) ? node709 : node706;
													assign node706 = (inp[1]) ? 4'b1011 : 4'b0111;
													assign node709 = (inp[13]) ? node713 : node710;
														assign node710 = (inp[2]) ? 4'b1010 : 4'b1011;
														assign node713 = (inp[1]) ? 4'b0010 : 4'b1010;
										assign node716 = (inp[8]) ? node720 : node717;
											assign node717 = (inp[2]) ? 4'b0010 : 4'b0011;
											assign node720 = (inp[2]) ? node734 : node721;
												assign node721 = (inp[13]) ? node727 : node722;
													assign node722 = (inp[10]) ? 4'b1010 : node723;
														assign node723 = (inp[11]) ? 4'b1010 : 4'b0110;
													assign node727 = (inp[1]) ? node731 : node728;
														assign node728 = (inp[10]) ? 4'b0010 : 4'b0110;
														assign node731 = (inp[6]) ? 4'b0010 : 4'b1010;
												assign node734 = (inp[1]) ? 4'b0011 : 4'b1011;
					assign node737 = (inp[15]) ? node1063 : node738;
						assign node738 = (inp[3]) ? node916 : node739;
							assign node739 = (inp[11]) ? node833 : node740;
								assign node740 = (inp[13]) ? node774 : node741;
									assign node741 = (inp[6]) ? node763 : node742;
										assign node742 = (inp[1]) ? node754 : node743;
											assign node743 = (inp[8]) ? node747 : node744;
												assign node744 = (inp[10]) ? 4'b1101 : 4'b1100;
												assign node747 = (inp[9]) ? node749 : 4'b1000;
													assign node749 = (inp[12]) ? 4'b1100 : node750;
														assign node750 = (inp[4]) ? 4'b1100 : 4'b1000;
											assign node754 = (inp[8]) ? node758 : node755;
												assign node755 = (inp[4]) ? 4'b1101 : 4'b1100;
												assign node758 = (inp[2]) ? node760 : 4'b1100;
													assign node760 = (inp[4]) ? 4'b0001 : 4'b0101;
										assign node763 = (inp[8]) ? node771 : node764;
											assign node764 = (inp[2]) ? node766 : 4'b0001;
												assign node766 = (inp[12]) ? node768 : 4'b0100;
													assign node768 = (inp[9]) ? 4'b0100 : 4'b0000;
											assign node771 = (inp[2]) ? 4'b1101 : 4'b0100;
									assign node774 = (inp[4]) ? node800 : node775;
										assign node775 = (inp[9]) ? node787 : node776;
											assign node776 = (inp[12]) ? node778 : 4'b0101;
												assign node778 = (inp[10]) ? 4'b0001 : node779;
													assign node779 = (inp[6]) ? node783 : node780;
														assign node780 = (inp[1]) ? 4'b0100 : 4'b1100;
														assign node783 = (inp[2]) ? 4'b0100 : 4'b0101;
											assign node787 = (inp[10]) ? node793 : node788;
												assign node788 = (inp[8]) ? node790 : 4'b1001;
													assign node790 = (inp[12]) ? 4'b0001 : 4'b0000;
												assign node793 = (inp[8]) ? node795 : 4'b0100;
													assign node795 = (inp[6]) ? 4'b1101 : node796;
														assign node796 = (inp[12]) ? 4'b0101 : 4'b0001;
										assign node800 = (inp[12]) ? node816 : node801;
											assign node801 = (inp[9]) ? node809 : node802;
												assign node802 = (inp[2]) ? node804 : 4'b0001;
													assign node804 = (inp[10]) ? 4'b0001 : node805;
														assign node805 = (inp[6]) ? 4'b0000 : 4'b1000;
												assign node809 = (inp[2]) ? 4'b1000 : node810;
													assign node810 = (inp[1]) ? 4'b1100 : node811;
														assign node811 = (inp[6]) ? 4'b0100 : 4'b1100;
											assign node816 = (inp[9]) ? node822 : node817;
												assign node817 = (inp[8]) ? 4'b1101 : node818;
													assign node818 = (inp[6]) ? 4'b0100 : 4'b1100;
												assign node822 = (inp[6]) ? node828 : node823;
													assign node823 = (inp[10]) ? 4'b0001 : node824;
														assign node824 = (inp[8]) ? 4'b0100 : 4'b1101;
													assign node828 = (inp[8]) ? node830 : 4'b0100;
														assign node830 = (inp[2]) ? 4'b1001 : 4'b1000;
								assign node833 = (inp[6]) ? node881 : node834;
									assign node834 = (inp[2]) ? node858 : node835;
										assign node835 = (inp[8]) ? node845 : node836;
											assign node836 = (inp[12]) ? 4'b0101 : node837;
												assign node837 = (inp[4]) ? 4'b0001 : node838;
													assign node838 = (inp[9]) ? 4'b0001 : node839;
														assign node839 = (inp[1]) ? 4'b0001 : 4'b0101;
											assign node845 = (inp[12]) ? node853 : node846;
												assign node846 = (inp[10]) ? node850 : node847;
													assign node847 = (inp[9]) ? 4'b0000 : 4'b0100;
													assign node850 = (inp[1]) ? 4'b1100 : 4'b0100;
												assign node853 = (inp[13]) ? node855 : 4'b0000;
													assign node855 = (inp[1]) ? 4'b1000 : 4'b0000;
										assign node858 = (inp[8]) ? node872 : node859;
											assign node859 = (inp[13]) ? node865 : node860;
												assign node860 = (inp[4]) ? 4'b0100 : node861;
													assign node861 = (inp[9]) ? 4'b0000 : 4'b0100;
												assign node865 = (inp[1]) ? node867 : 4'b0100;
													assign node867 = (inp[4]) ? node869 : 4'b1000;
														assign node869 = (inp[12]) ? 4'b1100 : 4'b1000;
											assign node872 = (inp[9]) ? node874 : 4'b1101;
												assign node874 = (inp[10]) ? 4'b0001 : node875;
													assign node875 = (inp[12]) ? node877 : 4'b1001;
														assign node877 = (inp[1]) ? 4'b1101 : 4'b1001;
									assign node881 = (inp[1]) ? node899 : node882;
										assign node882 = (inp[9]) ? node890 : node883;
											assign node883 = (inp[12]) ? node885 : 4'b1000;
												assign node885 = (inp[8]) ? 4'b1001 : node886;
													assign node886 = (inp[4]) ? 4'b1100 : 4'b1000;
											assign node890 = (inp[2]) ? 4'b1100 : node891;
												assign node891 = (inp[8]) ? node895 : node892;
													assign node892 = (inp[10]) ? 4'b1101 : 4'b1001;
													assign node895 = (inp[13]) ? 4'b1100 : 4'b1000;
										assign node899 = (inp[13]) ? node907 : node900;
											assign node900 = (inp[4]) ? 4'b0101 : node901;
												assign node901 = (inp[9]) ? 4'b1101 : node902;
													assign node902 = (inp[10]) ? 4'b1000 : 4'b1100;
											assign node907 = (inp[9]) ? 4'b0001 : node908;
												assign node908 = (inp[4]) ? 4'b0100 : node909;
													assign node909 = (inp[10]) ? 4'b0000 : node910;
														assign node910 = (inp[2]) ? 4'b0000 : 4'b0101;
							assign node916 = (inp[4]) ? node996 : node917;
								assign node917 = (inp[9]) ? node951 : node918;
									assign node918 = (inp[12]) ? node938 : node919;
										assign node919 = (inp[2]) ? node929 : node920;
											assign node920 = (inp[8]) ? node926 : node921;
												assign node921 = (inp[6]) ? node923 : 4'b0101;
													assign node923 = (inp[11]) ? 4'b1001 : 4'b0101;
												assign node926 = (inp[10]) ? 4'b0000 : 4'b0100;
											assign node929 = (inp[8]) ? node935 : node930;
												assign node930 = (inp[10]) ? node932 : 4'b1100;
													assign node932 = (inp[1]) ? 4'b0100 : 4'b1100;
												assign node935 = (inp[6]) ? 4'b0101 : 4'b1101;
										assign node938 = (inp[10]) ? node944 : node939;
											assign node939 = (inp[1]) ? 4'b1000 : node940;
												assign node940 = (inp[8]) ? 4'b1001 : 4'b0101;
											assign node944 = (inp[11]) ? 4'b0001 : node945;
												assign node945 = (inp[1]) ? 4'b0000 : node946;
													assign node946 = (inp[13]) ? 4'b0001 : 4'b0000;
									assign node951 = (inp[10]) ? node969 : node952;
										assign node952 = (inp[11]) ? node960 : node953;
											assign node953 = (inp[12]) ? node957 : node954;
												assign node954 = (inp[2]) ? 4'b0001 : 4'b1001;
												assign node957 = (inp[1]) ? 4'b0001 : 4'b0000;
											assign node960 = (inp[6]) ? node962 : 4'b0000;
												assign node962 = (inp[12]) ? 4'b1110 : node963;
													assign node963 = (inp[1]) ? node965 : 4'b1000;
														assign node965 = (inp[13]) ? 4'b0000 : 4'b0001;
										assign node969 = (inp[12]) ? node983 : node970;
											assign node970 = (inp[2]) ? node976 : node971;
												assign node971 = (inp[6]) ? node973 : 4'b0001;
													assign node973 = (inp[8]) ? 4'b1110 : 4'b1111;
												assign node976 = (inp[8]) ? 4'b0001 : node977;
													assign node977 = (inp[11]) ? node979 : 4'b0000;
														assign node979 = (inp[1]) ? 4'b0110 : 4'b0000;
											assign node983 = (inp[8]) ? node991 : node984;
												assign node984 = (inp[2]) ? node986 : 4'b0111;
													assign node986 = (inp[11]) ? 4'b0110 : node987;
														assign node987 = (inp[1]) ? 4'b1110 : 4'b0110;
												assign node991 = (inp[2]) ? node993 : 4'b1110;
													assign node993 = (inp[1]) ? 4'b0111 : 4'b1111;
								assign node996 = (inp[2]) ? node1024 : node997;
									assign node997 = (inp[8]) ? node1009 : node998;
										assign node998 = (inp[13]) ? node1004 : node999;
											assign node999 = (inp[12]) ? node1001 : 4'b1001;
												assign node1001 = (inp[10]) ? 4'b1111 : 4'b1011;
											assign node1004 = (inp[10]) ? node1006 : 4'b1111;
												assign node1006 = (inp[12]) ? 4'b1011 : 4'b1111;
										assign node1009 = (inp[9]) ? node1015 : node1010;
											assign node1010 = (inp[10]) ? node1012 : 4'b0000;
												assign node1012 = (inp[6]) ? 4'b0000 : 4'b1000;
											assign node1015 = (inp[13]) ? 4'b1010 : node1016;
												assign node1016 = (inp[6]) ? 4'b0110 : node1017;
													assign node1017 = (inp[10]) ? 4'b1010 : node1018;
														assign node1018 = (inp[1]) ? 4'b0110 : 4'b1110;
									assign node1024 = (inp[8]) ? node1044 : node1025;
										assign node1025 = (inp[11]) ? node1039 : node1026;
											assign node1026 = (inp[6]) ? node1032 : node1027;
												assign node1027 = (inp[13]) ? node1029 : 4'b1110;
													assign node1029 = (inp[9]) ? 4'b1010 : 4'b1110;
												assign node1032 = (inp[12]) ? node1036 : node1033;
													assign node1033 = (inp[9]) ? 4'b0110 : 4'b0000;
													assign node1036 = (inp[10]) ? 4'b1110 : 4'b0110;
											assign node1039 = (inp[6]) ? node1041 : 4'b0110;
												assign node1041 = (inp[1]) ? 4'b0110 : 4'b1110;
										assign node1044 = (inp[9]) ? node1052 : node1045;
											assign node1045 = (inp[11]) ? node1047 : 4'b1111;
												assign node1047 = (inp[12]) ? node1049 : 4'b0111;
													assign node1049 = (inp[13]) ? 4'b0111 : 4'b1111;
											assign node1052 = (inp[12]) ? node1060 : node1053;
												assign node1053 = (inp[1]) ? node1055 : 4'b0111;
													assign node1055 = (inp[10]) ? 4'b0011 : node1056;
														assign node1056 = (inp[11]) ? 4'b1111 : 4'b0111;
												assign node1060 = (inp[13]) ? 4'b0011 : 4'b1011;
						assign node1063 = (inp[3]) ? node1231 : node1064;
							assign node1064 = (inp[11]) ? node1154 : node1065;
								assign node1065 = (inp[6]) ? node1111 : node1066;
									assign node1066 = (inp[1]) ? node1088 : node1067;
										assign node1067 = (inp[9]) ? node1077 : node1068;
											assign node1068 = (inp[10]) ? 4'b1010 : node1069;
												assign node1069 = (inp[4]) ? node1071 : 4'b1111;
													assign node1071 = (inp[2]) ? 4'b1011 : node1072;
														assign node1072 = (inp[8]) ? 4'b1010 : 4'b1011;
											assign node1077 = (inp[12]) ? node1081 : node1078;
												assign node1078 = (inp[10]) ? 4'b1010 : 4'b1110;
												assign node1081 = (inp[4]) ? 4'b0111 : node1082;
													assign node1082 = (inp[10]) ? node1084 : 4'b1011;
														assign node1084 = (inp[13]) ? 4'b1110 : 4'b1111;
										assign node1088 = (inp[13]) ? node1102 : node1089;
											assign node1089 = (inp[9]) ? node1095 : node1090;
												assign node1090 = (inp[2]) ? 4'b0011 : node1091;
													assign node1091 = (inp[8]) ? 4'b1010 : 4'b1011;
												assign node1095 = (inp[2]) ? node1097 : 4'b1111;
													assign node1097 = (inp[12]) ? node1099 : 4'b1110;
														assign node1099 = (inp[4]) ? 4'b1010 : 4'b1110;
											assign node1102 = (inp[12]) ? node1104 : 4'b0010;
												assign node1104 = (inp[2]) ? node1108 : node1105;
													assign node1105 = (inp[8]) ? 4'b0110 : 4'b0111;
													assign node1108 = (inp[9]) ? 4'b0011 : 4'b0110;
									assign node1111 = (inp[13]) ? node1129 : node1112;
										assign node1112 = (inp[8]) ? node1122 : node1113;
											assign node1113 = (inp[2]) ? 4'b0010 : node1114;
												assign node1114 = (inp[10]) ? 4'b0011 : node1115;
													assign node1115 = (inp[12]) ? node1117 : 4'b0111;
														assign node1117 = (inp[9]) ? 4'b0011 : 4'b0111;
											assign node1122 = (inp[2]) ? node1126 : node1123;
												assign node1123 = (inp[9]) ? 4'b0110 : 4'b0010;
												assign node1126 = (inp[1]) ? 4'b1111 : 4'b0111;
										assign node1129 = (inp[1]) ? node1139 : node1130;
											assign node1130 = (inp[10]) ? 4'b0010 : node1131;
												assign node1131 = (inp[12]) ? node1135 : node1132;
													assign node1132 = (inp[4]) ? 4'b0110 : 4'b0010;
													assign node1135 = (inp[4]) ? 4'b0010 : 4'b0110;
											assign node1139 = (inp[9]) ? node1149 : node1140;
												assign node1140 = (inp[2]) ? node1146 : node1141;
													assign node1141 = (inp[12]) ? 4'b1011 : node1142;
														assign node1142 = (inp[4]) ? 4'b1011 : 4'b1111;
													assign node1146 = (inp[10]) ? 4'b1111 : 4'b1110;
												assign node1149 = (inp[4]) ? node1151 : 4'b1110;
													assign node1151 = (inp[10]) ? 4'b1010 : 4'b1110;
								assign node1154 = (inp[6]) ? node1190 : node1155;
									assign node1155 = (inp[8]) ? node1171 : node1156;
										assign node1156 = (inp[2]) ? node1166 : node1157;
											assign node1157 = (inp[12]) ? 4'b0011 : node1158;
												assign node1158 = (inp[10]) ? node1160 : 4'b0111;
													assign node1160 = (inp[1]) ? node1162 : 4'b0011;
														assign node1162 = (inp[9]) ? 4'b0011 : 4'b0111;
											assign node1166 = (inp[9]) ? 4'b0110 : node1167;
												assign node1167 = (inp[4]) ? 4'b0010 : 4'b0110;
										assign node1171 = (inp[2]) ? node1179 : node1172;
											assign node1172 = (inp[1]) ? node1176 : node1173;
												assign node1173 = (inp[4]) ? 4'b0010 : 4'b0110;
												assign node1176 = (inp[12]) ? 4'b1010 : 4'b0010;
											assign node1179 = (inp[1]) ? node1185 : node1180;
												assign node1180 = (inp[13]) ? node1182 : 4'b0111;
													assign node1182 = (inp[10]) ? 4'b1011 : 4'b1111;
												assign node1185 = (inp[13]) ? 4'b1111 : node1186;
													assign node1186 = (inp[9]) ? 4'b1011 : 4'b1111;
									assign node1190 = (inp[1]) ? node1200 : node1191;
										assign node1191 = (inp[2]) ? node1197 : node1192;
											assign node1192 = (inp[8]) ? 4'b1010 : node1193;
												assign node1193 = (inp[4]) ? 4'b1011 : 4'b1111;
											assign node1197 = (inp[13]) ? 4'b1010 : 4'b1110;
										assign node1200 = (inp[13]) ? node1216 : node1201;
											assign node1201 = (inp[8]) ? node1209 : node1202;
												assign node1202 = (inp[2]) ? 4'b1110 : node1203;
													assign node1203 = (inp[12]) ? 4'b1111 : node1204;
														assign node1204 = (inp[4]) ? 4'b1111 : 4'b1011;
												assign node1209 = (inp[2]) ? node1211 : 4'b1110;
													assign node1211 = (inp[10]) ? node1213 : 4'b0011;
														assign node1213 = (inp[9]) ? 4'b0011 : 4'b0111;
											assign node1216 = (inp[9]) ? node1224 : node1217;
												assign node1217 = (inp[4]) ? 4'b0111 : node1218;
													assign node1218 = (inp[12]) ? node1220 : 4'b0111;
														assign node1220 = (inp[8]) ? 4'b0011 : 4'b0010;
												assign node1224 = (inp[2]) ? node1228 : node1225;
													assign node1225 = (inp[8]) ? 4'b0010 : 4'b0011;
													assign node1228 = (inp[8]) ? 4'b0111 : 4'b0110;
							assign node1231 = (inp[9]) ? node1323 : node1232;
								assign node1232 = (inp[4]) ? node1276 : node1233;
									assign node1233 = (inp[11]) ? node1253 : node1234;
										assign node1234 = (inp[12]) ? node1242 : node1235;
											assign node1235 = (inp[8]) ? node1239 : node1236;
												assign node1236 = (inp[6]) ? 4'b0111 : 4'b1111;
												assign node1239 = (inp[2]) ? 4'b0111 : 4'b0110;
											assign node1242 = (inp[10]) ? 4'b1010 : node1243;
												assign node1243 = (inp[13]) ? node1249 : node1244;
													assign node1244 = (inp[6]) ? node1246 : 4'b1110;
														assign node1246 = (inp[8]) ? 4'b1011 : 4'b0110;
													assign node1249 = (inp[8]) ? 4'b0111 : 4'b0110;
										assign node1253 = (inp[13]) ? node1267 : node1254;
											assign node1254 = (inp[8]) ? node1258 : node1255;
												assign node1255 = (inp[10]) ? 4'b0010 : 4'b1010;
												assign node1258 = (inp[2]) ? node1260 : 4'b1010;
													assign node1260 = (inp[6]) ? node1264 : node1261;
														assign node1261 = (inp[12]) ? 4'b0011 : 4'b0111;
														assign node1264 = (inp[1]) ? 4'b0011 : 4'b1011;
											assign node1267 = (inp[12]) ? node1273 : node1268;
												assign node1268 = (inp[8]) ? node1270 : 4'b1110;
													assign node1270 = (inp[1]) ? 4'b0110 : 4'b1110;
												assign node1273 = (inp[6]) ? 4'b1011 : 4'b1010;
									assign node1276 = (inp[12]) ? node1306 : node1277;
										assign node1277 = (inp[11]) ? node1295 : node1278;
											assign node1278 = (inp[6]) ? node1286 : node1279;
												assign node1279 = (inp[2]) ? node1283 : node1280;
													assign node1280 = (inp[8]) ? 4'b1010 : 4'b1011;
													assign node1283 = (inp[1]) ? 4'b0010 : 4'b1010;
												assign node1286 = (inp[1]) ? node1290 : node1287;
													assign node1287 = (inp[10]) ? 4'b0010 : 4'b0011;
													assign node1290 = (inp[10]) ? node1292 : 4'b1010;
														assign node1292 = (inp[2]) ? 4'b1100 : 4'b1101;
											assign node1295 = (inp[10]) ? 4'b0010 : node1296;
												assign node1296 = (inp[8]) ? node1302 : node1297;
													assign node1297 = (inp[2]) ? 4'b0010 : node1298;
														assign node1298 = (inp[13]) ? 4'b0011 : 4'b1011;
													assign node1302 = (inp[1]) ? 4'b0011 : 4'b0010;
										assign node1306 = (inp[10]) ? node1314 : node1307;
											assign node1307 = (inp[8]) ? 4'b1011 : node1308;
												assign node1308 = (inp[1]) ? node1310 : 4'b1100;
													assign node1310 = (inp[13]) ? 4'b1100 : 4'b0010;
											assign node1314 = (inp[6]) ? node1316 : 4'b0100;
												assign node1316 = (inp[11]) ? node1320 : node1317;
													assign node1317 = (inp[1]) ? 4'b1100 : 4'b0100;
													assign node1320 = (inp[13]) ? 4'b0101 : 4'b1101;
								assign node1323 = (inp[4]) ? node1371 : node1324;
									assign node1324 = (inp[12]) ? node1344 : node1325;
										assign node1325 = (inp[1]) ? node1337 : node1326;
											assign node1326 = (inp[8]) ? node1328 : 4'b1010;
												assign node1328 = (inp[2]) ? node1334 : node1329;
													assign node1329 = (inp[11]) ? 4'b1100 : node1330;
														assign node1330 = (inp[10]) ? 4'b1010 : 4'b0010;
													assign node1334 = (inp[11]) ? 4'b0011 : 4'b1011;
											assign node1337 = (inp[8]) ? node1341 : node1338;
												assign node1338 = (inp[2]) ? 4'b0010 : 4'b0011;
												assign node1341 = (inp[6]) ? 4'b1010 : 4'b1011;
										assign node1344 = (inp[11]) ? node1360 : node1345;
											assign node1345 = (inp[10]) ? node1353 : node1346;
												assign node1346 = (inp[13]) ? 4'b1010 : node1347;
													assign node1347 = (inp[8]) ? 4'b0011 : node1348;
														assign node1348 = (inp[6]) ? 4'b0010 : 4'b1010;
												assign node1353 = (inp[6]) ? 4'b0100 : node1354;
													assign node1354 = (inp[8]) ? 4'b1100 : node1355;
														assign node1355 = (inp[2]) ? 4'b1100 : 4'b1101;
											assign node1360 = (inp[1]) ? node1364 : node1361;
												assign node1361 = (inp[6]) ? 4'b1100 : 4'b0100;
												assign node1364 = (inp[6]) ? node1368 : node1365;
													assign node1365 = (inp[2]) ? 4'b1101 : 4'b1100;
													assign node1368 = (inp[8]) ? 4'b0101 : 4'b1101;
									assign node1371 = (inp[10]) ? node1389 : node1372;
										assign node1372 = (inp[6]) ? node1384 : node1373;
											assign node1373 = (inp[13]) ? node1379 : node1374;
												assign node1374 = (inp[1]) ? node1376 : 4'b1100;
													assign node1376 = (inp[2]) ? 4'b1100 : 4'b1101;
												assign node1379 = (inp[11]) ? 4'b1101 : node1380;
													assign node1380 = (inp[2]) ? 4'b0101 : 4'b0100;
											assign node1384 = (inp[1]) ? 4'b1001 : node1385;
												assign node1385 = (inp[11]) ? 4'b0001 : 4'b0101;
										assign node1389 = (inp[6]) ? node1393 : node1390;
											assign node1390 = (inp[12]) ? 4'b0001 : 4'b0101;
											assign node1393 = (inp[11]) ? node1401 : node1394;
												assign node1394 = (inp[8]) ? node1398 : node1395;
													assign node1395 = (inp[1]) ? 4'b0001 : 4'b0101;
													assign node1398 = (inp[12]) ? 4'b0000 : 4'b0100;
												assign node1401 = (inp[13]) ? node1403 : 4'b1000;
													assign node1403 = (inp[12]) ? 4'b1000 : node1404;
														assign node1404 = (inp[1]) ? 4'b0000 : 4'b0001;
				assign node1408 = (inp[11]) ? node2090 : node1409;
					assign node1409 = (inp[6]) ? node1753 : node1410;
						assign node1410 = (inp[1]) ? node1564 : node1411;
							assign node1411 = (inp[2]) ? node1481 : node1412;
								assign node1412 = (inp[8]) ? node1450 : node1413;
									assign node1413 = (inp[3]) ? node1435 : node1414;
										assign node1414 = (inp[12]) ? node1426 : node1415;
											assign node1415 = (inp[13]) ? node1417 : 4'b1101;
												assign node1417 = (inp[10]) ? 4'b1101 : node1418;
													assign node1418 = (inp[9]) ? node1422 : node1419;
														assign node1419 = (inp[4]) ? 4'b1001 : 4'b1101;
														assign node1422 = (inp[4]) ? 4'b1101 : 4'b1001;
											assign node1426 = (inp[15]) ? node1432 : node1427;
												assign node1427 = (inp[13]) ? node1429 : 4'b1001;
													assign node1429 = (inp[0]) ? 4'b1111 : 4'b1101;
												assign node1432 = (inp[13]) ? 4'b1001 : 4'b1011;
										assign node1435 = (inp[15]) ? node1443 : node1436;
											assign node1436 = (inp[0]) ? node1438 : 4'b1001;
												assign node1438 = (inp[9]) ? node1440 : 4'b1111;
													assign node1440 = (inp[12]) ? 4'b1011 : 4'b1111;
											assign node1443 = (inp[0]) ? node1445 : 4'b1111;
												assign node1445 = (inp[12]) ? 4'b1101 : node1446;
													assign node1446 = (inp[13]) ? 4'b1101 : 4'b1001;
									assign node1450 = (inp[12]) ? node1468 : node1451;
										assign node1451 = (inp[15]) ? node1461 : node1452;
											assign node1452 = (inp[0]) ? node1458 : node1453;
												assign node1453 = (inp[9]) ? 4'b1000 : node1454;
													assign node1454 = (inp[4]) ? 4'b1000 : 4'b1100;
												assign node1458 = (inp[3]) ? 4'b1010 : 4'b1000;
											assign node1461 = (inp[0]) ? node1463 : 4'b1110;
												assign node1463 = (inp[4]) ? node1465 : 4'b1010;
													assign node1465 = (inp[13]) ? 4'b1100 : 4'b1000;
										assign node1468 = (inp[0]) ? node1478 : node1469;
											assign node1469 = (inp[15]) ? node1473 : node1470;
												assign node1470 = (inp[3]) ? 4'b1000 : 4'b1100;
												assign node1473 = (inp[3]) ? 4'b1110 : node1474;
													assign node1474 = (inp[10]) ? 4'b1010 : 4'b1000;
											assign node1478 = (inp[15]) ? 4'b1010 : 4'b1110;
								assign node1481 = (inp[8]) ? node1515 : node1482;
									assign node1482 = (inp[13]) ? node1496 : node1483;
										assign node1483 = (inp[12]) ? node1485 : 4'b1000;
											assign node1485 = (inp[10]) ? node1489 : node1486;
												assign node1486 = (inp[15]) ? 4'b1010 : 4'b1000;
												assign node1489 = (inp[15]) ? node1493 : node1490;
													assign node1490 = (inp[3]) ? 4'b1010 : 4'b1000;
													assign node1493 = (inp[9]) ? 4'b1100 : 4'b1000;
										assign node1496 = (inp[15]) ? node1506 : node1497;
											assign node1497 = (inp[0]) ? node1501 : node1498;
												assign node1498 = (inp[12]) ? 4'b1010 : 4'b1100;
												assign node1501 = (inp[12]) ? node1503 : 4'b1010;
													assign node1503 = (inp[9]) ? 4'b1110 : 4'b1010;
											assign node1506 = (inp[9]) ? node1508 : 4'b1000;
												assign node1508 = (inp[0]) ? 4'b1100 : node1509;
													assign node1509 = (inp[4]) ? node1511 : 4'b1000;
														assign node1511 = (inp[12]) ? 4'b1010 : 4'b1110;
									assign node1515 = (inp[13]) ? node1543 : node1516;
										assign node1516 = (inp[3]) ? node1530 : node1517;
											assign node1517 = (inp[10]) ? node1523 : node1518;
												assign node1518 = (inp[15]) ? 4'b1111 : node1519;
													assign node1519 = (inp[9]) ? 4'b1011 : 4'b1001;
												assign node1523 = (inp[4]) ? 4'b1011 : node1524;
													assign node1524 = (inp[0]) ? 4'b1011 : node1525;
														assign node1525 = (inp[15]) ? 4'b1001 : 4'b1011;
											assign node1530 = (inp[12]) ? node1534 : node1531;
												assign node1531 = (inp[0]) ? 4'b1001 : 4'b1011;
												assign node1534 = (inp[0]) ? node1540 : node1535;
													assign node1535 = (inp[10]) ? 4'b1101 : node1536;
														assign node1536 = (inp[9]) ? 4'b1101 : 4'b1001;
													assign node1540 = (inp[9]) ? 4'b1101 : 4'b1111;
										assign node1543 = (inp[10]) ? node1547 : node1544;
											assign node1544 = (inp[3]) ? 4'b0001 : 4'b0011;
											assign node1547 = (inp[15]) ? node1559 : node1548;
												assign node1548 = (inp[4]) ? node1554 : node1549;
													assign node1549 = (inp[9]) ? node1551 : 4'b0011;
														assign node1551 = (inp[0]) ? 4'b0001 : 4'b0011;
													assign node1554 = (inp[0]) ? node1556 : 4'b0101;
														assign node1556 = (inp[3]) ? 4'b0011 : 4'b0001;
												assign node1559 = (inp[3]) ? node1561 : 4'b0101;
													assign node1561 = (inp[0]) ? 4'b0101 : 4'b0111;
							assign node1564 = (inp[13]) ? node1654 : node1565;
								assign node1565 = (inp[8]) ? node1611 : node1566;
									assign node1566 = (inp[2]) ? node1586 : node1567;
										assign node1567 = (inp[0]) ? node1575 : node1568;
											assign node1568 = (inp[15]) ? node1570 : 4'b1001;
												assign node1570 = (inp[10]) ? 4'b1111 : node1571;
													assign node1571 = (inp[9]) ? 4'b1111 : 4'b1101;
											assign node1575 = (inp[12]) ? node1577 : 4'b1011;
												assign node1577 = (inp[15]) ? node1581 : node1578;
													assign node1578 = (inp[3]) ? 4'b1011 : 4'b1001;
													assign node1581 = (inp[4]) ? 4'b1101 : node1582;
														assign node1582 = (inp[9]) ? 4'b1001 : 4'b1001;
										assign node1586 = (inp[3]) ? node1598 : node1587;
											assign node1587 = (inp[12]) ? node1593 : node1588;
												assign node1588 = (inp[4]) ? 4'b1100 : node1589;
													assign node1589 = (inp[10]) ? 4'b1000 : 4'b1010;
												assign node1593 = (inp[15]) ? node1595 : 4'b1010;
													assign node1595 = (inp[10]) ? 4'b1010 : 4'b1110;
											assign node1598 = (inp[0]) ? node1606 : node1599;
												assign node1599 = (inp[15]) ? 4'b1110 : node1600;
													assign node1600 = (inp[10]) ? node1602 : 4'b1100;
														assign node1602 = (inp[9]) ? 4'b1100 : 4'b1000;
												assign node1606 = (inp[15]) ? node1608 : 4'b1010;
													assign node1608 = (inp[12]) ? 4'b1000 : 4'b1100;
									assign node1611 = (inp[2]) ? node1631 : node1612;
										assign node1612 = (inp[9]) ? node1622 : node1613;
											assign node1613 = (inp[12]) ? node1617 : node1614;
												assign node1614 = (inp[0]) ? 4'b1100 : 4'b1110;
												assign node1617 = (inp[4]) ? 4'b1000 : node1618;
													assign node1618 = (inp[10]) ? 4'b1010 : 4'b1110;
											assign node1622 = (inp[3]) ? node1626 : node1623;
												assign node1623 = (inp[4]) ? 4'b1110 : 4'b1010;
												assign node1626 = (inp[0]) ? 4'b1000 : node1627;
													assign node1627 = (inp[15]) ? 4'b1010 : 4'b1000;
										assign node1631 = (inp[15]) ? node1641 : node1632;
											assign node1632 = (inp[4]) ? node1638 : node1633;
												assign node1633 = (inp[3]) ? 4'b0111 : node1634;
													assign node1634 = (inp[0]) ? 4'b0101 : 4'b0111;
												assign node1638 = (inp[12]) ? 4'b0001 : 4'b0101;
											assign node1641 = (inp[0]) ? node1647 : node1642;
												assign node1642 = (inp[4]) ? node1644 : 4'b0011;
													assign node1644 = (inp[9]) ? 4'b0111 : 4'b0011;
												assign node1647 = (inp[12]) ? node1649 : 4'b0101;
													assign node1649 = (inp[9]) ? node1651 : 4'b0011;
														assign node1651 = (inp[4]) ? 4'b0001 : 4'b0101;
								assign node1654 = (inp[8]) ? node1704 : node1655;
									assign node1655 = (inp[2]) ? node1673 : node1656;
										assign node1656 = (inp[9]) ? node1664 : node1657;
											assign node1657 = (inp[4]) ? node1661 : node1658;
												assign node1658 = (inp[10]) ? 4'b0101 : 4'b0111;
												assign node1661 = (inp[12]) ? 4'b0111 : 4'b0011;
											assign node1664 = (inp[12]) ? node1666 : 4'b0111;
												assign node1666 = (inp[4]) ? 4'b0101 : node1667;
													assign node1667 = (inp[10]) ? node1669 : 4'b0011;
														assign node1669 = (inp[0]) ? 4'b0101 : 4'b0111;
										assign node1673 = (inp[4]) ? node1687 : node1674;
											assign node1674 = (inp[9]) ? node1678 : node1675;
												assign node1675 = (inp[0]) ? 4'b0110 : 4'b0010;
												assign node1678 = (inp[3]) ? 4'b0000 : node1679;
													assign node1679 = (inp[10]) ? node1683 : node1680;
														assign node1680 = (inp[12]) ? 4'b0010 : 4'b0000;
														assign node1683 = (inp[12]) ? 4'b0100 : 4'b0010;
											assign node1687 = (inp[9]) ? node1697 : node1688;
												assign node1688 = (inp[12]) ? node1692 : node1689;
													assign node1689 = (inp[15]) ? 4'b0000 : 4'b0010;
													assign node1692 = (inp[10]) ? node1694 : 4'b0000;
														assign node1694 = (inp[0]) ? 4'b0110 : 4'b0100;
												assign node1697 = (inp[12]) ? 4'b0100 : node1698;
													assign node1698 = (inp[3]) ? 4'b0110 : node1699;
														assign node1699 = (inp[0]) ? 4'b0110 : 4'b0100;
									assign node1704 = (inp[2]) ? node1726 : node1705;
										assign node1705 = (inp[9]) ? node1715 : node1706;
											assign node1706 = (inp[12]) ? 4'b0000 : node1707;
												assign node1707 = (inp[4]) ? node1711 : node1708;
													assign node1708 = (inp[10]) ? 4'b0110 : 4'b0100;
													assign node1711 = (inp[3]) ? 4'b0000 : 4'b0010;
											assign node1715 = (inp[15]) ? node1721 : node1716;
												assign node1716 = (inp[10]) ? node1718 : 4'b0100;
													assign node1718 = (inp[12]) ? 4'b0000 : 4'b0100;
												assign node1721 = (inp[0]) ? node1723 : 4'b0110;
													assign node1723 = (inp[12]) ? 4'b0100 : 4'b0000;
										assign node1726 = (inp[15]) ? node1742 : node1727;
											assign node1727 = (inp[0]) ? node1733 : node1728;
												assign node1728 = (inp[9]) ? node1730 : 4'b0111;
													assign node1730 = (inp[4]) ? 4'b0101 : 4'b0001;
												assign node1733 = (inp[10]) ? 4'b0111 : node1734;
													assign node1734 = (inp[4]) ? node1738 : node1735;
														assign node1735 = (inp[9]) ? 4'b0001 : 4'b0101;
														assign node1738 = (inp[3]) ? 4'b0011 : 4'b0111;
											assign node1742 = (inp[3]) ? node1750 : node1743;
												assign node1743 = (inp[4]) ? node1747 : node1744;
													assign node1744 = (inp[0]) ? 4'b0011 : 4'b0001;
													assign node1747 = (inp[0]) ? 4'b0101 : 4'b0111;
												assign node1750 = (inp[0]) ? 4'b0001 : 4'b0011;
						assign node1753 = (inp[1]) ? node1927 : node1754;
							assign node1754 = (inp[13]) ? node1836 : node1755;
								assign node1755 = (inp[4]) ? node1791 : node1756;
									assign node1756 = (inp[9]) ? node1766 : node1757;
										assign node1757 = (inp[10]) ? node1761 : node1758;
											assign node1758 = (inp[12]) ? 4'b0100 : 4'b0111;
											assign node1761 = (inp[2]) ? node1763 : 4'b0011;
												assign node1763 = (inp[3]) ? 4'b0000 : 4'b0001;
										assign node1766 = (inp[10]) ? node1784 : node1767;
											assign node1767 = (inp[0]) ? node1777 : node1768;
												assign node1768 = (inp[8]) ? node1774 : node1769;
													assign node1769 = (inp[2]) ? node1771 : 4'b0011;
														assign node1771 = (inp[15]) ? 4'b0010 : 4'b0000;
													assign node1774 = (inp[2]) ? 4'b0011 : 4'b0000;
												assign node1777 = (inp[2]) ? 4'b0000 : node1778;
													assign node1778 = (inp[8]) ? node1780 : 4'b0011;
														assign node1780 = (inp[15]) ? 4'b0000 : 4'b0000;
											assign node1784 = (inp[15]) ? node1786 : 4'b0001;
												assign node1786 = (inp[12]) ? 4'b0111 : node1787;
													assign node1787 = (inp[3]) ? 4'b0010 : 4'b0011;
									assign node1791 = (inp[15]) ? node1815 : node1792;
										assign node1792 = (inp[0]) ? node1806 : node1793;
											assign node1793 = (inp[3]) ? node1799 : node1794;
												assign node1794 = (inp[12]) ? node1796 : 4'b0101;
													assign node1796 = (inp[10]) ? 4'b0001 : 4'b0101;
												assign node1799 = (inp[9]) ? 4'b0100 : node1800;
													assign node1800 = (inp[8]) ? 4'b0000 : node1801;
														assign node1801 = (inp[12]) ? 4'b0101 : 4'b0001;
											assign node1806 = (inp[3]) ? 4'b0111 : node1807;
												assign node1807 = (inp[2]) ? 4'b0110 : node1808;
													assign node1808 = (inp[10]) ? node1810 : 4'b0001;
														assign node1810 = (inp[9]) ? 4'b0010 : 4'b0110;
										assign node1815 = (inp[0]) ? node1825 : node1816;
											assign node1816 = (inp[9]) ? 4'b0111 : node1817;
												assign node1817 = (inp[3]) ? node1821 : node1818;
													assign node1818 = (inp[2]) ? 4'b0111 : 4'b0110;
													assign node1821 = (inp[2]) ? 4'b0011 : 4'b0010;
											assign node1825 = (inp[12]) ? node1827 : 4'b0011;
												assign node1827 = (inp[3]) ? node1833 : node1828;
													assign node1828 = (inp[10]) ? node1830 : 4'b0011;
														assign node1830 = (inp[2]) ? 4'b0000 : 4'b0001;
													assign node1833 = (inp[2]) ? 4'b0101 : 4'b0000;
								assign node1836 = (inp[2]) ? node1888 : node1837;
									assign node1837 = (inp[8]) ? node1869 : node1838;
										assign node1838 = (inp[3]) ? node1850 : node1839;
											assign node1839 = (inp[9]) ? node1845 : node1840;
												assign node1840 = (inp[15]) ? node1842 : 4'b0111;
													assign node1842 = (inp[0]) ? 4'b0011 : 4'b0001;
												assign node1845 = (inp[15]) ? 4'b0111 : node1846;
													assign node1846 = (inp[0]) ? 4'b0111 : 4'b0011;
											assign node1850 = (inp[0]) ? node1858 : node1851;
												assign node1851 = (inp[15]) ? 4'b0011 : node1852;
													assign node1852 = (inp[10]) ? 4'b0001 : node1853;
														assign node1853 = (inp[4]) ? 4'b0101 : 4'b0001;
												assign node1858 = (inp[15]) ? node1864 : node1859;
													assign node1859 = (inp[4]) ? node1861 : 4'b0111;
														assign node1861 = (inp[10]) ? 4'b0011 : 4'b0011;
													assign node1864 = (inp[9]) ? node1866 : 4'b0101;
														assign node1866 = (inp[4]) ? 4'b0101 : 4'b0001;
										assign node1869 = (inp[3]) ? node1881 : node1870;
											assign node1870 = (inp[4]) ? node1878 : node1871;
												assign node1871 = (inp[9]) ? node1873 : 4'b0100;
													assign node1873 = (inp[10]) ? node1875 : 4'b0000;
														assign node1875 = (inp[15]) ? 4'b0110 : 4'b0010;
												assign node1878 = (inp[12]) ? 4'b0010 : 4'b0000;
											assign node1881 = (inp[15]) ? node1883 : 4'b0110;
												assign node1883 = (inp[0]) ? node1885 : 4'b0110;
													assign node1885 = (inp[9]) ? 4'b0000 : 4'b0100;
									assign node1888 = (inp[8]) ? node1908 : node1889;
										assign node1889 = (inp[3]) ? node1897 : node1890;
											assign node1890 = (inp[0]) ? node1892 : 4'b0010;
												assign node1892 = (inp[10]) ? node1894 : 4'b0110;
													assign node1894 = (inp[9]) ? 4'b0110 : 4'b0010;
											assign node1897 = (inp[12]) ? 4'b0010 : node1898;
												assign node1898 = (inp[10]) ? 4'b0000 : node1899;
													assign node1899 = (inp[15]) ? node1903 : node1900;
														assign node1900 = (inp[9]) ? 4'b0000 : 4'b0000;
														assign node1903 = (inp[4]) ? 4'b0110 : 4'b0100;
										assign node1908 = (inp[4]) ? node1922 : node1909;
											assign node1909 = (inp[9]) ? node1917 : node1910;
												assign node1910 = (inp[12]) ? node1912 : 4'b1111;
													assign node1912 = (inp[10]) ? 4'b1011 : node1913;
														assign node1913 = (inp[0]) ? 4'b1001 : 4'b1011;
												assign node1917 = (inp[12]) ? 4'b1111 : node1918;
													assign node1918 = (inp[10]) ? 4'b1111 : 4'b1001;
											assign node1922 = (inp[12]) ? node1924 : 4'b1011;
												assign node1924 = (inp[10]) ? 4'b1011 : 4'b1111;
							assign node1927 = (inp[13]) ? node2001 : node1928;
								assign node1928 = (inp[2]) ? node1968 : node1929;
									assign node1929 = (inp[8]) ? node1949 : node1930;
										assign node1930 = (inp[4]) ? node1936 : node1931;
											assign node1931 = (inp[10]) ? node1933 : 4'b0101;
												assign node1933 = (inp[15]) ? 4'b0111 : 4'b0101;
											assign node1936 = (inp[10]) ? node1940 : node1937;
												assign node1937 = (inp[15]) ? 4'b0011 : 4'b0001;
												assign node1940 = (inp[15]) ? node1944 : node1941;
													assign node1941 = (inp[12]) ? 4'b0111 : 4'b0011;
													assign node1944 = (inp[9]) ? node1946 : 4'b0101;
														assign node1946 = (inp[12]) ? 4'b0001 : 4'b0101;
										assign node1949 = (inp[10]) ? node1961 : node1950;
											assign node1950 = (inp[9]) ? node1954 : node1951;
												assign node1951 = (inp[15]) ? 4'b0000 : 4'b0110;
												assign node1954 = (inp[15]) ? 4'b0010 : node1955;
													assign node1955 = (inp[3]) ? node1957 : 4'b0000;
														assign node1957 = (inp[12]) ? 4'b0010 : 4'b0000;
											assign node1961 = (inp[4]) ? node1963 : 4'b0100;
												assign node1963 = (inp[12]) ? 4'b0000 : node1964;
													assign node1964 = (inp[9]) ? 4'b0100 : 4'b0000;
									assign node1968 = (inp[8]) ? node1982 : node1969;
										assign node1969 = (inp[4]) ? node1977 : node1970;
											assign node1970 = (inp[0]) ? node1972 : 4'b0000;
												assign node1972 = (inp[12]) ? node1974 : 4'b0110;
													assign node1974 = (inp[15]) ? 4'b0100 : 4'b0000;
											assign node1977 = (inp[0]) ? 4'b0110 : node1978;
												assign node1978 = (inp[15]) ? 4'b0110 : 4'b0010;
										assign node1982 = (inp[3]) ? node1988 : node1983;
											assign node1983 = (inp[4]) ? 4'b1011 : node1984;
												assign node1984 = (inp[0]) ? 4'b1011 : 4'b1001;
											assign node1988 = (inp[9]) ? node1996 : node1989;
												assign node1989 = (inp[4]) ? 4'b1101 : node1990;
													assign node1990 = (inp[12]) ? 4'b1001 : node1991;
														assign node1991 = (inp[0]) ? 4'b1011 : 4'b1001;
												assign node1996 = (inp[10]) ? node1998 : 4'b1101;
													assign node1998 = (inp[0]) ? 4'b1101 : 4'b1111;
								assign node2001 = (inp[10]) ? node2057 : node2002;
									assign node2002 = (inp[0]) ? node2022 : node2003;
										assign node2003 = (inp[15]) ? node2013 : node2004;
											assign node2004 = (inp[3]) ? node2010 : node2005;
												assign node2005 = (inp[4]) ? node2007 : 4'b1011;
													assign node2007 = (inp[12]) ? 4'b1100 : 4'b1010;
												assign node2010 = (inp[2]) ? 4'b1100 : 4'b1000;
											assign node2013 = (inp[9]) ? node2017 : node2014;
												assign node2014 = (inp[4]) ? 4'b1110 : 4'b1000;
												assign node2017 = (inp[4]) ? node2019 : 4'b1111;
													assign node2019 = (inp[3]) ? 4'b1011 : 4'b1010;
										assign node2022 = (inp[12]) ? node2044 : node2023;
											assign node2023 = (inp[2]) ? node2037 : node2024;
												assign node2024 = (inp[8]) ? node2030 : node2025;
													assign node2025 = (inp[4]) ? node2027 : 4'b1111;
														assign node2027 = (inp[15]) ? 4'b1011 : 4'b1001;
													assign node2030 = (inp[4]) ? node2034 : node2031;
														assign node2031 = (inp[15]) ? 4'b1000 : 4'b1010;
														assign node2034 = (inp[3]) ? 4'b1110 : 4'b1010;
												assign node2037 = (inp[3]) ? node2039 : 4'b1111;
													assign node2039 = (inp[9]) ? 4'b1111 : node2040;
														assign node2040 = (inp[4]) ? 4'b1011 : 4'b1111;
											assign node2044 = (inp[15]) ? node2050 : node2045;
												assign node2045 = (inp[8]) ? node2047 : 4'b1010;
													assign node2047 = (inp[4]) ? 4'b1111 : 4'b1001;
												assign node2050 = (inp[8]) ? node2052 : 4'b1001;
													assign node2052 = (inp[9]) ? node2054 : 4'b1101;
														assign node2054 = (inp[4]) ? 4'b1001 : 4'b1101;
									assign node2057 = (inp[15]) ? node2073 : node2058;
										assign node2058 = (inp[0]) ? node2064 : node2059;
											assign node2059 = (inp[8]) ? 4'b1101 : node2060;
												assign node2060 = (inp[12]) ? 4'b1001 : 4'b1101;
											assign node2064 = (inp[4]) ? node2068 : node2065;
												assign node2065 = (inp[3]) ? 4'b1011 : 4'b1111;
												assign node2068 = (inp[3]) ? node2070 : 4'b1111;
													assign node2070 = (inp[2]) ? 4'b1110 : 4'b1111;
										assign node2073 = (inp[0]) ? node2083 : node2074;
											assign node2074 = (inp[9]) ? node2076 : 4'b1110;
												assign node2076 = (inp[4]) ? node2080 : node2077;
													assign node2077 = (inp[12]) ? 4'b1111 : 4'b1110;
													assign node2080 = (inp[2]) ? 4'b1011 : 4'b1010;
											assign node2083 = (inp[2]) ? node2087 : node2084;
												assign node2084 = (inp[8]) ? 4'b1100 : 4'b1101;
												assign node2087 = (inp[8]) ? 4'b1001 : 4'b1100;
					assign node2090 = (inp[6]) ? node2458 : node2091;
						assign node2091 = (inp[13]) ? node2251 : node2092;
							assign node2092 = (inp[2]) ? node2168 : node2093;
								assign node2093 = (inp[8]) ? node2139 : node2094;
									assign node2094 = (inp[3]) ? node2118 : node2095;
										assign node2095 = (inp[12]) ? node2109 : node2096;
											assign node2096 = (inp[1]) ? node2102 : node2097;
												assign node2097 = (inp[4]) ? node2099 : 4'b0101;
													assign node2099 = (inp[9]) ? 4'b0101 : 4'b0001;
												assign node2102 = (inp[4]) ? 4'b0101 : node2103;
													assign node2103 = (inp[0]) ? 4'b0001 : node2104;
														assign node2104 = (inp[15]) ? 4'b0001 : 4'b0011;
											assign node2109 = (inp[4]) ? node2115 : node2110;
												assign node2110 = (inp[0]) ? node2112 : 4'b0001;
													assign node2112 = (inp[9]) ? 4'b0101 : 4'b0111;
												assign node2115 = (inp[0]) ? 4'b0001 : 4'b0011;
										assign node2118 = (inp[9]) ? node2124 : node2119;
											assign node2119 = (inp[4]) ? node2121 : 4'b0111;
												assign node2121 = (inp[10]) ? 4'b0111 : 4'b0011;
											assign node2124 = (inp[4]) ? node2134 : node2125;
												assign node2125 = (inp[0]) ? node2131 : node2126;
													assign node2126 = (inp[1]) ? 4'b0101 : node2127;
														assign node2127 = (inp[15]) ? 4'b0011 : 4'b0001;
													assign node2131 = (inp[15]) ? 4'b0001 : 4'b0011;
												assign node2134 = (inp[0]) ? node2136 : 4'b0101;
													assign node2136 = (inp[15]) ? 4'b0101 : 4'b0111;
									assign node2139 = (inp[10]) ? node2157 : node2140;
										assign node2140 = (inp[15]) ? node2152 : node2141;
											assign node2141 = (inp[3]) ? node2149 : node2142;
												assign node2142 = (inp[0]) ? 4'b0000 : node2143;
													assign node2143 = (inp[9]) ? 4'b0100 : node2144;
														assign node2144 = (inp[1]) ? 4'b0010 : 4'b0110;
												assign node2149 = (inp[0]) ? 4'b0110 : 4'b0100;
											assign node2152 = (inp[12]) ? 4'b0100 : node2153;
												assign node2153 = (inp[9]) ? 4'b0000 : 4'b0100;
										assign node2157 = (inp[4]) ? node2159 : 4'b0010;
											assign node2159 = (inp[3]) ? node2161 : 4'b0000;
												assign node2161 = (inp[15]) ? node2165 : node2162;
													assign node2162 = (inp[1]) ? 4'b0010 : 4'b0000;
													assign node2165 = (inp[1]) ? 4'b0000 : 4'b0010;
								assign node2168 = (inp[8]) ? node2218 : node2169;
									assign node2169 = (inp[4]) ? node2199 : node2170;
										assign node2170 = (inp[9]) ? node2178 : node2171;
											assign node2171 = (inp[12]) ? 4'b0010 : node2172;
												assign node2172 = (inp[0]) ? node2174 : 4'b0100;
													assign node2174 = (inp[1]) ? 4'b0110 : 4'b0100;
											assign node2178 = (inp[12]) ? node2188 : node2179;
												assign node2179 = (inp[3]) ? node2181 : 4'b0010;
													assign node2181 = (inp[10]) ? node2185 : node2182;
														assign node2182 = (inp[15]) ? 4'b0000 : 4'b0010;
														assign node2185 = (inp[1]) ? 4'b0010 : 4'b0000;
												assign node2188 = (inp[10]) ? node2194 : node2189;
													assign node2189 = (inp[3]) ? node2191 : 4'b0000;
														assign node2191 = (inp[0]) ? 4'b0010 : 4'b0000;
													assign node2194 = (inp[0]) ? 4'b0100 : node2195;
														assign node2195 = (inp[15]) ? 4'b0110 : 4'b0100;
										assign node2199 = (inp[9]) ? node2209 : node2200;
											assign node2200 = (inp[1]) ? node2206 : node2201;
												assign node2201 = (inp[12]) ? node2203 : 4'b0010;
													assign node2203 = (inp[0]) ? 4'b0000 : 4'b0110;
												assign node2206 = (inp[0]) ? 4'b0100 : 4'b0000;
											assign node2209 = (inp[10]) ? node2215 : node2210;
												assign node2210 = (inp[15]) ? 4'b0100 : node2211;
													assign node2211 = (inp[0]) ? 4'b0110 : 4'b0100;
												assign node2215 = (inp[12]) ? 4'b0000 : 4'b0100;
									assign node2218 = (inp[1]) ? node2240 : node2219;
										assign node2219 = (inp[3]) ? node2229 : node2220;
											assign node2220 = (inp[9]) ? node2222 : 4'b0011;
												assign node2222 = (inp[12]) ? node2226 : node2223;
													assign node2223 = (inp[4]) ? 4'b0111 : 4'b0001;
													assign node2226 = (inp[10]) ? 4'b0001 : 4'b0011;
											assign node2229 = (inp[9]) ? node2235 : node2230;
												assign node2230 = (inp[15]) ? 4'b0101 : node2231;
													assign node2231 = (inp[0]) ? 4'b0111 : 4'b0101;
												assign node2235 = (inp[4]) ? 4'b0111 : node2236;
													assign node2236 = (inp[12]) ? 4'b0111 : 4'b0011;
										assign node2240 = (inp[15]) ? 4'b1001 : node2241;
											assign node2241 = (inp[0]) ? node2245 : node2242;
												assign node2242 = (inp[9]) ? 4'b1101 : 4'b1001;
												assign node2245 = (inp[10]) ? node2247 : 4'b1111;
													assign node2247 = (inp[4]) ? 4'b1011 : 4'b1111;
							assign node2251 = (inp[1]) ? node2345 : node2252;
								assign node2252 = (inp[2]) ? node2300 : node2253;
									assign node2253 = (inp[8]) ? node2271 : node2254;
										assign node2254 = (inp[9]) ? node2268 : node2255;
											assign node2255 = (inp[4]) ? node2261 : node2256;
												assign node2256 = (inp[3]) ? 4'b0111 : node2257;
													assign node2257 = (inp[10]) ? 4'b0001 : 4'b0101;
												assign node2261 = (inp[3]) ? 4'b0001 : node2262;
													assign node2262 = (inp[10]) ? node2264 : 4'b0011;
														assign node2264 = (inp[12]) ? 4'b0111 : 4'b0011;
											assign node2268 = (inp[4]) ? 4'b0111 : 4'b0011;
										assign node2271 = (inp[12]) ? node2289 : node2272;
											assign node2272 = (inp[3]) ? node2280 : node2273;
												assign node2273 = (inp[0]) ? 4'b0010 : node2274;
													assign node2274 = (inp[9]) ? 4'b0010 : node2275;
														assign node2275 = (inp[4]) ? 4'b0000 : 4'b0100;
												assign node2280 = (inp[10]) ? node2284 : node2281;
													assign node2281 = (inp[4]) ? 4'b0100 : 4'b0010;
													assign node2284 = (inp[9]) ? 4'b0110 : node2285;
														assign node2285 = (inp[0]) ? 4'b0100 : 4'b0110;
											assign node2289 = (inp[10]) ? node2295 : node2290;
												assign node2290 = (inp[9]) ? 4'b0000 : node2291;
													assign node2291 = (inp[4]) ? 4'b0000 : 4'b0100;
												assign node2295 = (inp[0]) ? 4'b0010 : node2296;
													assign node2296 = (inp[4]) ? 4'b0010 : 4'b0100;
									assign node2300 = (inp[8]) ? node2322 : node2301;
										assign node2301 = (inp[4]) ? node2313 : node2302;
											assign node2302 = (inp[9]) ? node2306 : node2303;
												assign node2303 = (inp[0]) ? 4'b0110 : 4'b0100;
												assign node2306 = (inp[15]) ? node2310 : node2307;
													assign node2307 = (inp[12]) ? 4'b0010 : 4'b0000;
													assign node2310 = (inp[10]) ? 4'b0100 : 4'b0000;
											assign node2313 = (inp[3]) ? node2315 : 4'b0010;
												assign node2315 = (inp[15]) ? node2319 : node2316;
													assign node2316 = (inp[12]) ? 4'b0000 : 4'b0100;
													assign node2319 = (inp[0]) ? 4'b0000 : 4'b0010;
										assign node2322 = (inp[4]) ? node2340 : node2323;
											assign node2323 = (inp[9]) ? node2333 : node2324;
												assign node2324 = (inp[3]) ? node2326 : 4'b1001;
													assign node2326 = (inp[15]) ? node2330 : node2327;
														assign node2327 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node2330 = (inp[0]) ? 4'b1001 : 4'b1011;
												assign node2333 = (inp[12]) ? node2337 : node2334;
													assign node2334 = (inp[10]) ? 4'b1101 : 4'b1001;
													assign node2337 = (inp[10]) ? 4'b1111 : 4'b1101;
											assign node2340 = (inp[15]) ? 4'b1001 : node2341;
												assign node2341 = (inp[0]) ? 4'b1011 : 4'b1001;
								assign node2345 = (inp[10]) ? node2415 : node2346;
									assign node2346 = (inp[0]) ? node2382 : node2347;
										assign node2347 = (inp[4]) ? node2363 : node2348;
											assign node2348 = (inp[9]) ? node2358 : node2349;
												assign node2349 = (inp[12]) ? node2351 : 4'b1100;
													assign node2351 = (inp[2]) ? node2355 : node2352;
														assign node2352 = (inp[8]) ? 4'b1000 : 4'b1001;
														assign node2355 = (inp[8]) ? 4'b1001 : 4'b1010;
												assign node2358 = (inp[12]) ? 4'b1100 : node2359;
													assign node2359 = (inp[15]) ? 4'b1010 : 4'b1000;
											assign node2363 = (inp[9]) ? node2375 : node2364;
												assign node2364 = (inp[12]) ? node2372 : node2365;
													assign node2365 = (inp[2]) ? node2369 : node2366;
														assign node2366 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node2369 = (inp[15]) ? 4'b1000 : 4'b1010;
													assign node2372 = (inp[3]) ? 4'b1111 : 4'b1110;
												assign node2375 = (inp[15]) ? node2379 : node2376;
													assign node2376 = (inp[2]) ? 4'b1001 : 4'b1101;
													assign node2379 = (inp[2]) ? 4'b1111 : 4'b1010;
										assign node2382 = (inp[15]) ? node2398 : node2383;
											assign node2383 = (inp[12]) ? node2391 : node2384;
												assign node2384 = (inp[3]) ? node2388 : node2385;
													assign node2385 = (inp[8]) ? 4'b1000 : 4'b1101;
													assign node2388 = (inp[2]) ? 4'b1111 : 4'b1011;
												assign node2391 = (inp[2]) ? node2395 : node2392;
													assign node2392 = (inp[3]) ? 4'b1010 : 4'b1110;
													assign node2395 = (inp[3]) ? 4'b1010 : 4'b1011;
											assign node2398 = (inp[4]) ? node2404 : node2399;
												assign node2399 = (inp[12]) ? 4'b1011 : node2400;
													assign node2400 = (inp[3]) ? 4'b1101 : 4'b1110;
												assign node2404 = (inp[3]) ? node2412 : node2405;
													assign node2405 = (inp[2]) ? node2409 : node2406;
														assign node2406 = (inp[8]) ? 4'b1100 : 4'b1001;
														assign node2409 = (inp[8]) ? 4'b1101 : 4'b1100;
													assign node2412 = (inp[8]) ? 4'b1001 : 4'b1000;
									assign node2415 = (inp[4]) ? node2441 : node2416;
										assign node2416 = (inp[9]) ? node2424 : node2417;
											assign node2417 = (inp[0]) ? node2421 : node2418;
												assign node2418 = (inp[12]) ? 4'b1010 : 4'b1011;
												assign node2421 = (inp[15]) ? 4'b1010 : 4'b1000;
											assign node2424 = (inp[2]) ? node2432 : node2425;
												assign node2425 = (inp[8]) ? 4'b1110 : node2426;
													assign node2426 = (inp[3]) ? node2428 : 4'b1111;
														assign node2428 = (inp[0]) ? 4'b1101 : 4'b1111;
												assign node2432 = (inp[8]) ? node2438 : node2433;
													assign node2433 = (inp[0]) ? node2435 : 4'b1100;
														assign node2435 = (inp[15]) ? 4'b1100 : 4'b1110;
													assign node2438 = (inp[15]) ? 4'b1111 : 4'b1101;
										assign node2441 = (inp[9]) ? node2449 : node2442;
											assign node2442 = (inp[3]) ? node2444 : 4'b1110;
												assign node2444 = (inp[12]) ? node2446 : 4'b1100;
													assign node2446 = (inp[15]) ? 4'b1100 : 4'b1111;
											assign node2449 = (inp[3]) ? node2453 : node2450;
												assign node2450 = (inp[2]) ? 4'b1010 : 4'b1011;
												assign node2453 = (inp[2]) ? node2455 : 4'b1000;
													assign node2455 = (inp[8]) ? 4'b1001 : 4'b1000;
						assign node2458 = (inp[13]) ? node2668 : node2459;
							assign node2459 = (inp[1]) ? node2577 : node2460;
								assign node2460 = (inp[4]) ? node2518 : node2461;
									assign node2461 = (inp[2]) ? node2491 : node2462;
										assign node2462 = (inp[8]) ? node2468 : node2463;
											assign node2463 = (inp[15]) ? node2465 : 4'b1011;
												assign node2465 = (inp[12]) ? 4'b1001 : 4'b1101;
											assign node2468 = (inp[12]) ? node2484 : node2469;
												assign node2469 = (inp[0]) ? node2477 : node2470;
													assign node2470 = (inp[10]) ? node2474 : node2471;
														assign node2471 = (inp[9]) ? 4'b1000 : 4'b1100;
														assign node2474 = (inp[15]) ? 4'b1000 : 4'b1010;
													assign node2477 = (inp[9]) ? node2481 : node2478;
														assign node2478 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node2481 = (inp[15]) ? 4'b1000 : 4'b1010;
												assign node2484 = (inp[9]) ? 4'b1100 : node2485;
													assign node2485 = (inp[0]) ? 4'b1000 : node2486;
														assign node2486 = (inp[10]) ? 4'b1000 : 4'b1010;
										assign node2491 = (inp[8]) ? node2507 : node2492;
											assign node2492 = (inp[0]) ? node2500 : node2493;
												assign node2493 = (inp[12]) ? node2495 : 4'b1000;
													assign node2495 = (inp[10]) ? node2497 : 4'b1010;
														assign node2497 = (inp[15]) ? 4'b1000 : 4'b1000;
												assign node2500 = (inp[3]) ? node2502 : 4'b1010;
													assign node2502 = (inp[15]) ? node2504 : 4'b1110;
														assign node2504 = (inp[12]) ? 4'b1000 : 4'b1100;
											assign node2507 = (inp[9]) ? node2515 : node2508;
												assign node2508 = (inp[10]) ? node2512 : node2509;
													assign node2509 = (inp[12]) ? 4'b1001 : 4'b1101;
													assign node2512 = (inp[0]) ? 4'b1011 : 4'b1001;
												assign node2515 = (inp[12]) ? 4'b1111 : 4'b1011;
									assign node2518 = (inp[9]) ? node2548 : node2519;
										assign node2519 = (inp[12]) ? node2533 : node2520;
											assign node2520 = (inp[10]) ? node2526 : node2521;
												assign node2521 = (inp[2]) ? node2523 : 4'b1010;
													assign node2523 = (inp[15]) ? 4'b1001 : 4'b1000;
												assign node2526 = (inp[0]) ? node2530 : node2527;
													assign node2527 = (inp[2]) ? 4'b1100 : 4'b1101;
													assign node2530 = (inp[3]) ? 4'b1110 : 4'b1100;
											assign node2533 = (inp[3]) ? node2535 : 4'b1101;
												assign node2535 = (inp[10]) ? node2543 : node2536;
													assign node2536 = (inp[0]) ? node2540 : node2537;
														assign node2537 = (inp[8]) ? 4'b1111 : 4'b1110;
														assign node2540 = (inp[8]) ? 4'b1110 : 4'b1110;
													assign node2543 = (inp[8]) ? node2545 : 4'b1111;
														assign node2545 = (inp[2]) ? 4'b1111 : 4'b1110;
										assign node2548 = (inp[10]) ? node2562 : node2549;
											assign node2549 = (inp[12]) ? node2555 : node2550;
												assign node2550 = (inp[2]) ? 4'b1100 : node2551;
													assign node2551 = (inp[0]) ? 4'b1111 : 4'b1110;
												assign node2555 = (inp[3]) ? node2559 : node2556;
													assign node2556 = (inp[8]) ? 4'b1001 : 4'b1011;
													assign node2559 = (inp[0]) ? 4'b1010 : 4'b1000;
											assign node2562 = (inp[15]) ? node2570 : node2563;
												assign node2563 = (inp[0]) ? 4'b1011 : node2564;
													assign node2564 = (inp[8]) ? 4'b1001 : node2565;
														assign node2565 = (inp[3]) ? 4'b1001 : 4'b1000;
												assign node2570 = (inp[0]) ? 4'b1001 : node2571;
													assign node2571 = (inp[12]) ? 4'b1010 : node2572;
														assign node2572 = (inp[8]) ? 4'b1011 : 4'b1010;
								assign node2577 = (inp[2]) ? node2629 : node2578;
									assign node2578 = (inp[8]) ? node2606 : node2579;
										assign node2579 = (inp[4]) ? node2593 : node2580;
											assign node2580 = (inp[9]) ? node2586 : node2581;
												assign node2581 = (inp[10]) ? node2583 : 4'b1101;
													assign node2583 = (inp[15]) ? 4'b1011 : 4'b1001;
												assign node2586 = (inp[10]) ? 4'b1101 : node2587;
													assign node2587 = (inp[15]) ? node2589 : 4'b1111;
														assign node2589 = (inp[0]) ? 4'b1101 : 4'b1111;
											assign node2593 = (inp[10]) ? node2601 : node2594;
												assign node2594 = (inp[15]) ? node2596 : 4'b1011;
													assign node2596 = (inp[12]) ? 4'b1111 : node2597;
														assign node2597 = (inp[3]) ? 4'b1011 : 4'b1111;
												assign node2601 = (inp[9]) ? 4'b1011 : node2602;
													assign node2602 = (inp[12]) ? 4'b1101 : 4'b1111;
										assign node2606 = (inp[4]) ? node2620 : node2607;
											assign node2607 = (inp[0]) ? 4'b1110 : node2608;
												assign node2608 = (inp[10]) ? node2616 : node2609;
													assign node2609 = (inp[12]) ? node2613 : node2610;
														assign node2610 = (inp[9]) ? 4'b1010 : 4'b1110;
														assign node2613 = (inp[9]) ? 4'b1100 : 4'b1010;
													assign node2616 = (inp[15]) ? 4'b1000 : 4'b1100;
											assign node2620 = (inp[9]) ? node2622 : 4'b1000;
												assign node2622 = (inp[0]) ? node2626 : node2623;
													assign node2623 = (inp[15]) ? 4'b1010 : 4'b1000;
													assign node2626 = (inp[15]) ? 4'b1000 : 4'b1010;
									assign node2629 = (inp[8]) ? node2649 : node2630;
										assign node2630 = (inp[12]) ? node2642 : node2631;
											assign node2631 = (inp[10]) ? node2633 : 4'b1100;
												assign node2633 = (inp[15]) ? node2637 : node2634;
													assign node2634 = (inp[0]) ? 4'b1110 : 4'b1010;
													assign node2637 = (inp[9]) ? node2639 : 4'b1000;
														assign node2639 = (inp[4]) ? 4'b1000 : 4'b1100;
											assign node2642 = (inp[9]) ? node2646 : node2643;
												assign node2643 = (inp[4]) ? 4'b1110 : 4'b1010;
												assign node2646 = (inp[4]) ? 4'b1000 : 4'b1110;
										assign node2649 = (inp[15]) ? node2655 : node2650;
											assign node2650 = (inp[0]) ? 4'b0111 : node2651;
												assign node2651 = (inp[12]) ? 4'b0001 : 4'b0101;
											assign node2655 = (inp[9]) ? node2659 : node2656;
												assign node2656 = (inp[12]) ? 4'b0011 : 4'b0001;
												assign node2659 = (inp[0]) ? node2663 : node2660;
													assign node2660 = (inp[10]) ? 4'b0011 : 4'b0111;
													assign node2663 = (inp[12]) ? 4'b0101 : node2664;
														assign node2664 = (inp[4]) ? 4'b0001 : 4'b0001;
							assign node2668 = (inp[1]) ? node2736 : node2669;
								assign node2669 = (inp[8]) ? node2707 : node2670;
									assign node2670 = (inp[2]) ? node2694 : node2671;
										assign node2671 = (inp[9]) ? node2689 : node2672;
											assign node2672 = (inp[3]) ? node2680 : node2673;
												assign node2673 = (inp[15]) ? 4'b1111 : node2674;
													assign node2674 = (inp[12]) ? 4'b1011 : node2675;
														assign node2675 = (inp[4]) ? 4'b1011 : 4'b1111;
												assign node2680 = (inp[4]) ? node2686 : node2681;
													assign node2681 = (inp[12]) ? 4'b1011 : node2682;
														assign node2682 = (inp[0]) ? 4'b1001 : 4'b1011;
													assign node2686 = (inp[0]) ? 4'b1101 : 4'b1001;
											assign node2689 = (inp[12]) ? node2691 : 4'b1001;
												assign node2691 = (inp[4]) ? 4'b1001 : 4'b1101;
										assign node2694 = (inp[9]) ? node2704 : node2695;
											assign node2695 = (inp[3]) ? node2697 : 4'b1100;
												assign node2697 = (inp[15]) ? node2701 : node2698;
													assign node2698 = (inp[12]) ? 4'b1100 : 4'b1110;
													assign node2701 = (inp[10]) ? 4'b1010 : 4'b1000;
											assign node2704 = (inp[12]) ? 4'b1100 : 4'b1010;
									assign node2707 = (inp[2]) ? node2719 : node2708;
										assign node2708 = (inp[4]) ? node2716 : node2709;
											assign node2709 = (inp[10]) ? node2713 : node2710;
												assign node2710 = (inp[9]) ? 4'b1000 : 4'b1100;
												assign node2713 = (inp[9]) ? 4'b1110 : 4'b1010;
											assign node2716 = (inp[15]) ? 4'b1100 : 4'b1000;
										assign node2719 = (inp[3]) ? node2731 : node2720;
											assign node2720 = (inp[4]) ? node2724 : node2721;
												assign node2721 = (inp[0]) ? 4'b0011 : 4'b0111;
												assign node2724 = (inp[10]) ? 4'b0001 : node2725;
													assign node2725 = (inp[12]) ? node2727 : 4'b0001;
														assign node2727 = (inp[0]) ? 4'b0101 : 4'b0111;
											assign node2731 = (inp[4]) ? node2733 : 4'b0001;
												assign node2733 = (inp[0]) ? 4'b0101 : 4'b0011;
								assign node2736 = (inp[0]) ? node2776 : node2737;
									assign node2737 = (inp[15]) ? node2757 : node2738;
										assign node2738 = (inp[9]) ? node2750 : node2739;
											assign node2739 = (inp[3]) ? node2745 : node2740;
												assign node2740 = (inp[8]) ? node2742 : 4'b0011;
													assign node2742 = (inp[2]) ? 4'b0011 : 4'b0010;
												assign node2745 = (inp[10]) ? node2747 : 4'b0001;
													assign node2747 = (inp[8]) ? 4'b0100 : 4'b0101;
											assign node2750 = (inp[4]) ? node2752 : 4'b0100;
												assign node2752 = (inp[8]) ? 4'b0101 : node2753;
													assign node2753 = (inp[2]) ? 4'b0000 : 4'b0001;
										assign node2757 = (inp[9]) ? node2763 : node2758;
											assign node2758 = (inp[12]) ? node2760 : 4'b0000;
												assign node2760 = (inp[8]) ? 4'b0011 : 4'b0010;
											assign node2763 = (inp[4]) ? node2773 : node2764;
												assign node2764 = (inp[12]) ? node2768 : node2765;
													assign node2765 = (inp[8]) ? 4'b0011 : 4'b0010;
													assign node2768 = (inp[10]) ? 4'b0111 : node2769;
														assign node2769 = (inp[2]) ? 4'b0110 : 4'b0110;
												assign node2773 = (inp[10]) ? 4'b0010 : 4'b0011;
									assign node2776 = (inp[15]) ? node2800 : node2777;
										assign node2777 = (inp[3]) ? node2791 : node2778;
											assign node2778 = (inp[4]) ? node2782 : node2779;
												assign node2779 = (inp[2]) ? 4'b0000 : 4'b0001;
												assign node2782 = (inp[8]) ? node2788 : node2783;
													assign node2783 = (inp[12]) ? 4'b0011 : node2784;
														assign node2784 = (inp[9]) ? 4'b0111 : 4'b0001;
													assign node2788 = (inp[2]) ? 4'b0111 : 4'b0110;
											assign node2791 = (inp[10]) ? node2793 : 4'b0110;
												assign node2793 = (inp[4]) ? node2795 : 4'b0110;
													assign node2795 = (inp[8]) ? 4'b0111 : node2796;
														assign node2796 = (inp[2]) ? 4'b0110 : 4'b0111;
										assign node2800 = (inp[8]) ? node2810 : node2801;
											assign node2801 = (inp[2]) ? 4'b0000 : node2802;
												assign node2802 = (inp[12]) ? 4'b0101 : node2803;
													assign node2803 = (inp[10]) ? 4'b0001 : node2804;
														assign node2804 = (inp[3]) ? 4'b0001 : 4'b0101;
											assign node2810 = (inp[2]) ? node2820 : node2811;
												assign node2811 = (inp[9]) ? node2817 : node2812;
													assign node2812 = (inp[4]) ? 4'b0100 : node2813;
														assign node2813 = (inp[12]) ? 4'b0010 : 4'b0000;
													assign node2817 = (inp[4]) ? 4'b0000 : 4'b0100;
												assign node2820 = (inp[9]) ? 4'b0101 : 4'b0001;
			assign node2823 = (inp[2]) ? node4255 : node2824;
				assign node2824 = (inp[8]) ? node3518 : node2825;
					assign node2825 = (inp[12]) ? node3155 : node2826;
						assign node2826 = (inp[11]) ? node2988 : node2827;
							assign node2827 = (inp[6]) ? node2893 : node2828;
								assign node2828 = (inp[13]) ? node2854 : node2829;
									assign node2829 = (inp[5]) ? node2839 : node2830;
										assign node2830 = (inp[0]) ? node2836 : node2831;
											assign node2831 = (inp[10]) ? node2833 : 4'b1110;
												assign node2833 = (inp[9]) ? 4'b1100 : 4'b1000;
											assign node2836 = (inp[15]) ? 4'b1010 : 4'b1000;
										assign node2839 = (inp[4]) ? node2849 : node2840;
											assign node2840 = (inp[9]) ? 4'b1010 : node2841;
												assign node2841 = (inp[15]) ? node2843 : 4'b1110;
													assign node2843 = (inp[10]) ? 4'b1100 : node2844;
														assign node2844 = (inp[1]) ? 4'b1100 : 4'b1110;
											assign node2849 = (inp[9]) ? node2851 : 4'b1000;
												assign node2851 = (inp[15]) ? 4'b1100 : 4'b1110;
									assign node2854 = (inp[1]) ? node2870 : node2855;
										assign node2855 = (inp[9]) ? node2863 : node2856;
											assign node2856 = (inp[4]) ? 4'b1010 : node2857;
												assign node2857 = (inp[3]) ? node2859 : 4'b1100;
													assign node2859 = (inp[10]) ? 4'b1100 : 4'b1110;
											assign node2863 = (inp[4]) ? 4'b1110 : node2864;
												assign node2864 = (inp[5]) ? 4'b1010 : node2865;
													assign node2865 = (inp[15]) ? 4'b1010 : 4'b1000;
										assign node2870 = (inp[5]) ? node2882 : node2871;
											assign node2871 = (inp[9]) ? node2879 : node2872;
												assign node2872 = (inp[4]) ? node2876 : node2873;
													assign node2873 = (inp[3]) ? 4'b0100 : 4'b0110;
													assign node2876 = (inp[10]) ? 4'b0000 : 4'b0010;
												assign node2879 = (inp[4]) ? 4'b0110 : 4'b0010;
											assign node2882 = (inp[10]) ? node2888 : node2883;
												assign node2883 = (inp[9]) ? 4'b0100 : node2884;
													assign node2884 = (inp[0]) ? 4'b0010 : 4'b0110;
												assign node2888 = (inp[15]) ? 4'b0000 : node2889;
													assign node2889 = (inp[4]) ? 4'b0110 : 4'b0000;
								assign node2893 = (inp[13]) ? node2943 : node2894;
									assign node2894 = (inp[3]) ? node2922 : node2895;
										assign node2895 = (inp[15]) ? node2913 : node2896;
											assign node2896 = (inp[10]) ? node2902 : node2897;
												assign node2897 = (inp[0]) ? node2899 : 4'b0100;
													assign node2899 = (inp[5]) ? 4'b0110 : 4'b0100;
												assign node2902 = (inp[0]) ? node2910 : node2903;
													assign node2903 = (inp[4]) ? node2907 : node2904;
														assign node2904 = (inp[9]) ? 4'b0010 : 4'b0110;
														assign node2907 = (inp[1]) ? 4'b0110 : 4'b0100;
													assign node2910 = (inp[5]) ? 4'b0110 : 4'b0100;
											assign node2913 = (inp[0]) ? node2917 : node2914;
												assign node2914 = (inp[4]) ? 4'b0110 : 4'b0100;
												assign node2917 = (inp[9]) ? node2919 : 4'b0110;
													assign node2919 = (inp[4]) ? 4'b0110 : 4'b0010;
										assign node2922 = (inp[10]) ? node2932 : node2923;
											assign node2923 = (inp[15]) ? node2925 : 4'b0110;
												assign node2925 = (inp[1]) ? 4'b0100 : node2926;
													assign node2926 = (inp[5]) ? 4'b0110 : node2927;
														assign node2927 = (inp[0]) ? 4'b0110 : 4'b0000;
											assign node2932 = (inp[9]) ? node2940 : node2933;
												assign node2933 = (inp[4]) ? node2937 : node2934;
													assign node2934 = (inp[15]) ? 4'b0100 : 4'b0110;
													assign node2937 = (inp[1]) ? 4'b0000 : 4'b0010;
												assign node2940 = (inp[1]) ? 4'b0100 : 4'b0000;
									assign node2943 = (inp[1]) ? node2967 : node2944;
										assign node2944 = (inp[4]) ? node2956 : node2945;
											assign node2945 = (inp[9]) ? node2951 : node2946;
												assign node2946 = (inp[5]) ? node2948 : 4'b0110;
													assign node2948 = (inp[3]) ? 4'b0110 : 4'b0100;
												assign node2951 = (inp[0]) ? 4'b0000 : node2952;
													assign node2952 = (inp[15]) ? 4'b0000 : 4'b0010;
											assign node2956 = (inp[9]) ? node2964 : node2957;
												assign node2957 = (inp[15]) ? 4'b0010 : node2958;
													assign node2958 = (inp[3]) ? node2960 : 4'b0010;
														assign node2960 = (inp[5]) ? 4'b0000 : 4'b0010;
												assign node2964 = (inp[3]) ? 4'b0100 : 4'b0110;
										assign node2967 = (inp[10]) ? node2979 : node2968;
											assign node2968 = (inp[9]) ? node2972 : node2969;
												assign node2969 = (inp[5]) ? 4'b1000 : 4'b1010;
												assign node2972 = (inp[4]) ? node2974 : 4'b1000;
													assign node2974 = (inp[0]) ? node2976 : 4'b1100;
														assign node2976 = (inp[15]) ? 4'b1100 : 4'b1110;
											assign node2979 = (inp[0]) ? node2983 : node2980;
												assign node2980 = (inp[4]) ? 4'b1000 : 4'b1010;
												assign node2983 = (inp[9]) ? 4'b1010 : node2984;
													assign node2984 = (inp[4]) ? 4'b1110 : 4'b1010;
							assign node2988 = (inp[6]) ? node3076 : node2989;
								assign node2989 = (inp[13]) ? node3031 : node2990;
									assign node2990 = (inp[3]) ? node3012 : node2991;
										assign node2991 = (inp[5]) ? node3007 : node2992;
											assign node2992 = (inp[9]) ? node3000 : node2993;
												assign node2993 = (inp[1]) ? 4'b0100 : node2994;
													assign node2994 = (inp[15]) ? node2996 : 4'b0000;
														assign node2996 = (inp[0]) ? 4'b0010 : 4'b0000;
												assign node3000 = (inp[4]) ? node3004 : node3001;
													assign node3001 = (inp[10]) ? 4'b0000 : 4'b0010;
													assign node3004 = (inp[10]) ? 4'b0110 : 4'b0100;
											assign node3007 = (inp[4]) ? 4'b0010 : node3008;
												assign node3008 = (inp[15]) ? 4'b0110 : 4'b0010;
										assign node3012 = (inp[5]) ? node3020 : node3013;
											assign node3013 = (inp[9]) ? node3017 : node3014;
												assign node3014 = (inp[4]) ? 4'b0010 : 4'b0110;
												assign node3017 = (inp[4]) ? 4'b0110 : 4'b0010;
											assign node3020 = (inp[15]) ? node3028 : node3021;
												assign node3021 = (inp[0]) ? node3023 : 4'b0100;
													assign node3023 = (inp[4]) ? node3025 : 4'b0110;
														assign node3025 = (inp[9]) ? 4'b0110 : 4'b0010;
												assign node3028 = (inp[4]) ? 4'b0000 : 4'b0100;
									assign node3031 = (inp[1]) ? node3049 : node3032;
										assign node3032 = (inp[3]) ? node3036 : node3033;
											assign node3033 = (inp[0]) ? 4'b0010 : 4'b0110;
											assign node3036 = (inp[10]) ? 4'b0100 : node3037;
												assign node3037 = (inp[9]) ? node3043 : node3038;
													assign node3038 = (inp[15]) ? node3040 : 4'b0100;
														assign node3040 = (inp[5]) ? 4'b0110 : 4'b0100;
													assign node3043 = (inp[5]) ? node3045 : 4'b0110;
														assign node3045 = (inp[15]) ? 4'b0100 : 4'b0100;
										assign node3049 = (inp[10]) ? node3067 : node3050;
											assign node3050 = (inp[3]) ? node3064 : node3051;
												assign node3051 = (inp[9]) ? node3059 : node3052;
													assign node3052 = (inp[4]) ? node3056 : node3053;
														assign node3053 = (inp[0]) ? 4'b1100 : 4'b1110;
														assign node3056 = (inp[0]) ? 4'b1000 : 4'b1010;
													assign node3059 = (inp[4]) ? 4'b1100 : node3060;
														assign node3060 = (inp[15]) ? 4'b1000 : 4'b1010;
												assign node3064 = (inp[9]) ? 4'b1110 : 4'b1100;
											assign node3067 = (inp[9]) ? node3073 : node3068;
												assign node3068 = (inp[4]) ? 4'b1110 : node3069;
													assign node3069 = (inp[0]) ? 4'b1000 : 4'b1010;
												assign node3073 = (inp[5]) ? 4'b1100 : 4'b1000;
								assign node3076 = (inp[1]) ? node3110 : node3077;
									assign node3077 = (inp[15]) ? node3091 : node3078;
										assign node3078 = (inp[9]) ? node3086 : node3079;
											assign node3079 = (inp[10]) ? node3083 : node3080;
												assign node3080 = (inp[0]) ? 4'b1100 : 4'b1010;
												assign node3083 = (inp[4]) ? 4'b1100 : 4'b1000;
											assign node3086 = (inp[10]) ? node3088 : 4'b1010;
												assign node3088 = (inp[3]) ? 4'b1100 : 4'b1000;
										assign node3091 = (inp[9]) ? node3101 : node3092;
											assign node3092 = (inp[0]) ? 4'b1010 : node3093;
												assign node3093 = (inp[5]) ? node3095 : 4'b1100;
													assign node3095 = (inp[13]) ? node3097 : 4'b1010;
														assign node3097 = (inp[10]) ? 4'b1010 : 4'b1110;
											assign node3101 = (inp[5]) ? 4'b1110 : node3102;
												assign node3102 = (inp[0]) ? node3104 : 4'b1010;
													assign node3104 = (inp[3]) ? 4'b1100 : node3105;
														assign node3105 = (inp[10]) ? 4'b1110 : 4'b1010;
									assign node3110 = (inp[13]) ? node3130 : node3111;
										assign node3111 = (inp[15]) ? node3123 : node3112;
											assign node3112 = (inp[0]) ? node3120 : node3113;
												assign node3113 = (inp[4]) ? node3115 : 4'b1100;
													assign node3115 = (inp[10]) ? node3117 : 4'b1100;
														assign node3117 = (inp[3]) ? 4'b1000 : 4'b1010;
												assign node3120 = (inp[3]) ? 4'b1110 : 4'b1100;
											assign node3123 = (inp[9]) ? node3125 : 4'b1000;
												assign node3125 = (inp[5]) ? 4'b1010 : node3126;
													assign node3126 = (inp[10]) ? 4'b1010 : 4'b1110;
										assign node3130 = (inp[4]) ? node3142 : node3131;
											assign node3131 = (inp[9]) ? node3137 : node3132;
												assign node3132 = (inp[15]) ? 4'b0000 : node3133;
													assign node3133 = (inp[5]) ? 4'b0000 : 4'b0010;
												assign node3137 = (inp[10]) ? 4'b0110 : node3138;
													assign node3138 = (inp[3]) ? 4'b0010 : 4'b0000;
											assign node3142 = (inp[9]) ? node3146 : node3143;
												assign node3143 = (inp[15]) ? 4'b0110 : 4'b0100;
												assign node3146 = (inp[10]) ? node3152 : node3147;
													assign node3147 = (inp[0]) ? 4'b0100 : node3148;
														assign node3148 = (inp[15]) ? 4'b0110 : 4'b0100;
													assign node3152 = (inp[5]) ? 4'b0010 : 4'b0000;
						assign node3155 = (inp[3]) ? node3367 : node3156;
							assign node3156 = (inp[6]) ? node3256 : node3157;
								assign node3157 = (inp[11]) ? node3207 : node3158;
									assign node3158 = (inp[1]) ? node3184 : node3159;
										assign node3159 = (inp[15]) ? node3173 : node3160;
											assign node3160 = (inp[0]) ? node3162 : 4'b1100;
												assign node3162 = (inp[4]) ? node3168 : node3163;
													assign node3163 = (inp[13]) ? node3165 : 4'b1000;
														assign node3165 = (inp[10]) ? 4'b1000 : 4'b1100;
													assign node3168 = (inp[5]) ? 4'b1110 : node3169;
														assign node3169 = (inp[9]) ? 4'b1000 : 4'b1100;
											assign node3173 = (inp[9]) ? node3181 : node3174;
												assign node3174 = (inp[0]) ? node3176 : 4'b1100;
													assign node3176 = (inp[4]) ? node3178 : 4'b1110;
														assign node3178 = (inp[10]) ? 4'b1110 : 4'b1010;
												assign node3181 = (inp[0]) ? 4'b1100 : 4'b1110;
										assign node3184 = (inp[13]) ? node3194 : node3185;
											assign node3185 = (inp[5]) ? 4'b1100 : node3186;
												assign node3186 = (inp[15]) ? node3190 : node3187;
													assign node3187 = (inp[0]) ? 4'b1000 : 4'b1010;
													assign node3190 = (inp[0]) ? 4'b1110 : 4'b1100;
											assign node3194 = (inp[15]) ? node3200 : node3195;
												assign node3195 = (inp[4]) ? node3197 : 4'b0010;
													assign node3197 = (inp[5]) ? 4'b0100 : 4'b0110;
												assign node3200 = (inp[0]) ? node3204 : node3201;
													assign node3201 = (inp[4]) ? 4'b0000 : 4'b0100;
													assign node3204 = (inp[5]) ? 4'b0100 : 4'b0110;
									assign node3207 = (inp[1]) ? node3235 : node3208;
										assign node3208 = (inp[9]) ? node3228 : node3209;
											assign node3209 = (inp[0]) ? node3221 : node3210;
												assign node3210 = (inp[15]) ? node3218 : node3211;
													assign node3211 = (inp[10]) ? node3215 : node3212;
														assign node3212 = (inp[4]) ? 4'b0010 : 4'b0110;
														assign node3215 = (inp[4]) ? 4'b0100 : 4'b0010;
													assign node3218 = (inp[5]) ? 4'b0110 : 4'b0100;
												assign node3221 = (inp[15]) ? 4'b0110 : node3222;
													assign node3222 = (inp[5]) ? 4'b0000 : node3223;
														assign node3223 = (inp[4]) ? 4'b0100 : 4'b0000;
											assign node3228 = (inp[4]) ? node3232 : node3229;
												assign node3229 = (inp[10]) ? 4'b0110 : 4'b0010;
												assign node3232 = (inp[10]) ? 4'b0010 : 4'b0110;
										assign node3235 = (inp[13]) ? node3245 : node3236;
											assign node3236 = (inp[4]) ? node3242 : node3237;
												assign node3237 = (inp[5]) ? node3239 : 4'b0100;
													assign node3239 = (inp[0]) ? 4'b0100 : 4'b0000;
												assign node3242 = (inp[5]) ? 4'b0100 : 4'b0110;
											assign node3245 = (inp[0]) ? node3251 : node3246;
												assign node3246 = (inp[10]) ? node3248 : 4'b1110;
													assign node3248 = (inp[5]) ? 4'b1110 : 4'b1100;
												assign node3251 = (inp[15]) ? 4'b1010 : node3252;
													assign node3252 = (inp[4]) ? 4'b1000 : 4'b1100;
								assign node3256 = (inp[11]) ? node3316 : node3257;
									assign node3257 = (inp[1]) ? node3293 : node3258;
										assign node3258 = (inp[13]) ? node3274 : node3259;
											assign node3259 = (inp[10]) ? node3265 : node3260;
												assign node3260 = (inp[15]) ? 4'b0000 : node3261;
													assign node3261 = (inp[0]) ? 4'b0000 : 4'b0110;
												assign node3265 = (inp[15]) ? node3269 : node3266;
													assign node3266 = (inp[9]) ? 4'b0100 : 4'b0000;
													assign node3269 = (inp[5]) ? node3271 : 4'b0110;
														assign node3271 = (inp[0]) ? 4'b0100 : 4'b0110;
											assign node3274 = (inp[5]) ? node3278 : node3275;
												assign node3275 = (inp[10]) ? 4'b0010 : 4'b0110;
												assign node3278 = (inp[4]) ? node3286 : node3279;
													assign node3279 = (inp[9]) ? node3283 : node3280;
														assign node3280 = (inp[10]) ? 4'b0010 : 4'b0110;
														assign node3283 = (inp[0]) ? 4'b0100 : 4'b0100;
													assign node3286 = (inp[0]) ? node3290 : node3287;
														assign node3287 = (inp[10]) ? 4'b0000 : 4'b0100;
														assign node3290 = (inp[10]) ? 4'b0010 : 4'b0000;
										assign node3293 = (inp[13]) ? node3301 : node3294;
											assign node3294 = (inp[10]) ? 4'b0110 : node3295;
												assign node3295 = (inp[4]) ? node3297 : 4'b0000;
													assign node3297 = (inp[5]) ? 4'b0010 : 4'b0110;
											assign node3301 = (inp[4]) ? node3309 : node3302;
												assign node3302 = (inp[9]) ? 4'b1110 : node3303;
													assign node3303 = (inp[0]) ? 4'b1010 : node3304;
														assign node3304 = (inp[15]) ? 4'b1000 : 4'b1010;
												assign node3309 = (inp[9]) ? 4'b1000 : node3310;
													assign node3310 = (inp[10]) ? node3312 : 4'b1100;
														assign node3312 = (inp[0]) ? 4'b1110 : 4'b1100;
									assign node3316 = (inp[1]) ? node3338 : node3317;
										assign node3317 = (inp[13]) ? node3323 : node3318;
											assign node3318 = (inp[0]) ? 4'b1000 : node3319;
												assign node3319 = (inp[4]) ? 4'b1000 : 4'b1100;
											assign node3323 = (inp[0]) ? node3327 : node3324;
												assign node3324 = (inp[10]) ? 4'b1100 : 4'b1000;
												assign node3327 = (inp[5]) ? node3333 : node3328;
													assign node3328 = (inp[15]) ? node3330 : 4'b1100;
														assign node3330 = (inp[9]) ? 4'b1110 : 4'b1010;
													assign node3333 = (inp[15]) ? node3335 : 4'b1010;
														assign node3335 = (inp[10]) ? 4'b1100 : 4'b1000;
										assign node3338 = (inp[13]) ? node3346 : node3339;
											assign node3339 = (inp[5]) ? node3341 : 4'b1000;
												assign node3341 = (inp[4]) ? node3343 : 4'b1110;
													assign node3343 = (inp[15]) ? 4'b1010 : 4'b1000;
											assign node3346 = (inp[0]) ? node3358 : node3347;
												assign node3347 = (inp[5]) ? node3353 : node3348;
													assign node3348 = (inp[15]) ? node3350 : 4'b0110;
														assign node3350 = (inp[10]) ? 4'b0100 : 4'b0000;
													assign node3353 = (inp[4]) ? 4'b0000 : node3354;
														assign node3354 = (inp[15]) ? 4'b0000 : 4'b0010;
												assign node3358 = (inp[15]) ? node3364 : node3359;
													assign node3359 = (inp[9]) ? node3361 : 4'b0000;
														assign node3361 = (inp[4]) ? 4'b0010 : 4'b0110;
													assign node3364 = (inp[4]) ? 4'b0110 : 4'b0100;
							assign node3367 = (inp[1]) ? node3435 : node3368;
								assign node3368 = (inp[9]) ? node3404 : node3369;
									assign node3369 = (inp[5]) ? node3387 : node3370;
										assign node3370 = (inp[6]) ? node3380 : node3371;
											assign node3371 = (inp[4]) ? 4'b0010 : node3372;
												assign node3372 = (inp[10]) ? node3376 : node3373;
													assign node3373 = (inp[15]) ? 4'b0110 : 4'b0100;
													assign node3376 = (inp[0]) ? 4'b0010 : 4'b0000;
											assign node3380 = (inp[13]) ? node3384 : node3381;
												assign node3381 = (inp[0]) ? 4'b0000 : 4'b0100;
												assign node3384 = (inp[4]) ? 4'b1100 : 4'b1000;
										assign node3387 = (inp[13]) ? node3401 : node3388;
											assign node3388 = (inp[0]) ? node3394 : node3389;
												assign node3389 = (inp[4]) ? 4'b1110 : node3390;
													assign node3390 = (inp[15]) ? 4'b1010 : 4'b1000;
												assign node3394 = (inp[4]) ? node3398 : node3395;
													assign node3395 = (inp[11]) ? 4'b1000 : 4'b0000;
													assign node3398 = (inp[10]) ? 4'b1100 : 4'b1000;
											assign node3401 = (inp[0]) ? 4'b1100 : 4'b0100;
									assign node3404 = (inp[15]) ? node3420 : node3405;
										assign node3405 = (inp[0]) ? node3407 : 4'b0000;
											assign node3407 = (inp[10]) ? node3415 : node3408;
												assign node3408 = (inp[11]) ? node3412 : node3409;
													assign node3409 = (inp[6]) ? 4'b0110 : 4'b1110;
													assign node3412 = (inp[4]) ? 4'b1010 : 4'b0010;
												assign node3415 = (inp[5]) ? node3417 : 4'b0010;
													assign node3417 = (inp[6]) ? 4'b1010 : 4'b0010;
										assign node3420 = (inp[0]) ? node3428 : node3421;
											assign node3421 = (inp[6]) ? 4'b1110 : node3422;
												assign node3422 = (inp[4]) ? node3424 : 4'b1000;
													assign node3424 = (inp[11]) ? 4'b0010 : 4'b1010;
											assign node3428 = (inp[4]) ? node3432 : node3429;
												assign node3429 = (inp[6]) ? 4'b1100 : 4'b0010;
												assign node3432 = (inp[10]) ? 4'b0000 : 4'b0100;
								assign node3435 = (inp[9]) ? node3475 : node3436;
									assign node3436 = (inp[4]) ? node3458 : node3437;
										assign node3437 = (inp[11]) ? node3449 : node3438;
											assign node3438 = (inp[10]) ? 4'b1010 : node3439;
												assign node3439 = (inp[0]) ? node3445 : node3440;
													assign node3440 = (inp[5]) ? node3442 : 4'b0110;
														assign node3442 = (inp[6]) ? 4'b0100 : 4'b0110;
													assign node3445 = (inp[5]) ? 4'b1010 : 4'b0110;
											assign node3449 = (inp[15]) ? node3451 : 4'b0100;
												assign node3451 = (inp[6]) ? node3455 : node3452;
													assign node3452 = (inp[13]) ? 4'b1000 : 4'b0000;
													assign node3455 = (inp[5]) ? 4'b0000 : 4'b0010;
										assign node3458 = (inp[13]) ? node3468 : node3459;
											assign node3459 = (inp[10]) ? node3463 : node3460;
												assign node3460 = (inp[5]) ? 4'b0010 : 4'b0000;
												assign node3463 = (inp[5]) ? node3465 : 4'b1110;
													assign node3465 = (inp[11]) ? 4'b1110 : 4'b0110;
											assign node3468 = (inp[6]) ? node3472 : node3469;
												assign node3469 = (inp[11]) ? 4'b1110 : 4'b0110;
												assign node3472 = (inp[11]) ? 4'b0100 : 4'b1100;
									assign node3475 = (inp[4]) ? node3499 : node3476;
										assign node3476 = (inp[11]) ? node3488 : node3477;
											assign node3477 = (inp[5]) ? node3479 : 4'b0100;
												assign node3479 = (inp[15]) ? node3483 : node3480;
													assign node3480 = (inp[10]) ? 4'b1100 : 4'b1000;
													assign node3483 = (inp[13]) ? 4'b1110 : node3484;
														assign node3484 = (inp[10]) ? 4'b0110 : 4'b0010;
											assign node3488 = (inp[0]) ? node3492 : node3489;
												assign node3489 = (inp[15]) ? 4'b1110 : 4'b1100;
												assign node3492 = (inp[5]) ? 4'b1110 : node3493;
													assign node3493 = (inp[13]) ? node3495 : 4'b1110;
														assign node3495 = (inp[6]) ? 4'b0110 : 4'b1110;
										assign node3499 = (inp[10]) ? node3509 : node3500;
											assign node3500 = (inp[13]) ? node3506 : node3501;
												assign node3501 = (inp[15]) ? node3503 : 4'b0100;
													assign node3503 = (inp[5]) ? 4'b1110 : 4'b0110;
												assign node3506 = (inp[11]) ? 4'b0010 : 4'b1010;
											assign node3509 = (inp[11]) ? node3511 : 4'b1010;
												assign node3511 = (inp[15]) ? node3515 : node3512;
													assign node3512 = (inp[0]) ? 4'b1010 : 4'b1000;
													assign node3515 = (inp[13]) ? 4'b1000 : 4'b0000;
					assign node3518 = (inp[12]) ? node3898 : node3519;
						assign node3519 = (inp[0]) ? node3705 : node3520;
							assign node3520 = (inp[9]) ? node3610 : node3521;
								assign node3521 = (inp[4]) ? node3567 : node3522;
									assign node3522 = (inp[10]) ? node3546 : node3523;
										assign node3523 = (inp[15]) ? node3533 : node3524;
											assign node3524 = (inp[5]) ? node3528 : node3525;
												assign node3525 = (inp[13]) ? 4'b0111 : 4'b1111;
												assign node3528 = (inp[3]) ? node3530 : 4'b0111;
													assign node3530 = (inp[13]) ? 4'b1101 : 4'b0101;
											assign node3533 = (inp[13]) ? node3541 : node3534;
												assign node3534 = (inp[6]) ? 4'b0101 : node3535;
													assign node3535 = (inp[11]) ? node3537 : 4'b1101;
														assign node3537 = (inp[1]) ? 4'b1111 : 4'b0111;
												assign node3541 = (inp[1]) ? 4'b1101 : node3542;
													assign node3542 = (inp[6]) ? 4'b1101 : 4'b1111;
										assign node3546 = (inp[13]) ? node3562 : node3547;
											assign node3547 = (inp[11]) ? node3557 : node3548;
												assign node3548 = (inp[1]) ? node3552 : node3549;
													assign node3549 = (inp[3]) ? 4'b1101 : 4'b1111;
													assign node3552 = (inp[3]) ? 4'b0101 : node3553;
														assign node3553 = (inp[15]) ? 4'b0101 : 4'b0111;
												assign node3557 = (inp[3]) ? node3559 : 4'b0011;
													assign node3559 = (inp[15]) ? 4'b1001 : 4'b1011;
											assign node3562 = (inp[11]) ? 4'b1001 : node3563;
												assign node3563 = (inp[3]) ? 4'b1001 : 4'b1011;
									assign node3567 = (inp[10]) ? node3595 : node3568;
										assign node3568 = (inp[5]) ? node3578 : node3569;
											assign node3569 = (inp[15]) ? node3571 : 4'b1011;
												assign node3571 = (inp[1]) ? 4'b1001 : node3572;
													assign node3572 = (inp[3]) ? node3574 : 4'b0001;
														assign node3574 = (inp[11]) ? 4'b0001 : 4'b0001;
											assign node3578 = (inp[15]) ? node3586 : node3579;
												assign node3579 = (inp[3]) ? node3581 : 4'b0011;
													assign node3581 = (inp[1]) ? 4'b1001 : node3582;
														assign node3582 = (inp[11]) ? 4'b0001 : 4'b0001;
												assign node3586 = (inp[3]) ? node3590 : node3587;
													assign node3587 = (inp[13]) ? 4'b1001 : 4'b0001;
													assign node3590 = (inp[13]) ? 4'b0011 : node3591;
														assign node3591 = (inp[1]) ? 4'b0011 : 4'b1011;
										assign node3595 = (inp[15]) ? node3601 : node3596;
											assign node3596 = (inp[5]) ? 4'b1101 : node3597;
												assign node3597 = (inp[3]) ? 4'b1101 : 4'b1111;
											assign node3601 = (inp[1]) ? node3607 : node3602;
												assign node3602 = (inp[11]) ? node3604 : 4'b0001;
													assign node3604 = (inp[6]) ? 4'b1101 : 4'b0001;
												assign node3607 = (inp[3]) ? 4'b0111 : 4'b0101;
								assign node3610 = (inp[4]) ? node3640 : node3611;
									assign node3611 = (inp[10]) ? node3625 : node3612;
										assign node3612 = (inp[15]) ? node3618 : node3613;
											assign node3613 = (inp[5]) ? node3615 : 4'b1011;
												assign node3615 = (inp[6]) ? 4'b1001 : 4'b0011;
											assign node3618 = (inp[13]) ? node3622 : node3619;
												assign node3619 = (inp[6]) ? 4'b0001 : 4'b1001;
												assign node3622 = (inp[1]) ? 4'b0001 : 4'b0011;
										assign node3625 = (inp[6]) ? node3635 : node3626;
											assign node3626 = (inp[3]) ? 4'b0001 : node3627;
												assign node3627 = (inp[11]) ? 4'b1111 : node3628;
													assign node3628 = (inp[15]) ? 4'b0001 : node3629;
														assign node3629 = (inp[1]) ? 4'b0011 : 4'b1011;
											assign node3635 = (inp[11]) ? node3637 : 4'b1101;
												assign node3637 = (inp[15]) ? 4'b0111 : 4'b0101;
									assign node3640 = (inp[15]) ? node3674 : node3641;
										assign node3641 = (inp[10]) ? node3655 : node3642;
											assign node3642 = (inp[6]) ? node3644 : 4'b0101;
												assign node3644 = (inp[11]) ? node3648 : node3645;
													assign node3645 = (inp[1]) ? 4'b1101 : 4'b0101;
													assign node3648 = (inp[5]) ? node3652 : node3649;
														assign node3649 = (inp[3]) ? 4'b0101 : 4'b0111;
														assign node3652 = (inp[13]) ? 4'b0101 : 4'b1101;
											assign node3655 = (inp[6]) ? node3663 : node3656;
												assign node3656 = (inp[5]) ? node3658 : 4'b0101;
													assign node3658 = (inp[13]) ? 4'b1001 : node3659;
														assign node3659 = (inp[1]) ? 4'b0101 : 4'b1101;
												assign node3663 = (inp[3]) ? node3669 : node3664;
													assign node3664 = (inp[13]) ? 4'b0011 : node3665;
														assign node3665 = (inp[1]) ? 4'b1011 : 4'b0011;
													assign node3669 = (inp[1]) ? 4'b1001 : node3670;
														assign node3670 = (inp[5]) ? 4'b0001 : 4'b0101;
										assign node3674 = (inp[3]) ? node3690 : node3675;
											assign node3675 = (inp[5]) ? node3683 : node3676;
												assign node3676 = (inp[10]) ? node3680 : node3677;
													assign node3677 = (inp[11]) ? 4'b1101 : 4'b0101;
													assign node3680 = (inp[13]) ? 4'b1001 : 4'b0001;
												assign node3683 = (inp[13]) ? node3687 : node3684;
													assign node3684 = (inp[11]) ? 4'b1011 : 4'b1111;
													assign node3687 = (inp[10]) ? 4'b0011 : 4'b0111;
											assign node3690 = (inp[10]) ? node3702 : node3691;
												assign node3691 = (inp[6]) ? node3697 : node3692;
													assign node3692 = (inp[11]) ? node3694 : 4'b0111;
														assign node3694 = (inp[13]) ? 4'b1111 : 4'b0111;
													assign node3697 = (inp[11]) ? node3699 : 4'b1111;
														assign node3699 = (inp[13]) ? 4'b0111 : 4'b1111;
												assign node3702 = (inp[6]) ? 4'b0011 : 4'b0111;
							assign node3705 = (inp[15]) ? node3801 : node3706;
								assign node3706 = (inp[3]) ? node3752 : node3707;
									assign node3707 = (inp[5]) ? node3737 : node3708;
										assign node3708 = (inp[9]) ? node3720 : node3709;
											assign node3709 = (inp[10]) ? node3711 : 4'b0101;
												assign node3711 = (inp[1]) ? node3715 : node3712;
													assign node3712 = (inp[11]) ? 4'b0101 : 4'b0001;
													assign node3715 = (inp[13]) ? 4'b0001 : node3716;
														assign node3716 = (inp[6]) ? 4'b1101 : 4'b1001;
											assign node3720 = (inp[4]) ? node3728 : node3721;
												assign node3721 = (inp[6]) ? 4'b0101 : node3722;
													assign node3722 = (inp[1]) ? node3724 : 4'b1001;
														assign node3724 = (inp[11]) ? 4'b1001 : 4'b0001;
												assign node3728 = (inp[6]) ? node3734 : node3729;
													assign node3729 = (inp[10]) ? node3731 : 4'b1101;
														assign node3731 = (inp[1]) ? 4'b0101 : 4'b0101;
													assign node3734 = (inp[1]) ? 4'b1001 : 4'b1101;
										assign node3737 = (inp[10]) ? node3747 : node3738;
											assign node3738 = (inp[1]) ? 4'b0001 : node3739;
												assign node3739 = (inp[13]) ? node3743 : node3740;
													assign node3740 = (inp[11]) ? 4'b0001 : 4'b1001;
													assign node3743 = (inp[11]) ? 4'b1101 : 4'b1001;
											assign node3747 = (inp[11]) ? node3749 : 4'b0001;
												assign node3749 = (inp[4]) ? 4'b0111 : 4'b1111;
									assign node3752 = (inp[5]) ? node3782 : node3753;
										assign node3753 = (inp[4]) ? node3769 : node3754;
											assign node3754 = (inp[1]) ? node3764 : node3755;
												assign node3755 = (inp[9]) ? node3761 : node3756;
													assign node3756 = (inp[11]) ? node3758 : 4'b0101;
														assign node3758 = (inp[13]) ? 4'b1101 : 4'b0101;
													assign node3761 = (inp[11]) ? 4'b0001 : 4'b1001;
												assign node3764 = (inp[11]) ? node3766 : 4'b1001;
													assign node3766 = (inp[6]) ? 4'b0001 : 4'b1001;
											assign node3769 = (inp[6]) ? node3777 : node3770;
												assign node3770 = (inp[9]) ? node3774 : node3771;
													assign node3771 = (inp[1]) ? 4'b1001 : 4'b0001;
													assign node3774 = (inp[10]) ? 4'b1011 : 4'b1111;
												assign node3777 = (inp[11]) ? node3779 : 4'b1111;
													assign node3779 = (inp[1]) ? 4'b0111 : 4'b1111;
										assign node3782 = (inp[11]) ? node3796 : node3783;
											assign node3783 = (inp[6]) ? node3789 : node3784;
												assign node3784 = (inp[10]) ? node3786 : 4'b0111;
													assign node3786 = (inp[13]) ? 4'b0011 : 4'b1011;
												assign node3789 = (inp[1]) ? node3791 : 4'b0011;
													assign node3791 = (inp[9]) ? 4'b1011 : node3792;
														assign node3792 = (inp[4]) ? 4'b1111 : 4'b1011;
											assign node3796 = (inp[10]) ? 4'b1111 : node3797;
												assign node3797 = (inp[9]) ? 4'b1011 : 4'b1111;
								assign node3801 = (inp[3]) ? node3851 : node3802;
									assign node3802 = (inp[9]) ? node3822 : node3803;
										assign node3803 = (inp[11]) ? node3813 : node3804;
											assign node3804 = (inp[13]) ? node3808 : node3805;
												assign node3805 = (inp[5]) ? 4'b0111 : 4'b1111;
												assign node3808 = (inp[6]) ? 4'b1111 : node3809;
													assign node3809 = (inp[4]) ? 4'b0011 : 4'b0111;
											assign node3813 = (inp[13]) ? node3819 : node3814;
												assign node3814 = (inp[6]) ? 4'b1011 : node3815;
													assign node3815 = (inp[1]) ? 4'b1011 : 4'b0011;
												assign node3819 = (inp[10]) ? 4'b1111 : 4'b1011;
										assign node3822 = (inp[5]) ? node3836 : node3823;
											assign node3823 = (inp[4]) ? node3831 : node3824;
												assign node3824 = (inp[13]) ? node3828 : node3825;
													assign node3825 = (inp[10]) ? 4'b1111 : 4'b1011;
													assign node3828 = (inp[1]) ? 4'b0111 : 4'b0011;
												assign node3831 = (inp[10]) ? node3833 : 4'b0111;
													assign node3833 = (inp[6]) ? 4'b0011 : 4'b0111;
											assign node3836 = (inp[4]) ? node3844 : node3837;
												assign node3837 = (inp[6]) ? node3839 : 4'b0011;
													assign node3839 = (inp[10]) ? node3841 : 4'b0011;
														assign node3841 = (inp[1]) ? 4'b0101 : 4'b1101;
												assign node3844 = (inp[10]) ? node3846 : 4'b0101;
													assign node3846 = (inp[1]) ? 4'b0101 : node3847;
														assign node3847 = (inp[6]) ? 4'b0001 : 4'b1001;
									assign node3851 = (inp[5]) ? node3871 : node3852;
										assign node3852 = (inp[9]) ? node3858 : node3853;
											assign node3853 = (inp[4]) ? 4'b0011 : node3854;
												assign node3854 = (inp[10]) ? 4'b1011 : 4'b1111;
											assign node3858 = (inp[11]) ? node3864 : node3859;
												assign node3859 = (inp[1]) ? 4'b1001 : node3860;
													assign node3860 = (inp[13]) ? 4'b0011 : 4'b1011;
												assign node3864 = (inp[13]) ? node3866 : 4'b1101;
													assign node3866 = (inp[6]) ? node3868 : 4'b1001;
														assign node3868 = (inp[10]) ? 4'b0001 : 4'b0101;
										assign node3871 = (inp[1]) ? node3887 : node3872;
											assign node3872 = (inp[9]) ? node3878 : node3873;
												assign node3873 = (inp[11]) ? node3875 : 4'b1001;
													assign node3875 = (inp[10]) ? 4'b1001 : 4'b0001;
												assign node3878 = (inp[4]) ? node3880 : 4'b0001;
													assign node3880 = (inp[10]) ? node3884 : node3881;
														assign node3881 = (inp[11]) ? 4'b0101 : 4'b0101;
														assign node3884 = (inp[13]) ? 4'b1001 : 4'b1101;
											assign node3887 = (inp[4]) ? node3893 : node3888;
												assign node3888 = (inp[11]) ? 4'b1101 : node3889;
													assign node3889 = (inp[9]) ? 4'b0001 : 4'b0101;
												assign node3893 = (inp[11]) ? node3895 : 4'b0101;
													assign node3895 = (inp[10]) ? 4'b0001 : 4'b0101;
						assign node3898 = (inp[11]) ? node4070 : node3899;
							assign node3899 = (inp[6]) ? node3981 : node3900;
								assign node3900 = (inp[1]) ? node3948 : node3901;
									assign node3901 = (inp[13]) ? node3927 : node3902;
										assign node3902 = (inp[10]) ? node3920 : node3903;
											assign node3903 = (inp[4]) ? node3911 : node3904;
												assign node3904 = (inp[9]) ? node3908 : node3905;
													assign node3905 = (inp[0]) ? 4'b1111 : 4'b1101;
													assign node3908 = (inp[15]) ? 4'b1001 : 4'b1011;
												assign node3911 = (inp[9]) ? node3917 : node3912;
													assign node3912 = (inp[0]) ? node3914 : 4'b1001;
														assign node3914 = (inp[15]) ? 4'b1011 : 4'b1001;
													assign node3917 = (inp[3]) ? 4'b1101 : 4'b1111;
											assign node3920 = (inp[0]) ? node3924 : node3921;
												assign node3921 = (inp[3]) ? 4'b1001 : 4'b1111;
												assign node3924 = (inp[3]) ? 4'b1101 : 4'b1001;
										assign node3927 = (inp[9]) ? node3939 : node3928;
											assign node3928 = (inp[4]) ? node3934 : node3929;
												assign node3929 = (inp[0]) ? node3931 : 4'b0101;
													assign node3931 = (inp[15]) ? 4'b0111 : 4'b0101;
												assign node3934 = (inp[10]) ? 4'b0101 : node3935;
													assign node3935 = (inp[3]) ? 4'b0011 : 4'b0001;
											assign node3939 = (inp[0]) ? node3945 : node3940;
												assign node3940 = (inp[5]) ? 4'b0011 : node3941;
													assign node3941 = (inp[10]) ? 4'b0111 : 4'b0011;
												assign node3945 = (inp[15]) ? 4'b0001 : 4'b0011;
									assign node3948 = (inp[0]) ? node3964 : node3949;
										assign node3949 = (inp[15]) ? node3959 : node3950;
											assign node3950 = (inp[5]) ? node3952 : 4'b0011;
												assign node3952 = (inp[4]) ? 4'b0001 : node3953;
													assign node3953 = (inp[13]) ? 4'b0011 : node3954;
														assign node3954 = (inp[9]) ? 4'b0101 : 4'b0011;
											assign node3959 = (inp[5]) ? node3961 : 4'b0001;
												assign node3961 = (inp[13]) ? 4'b0011 : 4'b0111;
										assign node3964 = (inp[4]) ? node3976 : node3965;
											assign node3965 = (inp[9]) ? node3969 : node3966;
												assign node3966 = (inp[15]) ? 4'b0011 : 4'b0111;
												assign node3969 = (inp[13]) ? node3971 : 4'b0111;
													assign node3971 = (inp[15]) ? 4'b0101 : node3972;
														assign node3972 = (inp[3]) ? 4'b0111 : 4'b0101;
											assign node3976 = (inp[9]) ? 4'b0011 : node3977;
												assign node3977 = (inp[10]) ? 4'b0101 : 4'b0001;
								assign node3981 = (inp[1]) ? node4023 : node3982;
									assign node3982 = (inp[13]) ? node4010 : node3983;
										assign node3983 = (inp[3]) ? node3997 : node3984;
											assign node3984 = (inp[4]) ? node3994 : node3985;
												assign node3985 = (inp[10]) ? node3989 : node3986;
													assign node3986 = (inp[9]) ? 4'b0011 : 4'b0111;
													assign node3989 = (inp[15]) ? 4'b0101 : node3990;
														assign node3990 = (inp[0]) ? 4'b0001 : 4'b0011;
												assign node3994 = (inp[15]) ? 4'b0001 : 4'b0101;
											assign node3997 = (inp[5]) ? 4'b0011 : node3998;
												assign node3998 = (inp[4]) ? node4004 : node3999;
													assign node3999 = (inp[10]) ? 4'b0101 : node4000;
														assign node4000 = (inp[15]) ? 4'b0001 : 4'b0001;
													assign node4004 = (inp[10]) ? 4'b0011 : node4005;
														assign node4005 = (inp[0]) ? 4'b0011 : 4'b0001;
										assign node4010 = (inp[4]) ? node4016 : node4011;
											assign node4011 = (inp[9]) ? node4013 : 4'b1011;
												assign node4013 = (inp[10]) ? 4'b1111 : 4'b1101;
											assign node4016 = (inp[9]) ? node4018 : 4'b1101;
												assign node4018 = (inp[5]) ? node4020 : 4'b1001;
													assign node4020 = (inp[15]) ? 4'b1001 : 4'b1011;
									assign node4023 = (inp[5]) ? node4049 : node4024;
										assign node4024 = (inp[10]) ? node4034 : node4025;
											assign node4025 = (inp[13]) ? node4031 : node4026;
												assign node4026 = (inp[3]) ? node4028 : 4'b1011;
													assign node4028 = (inp[4]) ? 4'b1111 : 4'b1011;
												assign node4031 = (inp[0]) ? 4'b1001 : 4'b1011;
											assign node4034 = (inp[15]) ? node4040 : node4035;
												assign node4035 = (inp[9]) ? node4037 : 4'b1001;
													assign node4037 = (inp[0]) ? 4'b1011 : 4'b1001;
												assign node4040 = (inp[3]) ? node4044 : node4041;
													assign node4041 = (inp[13]) ? 4'b1001 : 4'b1011;
													assign node4044 = (inp[0]) ? node4046 : 4'b1111;
														assign node4046 = (inp[4]) ? 4'b1001 : 4'b1101;
										assign node4049 = (inp[10]) ? node4061 : node4050;
											assign node4050 = (inp[3]) ? node4056 : node4051;
												assign node4051 = (inp[13]) ? node4053 : 4'b1101;
													assign node4053 = (inp[9]) ? 4'b1011 : 4'b1111;
												assign node4056 = (inp[15]) ? 4'b1101 : node4057;
													assign node4057 = (inp[0]) ? 4'b1011 : 4'b1001;
											assign node4061 = (inp[15]) ? node4065 : node4062;
												assign node4062 = (inp[0]) ? 4'b1111 : 4'b1101;
												assign node4065 = (inp[0]) ? 4'b1101 : node4066;
													assign node4066 = (inp[3]) ? 4'b1111 : 4'b1001;
							assign node4070 = (inp[6]) ? node4154 : node4071;
								assign node4071 = (inp[1]) ? node4119 : node4072;
									assign node4072 = (inp[13]) ? node4106 : node4073;
										assign node4073 = (inp[4]) ? node4083 : node4074;
											assign node4074 = (inp[3]) ? node4078 : node4075;
												assign node4075 = (inp[0]) ? 4'b0001 : 4'b0011;
												assign node4078 = (inp[10]) ? 4'b0011 : node4079;
													assign node4079 = (inp[15]) ? 4'b0111 : 4'b0011;
											assign node4083 = (inp[5]) ? node4097 : node4084;
												assign node4084 = (inp[3]) ? node4092 : node4085;
													assign node4085 = (inp[0]) ? node4089 : node4086;
														assign node4086 = (inp[9]) ? 4'b0001 : 4'b0011;
														assign node4089 = (inp[9]) ? 4'b0011 : 4'b0111;
													assign node4092 = (inp[9]) ? node4094 : 4'b0111;
														assign node4094 = (inp[15]) ? 4'b0111 : 4'b0101;
												assign node4097 = (inp[10]) ? node4103 : node4098;
													assign node4098 = (inp[15]) ? node4100 : 4'b0011;
														assign node4100 = (inp[9]) ? 4'b0101 : 4'b0001;
													assign node4103 = (inp[0]) ? 4'b0101 : 4'b0111;
										assign node4106 = (inp[0]) ? node4114 : node4107;
											assign node4107 = (inp[15]) ? node4111 : node4108;
												assign node4108 = (inp[9]) ? 4'b1001 : 4'b1101;
												assign node4111 = (inp[4]) ? 4'b1011 : 4'b1001;
											assign node4114 = (inp[4]) ? node4116 : 4'b1111;
												assign node4116 = (inp[5]) ? 4'b1111 : 4'b1011;
									assign node4119 = (inp[9]) ? node4139 : node4120;
										assign node4120 = (inp[4]) ? node4126 : node4121;
											assign node4121 = (inp[15]) ? 4'b1001 : node4122;
												assign node4122 = (inp[13]) ? 4'b1001 : 4'b1011;
											assign node4126 = (inp[10]) ? node4134 : node4127;
												assign node4127 = (inp[15]) ? 4'b1101 : node4128;
													assign node4128 = (inp[13]) ? 4'b1111 : node4129;
														assign node4129 = (inp[0]) ? 4'b1111 : 4'b1101;
												assign node4134 = (inp[0]) ? 4'b1111 : node4135;
													assign node4135 = (inp[3]) ? 4'b1111 : 4'b1101;
										assign node4139 = (inp[4]) ? node4145 : node4140;
											assign node4140 = (inp[13]) ? node4142 : 4'b1111;
												assign node4142 = (inp[10]) ? 4'b1111 : 4'b1101;
											assign node4145 = (inp[5]) ? 4'b1011 : node4146;
												assign node4146 = (inp[0]) ? 4'b1011 : node4147;
													assign node4147 = (inp[10]) ? 4'b1011 : node4148;
														assign node4148 = (inp[3]) ? 4'b1001 : 4'b1001;
								assign node4154 = (inp[13]) ? node4198 : node4155;
									assign node4155 = (inp[1]) ? node4177 : node4156;
										assign node4156 = (inp[0]) ? node4166 : node4157;
											assign node4157 = (inp[15]) ? node4161 : node4158;
												assign node4158 = (inp[5]) ? 4'b1101 : 4'b1011;
												assign node4161 = (inp[9]) ? node4163 : 4'b1001;
													assign node4163 = (inp[3]) ? 4'b1011 : 4'b1001;
											assign node4166 = (inp[5]) ? 4'b1111 : node4167;
												assign node4167 = (inp[3]) ? node4171 : node4168;
													assign node4168 = (inp[15]) ? 4'b1111 : 4'b1101;
													assign node4171 = (inp[10]) ? 4'b1001 : node4172;
														assign node4172 = (inp[4]) ? 4'b1011 : 4'b1111;
										assign node4177 = (inp[5]) ? node4193 : node4178;
											assign node4178 = (inp[3]) ? node4186 : node4179;
												assign node4179 = (inp[15]) ? node4183 : node4180;
													assign node4180 = (inp[4]) ? 4'b0001 : 4'b0101;
													assign node4183 = (inp[10]) ? 4'b0011 : 4'b0111;
												assign node4186 = (inp[15]) ? node4190 : node4187;
													assign node4187 = (inp[0]) ? 4'b0111 : 4'b0101;
													assign node4190 = (inp[10]) ? 4'b0111 : 4'b0101;
											assign node4193 = (inp[0]) ? node4195 : 4'b0101;
												assign node4195 = (inp[3]) ? 4'b0001 : 4'b0011;
									assign node4198 = (inp[0]) ? node4224 : node4199;
										assign node4199 = (inp[10]) ? node4217 : node4200;
											assign node4200 = (inp[5]) ? node4212 : node4201;
												assign node4201 = (inp[15]) ? node4207 : node4202;
													assign node4202 = (inp[3]) ? node4204 : 4'b0111;
														assign node4204 = (inp[4]) ? 4'b0001 : 4'b0011;
													assign node4207 = (inp[1]) ? node4209 : 4'b0001;
														assign node4209 = (inp[3]) ? 4'b0111 : 4'b0101;
												assign node4212 = (inp[15]) ? 4'b0001 : node4213;
													assign node4213 = (inp[9]) ? 4'b0001 : 4'b0101;
											assign node4217 = (inp[9]) ? node4221 : node4218;
												assign node4218 = (inp[15]) ? 4'b0001 : 4'b0111;
												assign node4221 = (inp[15]) ? 4'b0111 : 4'b0101;
										assign node4224 = (inp[5]) ? node4238 : node4225;
											assign node4225 = (inp[4]) ? node4231 : node4226;
												assign node4226 = (inp[9]) ? 4'b0101 : node4227;
													assign node4227 = (inp[15]) ? 4'b0011 : 4'b0001;
												assign node4231 = (inp[9]) ? node4235 : node4232;
													assign node4232 = (inp[1]) ? 4'b0101 : 4'b0111;
													assign node4235 = (inp[3]) ? 4'b0011 : 4'b0001;
											assign node4238 = (inp[15]) ? node4250 : node4239;
												assign node4239 = (inp[1]) ? node4245 : node4240;
													assign node4240 = (inp[4]) ? node4242 : 4'b0111;
														assign node4242 = (inp[9]) ? 4'b0011 : 4'b0111;
													assign node4245 = (inp[3]) ? node4247 : 4'b0011;
														assign node4247 = (inp[9]) ? 4'b0111 : 4'b0011;
												assign node4250 = (inp[9]) ? node4252 : 4'b0011;
													assign node4252 = (inp[4]) ? 4'b0001 : 4'b0101;
				assign node4255 = (inp[8]) ? node5005 : node4256;
					assign node4256 = (inp[15]) ? node4636 : node4257;
						assign node4257 = (inp[13]) ? node4437 : node4258;
							assign node4258 = (inp[5]) ? node4350 : node4259;
								assign node4259 = (inp[0]) ? node4309 : node4260;
									assign node4260 = (inp[12]) ? node4284 : node4261;
										assign node4261 = (inp[1]) ? node4271 : node4262;
											assign node4262 = (inp[9]) ? node4266 : node4263;
												assign node4263 = (inp[4]) ? 4'b1011 : 4'b1111;
												assign node4266 = (inp[11]) ? node4268 : 4'b0111;
													assign node4268 = (inp[6]) ? 4'b1011 : 4'b0011;
											assign node4271 = (inp[10]) ? node4281 : node4272;
												assign node4272 = (inp[4]) ? node4278 : node4273;
													assign node4273 = (inp[9]) ? node4275 : 4'b1111;
														assign node4275 = (inp[3]) ? 4'b0011 : 4'b0011;
													assign node4278 = (inp[9]) ? 4'b1111 : 4'b1011;
												assign node4281 = (inp[3]) ? 4'b1101 : 4'b1111;
										assign node4284 = (inp[3]) ? node4298 : node4285;
											assign node4285 = (inp[4]) ? node4291 : node4286;
												assign node4286 = (inp[11]) ? 4'b1011 : node4287;
													assign node4287 = (inp[1]) ? 4'b1011 : 4'b0111;
												assign node4291 = (inp[9]) ? node4295 : node4292;
													assign node4292 = (inp[10]) ? 4'b0111 : 4'b0011;
													assign node4295 = (inp[11]) ? 4'b1011 : 4'b1111;
											assign node4298 = (inp[10]) ? node4306 : node4299;
												assign node4299 = (inp[9]) ? node4301 : 4'b0011;
													assign node4301 = (inp[6]) ? 4'b1101 : node4302;
														assign node4302 = (inp[1]) ? 4'b0011 : 4'b1011;
												assign node4306 = (inp[11]) ? 4'b0101 : 4'b0001;
									assign node4309 = (inp[3]) ? node4325 : node4310;
										assign node4310 = (inp[1]) ? node4316 : node4311;
											assign node4311 = (inp[6]) ? node4313 : 4'b0001;
												assign node4313 = (inp[11]) ? 4'b1001 : 4'b0001;
											assign node4316 = (inp[12]) ? 4'b1001 : node4317;
												assign node4317 = (inp[10]) ? node4321 : node4318;
													assign node4318 = (inp[9]) ? 4'b0101 : 4'b0001;
													assign node4321 = (inp[11]) ? 4'b1101 : 4'b0101;
										assign node4325 = (inp[9]) ? node4341 : node4326;
											assign node4326 = (inp[4]) ? node4334 : node4327;
												assign node4327 = (inp[12]) ? 4'b1001 : node4328;
													assign node4328 = (inp[10]) ? node4330 : 4'b1101;
														assign node4330 = (inp[1]) ? 4'b1001 : 4'b1101;
												assign node4334 = (inp[6]) ? 4'b1111 : node4335;
													assign node4335 = (inp[10]) ? 4'b0001 : node4336;
														assign node4336 = (inp[12]) ? 4'b0001 : 4'b1001;
											assign node4341 = (inp[11]) ? node4343 : 4'b0001;
												assign node4343 = (inp[12]) ? 4'b1011 : node4344;
													assign node4344 = (inp[1]) ? 4'b0111 : node4345;
														assign node4345 = (inp[10]) ? 4'b1011 : 4'b1111;
								assign node4350 = (inp[0]) ? node4392 : node4351;
									assign node4351 = (inp[9]) ? node4369 : node4352;
										assign node4352 = (inp[3]) ? node4362 : node4353;
											assign node4353 = (inp[1]) ? node4357 : node4354;
												assign node4354 = (inp[10]) ? 4'b0011 : 4'b1111;
												assign node4357 = (inp[4]) ? node4359 : 4'b1011;
													assign node4359 = (inp[6]) ? 4'b0101 : 4'b1101;
											assign node4362 = (inp[1]) ? 4'b0001 : node4363;
												assign node4363 = (inp[4]) ? node4365 : 4'b0101;
													assign node4365 = (inp[6]) ? 4'b1101 : 4'b0101;
										assign node4369 = (inp[3]) ? node4375 : node4370;
											assign node4370 = (inp[11]) ? node4372 : 4'b1101;
												assign node4372 = (inp[1]) ? 4'b1001 : 4'b0101;
											assign node4375 = (inp[6]) ? node4385 : node4376;
												assign node4376 = (inp[4]) ? node4378 : 4'b1101;
													assign node4378 = (inp[10]) ? node4382 : node4379;
														assign node4379 = (inp[11]) ? 4'b1001 : 4'b1101;
														assign node4382 = (inp[1]) ? 4'b0001 : 4'b1001;
												assign node4385 = (inp[4]) ? node4389 : node4386;
													assign node4386 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node4389 = (inp[1]) ? 4'b0101 : 4'b1001;
									assign node4392 = (inp[3]) ? node4418 : node4393;
										assign node4393 = (inp[4]) ? node4405 : node4394;
											assign node4394 = (inp[10]) ? node4396 : 4'b1001;
												assign node4396 = (inp[1]) ? 4'b1001 : node4397;
													assign node4397 = (inp[6]) ? node4401 : node4398;
														assign node4398 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node4401 = (inp[12]) ? 4'b0111 : 4'b0101;
											assign node4405 = (inp[9]) ? node4411 : node4406;
												assign node4406 = (inp[12]) ? 4'b1111 : node4407;
													assign node4407 = (inp[6]) ? 4'b0001 : 4'b1001;
												assign node4411 = (inp[10]) ? 4'b1011 : node4412;
													assign node4412 = (inp[11]) ? 4'b0111 : node4413;
														assign node4413 = (inp[1]) ? 4'b0111 : 4'b1111;
										assign node4418 = (inp[10]) ? node4430 : node4419;
											assign node4419 = (inp[1]) ? node4425 : node4420;
												assign node4420 = (inp[11]) ? 4'b1111 : node4421;
													assign node4421 = (inp[9]) ? 4'b1111 : 4'b1011;
												assign node4425 = (inp[6]) ? node4427 : 4'b1011;
													assign node4427 = (inp[9]) ? 4'b1011 : 4'b0111;
											assign node4430 = (inp[4]) ? node4434 : node4431;
												assign node4431 = (inp[11]) ? 4'b0011 : 4'b1011;
												assign node4434 = (inp[11]) ? 4'b0011 : 4'b0111;
							assign node4437 = (inp[0]) ? node4537 : node4438;
								assign node4438 = (inp[3]) ? node4490 : node4439;
									assign node4439 = (inp[5]) ? node4457 : node4440;
										assign node4440 = (inp[6]) ? node4450 : node4441;
											assign node4441 = (inp[11]) ? node4445 : node4442;
												assign node4442 = (inp[4]) ? 4'b0011 : 4'b0111;
												assign node4445 = (inp[1]) ? 4'b1111 : node4446;
													assign node4446 = (inp[4]) ? 4'b1111 : 4'b1011;
											assign node4450 = (inp[11]) ? node4452 : 4'b1111;
												assign node4452 = (inp[10]) ? 4'b0111 : node4453;
													assign node4453 = (inp[12]) ? 4'b0111 : 4'b0011;
										assign node4457 = (inp[10]) ? node4481 : node4458;
											assign node4458 = (inp[4]) ? node4468 : node4459;
												assign node4459 = (inp[11]) ? node4465 : node4460;
													assign node4460 = (inp[6]) ? node4462 : 4'b0111;
														assign node4462 = (inp[1]) ? 4'b1011 : 4'b1011;
													assign node4465 = (inp[1]) ? 4'b0011 : 4'b0101;
												assign node4468 = (inp[12]) ? node4476 : node4469;
													assign node4469 = (inp[6]) ? node4473 : node4470;
														assign node4470 = (inp[11]) ? 4'b1101 : 4'b0101;
														assign node4473 = (inp[11]) ? 4'b0101 : 4'b1101;
													assign node4476 = (inp[6]) ? node4478 : 4'b0011;
														assign node4478 = (inp[1]) ? 4'b1101 : 4'b0101;
											assign node4481 = (inp[11]) ? node4485 : node4482;
												assign node4482 = (inp[12]) ? 4'b0101 : 4'b1101;
												assign node4485 = (inp[4]) ? node4487 : 4'b1101;
													assign node4487 = (inp[9]) ? 4'b1001 : 4'b1101;
									assign node4490 = (inp[11]) ? node4516 : node4491;
										assign node4491 = (inp[6]) ? node4501 : node4492;
											assign node4492 = (inp[12]) ? node4494 : 4'b0011;
												assign node4494 = (inp[5]) ? 4'b0001 : node4495;
													assign node4495 = (inp[1]) ? 4'b0101 : node4496;
														assign node4496 = (inp[4]) ? 4'b0001 : 4'b0101;
											assign node4501 = (inp[9]) ? node4507 : node4502;
												assign node4502 = (inp[4]) ? 4'b1101 : node4503;
													assign node4503 = (inp[5]) ? 4'b1001 : 4'b1011;
												assign node4507 = (inp[4]) ? node4511 : node4508;
													assign node4508 = (inp[12]) ? 4'b1101 : 4'b1001;
													assign node4511 = (inp[10]) ? 4'b1001 : node4512;
														assign node4512 = (inp[1]) ? 4'b1101 : 4'b1001;
										assign node4516 = (inp[6]) ? node4522 : node4517;
											assign node4517 = (inp[5]) ? node4519 : 4'b1101;
												assign node4519 = (inp[9]) ? 4'b1001 : 4'b1101;
											assign node4522 = (inp[5]) ? node4532 : node4523;
												assign node4523 = (inp[1]) ? node4529 : node4524;
													assign node4524 = (inp[9]) ? node4526 : 4'b0101;
														assign node4526 = (inp[4]) ? 4'b0001 : 4'b0101;
													assign node4529 = (inp[9]) ? 4'b0101 : 4'b0011;
												assign node4532 = (inp[4]) ? 4'b0101 : node4533;
													assign node4533 = (inp[9]) ? 4'b0101 : 4'b0001;
								assign node4537 = (inp[3]) ? node4587 : node4538;
									assign node4538 = (inp[5]) ? node4566 : node4539;
										assign node4539 = (inp[12]) ? node4555 : node4540;
											assign node4540 = (inp[10]) ? node4552 : node4541;
												assign node4541 = (inp[9]) ? node4547 : node4542;
													assign node4542 = (inp[4]) ? 4'b1001 : node4543;
														assign node4543 = (inp[6]) ? 4'b0101 : 4'b0101;
													assign node4547 = (inp[6]) ? node4549 : 4'b0101;
														assign node4549 = (inp[11]) ? 4'b0101 : 4'b1101;
												assign node4552 = (inp[11]) ? 4'b1101 : 4'b1001;
											assign node4555 = (inp[4]) ? node4561 : node4556;
												assign node4556 = (inp[9]) ? node4558 : 4'b0001;
													assign node4558 = (inp[11]) ? 4'b1101 : 4'b0101;
												assign node4561 = (inp[9]) ? node4563 : 4'b1101;
													assign node4563 = (inp[1]) ? 4'b0001 : 4'b1001;
										assign node4566 = (inp[12]) ? node4578 : node4567;
											assign node4567 = (inp[4]) ? node4575 : node4568;
												assign node4568 = (inp[11]) ? node4570 : 4'b1001;
													assign node4570 = (inp[6]) ? node4572 : 4'b1001;
														assign node4572 = (inp[10]) ? 4'b0001 : 4'b0101;
												assign node4575 = (inp[10]) ? 4'b1111 : 4'b1001;
											assign node4578 = (inp[4]) ? node4582 : node4579;
												assign node4579 = (inp[11]) ? 4'b1111 : 4'b1001;
												assign node4582 = (inp[1]) ? 4'b0001 : node4583;
													assign node4583 = (inp[9]) ? 4'b0011 : 4'b0111;
									assign node4587 = (inp[9]) ? node4611 : node4588;
										assign node4588 = (inp[5]) ? node4598 : node4589;
											assign node4589 = (inp[1]) ? node4593 : node4590;
												assign node4590 = (inp[11]) ? 4'b0001 : 4'b1111;
												assign node4593 = (inp[10]) ? 4'b1001 : node4594;
													assign node4594 = (inp[4]) ? 4'b1001 : 4'b1101;
											assign node4598 = (inp[1]) ? node4606 : node4599;
												assign node4599 = (inp[12]) ? 4'b0011 : node4600;
													assign node4600 = (inp[6]) ? node4602 : 4'b1011;
														assign node4602 = (inp[10]) ? 4'b1111 : 4'b1011;
												assign node4606 = (inp[12]) ? node4608 : 4'b0111;
													assign node4608 = (inp[4]) ? 4'b1111 : 4'b1011;
										assign node4611 = (inp[1]) ? node4623 : node4612;
											assign node4612 = (inp[4]) ? node4618 : node4613;
												assign node4613 = (inp[12]) ? 4'b1111 : node4614;
													assign node4614 = (inp[10]) ? 4'b1111 : 4'b1011;
												assign node4618 = (inp[10]) ? 4'b0011 : node4619;
													assign node4619 = (inp[12]) ? 4'b1011 : 4'b1111;
											assign node4623 = (inp[5]) ? node4629 : node4624;
												assign node4624 = (inp[10]) ? node4626 : 4'b0001;
													assign node4626 = (inp[4]) ? 4'b0011 : 4'b0111;
												assign node4629 = (inp[10]) ? 4'b0011 : node4630;
													assign node4630 = (inp[11]) ? node4632 : 4'b1111;
														assign node4632 = (inp[12]) ? 4'b0111 : 4'b0011;
						assign node4636 = (inp[10]) ? node4816 : node4637;
							assign node4637 = (inp[11]) ? node4719 : node4638;
								assign node4638 = (inp[6]) ? node4670 : node4639;
									assign node4639 = (inp[1]) ? node4651 : node4640;
										assign node4640 = (inp[13]) ? node4648 : node4641;
											assign node4641 = (inp[0]) ? 4'b1011 : node4642;
												assign node4642 = (inp[4]) ? 4'b1001 : node4643;
													assign node4643 = (inp[9]) ? 4'b1001 : 4'b1101;
											assign node4648 = (inp[4]) ? 4'b0101 : 4'b0001;
										assign node4651 = (inp[4]) ? node4661 : node4652;
											assign node4652 = (inp[9]) ? node4658 : node4653;
												assign node4653 = (inp[13]) ? 4'b0111 : node4654;
													assign node4654 = (inp[5]) ? 4'b0111 : 4'b0101;
												assign node4658 = (inp[13]) ? 4'b0001 : 4'b0011;
											assign node4661 = (inp[9]) ? node4667 : node4662;
												assign node4662 = (inp[5]) ? 4'b0001 : node4663;
													assign node4663 = (inp[0]) ? 4'b0011 : 4'b0001;
												assign node4667 = (inp[13]) ? 4'b0111 : 4'b0101;
									assign node4670 = (inp[1]) ? node4696 : node4671;
										assign node4671 = (inp[13]) ? node4685 : node4672;
											assign node4672 = (inp[3]) ? node4678 : node4673;
												assign node4673 = (inp[5]) ? node4675 : 4'b0001;
													assign node4675 = (inp[12]) ? 4'b0001 : 4'b0101;
												assign node4678 = (inp[12]) ? node4680 : 4'b0101;
													assign node4680 = (inp[5]) ? node4682 : 4'b0111;
														assign node4682 = (inp[4]) ? 4'b0111 : 4'b0001;
											assign node4685 = (inp[3]) ? node4687 : 4'b1101;
												assign node4687 = (inp[4]) ? node4691 : node4688;
													assign node4688 = (inp[5]) ? 4'b1101 : 4'b1011;
													assign node4691 = (inp[5]) ? 4'b1011 : node4692;
														assign node4692 = (inp[12]) ? 4'b1001 : 4'b1001;
										assign node4696 = (inp[4]) ? node4702 : node4697;
											assign node4697 = (inp[0]) ? 4'b1101 : node4698;
												assign node4698 = (inp[12]) ? 4'b1001 : 4'b1101;
											assign node4702 = (inp[13]) ? node4712 : node4703;
												assign node4703 = (inp[3]) ? node4709 : node4704;
													assign node4704 = (inp[12]) ? node4706 : 4'b1101;
														assign node4706 = (inp[9]) ? 4'b1011 : 4'b1111;
													assign node4709 = (inp[12]) ? 4'b1101 : 4'b1001;
												assign node4712 = (inp[9]) ? node4716 : node4713;
													assign node4713 = (inp[3]) ? 4'b1011 : 4'b1001;
													assign node4716 = (inp[3]) ? 4'b1111 : 4'b1011;
								assign node4719 = (inp[6]) ? node4765 : node4720;
									assign node4720 = (inp[1]) ? node4748 : node4721;
										assign node4721 = (inp[13]) ? node4737 : node4722;
											assign node4722 = (inp[0]) ? node4730 : node4723;
												assign node4723 = (inp[3]) ? 4'b0001 : node4724;
													assign node4724 = (inp[4]) ? node4726 : 4'b0101;
														assign node4726 = (inp[12]) ? 4'b0101 : 4'b0001;
												assign node4730 = (inp[9]) ? node4734 : node4731;
													assign node4731 = (inp[5]) ? 4'b0101 : 4'b0111;
													assign node4734 = (inp[4]) ? 4'b0111 : 4'b0011;
											assign node4737 = (inp[3]) ? node4745 : node4738;
												assign node4738 = (inp[5]) ? node4740 : 4'b1101;
													assign node4740 = (inp[12]) ? 4'b1111 : node4741;
														assign node4741 = (inp[0]) ? 4'b1111 : 4'b1001;
												assign node4745 = (inp[12]) ? 4'b1001 : 4'b1101;
										assign node4748 = (inp[12]) ? node4754 : node4749;
											assign node4749 = (inp[5]) ? 4'b1111 : node4750;
												assign node4750 = (inp[0]) ? 4'b1011 : 4'b1111;
											assign node4754 = (inp[5]) ? node4762 : node4755;
												assign node4755 = (inp[9]) ? 4'b1101 : node4756;
													assign node4756 = (inp[4]) ? 4'b1101 : node4757;
														assign node4757 = (inp[0]) ? 4'b1011 : 4'b1001;
												assign node4762 = (inp[0]) ? 4'b1101 : 4'b1111;
									assign node4765 = (inp[13]) ? node4791 : node4766;
										assign node4766 = (inp[1]) ? node4778 : node4767;
											assign node4767 = (inp[5]) ? node4773 : node4768;
												assign node4768 = (inp[0]) ? node4770 : 4'b1001;
													assign node4770 = (inp[3]) ? 4'b1011 : 4'b1111;
												assign node4773 = (inp[0]) ? 4'b1101 : node4774;
													assign node4774 = (inp[3]) ? 4'b1111 : 4'b1101;
											assign node4778 = (inp[9]) ? node4788 : node4779;
												assign node4779 = (inp[12]) ? node4785 : node4780;
													assign node4780 = (inp[5]) ? 4'b0101 : node4781;
														assign node4781 = (inp[0]) ? 4'b0111 : 4'b0101;
													assign node4785 = (inp[4]) ? 4'b0101 : 4'b0001;
												assign node4788 = (inp[5]) ? 4'b0111 : 4'b0011;
										assign node4791 = (inp[9]) ? node4805 : node4792;
											assign node4792 = (inp[1]) ? node4798 : node4793;
												assign node4793 = (inp[0]) ? 4'b0011 : node4794;
													assign node4794 = (inp[5]) ? 4'b0011 : 4'b0001;
												assign node4798 = (inp[5]) ? 4'b0011 : node4799;
													assign node4799 = (inp[12]) ? node4801 : 4'b0111;
														assign node4801 = (inp[4]) ? 4'b0111 : 4'b0011;
											assign node4805 = (inp[3]) ? node4811 : node4806;
												assign node4806 = (inp[4]) ? node4808 : 4'b0101;
													assign node4808 = (inp[0]) ? 4'b0101 : 4'b0111;
												assign node4811 = (inp[12]) ? node4813 : 4'b0011;
													assign node4813 = (inp[0]) ? 4'b0101 : 4'b0011;
							assign node4816 = (inp[6]) ? node4924 : node4817;
								assign node4817 = (inp[11]) ? node4873 : node4818;
									assign node4818 = (inp[1]) ? node4848 : node4819;
										assign node4819 = (inp[13]) ? node4839 : node4820;
											assign node4820 = (inp[4]) ? node4832 : node4821;
												assign node4821 = (inp[12]) ? node4829 : node4822;
													assign node4822 = (inp[0]) ? node4826 : node4823;
														assign node4823 = (inp[5]) ? 4'b1111 : 4'b1101;
														assign node4826 = (inp[5]) ? 4'b1101 : 4'b1111;
													assign node4829 = (inp[9]) ? 4'b1111 : 4'b1001;
												assign node4832 = (inp[12]) ? 4'b1111 : node4833;
													assign node4833 = (inp[0]) ? node4835 : 4'b1011;
														assign node4835 = (inp[3]) ? 4'b1001 : 4'b1011;
											assign node4839 = (inp[5]) ? 4'b0001 : node4840;
												assign node4840 = (inp[0]) ? node4844 : node4841;
													assign node4841 = (inp[3]) ? 4'b0111 : 4'b0101;
													assign node4844 = (inp[9]) ? 4'b0011 : 4'b0111;
										assign node4848 = (inp[13]) ? node4860 : node4849;
											assign node4849 = (inp[5]) ? node4857 : node4850;
												assign node4850 = (inp[0]) ? node4852 : 4'b0101;
													assign node4852 = (inp[4]) ? node4854 : 4'b0011;
														assign node4854 = (inp[12]) ? 4'b0101 : 4'b0111;
												assign node4857 = (inp[9]) ? 4'b0101 : 4'b0001;
											assign node4860 = (inp[5]) ? node4870 : node4861;
												assign node4861 = (inp[0]) ? node4865 : node4862;
													assign node4862 = (inp[4]) ? 4'b0101 : 4'b0001;
													assign node4865 = (inp[3]) ? node4867 : 4'b0111;
														assign node4867 = (inp[9]) ? 4'b0101 : 4'b0111;
												assign node4870 = (inp[0]) ? 4'b0101 : 4'b0111;
									assign node4873 = (inp[13]) ? node4893 : node4874;
										assign node4874 = (inp[1]) ? node4886 : node4875;
											assign node4875 = (inp[12]) ? node4879 : node4876;
												assign node4876 = (inp[3]) ? 4'b0011 : 4'b0111;
												assign node4879 = (inp[0]) ? node4881 : 4'b0111;
													assign node4881 = (inp[4]) ? node4883 : 4'b0101;
														assign node4883 = (inp[3]) ? 4'b0101 : 4'b0111;
											assign node4886 = (inp[4]) ? node4890 : node4887;
												assign node4887 = (inp[9]) ? 4'b1111 : 4'b1011;
												assign node4890 = (inp[3]) ? 4'b1001 : 4'b1011;
										assign node4893 = (inp[0]) ? node4913 : node4894;
											assign node4894 = (inp[5]) ? node4900 : node4895;
												assign node4895 = (inp[3]) ? 4'b1111 : node4896;
													assign node4896 = (inp[4]) ? 4'b1101 : 4'b1001;
												assign node4900 = (inp[1]) ? node4908 : node4901;
													assign node4901 = (inp[4]) ? node4905 : node4902;
														assign node4902 = (inp[9]) ? 4'b1111 : 4'b1011;
														assign node4905 = (inp[9]) ? 4'b1011 : 4'b1111;
													assign node4908 = (inp[4]) ? 4'b1011 : node4909;
														assign node4909 = (inp[9]) ? 4'b1111 : 4'b1011;
											assign node4913 = (inp[3]) ? node4915 : 4'b1111;
												assign node4915 = (inp[5]) ? node4919 : node4916;
													assign node4916 = (inp[4]) ? 4'b1001 : 4'b1011;
													assign node4919 = (inp[1]) ? node4921 : 4'b1101;
														assign node4921 = (inp[9]) ? 4'b1001 : 4'b1101;
								assign node4924 = (inp[11]) ? node4964 : node4925;
									assign node4925 = (inp[1]) ? node4941 : node4926;
										assign node4926 = (inp[13]) ? node4938 : node4927;
											assign node4927 = (inp[5]) ? node4933 : node4928;
												assign node4928 = (inp[12]) ? node4930 : 4'b0001;
													assign node4930 = (inp[9]) ? 4'b0001 : 4'b0111;
												assign node4933 = (inp[9]) ? node4935 : 4'b0101;
													assign node4935 = (inp[12]) ? 4'b0011 : 4'b0111;
											assign node4938 = (inp[5]) ? 4'b1001 : 4'b1111;
										assign node4941 = (inp[12]) ? node4951 : node4942;
											assign node4942 = (inp[9]) ? node4948 : node4943;
												assign node4943 = (inp[4]) ? node4945 : 4'b1011;
													assign node4945 = (inp[3]) ? 4'b1101 : 4'b1111;
												assign node4948 = (inp[5]) ? 4'b1001 : 4'b1011;
											assign node4951 = (inp[3]) ? 4'b1101 : node4952;
												assign node4952 = (inp[0]) ? node4958 : node4953;
													assign node4953 = (inp[5]) ? 4'b1111 : node4954;
														assign node4954 = (inp[9]) ? 4'b1101 : 4'b1001;
													assign node4958 = (inp[5]) ? 4'b1001 : node4959;
														assign node4959 = (inp[13]) ? 4'b1111 : 4'b1011;
									assign node4964 = (inp[5]) ? node4986 : node4965;
										assign node4965 = (inp[3]) ? node4975 : node4966;
											assign node4966 = (inp[0]) ? 4'b0111 : node4967;
												assign node4967 = (inp[13]) ? node4969 : 4'b1101;
													assign node4969 = (inp[9]) ? 4'b0101 : node4970;
														assign node4970 = (inp[4]) ? 4'b0101 : 4'b0001;
											assign node4975 = (inp[12]) ? node4981 : node4976;
												assign node4976 = (inp[4]) ? 4'b0011 : node4977;
													assign node4977 = (inp[9]) ? 4'b0111 : 4'b0011;
												assign node4981 = (inp[9]) ? node4983 : 4'b1111;
													assign node4983 = (inp[4]) ? 4'b0011 : 4'b0101;
										assign node4986 = (inp[0]) ? node5000 : node4987;
											assign node4987 = (inp[1]) ? node4991 : node4988;
												assign node4988 = (inp[12]) ? 4'b0011 : 4'b1011;
												assign node4991 = (inp[3]) ? node4995 : node4992;
													assign node4992 = (inp[9]) ? 4'b0011 : 4'b0111;
													assign node4995 = (inp[4]) ? 4'b0011 : node4996;
														assign node4996 = (inp[9]) ? 4'b0111 : 4'b0011;
											assign node5000 = (inp[3]) ? 4'b0001 : node5001;
												assign node5001 = (inp[4]) ? 4'b0101 : 4'b0011;
					assign node5005 = (inp[11]) ? node5377 : node5006;
						assign node5006 = (inp[6]) ? node5184 : node5007;
							assign node5007 = (inp[1]) ? node5075 : node5008;
								assign node5008 = (inp[13]) ? node5046 : node5009;
									assign node5009 = (inp[4]) ? node5033 : node5010;
										assign node5010 = (inp[9]) ? node5024 : node5011;
											assign node5011 = (inp[5]) ? node5017 : node5012;
												assign node5012 = (inp[15]) ? node5014 : 4'b1100;
													assign node5014 = (inp[3]) ? 4'b1110 : 4'b1100;
												assign node5017 = (inp[3]) ? 4'b1110 : node5018;
													assign node5018 = (inp[12]) ? node5020 : 4'b1100;
														assign node5020 = (inp[15]) ? 4'b1100 : 4'b1110;
											assign node5024 = (inp[10]) ? node5030 : node5025;
												assign node5025 = (inp[0]) ? 4'b1010 : node5026;
													assign node5026 = (inp[15]) ? 4'b1000 : 4'b1010;
												assign node5030 = (inp[12]) ? 4'b1110 : 4'b1010;
										assign node5033 = (inp[9]) ? node5039 : node5034;
											assign node5034 = (inp[10]) ? 4'b1010 : node5035;
												assign node5035 = (inp[5]) ? 4'b1010 : 4'b1000;
											assign node5039 = (inp[12]) ? node5043 : node5040;
												assign node5040 = (inp[15]) ? 4'b1100 : 4'b1110;
												assign node5043 = (inp[5]) ? 4'b1010 : 4'b1000;
									assign node5046 = (inp[3]) ? node5054 : node5047;
										assign node5047 = (inp[4]) ? 4'b0010 : node5048;
											assign node5048 = (inp[15]) ? node5050 : 4'b0010;
												assign node5050 = (inp[10]) ? 4'b0110 : 4'b0100;
										assign node5054 = (inp[12]) ? node5068 : node5055;
											assign node5055 = (inp[0]) ? node5061 : node5056;
												assign node5056 = (inp[4]) ? 4'b0000 : node5057;
													assign node5057 = (inp[9]) ? 4'b0010 : 4'b0110;
												assign node5061 = (inp[10]) ? node5063 : 4'b0110;
													assign node5063 = (inp[9]) ? 4'b0000 : node5064;
														assign node5064 = (inp[4]) ? 4'b0000 : 4'b0100;
											assign node5068 = (inp[10]) ? 4'b0110 : node5069;
												assign node5069 = (inp[9]) ? node5071 : 4'b0100;
													assign node5071 = (inp[5]) ? 4'b0110 : 4'b0100;
								assign node5075 = (inp[13]) ? node5125 : node5076;
									assign node5076 = (inp[5]) ? node5102 : node5077;
										assign node5077 = (inp[3]) ? node5087 : node5078;
											assign node5078 = (inp[10]) ? node5082 : node5079;
												assign node5079 = (inp[9]) ? 4'b0100 : 4'b0000;
												assign node5082 = (inp[12]) ? 4'b0000 : node5083;
													assign node5083 = (inp[15]) ? 4'b0000 : 4'b0100;
											assign node5087 = (inp[4]) ? node5093 : node5088;
												assign node5088 = (inp[9]) ? node5090 : 4'b0100;
													assign node5090 = (inp[15]) ? 4'b0110 : 4'b0100;
												assign node5093 = (inp[12]) ? node5095 : 4'b0000;
													assign node5095 = (inp[15]) ? node5099 : node5096;
														assign node5096 = (inp[10]) ? 4'b0110 : 4'b0100;
														assign node5099 = (inp[10]) ? 4'b0100 : 4'b0000;
										assign node5102 = (inp[3]) ? node5114 : node5103;
											assign node5103 = (inp[15]) ? node5109 : node5104;
												assign node5104 = (inp[12]) ? 4'b0000 : node5105;
													assign node5105 = (inp[4]) ? 4'b0010 : 4'b0110;
												assign node5109 = (inp[12]) ? node5111 : 4'b0100;
													assign node5111 = (inp[10]) ? 4'b0110 : 4'b0100;
											assign node5114 = (inp[4]) ? node5120 : node5115;
												assign node5115 = (inp[15]) ? 4'b0010 : node5116;
													assign node5116 = (inp[0]) ? 4'b0010 : 4'b0000;
												assign node5120 = (inp[0]) ? node5122 : 4'b0000;
													assign node5122 = (inp[12]) ? 4'b0000 : 4'b0100;
									assign node5125 = (inp[12]) ? node5155 : node5126;
										assign node5126 = (inp[10]) ? node5136 : node5127;
											assign node5127 = (inp[5]) ? node5133 : node5128;
												assign node5128 = (inp[0]) ? node5130 : 4'b0000;
													assign node5130 = (inp[15]) ? 4'b0010 : 4'b0000;
												assign node5133 = (inp[15]) ? 4'b0100 : 4'b0010;
											assign node5136 = (inp[0]) ? node5144 : node5137;
												assign node5137 = (inp[9]) ? 4'b0100 : node5138;
													assign node5138 = (inp[4]) ? node5140 : 4'b0110;
														assign node5140 = (inp[15]) ? 4'b0000 : 4'b0010;
												assign node5144 = (inp[4]) ? node5148 : node5145;
													assign node5145 = (inp[9]) ? 4'b0000 : 4'b0100;
													assign node5148 = (inp[15]) ? node5152 : node5149;
														assign node5149 = (inp[3]) ? 4'b0110 : 4'b0100;
														assign node5152 = (inp[3]) ? 4'b0100 : 4'b0110;
										assign node5155 = (inp[4]) ? node5165 : node5156;
											assign node5156 = (inp[5]) ? node5158 : 4'b0110;
												assign node5158 = (inp[10]) ? 4'b0100 : node5159;
													assign node5159 = (inp[3]) ? 4'b0100 : node5160;
														assign node5160 = (inp[0]) ? 4'b0010 : 4'b0000;
											assign node5165 = (inp[0]) ? node5177 : node5166;
												assign node5166 = (inp[15]) ? node5172 : node5167;
													assign node5167 = (inp[3]) ? 4'b0100 : node5168;
														assign node5168 = (inp[5]) ? 4'b0100 : 4'b0110;
													assign node5172 = (inp[3]) ? 4'b0110 : node5173;
														assign node5173 = (inp[9]) ? 4'b0010 : 4'b0110;
												assign node5177 = (inp[3]) ? node5179 : 4'b0010;
													assign node5179 = (inp[10]) ? 4'b0010 : node5180;
														assign node5180 = (inp[15]) ? 4'b0100 : 4'b0110;
							assign node5184 = (inp[1]) ? node5282 : node5185;
								assign node5185 = (inp[13]) ? node5231 : node5186;
									assign node5186 = (inp[9]) ? node5212 : node5187;
										assign node5187 = (inp[4]) ? node5201 : node5188;
											assign node5188 = (inp[15]) ? node5196 : node5189;
												assign node5189 = (inp[10]) ? node5191 : 4'b0100;
													assign node5191 = (inp[0]) ? node5193 : 4'b0010;
														assign node5193 = (inp[12]) ? 4'b0000 : 4'b0100;
												assign node5196 = (inp[10]) ? 4'b0110 : node5197;
													assign node5197 = (inp[3]) ? 4'b0110 : 4'b0100;
											assign node5201 = (inp[10]) ? node5209 : node5202;
												assign node5202 = (inp[5]) ? 4'b0000 : node5203;
													assign node5203 = (inp[0]) ? 4'b0010 : node5204;
														assign node5204 = (inp[15]) ? 4'b0000 : 4'b0010;
												assign node5209 = (inp[12]) ? 4'b0100 : 4'b0000;
										assign node5212 = (inp[4]) ? node5216 : node5213;
											assign node5213 = (inp[12]) ? 4'b0100 : 4'b0010;
											assign node5216 = (inp[10]) ? node5224 : node5217;
												assign node5217 = (inp[5]) ? node5219 : 4'b0110;
													assign node5219 = (inp[3]) ? node5221 : 4'b0100;
														assign node5221 = (inp[0]) ? 4'b0100 : 4'b0110;
												assign node5224 = (inp[12]) ? 4'b0010 : node5225;
													assign node5225 = (inp[3]) ? node5227 : 4'b0110;
														assign node5227 = (inp[5]) ? 4'b0110 : 4'b0100;
									assign node5231 = (inp[10]) ? node5263 : node5232;
										assign node5232 = (inp[15]) ? node5246 : node5233;
											assign node5233 = (inp[0]) ? node5241 : node5234;
												assign node5234 = (inp[9]) ? 4'b1100 : node5235;
													assign node5235 = (inp[4]) ? 4'b1100 : node5236;
														assign node5236 = (inp[3]) ? 4'b1110 : 4'b1010;
												assign node5241 = (inp[12]) ? node5243 : 4'b1100;
													assign node5243 = (inp[4]) ? 4'b1100 : 4'b1000;
											assign node5246 = (inp[12]) ? node5258 : node5247;
												assign node5247 = (inp[3]) ? node5253 : node5248;
													assign node5248 = (inp[0]) ? 4'b1010 : node5249;
														assign node5249 = (inp[9]) ? 4'b1110 : 4'b1000;
													assign node5253 = (inp[9]) ? node5255 : 4'b1110;
														assign node5255 = (inp[4]) ? 4'b1100 : 4'b1000;
												assign node5258 = (inp[0]) ? 4'b1100 : node5259;
													assign node5259 = (inp[3]) ? 4'b1110 : 4'b1100;
										assign node5263 = (inp[15]) ? node5267 : node5264;
											assign node5264 = (inp[4]) ? 4'b1010 : 4'b1110;
											assign node5267 = (inp[0]) ? node5275 : node5268;
												assign node5268 = (inp[5]) ? 4'b1110 : node5269;
													assign node5269 = (inp[12]) ? 4'b1110 : node5270;
														assign node5270 = (inp[3]) ? 4'b1000 : 4'b1100;
												assign node5275 = (inp[5]) ? node5277 : 4'b1010;
													assign node5277 = (inp[9]) ? 4'b1000 : node5278;
														assign node5278 = (inp[3]) ? 4'b1000 : 4'b1100;
								assign node5282 = (inp[5]) ? node5336 : node5283;
									assign node5283 = (inp[0]) ? node5313 : node5284;
										assign node5284 = (inp[9]) ? node5296 : node5285;
											assign node5285 = (inp[4]) ? node5289 : node5286;
												assign node5286 = (inp[15]) ? 4'b1100 : 4'b1010;
												assign node5289 = (inp[10]) ? node5291 : 4'b1100;
													assign node5291 = (inp[15]) ? node5293 : 4'b1110;
														assign node5293 = (inp[3]) ? 4'b1110 : 4'b1100;
											assign node5296 = (inp[4]) ? node5304 : node5297;
												assign node5297 = (inp[3]) ? node5301 : node5298;
													assign node5298 = (inp[10]) ? 4'b1110 : 4'b1010;
													assign node5301 = (inp[15]) ? 4'b1110 : 4'b1100;
												assign node5304 = (inp[13]) ? node5308 : node5305;
													assign node5305 = (inp[12]) ? 4'b1000 : 4'b1010;
													assign node5308 = (inp[12]) ? 4'b1010 : node5309;
														assign node5309 = (inp[3]) ? 4'b1010 : 4'b1000;
										assign node5313 = (inp[10]) ? node5327 : node5314;
											assign node5314 = (inp[15]) ? node5318 : node5315;
												assign node5315 = (inp[13]) ? 4'b1100 : 4'b1110;
												assign node5318 = (inp[4]) ? node5322 : node5319;
													assign node5319 = (inp[9]) ? 4'b1010 : 4'b1110;
													assign node5322 = (inp[9]) ? node5324 : 4'b1010;
														assign node5324 = (inp[12]) ? 4'b1000 : 4'b1100;
											assign node5327 = (inp[15]) ? node5333 : node5328;
												assign node5328 = (inp[9]) ? node5330 : 4'b1000;
													assign node5330 = (inp[3]) ? 4'b1010 : 4'b1000;
												assign node5333 = (inp[4]) ? 4'b1110 : 4'b1010;
									assign node5336 = (inp[9]) ? node5358 : node5337;
										assign node5337 = (inp[4]) ? node5349 : node5338;
											assign node5338 = (inp[15]) ? node5344 : node5339;
												assign node5339 = (inp[10]) ? node5341 : 4'b1110;
													assign node5341 = (inp[13]) ? 4'b1000 : 4'b1010;
												assign node5344 = (inp[0]) ? node5346 : 4'b1000;
													assign node5346 = (inp[3]) ? 4'b1000 : 4'b1010;
											assign node5349 = (inp[12]) ? 4'b1100 : node5350;
												assign node5350 = (inp[10]) ? node5354 : node5351;
													assign node5351 = (inp[0]) ? 4'b1000 : 4'b1010;
													assign node5354 = (inp[0]) ? 4'b1100 : 4'b1110;
										assign node5358 = (inp[4]) ? node5370 : node5359;
											assign node5359 = (inp[10]) ? node5365 : node5360;
												assign node5360 = (inp[15]) ? 4'b1010 : node5361;
													assign node5361 = (inp[13]) ? 4'b1110 : 4'b1100;
												assign node5365 = (inp[0]) ? 4'b1100 : node5366;
													assign node5366 = (inp[15]) ? 4'b1110 : 4'b1100;
											assign node5370 = (inp[10]) ? 4'b1000 : node5371;
												assign node5371 = (inp[0]) ? 4'b1110 : node5372;
													assign node5372 = (inp[12]) ? 4'b1000 : 4'b1100;
						assign node5377 = (inp[6]) ? node5539 : node5378;
							assign node5378 = (inp[1]) ? node5458 : node5379;
								assign node5379 = (inp[13]) ? node5419 : node5380;
									assign node5380 = (inp[4]) ? node5394 : node5381;
										assign node5381 = (inp[9]) ? node5387 : node5382;
											assign node5382 = (inp[0]) ? 4'b0110 : node5383;
												assign node5383 = (inp[5]) ? 4'b0000 : 4'b0110;
											assign node5387 = (inp[5]) ? 4'b0110 : node5388;
												assign node5388 = (inp[15]) ? 4'b0010 : node5389;
													assign node5389 = (inp[0]) ? 4'b0000 : 4'b0010;
										assign node5394 = (inp[9]) ? node5404 : node5395;
											assign node5395 = (inp[10]) ? node5401 : node5396;
												assign node5396 = (inp[5]) ? node5398 : 4'b0000;
													assign node5398 = (inp[15]) ? 4'b0000 : 4'b0010;
												assign node5401 = (inp[5]) ? 4'b0100 : 4'b0110;
											assign node5404 = (inp[0]) ? node5414 : node5405;
												assign node5405 = (inp[10]) ? node5411 : node5406;
													assign node5406 = (inp[15]) ? node5408 : 4'b0100;
														assign node5408 = (inp[12]) ? 4'b0110 : 4'b0100;
													assign node5411 = (inp[12]) ? 4'b0000 : 4'b0100;
												assign node5414 = (inp[10]) ? node5416 : 4'b0110;
													assign node5416 = (inp[3]) ? 4'b0100 : 4'b0110;
									assign node5419 = (inp[5]) ? node5447 : node5420;
										assign node5420 = (inp[10]) ? node5438 : node5421;
											assign node5421 = (inp[0]) ? node5429 : node5422;
												assign node5422 = (inp[4]) ? node5424 : 4'b1010;
													assign node5424 = (inp[15]) ? 4'b1000 : node5425;
														assign node5425 = (inp[12]) ? 4'b1000 : 4'b1010;
												assign node5429 = (inp[9]) ? node5435 : node5430;
													assign node5430 = (inp[4]) ? 4'b1100 : node5431;
														assign node5431 = (inp[12]) ? 4'b1000 : 4'b1100;
													assign node5435 = (inp[3]) ? 4'b1010 : 4'b1000;
											assign node5438 = (inp[15]) ? node5444 : node5439;
												assign node5439 = (inp[4]) ? node5441 : 4'b1010;
													assign node5441 = (inp[9]) ? 4'b1010 : 4'b1110;
												assign node5444 = (inp[9]) ? 4'b1100 : 4'b1110;
										assign node5447 = (inp[12]) ? node5449 : 4'b1100;
											assign node5449 = (inp[0]) ? node5455 : node5450;
												assign node5450 = (inp[9]) ? 4'b1110 : node5451;
													assign node5451 = (inp[10]) ? 4'b1010 : 4'b1000;
												assign node5455 = (inp[15]) ? 4'b1100 : 4'b1110;
								assign node5458 = (inp[9]) ? node5500 : node5459;
									assign node5459 = (inp[4]) ? node5477 : node5460;
										assign node5460 = (inp[10]) ? node5468 : node5461;
											assign node5461 = (inp[12]) ? 4'b1010 : node5462;
												assign node5462 = (inp[13]) ? 4'b1110 : node5463;
													assign node5463 = (inp[15]) ? 4'b1110 : 4'b1100;
											assign node5468 = (inp[5]) ? node5470 : 4'b1010;
												assign node5470 = (inp[0]) ? node5472 : 4'b1000;
													assign node5472 = (inp[12]) ? 4'b1010 : node5473;
														assign node5473 = (inp[15]) ? 4'b1000 : 4'b1000;
										assign node5477 = (inp[10]) ? node5489 : node5478;
											assign node5478 = (inp[12]) ? node5484 : node5479;
												assign node5479 = (inp[0]) ? 4'b1010 : node5480;
													assign node5480 = (inp[13]) ? 4'b1000 : 4'b1010;
												assign node5484 = (inp[15]) ? node5486 : 4'b1100;
													assign node5486 = (inp[0]) ? 4'b1100 : 4'b1110;
											assign node5489 = (inp[3]) ? node5491 : 4'b1110;
												assign node5491 = (inp[13]) ? 4'b1100 : node5492;
													assign node5492 = (inp[0]) ? node5496 : node5493;
														assign node5493 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node5496 = (inp[15]) ? 4'b1100 : 4'b1110;
									assign node5500 = (inp[13]) ? node5520 : node5501;
										assign node5501 = (inp[0]) ? node5515 : node5502;
											assign node5502 = (inp[4]) ? node5508 : node5503;
												assign node5503 = (inp[15]) ? 4'b1110 : node5504;
													assign node5504 = (inp[10]) ? 4'b1100 : 4'b1000;
												assign node5508 = (inp[10]) ? node5512 : node5509;
													assign node5509 = (inp[12]) ? 4'b1010 : 4'b1110;
													assign node5512 = (inp[3]) ? 4'b1010 : 4'b1000;
											assign node5515 = (inp[15]) ? 4'b1010 : node5516;
												assign node5516 = (inp[12]) ? 4'b1100 : 4'b1110;
										assign node5520 = (inp[3]) ? node5530 : node5521;
											assign node5521 = (inp[15]) ? node5523 : 4'b1110;
												assign node5523 = (inp[10]) ? 4'b1110 : node5524;
													assign node5524 = (inp[4]) ? 4'b1100 : node5525;
														assign node5525 = (inp[0]) ? 4'b1110 : 4'b1100;
											assign node5530 = (inp[10]) ? node5534 : node5531;
												assign node5531 = (inp[12]) ? 4'b1100 : 4'b1000;
												assign node5534 = (inp[15]) ? 4'b1100 : node5535;
													assign node5535 = (inp[0]) ? 4'b1110 : 4'b1100;
							assign node5539 = (inp[13]) ? node5621 : node5540;
								assign node5540 = (inp[1]) ? node5584 : node5541;
									assign node5541 = (inp[0]) ? node5563 : node5542;
										assign node5542 = (inp[15]) ? node5554 : node5543;
											assign node5543 = (inp[3]) ? node5551 : node5544;
												assign node5544 = (inp[9]) ? node5548 : node5545;
													assign node5545 = (inp[5]) ? 4'b1010 : 4'b1110;
													assign node5548 = (inp[4]) ? 4'b1100 : 4'b1110;
												assign node5551 = (inp[5]) ? 4'b1100 : 4'b1000;
											assign node5554 = (inp[3]) ? 4'b1110 : node5555;
												assign node5555 = (inp[9]) ? node5557 : 4'b1100;
													assign node5557 = (inp[4]) ? 4'b1110 : node5558;
														assign node5558 = (inp[10]) ? 4'b1110 : 4'b1000;
										assign node5563 = (inp[9]) ? node5571 : node5564;
											assign node5564 = (inp[3]) ? 4'b1100 : node5565;
												assign node5565 = (inp[12]) ? node5567 : 4'b1100;
													assign node5567 = (inp[15]) ? 4'b1010 : 4'b1000;
											assign node5571 = (inp[4]) ? node5575 : node5572;
												assign node5572 = (inp[10]) ? 4'b1110 : 4'b1010;
												assign node5575 = (inp[10]) ? node5581 : node5576;
													assign node5576 = (inp[12]) ? 4'b1000 : node5577;
														assign node5577 = (inp[3]) ? 4'b1100 : 4'b1110;
													assign node5581 = (inp[3]) ? 4'b1000 : 4'b1010;
									assign node5584 = (inp[4]) ? node5604 : node5585;
										assign node5585 = (inp[9]) ? node5597 : node5586;
											assign node5586 = (inp[12]) ? node5592 : node5587;
												assign node5587 = (inp[15]) ? node5589 : 4'b0100;
													assign node5589 = (inp[3]) ? 4'b0000 : 4'b0010;
												assign node5592 = (inp[10]) ? node5594 : 4'b0010;
													assign node5594 = (inp[15]) ? 4'b0000 : 4'b0010;
											assign node5597 = (inp[10]) ? 4'b0110 : node5598;
												assign node5598 = (inp[5]) ? node5600 : 4'b0010;
													assign node5600 = (inp[15]) ? 4'b0000 : 4'b0100;
										assign node5604 = (inp[9]) ? node5612 : node5605;
											assign node5605 = (inp[5]) ? node5607 : 4'b0100;
												assign node5607 = (inp[10]) ? 4'b0110 : node5608;
													assign node5608 = (inp[0]) ? 4'b0100 : 4'b0110;
											assign node5612 = (inp[12]) ? node5616 : node5613;
												assign node5613 = (inp[10]) ? 4'b0000 : 4'b0100;
												assign node5616 = (inp[3]) ? node5618 : 4'b0010;
													assign node5618 = (inp[0]) ? 4'b0000 : 4'b0010;
								assign node5621 = (inp[12]) ? node5671 : node5622;
									assign node5622 = (inp[5]) ? node5638 : node5623;
										assign node5623 = (inp[3]) ? node5633 : node5624;
											assign node5624 = (inp[9]) ? node5626 : 4'b0000;
												assign node5626 = (inp[1]) ? 4'b0110 : node5627;
													assign node5627 = (inp[10]) ? 4'b0100 : node5628;
														assign node5628 = (inp[4]) ? 4'b0100 : 4'b0000;
											assign node5633 = (inp[4]) ? node5635 : 4'b0100;
												assign node5635 = (inp[15]) ? 4'b0110 : 4'b0100;
										assign node5638 = (inp[3]) ? node5656 : node5639;
											assign node5639 = (inp[0]) ? node5647 : node5640;
												assign node5640 = (inp[4]) ? node5642 : 4'b0010;
													assign node5642 = (inp[9]) ? node5644 : 4'b0010;
														assign node5644 = (inp[15]) ? 4'b0110 : 4'b0100;
												assign node5647 = (inp[4]) ? 4'b0100 : node5648;
													assign node5648 = (inp[10]) ? node5652 : node5649;
														assign node5649 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node5652 = (inp[9]) ? 4'b0110 : 4'b0010;
											assign node5656 = (inp[0]) ? node5662 : node5657;
												assign node5657 = (inp[10]) ? 4'b0000 : node5658;
													assign node5658 = (inp[15]) ? 4'b0110 : 4'b0100;
												assign node5662 = (inp[15]) ? node5668 : node5663;
													assign node5663 = (inp[4]) ? node5665 : 4'b0110;
														assign node5665 = (inp[10]) ? 4'b0010 : 4'b0010;
													assign node5668 = (inp[1]) ? 4'b0000 : 4'b0100;
									assign node5671 = (inp[3]) ? node5687 : node5672;
										assign node5672 = (inp[5]) ? node5680 : node5673;
											assign node5673 = (inp[10]) ? 4'b0000 : node5674;
												assign node5674 = (inp[15]) ? node5676 : 4'b0110;
													assign node5676 = (inp[0]) ? 4'b0110 : 4'b0000;
											assign node5680 = (inp[9]) ? node5684 : node5681;
												assign node5681 = (inp[4]) ? 4'b0110 : 4'b0000;
												assign node5684 = (inp[4]) ? 4'b0010 : 4'b0110;
										assign node5687 = (inp[1]) ? node5703 : node5688;
											assign node5688 = (inp[5]) ? node5698 : node5689;
												assign node5689 = (inp[4]) ? node5693 : node5690;
													assign node5690 = (inp[9]) ? 4'b0100 : 4'b0010;
													assign node5693 = (inp[9]) ? 4'b0010 : node5694;
														assign node5694 = (inp[15]) ? 4'b0110 : 4'b0100;
												assign node5698 = (inp[0]) ? 4'b0010 : node5699;
													assign node5699 = (inp[10]) ? 4'b0010 : 4'b0110;
											assign node5703 = (inp[9]) ? node5705 : 4'b0010;
												assign node5705 = (inp[4]) ? 4'b0010 : 4'b0110;
		assign node5708 = (inp[0]) ? node8310 : node5709;
			assign node5709 = (inp[7]) ? node7035 : node5710;
				assign node5710 = (inp[8]) ? node6338 : node5711;
					assign node5711 = (inp[6]) ? node6021 : node5712;
						assign node5712 = (inp[11]) ? node5862 : node5713;
							assign node5713 = (inp[1]) ? node5775 : node5714;
								assign node5714 = (inp[9]) ? node5740 : node5715;
									assign node5715 = (inp[4]) ? node5727 : node5716;
										assign node5716 = (inp[15]) ? node5722 : node5717;
											assign node5717 = (inp[10]) ? node5719 : 4'b1110;
												assign node5719 = (inp[5]) ? 4'b1110 : 4'b1010;
											assign node5722 = (inp[10]) ? node5724 : 4'b1100;
												assign node5724 = (inp[3]) ? 4'b1010 : 4'b1000;
										assign node5727 = (inp[13]) ? node5735 : node5728;
											assign node5728 = (inp[12]) ? node5730 : 4'b1010;
												assign node5730 = (inp[15]) ? node5732 : 4'b1000;
													assign node5732 = (inp[2]) ? 4'b1000 : 4'b1010;
											assign node5735 = (inp[15]) ? 4'b1000 : node5736;
												assign node5736 = (inp[2]) ? 4'b1000 : 4'b1010;
									assign node5740 = (inp[4]) ? node5756 : node5741;
										assign node5741 = (inp[3]) ? node5749 : node5742;
											assign node5742 = (inp[12]) ? node5744 : 4'b1010;
												assign node5744 = (inp[15]) ? node5746 : 4'b1100;
													assign node5746 = (inp[5]) ? 4'b1110 : 4'b1100;
											assign node5749 = (inp[13]) ? 4'b1010 : node5750;
												assign node5750 = (inp[5]) ? node5752 : 4'b1000;
													assign node5752 = (inp[15]) ? 4'b1010 : 4'b1000;
										assign node5756 = (inp[12]) ? node5768 : node5757;
											assign node5757 = (inp[15]) ? node5763 : node5758;
												assign node5758 = (inp[3]) ? 4'b1100 : node5759;
													assign node5759 = (inp[5]) ? 4'b1100 : 4'b1110;
												assign node5763 = (inp[5]) ? 4'b1110 : node5764;
													assign node5764 = (inp[10]) ? 4'b1100 : 4'b1110;
											assign node5768 = (inp[10]) ? node5772 : node5769;
												assign node5769 = (inp[13]) ? 4'b1110 : 4'b1100;
												assign node5772 = (inp[3]) ? 4'b1010 : 4'b1000;
								assign node5775 = (inp[13]) ? node5825 : node5776;
									assign node5776 = (inp[10]) ? node5802 : node5777;
										assign node5777 = (inp[15]) ? node5791 : node5778;
											assign node5778 = (inp[3]) ? node5788 : node5779;
												assign node5779 = (inp[9]) ? node5783 : node5780;
													assign node5780 = (inp[4]) ? 4'b1010 : 4'b1110;
													assign node5783 = (inp[4]) ? node5785 : 4'b1010;
														assign node5785 = (inp[12]) ? 4'b1110 : 4'b1100;
												assign node5788 = (inp[4]) ? 4'b1100 : 4'b1000;
											assign node5791 = (inp[5]) ? node5795 : node5792;
												assign node5792 = (inp[4]) ? 4'b1000 : 4'b1100;
												assign node5795 = (inp[3]) ? node5797 : 4'b1100;
													assign node5797 = (inp[9]) ? 4'b1110 : node5798;
														assign node5798 = (inp[2]) ? 4'b1010 : 4'b1110;
										assign node5802 = (inp[5]) ? node5818 : node5803;
											assign node5803 = (inp[15]) ? node5809 : node5804;
												assign node5804 = (inp[4]) ? 4'b1100 : node5805;
													assign node5805 = (inp[12]) ? 4'b1110 : 4'b1010;
												assign node5809 = (inp[3]) ? node5815 : node5810;
													assign node5810 = (inp[9]) ? node5812 : 4'b1000;
														assign node5812 = (inp[12]) ? 4'b1100 : 4'b1000;
													assign node5815 = (inp[12]) ? 4'b1010 : 4'b1000;
											assign node5818 = (inp[4]) ? node5820 : 4'b1100;
												assign node5820 = (inp[9]) ? node5822 : 4'b1110;
													assign node5822 = (inp[3]) ? 4'b1000 : 4'b1010;
									assign node5825 = (inp[9]) ? node5845 : node5826;
										assign node5826 = (inp[3]) ? node5836 : node5827;
											assign node5827 = (inp[15]) ? 4'b0100 : node5828;
												assign node5828 = (inp[4]) ? 4'b0100 : node5829;
													assign node5829 = (inp[2]) ? node5831 : 4'b0110;
														assign node5831 = (inp[12]) ? 4'b0010 : 4'b0110;
											assign node5836 = (inp[10]) ? node5840 : node5837;
												assign node5837 = (inp[4]) ? 4'b0010 : 4'b0110;
												assign node5840 = (inp[5]) ? node5842 : 4'b0010;
													assign node5842 = (inp[12]) ? 4'b0000 : 4'b0100;
										assign node5845 = (inp[4]) ? node5853 : node5846;
											assign node5846 = (inp[10]) ? node5848 : 4'b0000;
												assign node5848 = (inp[12]) ? 4'b0110 : node5849;
													assign node5849 = (inp[3]) ? 4'b0010 : 4'b0000;
											assign node5853 = (inp[10]) ? node5857 : node5854;
												assign node5854 = (inp[15]) ? 4'b0110 : 4'b0100;
												assign node5857 = (inp[3]) ? 4'b0010 : node5858;
													assign node5858 = (inp[12]) ? 4'b0000 : 4'b0100;
							assign node5862 = (inp[1]) ? node5930 : node5863;
								assign node5863 = (inp[9]) ? node5895 : node5864;
									assign node5864 = (inp[4]) ? node5878 : node5865;
										assign node5865 = (inp[10]) ? node5873 : node5866;
											assign node5866 = (inp[13]) ? node5868 : 4'b0100;
												assign node5868 = (inp[12]) ? node5870 : 4'b0110;
													assign node5870 = (inp[2]) ? 4'b0100 : 4'b0110;
											assign node5873 = (inp[12]) ? node5875 : 4'b0100;
												assign node5875 = (inp[15]) ? 4'b0000 : 4'b0010;
										assign node5878 = (inp[10]) ? node5890 : node5879;
											assign node5879 = (inp[15]) ? node5885 : node5880;
												assign node5880 = (inp[12]) ? node5882 : 4'b0010;
													assign node5882 = (inp[5]) ? 4'b0000 : 4'b0010;
												assign node5885 = (inp[5]) ? node5887 : 4'b0000;
													assign node5887 = (inp[3]) ? 4'b0010 : 4'b0000;
											assign node5890 = (inp[12]) ? node5892 : 4'b0010;
												assign node5892 = (inp[5]) ? 4'b0100 : 4'b0110;
									assign node5895 = (inp[4]) ? node5911 : node5896;
										assign node5896 = (inp[12]) ? node5900 : node5897;
											assign node5897 = (inp[15]) ? 4'b0000 : 4'b0010;
											assign node5900 = (inp[10]) ? node5904 : node5901;
												assign node5901 = (inp[3]) ? 4'b0000 : 4'b0010;
												assign node5904 = (inp[2]) ? 4'b0100 : node5905;
													assign node5905 = (inp[5]) ? node5907 : 4'b0100;
														assign node5907 = (inp[15]) ? 4'b0110 : 4'b0100;
										assign node5911 = (inp[10]) ? node5923 : node5912;
											assign node5912 = (inp[2]) ? node5914 : 4'b0100;
												assign node5914 = (inp[5]) ? node5920 : node5915;
													assign node5915 = (inp[15]) ? 4'b0100 : node5916;
														assign node5916 = (inp[3]) ? 4'b0100 : 4'b0110;
													assign node5920 = (inp[13]) ? 4'b0110 : 4'b0100;
											assign node5923 = (inp[15]) ? node5927 : node5924;
												assign node5924 = (inp[12]) ? 4'b0000 : 4'b0100;
												assign node5927 = (inp[12]) ? 4'b0010 : 4'b0110;
								assign node5930 = (inp[13]) ? node5964 : node5931;
									assign node5931 = (inp[15]) ? node5951 : node5932;
										assign node5932 = (inp[3]) ? node5938 : node5933;
											assign node5933 = (inp[9]) ? 4'b0010 : node5934;
												assign node5934 = (inp[4]) ? 4'b0010 : 4'b0110;
											assign node5938 = (inp[5]) ? node5942 : node5939;
												assign node5939 = (inp[9]) ? 4'b0010 : 4'b0110;
												assign node5942 = (inp[12]) ? node5948 : node5943;
													assign node5943 = (inp[9]) ? 4'b0000 : node5944;
														assign node5944 = (inp[4]) ? 4'b0000 : 4'b0100;
													assign node5948 = (inp[4]) ? 4'b0100 : 4'b0000;
										assign node5951 = (inp[2]) ? node5957 : node5952;
											assign node5952 = (inp[9]) ? 4'b0000 : node5953;
												assign node5953 = (inp[10]) ? 4'b0000 : 4'b0100;
											assign node5957 = (inp[9]) ? 4'b0110 : node5958;
												assign node5958 = (inp[12]) ? node5960 : 4'b0100;
													assign node5960 = (inp[10]) ? 4'b0100 : 4'b0000;
									assign node5964 = (inp[5]) ? node5990 : node5965;
										assign node5965 = (inp[15]) ? node5975 : node5966;
											assign node5966 = (inp[12]) ? node5968 : 4'b1110;
												assign node5968 = (inp[3]) ? node5970 : 4'b1010;
													assign node5970 = (inp[4]) ? node5972 : 4'b1010;
														assign node5972 = (inp[2]) ? 4'b1000 : 4'b1100;
											assign node5975 = (inp[12]) ? node5985 : node5976;
												assign node5976 = (inp[4]) ? node5980 : node5977;
													assign node5977 = (inp[9]) ? 4'b1110 : 4'b1100;
													assign node5980 = (inp[3]) ? 4'b1000 : node5981;
														assign node5981 = (inp[2]) ? 4'b1100 : 4'b1000;
												assign node5985 = (inp[4]) ? node5987 : 4'b1000;
													assign node5987 = (inp[9]) ? 4'b1000 : 4'b1100;
										assign node5990 = (inp[15]) ? node6006 : node5991;
											assign node5991 = (inp[4]) ? node6001 : node5992;
												assign node5992 = (inp[3]) ? node5998 : node5993;
													assign node5993 = (inp[10]) ? node5995 : 4'b1010;
														assign node5995 = (inp[9]) ? 4'b1100 : 4'b1010;
													assign node5998 = (inp[9]) ? 4'b1100 : 4'b1000;
												assign node6001 = (inp[12]) ? node6003 : 4'b1100;
													assign node6003 = (inp[9]) ? 4'b1000 : 4'b1100;
											assign node6006 = (inp[2]) ? node6014 : node6007;
												assign node6007 = (inp[4]) ? node6011 : node6008;
													assign node6008 = (inp[10]) ? 4'b1000 : 4'b1010;
													assign node6011 = (inp[9]) ? 4'b1010 : 4'b1110;
												assign node6014 = (inp[9]) ? 4'b1110 : node6015;
													assign node6015 = (inp[10]) ? 4'b1010 : node6016;
														assign node6016 = (inp[4]) ? 4'b1010 : 4'b1110;
						assign node6021 = (inp[11]) ? node6171 : node6022;
							assign node6022 = (inp[1]) ? node6102 : node6023;
								assign node6023 = (inp[2]) ? node6051 : node6024;
									assign node6024 = (inp[4]) ? node6042 : node6025;
										assign node6025 = (inp[9]) ? node6031 : node6026;
											assign node6026 = (inp[5]) ? 4'b0100 : node6027;
												assign node6027 = (inp[15]) ? 4'b0100 : 4'b0110;
											assign node6031 = (inp[10]) ? node6037 : node6032;
												assign node6032 = (inp[15]) ? node6034 : 4'b0010;
													assign node6034 = (inp[5]) ? 4'b0010 : 4'b0000;
												assign node6037 = (inp[12]) ? 4'b0100 : node6038;
													assign node6038 = (inp[15]) ? 4'b0000 : 4'b0010;
										assign node6042 = (inp[9]) ? node6044 : 4'b0010;
											assign node6044 = (inp[12]) ? node6046 : 4'b0110;
												assign node6046 = (inp[10]) ? node6048 : 4'b0110;
													assign node6048 = (inp[5]) ? 4'b0000 : 4'b0010;
									assign node6051 = (inp[10]) ? node6081 : node6052;
										assign node6052 = (inp[3]) ? node6070 : node6053;
											assign node6053 = (inp[15]) ? node6061 : node6054;
												assign node6054 = (inp[13]) ? 4'b0110 : node6055;
													assign node6055 = (inp[9]) ? 4'b0010 : node6056;
														assign node6056 = (inp[12]) ? 4'b0110 : 4'b0010;
												assign node6061 = (inp[13]) ? node6067 : node6062;
													assign node6062 = (inp[4]) ? 4'b0100 : node6063;
														assign node6063 = (inp[9]) ? 4'b0000 : 4'b0100;
													assign node6067 = (inp[12]) ? 4'b0100 : 4'b0110;
											assign node6070 = (inp[12]) ? node6072 : 4'b0100;
												assign node6072 = (inp[13]) ? node6078 : node6073;
													assign node6073 = (inp[9]) ? 4'b0110 : node6074;
														assign node6074 = (inp[5]) ? 4'b0100 : 4'b0000;
													assign node6078 = (inp[5]) ? 4'b0000 : 4'b0100;
										assign node6081 = (inp[12]) ? node6087 : node6082;
											assign node6082 = (inp[3]) ? 4'b0010 : node6083;
												assign node6083 = (inp[4]) ? 4'b0000 : 4'b0110;
											assign node6087 = (inp[15]) ? node6095 : node6088;
												assign node6088 = (inp[3]) ? 4'b0100 : node6089;
													assign node6089 = (inp[13]) ? node6091 : 4'b0100;
														assign node6091 = (inp[9]) ? 4'b0000 : 4'b0100;
												assign node6095 = (inp[3]) ? 4'b0010 : node6096;
													assign node6096 = (inp[9]) ? 4'b0110 : node6097;
														assign node6097 = (inp[4]) ? 4'b0110 : 4'b0000;
								assign node6102 = (inp[13]) ? node6136 : node6103;
									assign node6103 = (inp[15]) ? node6119 : node6104;
										assign node6104 = (inp[5]) ? node6110 : node6105;
											assign node6105 = (inp[3]) ? node6107 : 4'b0010;
												assign node6107 = (inp[4]) ? 4'b0100 : 4'b0010;
											assign node6110 = (inp[10]) ? 4'b0100 : node6111;
												assign node6111 = (inp[12]) ? 4'b0000 : node6112;
													assign node6112 = (inp[4]) ? node6114 : 4'b0100;
														assign node6114 = (inp[9]) ? 4'b0100 : 4'b0000;
										assign node6119 = (inp[4]) ? node6125 : node6120;
											assign node6120 = (inp[12]) ? node6122 : 4'b0100;
												assign node6122 = (inp[3]) ? 4'b0110 : 4'b0100;
											assign node6125 = (inp[5]) ? node6129 : node6126;
												assign node6126 = (inp[3]) ? 4'b0110 : 4'b0100;
												assign node6129 = (inp[2]) ? 4'b0010 : node6130;
													assign node6130 = (inp[3]) ? node6132 : 4'b0110;
														assign node6132 = (inp[9]) ? 4'b0010 : 4'b0010;
									assign node6136 = (inp[12]) ? node6152 : node6137;
										assign node6137 = (inp[4]) ? node6145 : node6138;
											assign node6138 = (inp[5]) ? 4'b1110 : node6139;
												assign node6139 = (inp[2]) ? node6141 : 4'b1100;
													assign node6141 = (inp[10]) ? 4'b1000 : 4'b1100;
											assign node6145 = (inp[9]) ? node6149 : node6146;
												assign node6146 = (inp[10]) ? 4'b1110 : 4'b1010;
												assign node6149 = (inp[5]) ? 4'b1100 : 4'b1000;
										assign node6152 = (inp[15]) ? node6160 : node6153;
											assign node6153 = (inp[5]) ? 4'b1000 : node6154;
												assign node6154 = (inp[3]) ? node6156 : 4'b1110;
													assign node6156 = (inp[10]) ? 4'b1010 : 4'b1000;
											assign node6160 = (inp[5]) ? node6162 : 4'b1000;
												assign node6162 = (inp[10]) ? 4'b1010 : node6163;
													assign node6163 = (inp[2]) ? node6167 : node6164;
														assign node6164 = (inp[4]) ? 4'b1010 : 4'b1110;
														assign node6167 = (inp[9]) ? 4'b1010 : 4'b1010;
							assign node6171 = (inp[13]) ? node6257 : node6172;
								assign node6172 = (inp[3]) ? node6224 : node6173;
									assign node6173 = (inp[15]) ? node6199 : node6174;
										assign node6174 = (inp[5]) ? node6188 : node6175;
											assign node6175 = (inp[2]) ? 4'b1010 : node6176;
												assign node6176 = (inp[1]) ? node6182 : node6177;
													assign node6177 = (inp[9]) ? 4'b1110 : node6178;
														assign node6178 = (inp[10]) ? 4'b1010 : 4'b1110;
													assign node6182 = (inp[10]) ? node6184 : 4'b1010;
														assign node6184 = (inp[12]) ? 4'b1110 : 4'b1010;
											assign node6188 = (inp[9]) ? node6196 : node6189;
												assign node6189 = (inp[4]) ? 4'b1100 : node6190;
													assign node6190 = (inp[12]) ? 4'b1010 : node6191;
														assign node6191 = (inp[10]) ? 4'b1010 : 4'b1110;
												assign node6196 = (inp[4]) ? 4'b1000 : 4'b1100;
										assign node6199 = (inp[5]) ? node6213 : node6200;
											assign node6200 = (inp[12]) ? node6206 : node6201;
												assign node6201 = (inp[1]) ? node6203 : 4'b1100;
													assign node6203 = (inp[9]) ? 4'b1000 : 4'b1100;
												assign node6206 = (inp[1]) ? node6208 : 4'b1000;
													assign node6208 = (inp[2]) ? 4'b1100 : node6209;
														assign node6209 = (inp[10]) ? 4'b1100 : 4'b1000;
											assign node6213 = (inp[2]) ? node6215 : 4'b1010;
												assign node6215 = (inp[10]) ? node6219 : node6216;
													assign node6216 = (inp[1]) ? 4'b1000 : 4'b1110;
													assign node6219 = (inp[9]) ? node6221 : 4'b1110;
														assign node6221 = (inp[4]) ? 4'b1010 : 4'b1110;
									assign node6224 = (inp[15]) ? node6244 : node6225;
										assign node6225 = (inp[5]) ? node6231 : node6226;
											assign node6226 = (inp[10]) ? node6228 : 4'b1100;
												assign node6228 = (inp[4]) ? 4'b1000 : 4'b1100;
											assign node6231 = (inp[1]) ? node6237 : node6232;
												assign node6232 = (inp[4]) ? node6234 : 4'b1000;
													assign node6234 = (inp[2]) ? 4'b1000 : 4'b1100;
												assign node6237 = (inp[9]) ? node6239 : 4'b1100;
													assign node6239 = (inp[4]) ? node6241 : 4'b1100;
														assign node6241 = (inp[10]) ? 4'b1000 : 4'b1000;
										assign node6244 = (inp[5]) ? node6252 : node6245;
											assign node6245 = (inp[12]) ? 4'b1110 : node6246;
												assign node6246 = (inp[10]) ? node6248 : 4'b1000;
													assign node6248 = (inp[4]) ? 4'b1110 : 4'b1000;
											assign node6252 = (inp[4]) ? 4'b1110 : node6253;
												assign node6253 = (inp[12]) ? 4'b1010 : 4'b1110;
								assign node6257 = (inp[1]) ? node6299 : node6258;
									assign node6258 = (inp[12]) ? node6276 : node6259;
										assign node6259 = (inp[4]) ? node6269 : node6260;
											assign node6260 = (inp[5]) ? 4'b1000 : node6261;
												assign node6261 = (inp[2]) ? node6263 : 4'b1110;
													assign node6263 = (inp[15]) ? 4'b1000 : node6264;
														assign node6264 = (inp[3]) ? 4'b1110 : 4'b1010;
											assign node6269 = (inp[10]) ? 4'b1000 : node6270;
												assign node6270 = (inp[3]) ? 4'b1110 : node6271;
													assign node6271 = (inp[9]) ? 4'b1100 : 4'b1000;
										assign node6276 = (inp[15]) ? node6290 : node6277;
											assign node6277 = (inp[3]) ? node6285 : node6278;
												assign node6278 = (inp[5]) ? 4'b1100 : node6279;
													assign node6279 = (inp[10]) ? 4'b1110 : node6280;
														assign node6280 = (inp[2]) ? 4'b1110 : 4'b1010;
												assign node6285 = (inp[2]) ? 4'b1000 : node6286;
													assign node6286 = (inp[4]) ? 4'b1100 : 4'b1000;
											assign node6290 = (inp[5]) ? node6292 : 4'b1000;
												assign node6292 = (inp[4]) ? node6296 : node6293;
													assign node6293 = (inp[9]) ? 4'b1110 : 4'b1010;
													assign node6296 = (inp[9]) ? 4'b1010 : 4'b1110;
									assign node6299 = (inp[4]) ? node6311 : node6300;
										assign node6300 = (inp[3]) ? node6302 : 4'b0000;
											assign node6302 = (inp[12]) ? node6308 : node6303;
												assign node6303 = (inp[5]) ? 4'b0110 : node6304;
													assign node6304 = (inp[2]) ? 4'b0000 : 4'b0010;
												assign node6308 = (inp[15]) ? 4'b0110 : 4'b0100;
										assign node6311 = (inp[9]) ? node6327 : node6312;
											assign node6312 = (inp[10]) ? node6320 : node6313;
												assign node6313 = (inp[12]) ? 4'b0100 : node6314;
													assign node6314 = (inp[5]) ? node6316 : 4'b0010;
														assign node6316 = (inp[3]) ? 4'b0010 : 4'b0000;
												assign node6320 = (inp[2]) ? node6322 : 4'b0110;
													assign node6322 = (inp[12]) ? 4'b0110 : node6323;
														assign node6323 = (inp[5]) ? 4'b0110 : 4'b0100;
											assign node6327 = (inp[12]) ? node6331 : node6328;
												assign node6328 = (inp[5]) ? 4'b0100 : 4'b0000;
												assign node6331 = (inp[5]) ? node6335 : node6332;
													assign node6332 = (inp[15]) ? 4'b0000 : 4'b0010;
													assign node6335 = (inp[15]) ? 4'b0010 : 4'b0000;
					assign node6338 = (inp[5]) ? node6702 : node6339;
						assign node6339 = (inp[15]) ? node6543 : node6340;
							assign node6340 = (inp[3]) ? node6438 : node6341;
								assign node6341 = (inp[1]) ? node6393 : node6342;
									assign node6342 = (inp[13]) ? node6362 : node6343;
										assign node6343 = (inp[11]) ? node6349 : node6344;
											assign node6344 = (inp[6]) ? 4'b0011 : node6345;
												assign node6345 = (inp[9]) ? 4'b1011 : 4'b1111;
											assign node6349 = (inp[6]) ? node6357 : node6350;
												assign node6350 = (inp[9]) ? 4'b0111 : node6351;
													assign node6351 = (inp[12]) ? node6353 : 4'b0111;
														assign node6353 = (inp[2]) ? 4'b0011 : 4'b0011;
												assign node6357 = (inp[12]) ? node6359 : 4'b1111;
													assign node6359 = (inp[10]) ? 4'b1111 : 4'b1011;
										assign node6362 = (inp[12]) ? node6378 : node6363;
											assign node6363 = (inp[2]) ? node6371 : node6364;
												assign node6364 = (inp[10]) ? node6366 : 4'b0011;
													assign node6366 = (inp[11]) ? 4'b0011 : node6367;
														assign node6367 = (inp[4]) ? 4'b0011 : 4'b0111;
												assign node6371 = (inp[6]) ? node6375 : node6372;
													assign node6372 = (inp[11]) ? 4'b1111 : 4'b0111;
													assign node6375 = (inp[9]) ? 4'b0111 : 4'b0011;
											assign node6378 = (inp[2]) ? 4'b0011 : node6379;
												assign node6379 = (inp[6]) ? node6385 : node6380;
													assign node6380 = (inp[10]) ? node6382 : 4'b1111;
														assign node6382 = (inp[9]) ? 4'b1011 : 4'b1111;
													assign node6385 = (inp[11]) ? node6389 : node6386;
														assign node6386 = (inp[4]) ? 4'b1111 : 4'b1011;
														assign node6389 = (inp[4]) ? 4'b0111 : 4'b0011;
									assign node6393 = (inp[10]) ? node6415 : node6394;
										assign node6394 = (inp[11]) ? node6402 : node6395;
											assign node6395 = (inp[6]) ? node6399 : node6396;
												assign node6396 = (inp[4]) ? 4'b0011 : 4'b0111;
												assign node6399 = (inp[12]) ? 4'b1011 : 4'b1111;
											assign node6402 = (inp[6]) ? node6408 : node6403;
												assign node6403 = (inp[12]) ? 4'b1011 : node6404;
													assign node6404 = (inp[4]) ? 4'b1111 : 4'b1011;
												assign node6408 = (inp[2]) ? node6410 : 4'b0011;
													assign node6410 = (inp[13]) ? node6412 : 4'b0011;
														assign node6412 = (inp[12]) ? 4'b0111 : 4'b0011;
										assign node6415 = (inp[9]) ? node6429 : node6416;
											assign node6416 = (inp[4]) ? node6420 : node6417;
												assign node6417 = (inp[6]) ? 4'b0011 : 4'b1011;
												assign node6420 = (inp[2]) ? node6424 : node6421;
													assign node6421 = (inp[12]) ? 4'b0111 : 4'b0011;
													assign node6424 = (inp[13]) ? node6426 : 4'b1111;
														assign node6426 = (inp[11]) ? 4'b0111 : 4'b1111;
											assign node6429 = (inp[4]) ? 4'b1011 : node6430;
												assign node6430 = (inp[12]) ? node6432 : 4'b1111;
													assign node6432 = (inp[13]) ? node6434 : 4'b0111;
														assign node6434 = (inp[11]) ? 4'b0111 : 4'b1111;
								assign node6438 = (inp[9]) ? node6488 : node6439;
									assign node6439 = (inp[4]) ? node6465 : node6440;
										assign node6440 = (inp[12]) ? node6458 : node6441;
											assign node6441 = (inp[6]) ? node6449 : node6442;
												assign node6442 = (inp[11]) ? node6444 : 4'b0111;
													assign node6444 = (inp[1]) ? 4'b1011 : node6445;
														assign node6445 = (inp[2]) ? 4'b0111 : 4'b1111;
												assign node6449 = (inp[10]) ? node6455 : node6450;
													assign node6450 = (inp[1]) ? 4'b0111 : node6451;
														assign node6451 = (inp[13]) ? 4'b0111 : 4'b1111;
													assign node6455 = (inp[11]) ? 4'b0011 : 4'b0111;
											assign node6458 = (inp[10]) ? node6460 : 4'b1011;
												assign node6460 = (inp[13]) ? 4'b0011 : node6461;
													assign node6461 = (inp[11]) ? 4'b0011 : 4'b1011;
										assign node6465 = (inp[12]) ? node6477 : node6466;
											assign node6466 = (inp[1]) ? node6472 : node6467;
												assign node6467 = (inp[11]) ? node6469 : 4'b0011;
													assign node6469 = (inp[6]) ? 4'b0101 : 4'b1101;
												assign node6472 = (inp[11]) ? node6474 : 4'b0011;
													assign node6474 = (inp[6]) ? 4'b0011 : 4'b1011;
											assign node6477 = (inp[13]) ? node6483 : node6478;
												assign node6478 = (inp[2]) ? node6480 : 4'b0011;
													assign node6480 = (inp[10]) ? 4'b1101 : 4'b0101;
												assign node6483 = (inp[10]) ? node6485 : 4'b1101;
													assign node6485 = (inp[6]) ? 4'b0101 : 4'b1101;
									assign node6488 = (inp[2]) ? node6518 : node6489;
										assign node6489 = (inp[10]) ? node6503 : node6490;
											assign node6490 = (inp[11]) ? node6496 : node6491;
												assign node6491 = (inp[4]) ? node6493 : 4'b0011;
													assign node6493 = (inp[13]) ? 4'b1101 : 4'b0101;
												assign node6496 = (inp[1]) ? node6498 : 4'b1101;
													assign node6498 = (inp[4]) ? node6500 : 4'b1011;
														assign node6500 = (inp[13]) ? 4'b1001 : 4'b1101;
											assign node6503 = (inp[12]) ? node6515 : node6504;
												assign node6504 = (inp[1]) ? node6510 : node6505;
													assign node6505 = (inp[4]) ? node6507 : 4'b0011;
														assign node6507 = (inp[13]) ? 4'b0101 : 4'b1101;
													assign node6510 = (inp[13]) ? node6512 : 4'b0101;
														assign node6512 = (inp[11]) ? 4'b0101 : 4'b1101;
												assign node6515 = (inp[6]) ? 4'b0101 : 4'b1101;
										assign node6518 = (inp[4]) ? node6530 : node6519;
											assign node6519 = (inp[12]) ? node6523 : node6520;
												assign node6520 = (inp[6]) ? 4'b1011 : 4'b0011;
												assign node6523 = (inp[1]) ? 4'b1101 : node6524;
													assign node6524 = (inp[6]) ? 4'b1101 : node6525;
														assign node6525 = (inp[13]) ? 4'b0101 : 4'b0011;
											assign node6530 = (inp[6]) ? node6538 : node6531;
												assign node6531 = (inp[12]) ? node6533 : 4'b1101;
													assign node6533 = (inp[11]) ? 4'b1001 : node6534;
														assign node6534 = (inp[13]) ? 4'b0001 : 4'b1001;
												assign node6538 = (inp[13]) ? 4'b0001 : node6539;
													assign node6539 = (inp[1]) ? 4'b0001 : 4'b1001;
							assign node6543 = (inp[3]) ? node6623 : node6544;
								assign node6544 = (inp[13]) ? node6584 : node6545;
									assign node6545 = (inp[11]) ? node6557 : node6546;
										assign node6546 = (inp[6]) ? node6552 : node6547;
											assign node6547 = (inp[1]) ? node6549 : 4'b1101;
												assign node6549 = (inp[12]) ? 4'b0101 : 4'b0001;
											assign node6552 = (inp[1]) ? 4'b1001 : node6553;
												assign node6553 = (inp[2]) ? 4'b0001 : 4'b0101;
										assign node6557 = (inp[9]) ? node6569 : node6558;
											assign node6558 = (inp[1]) ? node6564 : node6559;
												assign node6559 = (inp[6]) ? 4'b1101 : node6560;
													assign node6560 = (inp[12]) ? 4'b0101 : 4'b0001;
												assign node6564 = (inp[4]) ? node6566 : 4'b0001;
													assign node6566 = (inp[12]) ? 4'b0101 : 4'b0001;
											assign node6569 = (inp[12]) ? node6575 : node6570;
												assign node6570 = (inp[10]) ? 4'b0101 : node6571;
													assign node6571 = (inp[1]) ? 4'b0101 : 4'b1101;
												assign node6575 = (inp[4]) ? node6581 : node6576;
													assign node6576 = (inp[2]) ? 4'b1101 : node6577;
														assign node6577 = (inp[6]) ? 4'b1101 : 4'b0001;
													assign node6581 = (inp[6]) ? 4'b0001 : 4'b0101;
									assign node6584 = (inp[11]) ? node6606 : node6585;
										assign node6585 = (inp[6]) ? node6597 : node6586;
											assign node6586 = (inp[4]) ? node6592 : node6587;
												assign node6587 = (inp[12]) ? 4'b0101 : node6588;
													assign node6588 = (inp[2]) ? 4'b0101 : 4'b0001;
												assign node6592 = (inp[2]) ? node6594 : 4'b0001;
													assign node6594 = (inp[12]) ? 4'b0001 : 4'b0101;
											assign node6597 = (inp[9]) ? node6601 : node6598;
												assign node6598 = (inp[4]) ? 4'b1101 : 4'b1001;
												assign node6601 = (inp[4]) ? node6603 : 4'b1101;
													assign node6603 = (inp[2]) ? 4'b1101 : 4'b1001;
										assign node6606 = (inp[6]) ? node6618 : node6607;
											assign node6607 = (inp[12]) ? node6609 : 4'b1101;
												assign node6609 = (inp[10]) ? node6615 : node6610;
													assign node6610 = (inp[2]) ? 4'b1101 : node6611;
														assign node6611 = (inp[1]) ? 4'b1001 : 4'b1001;
													assign node6615 = (inp[2]) ? 4'b1001 : 4'b1101;
											assign node6618 = (inp[10]) ? node6620 : 4'b0101;
												assign node6620 = (inp[4]) ? 4'b0001 : 4'b0101;
								assign node6623 = (inp[4]) ? node6655 : node6624;
									assign node6624 = (inp[9]) ? node6638 : node6625;
										assign node6625 = (inp[6]) ? node6633 : node6626;
											assign node6626 = (inp[10]) ? node6630 : node6627;
												assign node6627 = (inp[2]) ? 4'b0101 : 4'b1101;
												assign node6630 = (inp[2]) ? 4'b0001 : 4'b0101;
											assign node6633 = (inp[13]) ? node6635 : 4'b0101;
												assign node6635 = (inp[11]) ? 4'b0001 : 4'b1001;
										assign node6638 = (inp[10]) ? node6650 : node6639;
											assign node6639 = (inp[12]) ? node6645 : node6640;
												assign node6640 = (inp[1]) ? 4'b0001 : node6641;
													assign node6641 = (inp[6]) ? 4'b0001 : 4'b1001;
												assign node6645 = (inp[11]) ? 4'b1111 : node6646;
													assign node6646 = (inp[6]) ? 4'b1111 : 4'b0001;
											assign node6650 = (inp[12]) ? 4'b0111 : node6651;
												assign node6651 = (inp[1]) ? 4'b0111 : 4'b1111;
									assign node6655 = (inp[9]) ? node6677 : node6656;
										assign node6656 = (inp[10]) ? node6674 : node6657;
											assign node6657 = (inp[12]) ? node6663 : node6658;
												assign node6658 = (inp[13]) ? 4'b0001 : node6659;
													assign node6659 = (inp[1]) ? 4'b1001 : 4'b0001;
												assign node6663 = (inp[6]) ? node6669 : node6664;
													assign node6664 = (inp[2]) ? 4'b0001 : node6665;
														assign node6665 = (inp[11]) ? 4'b1111 : 4'b0001;
													assign node6669 = (inp[11]) ? node6671 : 4'b1111;
														assign node6671 = (inp[13]) ? 4'b0111 : 4'b1111;
											assign node6674 = (inp[13]) ? 4'b1111 : 4'b0111;
										assign node6677 = (inp[10]) ? node6689 : node6678;
											assign node6678 = (inp[11]) ? node6686 : node6679;
												assign node6679 = (inp[2]) ? 4'b0111 : node6680;
													assign node6680 = (inp[1]) ? 4'b1011 : node6681;
														assign node6681 = (inp[13]) ? 4'b1111 : 4'b0111;
												assign node6686 = (inp[6]) ? 4'b0011 : 4'b1011;
											assign node6689 = (inp[12]) ? 4'b1011 : node6690;
												assign node6690 = (inp[2]) ? node6698 : node6691;
													assign node6691 = (inp[13]) ? node6695 : node6692;
														assign node6692 = (inp[6]) ? 4'b1011 : 4'b1111;
														assign node6695 = (inp[1]) ? 4'b1011 : 4'b0011;
													assign node6698 = (inp[6]) ? 4'b0011 : 4'b0111;
						assign node6702 = (inp[15]) ? node6880 : node6703;
							assign node6703 = (inp[3]) ? node6789 : node6704;
								assign node6704 = (inp[9]) ? node6742 : node6705;
									assign node6705 = (inp[4]) ? node6723 : node6706;
										assign node6706 = (inp[6]) ? node6714 : node6707;
											assign node6707 = (inp[10]) ? 4'b0011 : node6708;
												assign node6708 = (inp[11]) ? node6710 : 4'b0111;
													assign node6710 = (inp[13]) ? 4'b1111 : 4'b0111;
											assign node6714 = (inp[2]) ? 4'b1011 : node6715;
												assign node6715 = (inp[12]) ? node6717 : 4'b1011;
													assign node6717 = (inp[10]) ? node6719 : 4'b0011;
														assign node6719 = (inp[11]) ? 4'b1011 : 4'b0011;
										assign node6723 = (inp[10]) ? node6735 : node6724;
											assign node6724 = (inp[12]) ? node6728 : node6725;
												assign node6725 = (inp[2]) ? 4'b0011 : 4'b1011;
												assign node6728 = (inp[13]) ? node6732 : node6729;
													assign node6729 = (inp[6]) ? 4'b1101 : 4'b0011;
													assign node6732 = (inp[1]) ? 4'b0101 : 4'b1101;
											assign node6735 = (inp[11]) ? node6739 : node6736;
												assign node6736 = (inp[6]) ? 4'b1101 : 4'b0101;
												assign node6739 = (inp[6]) ? 4'b0101 : 4'b1101;
									assign node6742 = (inp[4]) ? node6772 : node6743;
										assign node6743 = (inp[10]) ? node6751 : node6744;
											assign node6744 = (inp[12]) ? node6746 : 4'b0011;
												assign node6746 = (inp[6]) ? node6748 : 4'b1011;
													assign node6748 = (inp[13]) ? 4'b1101 : 4'b0101;
											assign node6751 = (inp[12]) ? node6757 : node6752;
												assign node6752 = (inp[11]) ? node6754 : 4'b1101;
													assign node6754 = (inp[6]) ? 4'b0101 : 4'b1101;
												assign node6757 = (inp[2]) ? node6765 : node6758;
													assign node6758 = (inp[1]) ? node6762 : node6759;
														assign node6759 = (inp[11]) ? 4'b0101 : 4'b1101;
														assign node6762 = (inp[11]) ? 4'b1101 : 4'b0101;
													assign node6765 = (inp[13]) ? node6769 : node6766;
														assign node6766 = (inp[11]) ? 4'b0101 : 4'b1101;
														assign node6769 = (inp[11]) ? 4'b1101 : 4'b0101;
										assign node6772 = (inp[10]) ? node6778 : node6773;
											assign node6773 = (inp[11]) ? node6775 : 4'b0101;
												assign node6775 = (inp[12]) ? 4'b1001 : 4'b1101;
											assign node6778 = (inp[13]) ? node6780 : 4'b1001;
												assign node6780 = (inp[1]) ? node6786 : node6781;
													assign node6781 = (inp[6]) ? 4'b0001 : node6782;
														assign node6782 = (inp[11]) ? 4'b1001 : 4'b0001;
													assign node6786 = (inp[2]) ? 4'b1001 : 4'b0101;
								assign node6789 = (inp[6]) ? node6835 : node6790;
									assign node6790 = (inp[11]) ? node6810 : node6791;
										assign node6791 = (inp[13]) ? node6803 : node6792;
											assign node6792 = (inp[1]) ? node6796 : node6793;
												assign node6793 = (inp[10]) ? 4'b1101 : 4'b1001;
												assign node6796 = (inp[10]) ? node6798 : 4'b0101;
													assign node6798 = (inp[4]) ? 4'b0001 : node6799;
														assign node6799 = (inp[2]) ? 4'b0101 : 4'b0001;
											assign node6803 = (inp[9]) ? 4'b0001 : node6804;
												assign node6804 = (inp[2]) ? node6806 : 4'b0001;
													assign node6806 = (inp[10]) ? 4'b0101 : 4'b0001;
										assign node6810 = (inp[1]) ? node6824 : node6811;
											assign node6811 = (inp[13]) ? node6819 : node6812;
												assign node6812 = (inp[4]) ? node6814 : 4'b0101;
													assign node6814 = (inp[2]) ? 4'b0001 : node6815;
														assign node6815 = (inp[12]) ? 4'b0001 : 4'b0001;
												assign node6819 = (inp[10]) ? 4'b1001 : node6820;
													assign node6820 = (inp[4]) ? 4'b1101 : 4'b1001;
											assign node6824 = (inp[4]) ? node6828 : node6825;
												assign node6825 = (inp[9]) ? 4'b1101 : 4'b1001;
												assign node6828 = (inp[9]) ? node6830 : 4'b1101;
													assign node6830 = (inp[2]) ? 4'b1001 : node6831;
														assign node6831 = (inp[13]) ? 4'b1001 : 4'b1001;
									assign node6835 = (inp[11]) ? node6863 : node6836;
										assign node6836 = (inp[1]) ? node6850 : node6837;
											assign node6837 = (inp[13]) ? node6845 : node6838;
												assign node6838 = (inp[9]) ? node6840 : 4'b0001;
													assign node6840 = (inp[12]) ? node6842 : 4'b0001;
														assign node6842 = (inp[10]) ? 4'b0001 : 4'b0101;
												assign node6845 = (inp[12]) ? 4'b1101 : node6846;
													assign node6846 = (inp[9]) ? 4'b1101 : 4'b1001;
											assign node6850 = (inp[4]) ? node6860 : node6851;
												assign node6851 = (inp[2]) ? node6855 : node6852;
													assign node6852 = (inp[12]) ? 4'b1001 : 4'b1101;
													assign node6855 = (inp[10]) ? node6857 : 4'b1001;
														assign node6857 = (inp[12]) ? 4'b1101 : 4'b1001;
												assign node6860 = (inp[2]) ? 4'b1101 : 4'b1001;
										assign node6863 = (inp[13]) ? node6869 : node6864;
											assign node6864 = (inp[1]) ? node6866 : 4'b1101;
												assign node6866 = (inp[12]) ? 4'b0101 : 4'b0001;
											assign node6869 = (inp[1]) ? 4'b0101 : node6870;
												assign node6870 = (inp[12]) ? node6872 : 4'b0101;
													assign node6872 = (inp[2]) ? node6876 : node6873;
														assign node6873 = (inp[9]) ? 4'b0101 : 4'b0001;
														assign node6876 = (inp[9]) ? 4'b0001 : 4'b0101;
							assign node6880 = (inp[3]) ? node6956 : node6881;
								assign node6881 = (inp[9]) ? node6919 : node6882;
									assign node6882 = (inp[10]) ? node6902 : node6883;
										assign node6883 = (inp[4]) ? node6891 : node6884;
											assign node6884 = (inp[13]) ? node6886 : 4'b0101;
												assign node6886 = (inp[12]) ? 4'b0101 : node6887;
													assign node6887 = (inp[6]) ? 4'b0101 : 4'b1101;
											assign node6891 = (inp[12]) ? node6899 : node6892;
												assign node6892 = (inp[2]) ? 4'b1001 : node6893;
													assign node6893 = (inp[13]) ? 4'b0001 : node6894;
														assign node6894 = (inp[11]) ? 4'b1001 : 4'b0001;
												assign node6899 = (inp[6]) ? 4'b0111 : 4'b0001;
										assign node6902 = (inp[4]) ? node6912 : node6903;
											assign node6903 = (inp[6]) ? node6909 : node6904;
												assign node6904 = (inp[11]) ? 4'b1001 : node6905;
													assign node6905 = (inp[2]) ? 4'b1001 : 4'b0001;
												assign node6909 = (inp[11]) ? 4'b0001 : 4'b1001;
											assign node6912 = (inp[1]) ? node6916 : node6913;
												assign node6913 = (inp[2]) ? 4'b0111 : 4'b0001;
												assign node6916 = (inp[12]) ? 4'b0111 : 4'b1111;
									assign node6919 = (inp[1]) ? node6941 : node6920;
										assign node6920 = (inp[12]) ? node6932 : node6921;
											assign node6921 = (inp[4]) ? node6925 : node6922;
												assign node6922 = (inp[2]) ? 4'b1111 : 4'b0001;
												assign node6925 = (inp[11]) ? 4'b1111 : node6926;
													assign node6926 = (inp[10]) ? 4'b1111 : node6927;
														assign node6927 = (inp[13]) ? 4'b0111 : 4'b0111;
											assign node6932 = (inp[4]) ? node6938 : node6933;
												assign node6933 = (inp[13]) ? 4'b1111 : node6934;
													assign node6934 = (inp[10]) ? 4'b1111 : 4'b0001;
												assign node6938 = (inp[2]) ? 4'b1011 : 4'b1111;
										assign node6941 = (inp[12]) ? node6951 : node6942;
											assign node6942 = (inp[11]) ? node6948 : node6943;
												assign node6943 = (inp[6]) ? node6945 : 4'b0001;
													assign node6945 = (inp[10]) ? 4'b1111 : 4'b1001;
												assign node6948 = (inp[6]) ? 4'b0111 : 4'b1111;
											assign node6951 = (inp[4]) ? node6953 : 4'b0111;
												assign node6953 = (inp[10]) ? 4'b0011 : 4'b0111;
								assign node6956 = (inp[11]) ? node7000 : node6957;
									assign node6957 = (inp[1]) ? node6987 : node6958;
										assign node6958 = (inp[10]) ? node6972 : node6959;
											assign node6959 = (inp[4]) ? node6969 : node6960;
												assign node6960 = (inp[12]) ? node6964 : node6961;
													assign node6961 = (inp[9]) ? 4'b0011 : 4'b0111;
													assign node6964 = (inp[13]) ? node6966 : 4'b0011;
														assign node6966 = (inp[9]) ? 4'b1111 : 4'b1011;
												assign node6969 = (inp[12]) ? 4'b1011 : 4'b1111;
											assign node6972 = (inp[9]) ? node6974 : 4'b0011;
												assign node6974 = (inp[2]) ? node6980 : node6975;
													assign node6975 = (inp[4]) ? 4'b0111 : node6976;
														assign node6976 = (inp[12]) ? 4'b1111 : 4'b1011;
													assign node6980 = (inp[12]) ? node6984 : node6981;
														assign node6981 = (inp[4]) ? 4'b0111 : 4'b0011;
														assign node6984 = (inp[4]) ? 4'b0011 : 4'b0111;
										assign node6987 = (inp[6]) ? node6997 : node6988;
											assign node6988 = (inp[2]) ? node6990 : 4'b0111;
												assign node6990 = (inp[10]) ? node6992 : 4'b0111;
													assign node6992 = (inp[9]) ? 4'b0011 : node6993;
														assign node6993 = (inp[12]) ? 4'b0111 : 4'b0011;
											assign node6997 = (inp[9]) ? 4'b1111 : 4'b1011;
									assign node7000 = (inp[6]) ? node7020 : node7001;
										assign node7001 = (inp[13]) ? node7011 : node7002;
											assign node7002 = (inp[1]) ? node7008 : node7003;
												assign node7003 = (inp[10]) ? node7005 : 4'b0111;
													assign node7005 = (inp[4]) ? 4'b0111 : 4'b0011;
												assign node7008 = (inp[10]) ? 4'b1111 : 4'b1011;
											assign node7011 = (inp[2]) ? 4'b1011 : node7012;
												assign node7012 = (inp[9]) ? 4'b1011 : node7013;
													assign node7013 = (inp[1]) ? node7015 : 4'b1111;
														assign node7015 = (inp[4]) ? 4'b1111 : 4'b1011;
										assign node7020 = (inp[1]) ? node7028 : node7021;
											assign node7021 = (inp[13]) ? 4'b0011 : node7022;
												assign node7022 = (inp[9]) ? node7024 : 4'b1011;
													assign node7024 = (inp[4]) ? 4'b1011 : 4'b1111;
											assign node7028 = (inp[12]) ? 4'b0011 : node7029;
												assign node7029 = (inp[10]) ? node7031 : 4'b0111;
													assign node7031 = (inp[2]) ? 4'b0011 : 4'b0111;
				assign node7035 = (inp[8]) ? node7635 : node7036;
					assign node7036 = (inp[12]) ? node7348 : node7037;
						assign node7037 = (inp[15]) ? node7203 : node7038;
							assign node7038 = (inp[5]) ? node7126 : node7039;
								assign node7039 = (inp[3]) ? node7089 : node7040;
									assign node7040 = (inp[10]) ? node7066 : node7041;
										assign node7041 = (inp[6]) ? node7059 : node7042;
											assign node7042 = (inp[11]) ? node7048 : node7043;
												assign node7043 = (inp[4]) ? 4'b1111 : node7044;
													assign node7044 = (inp[9]) ? 4'b0011 : 4'b0111;
												assign node7048 = (inp[1]) ? node7054 : node7049;
													assign node7049 = (inp[4]) ? node7051 : 4'b1111;
														assign node7051 = (inp[2]) ? 4'b0011 : 4'b1011;
													assign node7054 = (inp[9]) ? node7056 : 4'b1011;
														assign node7056 = (inp[4]) ? 4'b1111 : 4'b1011;
											assign node7059 = (inp[13]) ? 4'b1011 : node7060;
												assign node7060 = (inp[1]) ? 4'b0011 : node7061;
													assign node7061 = (inp[11]) ? 4'b1011 : 4'b0011;
										assign node7066 = (inp[4]) ? node7086 : node7067;
											assign node7067 = (inp[2]) ? node7075 : node7068;
												assign node7068 = (inp[1]) ? node7070 : 4'b0011;
													assign node7070 = (inp[9]) ? 4'b1111 : node7071;
														assign node7071 = (inp[13]) ? 4'b0011 : 4'b1011;
												assign node7075 = (inp[9]) ? node7081 : node7076;
													assign node7076 = (inp[11]) ? node7078 : 4'b0111;
														assign node7078 = (inp[1]) ? 4'b0011 : 4'b0111;
													assign node7081 = (inp[6]) ? node7083 : 4'b1111;
														assign node7083 = (inp[1]) ? 4'b0111 : 4'b1111;
											assign node7086 = (inp[1]) ? 4'b0111 : 4'b1111;
									assign node7089 = (inp[9]) ? node7111 : node7090;
										assign node7090 = (inp[10]) ? node7098 : node7091;
											assign node7091 = (inp[4]) ? node7093 : 4'b1111;
												assign node7093 = (inp[6]) ? node7095 : 4'b1011;
													assign node7095 = (inp[13]) ? 4'b1011 : 4'b0011;
											assign node7098 = (inp[4]) ? node7106 : node7099;
												assign node7099 = (inp[1]) ? node7101 : 4'b0111;
													assign node7101 = (inp[2]) ? 4'b1011 : node7102;
														assign node7102 = (inp[11]) ? 4'b0011 : 4'b0111;
												assign node7106 = (inp[1]) ? 4'b1101 : node7107;
													assign node7107 = (inp[6]) ? 4'b0101 : 4'b0011;
										assign node7111 = (inp[2]) ? node7115 : node7112;
											assign node7112 = (inp[11]) ? 4'b1101 : 4'b1011;
											assign node7115 = (inp[11]) ? node7119 : node7116;
												assign node7116 = (inp[4]) ? 4'b0101 : 4'b0011;
												assign node7119 = (inp[13]) ? node7121 : 4'b0001;
													assign node7121 = (inp[4]) ? node7123 : 4'b0101;
														assign node7123 = (inp[10]) ? 4'b0001 : 4'b0101;
								assign node7126 = (inp[3]) ? node7156 : node7127;
									assign node7127 = (inp[9]) ? node7139 : node7128;
										assign node7128 = (inp[11]) ? node7134 : node7129;
											assign node7129 = (inp[6]) ? 4'b1011 : node7130;
												assign node7130 = (inp[4]) ? 4'b0011 : 4'b0111;
											assign node7134 = (inp[4]) ? node7136 : 4'b1011;
												assign node7136 = (inp[6]) ? 4'b0101 : 4'b1101;
										assign node7139 = (inp[4]) ? node7143 : node7140;
											assign node7140 = (inp[10]) ? 4'b1101 : 4'b1011;
											assign node7143 = (inp[2]) ? node7151 : node7144;
												assign node7144 = (inp[10]) ? node7146 : 4'b0101;
													assign node7146 = (inp[1]) ? 4'b0101 : node7147;
														assign node7147 = (inp[6]) ? 4'b0101 : 4'b1101;
												assign node7151 = (inp[11]) ? node7153 : 4'b1001;
													assign node7153 = (inp[6]) ? 4'b0101 : 4'b1101;
									assign node7156 = (inp[2]) ? node7180 : node7157;
										assign node7157 = (inp[13]) ? node7169 : node7158;
											assign node7158 = (inp[4]) ? node7164 : node7159;
												assign node7159 = (inp[1]) ? node7161 : 4'b0101;
													assign node7161 = (inp[11]) ? 4'b1001 : 4'b0001;
												assign node7164 = (inp[6]) ? node7166 : 4'b1001;
													assign node7166 = (inp[1]) ? 4'b1001 : 4'b0001;
											assign node7169 = (inp[6]) ? 4'b0001 : node7170;
												assign node7170 = (inp[11]) ? node7176 : node7171;
													assign node7171 = (inp[9]) ? node7173 : 4'b0001;
														assign node7173 = (inp[4]) ? 4'b0101 : 4'b0001;
													assign node7176 = (inp[9]) ? 4'b1001 : 4'b1101;
										assign node7180 = (inp[11]) ? node7194 : node7181;
											assign node7181 = (inp[4]) ? node7189 : node7182;
												assign node7182 = (inp[9]) ? node7184 : 4'b1101;
													assign node7184 = (inp[6]) ? node7186 : 4'b0001;
														assign node7186 = (inp[10]) ? 4'b1101 : 4'b1001;
												assign node7189 = (inp[9]) ? 4'b0101 : node7190;
													assign node7190 = (inp[6]) ? 4'b0001 : 4'b1001;
											assign node7194 = (inp[1]) ? 4'b0101 : node7195;
												assign node7195 = (inp[4]) ? node7197 : 4'b0001;
													assign node7197 = (inp[9]) ? 4'b0101 : node7198;
														assign node7198 = (inp[6]) ? 4'b0101 : 4'b0001;
							assign node7203 = (inp[3]) ? node7281 : node7204;
								assign node7204 = (inp[5]) ? node7244 : node7205;
									assign node7205 = (inp[11]) ? node7219 : node7206;
										assign node7206 = (inp[9]) ? node7210 : node7207;
											assign node7207 = (inp[13]) ? 4'b0101 : 4'b1101;
											assign node7210 = (inp[1]) ? node7212 : 4'b1001;
												assign node7212 = (inp[2]) ? node7214 : 4'b1001;
													assign node7214 = (inp[4]) ? node7216 : 4'b1101;
														assign node7216 = (inp[13]) ? 4'b1101 : 4'b1001;
										assign node7219 = (inp[4]) ? node7233 : node7220;
											assign node7220 = (inp[2]) ? node7226 : node7221;
												assign node7221 = (inp[10]) ? node7223 : 4'b0101;
													assign node7223 = (inp[9]) ? 4'b0001 : 4'b1001;
												assign node7226 = (inp[1]) ? 4'b0101 : node7227;
													assign node7227 = (inp[9]) ? 4'b1001 : node7228;
														assign node7228 = (inp[13]) ? 4'b1101 : 4'b0101;
											assign node7233 = (inp[9]) ? node7241 : node7234;
												assign node7234 = (inp[10]) ? 4'b1101 : node7235;
													assign node7235 = (inp[1]) ? 4'b1001 : node7236;
														assign node7236 = (inp[2]) ? 4'b0001 : 4'b1001;
												assign node7241 = (inp[6]) ? 4'b0101 : 4'b1101;
									assign node7244 = (inp[9]) ? node7258 : node7245;
										assign node7245 = (inp[4]) ? node7253 : node7246;
											assign node7246 = (inp[13]) ? node7250 : node7247;
												assign node7247 = (inp[11]) ? 4'b1001 : 4'b1101;
												assign node7250 = (inp[1]) ? 4'b0101 : 4'b1101;
											assign node7253 = (inp[6]) ? 4'b1111 : node7254;
												assign node7254 = (inp[11]) ? 4'b1001 : 4'b0001;
										assign node7258 = (inp[4]) ? node7268 : node7259;
											assign node7259 = (inp[1]) ? node7261 : 4'b0001;
												assign node7261 = (inp[10]) ? 4'b1111 : node7262;
													assign node7262 = (inp[2]) ? 4'b1001 : node7263;
														assign node7263 = (inp[13]) ? 4'b1001 : 4'b0001;
											assign node7268 = (inp[11]) ? node7276 : node7269;
												assign node7269 = (inp[10]) ? 4'b0111 : node7270;
													assign node7270 = (inp[6]) ? 4'b1111 : node7271;
														assign node7271 = (inp[1]) ? 4'b0111 : 4'b1111;
												assign node7276 = (inp[13]) ? node7278 : 4'b1011;
													assign node7278 = (inp[2]) ? 4'b1011 : 4'b0011;
								assign node7281 = (inp[5]) ? node7327 : node7282;
									assign node7282 = (inp[9]) ? node7310 : node7283;
										assign node7283 = (inp[10]) ? node7293 : node7284;
											assign node7284 = (inp[4]) ? node7288 : node7285;
												assign node7285 = (inp[1]) ? 4'b1101 : 4'b0101;
												assign node7288 = (inp[11]) ? node7290 : 4'b1001;
													assign node7290 = (inp[6]) ? 4'b0001 : 4'b1001;
											assign node7293 = (inp[6]) ? node7301 : node7294;
												assign node7294 = (inp[4]) ? 4'b0001 : node7295;
													assign node7295 = (inp[11]) ? node7297 : 4'b0101;
														assign node7297 = (inp[13]) ? 4'b1001 : 4'b0101;
												assign node7301 = (inp[4]) ? node7305 : node7302;
													assign node7302 = (inp[11]) ? 4'b0001 : 4'b0101;
													assign node7305 = (inp[11]) ? node7307 : 4'b1111;
														assign node7307 = (inp[1]) ? 4'b0111 : 4'b0111;
										assign node7310 = (inp[4]) ? node7314 : node7311;
											assign node7311 = (inp[11]) ? 4'b0001 : 4'b1111;
											assign node7314 = (inp[6]) ? node7322 : node7315;
												assign node7315 = (inp[13]) ? node7319 : node7316;
													assign node7316 = (inp[1]) ? 4'b1011 : 4'b1111;
													assign node7319 = (inp[11]) ? 4'b1111 : 4'b0111;
												assign node7322 = (inp[2]) ? node7324 : 4'b0111;
													assign node7324 = (inp[13]) ? 4'b1111 : 4'b0111;
									assign node7327 = (inp[6]) ? node7341 : node7328;
										assign node7328 = (inp[4]) ? node7338 : node7329;
											assign node7329 = (inp[1]) ? node7333 : node7330;
												assign node7330 = (inp[10]) ? 4'b1111 : 4'b0111;
												assign node7333 = (inp[13]) ? node7335 : 4'b1111;
													assign node7335 = (inp[9]) ? 4'b1011 : 4'b1111;
											assign node7338 = (inp[9]) ? 4'b1111 : 4'b1011;
										assign node7341 = (inp[11]) ? 4'b0011 : node7342;
											assign node7342 = (inp[2]) ? node7344 : 4'b1011;
												assign node7344 = (inp[1]) ? 4'b1111 : 4'b1011;
						assign node7348 = (inp[15]) ? node7486 : node7349;
							assign node7349 = (inp[5]) ? node7421 : node7350;
								assign node7350 = (inp[3]) ? node7386 : node7351;
									assign node7351 = (inp[1]) ? node7375 : node7352;
										assign node7352 = (inp[2]) ? node7370 : node7353;
											assign node7353 = (inp[13]) ? node7367 : node7354;
												assign node7354 = (inp[4]) ? node7360 : node7355;
													assign node7355 = (inp[6]) ? node7357 : 4'b1111;
														assign node7357 = (inp[11]) ? 4'b1011 : 4'b0011;
													assign node7360 = (inp[6]) ? node7364 : node7361;
														assign node7361 = (inp[9]) ? 4'b0011 : 4'b0111;
														assign node7364 = (inp[11]) ? 4'b1111 : 4'b0011;
												assign node7367 = (inp[11]) ? 4'b0011 : 4'b1011;
											assign node7370 = (inp[10]) ? node7372 : 4'b0111;
												assign node7372 = (inp[11]) ? 4'b0111 : 4'b1111;
										assign node7375 = (inp[11]) ? node7383 : node7376;
											assign node7376 = (inp[6]) ? node7380 : node7377;
												assign node7377 = (inp[2]) ? 4'b0011 : 4'b0111;
												assign node7380 = (inp[9]) ? 4'b1011 : 4'b1111;
											assign node7383 = (inp[6]) ? 4'b0011 : 4'b1011;
									assign node7386 = (inp[4]) ? node7406 : node7387;
										assign node7387 = (inp[9]) ? node7399 : node7388;
											assign node7388 = (inp[10]) ? node7392 : node7389;
												assign node7389 = (inp[11]) ? 4'b0011 : 4'b0111;
												assign node7392 = (inp[13]) ? node7394 : 4'b1011;
													assign node7394 = (inp[11]) ? 4'b1011 : node7395;
														assign node7395 = (inp[6]) ? 4'b1011 : 4'b0011;
											assign node7399 = (inp[6]) ? node7401 : 4'b0011;
												assign node7401 = (inp[10]) ? 4'b0101 : node7402;
													assign node7402 = (inp[2]) ? 4'b0101 : 4'b1101;
										assign node7406 = (inp[9]) ? node7414 : node7407;
											assign node7407 = (inp[13]) ? node7409 : 4'b1101;
												assign node7409 = (inp[6]) ? node7411 : 4'b1101;
													assign node7411 = (inp[2]) ? 4'b1101 : 4'b0101;
											assign node7414 = (inp[6]) ? node7416 : 4'b1001;
												assign node7416 = (inp[2]) ? 4'b0001 : node7417;
													assign node7417 = (inp[11]) ? 4'b1001 : 4'b0001;
								assign node7421 = (inp[4]) ? node7453 : node7422;
									assign node7422 = (inp[3]) ? node7436 : node7423;
										assign node7423 = (inp[9]) ? node7431 : node7424;
											assign node7424 = (inp[11]) ? node7428 : node7425;
												assign node7425 = (inp[10]) ? 4'b0011 : 4'b0111;
												assign node7428 = (inp[6]) ? 4'b0011 : 4'b1011;
											assign node7431 = (inp[10]) ? 4'b0101 : node7432;
												assign node7432 = (inp[2]) ? 4'b1011 : 4'b0011;
										assign node7436 = (inp[9]) ? node7450 : node7437;
											assign node7437 = (inp[10]) ? node7445 : node7438;
												assign node7438 = (inp[11]) ? node7440 : 4'b1101;
													assign node7440 = (inp[1]) ? 4'b1001 : node7441;
														assign node7441 = (inp[6]) ? 4'b0001 : 4'b0101;
												assign node7445 = (inp[1]) ? node7447 : 4'b0001;
													assign node7447 = (inp[13]) ? 4'b1001 : 4'b0001;
											assign node7450 = (inp[13]) ? 4'b0101 : 4'b1101;
									assign node7453 = (inp[9]) ? node7469 : node7454;
										assign node7454 = (inp[2]) ? node7462 : node7455;
											assign node7455 = (inp[13]) ? node7457 : 4'b1101;
												assign node7457 = (inp[10]) ? node7459 : 4'b1101;
													assign node7459 = (inp[11]) ? 4'b1101 : 4'b0101;
											assign node7462 = (inp[3]) ? node7464 : 4'b0101;
												assign node7464 = (inp[6]) ? node7466 : 4'b1101;
													assign node7466 = (inp[1]) ? 4'b0101 : 4'b1101;
										assign node7469 = (inp[10]) ? node7477 : node7470;
											assign node7470 = (inp[13]) ? 4'b1001 : node7471;
												assign node7471 = (inp[11]) ? 4'b0101 : node7472;
													assign node7472 = (inp[6]) ? 4'b0101 : 4'b1101;
											assign node7477 = (inp[6]) ? node7481 : node7478;
												assign node7478 = (inp[11]) ? 4'b1001 : 4'b0001;
												assign node7481 = (inp[11]) ? 4'b0001 : node7482;
													assign node7482 = (inp[13]) ? 4'b1001 : 4'b0001;
							assign node7486 = (inp[5]) ? node7570 : node7487;
								assign node7487 = (inp[3]) ? node7519 : node7488;
									assign node7488 = (inp[9]) ? node7504 : node7489;
										assign node7489 = (inp[4]) ? node7495 : node7490;
											assign node7490 = (inp[1]) ? 4'b1001 : node7491;
												assign node7491 = (inp[11]) ? 4'b0001 : 4'b0101;
											assign node7495 = (inp[10]) ? node7499 : node7496;
												assign node7496 = (inp[2]) ? 4'b0101 : 4'b1101;
												assign node7499 = (inp[13]) ? 4'b0101 : node7500;
													assign node7500 = (inp[2]) ? 4'b0101 : 4'b1101;
										assign node7504 = (inp[4]) ? node7514 : node7505;
											assign node7505 = (inp[1]) ? node7507 : 4'b0001;
												assign node7507 = (inp[2]) ? node7509 : 4'b1101;
													assign node7509 = (inp[6]) ? 4'b0101 : node7510;
														assign node7510 = (inp[11]) ? 4'b1101 : 4'b0101;
											assign node7514 = (inp[2]) ? 4'b1001 : node7515;
												assign node7515 = (inp[10]) ? 4'b0001 : 4'b0101;
									assign node7519 = (inp[10]) ? node7551 : node7520;
										assign node7520 = (inp[13]) ? node7538 : node7521;
											assign node7521 = (inp[11]) ? node7527 : node7522;
												assign node7522 = (inp[2]) ? node7524 : 4'b1001;
													assign node7524 = (inp[1]) ? 4'b1001 : 4'b0001;
												assign node7527 = (inp[2]) ? node7531 : node7528;
													assign node7528 = (inp[9]) ? 4'b0001 : 4'b0101;
													assign node7531 = (inp[6]) ? node7535 : node7532;
														assign node7532 = (inp[9]) ? 4'b1011 : 4'b1111;
														assign node7535 = (inp[4]) ? 4'b0111 : 4'b1111;
											assign node7538 = (inp[4]) ? node7546 : node7539;
												assign node7539 = (inp[9]) ? node7543 : node7540;
													assign node7540 = (inp[11]) ? 4'b0001 : 4'b0101;
													assign node7543 = (inp[1]) ? 4'b0111 : 4'b1111;
												assign node7546 = (inp[2]) ? node7548 : 4'b0111;
													assign node7548 = (inp[11]) ? 4'b0011 : 4'b0111;
										assign node7551 = (inp[6]) ? node7561 : node7552;
											assign node7552 = (inp[9]) ? node7556 : node7553;
												assign node7553 = (inp[4]) ? 4'b1111 : 4'b1001;
												assign node7556 = (inp[4]) ? 4'b1011 : node7557;
													assign node7557 = (inp[1]) ? 4'b1111 : 4'b0111;
											assign node7561 = (inp[11]) ? node7567 : node7562;
												assign node7562 = (inp[4]) ? node7564 : 4'b1111;
													assign node7564 = (inp[2]) ? 4'b1111 : 4'b1011;
												assign node7567 = (inp[2]) ? 4'b1111 : 4'b0111;
								assign node7570 = (inp[9]) ? node7596 : node7571;
									assign node7571 = (inp[4]) ? node7585 : node7572;
										assign node7572 = (inp[3]) ? node7576 : node7573;
											assign node7573 = (inp[10]) ? 4'b0001 : 4'b1001;
											assign node7576 = (inp[10]) ? node7578 : 4'b1011;
												assign node7578 = (inp[2]) ? 4'b1011 : node7579;
													assign node7579 = (inp[1]) ? 4'b0011 : node7580;
														assign node7580 = (inp[11]) ? 4'b0011 : 4'b0011;
										assign node7585 = (inp[6]) ? node7589 : node7586;
											assign node7586 = (inp[10]) ? 4'b1111 : 4'b0001;
											assign node7589 = (inp[11]) ? node7591 : 4'b1111;
												assign node7591 = (inp[1]) ? 4'b0111 : node7592;
													assign node7592 = (inp[13]) ? 4'b0111 : 4'b1111;
									assign node7596 = (inp[4]) ? node7622 : node7597;
										assign node7597 = (inp[10]) ? node7607 : node7598;
											assign node7598 = (inp[13]) ? node7604 : node7599;
												assign node7599 = (inp[1]) ? 4'b1111 : node7600;
													assign node7600 = (inp[3]) ? 4'b0011 : 4'b1111;
												assign node7604 = (inp[3]) ? 4'b0011 : 4'b0001;
											assign node7607 = (inp[3]) ? node7617 : node7608;
												assign node7608 = (inp[13]) ? node7614 : node7609;
													assign node7609 = (inp[11]) ? 4'b0111 : node7610;
														assign node7610 = (inp[2]) ? 4'b0111 : 4'b1111;
													assign node7614 = (inp[2]) ? 4'b1111 : 4'b0111;
												assign node7617 = (inp[1]) ? 4'b0111 : node7618;
													assign node7618 = (inp[11]) ? 4'b1111 : 4'b0111;
										assign node7622 = (inp[13]) ? node7630 : node7623;
											assign node7623 = (inp[1]) ? node7627 : node7624;
												assign node7624 = (inp[10]) ? 4'b0011 : 4'b0111;
												assign node7627 = (inp[3]) ? 4'b0011 : 4'b1011;
											assign node7630 = (inp[11]) ? node7632 : 4'b1011;
												assign node7632 = (inp[6]) ? 4'b0011 : 4'b1011;
					assign node7635 = (inp[1]) ? node8035 : node7636;
						assign node7636 = (inp[15]) ? node7844 : node7637;
							assign node7637 = (inp[5]) ? node7743 : node7638;
								assign node7638 = (inp[3]) ? node7696 : node7639;
									assign node7639 = (inp[12]) ? node7669 : node7640;
										assign node7640 = (inp[11]) ? node7654 : node7641;
											assign node7641 = (inp[10]) ? node7649 : node7642;
												assign node7642 = (inp[6]) ? node7646 : node7643;
													assign node7643 = (inp[4]) ? 4'b0110 : 4'b0010;
													assign node7646 = (inp[13]) ? 4'b1010 : 4'b0010;
												assign node7649 = (inp[13]) ? 4'b1110 : node7650;
													assign node7650 = (inp[9]) ? 4'b1110 : 4'b1010;
											assign node7654 = (inp[9]) ? node7664 : node7655;
												assign node7655 = (inp[4]) ? 4'b0010 : node7656;
													assign node7656 = (inp[2]) ? node7660 : node7657;
														assign node7657 = (inp[10]) ? 4'b0110 : 4'b1110;
														assign node7660 = (inp[6]) ? 4'b0010 : 4'b1010;
												assign node7664 = (inp[10]) ? 4'b1010 : node7665;
													assign node7665 = (inp[13]) ? 4'b0010 : 4'b1010;
										assign node7669 = (inp[9]) ? node7679 : node7670;
											assign node7670 = (inp[4]) ? node7672 : 4'b1010;
												assign node7672 = (inp[13]) ? 4'b1110 : node7673;
													assign node7673 = (inp[2]) ? node7675 : 4'b0010;
														assign node7675 = (inp[6]) ? 4'b1110 : 4'b0110;
											assign node7679 = (inp[13]) ? node7689 : node7680;
												assign node7680 = (inp[10]) ? node7686 : node7681;
													assign node7681 = (inp[4]) ? node7683 : 4'b1010;
														assign node7683 = (inp[11]) ? 4'b1010 : 4'b0110;
													assign node7686 = (inp[2]) ? 4'b1110 : 4'b0110;
												assign node7689 = (inp[2]) ? node7691 : 4'b1010;
													assign node7691 = (inp[11]) ? node7693 : 4'b0010;
														assign node7693 = (inp[6]) ? 4'b0010 : 4'b1010;
									assign node7696 = (inp[4]) ? node7716 : node7697;
										assign node7697 = (inp[12]) ? node7709 : node7698;
											assign node7698 = (inp[9]) ? 4'b0010 : node7699;
												assign node7699 = (inp[11]) ? 4'b1110 : node7700;
													assign node7700 = (inp[2]) ? node7704 : node7701;
														assign node7701 = (inp[10]) ? 4'b0110 : 4'b1110;
														assign node7704 = (inp[10]) ? 4'b1110 : 4'b0110;
											assign node7709 = (inp[10]) ? node7711 : 4'b0010;
												assign node7711 = (inp[9]) ? node7713 : 4'b1010;
													assign node7713 = (inp[13]) ? 4'b0100 : 4'b1100;
										assign node7716 = (inp[6]) ? node7734 : node7717;
											assign node7717 = (inp[9]) ? node7729 : node7718;
												assign node7718 = (inp[10]) ? node7724 : node7719;
													assign node7719 = (inp[13]) ? 4'b0010 : node7720;
														assign node7720 = (inp[2]) ? 4'b1010 : 4'b0010;
													assign node7724 = (inp[12]) ? node7726 : 4'b0010;
														assign node7726 = (inp[13]) ? 4'b0100 : 4'b1100;
												assign node7729 = (inp[12]) ? node7731 : 4'b1100;
													assign node7731 = (inp[2]) ? 4'b0000 : 4'b1000;
											assign node7734 = (inp[13]) ? node7738 : node7735;
												assign node7735 = (inp[11]) ? 4'b1000 : 4'b0100;
												assign node7738 = (inp[10]) ? 4'b1000 : node7739;
													assign node7739 = (inp[11]) ? 4'b0100 : 4'b1100;
								assign node7743 = (inp[3]) ? node7803 : node7744;
									assign node7744 = (inp[9]) ? node7778 : node7745;
										assign node7745 = (inp[4]) ? node7761 : node7746;
											assign node7746 = (inp[10]) ? node7752 : node7747;
												assign node7747 = (inp[12]) ? 4'b0110 : node7748;
													assign node7748 = (inp[11]) ? 4'b1110 : 4'b0110;
												assign node7752 = (inp[2]) ? node7756 : node7753;
													assign node7753 = (inp[11]) ? 4'b0110 : 4'b1110;
													assign node7756 = (inp[6]) ? node7758 : 4'b1010;
														assign node7758 = (inp[11]) ? 4'b0010 : 4'b1010;
											assign node7761 = (inp[10]) ? node7767 : node7762;
												assign node7762 = (inp[6]) ? 4'b1010 : node7763;
													assign node7763 = (inp[11]) ? 4'b0010 : 4'b1010;
												assign node7767 = (inp[2]) ? node7773 : node7768;
													assign node7768 = (inp[11]) ? 4'b1100 : node7769;
														assign node7769 = (inp[12]) ? 4'b1100 : 4'b1010;
													assign node7773 = (inp[11]) ? 4'b1100 : node7774;
														assign node7774 = (inp[6]) ? 4'b1100 : 4'b0100;
										assign node7778 = (inp[10]) ? node7792 : node7779;
											assign node7779 = (inp[4]) ? node7785 : node7780;
												assign node7780 = (inp[12]) ? 4'b0010 : node7781;
													assign node7781 = (inp[2]) ? 4'b0010 : 4'b1010;
												assign node7785 = (inp[12]) ? node7789 : node7786;
													assign node7786 = (inp[2]) ? 4'b1100 : 4'b0100;
													assign node7789 = (inp[6]) ? 4'b0000 : 4'b1000;
											assign node7792 = (inp[4]) ? node7798 : node7793;
												assign node7793 = (inp[13]) ? node7795 : 4'b0100;
													assign node7795 = (inp[12]) ? 4'b1100 : 4'b0100;
												assign node7798 = (inp[11]) ? 4'b0000 : node7799;
													assign node7799 = (inp[12]) ? 4'b1000 : 4'b1100;
									assign node7803 = (inp[2]) ? node7823 : node7804;
										assign node7804 = (inp[12]) ? node7816 : node7805;
											assign node7805 = (inp[10]) ? node7811 : node7806;
												assign node7806 = (inp[4]) ? 4'b1100 : node7807;
													assign node7807 = (inp[9]) ? 4'b1000 : 4'b1100;
												assign node7811 = (inp[6]) ? node7813 : 4'b0000;
													assign node7813 = (inp[11]) ? 4'b1100 : 4'b0000;
											assign node7816 = (inp[6]) ? node7820 : node7817;
												assign node7817 = (inp[13]) ? 4'b1100 : 4'b0100;
												assign node7820 = (inp[4]) ? 4'b1100 : 4'b1000;
										assign node7823 = (inp[13]) ? node7835 : node7824;
											assign node7824 = (inp[12]) ? 4'b0100 : node7825;
												assign node7825 = (inp[6]) ? node7831 : node7826;
													assign node7826 = (inp[9]) ? 4'b0100 : node7827;
														assign node7827 = (inp[4]) ? 4'b0000 : 4'b0100;
													assign node7831 = (inp[10]) ? 4'b1100 : 4'b1000;
											assign node7835 = (inp[10]) ? node7837 : 4'b1000;
												assign node7837 = (inp[11]) ? node7839 : 4'b0100;
													assign node7839 = (inp[12]) ? 4'b1000 : node7840;
														assign node7840 = (inp[9]) ? 4'b0100 : 4'b0000;
							assign node7844 = (inp[5]) ? node7944 : node7845;
								assign node7845 = (inp[3]) ? node7887 : node7846;
									assign node7846 = (inp[9]) ? node7858 : node7847;
										assign node7847 = (inp[10]) ? 4'b0100 : node7848;
											assign node7848 = (inp[6]) ? 4'b0000 : node7849;
												assign node7849 = (inp[12]) ? node7851 : 4'b0000;
													assign node7851 = (inp[4]) ? 4'b1100 : node7852;
														assign node7852 = (inp[13]) ? 4'b1000 : 4'b1100;
										assign node7858 = (inp[13]) ? node7872 : node7859;
											assign node7859 = (inp[2]) ? node7865 : node7860;
												assign node7860 = (inp[4]) ? node7862 : 4'b0000;
													assign node7862 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node7865 = (inp[12]) ? node7867 : 4'b0000;
													assign node7867 = (inp[6]) ? 4'b0100 : node7868;
														assign node7868 = (inp[11]) ? 4'b0100 : 4'b1000;
											assign node7872 = (inp[10]) ? node7882 : node7873;
												assign node7873 = (inp[4]) ? node7877 : node7874;
													assign node7874 = (inp[11]) ? 4'b0000 : 4'b1000;
													assign node7877 = (inp[12]) ? node7879 : 4'b0100;
														assign node7879 = (inp[6]) ? 4'b0000 : 4'b0100;
												assign node7882 = (inp[4]) ? node7884 : 4'b1100;
													assign node7884 = (inp[2]) ? 4'b1000 : 4'b0000;
									assign node7887 = (inp[9]) ? node7919 : node7888;
										assign node7888 = (inp[4]) ? node7906 : node7889;
											assign node7889 = (inp[12]) ? node7901 : node7890;
												assign node7890 = (inp[13]) ? node7896 : node7891;
													assign node7891 = (inp[11]) ? 4'b1100 : node7892;
														assign node7892 = (inp[2]) ? 4'b1100 : 4'b0100;
													assign node7896 = (inp[10]) ? node7898 : 4'b0100;
														assign node7898 = (inp[11]) ? 4'b0000 : 4'b0100;
												assign node7901 = (inp[13]) ? node7903 : 4'b1000;
													assign node7903 = (inp[2]) ? 4'b0000 : 4'b1000;
											assign node7906 = (inp[11]) ? node7914 : node7907;
												assign node7907 = (inp[13]) ? node7911 : node7908;
													assign node7908 = (inp[6]) ? 4'b0000 : 4'b1000;
													assign node7911 = (inp[12]) ? 4'b0110 : 4'b0000;
												assign node7914 = (inp[2]) ? node7916 : 4'b1110;
													assign node7916 = (inp[10]) ? 4'b0110 : 4'b0000;
										assign node7919 = (inp[4]) ? node7933 : node7920;
											assign node7920 = (inp[6]) ? node7924 : node7921;
												assign node7921 = (inp[2]) ? 4'b1000 : 4'b0000;
												assign node7924 = (inp[10]) ? node7926 : 4'b0000;
													assign node7926 = (inp[11]) ? node7930 : node7927;
														assign node7927 = (inp[13]) ? 4'b1110 : 4'b0000;
														assign node7930 = (inp[13]) ? 4'b0110 : 4'b1110;
											assign node7933 = (inp[11]) ? node7939 : node7934;
												assign node7934 = (inp[10]) ? 4'b0010 : node7935;
													assign node7935 = (inp[12]) ? 4'b0110 : 4'b1110;
												assign node7939 = (inp[6]) ? node7941 : 4'b1110;
													assign node7941 = (inp[13]) ? 4'b0010 : 4'b1010;
								assign node7944 = (inp[3]) ? node7998 : node7945;
									assign node7945 = (inp[4]) ? node7969 : node7946;
										assign node7946 = (inp[9]) ? node7958 : node7947;
											assign node7947 = (inp[10]) ? 4'b1000 : node7948;
												assign node7948 = (inp[12]) ? node7952 : node7949;
													assign node7949 = (inp[6]) ? 4'b0100 : 4'b1100;
													assign node7952 = (inp[11]) ? 4'b1000 : node7953;
														assign node7953 = (inp[6]) ? 4'b1000 : 4'b0100;
											assign node7958 = (inp[12]) ? node7962 : node7959;
												assign node7959 = (inp[2]) ? 4'b0000 : 4'b1000;
												assign node7962 = (inp[6]) ? 4'b0110 : node7963;
													assign node7963 = (inp[11]) ? 4'b1110 : node7964;
														assign node7964 = (inp[2]) ? 4'b1110 : 4'b1000;
										assign node7969 = (inp[9]) ? node7983 : node7970;
											assign node7970 = (inp[13]) ? node7980 : node7971;
												assign node7971 = (inp[12]) ? node7975 : node7972;
													assign node7972 = (inp[2]) ? 4'b0000 : 4'b1000;
													assign node7975 = (inp[11]) ? 4'b1110 : node7976;
														assign node7976 = (inp[6]) ? 4'b0000 : 4'b1110;
												assign node7980 = (inp[12]) ? 4'b1110 : 4'b0110;
											assign node7983 = (inp[12]) ? node7991 : node7984;
												assign node7984 = (inp[11]) ? node7988 : node7985;
													assign node7985 = (inp[13]) ? 4'b0110 : 4'b1110;
													assign node7988 = (inp[10]) ? 4'b1010 : 4'b1110;
												assign node7991 = (inp[13]) ? node7993 : 4'b0010;
													assign node7993 = (inp[10]) ? 4'b1010 : node7994;
														assign node7994 = (inp[6]) ? 4'b1010 : 4'b0010;
									assign node7998 = (inp[11]) ? node8026 : node7999;
										assign node7999 = (inp[4]) ? node8015 : node8000;
											assign node8000 = (inp[10]) ? node8004 : node8001;
												assign node8001 = (inp[6]) ? 4'b1110 : 4'b0010;
												assign node8004 = (inp[12]) ? node8008 : node8005;
													assign node8005 = (inp[2]) ? 4'b0010 : 4'b0110;
													assign node8008 = (inp[13]) ? node8012 : node8009;
														assign node8009 = (inp[6]) ? 4'b0110 : 4'b1110;
														assign node8012 = (inp[6]) ? 4'b1110 : 4'b0110;
											assign node8015 = (inp[2]) ? node8017 : 4'b1010;
												assign node8017 = (inp[10]) ? node8023 : node8018;
													assign node8018 = (inp[6]) ? 4'b1110 : node8019;
														assign node8019 = (inp[13]) ? 4'b0010 : 4'b1110;
													assign node8023 = (inp[9]) ? 4'b1010 : 4'b0010;
										assign node8026 = (inp[12]) ? node8030 : node8027;
											assign node8027 = (inp[13]) ? 4'b0010 : 4'b1010;
											assign node8030 = (inp[9]) ? 4'b0010 : node8031;
												assign node8031 = (inp[10]) ? 4'b1110 : 4'b0010;
						assign node8035 = (inp[10]) ? node8187 : node8036;
							assign node8036 = (inp[11]) ? node8116 : node8037;
								assign node8037 = (inp[6]) ? node8077 : node8038;
									assign node8038 = (inp[12]) ? node8060 : node8039;
										assign node8039 = (inp[3]) ? node8051 : node8040;
											assign node8040 = (inp[15]) ? node8046 : node8041;
												assign node8041 = (inp[2]) ? 4'b0010 : node8042;
													assign node8042 = (inp[13]) ? 4'b0010 : 4'b0110;
												assign node8046 = (inp[5]) ? node8048 : 4'b0000;
													assign node8048 = (inp[4]) ? 4'b0110 : 4'b0100;
											assign node8051 = (inp[15]) ? 4'b0110 : node8052;
												assign node8052 = (inp[5]) ? node8054 : 4'b0110;
													assign node8054 = (inp[4]) ? 4'b0100 : node8055;
														assign node8055 = (inp[13]) ? 4'b0000 : 4'b0100;
										assign node8060 = (inp[13]) ? node8072 : node8061;
											assign node8061 = (inp[9]) ? node8067 : node8062;
												assign node8062 = (inp[15]) ? 4'b0000 : node8063;
													assign node8063 = (inp[4]) ? 4'b0010 : 4'b0110;
												assign node8067 = (inp[4]) ? node8069 : 4'b0010;
													assign node8069 = (inp[2]) ? 4'b0110 : 4'b0100;
											assign node8072 = (inp[4]) ? 4'b0000 : node8073;
												assign node8073 = (inp[5]) ? 4'b0010 : 4'b0000;
									assign node8077 = (inp[5]) ? node8097 : node8078;
										assign node8078 = (inp[15]) ? node8086 : node8079;
											assign node8079 = (inp[13]) ? 4'b1010 : node8080;
												assign node8080 = (inp[3]) ? 4'b1100 : node8081;
													assign node8081 = (inp[9]) ? 4'b1110 : 4'b1010;
											assign node8086 = (inp[3]) ? node8094 : node8087;
												assign node8087 = (inp[2]) ? node8089 : 4'b1100;
													assign node8089 = (inp[4]) ? node8091 : 4'b1000;
														assign node8091 = (inp[13]) ? 4'b1000 : 4'b1100;
												assign node8094 = (inp[9]) ? 4'b1010 : 4'b1000;
										assign node8097 = (inp[15]) ? node8105 : node8098;
											assign node8098 = (inp[4]) ? 4'b1100 : node8099;
												assign node8099 = (inp[9]) ? node8101 : 4'b1010;
													assign node8101 = (inp[12]) ? 4'b1100 : 4'b1010;
											assign node8105 = (inp[9]) ? node8111 : node8106;
												assign node8106 = (inp[12]) ? node8108 : 4'b1010;
													assign node8108 = (inp[4]) ? 4'b1110 : 4'b1010;
												assign node8111 = (inp[13]) ? node8113 : 4'b1110;
													assign node8113 = (inp[2]) ? 4'b1110 : 4'b1010;
								assign node8116 = (inp[6]) ? node8158 : node8117;
									assign node8117 = (inp[4]) ? node8143 : node8118;
										assign node8118 = (inp[2]) ? node8130 : node8119;
											assign node8119 = (inp[5]) ? node8125 : node8120;
												assign node8120 = (inp[15]) ? node8122 : 4'b1010;
													assign node8122 = (inp[12]) ? 4'b1000 : 4'b1100;
												assign node8125 = (inp[15]) ? 4'b1110 : node8126;
													assign node8126 = (inp[12]) ? 4'b1100 : 4'b1000;
											assign node8130 = (inp[15]) ? node8136 : node8131;
												assign node8131 = (inp[3]) ? 4'b1100 : node8132;
													assign node8132 = (inp[9]) ? 4'b1100 : 4'b1110;
												assign node8136 = (inp[3]) ? node8140 : node8137;
													assign node8137 = (inp[13]) ? 4'b1100 : 4'b1000;
													assign node8140 = (inp[12]) ? 4'b1110 : 4'b1010;
										assign node8143 = (inp[2]) ? node8149 : node8144;
											assign node8144 = (inp[12]) ? 4'b1110 : node8145;
												assign node8145 = (inp[5]) ? 4'b1110 : 4'b1010;
											assign node8149 = (inp[12]) ? node8155 : node8150;
												assign node8150 = (inp[9]) ? node8152 : 4'b1010;
													assign node8152 = (inp[13]) ? 4'b1100 : 4'b1110;
												assign node8155 = (inp[9]) ? 4'b1000 : 4'b1100;
									assign node8158 = (inp[2]) ? node8170 : node8159;
										assign node8159 = (inp[15]) ? node8165 : node8160;
											assign node8160 = (inp[3]) ? node8162 : 4'b0110;
												assign node8162 = (inp[12]) ? 4'b0000 : 4'b0100;
											assign node8165 = (inp[5]) ? 4'b0110 : node8166;
												assign node8166 = (inp[12]) ? 4'b0010 : 4'b0110;
										assign node8170 = (inp[5]) ? node8180 : node8171;
											assign node8171 = (inp[15]) ? node8173 : 4'b0110;
												assign node8173 = (inp[13]) ? 4'b0110 : node8174;
													assign node8174 = (inp[9]) ? node8176 : 4'b0000;
														assign node8176 = (inp[3]) ? 4'b0110 : 4'b0100;
											assign node8180 = (inp[15]) ? node8182 : 4'b0000;
												assign node8182 = (inp[13]) ? node8184 : 4'b0010;
													assign node8184 = (inp[9]) ? 4'b0110 : 4'b0100;
							assign node8187 = (inp[9]) ? node8259 : node8188;
								assign node8188 = (inp[4]) ? node8222 : node8189;
									assign node8189 = (inp[15]) ? node8203 : node8190;
										assign node8190 = (inp[6]) ? node8200 : node8191;
											assign node8191 = (inp[11]) ? node8197 : node8192;
												assign node8192 = (inp[12]) ? 4'b0010 : node8193;
													assign node8193 = (inp[2]) ? 4'b0100 : 4'b0110;
												assign node8197 = (inp[3]) ? 4'b1000 : 4'b1010;
											assign node8200 = (inp[11]) ? 4'b0010 : 4'b1010;
										assign node8203 = (inp[3]) ? node8213 : node8204;
											assign node8204 = (inp[12]) ? 4'b1000 : node8205;
												assign node8205 = (inp[2]) ? node8207 : 4'b0000;
													assign node8207 = (inp[11]) ? node8209 : 4'b1000;
														assign node8209 = (inp[13]) ? 4'b0000 : 4'b1000;
											assign node8213 = (inp[5]) ? node8217 : node8214;
												assign node8214 = (inp[2]) ? 4'b1000 : 4'b0100;
												assign node8217 = (inp[11]) ? node8219 : 4'b1010;
													assign node8219 = (inp[6]) ? 4'b0010 : 4'b1010;
									assign node8222 = (inp[15]) ? node8242 : node8223;
										assign node8223 = (inp[5]) ? node8231 : node8224;
											assign node8224 = (inp[3]) ? node8226 : 4'b1110;
												assign node8226 = (inp[11]) ? node8228 : 4'b0010;
													assign node8228 = (inp[2]) ? 4'b0100 : 4'b1100;
											assign node8231 = (inp[13]) ? node8237 : node8232;
												assign node8232 = (inp[2]) ? node8234 : 4'b1100;
													assign node8234 = (inp[12]) ? 4'b1100 : 4'b0010;
												assign node8237 = (inp[6]) ? 4'b0100 : node8238;
													assign node8238 = (inp[11]) ? 4'b1100 : 4'b0100;
										assign node8242 = (inp[3]) ? node8254 : node8243;
											assign node8243 = (inp[5]) ? node8247 : node8244;
												assign node8244 = (inp[11]) ? 4'b0100 : 4'b1100;
												assign node8247 = (inp[13]) ? 4'b0110 : node8248;
													assign node8248 = (inp[11]) ? 4'b1110 : node8249;
														assign node8249 = (inp[6]) ? 4'b1110 : 4'b0110;
											assign node8254 = (inp[2]) ? node8256 : 4'b1110;
												assign node8256 = (inp[6]) ? 4'b0110 : 4'b1110;
								assign node8259 = (inp[4]) ? node8289 : node8260;
									assign node8260 = (inp[3]) ? node8282 : node8261;
										assign node8261 = (inp[2]) ? node8269 : node8262;
											assign node8262 = (inp[11]) ? node8266 : node8263;
												assign node8263 = (inp[15]) ? 4'b1100 : 4'b1110;
												assign node8266 = (inp[6]) ? 4'b0100 : 4'b1100;
											assign node8269 = (inp[12]) ? node8271 : 4'b1110;
												assign node8271 = (inp[13]) ? node8277 : node8272;
													assign node8272 = (inp[5]) ? node8274 : 4'b0100;
														assign node8274 = (inp[11]) ? 4'b1110 : 4'b0100;
													assign node8277 = (inp[11]) ? 4'b0100 : node8278;
														assign node8278 = (inp[6]) ? 4'b1110 : 4'b0110;
										assign node8282 = (inp[15]) ? 4'b1110 : node8283;
											assign node8283 = (inp[11]) ? 4'b1100 : node8284;
												assign node8284 = (inp[6]) ? 4'b1100 : 4'b0100;
									assign node8289 = (inp[15]) ? node8299 : node8290;
										assign node8290 = (inp[5]) ? node8294 : node8291;
											assign node8291 = (inp[3]) ? 4'b1000 : 4'b1010;
											assign node8294 = (inp[11]) ? node8296 : 4'b1000;
												assign node8296 = (inp[6]) ? 4'b0000 : 4'b1000;
										assign node8299 = (inp[3]) ? 4'b1010 : node8300;
											assign node8300 = (inp[5]) ? node8306 : node8301;
												assign node8301 = (inp[6]) ? 4'b1000 : node8302;
													assign node8302 = (inp[11]) ? 4'b1000 : 4'b0000;
												assign node8306 = (inp[11]) ? 4'b0010 : 4'b1010;
			assign node8310 = (inp[11]) ? node9572 : node8311;
				assign node8311 = (inp[6]) ? node8923 : node8312;
					assign node8312 = (inp[13]) ? node8646 : node8313;
						assign node8313 = (inp[1]) ? node8467 : node8314;
							assign node8314 = (inp[12]) ? node8386 : node8315;
								assign node8315 = (inp[7]) ? node8347 : node8316;
									assign node8316 = (inp[8]) ? node8338 : node8317;
										assign node8317 = (inp[5]) ? node8329 : node8318;
											assign node8318 = (inp[15]) ? node8326 : node8319;
												assign node8319 = (inp[3]) ? 4'b1100 : node8320;
													assign node8320 = (inp[4]) ? node8322 : 4'b1000;
														assign node8322 = (inp[9]) ? 4'b1100 : 4'b1000;
												assign node8326 = (inp[2]) ? 4'b1010 : 4'b1110;
											assign node8329 = (inp[15]) ? node8333 : node8330;
												assign node8330 = (inp[4]) ? 4'b1110 : 4'b1100;
												assign node8333 = (inp[2]) ? 4'b1100 : node8334;
													assign node8334 = (inp[9]) ? 4'b1010 : 4'b1110;
										assign node8338 = (inp[9]) ? node8344 : node8339;
											assign node8339 = (inp[4]) ? 4'b1011 : node8340;
												assign node8340 = (inp[10]) ? 4'b1111 : 4'b1101;
											assign node8344 = (inp[4]) ? 4'b1101 : 4'b1001;
									assign node8347 = (inp[8]) ? node8365 : node8348;
										assign node8348 = (inp[15]) ? node8356 : node8349;
											assign node8349 = (inp[3]) ? 4'b1011 : node8350;
												assign node8350 = (inp[10]) ? 4'b1001 : node8351;
													assign node8351 = (inp[9]) ? 4'b1111 : 4'b1001;
											assign node8356 = (inp[3]) ? node8362 : node8357;
												assign node8357 = (inp[10]) ? node8359 : 4'b1111;
													assign node8359 = (inp[9]) ? 4'b1111 : 4'b1011;
												assign node8362 = (inp[2]) ? 4'b1001 : 4'b1101;
										assign node8365 = (inp[5]) ? node8375 : node8366;
											assign node8366 = (inp[15]) ? node8368 : 4'b1000;
												assign node8368 = (inp[2]) ? 4'b1110 : node8369;
													assign node8369 = (inp[9]) ? 4'b1010 : node8370;
														assign node8370 = (inp[4]) ? 4'b1010 : 4'b1110;
											assign node8375 = (inp[3]) ? node8383 : node8376;
												assign node8376 = (inp[9]) ? node8380 : node8377;
													assign node8377 = (inp[2]) ? 4'b1110 : 4'b1010;
													assign node8380 = (inp[4]) ? 4'b1100 : 4'b1010;
												assign node8383 = (inp[15]) ? 4'b1100 : 4'b1110;
								assign node8386 = (inp[9]) ? node8428 : node8387;
									assign node8387 = (inp[8]) ? node8407 : node8388;
										assign node8388 = (inp[7]) ? node8402 : node8389;
											assign node8389 = (inp[4]) ? node8397 : node8390;
												assign node8390 = (inp[10]) ? node8394 : node8391;
													assign node8391 = (inp[5]) ? 4'b1110 : 4'b1100;
													assign node8394 = (inp[15]) ? 4'b1000 : 4'b1010;
												assign node8397 = (inp[5]) ? node8399 : 4'b1010;
													assign node8399 = (inp[10]) ? 4'b1100 : 4'b1000;
											assign node8402 = (inp[3]) ? node8404 : 4'b1011;
												assign node8404 = (inp[4]) ? 4'b1101 : 4'b1001;
										assign node8407 = (inp[7]) ? node8417 : node8408;
											assign node8408 = (inp[5]) ? node8414 : node8409;
												assign node8409 = (inp[3]) ? node8411 : 4'b1101;
													assign node8411 = (inp[4]) ? 4'b1001 : 4'b1101;
												assign node8414 = (inp[15]) ? 4'b1101 : 4'b1111;
											assign node8417 = (inp[15]) ? node8423 : node8418;
												assign node8418 = (inp[2]) ? 4'b1000 : node8419;
													assign node8419 = (inp[4]) ? 4'b1100 : 4'b1000;
												assign node8423 = (inp[4]) ? node8425 : 4'b1110;
													assign node8425 = (inp[3]) ? 4'b1000 : 4'b1100;
									assign node8428 = (inp[15]) ? node8452 : node8429;
										assign node8429 = (inp[5]) ? node8441 : node8430;
											assign node8430 = (inp[3]) ? node8438 : node8431;
												assign node8431 = (inp[7]) ? node8433 : 4'b1100;
													assign node8433 = (inp[4]) ? node8435 : 4'b1100;
														assign node8435 = (inp[8]) ? 4'b1000 : 4'b1001;
												assign node8438 = (inp[10]) ? 4'b1011 : 4'b1001;
											assign node8441 = (inp[2]) ? node8445 : node8442;
												assign node8442 = (inp[8]) ? 4'b1011 : 4'b1010;
												assign node8445 = (inp[10]) ? node8449 : node8446;
													assign node8446 = (inp[3]) ? 4'b1011 : 4'b1001;
													assign node8449 = (inp[8]) ? 4'b1011 : 4'b1111;
										assign node8452 = (inp[4]) ? node8464 : node8453;
											assign node8453 = (inp[10]) ? node8457 : node8454;
												assign node8454 = (inp[7]) ? 4'b1011 : 4'b1000;
												assign node8457 = (inp[2]) ? 4'b1100 : node8458;
													assign node8458 = (inp[8]) ? 4'b1111 : node8459;
														assign node8459 = (inp[7]) ? 4'b1101 : 4'b1100;
											assign node8464 = (inp[10]) ? 4'b1001 : 4'b1101;
							assign node8467 = (inp[7]) ? node8563 : node8468;
								assign node8468 = (inp[8]) ? node8530 : node8469;
									assign node8469 = (inp[2]) ? node8501 : node8470;
										assign node8470 = (inp[12]) ? node8480 : node8471;
											assign node8471 = (inp[10]) ? node8477 : node8472;
												assign node8472 = (inp[5]) ? 4'b1110 : node8473;
													assign node8473 = (inp[15]) ? 4'b1010 : 4'b1000;
												assign node8477 = (inp[9]) ? 4'b1100 : 4'b1000;
											assign node8480 = (inp[9]) ? node8492 : node8481;
												assign node8481 = (inp[15]) ? node8487 : node8482;
													assign node8482 = (inp[5]) ? node8484 : 4'b1100;
														assign node8484 = (inp[4]) ? 4'b1000 : 4'b1100;
													assign node8487 = (inp[4]) ? 4'b1100 : node8488;
														assign node8488 = (inp[3]) ? 4'b1100 : 4'b1110;
												assign node8492 = (inp[5]) ? node8496 : node8493;
													assign node8493 = (inp[4]) ? 4'b1110 : 4'b1000;
													assign node8496 = (inp[15]) ? node8498 : 4'b1110;
														assign node8498 = (inp[10]) ? 4'b1000 : 4'b1100;
										assign node8501 = (inp[15]) ? node8525 : node8502;
											assign node8502 = (inp[10]) ? node8514 : node8503;
												assign node8503 = (inp[12]) ? node8509 : node8504;
													assign node8504 = (inp[9]) ? 4'b1000 : node8505;
														assign node8505 = (inp[4]) ? 4'b1000 : 4'b1100;
													assign node8509 = (inp[3]) ? node8511 : 4'b1100;
														assign node8511 = (inp[9]) ? 4'b1110 : 4'b1000;
												assign node8514 = (inp[4]) ? node8520 : node8515;
													assign node8515 = (inp[5]) ? node8517 : 4'b1000;
														assign node8517 = (inp[3]) ? 4'b1010 : 4'b1000;
													assign node8520 = (inp[3]) ? node8522 : 4'b1010;
														assign node8522 = (inp[9]) ? 4'b1110 : 4'b1010;
											assign node8525 = (inp[3]) ? 4'b1000 : node8526;
												assign node8526 = (inp[12]) ? 4'b1010 : 4'b1110;
									assign node8530 = (inp[15]) ? node8552 : node8531;
										assign node8531 = (inp[9]) ? node8543 : node8532;
											assign node8532 = (inp[4]) ? node8538 : node8533;
												assign node8533 = (inp[10]) ? node8535 : 4'b0101;
													assign node8535 = (inp[12]) ? 4'b0001 : 4'b0101;
												assign node8538 = (inp[12]) ? node8540 : 4'b0001;
													assign node8540 = (inp[2]) ? 4'b0001 : 4'b0111;
											assign node8543 = (inp[3]) ? node8545 : 4'b0001;
												assign node8545 = (inp[5]) ? node8547 : 4'b0001;
													assign node8547 = (inp[10]) ? node8549 : 4'b0011;
														assign node8549 = (inp[2]) ? 4'b0011 : 4'b0111;
										assign node8552 = (inp[4]) ? node8556 : node8553;
											assign node8553 = (inp[9]) ? 4'b0011 : 4'b0111;
											assign node8556 = (inp[5]) ? 4'b0001 : node8557;
												assign node8557 = (inp[10]) ? node8559 : 4'b0011;
													assign node8559 = (inp[2]) ? 4'b0111 : 4'b0101;
								assign node8563 = (inp[8]) ? node8599 : node8564;
									assign node8564 = (inp[15]) ? node8580 : node8565;
										assign node8565 = (inp[3]) ? node8573 : node8566;
											assign node8566 = (inp[5]) ? 4'b0001 : node8567;
												assign node8567 = (inp[2]) ? 4'b0101 : node8568;
													assign node8568 = (inp[9]) ? 4'b0001 : 4'b0101;
											assign node8573 = (inp[12]) ? 4'b0111 : node8574;
												assign node8574 = (inp[9]) ? 4'b0011 : node8575;
													assign node8575 = (inp[4]) ? 4'b0001 : 4'b0101;
										assign node8580 = (inp[5]) ? node8590 : node8581;
											assign node8581 = (inp[10]) ? node8587 : node8582;
												assign node8582 = (inp[9]) ? node8584 : 4'b0111;
													assign node8584 = (inp[4]) ? 4'b0111 : 4'b0011;
												assign node8587 = (inp[12]) ? 4'b0001 : 4'b0011;
											assign node8590 = (inp[3]) ? node8594 : node8591;
												assign node8591 = (inp[9]) ? 4'b0101 : 4'b0111;
												assign node8594 = (inp[2]) ? 4'b0001 : node8595;
													assign node8595 = (inp[4]) ? 4'b0101 : 4'b0001;
									assign node8599 = (inp[12]) ? node8625 : node8600;
										assign node8600 = (inp[15]) ? node8606 : node8601;
											assign node8601 = (inp[3]) ? node8603 : 4'b0000;
												assign node8603 = (inp[9]) ? 4'b0010 : 4'b0110;
											assign node8606 = (inp[2]) ? node8614 : node8607;
												assign node8607 = (inp[5]) ? 4'b0100 : node8608;
													assign node8608 = (inp[10]) ? 4'b0110 : node8609;
														assign node8609 = (inp[9]) ? 4'b0010 : 4'b0110;
												assign node8614 = (inp[10]) ? node8620 : node8615;
													assign node8615 = (inp[3]) ? 4'b0110 : node8616;
														assign node8616 = (inp[4]) ? 4'b0110 : 4'b0010;
													assign node8620 = (inp[4]) ? 4'b0010 : node8621;
														assign node8621 = (inp[5]) ? 4'b0110 : 4'b0010;
										assign node8625 = (inp[3]) ? node8635 : node8626;
											assign node8626 = (inp[10]) ? node8628 : 4'b0100;
												assign node8628 = (inp[5]) ? node8630 : 4'b0000;
													assign node8630 = (inp[15]) ? node8632 : 4'b0110;
														assign node8632 = (inp[2]) ? 4'b0100 : 4'b0000;
											assign node8635 = (inp[10]) ? node8637 : 4'b0000;
												assign node8637 = (inp[2]) ? node8643 : node8638;
													assign node8638 = (inp[4]) ? node8640 : 4'b0000;
														assign node8640 = (inp[9]) ? 4'b0000 : 4'b0100;
													assign node8643 = (inp[4]) ? 4'b0000 : 4'b0100;
						assign node8646 = (inp[7]) ? node8796 : node8647;
							assign node8647 = (inp[8]) ? node8739 : node8648;
								assign node8648 = (inp[1]) ? node8702 : node8649;
									assign node8649 = (inp[10]) ? node8675 : node8650;
										assign node8650 = (inp[5]) ? node8666 : node8651;
											assign node8651 = (inp[15]) ? node8661 : node8652;
												assign node8652 = (inp[2]) ? 4'b1000 : node8653;
													assign node8653 = (inp[9]) ? node8657 : node8654;
														assign node8654 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node8657 = (inp[3]) ? 4'b1110 : 4'b1100;
												assign node8661 = (inp[12]) ? 4'b1010 : node8662;
													assign node8662 = (inp[9]) ? 4'b1100 : 4'b1110;
											assign node8666 = (inp[2]) ? node8672 : node8667;
												assign node8667 = (inp[15]) ? 4'b1100 : node8668;
													assign node8668 = (inp[4]) ? 4'b1000 : 4'b1100;
												assign node8672 = (inp[15]) ? 4'b1100 : 4'b1110;
										assign node8675 = (inp[5]) ? node8691 : node8676;
											assign node8676 = (inp[15]) ? node8682 : node8677;
												assign node8677 = (inp[12]) ? 4'b1110 : node8678;
													assign node8678 = (inp[3]) ? 4'b1000 : 4'b1100;
												assign node8682 = (inp[12]) ? node8688 : node8683;
													assign node8683 = (inp[2]) ? 4'b1010 : node8684;
														assign node8684 = (inp[9]) ? 4'b1010 : 4'b1110;
													assign node8688 = (inp[3]) ? 4'b1000 : 4'b1010;
											assign node8691 = (inp[9]) ? node8697 : node8692;
												assign node8692 = (inp[15]) ? node8694 : 4'b1000;
													assign node8694 = (inp[4]) ? 4'b1000 : 4'b1100;
												assign node8697 = (inp[3]) ? 4'b1110 : node8698;
													assign node8698 = (inp[15]) ? 4'b1000 : 4'b1010;
									assign node8702 = (inp[5]) ? node8718 : node8703;
										assign node8703 = (inp[15]) ? node8715 : node8704;
											assign node8704 = (inp[9]) ? node8710 : node8705;
												assign node8705 = (inp[4]) ? 4'b0000 : node8706;
													assign node8706 = (inp[2]) ? 4'b0000 : 4'b0100;
												assign node8710 = (inp[4]) ? node8712 : 4'b0000;
													assign node8712 = (inp[3]) ? 4'b0110 : 4'b0100;
											assign node8715 = (inp[2]) ? 4'b0010 : 4'b0000;
										assign node8718 = (inp[4]) ? node8732 : node8719;
											assign node8719 = (inp[2]) ? node8729 : node8720;
												assign node8720 = (inp[9]) ? node8726 : node8721;
													assign node8721 = (inp[10]) ? 4'b0010 : node8722;
														assign node8722 = (inp[12]) ? 4'b0100 : 4'b0110;
													assign node8726 = (inp[10]) ? 4'b0110 : 4'b0010;
												assign node8729 = (inp[15]) ? 4'b0010 : 4'b0000;
											assign node8732 = (inp[9]) ? node8736 : node8733;
												assign node8733 = (inp[15]) ? 4'b0010 : 4'b0110;
												assign node8736 = (inp[15]) ? 4'b0100 : 4'b0110;
								assign node8739 = (inp[4]) ? node8775 : node8740;
									assign node8740 = (inp[15]) ? node8760 : node8741;
										assign node8741 = (inp[5]) ? node8747 : node8742;
											assign node8742 = (inp[2]) ? node8744 : 4'b0001;
												assign node8744 = (inp[9]) ? 4'b0001 : 4'b0101;
											assign node8747 = (inp[3]) ? node8753 : node8748;
												assign node8748 = (inp[2]) ? 4'b0001 : node8749;
													assign node8749 = (inp[1]) ? 4'b0101 : 4'b0111;
												assign node8753 = (inp[1]) ? node8755 : 4'b0111;
													assign node8755 = (inp[12]) ? 4'b0011 : node8756;
														assign node8756 = (inp[9]) ? 4'b0011 : 4'b0111;
										assign node8760 = (inp[3]) ? node8768 : node8761;
											assign node8761 = (inp[5]) ? node8763 : 4'b0111;
												assign node8763 = (inp[12]) ? 4'b0101 : node8764;
													assign node8764 = (inp[2]) ? 4'b0111 : 4'b0011;
											assign node8768 = (inp[10]) ? node8770 : 4'b0011;
												assign node8770 = (inp[12]) ? 4'b0101 : node8771;
													assign node8771 = (inp[5]) ? 4'b0001 : 4'b0011;
									assign node8775 = (inp[9]) ? node8785 : node8776;
										assign node8776 = (inp[10]) ? node8782 : node8777;
											assign node8777 = (inp[15]) ? node8779 : 4'b0001;
												assign node8779 = (inp[5]) ? 4'b0001 : 4'b0011;
											assign node8782 = (inp[12]) ? 4'b0111 : 4'b0011;
										assign node8785 = (inp[10]) ? node8791 : node8786;
											assign node8786 = (inp[15]) ? 4'b0101 : node8787;
												assign node8787 = (inp[1]) ? 4'b0111 : 4'b0101;
											assign node8791 = (inp[12]) ? node8793 : 4'b0111;
												assign node8793 = (inp[2]) ? 4'b0011 : 4'b0001;
							assign node8796 = (inp[8]) ? node8862 : node8797;
								assign node8797 = (inp[9]) ? node8833 : node8798;
									assign node8798 = (inp[4]) ? node8820 : node8799;
										assign node8799 = (inp[12]) ? node8811 : node8800;
											assign node8800 = (inp[15]) ? node8806 : node8801;
												assign node8801 = (inp[3]) ? node8803 : 4'b0101;
													assign node8803 = (inp[10]) ? 4'b0111 : 4'b0101;
												assign node8806 = (inp[3]) ? node8808 : 4'b0111;
													assign node8808 = (inp[1]) ? 4'b0101 : 4'b0111;
											assign node8811 = (inp[10]) ? node8813 : 4'b0111;
												assign node8813 = (inp[2]) ? 4'b0001 : node8814;
													assign node8814 = (inp[15]) ? 4'b0011 : node8815;
														assign node8815 = (inp[5]) ? 4'b0011 : 4'b0001;
										assign node8820 = (inp[12]) ? 4'b0101 : node8821;
											assign node8821 = (inp[5]) ? node8825 : node8822;
												assign node8822 = (inp[15]) ? 4'b0011 : 4'b0001;
												assign node8825 = (inp[10]) ? node8827 : 4'b0001;
													assign node8827 = (inp[2]) ? 4'b0001 : node8828;
														assign node8828 = (inp[3]) ? 4'b0011 : 4'b0001;
									assign node8833 = (inp[4]) ? node8849 : node8834;
										assign node8834 = (inp[12]) ? node8838 : node8835;
											assign node8835 = (inp[15]) ? 4'b0011 : 4'b0001;
											assign node8838 = (inp[10]) ? node8840 : 4'b0011;
												assign node8840 = (inp[3]) ? node8846 : node8841;
													assign node8841 = (inp[15]) ? 4'b0111 : node8842;
														assign node8842 = (inp[5]) ? 4'b0111 : 4'b0101;
													assign node8846 = (inp[15]) ? 4'b0101 : 4'b0111;
										assign node8849 = (inp[15]) ? node8857 : node8850;
											assign node8850 = (inp[10]) ? 4'b0011 : node8851;
												assign node8851 = (inp[1]) ? 4'b0111 : node8852;
													assign node8852 = (inp[12]) ? 4'b0111 : 4'b0101;
											assign node8857 = (inp[5]) ? 4'b0101 : node8858;
												assign node8858 = (inp[3]) ? 4'b0101 : 4'b0111;
								assign node8862 = (inp[4]) ? node8894 : node8863;
									assign node8863 = (inp[9]) ? node8875 : node8864;
										assign node8864 = (inp[5]) ? 4'b0110 : node8865;
											assign node8865 = (inp[15]) ? node8871 : node8866;
												assign node8866 = (inp[12]) ? node8868 : 4'b0100;
													assign node8868 = (inp[10]) ? 4'b0000 : 4'b0100;
												assign node8871 = (inp[12]) ? 4'b0010 : 4'b0110;
										assign node8875 = (inp[12]) ? node8889 : node8876;
											assign node8876 = (inp[15]) ? node8884 : node8877;
												assign node8877 = (inp[2]) ? node8879 : 4'b0000;
													assign node8879 = (inp[5]) ? node8881 : 4'b0000;
														assign node8881 = (inp[3]) ? 4'b0010 : 4'b0000;
												assign node8884 = (inp[10]) ? node8886 : 4'b0010;
													assign node8886 = (inp[1]) ? 4'b0000 : 4'b0010;
											assign node8889 = (inp[1]) ? 4'b0010 : node8890;
												assign node8890 = (inp[15]) ? 4'b0100 : 4'b0110;
									assign node8894 = (inp[9]) ? node8902 : node8895;
										assign node8895 = (inp[10]) ? node8897 : 4'b0000;
											assign node8897 = (inp[12]) ? 4'b0110 : node8898;
												assign node8898 = (inp[5]) ? 4'b0010 : 4'b0000;
										assign node8902 = (inp[15]) ? node8912 : node8903;
											assign node8903 = (inp[12]) ? node8909 : node8904;
												assign node8904 = (inp[3]) ? 4'b0110 : node8905;
													assign node8905 = (inp[1]) ? 4'b0100 : 4'b0110;
												assign node8909 = (inp[1]) ? 4'b0010 : 4'b0110;
											assign node8912 = (inp[1]) ? node8918 : node8913;
												assign node8913 = (inp[3]) ? 4'b0100 : node8914;
													assign node8914 = (inp[12]) ? 4'b0010 : 4'b0110;
												assign node8918 = (inp[12]) ? node8920 : 4'b0100;
													assign node8920 = (inp[10]) ? 4'b0000 : 4'b0100;
					assign node8923 = (inp[13]) ? node9277 : node8924;
						assign node8924 = (inp[1]) ? node9098 : node8925;
							assign node8925 = (inp[12]) ? node9001 : node8926;
								assign node8926 = (inp[15]) ? node8960 : node8927;
									assign node8927 = (inp[5]) ? node8943 : node8928;
										assign node8928 = (inp[9]) ? node8932 : node8929;
											assign node8929 = (inp[4]) ? 4'b0000 : 4'b0100;
											assign node8932 = (inp[4]) ? node8936 : node8933;
												assign node8933 = (inp[10]) ? 4'b0000 : 4'b0001;
												assign node8936 = (inp[3]) ? node8940 : node8937;
													assign node8937 = (inp[8]) ? 4'b0101 : 4'b0100;
													assign node8940 = (inp[2]) ? 4'b0110 : 4'b0111;
										assign node8943 = (inp[3]) ? node8951 : node8944;
											assign node8944 = (inp[9]) ? 4'b0110 : node8945;
												assign node8945 = (inp[7]) ? 4'b0101 : node8946;
													assign node8946 = (inp[8]) ? 4'b0101 : 4'b0100;
											assign node8951 = (inp[2]) ? node8953 : 4'b0111;
												assign node8953 = (inp[4]) ? 4'b0011 : node8954;
													assign node8954 = (inp[9]) ? 4'b0010 : node8955;
														assign node8955 = (inp[10]) ? 4'b0111 : 4'b0110;
									assign node8960 = (inp[3]) ? node8982 : node8961;
										assign node8961 = (inp[2]) ? node8969 : node8962;
											assign node8962 = (inp[7]) ? node8966 : node8963;
												assign node8963 = (inp[8]) ? 4'b0111 : 4'b0110;
												assign node8966 = (inp[4]) ? 4'b0100 : 4'b0110;
											assign node8969 = (inp[9]) ? node8975 : node8970;
												assign node8970 = (inp[4]) ? 4'b0011 : node8971;
													assign node8971 = (inp[10]) ? 4'b0110 : 4'b0111;
												assign node8975 = (inp[4]) ? 4'b0111 : node8976;
													assign node8976 = (inp[7]) ? 4'b0010 : node8977;
														assign node8977 = (inp[8]) ? 4'b0011 : 4'b0010;
										assign node8982 = (inp[5]) ? node8992 : node8983;
											assign node8983 = (inp[9]) ? node8989 : node8984;
												assign node8984 = (inp[4]) ? node8986 : 4'b0111;
													assign node8986 = (inp[8]) ? 4'b0011 : 4'b0010;
												assign node8989 = (inp[2]) ? 4'b0100 : 4'b0101;
											assign node8992 = (inp[10]) ? node8994 : 4'b0101;
												assign node8994 = (inp[2]) ? node8996 : 4'b0000;
													assign node8996 = (inp[4]) ? node8998 : 4'b0100;
														assign node8998 = (inp[9]) ? 4'b0100 : 4'b0000;
								assign node9001 = (inp[3]) ? node9053 : node9002;
									assign node9002 = (inp[15]) ? node9030 : node9003;
										assign node9003 = (inp[4]) ? node9019 : node9004;
											assign node9004 = (inp[10]) ? node9012 : node9005;
												assign node9005 = (inp[9]) ? node9007 : 4'b0100;
													assign node9007 = (inp[8]) ? node9009 : 4'b0000;
														assign node9009 = (inp[2]) ? 4'b0000 : 4'b0001;
												assign node9012 = (inp[9]) ? node9014 : 4'b0000;
													assign node9014 = (inp[7]) ? 4'b0101 : node9015;
														assign node9015 = (inp[5]) ? 4'b0110 : 4'b0100;
											assign node9019 = (inp[9]) ? node9027 : node9020;
												assign node9020 = (inp[10]) ? node9022 : 4'b0000;
													assign node9022 = (inp[2]) ? 4'b0101 : node9023;
														assign node9023 = (inp[8]) ? 4'b0111 : 4'b0110;
												assign node9027 = (inp[2]) ? 4'b0101 : 4'b0111;
										assign node9030 = (inp[5]) ? node9044 : node9031;
											assign node9031 = (inp[9]) ? node9037 : node9032;
												assign node9032 = (inp[2]) ? 4'b0110 : node9033;
													assign node9033 = (inp[10]) ? 4'b0010 : 4'b0110;
												assign node9037 = (inp[8]) ? node9041 : node9038;
													assign node9038 = (inp[7]) ? 4'b0011 : 4'b0010;
													assign node9041 = (inp[7]) ? 4'b0110 : 4'b0011;
											assign node9044 = (inp[10]) ? node9046 : 4'b0110;
												assign node9046 = (inp[7]) ? node9050 : node9047;
													assign node9047 = (inp[8]) ? 4'b0001 : 4'b0100;
													assign node9050 = (inp[9]) ? 4'b0101 : 4'b0011;
									assign node9053 = (inp[4]) ? node9073 : node9054;
										assign node9054 = (inp[8]) ? node9062 : node9055;
											assign node9055 = (inp[7]) ? node9057 : 4'b0010;
												assign node9057 = (inp[5]) ? 4'b0011 : node9058;
													assign node9058 = (inp[15]) ? 4'b0011 : 4'b0001;
											assign node9062 = (inp[7]) ? node9066 : node9063;
												assign node9063 = (inp[10]) ? 4'b0001 : 4'b0101;
												assign node9066 = (inp[2]) ? node9068 : 4'b0010;
													assign node9068 = (inp[15]) ? 4'b0100 : node9069;
														assign node9069 = (inp[5]) ? 4'b0010 : 4'b0000;
										assign node9073 = (inp[8]) ? node9087 : node9074;
											assign node9074 = (inp[7]) ? node9082 : node9075;
												assign node9075 = (inp[9]) ? node9079 : node9076;
													assign node9076 = (inp[10]) ? 4'b0110 : 4'b0000;
													assign node9079 = (inp[10]) ? 4'b0000 : 4'b0100;
												assign node9082 = (inp[9]) ? node9084 : 4'b0111;
													assign node9084 = (inp[5]) ? 4'b0001 : 4'b0101;
											assign node9087 = (inp[15]) ? node9091 : node9088;
												assign node9088 = (inp[5]) ? 4'b0011 : 4'b0001;
												assign node9091 = (inp[2]) ? 4'b0101 : node9092;
													assign node9092 = (inp[10]) ? node9094 : 4'b0001;
														assign node9094 = (inp[9]) ? 4'b0001 : 4'b0101;
							assign node9098 = (inp[7]) ? node9186 : node9099;
								assign node9099 = (inp[8]) ? node9143 : node9100;
									assign node9100 = (inp[10]) ? node9118 : node9101;
										assign node9101 = (inp[2]) ? node9109 : node9102;
											assign node9102 = (inp[5]) ? node9106 : node9103;
												assign node9103 = (inp[15]) ? 4'b0010 : 4'b0000;
												assign node9106 = (inp[4]) ? 4'b0100 : 4'b0110;
											assign node9109 = (inp[3]) ? node9113 : node9110;
												assign node9110 = (inp[12]) ? 4'b0100 : 4'b0000;
												assign node9113 = (inp[9]) ? 4'b0100 : node9114;
													assign node9114 = (inp[4]) ? 4'b0000 : 4'b0100;
										assign node9118 = (inp[3]) ? node9126 : node9119;
											assign node9119 = (inp[15]) ? 4'b0010 : node9120;
												assign node9120 = (inp[9]) ? node9122 : 4'b0000;
													assign node9122 = (inp[2]) ? 4'b0100 : 4'b0000;
											assign node9126 = (inp[15]) ? node9134 : node9127;
												assign node9127 = (inp[5]) ? node9129 : 4'b0000;
													assign node9129 = (inp[4]) ? node9131 : 4'b0010;
														assign node9131 = (inp[2]) ? 4'b0010 : 4'b0110;
												assign node9134 = (inp[12]) ? node9136 : 4'b0110;
													assign node9136 = (inp[9]) ? node9140 : node9137;
														assign node9137 = (inp[5]) ? 4'b0000 : 4'b0010;
														assign node9140 = (inp[4]) ? 4'b0000 : 4'b0100;
									assign node9143 = (inp[12]) ? node9165 : node9144;
										assign node9144 = (inp[2]) ? node9156 : node9145;
											assign node9145 = (inp[3]) ? node9151 : node9146;
												assign node9146 = (inp[5]) ? 4'b1111 : node9147;
													assign node9147 = (inp[15]) ? 4'b1111 : 4'b1101;
												assign node9151 = (inp[5]) ? node9153 : 4'b1111;
													assign node9153 = (inp[15]) ? 4'b1101 : 4'b1111;
											assign node9156 = (inp[15]) ? node9160 : node9157;
												assign node9157 = (inp[9]) ? 4'b1011 : 4'b1001;
												assign node9160 = (inp[3]) ? 4'b1101 : node9161;
													assign node9161 = (inp[9]) ? 4'b1011 : 4'b1111;
										assign node9165 = (inp[2]) ? node9175 : node9166;
											assign node9166 = (inp[9]) ? node9172 : node9167;
												assign node9167 = (inp[15]) ? node9169 : 4'b1001;
													assign node9169 = (inp[10]) ? 4'b1011 : 4'b1001;
												assign node9172 = (inp[4]) ? 4'b1011 : 4'b1111;
											assign node9175 = (inp[15]) ? node9181 : node9176;
												assign node9176 = (inp[3]) ? node9178 : 4'b1101;
													assign node9178 = (inp[9]) ? 4'b1011 : 4'b1111;
												assign node9181 = (inp[4]) ? node9183 : 4'b1101;
													assign node9183 = (inp[9]) ? 4'b1001 : 4'b1101;
								assign node9186 = (inp[8]) ? node9236 : node9187;
									assign node9187 = (inp[10]) ? node9223 : node9188;
										assign node9188 = (inp[9]) ? node9206 : node9189;
											assign node9189 = (inp[12]) ? node9199 : node9190;
												assign node9190 = (inp[4]) ? node9194 : node9191;
													assign node9191 = (inp[15]) ? 4'b1111 : 4'b1101;
													assign node9194 = (inp[2]) ? node9196 : 4'b1011;
														assign node9196 = (inp[5]) ? 4'b1001 : 4'b1011;
												assign node9199 = (inp[4]) ? 4'b1101 : node9200;
													assign node9200 = (inp[5]) ? node9202 : 4'b1001;
														assign node9202 = (inp[2]) ? 4'b1011 : 4'b1001;
											assign node9206 = (inp[15]) ? node9214 : node9207;
												assign node9207 = (inp[3]) ? node9209 : 4'b1001;
													assign node9209 = (inp[5]) ? 4'b1111 : node9210;
														assign node9210 = (inp[2]) ? 4'b1111 : 4'b1001;
												assign node9214 = (inp[5]) ? node9218 : node9215;
													assign node9215 = (inp[3]) ? 4'b1101 : 4'b1111;
													assign node9218 = (inp[3]) ? 4'b1101 : node9219;
														assign node9219 = (inp[4]) ? 4'b1001 : 4'b1101;
										assign node9223 = (inp[15]) ? node9229 : node9224;
											assign node9224 = (inp[5]) ? 4'b1111 : node9225;
												assign node9225 = (inp[3]) ? 4'b1011 : 4'b1001;
											assign node9229 = (inp[5]) ? node9231 : 4'b1111;
												assign node9231 = (inp[4]) ? 4'b1001 : node9232;
													assign node9232 = (inp[9]) ? 4'b1101 : 4'b1001;
									assign node9236 = (inp[15]) ? node9258 : node9237;
										assign node9237 = (inp[3]) ? node9249 : node9238;
											assign node9238 = (inp[5]) ? node9242 : node9239;
												assign node9239 = (inp[4]) ? 4'b1100 : 4'b1000;
												assign node9242 = (inp[4]) ? node9244 : 4'b1000;
													assign node9244 = (inp[12]) ? 4'b1010 : node9245;
														assign node9245 = (inp[10]) ? 4'b1010 : 4'b1110;
											assign node9249 = (inp[12]) ? 4'b1110 : node9250;
												assign node9250 = (inp[2]) ? node9252 : 4'b1000;
													assign node9252 = (inp[5]) ? node9254 : 4'b1010;
														assign node9254 = (inp[4]) ? 4'b1110 : 4'b1010;
										assign node9258 = (inp[12]) ? node9266 : node9259;
											assign node9259 = (inp[9]) ? 4'b1100 : node9260;
												assign node9260 = (inp[4]) ? 4'b1100 : node9261;
													assign node9261 = (inp[3]) ? 4'b1000 : 4'b1010;
											assign node9266 = (inp[4]) ? node9272 : node9267;
												assign node9267 = (inp[9]) ? node9269 : 4'b1010;
													assign node9269 = (inp[3]) ? 4'b1100 : 4'b1110;
												assign node9272 = (inp[5]) ? 4'b1000 : node9273;
													assign node9273 = (inp[3]) ? 4'b1000 : 4'b1010;
						assign node9277 = (inp[7]) ? node9423 : node9278;
							assign node9278 = (inp[8]) ? node9358 : node9279;
								assign node9279 = (inp[1]) ? node9315 : node9280;
									assign node9280 = (inp[4]) ? node9294 : node9281;
										assign node9281 = (inp[15]) ? node9287 : node9282;
											assign node9282 = (inp[5]) ? node9284 : 4'b0000;
												assign node9284 = (inp[10]) ? 4'b0000 : 4'b0010;
											assign node9287 = (inp[9]) ? 4'b0010 : node9288;
												assign node9288 = (inp[12]) ? node9290 : 4'b0100;
													assign node9290 = (inp[10]) ? 4'b0010 : 4'b0110;
										assign node9294 = (inp[5]) ? node9306 : node9295;
											assign node9295 = (inp[2]) ? node9301 : node9296;
												assign node9296 = (inp[10]) ? 4'b0110 : node9297;
													assign node9297 = (inp[12]) ? 4'b0100 : 4'b0110;
												assign node9301 = (inp[9]) ? 4'b0100 : node9302;
													assign node9302 = (inp[10]) ? 4'b0100 : 4'b0000;
											assign node9306 = (inp[9]) ? 4'b0110 : node9307;
												assign node9307 = (inp[15]) ? 4'b0000 : node9308;
													assign node9308 = (inp[12]) ? 4'b0110 : node9309;
														assign node9309 = (inp[2]) ? 4'b0000 : 4'b0010;
									assign node9315 = (inp[10]) ? node9347 : node9316;
										assign node9316 = (inp[2]) ? node9336 : node9317;
											assign node9317 = (inp[3]) ? node9325 : node9318;
												assign node9318 = (inp[12]) ? 4'b1110 : node9319;
													assign node9319 = (inp[15]) ? node9321 : 4'b1100;
														assign node9321 = (inp[4]) ? 4'b1100 : 4'b1010;
												assign node9325 = (inp[15]) ? node9333 : node9326;
													assign node9326 = (inp[9]) ? node9330 : node9327;
														assign node9327 = (inp[5]) ? 4'b1010 : 4'b1000;
														assign node9330 = (inp[4]) ? 4'b1010 : 4'b1110;
													assign node9333 = (inp[9]) ? 4'b1000 : 4'b1100;
											assign node9336 = (inp[3]) ? node9342 : node9337;
												assign node9337 = (inp[15]) ? 4'b1010 : node9338;
													assign node9338 = (inp[4]) ? 4'b1110 : 4'b1000;
												assign node9342 = (inp[12]) ? 4'b1100 : node9343;
													assign node9343 = (inp[9]) ? 4'b1010 : 4'b1110;
										assign node9347 = (inp[15]) ? node9353 : node9348;
											assign node9348 = (inp[12]) ? node9350 : 4'b1110;
												assign node9350 = (inp[4]) ? 4'b1010 : 4'b1110;
											assign node9353 = (inp[3]) ? 4'b1100 : node9354;
												assign node9354 = (inp[5]) ? 4'b1010 : 4'b1110;
								assign node9358 = (inp[3]) ? node9400 : node9359;
									assign node9359 = (inp[9]) ? node9377 : node9360;
										assign node9360 = (inp[15]) ? node9366 : node9361;
											assign node9361 = (inp[5]) ? node9363 : 4'b1101;
												assign node9363 = (inp[1]) ? 4'b1001 : 4'b1111;
											assign node9366 = (inp[12]) ? node9372 : node9367;
												assign node9367 = (inp[10]) ? node9369 : 4'b1011;
													assign node9369 = (inp[4]) ? 4'b1111 : 4'b1011;
												assign node9372 = (inp[2]) ? node9374 : 4'b1011;
													assign node9374 = (inp[5]) ? 4'b1101 : 4'b1111;
										assign node9377 = (inp[1]) ? node9387 : node9378;
											assign node9378 = (inp[5]) ? node9380 : 4'b1001;
												assign node9380 = (inp[10]) ? 4'b1011 : node9381;
													assign node9381 = (inp[2]) ? node9383 : 4'b1001;
														assign node9383 = (inp[15]) ? 4'b1011 : 4'b1001;
											assign node9387 = (inp[4]) ? node9393 : node9388;
												assign node9388 = (inp[12]) ? 4'b1111 : node9389;
													assign node9389 = (inp[10]) ? 4'b1101 : 4'b1001;
												assign node9393 = (inp[12]) ? node9395 : 4'b1101;
													assign node9395 = (inp[15]) ? 4'b1001 : node9396;
														assign node9396 = (inp[5]) ? 4'b1011 : 4'b1001;
									assign node9400 = (inp[15]) ? node9410 : node9401;
										assign node9401 = (inp[4]) ? 4'b1111 : node9402;
											assign node9402 = (inp[5]) ? node9406 : node9403;
												assign node9403 = (inp[10]) ? 4'b1001 : 4'b1101;
												assign node9406 = (inp[9]) ? 4'b1111 : 4'b1011;
										assign node9410 = (inp[10]) ? node9418 : node9411;
											assign node9411 = (inp[5]) ? 4'b1101 : node9412;
												assign node9412 = (inp[2]) ? node9414 : 4'b1101;
													assign node9414 = (inp[1]) ? 4'b1111 : 4'b1011;
											assign node9418 = (inp[1]) ? 4'b1101 : node9419;
												assign node9419 = (inp[4]) ? 4'b1001 : 4'b1101;
							assign node9423 = (inp[8]) ? node9489 : node9424;
								assign node9424 = (inp[15]) ? node9460 : node9425;
									assign node9425 = (inp[5]) ? node9441 : node9426;
										assign node9426 = (inp[3]) ? node9434 : node9427;
											assign node9427 = (inp[2]) ? node9429 : 4'b1101;
												assign node9429 = (inp[12]) ? node9431 : 4'b1001;
													assign node9431 = (inp[4]) ? 4'b1101 : 4'b1001;
											assign node9434 = (inp[1]) ? 4'b1001 : node9435;
												assign node9435 = (inp[4]) ? node9437 : 4'b1111;
													assign node9437 = (inp[10]) ? 4'b1011 : 4'b1111;
										assign node9441 = (inp[10]) ? node9449 : node9442;
											assign node9442 = (inp[4]) ? 4'b1111 : node9443;
												assign node9443 = (inp[12]) ? node9445 : 4'b1001;
													assign node9445 = (inp[9]) ? 4'b1111 : 4'b1011;
											assign node9449 = (inp[2]) ? node9451 : 4'b1111;
												assign node9451 = (inp[1]) ? 4'b1011 : node9452;
													assign node9452 = (inp[4]) ? node9456 : node9453;
														assign node9453 = (inp[9]) ? 4'b1111 : 4'b1011;
														assign node9456 = (inp[3]) ? 4'b1111 : 4'b1011;
									assign node9460 = (inp[3]) ? node9476 : node9461;
										assign node9461 = (inp[9]) ? node9471 : node9462;
											assign node9462 = (inp[10]) ? node9466 : node9463;
												assign node9463 = (inp[2]) ? 4'b1111 : 4'b1011;
												assign node9466 = (inp[5]) ? 4'b1101 : node9467;
													assign node9467 = (inp[12]) ? 4'b1111 : 4'b1011;
											assign node9471 = (inp[4]) ? 4'b1001 : node9472;
												assign node9472 = (inp[12]) ? 4'b1101 : 4'b1011;
										assign node9476 = (inp[5]) ? node9484 : node9477;
											assign node9477 = (inp[10]) ? node9479 : 4'b1011;
												assign node9479 = (inp[9]) ? node9481 : 4'b1101;
													assign node9481 = (inp[4]) ? 4'b1001 : 4'b1101;
											assign node9484 = (inp[2]) ? node9486 : 4'b1101;
												assign node9486 = (inp[1]) ? 4'b1001 : 4'b1101;
								assign node9489 = (inp[15]) ? node9539 : node9490;
									assign node9490 = (inp[10]) ? node9516 : node9491;
										assign node9491 = (inp[5]) ? node9505 : node9492;
											assign node9492 = (inp[12]) ? node9500 : node9493;
												assign node9493 = (inp[4]) ? node9497 : node9494;
													assign node9494 = (inp[9]) ? 4'b1000 : 4'b1100;
													assign node9497 = (inp[9]) ? 4'b1100 : 4'b1000;
												assign node9500 = (inp[3]) ? 4'b1110 : node9501;
													assign node9501 = (inp[2]) ? 4'b1100 : 4'b1000;
											assign node9505 = (inp[3]) ? 4'b1110 : node9506;
												assign node9506 = (inp[9]) ? 4'b1110 : node9507;
													assign node9507 = (inp[12]) ? node9511 : node9508;
														assign node9508 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node9511 = (inp[1]) ? 4'b1000 : 4'b1110;
										assign node9516 = (inp[3]) ? node9530 : node9517;
											assign node9517 = (inp[2]) ? node9523 : node9518;
												assign node9518 = (inp[1]) ? node9520 : 4'b1000;
													assign node9520 = (inp[12]) ? 4'b1000 : 4'b1100;
												assign node9523 = (inp[9]) ? node9527 : node9524;
													assign node9524 = (inp[4]) ? 4'b1100 : 4'b1000;
													assign node9527 = (inp[4]) ? 4'b1010 : 4'b1110;
											assign node9530 = (inp[4]) ? node9536 : node9531;
												assign node9531 = (inp[9]) ? 4'b1110 : node9532;
													assign node9532 = (inp[5]) ? 4'b1010 : 4'b1000;
												assign node9536 = (inp[9]) ? 4'b1010 : 4'b1110;
									assign node9539 = (inp[3]) ? node9551 : node9540;
										assign node9540 = (inp[9]) ? node9542 : 4'b1010;
											assign node9542 = (inp[5]) ? node9546 : node9543;
												assign node9543 = (inp[4]) ? 4'b1010 : 4'b1110;
												assign node9546 = (inp[1]) ? 4'b1100 : node9547;
													assign node9547 = (inp[10]) ? 4'b1000 : 4'b1010;
										assign node9551 = (inp[9]) ? node9563 : node9552;
											assign node9552 = (inp[4]) ? node9556 : node9553;
												assign node9553 = (inp[12]) ? 4'b1010 : 4'b1110;
												assign node9556 = (inp[2]) ? node9558 : 4'b1100;
													assign node9558 = (inp[10]) ? 4'b1100 : node9559;
														assign node9559 = (inp[12]) ? 4'b1100 : 4'b1000;
											assign node9563 = (inp[2]) ? node9569 : node9564;
												assign node9564 = (inp[4]) ? 4'b1000 : node9565;
													assign node9565 = (inp[10]) ? 4'b1100 : 4'b1000;
												assign node9569 = (inp[10]) ? 4'b1000 : 4'b1010;
				assign node9572 = (inp[6]) ? node10214 : node9573;
					assign node9573 = (inp[13]) ? node9923 : node9574;
						assign node9574 = (inp[1]) ? node9778 : node9575;
							assign node9575 = (inp[10]) ? node9663 : node9576;
								assign node9576 = (inp[5]) ? node9610 : node9577;
									assign node9577 = (inp[15]) ? node9597 : node9578;
										assign node9578 = (inp[3]) ? node9586 : node9579;
											assign node9579 = (inp[4]) ? node9581 : 4'b0001;
												assign node9581 = (inp[2]) ? node9583 : 4'b0001;
													assign node9583 = (inp[12]) ? 4'b0101 : 4'b0100;
											assign node9586 = (inp[4]) ? node9592 : node9587;
												assign node9587 = (inp[9]) ? node9589 : 4'b0100;
													assign node9589 = (inp[2]) ? 4'b0001 : 4'b0000;
												assign node9592 = (inp[9]) ? node9594 : 4'b0001;
													assign node9594 = (inp[12]) ? 4'b0110 : 4'b0111;
										assign node9597 = (inp[7]) ? node9603 : node9598;
											assign node9598 = (inp[8]) ? 4'b0111 : node9599;
												assign node9599 = (inp[3]) ? 4'b0010 : 4'b0110;
											assign node9603 = (inp[8]) ? 4'b0010 : node9604;
												assign node9604 = (inp[4]) ? node9606 : 4'b0011;
													assign node9606 = (inp[9]) ? 4'b0101 : 4'b0011;
									assign node9610 = (inp[15]) ? node9642 : node9611;
										assign node9611 = (inp[3]) ? node9625 : node9612;
											assign node9612 = (inp[12]) ? node9618 : node9613;
												assign node9613 = (inp[9]) ? 4'b0001 : node9614;
													assign node9614 = (inp[4]) ? 4'b0001 : 4'b0101;
												assign node9618 = (inp[9]) ? 4'b0110 : node9619;
													assign node9619 = (inp[4]) ? node9621 : 4'b0100;
														assign node9621 = (inp[7]) ? 4'b0001 : 4'b0000;
											assign node9625 = (inp[2]) ? node9635 : node9626;
												assign node9626 = (inp[4]) ? node9630 : node9627;
													assign node9627 = (inp[12]) ? 4'b0110 : 4'b0011;
													assign node9630 = (inp[8]) ? node9632 : 4'b0011;
														assign node9632 = (inp[7]) ? 4'b0010 : 4'b0011;
												assign node9635 = (inp[12]) ? node9637 : 4'b0110;
													assign node9637 = (inp[9]) ? 4'b0111 : node9638;
														assign node9638 = (inp[4]) ? 4'b0011 : 4'b0111;
										assign node9642 = (inp[4]) ? node9656 : node9643;
											assign node9643 = (inp[9]) ? node9649 : node9644;
												assign node9644 = (inp[12]) ? 4'b0101 : node9645;
													assign node9645 = (inp[8]) ? 4'b0100 : 4'b0110;
												assign node9649 = (inp[3]) ? node9651 : 4'b0011;
													assign node9651 = (inp[7]) ? node9653 : 4'b0000;
														assign node9653 = (inp[8]) ? 4'b0000 : 4'b0001;
											assign node9656 = (inp[7]) ? node9660 : node9657;
												assign node9657 = (inp[9]) ? 4'b0100 : 4'b0000;
												assign node9660 = (inp[8]) ? 4'b0100 : 4'b0101;
								assign node9663 = (inp[9]) ? node9721 : node9664;
									assign node9664 = (inp[8]) ? node9692 : node9665;
										assign node9665 = (inp[7]) ? node9681 : node9666;
											assign node9666 = (inp[3]) ? node9672 : node9667;
												assign node9667 = (inp[4]) ? 4'b0110 : node9668;
													assign node9668 = (inp[12]) ? 4'b0010 : 4'b0110;
												assign node9672 = (inp[5]) ? node9676 : node9673;
													assign node9673 = (inp[12]) ? 4'b0000 : 4'b0100;
													assign node9676 = (inp[15]) ? 4'b0000 : node9677;
														assign node9677 = (inp[12]) ? 4'b0110 : 4'b0010;
											assign node9681 = (inp[12]) ? node9685 : node9682;
												assign node9682 = (inp[15]) ? 4'b0011 : 4'b0001;
												assign node9685 = (inp[4]) ? node9687 : 4'b0011;
													assign node9687 = (inp[3]) ? node9689 : 4'b0101;
														assign node9689 = (inp[15]) ? 4'b0101 : 4'b0111;
										assign node9692 = (inp[7]) ? node9710 : node9693;
											assign node9693 = (inp[2]) ? node9705 : node9694;
												assign node9694 = (inp[5]) ? node9700 : node9695;
													assign node9695 = (inp[4]) ? 4'b0111 : node9696;
														assign node9696 = (inp[15]) ? 4'b0111 : 4'b0001;
													assign node9700 = (inp[3]) ? node9702 : 4'b0011;
														assign node9702 = (inp[4]) ? 4'b0011 : 4'b0001;
												assign node9705 = (inp[15]) ? 4'b0101 : node9706;
													assign node9706 = (inp[3]) ? 4'b0011 : 4'b0001;
											assign node9710 = (inp[15]) ? node9718 : node9711;
												assign node9711 = (inp[3]) ? node9713 : 4'b0100;
													assign node9713 = (inp[4]) ? 4'b0000 : node9714;
														assign node9714 = (inp[2]) ? 4'b0000 : 4'b0100;
												assign node9718 = (inp[12]) ? 4'b0010 : 4'b0100;
									assign node9721 = (inp[15]) ? node9757 : node9722;
										assign node9722 = (inp[3]) ? node9734 : node9723;
											assign node9723 = (inp[12]) ? node9731 : node9724;
												assign node9724 = (inp[4]) ? 4'b0100 : node9725;
													assign node9725 = (inp[8]) ? 4'b0000 : node9726;
														assign node9726 = (inp[7]) ? 4'b0001 : 4'b0000;
												assign node9731 = (inp[8]) ? 4'b0010 : 4'b0110;
											assign node9734 = (inp[12]) ? node9744 : node9735;
												assign node9735 = (inp[4]) ? node9739 : node9736;
													assign node9736 = (inp[5]) ? 4'b0010 : 4'b0000;
													assign node9739 = (inp[7]) ? node9741 : 4'b0110;
														assign node9741 = (inp[8]) ? 4'b0110 : 4'b0111;
												assign node9744 = (inp[4]) ? node9750 : node9745;
													assign node9745 = (inp[7]) ? node9747 : 4'b0111;
														assign node9747 = (inp[8]) ? 4'b0110 : 4'b0111;
													assign node9750 = (inp[8]) ? node9754 : node9751;
														assign node9751 = (inp[7]) ? 4'b0011 : 4'b0010;
														assign node9754 = (inp[7]) ? 4'b0010 : 4'b0011;
										assign node9757 = (inp[5]) ? node9767 : node9758;
											assign node9758 = (inp[4]) ? node9764 : node9759;
												assign node9759 = (inp[12]) ? 4'b0111 : node9760;
													assign node9760 = (inp[2]) ? 4'b0011 : 4'b0010;
												assign node9764 = (inp[3]) ? 4'b0100 : 4'b0111;
											assign node9767 = (inp[4]) ? node9773 : node9768;
												assign node9768 = (inp[8]) ? node9770 : 4'b0101;
													assign node9770 = (inp[3]) ? 4'b0001 : 4'b0010;
												assign node9773 = (inp[8]) ? node9775 : 4'b0000;
													assign node9775 = (inp[7]) ? 4'b0000 : 4'b0001;
							assign node9778 = (inp[8]) ? node9850 : node9779;
								assign node9779 = (inp[7]) ? node9825 : node9780;
									assign node9780 = (inp[2]) ? node9804 : node9781;
										assign node9781 = (inp[12]) ? node9797 : node9782;
											assign node9782 = (inp[15]) ? node9790 : node9783;
												assign node9783 = (inp[5]) ? 4'b0110 : node9784;
													assign node9784 = (inp[3]) ? 4'b0000 : node9785;
														assign node9785 = (inp[9]) ? 4'b0000 : 4'b0100;
												assign node9790 = (inp[9]) ? node9792 : 4'b0110;
													assign node9792 = (inp[4]) ? 4'b0100 : node9793;
														assign node9793 = (inp[3]) ? 4'b0000 : 4'b0010;
											assign node9797 = (inp[9]) ? 4'b0000 : node9798;
												assign node9798 = (inp[4]) ? node9800 : 4'b0110;
													assign node9800 = (inp[5]) ? 4'b0000 : 4'b0010;
										assign node9804 = (inp[15]) ? node9814 : node9805;
											assign node9805 = (inp[4]) ? node9809 : node9806;
												assign node9806 = (inp[12]) ? 4'b0000 : 4'b0100;
												assign node9809 = (inp[12]) ? 4'b0110 : node9810;
													assign node9810 = (inp[3]) ? 4'b0110 : 4'b0100;
											assign node9814 = (inp[3]) ? node9820 : node9815;
												assign node9815 = (inp[9]) ? 4'b0010 : node9816;
													assign node9816 = (inp[12]) ? 4'b0010 : 4'b0110;
												assign node9820 = (inp[5]) ? 4'b0100 : node9821;
													assign node9821 = (inp[9]) ? 4'b0010 : 4'b0110;
									assign node9825 = (inp[2]) ? node9843 : node9826;
										assign node9826 = (inp[9]) ? node9834 : node9827;
											assign node9827 = (inp[15]) ? node9831 : node9828;
												assign node9828 = (inp[3]) ? 4'b1011 : 4'b1001;
												assign node9831 = (inp[4]) ? 4'b1111 : 4'b1011;
											assign node9834 = (inp[15]) ? node9840 : node9835;
												assign node9835 = (inp[5]) ? node9837 : 4'b1111;
													assign node9837 = (inp[4]) ? 4'b1111 : 4'b1011;
												assign node9840 = (inp[4]) ? 4'b1111 : 4'b1101;
										assign node9843 = (inp[10]) ? 4'b1101 : node9844;
											assign node9844 = (inp[15]) ? node9846 : 4'b1111;
												assign node9846 = (inp[4]) ? 4'b1001 : 4'b1011;
								assign node9850 = (inp[7]) ? node9888 : node9851;
									assign node9851 = (inp[2]) ? node9865 : node9852;
										assign node9852 = (inp[5]) ? node9860 : node9853;
											assign node9853 = (inp[4]) ? node9855 : 4'b1001;
												assign node9855 = (inp[12]) ? node9857 : 4'b1011;
													assign node9857 = (inp[10]) ? 4'b1111 : 4'b1011;
											assign node9860 = (inp[15]) ? node9862 : 4'b1011;
												assign node9862 = (inp[4]) ? 4'b1001 : 4'b1101;
										assign node9865 = (inp[10]) ? node9879 : node9866;
											assign node9866 = (inp[5]) ? node9876 : node9867;
												assign node9867 = (inp[12]) ? node9871 : node9868;
													assign node9868 = (inp[15]) ? 4'b1011 : 4'b1001;
													assign node9871 = (inp[15]) ? node9873 : 4'b1111;
														assign node9873 = (inp[9]) ? 4'b1001 : 4'b1111;
												assign node9876 = (inp[12]) ? 4'b1101 : 4'b1111;
											assign node9879 = (inp[15]) ? node9885 : node9880;
												assign node9880 = (inp[9]) ? node9882 : 4'b1111;
													assign node9882 = (inp[4]) ? 4'b1011 : 4'b1111;
												assign node9885 = (inp[9]) ? 4'b1101 : 4'b1011;
									assign node9888 = (inp[9]) ? node9904 : node9889;
										assign node9889 = (inp[15]) ? node9899 : node9890;
											assign node9890 = (inp[5]) ? node9896 : node9891;
												assign node9891 = (inp[3]) ? 4'b1000 : node9892;
													assign node9892 = (inp[10]) ? 4'b1000 : 4'b1100;
												assign node9896 = (inp[3]) ? 4'b1010 : 4'b1000;
											assign node9899 = (inp[4]) ? node9901 : 4'b1010;
												assign node9901 = (inp[3]) ? 4'b1100 : 4'b1010;
										assign node9904 = (inp[4]) ? node9916 : node9905;
											assign node9905 = (inp[12]) ? node9911 : node9906;
												assign node9906 = (inp[2]) ? node9908 : 4'b1000;
													assign node9908 = (inp[10]) ? 4'b1110 : 4'b1010;
												assign node9911 = (inp[15]) ? 4'b1100 : node9912;
													assign node9912 = (inp[3]) ? 4'b1110 : 4'b1100;
											assign node9916 = (inp[10]) ? node9920 : node9917;
												assign node9917 = (inp[12]) ? 4'b1010 : 4'b1110;
												assign node9920 = (inp[12]) ? 4'b1010 : 4'b1000;
						assign node9923 = (inp[7]) ? node10063 : node9924;
							assign node9924 = (inp[8]) ? node9994 : node9925;
								assign node9925 = (inp[1]) ? node9963 : node9926;
									assign node9926 = (inp[4]) ? node9948 : node9927;
										assign node9927 = (inp[9]) ? node9939 : node9928;
											assign node9928 = (inp[5]) ? node9930 : 4'b0110;
												assign node9930 = (inp[10]) ? node9932 : 4'b0100;
													assign node9932 = (inp[12]) ? node9936 : node9933;
														assign node9933 = (inp[2]) ? 4'b0100 : 4'b0110;
														assign node9936 = (inp[3]) ? 4'b0000 : 4'b0000;
											assign node9939 = (inp[3]) ? node9943 : node9940;
												assign node9940 = (inp[12]) ? 4'b0110 : 4'b0010;
												assign node9943 = (inp[5]) ? node9945 : 4'b0000;
													assign node9945 = (inp[15]) ? 4'b0000 : 4'b0010;
										assign node9948 = (inp[9]) ? node9958 : node9949;
											assign node9949 = (inp[12]) ? node9955 : node9950;
												assign node9950 = (inp[3]) ? node9952 : 4'b0010;
													assign node9952 = (inp[15]) ? 4'b0000 : 4'b0010;
												assign node9955 = (inp[15]) ? 4'b0010 : 4'b0000;
											assign node9958 = (inp[10]) ? 4'b0010 : node9959;
												assign node9959 = (inp[2]) ? 4'b0110 : 4'b0100;
									assign node9963 = (inp[3]) ? node9985 : node9964;
										assign node9964 = (inp[15]) ? node9978 : node9965;
											assign node9965 = (inp[5]) ? node9971 : node9966;
												assign node9966 = (inp[4]) ? 4'b1000 : node9967;
													assign node9967 = (inp[9]) ? 4'b1100 : 4'b1000;
												assign node9971 = (inp[2]) ? node9973 : 4'b1000;
													assign node9973 = (inp[10]) ? node9975 : 4'b1010;
														assign node9975 = (inp[4]) ? 4'b1110 : 4'b1000;
											assign node9978 = (inp[5]) ? 4'b1000 : node9979;
												assign node9979 = (inp[2]) ? node9981 : 4'b1110;
													assign node9981 = (inp[10]) ? 4'b1110 : 4'b1010;
										assign node9985 = (inp[15]) ? node9987 : 4'b1110;
											assign node9987 = (inp[9]) ? node9991 : node9988;
												assign node9988 = (inp[12]) ? 4'b1010 : 4'b1100;
												assign node9991 = (inp[5]) ? 4'b1000 : 4'b1100;
								assign node9994 = (inp[4]) ? node10032 : node9995;
									assign node9995 = (inp[9]) ? node10015 : node9996;
										assign node9996 = (inp[15]) ? node10008 : node9997;
											assign node9997 = (inp[10]) ? node10003 : node9998;
												assign node9998 = (inp[12]) ? node10000 : 4'b1101;
													assign node10000 = (inp[5]) ? 4'b1011 : 4'b1001;
												assign node10003 = (inp[5]) ? node10005 : 4'b1001;
													assign node10005 = (inp[3]) ? 4'b1011 : 4'b1001;
											assign node10008 = (inp[10]) ? 4'b1011 : node10009;
												assign node10009 = (inp[12]) ? 4'b1011 : node10010;
													assign node10010 = (inp[5]) ? 4'b1101 : 4'b1111;
										assign node10015 = (inp[12]) ? node10021 : node10016;
											assign node10016 = (inp[10]) ? 4'b1111 : node10017;
												assign node10017 = (inp[5]) ? 4'b1001 : 4'b1011;
											assign node10021 = (inp[15]) ? node10027 : node10022;
												assign node10022 = (inp[3]) ? 4'b1111 : node10023;
													assign node10023 = (inp[5]) ? 4'b1111 : 4'b1101;
												assign node10027 = (inp[3]) ? 4'b1101 : node10028;
													assign node10028 = (inp[5]) ? 4'b1101 : 4'b1111;
									assign node10032 = (inp[9]) ? node10050 : node10033;
										assign node10033 = (inp[10]) ? node10041 : node10034;
											assign node10034 = (inp[12]) ? 4'b1101 : node10035;
												assign node10035 = (inp[3]) ? node10037 : 4'b1011;
													assign node10037 = (inp[5]) ? 4'b1011 : 4'b1001;
											assign node10041 = (inp[3]) ? 4'b1111 : node10042;
												assign node10042 = (inp[1]) ? node10044 : 4'b1111;
													assign node10044 = (inp[5]) ? node10046 : 4'b1101;
														assign node10046 = (inp[12]) ? 4'b1111 : 4'b1101;
										assign node10050 = (inp[15]) ? node10056 : node10051;
											assign node10051 = (inp[12]) ? 4'b1011 : node10052;
												assign node10052 = (inp[10]) ? 4'b1011 : 4'b1111;
											assign node10056 = (inp[5]) ? node10060 : node10057;
												assign node10057 = (inp[3]) ? 4'b1001 : 4'b1011;
												assign node10060 = (inp[12]) ? 4'b1001 : 4'b1101;
							assign node10063 = (inp[8]) ? node10139 : node10064;
								assign node10064 = (inp[15]) ? node10098 : node10065;
									assign node10065 = (inp[3]) ? node10077 : node10066;
										assign node10066 = (inp[4]) ? node10068 : 4'b1001;
											assign node10068 = (inp[9]) ? node10072 : node10069;
												assign node10069 = (inp[12]) ? 4'b1111 : 4'b1001;
												assign node10072 = (inp[12]) ? 4'b1011 : node10073;
													assign node10073 = (inp[10]) ? 4'b1011 : 4'b1111;
										assign node10077 = (inp[5]) ? node10087 : node10078;
											assign node10078 = (inp[10]) ? node10080 : 4'b1001;
												assign node10080 = (inp[9]) ? node10084 : node10081;
													assign node10081 = (inp[4]) ? 4'b1111 : 4'b1001;
													assign node10084 = (inp[2]) ? 4'b1111 : 4'b1011;
											assign node10087 = (inp[9]) ? node10093 : node10088;
												assign node10088 = (inp[4]) ? node10090 : 4'b1011;
													assign node10090 = (inp[12]) ? 4'b1111 : 4'b1011;
												assign node10093 = (inp[10]) ? 4'b1111 : node10094;
													assign node10094 = (inp[4]) ? 4'b1111 : 4'b1011;
									assign node10098 = (inp[5]) ? node10122 : node10099;
										assign node10099 = (inp[3]) ? node10113 : node10100;
											assign node10100 = (inp[1]) ? node10106 : node10101;
												assign node10101 = (inp[9]) ? node10103 : 4'b1111;
													assign node10103 = (inp[4]) ? 4'b1011 : 4'b1111;
												assign node10106 = (inp[2]) ? node10108 : 4'b1011;
													assign node10108 = (inp[10]) ? 4'b1011 : node10109;
														assign node10109 = (inp[12]) ? 4'b1011 : 4'b1111;
											assign node10113 = (inp[9]) ? 4'b1101 : node10114;
												assign node10114 = (inp[2]) ? 4'b1101 : node10115;
													assign node10115 = (inp[10]) ? 4'b1011 : node10116;
														assign node10116 = (inp[12]) ? 4'b1011 : 4'b1111;
										assign node10122 = (inp[3]) ? node10130 : node10123;
											assign node10123 = (inp[4]) ? node10127 : node10124;
												assign node10124 = (inp[9]) ? 4'b1011 : 4'b1111;
												assign node10127 = (inp[1]) ? 4'b1001 : 4'b1101;
											assign node10130 = (inp[12]) ? 4'b1001 : node10131;
												assign node10131 = (inp[1]) ? node10133 : 4'b1001;
													assign node10133 = (inp[4]) ? node10135 : 4'b1101;
														assign node10135 = (inp[10]) ? 4'b1101 : 4'b1001;
								assign node10139 = (inp[4]) ? node10179 : node10140;
									assign node10140 = (inp[9]) ? node10158 : node10141;
										assign node10141 = (inp[10]) ? node10151 : node10142;
											assign node10142 = (inp[12]) ? node10148 : node10143;
												assign node10143 = (inp[15]) ? 4'b1110 : node10144;
													assign node10144 = (inp[3]) ? 4'b1110 : 4'b1100;
												assign node10148 = (inp[3]) ? 4'b1000 : 4'b1010;
											assign node10151 = (inp[1]) ? node10155 : node10152;
												assign node10152 = (inp[2]) ? 4'b1010 : 4'b1000;
												assign node10155 = (inp[2]) ? 4'b1000 : 4'b1010;
										assign node10158 = (inp[12]) ? node10170 : node10159;
											assign node10159 = (inp[10]) ? node10167 : node10160;
												assign node10160 = (inp[3]) ? node10162 : 4'b1000;
													assign node10162 = (inp[2]) ? node10164 : 4'b1010;
														assign node10164 = (inp[5]) ? 4'b1000 : 4'b1010;
												assign node10167 = (inp[15]) ? 4'b1100 : 4'b1110;
											assign node10170 = (inp[2]) ? node10172 : 4'b1100;
												assign node10172 = (inp[5]) ? 4'b1100 : node10173;
													assign node10173 = (inp[3]) ? node10175 : 4'b1110;
														assign node10175 = (inp[15]) ? 4'b1100 : 4'b1110;
									assign node10179 = (inp[1]) ? node10205 : node10180;
										assign node10180 = (inp[3]) ? node10194 : node10181;
											assign node10181 = (inp[15]) ? node10191 : node10182;
												assign node10182 = (inp[5]) ? node10188 : node10183;
													assign node10183 = (inp[10]) ? 4'b1000 : node10184;
														assign node10184 = (inp[9]) ? 4'b1100 : 4'b1000;
													assign node10188 = (inp[10]) ? 4'b1110 : 4'b1000;
												assign node10191 = (inp[10]) ? 4'b1000 : 4'b1010;
											assign node10194 = (inp[15]) ? node10200 : node10195;
												assign node10195 = (inp[12]) ? 4'b1110 : node10196;
													assign node10196 = (inp[9]) ? 4'b1110 : 4'b1000;
												assign node10200 = (inp[10]) ? 4'b1100 : node10201;
													assign node10201 = (inp[5]) ? 4'b1100 : 4'b1010;
										assign node10205 = (inp[10]) ? node10207 : 4'b1110;
											assign node10207 = (inp[9]) ? 4'b1000 : node10208;
												assign node10208 = (inp[15]) ? node10210 : 4'b1110;
													assign node10210 = (inp[5]) ? 4'b1100 : 4'b1110;
					assign node10214 = (inp[1]) ? node10586 : node10215;
						assign node10215 = (inp[13]) ? node10407 : node10216;
							assign node10216 = (inp[15]) ? node10328 : node10217;
								assign node10217 = (inp[3]) ? node10265 : node10218;
									assign node10218 = (inp[5]) ? node10248 : node10219;
										assign node10219 = (inp[10]) ? node10239 : node10220;
											assign node10220 = (inp[9]) ? node10230 : node10221;
												assign node10221 = (inp[8]) ? node10225 : node10222;
													assign node10222 = (inp[7]) ? 4'b1101 : 4'b1000;
													assign node10225 = (inp[12]) ? 4'b1101 : node10226;
														assign node10226 = (inp[4]) ? 4'b1001 : 4'b1101;
												assign node10230 = (inp[4]) ? node10236 : node10231;
													assign node10231 = (inp[2]) ? node10233 : 4'b1100;
														assign node10233 = (inp[7]) ? 4'b1000 : 4'b1001;
													assign node10236 = (inp[12]) ? 4'b1001 : 4'b1100;
											assign node10239 = (inp[4]) ? node10243 : node10240;
												assign node10240 = (inp[9]) ? 4'b1101 : 4'b1001;
												assign node10243 = (inp[9]) ? node10245 : 4'b1100;
													assign node10245 = (inp[12]) ? 4'b1001 : 4'b1000;
										assign node10248 = (inp[4]) ? node10258 : node10249;
											assign node10249 = (inp[10]) ? 4'b1000 : node10250;
												assign node10250 = (inp[12]) ? 4'b1111 : node10251;
													assign node10251 = (inp[9]) ? node10253 : 4'b1100;
														assign node10253 = (inp[8]) ? 4'b1001 : 4'b1000;
											assign node10258 = (inp[8]) ? node10262 : node10259;
												assign node10259 = (inp[7]) ? 4'b1011 : 4'b1010;
												assign node10262 = (inp[9]) ? 4'b1111 : 4'b1110;
									assign node10265 = (inp[5]) ? node10299 : node10266;
										assign node10266 = (inp[9]) ? node10282 : node10267;
											assign node10267 = (inp[4]) ? node10275 : node10268;
												assign node10268 = (inp[2]) ? 4'b1001 : node10269;
													assign node10269 = (inp[10]) ? node10271 : 4'b1001;
														assign node10271 = (inp[12]) ? 4'b1000 : 4'b1000;
												assign node10275 = (inp[12]) ? node10277 : 4'b1001;
													assign node10277 = (inp[2]) ? node10279 : 4'b1111;
														assign node10279 = (inp[7]) ? 4'b1110 : 4'b1110;
											assign node10282 = (inp[4]) ? node10292 : node10283;
												assign node10283 = (inp[10]) ? node10287 : node10284;
													assign node10284 = (inp[12]) ? 4'b1110 : 4'b1000;
													assign node10287 = (inp[7]) ? 4'b1111 : node10288;
														assign node10288 = (inp[8]) ? 4'b1111 : 4'b1110;
												assign node10292 = (inp[7]) ? 4'b1010 : node10293;
													assign node10293 = (inp[8]) ? node10295 : 4'b1010;
														assign node10295 = (inp[10]) ? 4'b1011 : 4'b1111;
										assign node10299 = (inp[10]) ? node10313 : node10300;
											assign node10300 = (inp[9]) ? node10306 : node10301;
												assign node10301 = (inp[12]) ? node10303 : 4'b1110;
													assign node10303 = (inp[2]) ? 4'b1011 : 4'b1010;
												assign node10306 = (inp[12]) ? node10310 : node10307;
													assign node10307 = (inp[4]) ? 4'b1111 : 4'b1011;
													assign node10310 = (inp[7]) ? 4'b1010 : 4'b1011;
											assign node10313 = (inp[12]) ? node10321 : node10314;
												assign node10314 = (inp[7]) ? node10316 : 4'b1010;
													assign node10316 = (inp[4]) ? node10318 : 4'b1110;
														assign node10318 = (inp[9]) ? 4'b1010 : 4'b1110;
												assign node10321 = (inp[9]) ? node10325 : node10322;
													assign node10322 = (inp[2]) ? 4'b1011 : 4'b1111;
													assign node10325 = (inp[4]) ? 4'b1011 : 4'b1110;
								assign node10328 = (inp[5]) ? node10360 : node10329;
									assign node10329 = (inp[3]) ? node10347 : node10330;
										assign node10330 = (inp[12]) ? node10340 : node10331;
											assign node10331 = (inp[4]) ? node10335 : node10332;
												assign node10332 = (inp[2]) ? 4'b1010 : 4'b1011;
												assign node10335 = (inp[9]) ? 4'b1111 : node10336;
													assign node10336 = (inp[10]) ? 4'b1110 : 4'b1010;
											assign node10340 = (inp[10]) ? 4'b1011 : node10341;
												assign node10341 = (inp[8]) ? node10343 : 4'b1111;
													assign node10343 = (inp[2]) ? 4'b1111 : 4'b1110;
										assign node10347 = (inp[8]) ? node10353 : node10348;
											assign node10348 = (inp[12]) ? node10350 : 4'b1100;
												assign node10350 = (inp[7]) ? 4'b1001 : 4'b1000;
											assign node10353 = (inp[2]) ? 4'b1011 : node10354;
												assign node10354 = (inp[4]) ? node10356 : 4'b1010;
													assign node10356 = (inp[7]) ? 4'b1100 : 4'b1101;
									assign node10360 = (inp[3]) ? node10378 : node10361;
										assign node10361 = (inp[12]) ? node10367 : node10362;
											assign node10362 = (inp[10]) ? 4'b1101 : node10363;
												assign node10363 = (inp[4]) ? 4'b1010 : 4'b1111;
											assign node10367 = (inp[4]) ? node10371 : node10368;
												assign node10368 = (inp[9]) ? 4'b1100 : 4'b1010;
												assign node10371 = (inp[9]) ? 4'b1000 : node10372;
													assign node10372 = (inp[2]) ? node10374 : 4'b1100;
														assign node10374 = (inp[8]) ? 4'b1100 : 4'b1101;
										assign node10378 = (inp[9]) ? node10386 : node10379;
											assign node10379 = (inp[10]) ? 4'b1000 : node10380;
												assign node10380 = (inp[2]) ? 4'b1001 : node10381;
													assign node10381 = (inp[4]) ? 4'b1101 : 4'b1001;
											assign node10386 = (inp[4]) ? node10400 : node10387;
												assign node10387 = (inp[10]) ? node10395 : node10388;
													assign node10388 = (inp[12]) ? node10392 : node10389;
														assign node10389 = (inp[8]) ? 4'b1000 : 4'b1000;
														assign node10392 = (inp[7]) ? 4'b1100 : 4'b1101;
													assign node10395 = (inp[2]) ? 4'b1101 : node10396;
														assign node10396 = (inp[7]) ? 4'b1101 : 4'b1100;
												assign node10400 = (inp[10]) ? node10402 : 4'b1100;
													assign node10402 = (inp[7]) ? 4'b1000 : node10403;
														assign node10403 = (inp[8]) ? 4'b1001 : 4'b1000;
							assign node10407 = (inp[8]) ? node10483 : node10408;
								assign node10408 = (inp[7]) ? node10444 : node10409;
									assign node10409 = (inp[4]) ? node10429 : node10410;
										assign node10410 = (inp[10]) ? node10422 : node10411;
											assign node10411 = (inp[15]) ? node10413 : 4'b1000;
												assign node10413 = (inp[12]) ? node10417 : node10414;
													assign node10414 = (inp[9]) ? 4'b1010 : 4'b1110;
													assign node10417 = (inp[5]) ? node10419 : 4'b1010;
														assign node10419 = (inp[2]) ? 4'b1000 : 4'b1010;
											assign node10422 = (inp[9]) ? node10426 : node10423;
												assign node10423 = (inp[2]) ? 4'b1000 : 4'b1010;
												assign node10426 = (inp[12]) ? 4'b1100 : 4'b1110;
										assign node10429 = (inp[9]) ? node10435 : node10430;
											assign node10430 = (inp[12]) ? 4'b1100 : node10431;
												assign node10431 = (inp[10]) ? 4'b1100 : 4'b1000;
											assign node10435 = (inp[15]) ? node10439 : node10436;
												assign node10436 = (inp[3]) ? 4'b1010 : 4'b1000;
												assign node10439 = (inp[12]) ? 4'b1000 : node10440;
													assign node10440 = (inp[2]) ? 4'b1000 : 4'b1100;
									assign node10444 = (inp[10]) ? node10462 : node10445;
										assign node10445 = (inp[2]) ? 4'b0111 : node10446;
											assign node10446 = (inp[12]) ? node10456 : node10447;
												assign node10447 = (inp[5]) ? node10451 : node10448;
													assign node10448 = (inp[15]) ? 4'b0111 : 4'b0101;
													assign node10451 = (inp[3]) ? 4'b0011 : node10452;
														assign node10452 = (inp[4]) ? 4'b0011 : 4'b0111;
												assign node10456 = (inp[5]) ? 4'b0101 : node10457;
													assign node10457 = (inp[15]) ? 4'b0011 : 4'b0001;
										assign node10462 = (inp[15]) ? node10468 : node10463;
											assign node10463 = (inp[5]) ? node10465 : 4'b0001;
												assign node10465 = (inp[12]) ? 4'b0111 : 4'b0001;
											assign node10468 = (inp[5]) ? node10476 : node10469;
												assign node10469 = (inp[9]) ? 4'b0001 : node10470;
													assign node10470 = (inp[4]) ? node10472 : 4'b0011;
														assign node10472 = (inp[12]) ? 4'b0101 : 4'b0111;
												assign node10476 = (inp[2]) ? node10478 : 4'b0001;
													assign node10478 = (inp[12]) ? node10480 : 4'b0101;
														assign node10480 = (inp[4]) ? 4'b0001 : 4'b0101;
								assign node10483 = (inp[7]) ? node10547 : node10484;
									assign node10484 = (inp[5]) ? node10518 : node10485;
										assign node10485 = (inp[3]) ? node10497 : node10486;
											assign node10486 = (inp[15]) ? node10490 : node10487;
												assign node10487 = (inp[2]) ? 4'b0101 : 4'b0001;
												assign node10490 = (inp[12]) ? node10492 : 4'b0011;
													assign node10492 = (inp[10]) ? 4'b0011 : node10493;
														assign node10493 = (inp[2]) ? 4'b0111 : 4'b0011;
											assign node10497 = (inp[9]) ? node10507 : node10498;
												assign node10498 = (inp[2]) ? node10504 : node10499;
													assign node10499 = (inp[15]) ? node10501 : 4'b0101;
														assign node10501 = (inp[12]) ? 4'b0101 : 4'b0111;
													assign node10504 = (inp[4]) ? 4'b0111 : 4'b0011;
												assign node10507 = (inp[15]) ? node10513 : node10508;
													assign node10508 = (inp[4]) ? node10510 : 4'b0001;
														assign node10510 = (inp[10]) ? 4'b0011 : 4'b0011;
													assign node10513 = (inp[2]) ? node10515 : 4'b0101;
														assign node10515 = (inp[4]) ? 4'b0101 : 4'b0011;
										assign node10518 = (inp[15]) ? node10530 : node10519;
											assign node10519 = (inp[3]) ? node10527 : node10520;
												assign node10520 = (inp[4]) ? node10522 : 4'b0001;
													assign node10522 = (inp[12]) ? 4'b0111 : node10523;
														assign node10523 = (inp[9]) ? 4'b0011 : 4'b0001;
												assign node10527 = (inp[10]) ? 4'b0111 : 4'b0011;
											assign node10530 = (inp[3]) ? node10536 : node10531;
												assign node10531 = (inp[2]) ? node10533 : 4'b0101;
													assign node10533 = (inp[12]) ? 4'b0101 : 4'b0011;
												assign node10536 = (inp[12]) ? node10542 : node10537;
													assign node10537 = (inp[2]) ? 4'b0101 : node10538;
														assign node10538 = (inp[4]) ? 4'b0001 : 4'b0101;
													assign node10542 = (inp[4]) ? node10544 : 4'b0001;
														assign node10544 = (inp[9]) ? 4'b0001 : 4'b0101;
									assign node10547 = (inp[10]) ? node10563 : node10548;
										assign node10548 = (inp[12]) ? node10554 : node10549;
											assign node10549 = (inp[9]) ? 4'b0110 : node10550;
												assign node10550 = (inp[4]) ? 4'b0000 : 4'b0100;
											assign node10554 = (inp[5]) ? node10560 : node10555;
												assign node10555 = (inp[2]) ? 4'b0000 : node10556;
													assign node10556 = (inp[4]) ? 4'b0000 : 4'b0100;
												assign node10560 = (inp[2]) ? 4'b0110 : 4'b0010;
										assign node10563 = (inp[3]) ? node10577 : node10564;
											assign node10564 = (inp[4]) ? node10572 : node10565;
												assign node10565 = (inp[9]) ? node10567 : 4'b0010;
													assign node10567 = (inp[2]) ? node10569 : 4'b0110;
														assign node10569 = (inp[5]) ? 4'b0110 : 4'b0100;
												assign node10572 = (inp[9]) ? node10574 : 4'b0110;
													assign node10574 = (inp[12]) ? 4'b0010 : 4'b0000;
											assign node10577 = (inp[15]) ? node10583 : node10578;
												assign node10578 = (inp[12]) ? node10580 : 4'b0010;
													assign node10580 = (inp[5]) ? 4'b0010 : 4'b0000;
												assign node10583 = (inp[2]) ? 4'b0100 : 4'b0000;
						assign node10586 = (inp[8]) ? node10718 : node10587;
							assign node10587 = (inp[7]) ? node10653 : node10588;
								assign node10588 = (inp[13]) ? node10632 : node10589;
									assign node10589 = (inp[5]) ? node10615 : node10590;
										assign node10590 = (inp[12]) ? node10602 : node10591;
											assign node10591 = (inp[10]) ? node10595 : node10592;
												assign node10592 = (inp[15]) ? 4'b1110 : 4'b1100;
												assign node10595 = (inp[4]) ? node10599 : node10596;
													assign node10596 = (inp[15]) ? 4'b1010 : 4'b1000;
													assign node10599 = (inp[9]) ? 4'b1010 : 4'b1110;
											assign node10602 = (inp[2]) ? node10610 : node10603;
												assign node10603 = (inp[15]) ? node10607 : node10604;
													assign node10604 = (inp[3]) ? 4'b1110 : 4'b1100;
													assign node10607 = (inp[3]) ? 4'b1100 : 4'b1110;
												assign node10610 = (inp[9]) ? node10612 : 4'b1010;
													assign node10612 = (inp[4]) ? 4'b1000 : 4'b1100;
										assign node10615 = (inp[4]) ? node10627 : node10616;
											assign node10616 = (inp[10]) ? node10618 : 4'b1010;
												assign node10618 = (inp[2]) ? node10624 : node10619;
													assign node10619 = (inp[15]) ? node10621 : 4'b1000;
														assign node10621 = (inp[3]) ? 4'b1000 : 4'b1010;
													assign node10624 = (inp[3]) ? 4'b1010 : 4'b1000;
											assign node10627 = (inp[10]) ? node10629 : 4'b1000;
												assign node10629 = (inp[9]) ? 4'b1010 : 4'b1100;
									assign node10632 = (inp[5]) ? node10644 : node10633;
										assign node10633 = (inp[3]) ? node10639 : node10634;
											assign node10634 = (inp[15]) ? 4'b0010 : node10635;
												assign node10635 = (inp[12]) ? 4'b0100 : 4'b0000;
											assign node10639 = (inp[4]) ? 4'b0000 : node10640;
												assign node10640 = (inp[15]) ? 4'b0100 : 4'b0000;
										assign node10644 = (inp[15]) ? node10650 : node10645;
											assign node10645 = (inp[12]) ? 4'b0110 : node10646;
												assign node10646 = (inp[9]) ? 4'b0110 : 4'b0010;
											assign node10650 = (inp[2]) ? 4'b0100 : 4'b0000;
								assign node10653 = (inp[4]) ? node10699 : node10654;
									assign node10654 = (inp[2]) ? node10680 : node10655;
										assign node10655 = (inp[12]) ? node10669 : node10656;
											assign node10656 = (inp[9]) ? node10664 : node10657;
												assign node10657 = (inp[10]) ? 4'b0001 : node10658;
													assign node10658 = (inp[15]) ? node10660 : 4'b0101;
														assign node10660 = (inp[5]) ? 4'b0101 : 4'b0111;
												assign node10664 = (inp[5]) ? node10666 : 4'b0001;
													assign node10666 = (inp[15]) ? 4'b0001 : 4'b0011;
											assign node10669 = (inp[9]) ? node10673 : node10670;
												assign node10670 = (inp[15]) ? 4'b0011 : 4'b0001;
												assign node10673 = (inp[13]) ? node10675 : 4'b0101;
													assign node10675 = (inp[3]) ? 4'b0101 : node10676;
														assign node10676 = (inp[15]) ? 4'b0111 : 4'b0101;
										assign node10680 = (inp[9]) ? node10690 : node10681;
											assign node10681 = (inp[10]) ? node10687 : node10682;
												assign node10682 = (inp[12]) ? node10684 : 4'b0111;
													assign node10684 = (inp[5]) ? 4'b0001 : 4'b0011;
												assign node10687 = (inp[12]) ? 4'b0011 : 4'b0001;
											assign node10690 = (inp[10]) ? node10696 : node10691;
												assign node10691 = (inp[12]) ? 4'b0111 : node10692;
													assign node10692 = (inp[15]) ? 4'b0011 : 4'b0001;
												assign node10696 = (inp[15]) ? 4'b0101 : 4'b0111;
									assign node10699 = (inp[15]) ? node10709 : node10700;
										assign node10700 = (inp[2]) ? node10704 : node10701;
											assign node10701 = (inp[5]) ? 4'b0011 : 4'b0001;
											assign node10704 = (inp[9]) ? node10706 : 4'b0111;
												assign node10706 = (inp[12]) ? 4'b0011 : 4'b0111;
										assign node10709 = (inp[5]) ? node10715 : node10710;
											assign node10710 = (inp[3]) ? node10712 : 4'b0011;
												assign node10712 = (inp[9]) ? 4'b0001 : 4'b0011;
											assign node10715 = (inp[9]) ? 4'b0001 : 4'b0101;
							assign node10718 = (inp[7]) ? node10792 : node10719;
								assign node10719 = (inp[5]) ? node10771 : node10720;
									assign node10720 = (inp[3]) ? node10744 : node10721;
										assign node10721 = (inp[15]) ? node10741 : node10722;
											assign node10722 = (inp[13]) ? node10734 : node10723;
												assign node10723 = (inp[12]) ? node10729 : node10724;
													assign node10724 = (inp[9]) ? 4'b0001 : node10725;
														assign node10725 = (inp[4]) ? 4'b0001 : 4'b0001;
													assign node10729 = (inp[9]) ? 4'b0101 : node10730;
														assign node10730 = (inp[4]) ? 4'b0101 : 4'b0001;
												assign node10734 = (inp[2]) ? node10736 : 4'b0101;
													assign node10736 = (inp[10]) ? 4'b0101 : node10737;
														assign node10737 = (inp[12]) ? 4'b0101 : 4'b0001;
											assign node10741 = (inp[10]) ? 4'b0111 : 4'b0011;
										assign node10744 = (inp[12]) ? node10760 : node10745;
											assign node10745 = (inp[13]) ? node10755 : node10746;
												assign node10746 = (inp[9]) ? node10748 : 4'b0001;
													assign node10748 = (inp[15]) ? node10752 : node10749;
														assign node10749 = (inp[10]) ? 4'b0011 : 4'b0111;
														assign node10752 = (inp[10]) ? 4'b0101 : 4'b0011;
												assign node10755 = (inp[15]) ? node10757 : 4'b0111;
													assign node10757 = (inp[9]) ? 4'b0101 : 4'b0111;
											assign node10760 = (inp[13]) ? 4'b0011 : node10761;
												assign node10761 = (inp[4]) ? node10765 : node10762;
													assign node10762 = (inp[15]) ? 4'b0011 : 4'b0001;
													assign node10765 = (inp[15]) ? node10767 : 4'b0111;
														assign node10767 = (inp[2]) ? 4'b0001 : 4'b0101;
									assign node10771 = (inp[15]) ? node10783 : node10772;
										assign node10772 = (inp[4]) ? node10776 : node10773;
											assign node10773 = (inp[2]) ? 4'b0001 : 4'b0011;
											assign node10776 = (inp[10]) ? node10780 : node10777;
												assign node10777 = (inp[2]) ? 4'b0111 : 4'b0011;
												assign node10780 = (inp[9]) ? 4'b0011 : 4'b0111;
										assign node10783 = (inp[4]) ? node10787 : node10784;
											assign node10784 = (inp[3]) ? 4'b0001 : 4'b0011;
											assign node10787 = (inp[10]) ? 4'b0001 : node10788;
												assign node10788 = (inp[13]) ? 4'b0001 : 4'b0101;
								assign node10792 = (inp[15]) ? node10852 : node10793;
									assign node10793 = (inp[3]) ? node10827 : node10794;
										assign node10794 = (inp[5]) ? node10816 : node10795;
											assign node10795 = (inp[2]) ? node10805 : node10796;
												assign node10796 = (inp[9]) ? node10798 : 4'b0100;
													assign node10798 = (inp[10]) ? node10802 : node10799;
														assign node10799 = (inp[13]) ? 4'b0000 : 4'b0100;
														assign node10802 = (inp[12]) ? 4'b0100 : 4'b0000;
												assign node10805 = (inp[10]) ? node10811 : node10806;
													assign node10806 = (inp[12]) ? 4'b0100 : node10807;
														assign node10807 = (inp[4]) ? 4'b0000 : 4'b0100;
													assign node10811 = (inp[12]) ? 4'b0000 : node10812;
														assign node10812 = (inp[9]) ? 4'b0100 : 4'b0000;
											assign node10816 = (inp[4]) ? node10824 : node10817;
												assign node10817 = (inp[12]) ? 4'b0000 : node10818;
													assign node10818 = (inp[9]) ? 4'b0000 : node10819;
														assign node10819 = (inp[10]) ? 4'b0000 : 4'b0100;
												assign node10824 = (inp[13]) ? 4'b0110 : 4'b0010;
										assign node10827 = (inp[5]) ? node10841 : node10828;
											assign node10828 = (inp[4]) ? node10834 : node10829;
												assign node10829 = (inp[13]) ? node10831 : 4'b0000;
													assign node10831 = (inp[2]) ? 4'b0100 : 4'b0000;
												assign node10834 = (inp[12]) ? 4'b0010 : node10835;
													assign node10835 = (inp[13]) ? 4'b0110 : node10836;
														assign node10836 = (inp[9]) ? 4'b0010 : 4'b0110;
											assign node10841 = (inp[10]) ? node10843 : 4'b0010;
												assign node10843 = (inp[2]) ? node10849 : node10844;
													assign node10844 = (inp[4]) ? node10846 : 4'b0110;
														assign node10846 = (inp[9]) ? 4'b0010 : 4'b0110;
													assign node10849 = (inp[9]) ? 4'b0110 : 4'b0010;
									assign node10852 = (inp[3]) ? node10870 : node10853;
										assign node10853 = (inp[5]) ? node10861 : node10854;
											assign node10854 = (inp[12]) ? node10856 : 4'b0110;
												assign node10856 = (inp[4]) ? node10858 : 4'b0010;
													assign node10858 = (inp[9]) ? 4'b0010 : 4'b0110;
											assign node10861 = (inp[9]) ? node10867 : node10862;
												assign node10862 = (inp[4]) ? 4'b0100 : node10863;
													assign node10863 = (inp[10]) ? 4'b0010 : 4'b0110;
												assign node10867 = (inp[4]) ? 4'b0000 : 4'b0100;
										assign node10870 = (inp[12]) ? 4'b0100 : node10871;
											assign node10871 = (inp[4]) ? node10879 : node10872;
												assign node10872 = (inp[2]) ? node10874 : 4'b0100;
													assign node10874 = (inp[13]) ? node10876 : 4'b0000;
														assign node10876 = (inp[9]) ? 4'b0100 : 4'b0000;
												assign node10879 = (inp[5]) ? node10881 : 4'b0000;
													assign node10881 = (inp[10]) ? 4'b0100 : 4'b0000;

endmodule