module dtc_split05_bm89 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node9;
	wire [3-1:0] node10;
	wire [3-1:0] node13;
	wire [3-1:0] node16;
	wire [3-1:0] node17;
	wire [3-1:0] node18;
	wire [3-1:0] node21;
	wire [3-1:0] node24;
	wire [3-1:0] node26;
	wire [3-1:0] node29;
	wire [3-1:0] node30;
	wire [3-1:0] node32;
	wire [3-1:0] node34;
	wire [3-1:0] node37;
	wire [3-1:0] node38;
	wire [3-1:0] node39;
	wire [3-1:0] node42;
	wire [3-1:0] node45;
	wire [3-1:0] node46;
	wire [3-1:0] node49;
	wire [3-1:0] node52;
	wire [3-1:0] node53;
	wire [3-1:0] node54;
	wire [3-1:0] node55;
	wire [3-1:0] node56;
	wire [3-1:0] node59;
	wire [3-1:0] node62;
	wire [3-1:0] node64;
	wire [3-1:0] node67;
	wire [3-1:0] node68;
	wire [3-1:0] node69;
	wire [3-1:0] node72;
	wire [3-1:0] node75;
	wire [3-1:0] node76;
	wire [3-1:0] node79;
	wire [3-1:0] node82;
	wire [3-1:0] node84;
	wire [3-1:0] node85;
	wire [3-1:0] node86;
	wire [3-1:0] node89;
	wire [3-1:0] node92;
	wire [3-1:0] node93;
	wire [3-1:0] node96;

	assign outp = (inp[6]) ? node52 : node1;
		assign node1 = (inp[9]) ? node29 : node2;
			assign node2 = (inp[3]) ? node16 : node3;
				assign node3 = (inp[8]) ? node9 : node4;
					assign node4 = (inp[5]) ? 3'b011 : node5;
						assign node5 = (inp[7]) ? 3'b100 : 3'b101;
					assign node9 = (inp[0]) ? node13 : node10;
						assign node10 = (inp[10]) ? 3'b010 : 3'b100;
						assign node13 = (inp[10]) ? 3'b101 : 3'b000;
				assign node16 = (inp[7]) ? node24 : node17;
					assign node17 = (inp[10]) ? node21 : node18;
						assign node18 = (inp[4]) ? 3'b000 : 3'b100;
						assign node21 = (inp[4]) ? 3'b100 : 3'b011;
					assign node24 = (inp[10]) ? node26 : 3'b000;
						assign node26 = (inp[0]) ? 3'b000 : 3'b000;
			assign node29 = (inp[7]) ? node37 : node30;
				assign node30 = (inp[3]) ? node32 : 3'b111;
					assign node32 = (inp[10]) ? node34 : 3'b010;
						assign node34 = (inp[8]) ? 3'b001 : 3'b011;
				assign node37 = (inp[4]) ? node45 : node38;
					assign node38 = (inp[10]) ? node42 : node39;
						assign node39 = (inp[5]) ? 3'b110 : 3'b010;
						assign node42 = (inp[3]) ? 3'b001 : 3'b100;
					assign node45 = (inp[8]) ? node49 : node46;
						assign node46 = (inp[5]) ? 3'b010 : 3'b001;
						assign node49 = (inp[3]) ? 3'b110 : 3'b111;
		assign node52 = (inp[3]) ? node82 : node53;
			assign node53 = (inp[9]) ? node67 : node54;
				assign node54 = (inp[4]) ? node62 : node55;
					assign node55 = (inp[11]) ? node59 : node56;
						assign node56 = (inp[0]) ? 3'b100 : 3'b000;
						assign node59 = (inp[5]) ? 3'b010 : 3'b110;
					assign node62 = (inp[10]) ? node64 : 3'b000;
						assign node64 = (inp[7]) ? 3'b000 : 3'b010;
				assign node67 = (inp[4]) ? node75 : node68;
					assign node68 = (inp[7]) ? node72 : node69;
						assign node69 = (inp[8]) ? 3'b001 : 3'b011;
						assign node72 = (inp[11]) ? 3'b101 : 3'b000;
					assign node75 = (inp[10]) ? node79 : node76;
						assign node76 = (inp[7]) ? 3'b010 : 3'b010;
						assign node79 = (inp[7]) ? 3'b110 : 3'b101;
			assign node82 = (inp[9]) ? node84 : 3'b000;
				assign node84 = (inp[11]) ? node92 : node85;
					assign node85 = (inp[0]) ? node89 : node86;
						assign node86 = (inp[10]) ? 3'b100 : 3'b000;
						assign node89 = (inp[2]) ? 3'b000 : 3'b000;
					assign node92 = (inp[4]) ? node96 : node93;
						assign node93 = (inp[5]) ? 3'b000 : 3'b010;
						assign node96 = (inp[5]) ? 3'b000 : 3'b000;

endmodule