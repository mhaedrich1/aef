module dtc_split125_bm80 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node9;
	wire [3-1:0] node11;
	wire [3-1:0] node14;
	wire [3-1:0] node15;
	wire [3-1:0] node16;
	wire [3-1:0] node20;
	wire [3-1:0] node21;
	wire [3-1:0] node24;
	wire [3-1:0] node27;
	wire [3-1:0] node28;
	wire [3-1:0] node29;
	wire [3-1:0] node31;
	wire [3-1:0] node34;
	wire [3-1:0] node35;
	wire [3-1:0] node39;
	wire [3-1:0] node40;
	wire [3-1:0] node41;
	wire [3-1:0] node44;
	wire [3-1:0] node47;
	wire [3-1:0] node49;
	wire [3-1:0] node52;
	wire [3-1:0] node53;
	wire [3-1:0] node54;
	wire [3-1:0] node55;
	wire [3-1:0] node56;
	wire [3-1:0] node59;
	wire [3-1:0] node62;
	wire [3-1:0] node64;
	wire [3-1:0] node67;
	wire [3-1:0] node68;
	wire [3-1:0] node69;
	wire [3-1:0] node73;
	wire [3-1:0] node74;
	wire [3-1:0] node77;
	wire [3-1:0] node80;
	wire [3-1:0] node81;
	wire [3-1:0] node82;
	wire [3-1:0] node84;
	wire [3-1:0] node87;
	wire [3-1:0] node88;
	wire [3-1:0] node91;
	wire [3-1:0] node94;
	wire [3-1:0] node95;
	wire [3-1:0] node98;
	wire [3-1:0] node100;
	wire [3-1:0] node103;
	wire [3-1:0] node104;
	wire [3-1:0] node105;
	wire [3-1:0] node106;
	wire [3-1:0] node107;
	wire [3-1:0] node108;
	wire [3-1:0] node113;
	wire [3-1:0] node115;
	wire [3-1:0] node117;
	wire [3-1:0] node120;
	wire [3-1:0] node121;
	wire [3-1:0] node122;
	wire [3-1:0] node123;
	wire [3-1:0] node126;
	wire [3-1:0] node129;
	wire [3-1:0] node132;
	wire [3-1:0] node133;
	wire [3-1:0] node135;
	wire [3-1:0] node138;
	wire [3-1:0] node139;
	wire [3-1:0] node143;
	wire [3-1:0] node144;
	wire [3-1:0] node145;
	wire [3-1:0] node146;
	wire [3-1:0] node149;
	wire [3-1:0] node151;
	wire [3-1:0] node156;
	wire [3-1:0] node157;
	wire [3-1:0] node158;
	wire [3-1:0] node159;
	wire [3-1:0] node160;
	wire [3-1:0] node161;
	wire [3-1:0] node165;
	wire [3-1:0] node167;
	wire [3-1:0] node168;
	wire [3-1:0] node172;
	wire [3-1:0] node173;
	wire [3-1:0] node174;
	wire [3-1:0] node176;
	wire [3-1:0] node179;
	wire [3-1:0] node182;
	wire [3-1:0] node183;
	wire [3-1:0] node184;
	wire [3-1:0] node187;
	wire [3-1:0] node190;
	wire [3-1:0] node191;
	wire [3-1:0] node194;
	wire [3-1:0] node197;
	wire [3-1:0] node198;
	wire [3-1:0] node199;
	wire [3-1:0] node200;
	wire [3-1:0] node201;
	wire [3-1:0] node204;
	wire [3-1:0] node208;
	wire [3-1:0] node209;
	wire [3-1:0] node210;
	wire [3-1:0] node213;
	wire [3-1:0] node216;
	wire [3-1:0] node217;
	wire [3-1:0] node221;
	wire [3-1:0] node222;
	wire [3-1:0] node223;
	wire [3-1:0] node224;
	wire [3-1:0] node228;
	wire [3-1:0] node229;
	wire [3-1:0] node232;
	wire [3-1:0] node235;
	wire [3-1:0] node236;
	wire [3-1:0] node237;
	wire [3-1:0] node241;
	wire [3-1:0] node243;
	wire [3-1:0] node246;
	wire [3-1:0] node247;
	wire [3-1:0] node248;
	wire [3-1:0] node249;
	wire [3-1:0] node250;
	wire [3-1:0] node251;
	wire [3-1:0] node255;
	wire [3-1:0] node256;
	wire [3-1:0] node259;
	wire [3-1:0] node262;
	wire [3-1:0] node263;
	wire [3-1:0] node264;
	wire [3-1:0] node268;
	wire [3-1:0] node269;
	wire [3-1:0] node273;
	wire [3-1:0] node274;
	wire [3-1:0] node275;
	wire [3-1:0] node277;
	wire [3-1:0] node280;
	wire [3-1:0] node282;
	wire [3-1:0] node285;
	wire [3-1:0] node286;
	wire [3-1:0] node288;
	wire [3-1:0] node291;
	wire [3-1:0] node292;
	wire [3-1:0] node295;
	wire [3-1:0] node298;
	wire [3-1:0] node299;
	wire [3-1:0] node300;
	wire [3-1:0] node301;
	wire [3-1:0] node303;
	wire [3-1:0] node306;
	wire [3-1:0] node307;
	wire [3-1:0] node310;
	wire [3-1:0] node313;
	wire [3-1:0] node314;
	wire [3-1:0] node315;
	wire [3-1:0] node318;
	wire [3-1:0] node321;
	wire [3-1:0] node322;
	wire [3-1:0] node325;
	wire [3-1:0] node328;
	wire [3-1:0] node329;
	wire [3-1:0] node330;
	wire [3-1:0] node331;
	wire [3-1:0] node334;
	wire [3-1:0] node337;
	wire [3-1:0] node339;
	wire [3-1:0] node342;
	wire [3-1:0] node343;
	wire [3-1:0] node344;
	wire [3-1:0] node347;

	assign outp = (inp[6]) ? node156 : node1;
		assign node1 = (inp[3]) ? node103 : node2;
			assign node2 = (inp[9]) ? node52 : node3;
				assign node3 = (inp[7]) ? node27 : node4;
					assign node4 = (inp[2]) ? node14 : node5;
						assign node5 = (inp[1]) ? node9 : node6;
							assign node6 = (inp[0]) ? 3'b010 : 3'b011;
							assign node9 = (inp[4]) ? node11 : 3'b110;
								assign node11 = (inp[0]) ? 3'b000 : 3'b010;
						assign node14 = (inp[4]) ? node20 : node15;
							assign node15 = (inp[8]) ? 3'b001 : node16;
								assign node16 = (inp[0]) ? 3'b010 : 3'b101;
							assign node20 = (inp[5]) ? node24 : node21;
								assign node21 = (inp[11]) ? 3'b110 : 3'b100;
								assign node24 = (inp[8]) ? 3'b000 : 3'b000;
					assign node27 = (inp[0]) ? node39 : node28;
						assign node28 = (inp[10]) ? node34 : node29;
							assign node29 = (inp[2]) ? node31 : 3'b111;
								assign node31 = (inp[1]) ? 3'b001 : 3'b001;
							assign node34 = (inp[1]) ? 3'b101 : node35;
								assign node35 = (inp[2]) ? 3'b001 : 3'b000;
						assign node39 = (inp[4]) ? node47 : node40;
							assign node40 = (inp[11]) ? node44 : node41;
								assign node41 = (inp[8]) ? 3'b001 : 3'b100;
								assign node44 = (inp[10]) ? 3'b110 : 3'b001;
							assign node47 = (inp[2]) ? node49 : 3'b010;
								assign node49 = (inp[5]) ? 3'b010 : 3'b110;
				assign node52 = (inp[4]) ? node80 : node53;
					assign node53 = (inp[5]) ? node67 : node54;
						assign node54 = (inp[0]) ? node62 : node55;
							assign node55 = (inp[7]) ? node59 : node56;
								assign node56 = (inp[2]) ? 3'b010 : 3'b111;
								assign node59 = (inp[11]) ? 3'b001 : 3'b101;
							assign node62 = (inp[8]) ? node64 : 3'b110;
								assign node64 = (inp[10]) ? 3'b110 : 3'b010;
						assign node67 = (inp[0]) ? node73 : node68;
							assign node68 = (inp[1]) ? 3'b010 : node69;
								assign node69 = (inp[11]) ? 3'b000 : 3'b101;
							assign node73 = (inp[7]) ? node77 : node74;
								assign node74 = (inp[10]) ? 3'b100 : 3'b100;
								assign node77 = (inp[1]) ? 3'b000 : 3'b010;
					assign node80 = (inp[5]) ? node94 : node81;
						assign node81 = (inp[1]) ? node87 : node82;
							assign node82 = (inp[11]) ? node84 : 3'b010;
								assign node84 = (inp[2]) ? 3'b000 : 3'b000;
							assign node87 = (inp[2]) ? node91 : node88;
								assign node88 = (inp[10]) ? 3'b000 : 3'b000;
								assign node91 = (inp[10]) ? 3'b000 : 3'b100;
						assign node94 = (inp[10]) ? node98 : node95;
							assign node95 = (inp[11]) ? 3'b000 : 3'b010;
							assign node98 = (inp[8]) ? node100 : 3'b000;
								assign node100 = (inp[1]) ? 3'b000 : 3'b100;
			assign node103 = (inp[9]) ? node143 : node104;
				assign node104 = (inp[7]) ? node120 : node105;
					assign node105 = (inp[5]) ? node113 : node106;
						assign node106 = (inp[4]) ? 3'b000 : node107;
							assign node107 = (inp[8]) ? 3'b100 : node108;
								assign node108 = (inp[10]) ? 3'b000 : 3'b000;
						assign node113 = (inp[8]) ? node115 : 3'b000;
							assign node115 = (inp[1]) ? node117 : 3'b000;
								assign node117 = (inp[0]) ? 3'b000 : 3'b010;
					assign node120 = (inp[4]) ? node132 : node121;
						assign node121 = (inp[5]) ? node129 : node122;
							assign node122 = (inp[1]) ? node126 : node123;
								assign node123 = (inp[11]) ? 3'b010 : 3'b100;
								assign node126 = (inp[11]) ? 3'b100 : 3'b100;
							assign node129 = (inp[1]) ? 3'b000 : 3'b100;
						assign node132 = (inp[10]) ? node138 : node133;
							assign node133 = (inp[8]) ? node135 : 3'b000;
								assign node135 = (inp[0]) ? 3'b100 : 3'b110;
							assign node138 = (inp[0]) ? 3'b000 : node139;
								assign node139 = (inp[5]) ? 3'b000 : 3'b000;
				assign node143 = (inp[10]) ? 3'b000 : node144;
					assign node144 = (inp[4]) ? 3'b000 : node145;
						assign node145 = (inp[1]) ? node149 : node146;
							assign node146 = (inp[0]) ? 3'b000 : 3'b010;
							assign node149 = (inp[7]) ? node151 : 3'b000;
								assign node151 = (inp[11]) ? 3'b000 : 3'b100;
		assign node156 = (inp[3]) ? node246 : node157;
			assign node157 = (inp[9]) ? node197 : node158;
				assign node158 = (inp[0]) ? node172 : node159;
					assign node159 = (inp[4]) ? node165 : node160;
						assign node160 = (inp[8]) ? 3'b111 : node161;
							assign node161 = (inp[2]) ? 3'b111 : 3'b010;
						assign node165 = (inp[1]) ? node167 : 3'b111;
							assign node167 = (inp[11]) ? 3'b101 : node168;
								assign node168 = (inp[10]) ? 3'b101 : 3'b111;
					assign node172 = (inp[4]) ? node182 : node173;
						assign node173 = (inp[7]) ? node179 : node174;
							assign node174 = (inp[5]) ? node176 : 3'b101;
								assign node176 = (inp[8]) ? 3'b011 : 3'b101;
							assign node179 = (inp[11]) ? 3'b011 : 3'b111;
						assign node182 = (inp[1]) ? node190 : node183;
							assign node183 = (inp[11]) ? node187 : node184;
								assign node184 = (inp[2]) ? 3'b011 : 3'b011;
								assign node187 = (inp[8]) ? 3'b011 : 3'b101;
							assign node190 = (inp[5]) ? node194 : node191;
								assign node191 = (inp[2]) ? 3'b001 : 3'b101;
								assign node194 = (inp[7]) ? 3'b001 : 3'b110;
				assign node197 = (inp[0]) ? node221 : node198;
					assign node198 = (inp[7]) ? node208 : node199;
						assign node199 = (inp[2]) ? 3'b001 : node200;
							assign node200 = (inp[5]) ? node204 : node201;
								assign node201 = (inp[11]) ? 3'b001 : 3'b101;
								assign node204 = (inp[8]) ? 3'b110 : 3'b101;
						assign node208 = (inp[4]) ? node216 : node209;
							assign node209 = (inp[2]) ? node213 : node210;
								assign node210 = (inp[8]) ? 3'b111 : 3'b011;
								assign node213 = (inp[5]) ? 3'b111 : 3'b111;
							assign node216 = (inp[2]) ? 3'b011 : node217;
								assign node217 = (inp[8]) ? 3'b101 : 3'b001;
					assign node221 = (inp[11]) ? node235 : node222;
						assign node222 = (inp[10]) ? node228 : node223;
							assign node223 = (inp[2]) ? 3'b001 : node224;
								assign node224 = (inp[4]) ? 3'b001 : 3'b101;
							assign node228 = (inp[8]) ? node232 : node229;
								assign node229 = (inp[4]) ? 3'b100 : 3'b110;
								assign node232 = (inp[4]) ? 3'b100 : 3'b101;
						assign node235 = (inp[4]) ? node241 : node236;
							assign node236 = (inp[5]) ? 3'b110 : node237;
								assign node237 = (inp[10]) ? 3'b010 : 3'b001;
							assign node241 = (inp[7]) ? node243 : 3'b100;
								assign node243 = (inp[8]) ? 3'b000 : 3'b000;
			assign node246 = (inp[9]) ? node298 : node247;
				assign node247 = (inp[7]) ? node273 : node248;
					assign node248 = (inp[4]) ? node262 : node249;
						assign node249 = (inp[1]) ? node255 : node250;
							assign node250 = (inp[2]) ? 3'b101 : node251;
								assign node251 = (inp[0]) ? 3'b100 : 3'b110;
							assign node255 = (inp[0]) ? node259 : node256;
								assign node256 = (inp[5]) ? 3'b101 : 3'b001;
								assign node259 = (inp[8]) ? 3'b110 : 3'b010;
						assign node262 = (inp[0]) ? node268 : node263;
							assign node263 = (inp[8]) ? 3'b110 : node264;
								assign node264 = (inp[1]) ? 3'b000 : 3'b110;
							assign node268 = (inp[1]) ? 3'b100 : node269;
								assign node269 = (inp[8]) ? 3'b110 : 3'b100;
					assign node273 = (inp[0]) ? node285 : node274;
						assign node274 = (inp[4]) ? node280 : node275;
							assign node275 = (inp[1]) ? node277 : 3'b111;
								assign node277 = (inp[10]) ? 3'b001 : 3'b101;
							assign node280 = (inp[8]) ? node282 : 3'b001;
								assign node282 = (inp[2]) ? 3'b001 : 3'b101;
						assign node285 = (inp[4]) ? node291 : node286;
							assign node286 = (inp[11]) ? node288 : 3'b001;
								assign node288 = (inp[2]) ? 3'b110 : 3'b001;
							assign node291 = (inp[10]) ? node295 : node292;
								assign node292 = (inp[8]) ? 3'b110 : 3'b010;
								assign node295 = (inp[8]) ? 3'b110 : 3'b100;
				assign node298 = (inp[0]) ? node328 : node299;
					assign node299 = (inp[8]) ? node313 : node300;
						assign node300 = (inp[4]) ? node306 : node301;
							assign node301 = (inp[7]) ? node303 : 3'b010;
								assign node303 = (inp[11]) ? 3'b010 : 3'b001;
							assign node306 = (inp[10]) ? node310 : node307;
								assign node307 = (inp[11]) ? 3'b110 : 3'b000;
								assign node310 = (inp[7]) ? 3'b100 : 3'b000;
						assign node313 = (inp[4]) ? node321 : node314;
							assign node314 = (inp[7]) ? node318 : node315;
								assign node315 = (inp[10]) ? 3'b110 : 3'b000;
								assign node318 = (inp[5]) ? 3'b001 : 3'b101;
							assign node321 = (inp[1]) ? node325 : node322;
								assign node322 = (inp[2]) ? 3'b010 : 3'b110;
								assign node325 = (inp[7]) ? 3'b010 : 3'b100;
					assign node328 = (inp[4]) ? node342 : node329;
						assign node329 = (inp[5]) ? node337 : node330;
							assign node330 = (inp[7]) ? node334 : node331;
								assign node331 = (inp[8]) ? 3'b000 : 3'b100;
								assign node334 = (inp[8]) ? 3'b110 : 3'b010;
							assign node337 = (inp[7]) ? node339 : 3'b000;
								assign node339 = (inp[10]) ? 3'b000 : 3'b010;
						assign node342 = (inp[10]) ? 3'b000 : node343;
							assign node343 = (inp[5]) ? node347 : node344;
								assign node344 = (inp[2]) ? 3'b010 : 3'b000;
								assign node347 = (inp[11]) ? 3'b000 : 3'b100;

endmodule