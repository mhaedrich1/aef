module dtc_split05_bm45 (
	input  wire [16-1:0] inp,
	output wire [46-1:0] outp
);

	wire [46-1:0] node1;
	wire [46-1:0] node2;
	wire [46-1:0] node4;
	wire [46-1:0] node5;
	wire [46-1:0] node6;
	wire [46-1:0] node8;
	wire [46-1:0] node10;
	wire [46-1:0] node12;
	wire [46-1:0] node14;
	wire [46-1:0] node16;
	wire [46-1:0] node21;
	wire [46-1:0] node23;
	wire [46-1:0] node24;
	wire [46-1:0] node25;
	wire [46-1:0] node26;
	wire [46-1:0] node27;
	wire [46-1:0] node32;
	wire [46-1:0] node33;
	wire [46-1:0] node34;
	wire [46-1:0] node38;
	wire [46-1:0] node39;
	wire [46-1:0] node42;
	wire [46-1:0] node45;
	wire [46-1:0] node46;
	wire [46-1:0] node47;
	wire [46-1:0] node48;
	wire [46-1:0] node52;
	wire [46-1:0] node53;
	wire [46-1:0] node55;
	wire [46-1:0] node57;
	wire [46-1:0] node61;
	wire [46-1:0] node62;
	wire [46-1:0] node63;
	wire [46-1:0] node65;
	wire [46-1:0] node66;
	wire [46-1:0] node72;
	wire [46-1:0] node73;
	wire [46-1:0] node74;
	wire [46-1:0] node77;
	wire [46-1:0] node78;
	wire [46-1:0] node79;
	wire [46-1:0] node80;
	wire [46-1:0] node81;
	wire [46-1:0] node84;
	wire [46-1:0] node87;
	wire [46-1:0] node88;
	wire [46-1:0] node91;
	wire [46-1:0] node94;
	wire [46-1:0] node95;
	wire [46-1:0] node96;
	wire [46-1:0] node99;
	wire [46-1:0] node102;
	wire [46-1:0] node103;
	wire [46-1:0] node106;
	wire [46-1:0] node109;
	wire [46-1:0] node110;
	wire [46-1:0] node111;
	wire [46-1:0] node112;
	wire [46-1:0] node115;
	wire [46-1:0] node118;
	wire [46-1:0] node119;
	wire [46-1:0] node122;
	wire [46-1:0] node125;
	wire [46-1:0] node126;
	wire [46-1:0] node127;
	wire [46-1:0] node130;
	wire [46-1:0] node133;
	wire [46-1:0] node134;
	wire [46-1:0] node137;
	wire [46-1:0] node140;
	wire [46-1:0] node141;
	wire [46-1:0] node144;
	wire [46-1:0] node146;
	wire [46-1:0] node147;
	wire [46-1:0] node148;
	wire [46-1:0] node149;
	wire [46-1:0] node150;
	wire [46-1:0] node151;
	wire [46-1:0] node152;
	wire [46-1:0] node153;
	wire [46-1:0] node157;
	wire [46-1:0] node159;
	wire [46-1:0] node162;
	wire [46-1:0] node163;
	wire [46-1:0] node166;
	wire [46-1:0] node169;
	wire [46-1:0] node170;
	wire [46-1:0] node171;
	wire [46-1:0] node174;
	wire [46-1:0] node177;
	wire [46-1:0] node178;
	wire [46-1:0] node181;
	wire [46-1:0] node184;
	wire [46-1:0] node185;
	wire [46-1:0] node186;
	wire [46-1:0] node188;
	wire [46-1:0] node191;
	wire [46-1:0] node192;
	wire [46-1:0] node193;
	wire [46-1:0] node199;
	wire [46-1:0] node200;
	wire [46-1:0] node201;
	wire [46-1:0] node203;
	wire [46-1:0] node206;
	wire [46-1:0] node207;
	wire [46-1:0] node208;
	wire [46-1:0] node210;
	wire [46-1:0] node213;
	wire [46-1:0] node214;
	wire [46-1:0] node218;
	wire [46-1:0] node219;
	wire [46-1:0] node220;
	wire [46-1:0] node224;
	wire [46-1:0] node225;
	wire [46-1:0] node229;
	wire [46-1:0] node230;
	wire [46-1:0] node231;
	wire [46-1:0] node232;
	wire [46-1:0] node233;
	wire [46-1:0] node237;
	wire [46-1:0] node240;
	wire [46-1:0] node241;
	wire [46-1:0] node244;
	wire [46-1:0] node245;
	wire [46-1:0] node248;
	wire [46-1:0] node251;
	wire [46-1:0] node252;
	wire [46-1:0] node253;
	wire [46-1:0] node254;
	wire [46-1:0] node258;
	wire [46-1:0] node261;
	wire [46-1:0] node262;
	wire [46-1:0] node263;
	wire [46-1:0] node266;
	wire [46-1:0] node269;
	wire [46-1:0] node271;
	wire [46-1:0] node274;
	wire [46-1:0] node275;
	wire [46-1:0] node276;
	wire [46-1:0] node278;
	wire [46-1:0] node279;
	wire [46-1:0] node281;
	wire [46-1:0] node283;
	wire [46-1:0] node286;
	wire [46-1:0] node287;
	wire [46-1:0] node288;
	wire [46-1:0] node293;
	wire [46-1:0] node294;
	wire [46-1:0] node295;
	wire [46-1:0] node296;
	wire [46-1:0] node298;
	wire [46-1:0] node301;
	wire [46-1:0] node302;
	wire [46-1:0] node305;
	wire [46-1:0] node308;
	wire [46-1:0] node309;
	wire [46-1:0] node310;
	wire [46-1:0] node313;
	wire [46-1:0] node316;
	wire [46-1:0] node318;
	wire [46-1:0] node321;
	wire [46-1:0] node322;
	wire [46-1:0] node323;
	wire [46-1:0] node325;
	wire [46-1:0] node328;
	wire [46-1:0] node330;
	wire [46-1:0] node333;
	wire [46-1:0] node334;
	wire [46-1:0] node336;
	wire [46-1:0] node339;
	wire [46-1:0] node341;
	wire [46-1:0] node344;
	wire [46-1:0] node345;
	wire [46-1:0] node347;
	wire [46-1:0] node348;
	wire [46-1:0] node349;
	wire [46-1:0] node352;
	wire [46-1:0] node355;
	wire [46-1:0] node356;
	wire [46-1:0] node357;
	wire [46-1:0] node360;
	wire [46-1:0] node363;
	wire [46-1:0] node366;
	wire [46-1:0] node367;
	wire [46-1:0] node368;
	wire [46-1:0] node369;
	wire [46-1:0] node370;
	wire [46-1:0] node373;
	wire [46-1:0] node376;
	wire [46-1:0] node377;
	wire [46-1:0] node380;

	assign outp = (inp[1]) ? node72 : node1;
		assign node1 = (inp[15]) ? node21 : node2;
			assign node2 = (inp[6]) ? node4 : 46'b0000000000000000000000000000000000000000000000;
				assign node4 = (inp[9]) ? 46'b0000000000000000000000000000000000000000000000 : node5;
					assign node5 = (inp[11]) ? 46'b0000000000000000000000000000000000000000000000 : node6;
						assign node6 = (inp[5]) ? node8 : 46'b0000000000000000000000000000000000000000000000;
							assign node8 = (inp[12]) ? node10 : 46'b0000000000000000000000000000000000000000000000;
								assign node10 = (inp[7]) ? node12 : 46'b0000000000000000000000000000000000000000000000;
									assign node12 = (inp[3]) ? node14 : 46'b0000000000000000000000000000000000000000000000;
										assign node14 = (inp[13]) ? node16 : 46'b0000000000000000000000000000000000000000000000;
											assign node16 = (inp[2]) ? 46'b0000000000000000000000000000000000000100000000 : 46'b0000000000000000000000000000000000000000000000;
			assign node21 = (inp[3]) ? node23 : 46'b0000000000000000000000000000001000000000000000;
				assign node23 = (inp[9]) ? node45 : node24;
					assign node24 = (inp[11]) ? node32 : node25;
						assign node25 = (inp[2]) ? 46'b0000000000000000000000000000000000000000000000 : node26;
							assign node26 = (inp[13]) ? 46'b0000000000000000000000000000000000000000000000 : node27;
								assign node27 = (inp[0]) ? 46'b0000000000001000000000000010000000000000000000 : 46'b0000001000001000000000000000000000000000000000;
						assign node32 = (inp[13]) ? node38 : node33;
							assign node33 = (inp[2]) ? 46'b0000000000000000000000000000000000000000000000 : node34;
								assign node34 = (inp[0]) ? 46'b0000010000000000000000000010000000000000000000 : 46'b0000011000000000000000000000000000000000000000;
							assign node38 = (inp[2]) ? node42 : node39;
								assign node39 = (inp[0]) ? 46'b0000001000000000011000000100000000000000010000 : 46'b0000001000000000010000000100000000000000010010;
								assign node42 = (inp[0]) ? 46'b0000001000000000010010000000010000000010000000 : 46'b0000001000000000010010100000000000000010000000;
					assign node45 = (inp[2]) ? node61 : node46;
						assign node46 = (inp[0]) ? node52 : node47;
							assign node47 = (inp[13]) ? 46'b0000000000000000000000000000000000000000000000 : node48;
								assign node48 = (inp[11]) ? 46'b0000010100000000000000000000000000000000000000 : 46'b0000000100001000000000000000000000000000000000;
							assign node52 = (inp[11]) ? 46'b0000000000000000000000000000000000000000000000 : node53;
								assign node53 = (inp[13]) ? node55 : 46'b0010001000000000000000000000000000000000010000;
									assign node55 = (inp[12]) ? node57 : 46'b0000000000000000000000000000000000000000000000;
										assign node57 = (inp[10]) ? 46'b0000010000000000010000010000000000000000010100 : 46'b0000000000000000000000000000000000000000000000;
						assign node61 = (inp[0]) ? 46'b0000000000000000000000000000000000000000000000 : node62;
							assign node62 = (inp[11]) ? 46'b0000000000000000000000000000000000000000000000 : node63;
								assign node63 = (inp[14]) ? node65 : 46'b0000000000000000000000000000000000000000000000;
									assign node65 = (inp[12]) ? 46'b0000000000000000000000000000000000000000000000 : node66;
										assign node66 = (inp[5]) ? 46'b0000000000001000010000000000000100000010000000 : 46'b0000000000000000000000000000000000000000000000;
		assign node72 = (inp[15]) ? node140 : node73;
			assign node73 = (inp[13]) ? node77 : node74;
				assign node74 = (inp[3]) ? 46'b0000100000000000000000000000001000000000000000 : 46'b0000100000000000000000000000000000000000000000;
				assign node77 = (inp[2]) ? node109 : node78;
					assign node78 = (inp[9]) ? node94 : node79;
						assign node79 = (inp[0]) ? node87 : node80;
							assign node80 = (inp[11]) ? node84 : node81;
								assign node81 = (inp[3]) ? 46'b0000100000001000010000010100001000000000010010 : 46'b0000100000001000010000010100000000000000010010;
								assign node84 = (inp[3]) ? 46'b0000100000001000011000010100001000000000010000 : 46'b0000100000001000011000010100000000000000010000;
							assign node87 = (inp[11]) ? node91 : node88;
								assign node88 = (inp[3]) ? 46'b0000100000001000010000000100001100000000010010 : 46'b0000100000001000010000000100000100000000010010;
								assign node91 = (inp[3]) ? 46'b0000100000001000011000000100001100000000010000 : 46'b0000100000001000011000000100000100000000010000;
						assign node94 = (inp[0]) ? node102 : node95;
							assign node95 = (inp[11]) ? node99 : node96;
								assign node96 = (inp[3]) ? 46'b0000110000000000010000010100001000000000010010 : 46'b0000110000000000010000010100000000000000010010;
								assign node99 = (inp[3]) ? 46'b0000110000000000011000010100001000000000010000 : 46'b0000110000000000011000010100000000000000010000;
							assign node102 = (inp[11]) ? node106 : node103;
								assign node103 = (inp[3]) ? 46'b0000110000000000010000000100001100000000010010 : 46'b0000110000000000010000000100000100000000010010;
								assign node106 = (inp[3]) ? 46'b0000110000000000011000000100001100000000010000 : 46'b0000110000000000011000000100000100000000010000;
					assign node109 = (inp[0]) ? node125 : node110;
						assign node110 = (inp[9]) ? node118 : node111;
							assign node111 = (inp[11]) ? node115 : node112;
								assign node112 = (inp[3]) ? 46'b0000100000001000010010110000001000000010000000 : 46'b0000100000001000010010110000000000000010000000;
								assign node115 = (inp[3]) ? 46'b0000100000001000010010010000011000000010000000 : 46'b0000100000001000010010010000010000000010000000;
							assign node118 = (inp[11]) ? node122 : node119;
								assign node119 = (inp[3]) ? 46'b0000110000000000010010110000001000000010000000 : 46'b0000110000000000010010110000000000000010000000;
								assign node122 = (inp[3]) ? 46'b0000110000000000010010010000011000000010000000 : 46'b0000110000000000010010010000010000000010000000;
						assign node125 = (inp[9]) ? node133 : node126;
							assign node126 = (inp[11]) ? node130 : node127;
								assign node127 = (inp[3]) ? 46'b0000100000001000010010100000001100000010000000 : 46'b0000100000001000010010100000000100000010000000;
								assign node130 = (inp[3]) ? 46'b0000100000001000010010000000011100000010000000 : 46'b0000100000001000010010000000010100000010000000;
							assign node133 = (inp[11]) ? node137 : node134;
								assign node134 = (inp[3]) ? 46'b0000110000000000010010100000001100000010000000 : 46'b0000110000000000010010100000000100000010000000;
								assign node137 = (inp[3]) ? 46'b0000110000000000010010000000011100000010000000 : 46'b0000110000000000010010000000010100000010000000;
			assign node140 = (inp[13]) ? node144 : node141;
				assign node141 = (inp[3]) ? 46'b0000000000000000000000000000000000000000001000 : 46'b0000000000000000000000000000001000000000001000;
				assign node144 = (inp[3]) ? node146 : 46'b0000000000000000000000000000001000000000000000;
					assign node146 = (inp[2]) ? node274 : node147;
						assign node147 = (inp[11]) ? node199 : node148;
							assign node148 = (inp[9]) ? node184 : node149;
								assign node149 = (inp[6]) ? node169 : node150;
									assign node150 = (inp[5]) ? node162 : node151;
										assign node151 = (inp[8]) ? node157 : node152;
											assign node152 = (inp[0]) ? 46'b0011000000000100000000010000100000110000010000 : node153;
												assign node153 = (inp[14]) ? 46'b0011000000000000001000010001100000110001010010 : 46'b0011000000000100001000010001000010110001010000;
											assign node157 = (inp[12]) ? node159 : 46'b0011000000000010000000010001100010110000010010;
												assign node159 = (inp[4]) ? 46'b0011000000000010000000010000000000110001010000 : 46'b0011000000000010000000010001000000110001010010;
										assign node162 = (inp[12]) ? node166 : node163;
											assign node163 = (inp[14]) ? 46'b0010000000000010000000010001000010110001010010 : 46'b0010000000000100000000010001000010110001010010;
											assign node166 = (inp[10]) ? 46'b0010000000000000000000010001000000110000010010 : 46'b0010000000000100000000010001000000110001010010;
									assign node169 = (inp[5]) ? node177 : node170;
										assign node170 = (inp[12]) ? node174 : node171;
											assign node171 = (inp[4]) ? 46'b0011000000000110000000010000000010010001010000 : 46'b0011000000000100000000010001000010010001010010;
											assign node174 = (inp[4]) ? 46'b0011000000000010001000010001000000010001010000 : 46'b0011000000000110000000010000100000010001010000;
										assign node177 = (inp[0]) ? node181 : node178;
											assign node178 = (inp[12]) ? 46'b0010000000000010001000010001100000010001010000 : 46'b0010000000000110000000010000100010010001010000;
											assign node181 = (inp[8]) ? 46'b0010000000000010000000010001100010010000010010 : 46'b0010000000000100001000010001100010010000010000;
								assign node184 = (inp[0]) ? 46'b0000000000000000000000000000000000000000000000 : node185;
									assign node185 = (inp[6]) ? node191 : node186;
										assign node186 = (inp[7]) ? node188 : 46'b0000000000000000000000000000000000000000000000;
											assign node188 = (inp[10]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0001000000000100001000001001000000100000000000;
										assign node191 = (inp[4]) ? 46'b0000000000000000000000000000000000000000000000 : node192;
											assign node192 = (inp[14]) ? 46'b0000000000000010000000001001100010000000000010 : node193;
												assign node193 = (inp[10]) ? 46'b0001000000000100000000001001000010000000000010 : 46'b0000000000000100000000001001100010000000000010;
							assign node199 = (inp[9]) ? node229 : node200;
								assign node200 = (inp[0]) ? node206 : node201;
									assign node201 = (inp[7]) ? node203 : 46'b0000000000000000000000000000000000000000000000;
										assign node203 = (inp[5]) ? 46'b0000000000000000001001000001000010000000000000 : 46'b0000000000000000000000000000000000000000000000;
									assign node206 = (inp[6]) ? node218 : node207;
										assign node207 = (inp[12]) ? node213 : node208;
											assign node208 = (inp[4]) ? node210 : 46'b0100000000000100000000000000100010100000000000;
												assign node210 = (inp[7]) ? 46'b0100000000000100001000000001000010100000000000 : 46'b0100000000000100001000000001100010100000000000;
											assign node213 = (inp[7]) ? 46'b0100000000000110000000000000000000100000000000 : node214;
												assign node214 = (inp[4]) ? 46'b0100000000000000001000000001100000100000000000 : 46'b0100000000000110000000000000100000100000000000;
										assign node218 = (inp[10]) ? node224 : node219;
											assign node219 = (inp[14]) ? 46'b0101000000000110000000000000100010000000000000 : node220;
												assign node220 = (inp[4]) ? 46'b0101000000000100001000000001000010000000000000 : 46'b0101000000000100000000000000000000000000000000;
											assign node224 = (inp[12]) ? 46'b0101000000000000001000000001000000000000000010 : node225;
												assign node225 = (inp[8]) ? 46'b0101000000000010000000000000000010000000000000 : 46'b0101000000000010001000000001000010000000000000;
								assign node229 = (inp[0]) ? node251 : node230;
									assign node230 = (inp[4]) ? node240 : node231;
										assign node231 = (inp[6]) ? node237 : node232;
											assign node232 = (inp[5]) ? 46'b1000000000000100000000000001000010100000000010 : node233;
												assign node233 = (inp[12]) ? 46'b1001000000000110000000000000000000100000000000 : 46'b1001000000000110000000000000000010100000000000;
											assign node237 = (inp[8]) ? 46'b1001000000000100000000000001000010000000000010 : 46'b1001000000000000001000000001000000000000000010;
										assign node240 = (inp[6]) ? node244 : node241;
											assign node241 = (inp[8]) ? 46'b1000000000000000001000000001100000100000000010 : 46'b1001000000000100001000000001100000100000000000;
											assign node244 = (inp[14]) ? node248 : node245;
												assign node245 = (inp[5]) ? 46'b1000000000000100001000000001000000000000000000 : 46'b1001000000000100001000000001000010000000000000;
												assign node248 = (inp[12]) ? 46'b1000000000000010001000000001000000000000000000 : 46'b1000000000000010001000000001000010000000000000;
									assign node251 = (inp[12]) ? node261 : node252;
										assign node252 = (inp[6]) ? node258 : node253;
											assign node253 = (inp[8]) ? 46'b0001000000000010000000000001100010101000000010 : node254;
												assign node254 = (inp[7]) ? 46'b0001000000000100000000000001000010101000000010 : 46'b0001000000000100000000000001100010101000000010;
											assign node258 = (inp[10]) ? 46'b0000000000000000000000000001100010001000000010 : 46'b0000000000000100000000000001100010001000000010;
										assign node261 = (inp[7]) ? node269 : node262;
											assign node262 = (inp[8]) ? node266 : node263;
												assign node263 = (inp[4]) ? 46'b0000000000000100001000000001100000101000000000 : 46'b0000000000000100001000000001100000001000000000;
												assign node266 = (inp[10]) ? 46'b0001000000000000000000000001100000001000000010 : 46'b0000000000000100000000000001100000001000000010;
											assign node269 = (inp[5]) ? node271 : 46'b0001000000000000001000000001000000101000000000;
												assign node271 = (inp[4]) ? 46'b0000000000000110000000000000000000101000000000 : 46'b0000000000000000000000000000000000101000000000;
						assign node274 = (inp[11]) ? node344 : node275;
							assign node275 = (inp[9]) ? node293 : node276;
								assign node276 = (inp[7]) ? node278 : 46'b0000000000000000000000000000000000000000000000;
									assign node278 = (inp[5]) ? node286 : node279;
										assign node279 = (inp[0]) ? node281 : 46'b0000000000000000000000000000000000000000000000;
											assign node281 = (inp[12]) ? node283 : 46'b0000000000000000000000000000000000000000000000;
												assign node283 = (inp[4]) ? 46'b0001000000000011001000000001000000000000100000 : 46'b0001000000000001001000000001000000000000100010;
										assign node286 = (inp[0]) ? 46'b0000000000000000000000000000000000000000000000 : node287;
											assign node287 = (inp[8]) ? 46'b0000000000100110000001000000000010100000000000 : node288;
												assign node288 = (inp[12]) ? 46'b0000000000100100001001000001000000000000000000 : 46'b0000000000100100001001000001000010100000000000;
								assign node293 = (inp[5]) ? node321 : node294;
									assign node294 = (inp[0]) ? node308 : node295;
										assign node295 = (inp[6]) ? node301 : node296;
											assign node296 = (inp[4]) ? node298 : 46'b0001000000100010000000000001000000100000100010;
												assign node298 = (inp[10]) ? 46'b0001000000100010001000000001000010100000100000 : 46'b0001000000100010001000000001000000100000100000;
											assign node301 = (inp[10]) ? node305 : node302;
												assign node302 = (inp[4]) ? 46'b0001000000100000001000000001100000000000100000 : 46'b0001000000100100001000000001100000000000100000;
												assign node305 = (inp[7]) ? 46'b0001000000100110000000000000000000000000100000 : 46'b0001000000100110000000000000100010000000100000;
										assign node308 = (inp[12]) ? node316 : node309;
											assign node309 = (inp[7]) ? node313 : node310;
												assign node310 = (inp[6]) ? 46'b0001000000000000001000000001100010000000100010 : 46'b0001000000000100001000000001100010100000100000;
												assign node313 = (inp[10]) ? 46'b0001000000000000001000000001000010100000100010 : 46'b0001000000000100000000000001000010000000100000;
											assign node316 = (inp[10]) ? node318 : 46'b0001000000000000001000000001000000100000100000;
												assign node318 = (inp[6]) ? 46'b0001000000000010000000000001000000000000100010 : 46'b0001000000000000000000000001000000100000100010;
									assign node321 = (inp[0]) ? node333 : node322;
										assign node322 = (inp[12]) ? node328 : node323;
											assign node323 = (inp[8]) ? node325 : 46'b0000000000100000001000000001100010000000100010;
												assign node325 = (inp[4]) ? 46'b0000000000100010000000000001000010100000100010 : 46'b0000000000100010000000000001000010000000100010;
											assign node328 = (inp[8]) ? node330 : 46'b0000000000100110000000000000100000000000100000;
												assign node330 = (inp[4]) ? 46'b0000000000100000001000000001100000100000100010 : 46'b0000000000100110000000000000000000100000100000;
										assign node333 = (inp[7]) ? node339 : node334;
											assign node334 = (inp[12]) ? node336 : 46'b0000000000000110000000000000100010000000100000;
												assign node336 = (inp[10]) ? 46'b0000000000000010000000000000100000000000100000 : 46'b0000000000000000001000000001100000000000100010;
											assign node339 = (inp[8]) ? node341 : 46'b0000000000000100001000000001000000100000100000;
												assign node341 = (inp[4]) ? 46'b0000000000000010001000000001000000000000100000 : 46'b0000000000000000000000000001000000000000100010;
							assign node344 = (inp[7]) ? node366 : node345;
								assign node345 = (inp[5]) ? node347 : 46'b0000000000000000000000000000000000000000000000;
									assign node347 = (inp[12]) ? node355 : node348;
										assign node348 = (inp[9]) ? node352 : node349;
											assign node349 = (inp[6]) ? 46'b0000000000100010000000000000100010000000100000 : 46'b0000000000000000000000000000000000000000000000;
											assign node352 = (inp[8]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0000000010000000000000000001100010100001000010;
										assign node355 = (inp[9]) ? node363 : node356;
											assign node356 = (inp[0]) ? node360 : node357;
												assign node357 = (inp[10]) ? 46'b0000000000100000001000000001100000100000100000 : 46'b0000000000000000000000000000000000000000000000;
												assign node360 = (inp[6]) ? 46'b0000000010000000000000000001100000000000000010 : 46'b0000000010000000000000000001100000100000000010;
											assign node363 = (inp[0]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0000000010000000000000000001100000000001000010;
								assign node366 = (inp[5]) ? 46'b0000000000000000000000000000000000000000000000 : node367;
									assign node367 = (inp[10]) ? 46'b0001000000100000001000000001000000100000100000 : node368;
										assign node368 = (inp[12]) ? node376 : node369;
											assign node369 = (inp[6]) ? node373 : node370;
												assign node370 = (inp[0]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0001000010000100000000000000000010100001000000;
												assign node373 = (inp[9]) ? 46'b0001000010000100000000000000000010000001000000 : 46'b0001000000100010000000000000000010000000100000;
											assign node376 = (inp[0]) ? node380 : node377;
												assign node377 = (inp[9]) ? 46'b0001000010000100000000000000000000000001000000 : 46'b0000000000000000000000000000000000000000000000;
												assign node380 = (inp[9]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0001000010000100000000000000000000100000000000;

endmodule