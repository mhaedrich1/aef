module dtc_split125_bm83 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node8;
	wire [3-1:0] node11;
	wire [3-1:0] node12;
	wire [3-1:0] node15;
	wire [3-1:0] node18;
	wire [3-1:0] node19;
	wire [3-1:0] node20;
	wire [3-1:0] node23;
	wire [3-1:0] node26;
	wire [3-1:0] node27;
	wire [3-1:0] node30;
	wire [3-1:0] node33;
	wire [3-1:0] node34;
	wire [3-1:0] node35;
	wire [3-1:0] node36;
	wire [3-1:0] node39;
	wire [3-1:0] node42;
	wire [3-1:0] node43;
	wire [3-1:0] node46;
	wire [3-1:0] node49;
	wire [3-1:0] node50;
	wire [3-1:0] node51;
	wire [3-1:0] node54;
	wire [3-1:0] node57;
	wire [3-1:0] node58;
	wire [3-1:0] node61;
	wire [3-1:0] node64;
	wire [3-1:0] node65;
	wire [3-1:0] node66;
	wire [3-1:0] node67;
	wire [3-1:0] node68;
	wire [3-1:0] node71;
	wire [3-1:0] node74;
	wire [3-1:0] node75;
	wire [3-1:0] node78;
	wire [3-1:0] node81;
	wire [3-1:0] node82;
	wire [3-1:0] node83;
	wire [3-1:0] node86;
	wire [3-1:0] node89;
	wire [3-1:0] node90;
	wire [3-1:0] node93;
	wire [3-1:0] node96;
	wire [3-1:0] node97;
	wire [3-1:0] node98;
	wire [3-1:0] node99;
	wire [3-1:0] node102;
	wire [3-1:0] node105;
	wire [3-1:0] node106;
	wire [3-1:0] node109;
	wire [3-1:0] node112;
	wire [3-1:0] node114;
	wire [3-1:0] node115;

	assign outp = (inp[3]) ? node64 : node1;
		assign node1 = (inp[4]) ? node33 : node2;
			assign node2 = (inp[9]) ? node18 : node3;
				assign node3 = (inp[7]) ? node11 : node4;
					assign node4 = (inp[1]) ? node8 : node5;
						assign node5 = (inp[5]) ? 3'b101 : 3'b111;
						assign node8 = (inp[11]) ? 3'b111 : 3'b011;
					assign node11 = (inp[5]) ? node15 : node12;
						assign node12 = (inp[11]) ? 3'b111 : 3'b111;
						assign node15 = (inp[1]) ? 3'b111 : 3'b011;
				assign node18 = (inp[0]) ? node26 : node19;
					assign node19 = (inp[6]) ? node23 : node20;
						assign node20 = (inp[10]) ? 3'b010 : 3'b001;
						assign node23 = (inp[10]) ? 3'b101 : 3'b001;
					assign node26 = (inp[6]) ? node30 : node27;
						assign node27 = (inp[7]) ? 3'b001 : 3'b101;
						assign node30 = (inp[1]) ? 3'b111 : 3'b111;
			assign node33 = (inp[0]) ? node49 : node34;
				assign node34 = (inp[8]) ? node42 : node35;
					assign node35 = (inp[11]) ? node39 : node36;
						assign node36 = (inp[7]) ? 3'b001 : 3'b100;
						assign node39 = (inp[5]) ? 3'b000 : 3'b010;
					assign node42 = (inp[5]) ? node46 : node43;
						assign node43 = (inp[2]) ? 3'b100 : 3'b101;
						assign node46 = (inp[7]) ? 3'b110 : 3'b000;
				assign node49 = (inp[6]) ? node57 : node50;
					assign node50 = (inp[5]) ? node54 : node51;
						assign node51 = (inp[8]) ? 3'b111 : 3'b001;
						assign node54 = (inp[7]) ? 3'b101 : 3'b100;
					assign node57 = (inp[7]) ? node61 : node58;
						assign node58 = (inp[1]) ? 3'b101 : 3'b011;
						assign node61 = (inp[5]) ? 3'b001 : 3'b011;
		assign node64 = (inp[9]) ? node96 : node65;
			assign node65 = (inp[4]) ? node81 : node66;
				assign node66 = (inp[6]) ? node74 : node67;
					assign node67 = (inp[11]) ? node71 : node68;
						assign node68 = (inp[0]) ? 3'b110 : 3'b000;
						assign node71 = (inp[1]) ? 3'b000 : 3'b100;
					assign node74 = (inp[0]) ? node78 : node75;
						assign node75 = (inp[2]) ? 3'b000 : 3'b110;
						assign node78 = (inp[7]) ? 3'b001 : 3'b100;
				assign node81 = (inp[6]) ? node89 : node82;
					assign node82 = (inp[7]) ? node86 : node83;
						assign node83 = (inp[0]) ? 3'b000 : 3'b000;
						assign node86 = (inp[1]) ? 3'b100 : 3'b000;
					assign node89 = (inp[10]) ? node93 : node90;
						assign node90 = (inp[8]) ? 3'b110 : 3'b010;
						assign node93 = (inp[0]) ? 3'b010 : 3'b000;
			assign node96 = (inp[4]) ? node112 : node97;
				assign node97 = (inp[0]) ? node105 : node98;
					assign node98 = (inp[10]) ? node102 : node99;
						assign node99 = (inp[2]) ? 3'b010 : 3'b000;
						assign node102 = (inp[6]) ? 3'b000 : 3'b000;
					assign node105 = (inp[6]) ? node109 : node106;
						assign node106 = (inp[10]) ? 3'b000 : 3'b100;
						assign node109 = (inp[1]) ? 3'b010 : 3'b010;
				assign node112 = (inp[7]) ? node114 : 3'b000;
					assign node114 = (inp[10]) ? 3'b000 : node115;
						assign node115 = (inp[6]) ? 3'b100 : 3'b000;

endmodule