module dtc_split75_bm76 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node6;
	wire [3-1:0] node8;
	wire [3-1:0] node10;
	wire [3-1:0] node11;
	wire [3-1:0] node13;
	wire [3-1:0] node17;
	wire [3-1:0] node18;
	wire [3-1:0] node19;
	wire [3-1:0] node21;
	wire [3-1:0] node23;
	wire [3-1:0] node24;
	wire [3-1:0] node26;
	wire [3-1:0] node28;
	wire [3-1:0] node31;
	wire [3-1:0] node32;
	wire [3-1:0] node36;
	wire [3-1:0] node37;
	wire [3-1:0] node39;
	wire [3-1:0] node40;
	wire [3-1:0] node42;
	wire [3-1:0] node43;
	wire [3-1:0] node47;
	wire [3-1:0] node48;
	wire [3-1:0] node49;
	wire [3-1:0] node55;
	wire [3-1:0] node56;
	wire [3-1:0] node57;
	wire [3-1:0] node58;
	wire [3-1:0] node60;
	wire [3-1:0] node64;
	wire [3-1:0] node66;
	wire [3-1:0] node67;
	wire [3-1:0] node69;
	wire [3-1:0] node70;
	wire [3-1:0] node75;
	wire [3-1:0] node76;
	wire [3-1:0] node78;
	wire [3-1:0] node79;
	wire [3-1:0] node83;
	wire [3-1:0] node85;
	wire [3-1:0] node87;
	wire [3-1:0] node89;
	wire [3-1:0] node92;
	wire [3-1:0] node93;
	wire [3-1:0] node94;
	wire [3-1:0] node95;
	wire [3-1:0] node98;
	wire [3-1:0] node100;
	wire [3-1:0] node101;
	wire [3-1:0] node102;
	wire [3-1:0] node104;
	wire [3-1:0] node106;
	wire [3-1:0] node109;
	wire [3-1:0] node110;
	wire [3-1:0] node112;
	wire [3-1:0] node117;
	wire [3-1:0] node118;
	wire [3-1:0] node119;
	wire [3-1:0] node121;
	wire [3-1:0] node123;
	wire [3-1:0] node127;
	wire [3-1:0] node129;
	wire [3-1:0] node130;
	wire [3-1:0] node131;
	wire [3-1:0] node133;
	wire [3-1:0] node136;
	wire [3-1:0] node137;
	wire [3-1:0] node142;
	wire [3-1:0] node143;
	wire [3-1:0] node144;
	wire [3-1:0] node145;
	wire [3-1:0] node146;
	wire [3-1:0] node147;
	wire [3-1:0] node149;
	wire [3-1:0] node152;
	wire [3-1:0] node153;
	wire [3-1:0] node158;
	wire [3-1:0] node160;
	wire [3-1:0] node161;
	wire [3-1:0] node165;
	wire [3-1:0] node166;
	wire [3-1:0] node167;
	wire [3-1:0] node169;
	wire [3-1:0] node171;
	wire [3-1:0] node174;
	wire [3-1:0] node175;
	wire [3-1:0] node176;
	wire [3-1:0] node181;
	wire [3-1:0] node183;
	wire [3-1:0] node184;
	wire [3-1:0] node188;
	wire [3-1:0] node189;
	wire [3-1:0] node190;
	wire [3-1:0] node191;
	wire [3-1:0] node192;
	wire [3-1:0] node197;
	wire [3-1:0] node199;
	wire [3-1:0] node200;
	wire [3-1:0] node201;
	wire [3-1:0] node203;
	wire [3-1:0] node208;
	wire [3-1:0] node209;
	wire [3-1:0] node210;
	wire [3-1:0] node212;
	wire [3-1:0] node214;
	wire [3-1:0] node217;
	wire [3-1:0] node218;
	wire [3-1:0] node219;
	wire [3-1:0] node224;
	wire [3-1:0] node226;
	wire [3-1:0] node228;
	wire [3-1:0] node231;
	wire [3-1:0] node232;
	wire [3-1:0] node233;
	wire [3-1:0] node234;
	wire [3-1:0] node235;
	wire [3-1:0] node236;
	wire [3-1:0] node238;
	wire [3-1:0] node240;
	wire [3-1:0] node242;
	wire [3-1:0] node245;
	wire [3-1:0] node246;
	wire [3-1:0] node247;
	wire [3-1:0] node252;
	wire [3-1:0] node253;
	wire [3-1:0] node255;
	wire [3-1:0] node256;
	wire [3-1:0] node260;
	wire [3-1:0] node261;
	wire [3-1:0] node263;
	wire [3-1:0] node267;
	wire [3-1:0] node268;
	wire [3-1:0] node269;
	wire [3-1:0] node271;
	wire [3-1:0] node273;
	wire [3-1:0] node276;
	wire [3-1:0] node277;
	wire [3-1:0] node278;
	wire [3-1:0] node279;
	wire [3-1:0] node285;
	wire [3-1:0] node287;
	wire [3-1:0] node288;
	wire [3-1:0] node289;
	wire [3-1:0] node291;
	wire [3-1:0] node294;
	wire [3-1:0] node295;
	wire [3-1:0] node300;
	wire [3-1:0] node301;
	wire [3-1:0] node302;
	wire [3-1:0] node303;
	wire [3-1:0] node304;
	wire [3-1:0] node305;
	wire [3-1:0] node307;
	wire [3-1:0] node310;
	wire [3-1:0] node311;
	wire [3-1:0] node316;
	wire [3-1:0] node318;
	wire [3-1:0] node319;
	wire [3-1:0] node321;
	wire [3-1:0] node324;
	wire [3-1:0] node325;
	wire [3-1:0] node326;
	wire [3-1:0] node331;
	wire [3-1:0] node332;
	wire [3-1:0] node334;
	wire [3-1:0] node335;
	wire [3-1:0] node339;
	wire [3-1:0] node341;
	wire [3-1:0] node343;
	wire [3-1:0] node345;
	wire [3-1:0] node346;
	wire [3-1:0] node350;
	wire [3-1:0] node351;
	wire [3-1:0] node352;
	wire [3-1:0] node353;
	wire [3-1:0] node354;
	wire [3-1:0] node356;
	wire [3-1:0] node359;
	wire [3-1:0] node360;
	wire [3-1:0] node365;
	wire [3-1:0] node366;
	wire [3-1:0] node367;
	wire [3-1:0] node369;
	wire [3-1:0] node373;
	wire [3-1:0] node374;
	wire [3-1:0] node376;
	wire [3-1:0] node380;
	wire [3-1:0] node381;
	wire [3-1:0] node383;
	wire [3-1:0] node384;
	wire [3-1:0] node388;
	wire [3-1:0] node390;
	wire [3-1:0] node392;
	wire [3-1:0] node393;
	wire [3-1:0] node395;
	wire [3-1:0] node399;
	wire [3-1:0] node400;
	wire [3-1:0] node401;
	wire [3-1:0] node402;
	wire [3-1:0] node403;
	wire [3-1:0] node405;
	wire [3-1:0] node407;
	wire [3-1:0] node411;
	wire [3-1:0] node413;
	wire [3-1:0] node414;
	wire [3-1:0] node415;
	wire [3-1:0] node417;
	wire [3-1:0] node418;
	wire [3-1:0] node422;
	wire [3-1:0] node423;
	wire [3-1:0] node424;
	wire [3-1:0] node430;
	wire [3-1:0] node431;
	wire [3-1:0] node432;
	wire [3-1:0] node434;
	wire [3-1:0] node438;
	wire [3-1:0] node440;
	wire [3-1:0] node441;
	wire [3-1:0] node442;
	wire [3-1:0] node447;
	wire [3-1:0] node448;
	wire [3-1:0] node449;
	wire [3-1:0] node450;
	wire [3-1:0] node451;
	wire [3-1:0] node452;
	wire [3-1:0] node457;
	wire [3-1:0] node458;
	wire [3-1:0] node460;
	wire [3-1:0] node462;
	wire [3-1:0] node466;
	wire [3-1:0] node467;
	wire [3-1:0] node468;
	wire [3-1:0] node470;
	wire [3-1:0] node472;
	wire [3-1:0] node475;
	wire [3-1:0] node476;
	wire [3-1:0] node480;
	wire [3-1:0] node482;
	wire [3-1:0] node484;
	wire [3-1:0] node487;
	wire [3-1:0] node488;
	wire [3-1:0] node489;
	wire [3-1:0] node490;
	wire [3-1:0] node491;
	wire [3-1:0] node496;
	wire [3-1:0] node497;
	wire [3-1:0] node499;
	wire [3-1:0] node501;
	wire [3-1:0] node504;
	wire [3-1:0] node505;
	wire [3-1:0] node506;
	wire [3-1:0] node511;
	wire [3-1:0] node512;
	wire [3-1:0] node513;
	wire [3-1:0] node515;
	wire [3-1:0] node520;
	wire [3-1:0] node521;
	wire [3-1:0] node522;
	wire [3-1:0] node523;
	wire [3-1:0] node524;
	wire [3-1:0] node525;
	wire [3-1:0] node526;
	wire [3-1:0] node528;
	wire [3-1:0] node530;
	wire [3-1:0] node531;
	wire [3-1:0] node536;
	wire [3-1:0] node538;
	wire [3-1:0] node539;
	wire [3-1:0] node540;
	wire [3-1:0] node545;
	wire [3-1:0] node546;
	wire [3-1:0] node547;
	wire [3-1:0] node549;
	wire [3-1:0] node550;
	wire [3-1:0] node555;
	wire [3-1:0] node557;
	wire [3-1:0] node558;
	wire [3-1:0] node559;
	wire [3-1:0] node564;
	wire [3-1:0] node565;
	wire [3-1:0] node566;
	wire [3-1:0] node567;
	wire [3-1:0] node568;
	wire [3-1:0] node569;
	wire [3-1:0] node574;
	wire [3-1:0] node575;
	wire [3-1:0] node577;
	wire [3-1:0] node579;
	wire [3-1:0] node582;
	wire [3-1:0] node583;
	wire [3-1:0] node584;
	wire [3-1:0] node589;
	wire [3-1:0] node590;
	wire [3-1:0] node591;
	wire [3-1:0] node593;
	wire [3-1:0] node597;
	wire [3-1:0] node599;
	wire [3-1:0] node600;
	wire [3-1:0] node602;
	wire [3-1:0] node605;
	wire [3-1:0] node606;
	wire [3-1:0] node610;
	wire [3-1:0] node611;
	wire [3-1:0] node612;
	wire [3-1:0] node615;
	wire [3-1:0] node616;
	wire [3-1:0] node618;
	wire [3-1:0] node620;
	wire [3-1:0] node624;
	wire [3-1:0] node625;
	wire [3-1:0] node626;
	wire [3-1:0] node628;
	wire [3-1:0] node632;
	wire [3-1:0] node634;
	wire [3-1:0] node636;
	wire [3-1:0] node637;
	wire [3-1:0] node641;
	wire [3-1:0] node642;
	wire [3-1:0] node643;
	wire [3-1:0] node644;
	wire [3-1:0] node645;
	wire [3-1:0] node647;
	wire [3-1:0] node651;
	wire [3-1:0] node652;
	wire [3-1:0] node654;
	wire [3-1:0] node656;
	wire [3-1:0] node658;
	wire [3-1:0] node660;
	wire [3-1:0] node663;
	wire [3-1:0] node664;
	wire [3-1:0] node665;
	wire [3-1:0] node666;
	wire [3-1:0] node672;
	wire [3-1:0] node673;
	wire [3-1:0] node674;
	wire [3-1:0] node677;
	wire [3-1:0] node679;
	wire [3-1:0] node681;
	wire [3-1:0] node684;
	wire [3-1:0] node685;
	wire [3-1:0] node687;
	wire [3-1:0] node689;
	wire [3-1:0] node691;
	wire [3-1:0] node694;
	wire [3-1:0] node695;
	wire [3-1:0] node696;
	wire [3-1:0] node697;
	wire [3-1:0] node703;
	wire [3-1:0] node704;
	wire [3-1:0] node705;
	wire [3-1:0] node706;
	wire [3-1:0] node707;
	wire [3-1:0] node708;
	wire [3-1:0] node713;
	wire [3-1:0] node714;
	wire [3-1:0] node716;
	wire [3-1:0] node720;
	wire [3-1:0] node721;
	wire [3-1:0] node722;
	wire [3-1:0] node728;
	wire [3-1:0] node729;
	wire [3-1:0] node730;
	wire [3-1:0] node731;
	wire [3-1:0] node732;
	wire [3-1:0] node733;
	wire [3-1:0] node735;
	wire [3-1:0] node739;
	wire [3-1:0] node740;
	wire [3-1:0] node742;
	wire [3-1:0] node744;
	wire [3-1:0] node746;
	wire [3-1:0] node748;
	wire [3-1:0] node751;
	wire [3-1:0] node752;
	wire [3-1:0] node753;
	wire [3-1:0] node754;
	wire [3-1:0] node760;
	wire [3-1:0] node761;
	wire [3-1:0] node762;
	wire [3-1:0] node764;

	assign outp = (inp[9]) ? node520 : node1;
		assign node1 = (inp[6]) ? node231 : node2;
			assign node2 = (inp[10]) ? node92 : node3;
				assign node3 = (inp[7]) ? node17 : node4;
					assign node4 = (inp[11]) ? node6 : 3'b111;
						assign node6 = (inp[8]) ? node8 : 3'b111;
							assign node8 = (inp[3]) ? node10 : 3'b111;
								assign node10 = (inp[4]) ? 3'b011 : node11;
									assign node11 = (inp[5]) ? node13 : 3'b111;
										assign node13 = (inp[0]) ? 3'b011 : 3'b111;
					assign node17 = (inp[11]) ? node55 : node18;
						assign node18 = (inp[8]) ? node36 : node19;
							assign node19 = (inp[4]) ? node21 : 3'b111;
								assign node21 = (inp[3]) ? node23 : 3'b111;
									assign node23 = (inp[5]) ? node31 : node24;
										assign node24 = (inp[0]) ? node26 : 3'b111;
											assign node26 = (inp[1]) ? node28 : 3'b111;
												assign node28 = (inp[2]) ? 3'b011 : 3'b111;
										assign node31 = (inp[0]) ? 3'b011 : node32;
											assign node32 = (inp[1]) ? 3'b011 : 3'b111;
							assign node36 = (inp[3]) ? 3'b011 : node37;
								assign node37 = (inp[4]) ? node39 : 3'b111;
									assign node39 = (inp[0]) ? node47 : node40;
										assign node40 = (inp[5]) ? node42 : 3'b111;
											assign node42 = (inp[1]) ? 3'b011 : node43;
												assign node43 = (inp[2]) ? 3'b011 : 3'b111;
										assign node47 = (inp[1]) ? 3'b011 : node48;
											assign node48 = (inp[2]) ? 3'b011 : node49;
												assign node49 = (inp[5]) ? 3'b011 : 3'b111;
						assign node55 = (inp[8]) ? node75 : node56;
							assign node56 = (inp[4]) ? node64 : node57;
								assign node57 = (inp[3]) ? 3'b011 : node58;
									assign node58 = (inp[5]) ? node60 : 3'b111;
										assign node60 = (inp[0]) ? 3'b011 : 3'b111;
								assign node64 = (inp[3]) ? node66 : 3'b011;
									assign node66 = (inp[5]) ? 3'b101 : node67;
										assign node67 = (inp[0]) ? node69 : 3'b011;
											assign node69 = (inp[2]) ? 3'b101 : node70;
												assign node70 = (inp[1]) ? 3'b101 : 3'b011;
							assign node75 = (inp[3]) ? node83 : node76;
								assign node76 = (inp[4]) ? node78 : 3'b011;
									assign node78 = (inp[5]) ? 3'b101 : node79;
										assign node79 = (inp[0]) ? 3'b101 : 3'b011;
								assign node83 = (inp[5]) ? node85 : 3'b101;
									assign node85 = (inp[2]) ? node87 : 3'b101;
										assign node87 = (inp[1]) ? node89 : 3'b101;
											assign node89 = (inp[4]) ? 3'b001 : 3'b101;
				assign node92 = (inp[7]) ? node142 : node93;
					assign node93 = (inp[11]) ? node117 : node94;
						assign node94 = (inp[3]) ? node98 : node95;
							assign node95 = (inp[8]) ? 3'b011 : 3'b111;
							assign node98 = (inp[8]) ? node100 : 3'b011;
								assign node100 = (inp[4]) ? 3'b101 : node101;
									assign node101 = (inp[0]) ? node109 : node102;
										assign node102 = (inp[5]) ? node104 : 3'b011;
											assign node104 = (inp[2]) ? node106 : 3'b011;
												assign node106 = (inp[1]) ? 3'b101 : 3'b011;
										assign node109 = (inp[5]) ? 3'b101 : node110;
											assign node110 = (inp[1]) ? node112 : 3'b011;
												assign node112 = (inp[2]) ? 3'b101 : 3'b011;
						assign node117 = (inp[8]) ? node127 : node118;
							assign node118 = (inp[3]) ? 3'b101 : node119;
								assign node119 = (inp[0]) ? node121 : 3'b011;
									assign node121 = (inp[4]) ? node123 : 3'b011;
										assign node123 = (inp[5]) ? 3'b101 : 3'b011;
							assign node127 = (inp[3]) ? node129 : 3'b101;
								assign node129 = (inp[4]) ? 3'b001 : node130;
									assign node130 = (inp[5]) ? node136 : node131;
										assign node131 = (inp[1]) ? node133 : 3'b101;
											assign node133 = (inp[2]) ? 3'b101 : 3'b001;
										assign node136 = (inp[0]) ? 3'b001 : node137;
											assign node137 = (inp[1]) ? 3'b001 : 3'b101;
					assign node142 = (inp[11]) ? node188 : node143;
						assign node143 = (inp[8]) ? node165 : node144;
							assign node144 = (inp[4]) ? node158 : node145;
								assign node145 = (inp[3]) ? 3'b101 : node146;
									assign node146 = (inp[0]) ? node152 : node147;
										assign node147 = (inp[1]) ? node149 : 3'b011;
											assign node149 = (inp[5]) ? 3'b111 : 3'b011;
										assign node152 = (inp[5]) ? 3'b101 : node153;
											assign node153 = (inp[1]) ? 3'b111 : 3'b011;
								assign node158 = (inp[3]) ? node160 : 3'b101;
									assign node160 = (inp[5]) ? 3'b001 : node161;
										assign node161 = (inp[0]) ? 3'b001 : 3'b101;
							assign node165 = (inp[3]) ? node181 : node166;
								assign node166 = (inp[4]) ? node174 : node167;
									assign node167 = (inp[5]) ? node169 : 3'b101;
										assign node169 = (inp[0]) ? node171 : 3'b101;
											assign node171 = (inp[2]) ? 3'b001 : 3'b101;
									assign node174 = (inp[0]) ? 3'b001 : node175;
										assign node175 = (inp[5]) ? 3'b001 : node176;
											assign node176 = (inp[2]) ? 3'b001 : 3'b101;
								assign node181 = (inp[1]) ? node183 : 3'b001;
									assign node183 = (inp[2]) ? 3'b001 : node184;
										assign node184 = (inp[5]) ? 3'b110 : 3'b001;
						assign node188 = (inp[8]) ? node208 : node189;
							assign node189 = (inp[4]) ? node197 : node190;
								assign node190 = (inp[5]) ? 3'b001 : node191;
									assign node191 = (inp[3]) ? 3'b001 : node192;
										assign node192 = (inp[0]) ? 3'b001 : 3'b101;
								assign node197 = (inp[3]) ? node199 : 3'b001;
									assign node199 = (inp[5]) ? 3'b110 : node200;
										assign node200 = (inp[0]) ? 3'b110 : node201;
											assign node201 = (inp[2]) ? node203 : 3'b001;
												assign node203 = (inp[1]) ? 3'b110 : 3'b001;
							assign node208 = (inp[3]) ? node224 : node209;
								assign node209 = (inp[4]) ? node217 : node210;
									assign node210 = (inp[5]) ? node212 : 3'b001;
										assign node212 = (inp[2]) ? node214 : 3'b001;
											assign node214 = (inp[0]) ? 3'b110 : 3'b001;
									assign node217 = (inp[2]) ? 3'b110 : node218;
										assign node218 = (inp[5]) ? 3'b110 : node219;
											assign node219 = (inp[1]) ? 3'b110 : 3'b001;
								assign node224 = (inp[5]) ? node226 : 3'b110;
									assign node226 = (inp[0]) ? node228 : 3'b110;
										assign node228 = (inp[4]) ? 3'b010 : 3'b110;
			assign node231 = (inp[10]) ? node399 : node232;
				assign node232 = (inp[7]) ? node300 : node233;
					assign node233 = (inp[11]) ? node267 : node234;
						assign node234 = (inp[3]) ? node252 : node235;
							assign node235 = (inp[8]) ? node245 : node236;
								assign node236 = (inp[2]) ? node238 : 3'b011;
									assign node238 = (inp[1]) ? node240 : 3'b101;
										assign node240 = (inp[0]) ? node242 : 3'b011;
											assign node242 = (inp[4]) ? 3'b101 : 3'b011;
								assign node245 = (inp[4]) ? 3'b101 : node246;
									assign node246 = (inp[0]) ? 3'b101 : node247;
										assign node247 = (inp[5]) ? 3'b101 : 3'b011;
							assign node252 = (inp[8]) ? node260 : node253;
								assign node253 = (inp[2]) ? node255 : 3'b101;
									assign node255 = (inp[0]) ? 3'b101 : node256;
										assign node256 = (inp[5]) ? 3'b101 : 3'b011;
								assign node260 = (inp[4]) ? 3'b001 : node261;
									assign node261 = (inp[0]) ? node263 : 3'b101;
										assign node263 = (inp[5]) ? 3'b001 : 3'b101;
						assign node267 = (inp[8]) ? node285 : node268;
							assign node268 = (inp[3]) ? node276 : node269;
								assign node269 = (inp[4]) ? node271 : 3'b101;
									assign node271 = (inp[5]) ? node273 : 3'b101;
										assign node273 = (inp[0]) ? 3'b001 : 3'b101;
								assign node276 = (inp[0]) ? 3'b001 : node277;
									assign node277 = (inp[1]) ? 3'b001 : node278;
										assign node278 = (inp[2]) ? 3'b001 : node279;
											assign node279 = (inp[4]) ? 3'b001 : 3'b101;
							assign node285 = (inp[3]) ? node287 : 3'b001;
								assign node287 = (inp[4]) ? 3'b110 : node288;
									assign node288 = (inp[0]) ? node294 : node289;
										assign node289 = (inp[5]) ? node291 : 3'b001;
											assign node291 = (inp[2]) ? 3'b110 : 3'b001;
										assign node294 = (inp[5]) ? 3'b110 : node295;
											assign node295 = (inp[2]) ? 3'b110 : 3'b001;
					assign node300 = (inp[11]) ? node350 : node301;
						assign node301 = (inp[8]) ? node331 : node302;
							assign node302 = (inp[3]) ? node316 : node303;
								assign node303 = (inp[4]) ? 3'b001 : node304;
									assign node304 = (inp[5]) ? node310 : node305;
										assign node305 = (inp[1]) ? node307 : 3'b101;
											assign node307 = (inp[0]) ? 3'b001 : 3'b101;
										assign node310 = (inp[0]) ? 3'b001 : node311;
											assign node311 = (inp[1]) ? 3'b001 : 3'b101;
								assign node316 = (inp[4]) ? node318 : 3'b001;
									assign node318 = (inp[0]) ? node324 : node319;
										assign node319 = (inp[5]) ? node321 : 3'b001;
											assign node321 = (inp[1]) ? 3'b110 : 3'b111;
										assign node324 = (inp[1]) ? 3'b110 : node325;
											assign node325 = (inp[2]) ? 3'b110 : node326;
												assign node326 = (inp[5]) ? 3'b110 : 3'b111;
							assign node331 = (inp[3]) ? node339 : node332;
								assign node332 = (inp[4]) ? node334 : 3'b001;
									assign node334 = (inp[5]) ? 3'b110 : node335;
										assign node335 = (inp[0]) ? 3'b110 : 3'b001;
								assign node339 = (inp[5]) ? node341 : 3'b110;
									assign node341 = (inp[0]) ? node343 : 3'b110;
										assign node343 = (inp[4]) ? node345 : 3'b110;
											assign node345 = (inp[2]) ? 3'b010 : node346;
												assign node346 = (inp[1]) ? 3'b010 : 3'b110;
						assign node350 = (inp[3]) ? node380 : node351;
							assign node351 = (inp[8]) ? node365 : node352;
								assign node352 = (inp[4]) ? 3'b110 : node353;
									assign node353 = (inp[0]) ? node359 : node354;
										assign node354 = (inp[5]) ? node356 : 3'b001;
											assign node356 = (inp[1]) ? 3'b110 : 3'b001;
										assign node359 = (inp[1]) ? 3'b110 : node360;
											assign node360 = (inp[5]) ? 3'b110 : 3'b001;
								assign node365 = (inp[1]) ? node373 : node366;
									assign node366 = (inp[2]) ? 3'b110 : node367;
										assign node367 = (inp[4]) ? node369 : 3'b110;
											assign node369 = (inp[5]) ? 3'b010 : 3'b110;
									assign node373 = (inp[2]) ? 3'b010 : node374;
										assign node374 = (inp[4]) ? node376 : 3'b110;
											assign node376 = (inp[5]) ? 3'b010 : 3'b110;
							assign node380 = (inp[8]) ? node388 : node381;
								assign node381 = (inp[4]) ? node383 : 3'b110;
									assign node383 = (inp[5]) ? 3'b010 : node384;
										assign node384 = (inp[0]) ? 3'b010 : 3'b110;
								assign node388 = (inp[5]) ? node390 : 3'b010;
									assign node390 = (inp[0]) ? node392 : 3'b010;
										assign node392 = (inp[1]) ? 3'b100 : node393;
											assign node393 = (inp[2]) ? node395 : 3'b010;
												assign node395 = (inp[4]) ? 3'b100 : 3'b010;
				assign node399 = (inp[7]) ? node447 : node400;
					assign node400 = (inp[11]) ? node430 : node401;
						assign node401 = (inp[8]) ? node411 : node402;
							assign node402 = (inp[3]) ? 3'b110 : node403;
								assign node403 = (inp[5]) ? node405 : 3'b001;
									assign node405 = (inp[4]) ? node407 : 3'b001;
										assign node407 = (inp[0]) ? 3'b110 : 3'b001;
							assign node411 = (inp[3]) ? node413 : 3'b110;
								assign node413 = (inp[4]) ? 3'b010 : node414;
									assign node414 = (inp[0]) ? node422 : node415;
										assign node415 = (inp[5]) ? node417 : 3'b110;
											assign node417 = (inp[1]) ? 3'b010 : node418;
												assign node418 = (inp[2]) ? 3'b010 : 3'b110;
										assign node422 = (inp[1]) ? 3'b010 : node423;
											assign node423 = (inp[2]) ? 3'b010 : node424;
												assign node424 = (inp[5]) ? 3'b010 : 3'b110;
						assign node430 = (inp[8]) ? node438 : node431;
							assign node431 = (inp[3]) ? 3'b010 : node432;
								assign node432 = (inp[2]) ? node434 : 3'b110;
									assign node434 = (inp[4]) ? 3'b010 : 3'b110;
							assign node438 = (inp[3]) ? node440 : 3'b010;
								assign node440 = (inp[4]) ? 3'b100 : node441;
									assign node441 = (inp[5]) ? 3'b100 : node442;
										assign node442 = (inp[0]) ? 3'b100 : 3'b010;
					assign node447 = (inp[11]) ? node487 : node448;
						assign node448 = (inp[3]) ? node466 : node449;
							assign node449 = (inp[8]) ? node457 : node450;
								assign node450 = (inp[4]) ? 3'b010 : node451;
									assign node451 = (inp[5]) ? 3'b010 : node452;
										assign node452 = (inp[2]) ? 3'b110 : 3'b010;
								assign node457 = (inp[4]) ? 3'b100 : node458;
									assign node458 = (inp[0]) ? node460 : 3'b010;
										assign node460 = (inp[5]) ? node462 : 3'b010;
											assign node462 = (inp[2]) ? 3'b100 : 3'b010;
							assign node466 = (inp[8]) ? node480 : node467;
								assign node467 = (inp[4]) ? node475 : node468;
									assign node468 = (inp[0]) ? node470 : 3'b010;
										assign node470 = (inp[2]) ? node472 : 3'b010;
											assign node472 = (inp[5]) ? 3'b100 : 3'b010;
									assign node475 = (inp[0]) ? 3'b100 : node476;
										assign node476 = (inp[5]) ? 3'b100 : 3'b010;
								assign node480 = (inp[0]) ? node482 : 3'b100;
									assign node482 = (inp[5]) ? node484 : 3'b100;
										assign node484 = (inp[4]) ? 3'b000 : 3'b100;
						assign node487 = (inp[8]) ? node511 : node488;
							assign node488 = (inp[3]) ? node496 : node489;
								assign node489 = (inp[5]) ? 3'b100 : node490;
									assign node490 = (inp[4]) ? 3'b100 : node491;
										assign node491 = (inp[0]) ? 3'b100 : 3'b010;
								assign node496 = (inp[4]) ? node504 : node497;
									assign node497 = (inp[2]) ? node499 : 3'b100;
										assign node499 = (inp[0]) ? node501 : 3'b100;
											assign node501 = (inp[5]) ? 3'b000 : 3'b100;
									assign node504 = (inp[5]) ? 3'b000 : node505;
										assign node505 = (inp[1]) ? 3'b000 : node506;
											assign node506 = (inp[0]) ? 3'b000 : 3'b100;
							assign node511 = (inp[4]) ? 3'b000 : node512;
								assign node512 = (inp[3]) ? 3'b000 : node513;
									assign node513 = (inp[0]) ? node515 : 3'b100;
										assign node515 = (inp[5]) ? 3'b000 : 3'b100;
		assign node520 = (inp[6]) ? node728 : node521;
			assign node521 = (inp[10]) ? node641 : node522;
				assign node522 = (inp[7]) ? node564 : node523;
					assign node523 = (inp[11]) ? node545 : node524;
						assign node524 = (inp[3]) ? node536 : node525;
							assign node525 = (inp[8]) ? 3'b001 : node526;
								assign node526 = (inp[5]) ? node528 : 3'b101;
									assign node528 = (inp[4]) ? node530 : 3'b101;
										assign node530 = (inp[2]) ? 3'b001 : node531;
											assign node531 = (inp[0]) ? 3'b001 : 3'b101;
							assign node536 = (inp[8]) ? node538 : 3'b001;
								assign node538 = (inp[4]) ? 3'b110 : node539;
									assign node539 = (inp[0]) ? 3'b110 : node540;
										assign node540 = (inp[5]) ? 3'b110 : 3'b001;
						assign node545 = (inp[8]) ? node555 : node546;
							assign node546 = (inp[3]) ? 3'b110 : node547;
								assign node547 = (inp[4]) ? node549 : 3'b001;
									assign node549 = (inp[0]) ? 3'b110 : node550;
										assign node550 = (inp[5]) ? 3'b110 : 3'b001;
							assign node555 = (inp[3]) ? node557 : 3'b110;
								assign node557 = (inp[5]) ? 3'b010 : node558;
									assign node558 = (inp[0]) ? 3'b010 : node559;
										assign node559 = (inp[4]) ? 3'b010 : 3'b110;
					assign node564 = (inp[11]) ? node610 : node565;
						assign node565 = (inp[8]) ? node589 : node566;
							assign node566 = (inp[3]) ? node574 : node567;
								assign node567 = (inp[4]) ? 3'b110 : node568;
									assign node568 = (inp[0]) ? 3'b110 : node569;
										assign node569 = (inp[5]) ? 3'b110 : 3'b001;
								assign node574 = (inp[4]) ? node582 : node575;
									assign node575 = (inp[5]) ? node577 : 3'b110;
										assign node577 = (inp[0]) ? node579 : 3'b110;
											assign node579 = (inp[1]) ? 3'b010 : 3'b110;
									assign node582 = (inp[5]) ? 3'b010 : node583;
										assign node583 = (inp[0]) ? 3'b010 : node584;
											assign node584 = (inp[1]) ? 3'b010 : 3'b110;
							assign node589 = (inp[4]) ? node597 : node590;
								assign node590 = (inp[3]) ? 3'b010 : node591;
									assign node591 = (inp[0]) ? node593 : 3'b110;
										assign node593 = (inp[5]) ? 3'b010 : 3'b110;
								assign node597 = (inp[3]) ? node599 : 3'b010;
									assign node599 = (inp[2]) ? node605 : node600;
										assign node600 = (inp[5]) ? node602 : 3'b010;
											assign node602 = (inp[0]) ? 3'b100 : 3'b010;
										assign node605 = (inp[5]) ? 3'b100 : node606;
											assign node606 = (inp[0]) ? 3'b100 : 3'b010;
						assign node610 = (inp[8]) ? node624 : node611;
							assign node611 = (inp[3]) ? node615 : node612;
								assign node612 = (inp[4]) ? 3'b010 : 3'b110;
								assign node615 = (inp[4]) ? 3'b100 : node616;
									assign node616 = (inp[2]) ? node618 : 3'b010;
										assign node618 = (inp[0]) ? node620 : 3'b010;
											assign node620 = (inp[5]) ? 3'b100 : 3'b010;
							assign node624 = (inp[4]) ? node632 : node625;
								assign node625 = (inp[3]) ? 3'b100 : node626;
									assign node626 = (inp[5]) ? node628 : 3'b010;
										assign node628 = (inp[0]) ? 3'b100 : 3'b010;
								assign node632 = (inp[3]) ? node634 : 3'b100;
									assign node634 = (inp[0]) ? node636 : 3'b100;
										assign node636 = (inp[5]) ? 3'b000 : node637;
											assign node637 = (inp[2]) ? 3'b000 : 3'b100;
				assign node641 = (inp[7]) ? node703 : node642;
					assign node642 = (inp[11]) ? node672 : node643;
						assign node643 = (inp[8]) ? node651 : node644;
							assign node644 = (inp[3]) ? 3'b010 : node645;
								assign node645 = (inp[4]) ? node647 : 3'b110;
									assign node647 = (inp[1]) ? 3'b010 : 3'b110;
							assign node651 = (inp[3]) ? node663 : node652;
								assign node652 = (inp[2]) ? node654 : 3'b010;
									assign node654 = (inp[1]) ? node656 : 3'b100;
										assign node656 = (inp[0]) ? node658 : 3'b010;
											assign node658 = (inp[4]) ? node660 : 3'b010;
												assign node660 = (inp[5]) ? 3'b100 : 3'b010;
								assign node663 = (inp[2]) ? 3'b100 : node664;
									assign node664 = (inp[4]) ? 3'b100 : node665;
										assign node665 = (inp[5]) ? 3'b100 : node666;
											assign node666 = (inp[0]) ? 3'b100 : 3'b010;
						assign node672 = (inp[8]) ? node684 : node673;
							assign node673 = (inp[3]) ? node677 : node674;
								assign node674 = (inp[4]) ? 3'b100 : 3'b000;
								assign node677 = (inp[4]) ? node679 : 3'b100;
									assign node679 = (inp[5]) ? node681 : 3'b100;
										assign node681 = (inp[0]) ? 3'b000 : 3'b100;
							assign node684 = (inp[3]) ? node694 : node685;
								assign node685 = (inp[2]) ? node687 : 3'b100;
									assign node687 = (inp[1]) ? node689 : 3'b000;
										assign node689 = (inp[0]) ? node691 : 3'b100;
											assign node691 = (inp[4]) ? 3'b000 : 3'b100;
								assign node694 = (inp[2]) ? 3'b000 : node695;
									assign node695 = (inp[5]) ? 3'b000 : node696;
										assign node696 = (inp[4]) ? 3'b000 : node697;
											assign node697 = (inp[0]) ? 3'b000 : 3'b100;
					assign node703 = (inp[11]) ? 3'b000 : node704;
						assign node704 = (inp[8]) ? node720 : node705;
							assign node705 = (inp[3]) ? node713 : node706;
								assign node706 = (inp[5]) ? 3'b100 : node707;
									assign node707 = (inp[4]) ? 3'b100 : node708;
										assign node708 = (inp[0]) ? 3'b100 : 3'b000;
								assign node713 = (inp[4]) ? 3'b000 : node714;
									assign node714 = (inp[0]) ? node716 : 3'b100;
										assign node716 = (inp[5]) ? 3'b000 : 3'b100;
							assign node720 = (inp[5]) ? 3'b000 : node721;
								assign node721 = (inp[4]) ? 3'b000 : node722;
									assign node722 = (inp[0]) ? 3'b000 : 3'b100;
			assign node728 = (inp[7]) ? 3'b000 : node729;
				assign node729 = (inp[10]) ? 3'b000 : node730;
					assign node730 = (inp[11]) ? node760 : node731;
						assign node731 = (inp[8]) ? node739 : node732;
							assign node732 = (inp[3]) ? 3'b100 : node733;
								assign node733 = (inp[1]) ? node735 : 3'b010;
									assign node735 = (inp[4]) ? 3'b100 : 3'b010;
							assign node739 = (inp[3]) ? node751 : node740;
								assign node740 = (inp[2]) ? node742 : 3'b100;
									assign node742 = (inp[1]) ? node744 : 3'b000;
										assign node744 = (inp[5]) ? node746 : 3'b100;
											assign node746 = (inp[0]) ? node748 : 3'b100;
												assign node748 = (inp[4]) ? 3'b000 : 3'b100;
								assign node751 = (inp[2]) ? 3'b000 : node752;
									assign node752 = (inp[4]) ? 3'b000 : node753;
										assign node753 = (inp[0]) ? 3'b000 : node754;
											assign node754 = (inp[5]) ? 3'b000 : 3'b100;
						assign node760 = (inp[3]) ? 3'b000 : node761;
							assign node761 = (inp[8]) ? 3'b000 : node762;
								assign node762 = (inp[4]) ? node764 : 3'b100;
									assign node764 = (inp[2]) ? 3'b000 : 3'b100;

endmodule