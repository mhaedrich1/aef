module dtc_split05_bm48 (
	input  wire [14-1:0] inp,
	output wire [14-1:0] outp
);

	wire [14-1:0] node1;
	wire [14-1:0] node2;
	wire [14-1:0] node3;
	wire [14-1:0] node4;
	wire [14-1:0] node7;
	wire [14-1:0] node8;
	wire [14-1:0] node12;
	wire [14-1:0] node13;
	wire [14-1:0] node14;
	wire [14-1:0] node18;
	wire [14-1:0] node19;
	wire [14-1:0] node22;
	wire [14-1:0] node25;
	wire [14-1:0] node26;
	wire [14-1:0] node27;
	wire [14-1:0] node28;
	wire [14-1:0] node31;
	wire [14-1:0] node34;
	wire [14-1:0] node35;
	wire [14-1:0] node38;
	wire [14-1:0] node41;
	wire [14-1:0] node42;
	wire [14-1:0] node43;
	wire [14-1:0] node46;
	wire [14-1:0] node49;
	wire [14-1:0] node50;
	wire [14-1:0] node54;
	wire [14-1:0] node55;
	wire [14-1:0] node56;
	wire [14-1:0] node57;
	wire [14-1:0] node60;
	wire [14-1:0] node62;
	wire [14-1:0] node65;
	wire [14-1:0] node66;
	wire [14-1:0] node67;
	wire [14-1:0] node71;
	wire [14-1:0] node72;
	wire [14-1:0] node75;
	wire [14-1:0] node78;
	wire [14-1:0] node79;
	wire [14-1:0] node80;
	wire [14-1:0] node81;
	wire [14-1:0] node85;
	wire [14-1:0] node86;
	wire [14-1:0] node89;
	wire [14-1:0] node92;
	wire [14-1:0] node93;
	wire [14-1:0] node94;
	wire [14-1:0] node98;
	wire [14-1:0] node99;

	assign outp = (inp[10]) ? node54 : node1;
		assign node1 = (inp[8]) ? node25 : node2;
			assign node2 = (inp[13]) ? node12 : node3;
				assign node3 = (inp[11]) ? node7 : node4;
					assign node4 = (inp[12]) ? 14'b00000000000000 : 14'b00000100000011;
					assign node7 = (inp[9]) ? 14'b00000000000000 : node8;
						assign node8 = (inp[2]) ? 14'b00000000000000 : 14'b00000000000000;
				assign node12 = (inp[7]) ? node18 : node13;
					assign node13 = (inp[4]) ? 14'b00000000000000 : node14;
						assign node14 = (inp[5]) ? 14'b00000000000000 : 14'b00000000000000;
					assign node18 = (inp[3]) ? node22 : node19;
						assign node19 = (inp[1]) ? 14'b00000000000000 : 14'b00000000000000;
						assign node22 = (inp[11]) ? 14'b00000000000000 : 14'b00000000000000;
			assign node25 = (inp[11]) ? node41 : node26;
				assign node26 = (inp[12]) ? node34 : node27;
					assign node27 = (inp[5]) ? node31 : node28;
						assign node28 = (inp[4]) ? 14'b00000000000000 : 14'b00000000000000;
						assign node31 = (inp[3]) ? 14'b00000000000000 : 14'b00000000000000;
					assign node34 = (inp[6]) ? node38 : node35;
						assign node35 = (inp[4]) ? 14'b00000000000000 : 14'b00000000000000;
						assign node38 = (inp[13]) ? 14'b00000000000000 : 14'b00000000000000;
				assign node41 = (inp[13]) ? node49 : node42;
					assign node42 = (inp[0]) ? node46 : node43;
						assign node43 = (inp[5]) ? 14'b00000000000000 : 14'b00000000000000;
						assign node46 = (inp[3]) ? 14'b00000000000000 : 14'b00000000000000;
					assign node49 = (inp[12]) ? 14'b01000000010100 : node50;
						assign node50 = (inp[0]) ? 14'b00000000000000 : 14'b00000000001100;
		assign node54 = (inp[11]) ? node78 : node55;
			assign node55 = (inp[8]) ? node65 : node56;
				assign node56 = (inp[12]) ? node60 : node57;
					assign node57 = (inp[13]) ? 14'b00000000000000 : 14'b10000100001000;
					assign node60 = (inp[1]) ? node62 : 14'b00000000000000;
						assign node62 = (inp[9]) ? 14'b00000000000000 : 14'b00000000000000;
				assign node65 = (inp[6]) ? node71 : node66;
					assign node66 = (inp[2]) ? 14'b00000000000000 : node67;
						assign node67 = (inp[0]) ? 14'b00000000000000 : 14'b00000000000000;
					assign node71 = (inp[12]) ? node75 : node72;
						assign node72 = (inp[5]) ? 14'b00000000000000 : 14'b00000000000000;
						assign node75 = (inp[13]) ? 14'b00000000000000 : 14'b00000000000000;
			assign node78 = (inp[8]) ? node92 : node79;
				assign node79 = (inp[1]) ? node85 : node80;
					assign node80 = (inp[13]) ? 14'b00000000000000 : node81;
						assign node81 = (inp[12]) ? 14'b00000000000000 : 14'b00000000000000;
					assign node85 = (inp[12]) ? node89 : node86;
						assign node86 = (inp[5]) ? 14'b00000000000000 : 14'b00000000000000;
						assign node89 = (inp[2]) ? 14'b00000000000000 : 14'b00000000000000;
				assign node92 = (inp[13]) ? node98 : node93;
					assign node93 = (inp[6]) ? 14'b00000000000000 : node94;
						assign node94 = (inp[2]) ? 14'b00000000000000 : 14'b00000000000000;
					assign node98 = (inp[12]) ? 14'b10000100001000 : node99;
						assign node99 = (inp[1]) ? 14'b00000000000000 : 14'b00000000000000;

endmodule