module dtc_split33_bm87 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node7;
	wire [3-1:0] node9;
	wire [3-1:0] node10;
	wire [3-1:0] node17;
	wire [3-1:0] node18;
	wire [3-1:0] node19;
	wire [3-1:0] node20;
	wire [3-1:0] node21;
	wire [3-1:0] node24;
	wire [3-1:0] node25;
	wire [3-1:0] node27;
	wire [3-1:0] node28;
	wire [3-1:0] node30;
	wire [3-1:0] node32;
	wire [3-1:0] node35;
	wire [3-1:0] node38;
	wire [3-1:0] node39;
	wire [3-1:0] node40;
	wire [3-1:0] node42;
	wire [3-1:0] node43;
	wire [3-1:0] node48;
	wire [3-1:0] node51;
	wire [3-1:0] node53;
	wire [3-1:0] node54;
	wire [3-1:0] node55;
	wire [3-1:0] node58;
	wire [3-1:0] node60;
	wire [3-1:0] node61;
	wire [3-1:0] node64;
	wire [3-1:0] node67;
	wire [3-1:0] node69;
	wire [3-1:0] node70;
	wire [3-1:0] node73;
	wire [3-1:0] node76;
	wire [3-1:0] node77;
	wire [3-1:0] node78;
	wire [3-1:0] node79;
	wire [3-1:0] node80;
	wire [3-1:0] node83;
	wire [3-1:0] node85;
	wire [3-1:0] node88;
	wire [3-1:0] node89;
	wire [3-1:0] node92;
	wire [3-1:0] node94;
	wire [3-1:0] node97;
	wire [3-1:0] node98;
	wire [3-1:0] node99;
	wire [3-1:0] node103;
	wire [3-1:0] node104;
	wire [3-1:0] node105;
	wire [3-1:0] node108;
	wire [3-1:0] node110;
	wire [3-1:0] node113;
	wire [3-1:0] node115;
	wire [3-1:0] node118;
	wire [3-1:0] node119;
	wire [3-1:0] node120;
	wire [3-1:0] node122;
	wire [3-1:0] node124;
	wire [3-1:0] node129;
	wire [3-1:0] node130;
	wire [3-1:0] node131;
	wire [3-1:0] node132;
	wire [3-1:0] node133;
	wire [3-1:0] node136;
	wire [3-1:0] node139;
	wire [3-1:0] node141;
	wire [3-1:0] node142;
	wire [3-1:0] node143;
	wire [3-1:0] node147;
	wire [3-1:0] node148;
	wire [3-1:0] node151;
	wire [3-1:0] node156;
	wire [3-1:0] node157;
	wire [3-1:0] node158;
	wire [3-1:0] node159;
	wire [3-1:0] node160;
	wire [3-1:0] node161;
	wire [3-1:0] node162;
	wire [3-1:0] node163;
	wire [3-1:0] node164;
	wire [3-1:0] node168;
	wire [3-1:0] node169;
	wire [3-1:0] node173;
	wire [3-1:0] node174;
	wire [3-1:0] node177;
	wire [3-1:0] node178;
	wire [3-1:0] node182;
	wire [3-1:0] node183;
	wire [3-1:0] node184;
	wire [3-1:0] node185;
	wire [3-1:0] node187;
	wire [3-1:0] node191;
	wire [3-1:0] node192;
	wire [3-1:0] node196;
	wire [3-1:0] node197;
	wire [3-1:0] node199;
	wire [3-1:0] node203;
	wire [3-1:0] node204;
	wire [3-1:0] node205;
	wire [3-1:0] node206;
	wire [3-1:0] node207;
	wire [3-1:0] node211;
	wire [3-1:0] node213;
	wire [3-1:0] node214;
	wire [3-1:0] node215;
	wire [3-1:0] node220;
	wire [3-1:0] node221;
	wire [3-1:0] node224;
	wire [3-1:0] node225;
	wire [3-1:0] node228;
	wire [3-1:0] node230;
	wire [3-1:0] node233;
	wire [3-1:0] node234;
	wire [3-1:0] node235;
	wire [3-1:0] node236;
	wire [3-1:0] node237;
	wire [3-1:0] node241;
	wire [3-1:0] node244;
	wire [3-1:0] node246;
	wire [3-1:0] node249;
	wire [3-1:0] node250;
	wire [3-1:0] node253;
	wire [3-1:0] node254;
	wire [3-1:0] node256;
	wire [3-1:0] node260;
	wire [3-1:0] node261;
	wire [3-1:0] node262;
	wire [3-1:0] node263;
	wire [3-1:0] node264;
	wire [3-1:0] node267;
	wire [3-1:0] node270;
	wire [3-1:0] node271;
	wire [3-1:0] node273;
	wire [3-1:0] node274;
	wire [3-1:0] node278;
	wire [3-1:0] node280;
	wire [3-1:0] node283;
	wire [3-1:0] node284;
	wire [3-1:0] node286;
	wire [3-1:0] node288;
	wire [3-1:0] node291;
	wire [3-1:0] node293;
	wire [3-1:0] node294;
	wire [3-1:0] node298;
	wire [3-1:0] node299;
	wire [3-1:0] node300;
	wire [3-1:0] node301;
	wire [3-1:0] node305;
	wire [3-1:0] node307;
	wire [3-1:0] node308;
	wire [3-1:0] node311;
	wire [3-1:0] node314;
	wire [3-1:0] node315;
	wire [3-1:0] node316;
	wire [3-1:0] node317;
	wire [3-1:0] node320;
	wire [3-1:0] node324;
	wire [3-1:0] node325;
	wire [3-1:0] node326;
	wire [3-1:0] node329;
	wire [3-1:0] node330;
	wire [3-1:0] node334;
	wire [3-1:0] node335;
	wire [3-1:0] node339;
	wire [3-1:0] node340;
	wire [3-1:0] node341;
	wire [3-1:0] node343;
	wire [3-1:0] node344;
	wire [3-1:0] node345;
	wire [3-1:0] node347;
	wire [3-1:0] node352;
	wire [3-1:0] node353;
	wire [3-1:0] node354;
	wire [3-1:0] node356;
	wire [3-1:0] node357;
	wire [3-1:0] node361;
	wire [3-1:0] node362;
	wire [3-1:0] node365;
	wire [3-1:0] node366;
	wire [3-1:0] node367;
	wire [3-1:0] node372;
	wire [3-1:0] node373;
	wire [3-1:0] node374;
	wire [3-1:0] node375;
	wire [3-1:0] node379;
	wire [3-1:0] node382;
	wire [3-1:0] node383;
	wire [3-1:0] node386;
	wire [3-1:0] node387;
	wire [3-1:0] node389;
	wire [3-1:0] node390;
	wire [3-1:0] node395;
	wire [3-1:0] node396;
	wire [3-1:0] node397;
	wire [3-1:0] node398;
	wire [3-1:0] node399;
	wire [3-1:0] node402;
	wire [3-1:0] node403;
	wire [3-1:0] node407;
	wire [3-1:0] node408;
	wire [3-1:0] node409;
	wire [3-1:0] node413;
	wire [3-1:0] node415;
	wire [3-1:0] node417;
	wire [3-1:0] node420;
	wire [3-1:0] node421;
	wire [3-1:0] node423;
	wire [3-1:0] node424;
	wire [3-1:0] node425;
	wire [3-1:0] node428;
	wire [3-1:0] node432;
	wire [3-1:0] node433;
	wire [3-1:0] node434;
	wire [3-1:0] node437;
	wire [3-1:0] node439;
	wire [3-1:0] node442;
	wire [3-1:0] node443;
	wire [3-1:0] node446;
	wire [3-1:0] node449;
	wire [3-1:0] node450;
	wire [3-1:0] node451;
	wire [3-1:0] node452;
	wire [3-1:0] node453;
	wire [3-1:0] node455;
	wire [3-1:0] node460;
	wire [3-1:0] node461;
	wire [3-1:0] node462;
	wire [3-1:0] node463;
	wire [3-1:0] node468;
	wire [3-1:0] node470;
	wire [3-1:0] node473;
	wire [3-1:0] node474;
	wire [3-1:0] node475;
	wire [3-1:0] node476;
	wire [3-1:0] node477;
	wire [3-1:0] node482;
	wire [3-1:0] node483;
	wire [3-1:0] node487;
	wire [3-1:0] node489;
	wire [3-1:0] node490;
	wire [3-1:0] node491;
	wire [3-1:0] node496;
	wire [3-1:0] node497;
	wire [3-1:0] node498;
	wire [3-1:0] node499;
	wire [3-1:0] node500;
	wire [3-1:0] node501;
	wire [3-1:0] node502;
	wire [3-1:0] node504;
	wire [3-1:0] node505;
	wire [3-1:0] node509;
	wire [3-1:0] node510;
	wire [3-1:0] node514;
	wire [3-1:0] node515;
	wire [3-1:0] node517;
	wire [3-1:0] node518;
	wire [3-1:0] node522;
	wire [3-1:0] node524;
	wire [3-1:0] node525;
	wire [3-1:0] node526;
	wire [3-1:0] node531;
	wire [3-1:0] node532;
	wire [3-1:0] node533;
	wire [3-1:0] node535;
	wire [3-1:0] node536;
	wire [3-1:0] node537;
	wire [3-1:0] node542;
	wire [3-1:0] node544;
	wire [3-1:0] node545;
	wire [3-1:0] node549;
	wire [3-1:0] node550;
	wire [3-1:0] node553;
	wire [3-1:0] node556;
	wire [3-1:0] node557;
	wire [3-1:0] node558;
	wire [3-1:0] node559;
	wire [3-1:0] node562;
	wire [3-1:0] node563;
	wire [3-1:0] node567;
	wire [3-1:0] node569;
	wire [3-1:0] node570;
	wire [3-1:0] node573;
	wire [3-1:0] node576;
	wire [3-1:0] node578;
	wire [3-1:0] node579;
	wire [3-1:0] node580;
	wire [3-1:0] node585;
	wire [3-1:0] node586;
	wire [3-1:0] node587;
	wire [3-1:0] node588;
	wire [3-1:0] node589;
	wire [3-1:0] node591;
	wire [3-1:0] node593;
	wire [3-1:0] node596;
	wire [3-1:0] node599;
	wire [3-1:0] node600;
	wire [3-1:0] node604;
	wire [3-1:0] node605;
	wire [3-1:0] node607;
	wire [3-1:0] node609;
	wire [3-1:0] node612;
	wire [3-1:0] node613;
	wire [3-1:0] node616;
	wire [3-1:0] node618;
	wire [3-1:0] node621;
	wire [3-1:0] node622;
	wire [3-1:0] node623;
	wire [3-1:0] node624;
	wire [3-1:0] node627;
	wire [3-1:0] node629;
	wire [3-1:0] node630;
	wire [3-1:0] node634;
	wire [3-1:0] node635;
	wire [3-1:0] node638;
	wire [3-1:0] node641;
	wire [3-1:0] node642;
	wire [3-1:0] node643;
	wire [3-1:0] node644;
	wire [3-1:0] node648;
	wire [3-1:0] node651;
	wire [3-1:0] node652;
	wire [3-1:0] node654;
	wire [3-1:0] node655;
	wire [3-1:0] node659;
	wire [3-1:0] node662;
	wire [3-1:0] node663;
	wire [3-1:0] node664;
	wire [3-1:0] node666;
	wire [3-1:0] node667;
	wire [3-1:0] node668;
	wire [3-1:0] node669;
	wire [3-1:0] node670;
	wire [3-1:0] node674;
	wire [3-1:0] node676;
	wire [3-1:0] node679;
	wire [3-1:0] node680;
	wire [3-1:0] node681;
	wire [3-1:0] node687;
	wire [3-1:0] node688;
	wire [3-1:0] node689;
	wire [3-1:0] node690;
	wire [3-1:0] node693;
	wire [3-1:0] node696;
	wire [3-1:0] node698;
	wire [3-1:0] node699;
	wire [3-1:0] node702;
	wire [3-1:0] node705;
	wire [3-1:0] node706;
	wire [3-1:0] node707;
	wire [3-1:0] node709;
	wire [3-1:0] node710;
	wire [3-1:0] node714;
	wire [3-1:0] node716;
	wire [3-1:0] node718;
	wire [3-1:0] node721;
	wire [3-1:0] node722;
	wire [3-1:0] node725;
	wire [3-1:0] node728;
	wire [3-1:0] node730;
	wire [3-1:0] node732;
	wire [3-1:0] node733;
	wire [3-1:0] node735;
	wire [3-1:0] node737;

	assign outp = (inp[6]) ? node156 : node1;
		assign node1 = (inp[7]) ? node17 : node2;
			assign node2 = (inp[1]) ? 3'b000 : node3;
				assign node3 = (inp[10]) ? 3'b000 : node4;
					assign node4 = (inp[9]) ? 3'b000 : node5;
						assign node5 = (inp[0]) ? node7 : 3'b000;
							assign node7 = (inp[8]) ? node9 : 3'b000;
								assign node9 = (inp[11]) ? 3'b100 : node10;
									assign node10 = (inp[2]) ? 3'b000 : 3'b100;
			assign node17 = (inp[9]) ? node129 : node18;
				assign node18 = (inp[0]) ? node76 : node19;
					assign node19 = (inp[10]) ? node51 : node20;
						assign node20 = (inp[1]) ? node24 : node21;
							assign node21 = (inp[11]) ? 3'b001 : 3'b101;
							assign node24 = (inp[8]) ? node38 : node25;
								assign node25 = (inp[5]) ? node27 : 3'b010;
									assign node27 = (inp[4]) ? node35 : node28;
										assign node28 = (inp[3]) ? node30 : 3'b110;
											assign node30 = (inp[2]) ? node32 : 3'b010;
												assign node32 = (inp[11]) ? 3'b110 : 3'b010;
										assign node35 = (inp[3]) ? 3'b110 : 3'b010;
								assign node38 = (inp[11]) ? node48 : node39;
									assign node39 = (inp[4]) ? 3'b001 : node40;
										assign node40 = (inp[2]) ? node42 : 3'b001;
											assign node42 = (inp[5]) ? 3'b110 : node43;
												assign node43 = (inp[3]) ? 3'b110 : 3'b001;
									assign node48 = (inp[4]) ? 3'b110 : 3'b010;
						assign node51 = (inp[1]) ? node53 : 3'b110;
							assign node53 = (inp[4]) ? node67 : node54;
								assign node54 = (inp[8]) ? node58 : node55;
									assign node55 = (inp[3]) ? 3'b100 : 3'b000;
									assign node58 = (inp[11]) ? node60 : 3'b010;
										assign node60 = (inp[5]) ? node64 : node61;
											assign node61 = (inp[2]) ? 3'b110 : 3'b010;
											assign node64 = (inp[2]) ? 3'b010 : 3'b110;
								assign node67 = (inp[5]) ? node69 : 3'b100;
									assign node69 = (inp[8]) ? node73 : node70;
										assign node70 = (inp[11]) ? 3'b000 : 3'b100;
										assign node73 = (inp[11]) ? 3'b100 : 3'b010;
					assign node76 = (inp[10]) ? node118 : node77;
						assign node77 = (inp[1]) ? node97 : node78;
							assign node78 = (inp[11]) ? node88 : node79;
								assign node79 = (inp[8]) ? node83 : node80;
									assign node80 = (inp[2]) ? 3'b100 : 3'b010;
									assign node83 = (inp[2]) ? node85 : 3'b110;
										assign node85 = (inp[5]) ? 3'b010 : 3'b110;
								assign node88 = (inp[2]) ? node92 : node89;
									assign node89 = (inp[8]) ? 3'b010 : 3'b100;
									assign node92 = (inp[8]) ? node94 : 3'b010;
										assign node94 = (inp[5]) ? 3'b010 : 3'b100;
							assign node97 = (inp[8]) ? node103 : node98;
								assign node98 = (inp[2]) ? 3'b000 : node99;
									assign node99 = (inp[11]) ? 3'b000 : 3'b100;
								assign node103 = (inp[2]) ? node113 : node104;
									assign node104 = (inp[11]) ? node108 : node105;
										assign node105 = (inp[5]) ? 3'b100 : 3'b010;
										assign node108 = (inp[3]) ? node110 : 3'b100;
											assign node110 = (inp[4]) ? 3'b000 : 3'b100;
									assign node113 = (inp[5]) ? node115 : 3'b100;
										assign node115 = (inp[4]) ? 3'b000 : 3'b100;
						assign node118 = (inp[11]) ? 3'b000 : node119;
							assign node119 = (inp[1]) ? 3'b000 : node120;
								assign node120 = (inp[8]) ? node122 : 3'b000;
									assign node122 = (inp[2]) ? node124 : 3'b100;
										assign node124 = (inp[4]) ? 3'b000 : 3'b100;
				assign node129 = (inp[0]) ? 3'b000 : node130;
					assign node130 = (inp[10]) ? 3'b000 : node131;
						assign node131 = (inp[1]) ? node139 : node132;
							assign node132 = (inp[2]) ? node136 : node133;
								assign node133 = (inp[11]) ? 3'b110 : 3'b010;
								assign node136 = (inp[11]) ? 3'b000 : 3'b100;
							assign node139 = (inp[8]) ? node141 : 3'b000;
								assign node141 = (inp[3]) ? node147 : node142;
									assign node142 = (inp[4]) ? 3'b000 : node143;
										assign node143 = (inp[2]) ? 3'b000 : 3'b100;
									assign node147 = (inp[11]) ? node151 : node148;
										assign node148 = (inp[2]) ? 3'b100 : 3'b000;
										assign node151 = (inp[5]) ? 3'b100 : 3'b000;
		assign node156 = (inp[9]) ? node496 : node157;
			assign node157 = (inp[7]) ? node339 : node158;
				assign node158 = (inp[0]) ? node260 : node159;
					assign node159 = (inp[10]) ? node203 : node160;
						assign node160 = (inp[8]) ? node182 : node161;
							assign node161 = (inp[11]) ? node173 : node162;
								assign node162 = (inp[1]) ? node168 : node163;
									assign node163 = (inp[2]) ? 3'b011 : node164;
										assign node164 = (inp[5]) ? 3'b011 : 3'b111;
									assign node168 = (inp[3]) ? 3'b001 : node169;
										assign node169 = (inp[4]) ? 3'b101 : 3'b110;
								assign node173 = (inp[1]) ? node177 : node174;
									assign node174 = (inp[3]) ? 3'b101 : 3'b001;
									assign node177 = (inp[3]) ? 3'b001 : node178;
										assign node178 = (inp[2]) ? 3'b001 : 3'b101;
							assign node182 = (inp[1]) ? node196 : node183;
								assign node183 = (inp[11]) ? node191 : node184;
									assign node184 = (inp[2]) ? 3'b111 : node185;
										assign node185 = (inp[5]) ? node187 : 3'b011;
											assign node187 = (inp[3]) ? 3'b111 : 3'b011;
									assign node191 = (inp[2]) ? 3'b011 : node192;
										assign node192 = (inp[3]) ? 3'b011 : 3'b111;
								assign node196 = (inp[11]) ? 3'b101 : node197;
									assign node197 = (inp[4]) ? node199 : 3'b011;
										assign node199 = (inp[5]) ? 3'b101 : 3'b011;
						assign node203 = (inp[1]) ? node233 : node204;
							assign node204 = (inp[8]) ? node220 : node205;
								assign node205 = (inp[5]) ? node211 : node206;
									assign node206 = (inp[4]) ? 3'b001 : node207;
										assign node207 = (inp[11]) ? 3'b001 : 3'b101;
									assign node211 = (inp[11]) ? node213 : 3'b001;
										assign node213 = (inp[4]) ? 3'b110 : node214;
											assign node214 = (inp[2]) ? 3'b010 : node215;
												assign node215 = (inp[3]) ? 3'b000 : 3'b001;
								assign node220 = (inp[11]) ? node224 : node221;
									assign node221 = (inp[2]) ? 3'b101 : 3'b011;
									assign node224 = (inp[2]) ? node228 : node225;
										assign node225 = (inp[4]) ? 3'b001 : 3'b101;
										assign node228 = (inp[3]) ? node230 : 3'b001;
											assign node230 = (inp[5]) ? 3'b001 : 3'b011;
							assign node233 = (inp[8]) ? node249 : node234;
								assign node234 = (inp[11]) ? node244 : node235;
									assign node235 = (inp[4]) ? node241 : node236;
										assign node236 = (inp[2]) ? 3'b110 : node237;
											assign node237 = (inp[3]) ? 3'b110 : 3'b001;
										assign node241 = (inp[2]) ? 3'b010 : 3'b110;
									assign node244 = (inp[4]) ? node246 : 3'b010;
										assign node246 = (inp[3]) ? 3'b100 : 3'b010;
								assign node249 = (inp[11]) ? node253 : node250;
									assign node250 = (inp[3]) ? 3'b001 : 3'b101;
									assign node253 = (inp[4]) ? 3'b001 : node254;
										assign node254 = (inp[5]) ? node256 : 3'b110;
											assign node256 = (inp[3]) ? 3'b110 : 3'b010;
					assign node260 = (inp[10]) ? node298 : node261;
						assign node261 = (inp[1]) ? node283 : node262;
							assign node262 = (inp[2]) ? node270 : node263;
								assign node263 = (inp[11]) ? node267 : node264;
									assign node264 = (inp[8]) ? 3'b101 : 3'b001;
									assign node267 = (inp[8]) ? 3'b001 : 3'b110;
								assign node270 = (inp[8]) ? node278 : node271;
									assign node271 = (inp[11]) ? node273 : 3'b110;
										assign node273 = (inp[3]) ? 3'b010 : node274;
											assign node274 = (inp[4]) ? 3'b010 : 3'b110;
									assign node278 = (inp[11]) ? node280 : 3'b001;
										assign node280 = (inp[3]) ? 3'b110 : 3'b101;
							assign node283 = (inp[5]) ? node291 : node284;
								assign node284 = (inp[2]) ? node286 : 3'b110;
									assign node286 = (inp[11]) ? node288 : 3'b110;
										assign node288 = (inp[8]) ? 3'b001 : 3'b010;
								assign node291 = (inp[2]) ? node293 : 3'b010;
									assign node293 = (inp[8]) ? 3'b010 : node294;
										assign node294 = (inp[11]) ? 3'b100 : 3'b010;
						assign node298 = (inp[11]) ? node314 : node299;
							assign node299 = (inp[8]) ? node305 : node300;
								assign node300 = (inp[1]) ? 3'b100 : node301;
									assign node301 = (inp[2]) ? 3'b100 : 3'b010;
								assign node305 = (inp[5]) ? node307 : 3'b110;
									assign node307 = (inp[2]) ? node311 : node308;
										assign node308 = (inp[1]) ? 3'b010 : 3'b110;
										assign node311 = (inp[1]) ? 3'b110 : 3'b010;
							assign node314 = (inp[2]) ? node324 : node315;
								assign node315 = (inp[3]) ? 3'b100 : node316;
									assign node316 = (inp[8]) ? node320 : node317;
										assign node317 = (inp[1]) ? 3'b100 : 3'b000;
										assign node320 = (inp[4]) ? 3'b010 : 3'b110;
								assign node324 = (inp[4]) ? node334 : node325;
									assign node325 = (inp[5]) ? node329 : node326;
										assign node326 = (inp[8]) ? 3'b000 : 3'b100;
										assign node329 = (inp[1]) ? 3'b100 : node330;
											assign node330 = (inp[8]) ? 3'b100 : 3'b000;
									assign node334 = (inp[1]) ? 3'b000 : node335;
										assign node335 = (inp[8]) ? 3'b100 : 3'b000;
				assign node339 = (inp[0]) ? node395 : node340;
					assign node340 = (inp[10]) ? node352 : node341;
						assign node341 = (inp[1]) ? node343 : 3'b111;
							assign node343 = (inp[8]) ? 3'b111 : node344;
								assign node344 = (inp[11]) ? 3'b011 : node345;
									assign node345 = (inp[5]) ? node347 : 3'b111;
										assign node347 = (inp[3]) ? 3'b011 : 3'b111;
						assign node352 = (inp[11]) ? node372 : node353;
							assign node353 = (inp[4]) ? node361 : node354;
								assign node354 = (inp[1]) ? node356 : 3'b111;
									assign node356 = (inp[2]) ? 3'b011 : node357;
										assign node357 = (inp[8]) ? 3'b111 : 3'b011;
								assign node361 = (inp[1]) ? node365 : node362;
									assign node362 = (inp[8]) ? 3'b111 : 3'b011;
									assign node365 = (inp[2]) ? 3'b101 : node366;
										assign node366 = (inp[5]) ? 3'b011 : node367;
											assign node367 = (inp[8]) ? 3'b011 : 3'b101;
							assign node372 = (inp[1]) ? node382 : node373;
								assign node373 = (inp[8]) ? node379 : node374;
									assign node374 = (inp[4]) ? 3'b101 : node375;
										assign node375 = (inp[3]) ? 3'b001 : 3'b011;
									assign node379 = (inp[2]) ? 3'b011 : 3'b111;
								assign node382 = (inp[8]) ? node386 : node383;
									assign node383 = (inp[2]) ? 3'b001 : 3'b101;
									assign node386 = (inp[2]) ? 3'b101 : node387;
										assign node387 = (inp[3]) ? node389 : 3'b001;
											assign node389 = (inp[5]) ? 3'b101 : node390;
												assign node390 = (inp[4]) ? 3'b101 : 3'b001;
					assign node395 = (inp[10]) ? node449 : node396;
						assign node396 = (inp[1]) ? node420 : node397;
							assign node397 = (inp[2]) ? node407 : node398;
								assign node398 = (inp[11]) ? node402 : node399;
									assign node399 = (inp[8]) ? 3'b111 : 3'b011;
									assign node402 = (inp[8]) ? 3'b011 : node403;
										assign node403 = (inp[5]) ? 3'b101 : 3'b011;
								assign node407 = (inp[4]) ? node413 : node408;
									assign node408 = (inp[8]) ? 3'b011 : node409;
										assign node409 = (inp[5]) ? 3'b001 : 3'b011;
									assign node413 = (inp[5]) ? node415 : 3'b101;
										assign node415 = (inp[8]) ? node417 : 3'b101;
											assign node417 = (inp[11]) ? 3'b101 : 3'b011;
							assign node420 = (inp[4]) ? node432 : node421;
								assign node421 = (inp[8]) ? node423 : 3'b001;
									assign node423 = (inp[3]) ? 3'b101 : node424;
										assign node424 = (inp[11]) ? node428 : node425;
											assign node425 = (inp[2]) ? 3'b101 : 3'b011;
											assign node428 = (inp[2]) ? 3'b001 : 3'b101;
								assign node432 = (inp[8]) ? node442 : node433;
									assign node433 = (inp[2]) ? node437 : node434;
										assign node434 = (inp[11]) ? 3'b001 : 3'b101;
										assign node437 = (inp[3]) ? node439 : 3'b111;
											assign node439 = (inp[5]) ? 3'b110 : 3'b111;
									assign node442 = (inp[11]) ? node446 : node443;
										assign node443 = (inp[2]) ? 3'b101 : 3'b011;
										assign node446 = (inp[2]) ? 3'b001 : 3'b101;
						assign node449 = (inp[1]) ? node473 : node450;
							assign node450 = (inp[2]) ? node460 : node451;
								assign node451 = (inp[3]) ? 3'b001 : node452;
									assign node452 = (inp[5]) ? 3'b101 : node453;
										assign node453 = (inp[4]) ? node455 : 3'b101;
											assign node455 = (inp[8]) ? 3'b101 : 3'b001;
								assign node460 = (inp[4]) ? node468 : node461;
									assign node461 = (inp[5]) ? 3'b101 : node462;
										assign node462 = (inp[11]) ? 3'b010 : node463;
											assign node463 = (inp[8]) ? 3'b101 : 3'b001;
									assign node468 = (inp[11]) ? node470 : 3'b110;
										assign node470 = (inp[8]) ? 3'b110 : 3'b010;
							assign node473 = (inp[8]) ? node487 : node474;
								assign node474 = (inp[4]) ? node482 : node475;
									assign node475 = (inp[3]) ? 3'b010 : node476;
										assign node476 = (inp[11]) ? 3'b010 : node477;
											assign node477 = (inp[5]) ? 3'b110 : 3'b010;
									assign node482 = (inp[2]) ? 3'b100 : node483;
										assign node483 = (inp[11]) ? 3'b010 : 3'b110;
								assign node487 = (inp[5]) ? node489 : 3'b110;
									assign node489 = (inp[11]) ? 3'b111 : node490;
										assign node490 = (inp[2]) ? 3'b111 : node491;
											assign node491 = (inp[4]) ? 3'b001 : 3'b000;
			assign node496 = (inp[0]) ? node662 : node497;
				assign node497 = (inp[7]) ? node585 : node498;
					assign node498 = (inp[10]) ? node556 : node499;
						assign node499 = (inp[8]) ? node531 : node500;
							assign node500 = (inp[11]) ? node514 : node501;
								assign node501 = (inp[1]) ? node509 : node502;
									assign node502 = (inp[3]) ? node504 : 3'b110;
										assign node504 = (inp[4]) ? 3'b010 : node505;
											assign node505 = (inp[2]) ? 3'b010 : 3'b110;
									assign node509 = (inp[2]) ? 3'b100 : node510;
										assign node510 = (inp[4]) ? 3'b000 : 3'b010;
								assign node514 = (inp[4]) ? node522 : node515;
									assign node515 = (inp[5]) ? node517 : 3'b000;
										assign node517 = (inp[2]) ? 3'b100 : node518;
											assign node518 = (inp[3]) ? 3'b000 : 3'b100;
									assign node522 = (inp[5]) ? node524 : 3'b100;
										assign node524 = (inp[1]) ? 3'b000 : node525;
											assign node525 = (inp[2]) ? 3'b100 : node526;
												assign node526 = (inp[3]) ? 3'b100 : 3'b000;
							assign node531 = (inp[3]) ? node549 : node532;
								assign node532 = (inp[11]) ? node542 : node533;
									assign node533 = (inp[2]) ? node535 : 3'b110;
										assign node535 = (inp[1]) ? 3'b010 : node536;
											assign node536 = (inp[5]) ? 3'b110 : node537;
												assign node537 = (inp[4]) ? 3'b010 : 3'b110;
									assign node542 = (inp[4]) ? node544 : 3'b010;
										assign node544 = (inp[2]) ? 3'b100 : node545;
											assign node545 = (inp[1]) ? 3'b010 : 3'b110;
								assign node549 = (inp[11]) ? node553 : node550;
									assign node550 = (inp[1]) ? 3'b010 : 3'b001;
									assign node553 = (inp[1]) ? 3'b100 : 3'b010;
						assign node556 = (inp[1]) ? node576 : node557;
							assign node557 = (inp[3]) ? node567 : node558;
								assign node558 = (inp[11]) ? node562 : node559;
									assign node559 = (inp[2]) ? 3'b000 : 3'b010;
									assign node562 = (inp[2]) ? 3'b100 : node563;
										assign node563 = (inp[8]) ? 3'b100 : 3'b000;
								assign node567 = (inp[11]) ? node569 : 3'b100;
									assign node569 = (inp[8]) ? node573 : node570;
										assign node570 = (inp[2]) ? 3'b100 : 3'b000;
										assign node573 = (inp[2]) ? 3'b000 : 3'b100;
							assign node576 = (inp[8]) ? node578 : 3'b000;
								assign node578 = (inp[2]) ? 3'b000 : node579;
									assign node579 = (inp[3]) ? 3'b000 : node580;
										assign node580 = (inp[11]) ? 3'b000 : 3'b100;
					assign node585 = (inp[10]) ? node621 : node586;
						assign node586 = (inp[1]) ? node604 : node587;
							assign node587 = (inp[8]) ? node599 : node588;
								assign node588 = (inp[2]) ? node596 : node589;
									assign node589 = (inp[11]) ? node591 : 3'b101;
										assign node591 = (inp[3]) ? node593 : 3'b101;
											assign node593 = (inp[4]) ? 3'b101 : 3'b001;
									assign node596 = (inp[11]) ? 3'b110 : 3'b001;
								assign node599 = (inp[11]) ? 3'b001 : node600;
									assign node600 = (inp[3]) ? 3'b101 : 3'b011;
							assign node604 = (inp[11]) ? node612 : node605;
								assign node605 = (inp[8]) ? node607 : 3'b110;
									assign node607 = (inp[4]) ? node609 : 3'b101;
										assign node609 = (inp[3]) ? 3'b001 : 3'b101;
								assign node612 = (inp[2]) ? node616 : node613;
									assign node613 = (inp[8]) ? 3'b010 : 3'b110;
									assign node616 = (inp[4]) ? node618 : 3'b110;
										assign node618 = (inp[5]) ? 3'b110 : 3'b010;
						assign node621 = (inp[1]) ? node641 : node622;
							assign node622 = (inp[11]) ? node634 : node623;
								assign node623 = (inp[2]) ? node627 : node624;
									assign node624 = (inp[8]) ? 3'b001 : 3'b110;
									assign node627 = (inp[8]) ? node629 : 3'b010;
										assign node629 = (inp[5]) ? 3'b110 : node630;
											assign node630 = (inp[3]) ? 3'b110 : 3'b111;
								assign node634 = (inp[8]) ? node638 : node635;
									assign node635 = (inp[2]) ? 3'b100 : 3'b010;
									assign node638 = (inp[2]) ? 3'b010 : 3'b110;
							assign node641 = (inp[8]) ? node651 : node642;
								assign node642 = (inp[2]) ? node648 : node643;
									assign node643 = (inp[11]) ? 3'b100 : node644;
										assign node644 = (inp[3]) ? 3'b100 : 3'b010;
									assign node648 = (inp[11]) ? 3'b000 : 3'b100;
								assign node651 = (inp[11]) ? node659 : node652;
									assign node652 = (inp[4]) ? node654 : 3'b010;
										assign node654 = (inp[5]) ? 3'b010 : node655;
											assign node655 = (inp[2]) ? 3'b100 : 3'b010;
									assign node659 = (inp[3]) ? 3'b010 : 3'b100;
				assign node662 = (inp[10]) ? node728 : node663;
					assign node663 = (inp[7]) ? node687 : node664;
						assign node664 = (inp[8]) ? node666 : 3'b000;
							assign node666 = (inp[1]) ? 3'b000 : node667;
								assign node667 = (inp[11]) ? node679 : node668;
									assign node668 = (inp[2]) ? node674 : node669;
										assign node669 = (inp[5]) ? 3'b100 : node670;
											assign node670 = (inp[4]) ? 3'b100 : 3'b010;
										assign node674 = (inp[4]) ? node676 : 3'b100;
											assign node676 = (inp[3]) ? 3'b000 : 3'b100;
									assign node679 = (inp[4]) ? 3'b000 : node680;
										assign node680 = (inp[3]) ? 3'b010 : node681;
											assign node681 = (inp[2]) ? 3'b010 : 3'b100;
						assign node687 = (inp[11]) ? node705 : node688;
							assign node688 = (inp[8]) ? node696 : node689;
								assign node689 = (inp[5]) ? node693 : node690;
									assign node690 = (inp[2]) ? 3'b000 : 3'b100;
									assign node693 = (inp[2]) ? 3'b100 : 3'b010;
								assign node696 = (inp[4]) ? node698 : 3'b110;
									assign node698 = (inp[2]) ? node702 : node699;
										assign node699 = (inp[1]) ? 3'b010 : 3'b110;
										assign node702 = (inp[1]) ? 3'b110 : 3'b010;
							assign node705 = (inp[2]) ? node721 : node706;
								assign node706 = (inp[1]) ? node714 : node707;
									assign node707 = (inp[3]) ? node709 : 3'b010;
										assign node709 = (inp[4]) ? 3'b100 : node710;
											assign node710 = (inp[8]) ? 3'b110 : 3'b010;
									assign node714 = (inp[8]) ? node716 : 3'b000;
										assign node716 = (inp[5]) ? node718 : 3'b100;
											assign node718 = (inp[3]) ? 3'b100 : 3'b110;
								assign node721 = (inp[1]) ? node725 : node722;
									assign node722 = (inp[8]) ? 3'b100 : 3'b000;
									assign node725 = (inp[8]) ? 3'b000 : 3'b100;
					assign node728 = (inp[8]) ? node730 : 3'b000;
						assign node730 = (inp[7]) ? node732 : 3'b000;
							assign node732 = (inp[1]) ? 3'b000 : node733;
								assign node733 = (inp[4]) ? node735 : 3'b100;
									assign node735 = (inp[3]) ? node737 : 3'b010;
										assign node737 = (inp[11]) ? 3'b000 : 3'b100;

endmodule