module dtc_split33_bm59 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node7;
	wire [3-1:0] node9;
	wire [3-1:0] node11;
	wire [3-1:0] node14;
	wire [3-1:0] node15;
	wire [3-1:0] node17;
	wire [3-1:0] node18;
	wire [3-1:0] node22;
	wire [3-1:0] node23;
	wire [3-1:0] node26;
	wire [3-1:0] node30;
	wire [3-1:0] node31;
	wire [3-1:0] node32;
	wire [3-1:0] node34;
	wire [3-1:0] node35;
	wire [3-1:0] node39;
	wire [3-1:0] node40;
	wire [3-1:0] node41;
	wire [3-1:0] node42;
	wire [3-1:0] node47;
	wire [3-1:0] node50;
	wire [3-1:0] node51;
	wire [3-1:0] node53;
	wire [3-1:0] node54;
	wire [3-1:0] node56;
	wire [3-1:0] node57;
	wire [3-1:0] node62;
	wire [3-1:0] node63;
	wire [3-1:0] node65;
	wire [3-1:0] node70;
	wire [3-1:0] node71;
	wire [3-1:0] node72;
	wire [3-1:0] node73;
	wire [3-1:0] node74;
	wire [3-1:0] node75;
	wire [3-1:0] node78;
	wire [3-1:0] node79;
	wire [3-1:0] node83;
	wire [3-1:0] node84;
	wire [3-1:0] node88;
	wire [3-1:0] node89;
	wire [3-1:0] node90;
	wire [3-1:0] node91;
	wire [3-1:0] node96;
	wire [3-1:0] node97;
	wire [3-1:0] node98;
	wire [3-1:0] node99;
	wire [3-1:0] node100;
	wire [3-1:0] node105;
	wire [3-1:0] node106;
	wire [3-1:0] node111;
	wire [3-1:0] node112;
	wire [3-1:0] node113;
	wire [3-1:0] node114;
	wire [3-1:0] node117;
	wire [3-1:0] node118;
	wire [3-1:0] node120;
	wire [3-1:0] node123;
	wire [3-1:0] node126;
	wire [3-1:0] node127;
	wire [3-1:0] node130;
	wire [3-1:0] node131;
	wire [3-1:0] node132;
	wire [3-1:0] node134;
	wire [3-1:0] node138;
	wire [3-1:0] node139;
	wire [3-1:0] node144;
	wire [3-1:0] node145;
	wire [3-1:0] node146;
	wire [3-1:0] node147;
	wire [3-1:0] node148;
	wire [3-1:0] node149;
	wire [3-1:0] node151;
	wire [3-1:0] node153;
	wire [3-1:0] node156;
	wire [3-1:0] node159;
	wire [3-1:0] node160;
	wire [3-1:0] node163;
	wire [3-1:0] node165;
	wire [3-1:0] node168;
	wire [3-1:0] node169;
	wire [3-1:0] node170;
	wire [3-1:0] node173;
	wire [3-1:0] node175;
	wire [3-1:0] node178;
	wire [3-1:0] node179;
	wire [3-1:0] node182;
	wire [3-1:0] node185;
	wire [3-1:0] node186;
	wire [3-1:0] node187;
	wire [3-1:0] node188;
	wire [3-1:0] node190;
	wire [3-1:0] node193;
	wire [3-1:0] node194;
	wire [3-1:0] node198;
	wire [3-1:0] node199;
	wire [3-1:0] node202;
	wire [3-1:0] node203;
	wire [3-1:0] node207;
	wire [3-1:0] node208;
	wire [3-1:0] node209;
	wire [3-1:0] node210;
	wire [3-1:0] node213;
	wire [3-1:0] node218;
	wire [3-1:0] node219;
	wire [3-1:0] node220;
	wire [3-1:0] node221;
	wire [3-1:0] node223;
	wire [3-1:0] node225;
	wire [3-1:0] node228;
	wire [3-1:0] node230;
	wire [3-1:0] node233;
	wire [3-1:0] node234;
	wire [3-1:0] node238;
	wire [3-1:0] node239;
	wire [3-1:0] node241;
	wire [3-1:0] node242;
	wire [3-1:0] node243;
	wire [3-1:0] node244;
	wire [3-1:0] node251;
	wire [3-1:0] node252;
	wire [3-1:0] node253;
	wire [3-1:0] node254;
	wire [3-1:0] node255;
	wire [3-1:0] node257;
	wire [3-1:0] node258;
	wire [3-1:0] node261;
	wire [3-1:0] node265;
	wire [3-1:0] node266;
	wire [3-1:0] node267;
	wire [3-1:0] node268;
	wire [3-1:0] node269;
	wire [3-1:0] node270;
	wire [3-1:0] node275;
	wire [3-1:0] node276;
	wire [3-1:0] node279;
	wire [3-1:0] node282;
	wire [3-1:0] node283;
	wire [3-1:0] node284;
	wire [3-1:0] node286;
	wire [3-1:0] node289;
	wire [3-1:0] node292;
	wire [3-1:0] node293;
	wire [3-1:0] node296;
	wire [3-1:0] node299;
	wire [3-1:0] node301;
	wire [3-1:0] node302;
	wire [3-1:0] node304;
	wire [3-1:0] node307;
	wire [3-1:0] node309;
	wire [3-1:0] node311;
	wire [3-1:0] node315;
	wire [3-1:0] node316;
	wire [3-1:0] node317;
	wire [3-1:0] node318;
	wire [3-1:0] node319;
	wire [3-1:0] node320;
	wire [3-1:0] node321;
	wire [3-1:0] node324;
	wire [3-1:0] node325;
	wire [3-1:0] node326;
	wire [3-1:0] node331;
	wire [3-1:0] node333;
	wire [3-1:0] node336;
	wire [3-1:0] node337;
	wire [3-1:0] node339;
	wire [3-1:0] node342;
	wire [3-1:0] node344;
	wire [3-1:0] node347;
	wire [3-1:0] node348;
	wire [3-1:0] node349;
	wire [3-1:0] node350;
	wire [3-1:0] node354;
	wire [3-1:0] node357;
	wire [3-1:0] node358;
	wire [3-1:0] node362;
	wire [3-1:0] node364;
	wire [3-1:0] node365;
	wire [3-1:0] node366;
	wire [3-1:0] node368;
	wire [3-1:0] node369;
	wire [3-1:0] node373;
	wire [3-1:0] node375;
	wire [3-1:0] node379;
	wire [3-1:0] node380;
	wire [3-1:0] node381;
	wire [3-1:0] node382;
	wire [3-1:0] node384;
	wire [3-1:0] node385;
	wire [3-1:0] node389;
	wire [3-1:0] node390;
	wire [3-1:0] node391;
	wire [3-1:0] node393;
	wire [3-1:0] node396;
	wire [3-1:0] node399;
	wire [3-1:0] node400;
	wire [3-1:0] node402;
	wire [3-1:0] node405;
	wire [3-1:0] node408;
	wire [3-1:0] node409;
	wire [3-1:0] node411;
	wire [3-1:0] node414;
	wire [3-1:0] node416;
	wire [3-1:0] node417;
	wire [3-1:0] node421;
	wire [3-1:0] node422;
	wire [3-1:0] node423;
	wire [3-1:0] node424;
	wire [3-1:0] node425;
	wire [3-1:0] node427;
	wire [3-1:0] node428;
	wire [3-1:0] node431;
	wire [3-1:0] node435;
	wire [3-1:0] node436;
	wire [3-1:0] node437;
	wire [3-1:0] node438;
	wire [3-1:0] node444;
	wire [3-1:0] node445;
	wire [3-1:0] node447;
	wire [3-1:0] node448;
	wire [3-1:0] node453;
	wire [3-1:0] node454;
	wire [3-1:0] node455;
	wire [3-1:0] node457;
	wire [3-1:0] node462;
	wire [3-1:0] node463;
	wire [3-1:0] node464;
	wire [3-1:0] node465;
	wire [3-1:0] node466;
	wire [3-1:0] node467;
	wire [3-1:0] node468;
	wire [3-1:0] node469;
	wire [3-1:0] node471;
	wire [3-1:0] node474;
	wire [3-1:0] node475;
	wire [3-1:0] node477;
	wire [3-1:0] node480;
	wire [3-1:0] node483;
	wire [3-1:0] node484;
	wire [3-1:0] node487;
	wire [3-1:0] node490;
	wire [3-1:0] node491;
	wire [3-1:0] node492;
	wire [3-1:0] node493;
	wire [3-1:0] node494;
	wire [3-1:0] node499;
	wire [3-1:0] node502;
	wire [3-1:0] node503;
	wire [3-1:0] node505;
	wire [3-1:0] node508;
	wire [3-1:0] node510;
	wire [3-1:0] node513;
	wire [3-1:0] node515;
	wire [3-1:0] node516;
	wire [3-1:0] node517;
	wire [3-1:0] node521;
	wire [3-1:0] node522;
	wire [3-1:0] node523;
	wire [3-1:0] node525;
	wire [3-1:0] node529;
	wire [3-1:0] node530;
	wire [3-1:0] node535;
	wire [3-1:0] node536;
	wire [3-1:0] node537;
	wire [3-1:0] node538;
	wire [3-1:0] node539;
	wire [3-1:0] node540;
	wire [3-1:0] node542;
	wire [3-1:0] node543;
	wire [3-1:0] node547;
	wire [3-1:0] node548;
	wire [3-1:0] node552;
	wire [3-1:0] node553;
	wire [3-1:0] node554;
	wire [3-1:0] node555;
	wire [3-1:0] node559;
	wire [3-1:0] node562;
	wire [3-1:0] node564;
	wire [3-1:0] node567;
	wire [3-1:0] node569;
	wire [3-1:0] node570;
	wire [3-1:0] node572;
	wire [3-1:0] node574;
	wire [3-1:0] node577;
	wire [3-1:0] node578;
	wire [3-1:0] node582;
	wire [3-1:0] node583;
	wire [3-1:0] node584;
	wire [3-1:0] node585;
	wire [3-1:0] node586;
	wire [3-1:0] node590;
	wire [3-1:0] node591;
	wire [3-1:0] node594;
	wire [3-1:0] node596;
	wire [3-1:0] node599;
	wire [3-1:0] node600;
	wire [3-1:0] node601;
	wire [3-1:0] node602;
	wire [3-1:0] node607;
	wire [3-1:0] node609;
	wire [3-1:0] node611;
	wire [3-1:0] node615;
	wire [3-1:0] node616;
	wire [3-1:0] node617;
	wire [3-1:0] node618;
	wire [3-1:0] node619;
	wire [3-1:0] node621;
	wire [3-1:0] node624;
	wire [3-1:0] node625;
	wire [3-1:0] node627;
	wire [3-1:0] node631;
	wire [3-1:0] node632;
	wire [3-1:0] node633;
	wire [3-1:0] node637;
	wire [3-1:0] node638;
	wire [3-1:0] node642;
	wire [3-1:0] node643;
	wire [3-1:0] node646;
	wire [3-1:0] node647;
	wire [3-1:0] node650;
	wire [3-1:0] node651;
	wire [3-1:0] node653;
	wire [3-1:0] node656;
	wire [3-1:0] node658;
	wire [3-1:0] node661;
	wire [3-1:0] node662;
	wire [3-1:0] node663;
	wire [3-1:0] node664;
	wire [3-1:0] node665;
	wire [3-1:0] node667;
	wire [3-1:0] node672;
	wire [3-1:0] node674;
	wire [3-1:0] node675;
	wire [3-1:0] node679;
	wire [3-1:0] node681;
	wire [3-1:0] node682;
	wire [3-1:0] node684;
	wire [3-1:0] node685;
	wire [3-1:0] node690;
	wire [3-1:0] node691;
	wire [3-1:0] node692;
	wire [3-1:0] node693;
	wire [3-1:0] node695;
	wire [3-1:0] node697;
	wire [3-1:0] node698;
	wire [3-1:0] node699;
	wire [3-1:0] node701;
	wire [3-1:0] node706;
	wire [3-1:0] node707;
	wire [3-1:0] node708;
	wire [3-1:0] node709;
	wire [3-1:0] node710;
	wire [3-1:0] node713;
	wire [3-1:0] node714;
	wire [3-1:0] node718;
	wire [3-1:0] node719;
	wire [3-1:0] node720;
	wire [3-1:0] node724;
	wire [3-1:0] node727;
	wire [3-1:0] node728;
	wire [3-1:0] node729;
	wire [3-1:0] node730;
	wire [3-1:0] node735;
	wire [3-1:0] node737;
	wire [3-1:0] node740;
	wire [3-1:0] node742;
	wire [3-1:0] node743;
	wire [3-1:0] node744;
	wire [3-1:0] node747;
	wire [3-1:0] node750;
	wire [3-1:0] node753;
	wire [3-1:0] node754;
	wire [3-1:0] node755;
	wire [3-1:0] node756;
	wire [3-1:0] node758;
	wire [3-1:0] node759;
	wire [3-1:0] node762;
	wire [3-1:0] node763;
	wire [3-1:0] node767;
	wire [3-1:0] node768;
	wire [3-1:0] node770;
	wire [3-1:0] node773;
	wire [3-1:0] node774;
	wire [3-1:0] node775;
	wire [3-1:0] node778;
	wire [3-1:0] node782;
	wire [3-1:0] node783;
	wire [3-1:0] node785;
	wire [3-1:0] node786;
	wire [3-1:0] node787;
	wire [3-1:0] node791;
	wire [3-1:0] node792;
	wire [3-1:0] node796;
	wire [3-1:0] node797;
	wire [3-1:0] node801;
	wire [3-1:0] node802;
	wire [3-1:0] node803;
	wire [3-1:0] node804;
	wire [3-1:0] node807;
	wire [3-1:0] node808;
	wire [3-1:0] node809;
	wire [3-1:0] node814;
	wire [3-1:0] node815;
	wire [3-1:0] node817;
	wire [3-1:0] node818;
	wire [3-1:0] node822;
	wire [3-1:0] node823;
	wire [3-1:0] node826;
	wire [3-1:0] node829;
	wire [3-1:0] node831;
	wire [3-1:0] node832;
	wire [3-1:0] node834;
	wire [3-1:0] node838;
	wire [3-1:0] node840;
	wire [3-1:0] node841;
	wire [3-1:0] node842;
	wire [3-1:0] node844;
	wire [3-1:0] node846;
	wire [3-1:0] node847;
	wire [3-1:0] node852;
	wire [3-1:0] node853;
	wire [3-1:0] node854;
	wire [3-1:0] node855;
	wire [3-1:0] node856;
	wire [3-1:0] node858;
	wire [3-1:0] node859;
	wire [3-1:0] node863;
	wire [3-1:0] node866;
	wire [3-1:0] node867;
	wire [3-1:0] node868;
	wire [3-1:0] node873;
	wire [3-1:0] node874;
	wire [3-1:0] node875;
	wire [3-1:0] node880;
	wire [3-1:0] node881;
	wire [3-1:0] node882;

	assign outp = (inp[10]) ? node462 : node1;
		assign node1 = (inp[9]) ? node251 : node2;
			assign node2 = (inp[2]) ? node70 : node3;
				assign node3 = (inp[0]) ? 3'b110 : node4;
					assign node4 = (inp[1]) ? node30 : node5;
						assign node5 = (inp[3]) ? 3'b111 : node6;
							assign node6 = (inp[7]) ? node14 : node7;
								assign node7 = (inp[4]) ? node9 : 3'b111;
									assign node9 = (inp[5]) ? node11 : 3'b000;
										assign node11 = (inp[6]) ? 3'b000 : 3'b010;
								assign node14 = (inp[8]) ? node22 : node15;
									assign node15 = (inp[6]) ? node17 : 3'b110;
										assign node17 = (inp[5]) ? 3'b100 : node18;
											assign node18 = (inp[4]) ? 3'b110 : 3'b100;
									assign node22 = (inp[6]) ? node26 : node23;
										assign node23 = (inp[5]) ? 3'b110 : 3'b100;
										assign node26 = (inp[5]) ? 3'b000 : 3'b010;
						assign node30 = (inp[5]) ? node50 : node31;
							assign node31 = (inp[6]) ? node39 : node32;
								assign node32 = (inp[7]) ? node34 : 3'b000;
									assign node34 = (inp[4]) ? 3'b100 : node35;
										assign node35 = (inp[8]) ? 3'b000 : 3'b100;
								assign node39 = (inp[11]) ? node47 : node40;
									assign node40 = (inp[8]) ? 3'b110 : node41;
										assign node41 = (inp[4]) ? 3'b010 : node42;
											assign node42 = (inp[7]) ? 3'b010 : 3'b111;
									assign node47 = (inp[7]) ? 3'b100 : 3'b000;
							assign node50 = (inp[7]) ? node62 : node51;
								assign node51 = (inp[6]) ? node53 : 3'b010;
									assign node53 = (inp[4]) ? 3'b000 : node54;
										assign node54 = (inp[8]) ? node56 : 3'b010;
											assign node56 = (inp[3]) ? 3'b111 : node57;
												assign node57 = (inp[11]) ? 3'b110 : 3'b100;
								assign node62 = (inp[4]) ? 3'b110 : node63;
									assign node63 = (inp[3]) ? node65 : 3'b000;
										assign node65 = (inp[8]) ? 3'b010 : 3'b110;
				assign node70 = (inp[1]) ? node144 : node71;
					assign node71 = (inp[0]) ? node111 : node72;
						assign node72 = (inp[11]) ? node88 : node73;
							assign node73 = (inp[4]) ? node83 : node74;
								assign node74 = (inp[5]) ? node78 : node75;
									assign node75 = (inp[6]) ? 3'b100 : 3'b000;
									assign node78 = (inp[6]) ? 3'b000 : node79;
										assign node79 = (inp[7]) ? 3'b000 : 3'b010;
								assign node83 = (inp[5]) ? 3'b100 : node84;
									assign node84 = (inp[8]) ? 3'b000 : 3'b010;
							assign node88 = (inp[4]) ? node96 : node89;
								assign node89 = (inp[5]) ? 3'b010 : node90;
									assign node90 = (inp[3]) ? 3'b000 : node91;
										assign node91 = (inp[8]) ? 3'b110 : 3'b010;
								assign node96 = (inp[5]) ? 3'b110 : node97;
									assign node97 = (inp[8]) ? node105 : node98;
										assign node98 = (inp[6]) ? 3'b000 : node99;
											assign node99 = (inp[3]) ? 3'b110 : node100;
												assign node100 = (inp[7]) ? 3'b100 : 3'b110;
										assign node105 = (inp[3]) ? 3'b010 : node106;
											assign node106 = (inp[7]) ? 3'b000 : 3'b010;
						assign node111 = (inp[3]) ? 3'b110 : node112;
							assign node112 = (inp[5]) ? node126 : node113;
								assign node113 = (inp[6]) ? node117 : node114;
									assign node114 = (inp[7]) ? 3'b100 : 3'b000;
									assign node117 = (inp[11]) ? node123 : node118;
										assign node118 = (inp[8]) ? node120 : 3'b110;
											assign node120 = (inp[7]) ? 3'b010 : 3'b110;
										assign node123 = (inp[7]) ? 3'b100 : 3'b110;
								assign node126 = (inp[11]) ? node130 : node127;
									assign node127 = (inp[6]) ? 3'b100 : 3'b110;
									assign node130 = (inp[6]) ? node138 : node131;
										assign node131 = (inp[4]) ? 3'b110 : node132;
											assign node132 = (inp[8]) ? node134 : 3'b110;
												assign node134 = (inp[7]) ? 3'b010 : 3'b110;
										assign node138 = (inp[4]) ? 3'b010 : node139;
											assign node139 = (inp[8]) ? 3'b010 : 3'b110;
					assign node144 = (inp[7]) ? node218 : node145;
						assign node145 = (inp[11]) ? node185 : node146;
							assign node146 = (inp[0]) ? node168 : node147;
								assign node147 = (inp[4]) ? node159 : node148;
									assign node148 = (inp[8]) ? node156 : node149;
										assign node149 = (inp[5]) ? node151 : 3'b010;
											assign node151 = (inp[3]) ? node153 : 3'b110;
												assign node153 = (inp[6]) ? 3'b010 : 3'b100;
										assign node156 = (inp[6]) ? 3'b100 : 3'b110;
									assign node159 = (inp[3]) ? node163 : node160;
										assign node160 = (inp[5]) ? 3'b000 : 3'b010;
										assign node163 = (inp[8]) ? node165 : 3'b010;
											assign node165 = (inp[5]) ? 3'b010 : 3'b110;
								assign node168 = (inp[5]) ? node178 : node169;
									assign node169 = (inp[6]) ? node173 : node170;
										assign node170 = (inp[8]) ? 3'b100 : 3'b000;
										assign node173 = (inp[4]) ? node175 : 3'b110;
											assign node175 = (inp[8]) ? 3'b000 : 3'b100;
									assign node178 = (inp[8]) ? node182 : node179;
										assign node179 = (inp[4]) ? 3'b010 : 3'b000;
										assign node182 = (inp[4]) ? 3'b100 : 3'b000;
							assign node185 = (inp[5]) ? node207 : node186;
								assign node186 = (inp[8]) ? node198 : node187;
									assign node187 = (inp[0]) ? node193 : node188;
										assign node188 = (inp[3]) ? node190 : 3'b010;
											assign node190 = (inp[4]) ? 3'b010 : 3'b000;
										assign node193 = (inp[4]) ? 3'b000 : node194;
											assign node194 = (inp[3]) ? 3'b000 : 3'b010;
									assign node198 = (inp[6]) ? node202 : node199;
										assign node199 = (inp[3]) ? 3'b000 : 3'b100;
										assign node202 = (inp[4]) ? 3'b010 : node203;
											assign node203 = (inp[0]) ? 3'b100 : 3'b010;
								assign node207 = (inp[4]) ? 3'b010 : node208;
									assign node208 = (inp[0]) ? 3'b010 : node209;
										assign node209 = (inp[8]) ? node213 : node210;
											assign node210 = (inp[6]) ? 3'b110 : 3'b010;
											assign node213 = (inp[3]) ? 3'b010 : 3'b110;
						assign node218 = (inp[4]) ? node238 : node219;
							assign node219 = (inp[5]) ? node233 : node220;
								assign node220 = (inp[3]) ? node228 : node221;
									assign node221 = (inp[8]) ? node223 : 3'b010;
										assign node223 = (inp[11]) ? node225 : 3'b010;
											assign node225 = (inp[0]) ? 3'b010 : 3'b000;
									assign node228 = (inp[0]) ? node230 : 3'b000;
										assign node230 = (inp[11]) ? 3'b000 : 3'b010;
								assign node233 = (inp[11]) ? 3'b010 : node234;
									assign node234 = (inp[8]) ? 3'b010 : 3'b000;
							assign node238 = (inp[11]) ? 3'b000 : node239;
								assign node239 = (inp[3]) ? node241 : 3'b000;
									assign node241 = (inp[0]) ? 3'b010 : node242;
										assign node242 = (inp[8]) ? 3'b000 : node243;
											assign node243 = (inp[6]) ? 3'b000 : node244;
												assign node244 = (inp[5]) ? 3'b000 : 3'b010;
			assign node251 = (inp[2]) ? node315 : node252;
				assign node252 = (inp[0]) ? 3'b010 : node253;
					assign node253 = (inp[1]) ? node265 : node254;
						assign node254 = (inp[3]) ? 3'b011 : node255;
							assign node255 = (inp[7]) ? node257 : 3'b011;
								assign node257 = (inp[6]) ? node261 : node258;
									assign node258 = (inp[5]) ? 3'b010 : 3'b000;
									assign node261 = (inp[4]) ? 3'b010 : 3'b011;
						assign node265 = (inp[3]) ? node299 : node266;
							assign node266 = (inp[5]) ? node282 : node267;
								assign node267 = (inp[6]) ? node275 : node268;
									assign node268 = (inp[11]) ? 3'b000 : node269;
										assign node269 = (inp[4]) ? 3'b000 : node270;
											assign node270 = (inp[8]) ? 3'b100 : 3'b000;
									assign node275 = (inp[11]) ? node279 : node276;
										assign node276 = (inp[8]) ? 3'b010 : 3'b110;
										assign node279 = (inp[7]) ? 3'b000 : 3'b100;
								assign node282 = (inp[6]) ? node292 : node283;
									assign node283 = (inp[11]) ? node289 : node284;
										assign node284 = (inp[7]) ? node286 : 3'b010;
											assign node286 = (inp[4]) ? 3'b010 : 3'b110;
										assign node289 = (inp[7]) ? 3'b010 : 3'b110;
									assign node292 = (inp[11]) ? node296 : node293;
										assign node293 = (inp[4]) ? 3'b000 : 3'b100;
										assign node296 = (inp[7]) ? 3'b010 : 3'b110;
							assign node299 = (inp[7]) ? node301 : 3'b011;
								assign node301 = (inp[8]) ? node307 : node302;
									assign node302 = (inp[4]) ? node304 : 3'b000;
										assign node304 = (inp[5]) ? 3'b010 : 3'b000;
									assign node307 = (inp[4]) ? node309 : 3'b011;
										assign node309 = (inp[11]) ? node311 : 3'b011;
											assign node311 = (inp[6]) ? 3'b000 : 3'b010;
				assign node315 = (inp[1]) ? node379 : node316;
					assign node316 = (inp[0]) ? node362 : node317;
						assign node317 = (inp[5]) ? node347 : node318;
							assign node318 = (inp[8]) ? node336 : node319;
								assign node319 = (inp[6]) ? node331 : node320;
									assign node320 = (inp[4]) ? node324 : node321;
										assign node321 = (inp[7]) ? 3'b000 : 3'b100;
										assign node324 = (inp[3]) ? 3'b010 : node325;
											assign node325 = (inp[7]) ? 3'b000 : node326;
												assign node326 = (inp[11]) ? 3'b010 : 3'b000;
									assign node331 = (inp[4]) ? node333 : 3'b010;
										assign node333 = (inp[11]) ? 3'b010 : 3'b000;
								assign node336 = (inp[4]) ? node342 : node337;
									assign node337 = (inp[7]) ? node339 : 3'b000;
										assign node339 = (inp[3]) ? 3'b100 : 3'b010;
									assign node342 = (inp[7]) ? node344 : 3'b100;
										assign node344 = (inp[6]) ? 3'b100 : 3'b000;
							assign node347 = (inp[8]) ? node357 : node348;
								assign node348 = (inp[7]) ? node354 : node349;
									assign node349 = (inp[11]) ? 3'b110 : node350;
										assign node350 = (inp[6]) ? 3'b100 : 3'b110;
									assign node354 = (inp[4]) ? 3'b000 : 3'b010;
								assign node357 = (inp[7]) ? 3'b110 : node358;
									assign node358 = (inp[4]) ? 3'b110 : 3'b010;
						assign node362 = (inp[7]) ? node364 : 3'b010;
							assign node364 = (inp[3]) ? 3'b010 : node365;
								assign node365 = (inp[5]) ? node373 : node366;
									assign node366 = (inp[4]) ? node368 : 3'b010;
										assign node368 = (inp[11]) ? 3'b000 : node369;
											assign node369 = (inp[8]) ? 3'b000 : 3'b010;
									assign node373 = (inp[6]) ? node375 : 3'b010;
										assign node375 = (inp[4]) ? 3'b010 : 3'b000;
					assign node379 = (inp[7]) ? node421 : node380;
						assign node380 = (inp[5]) ? node408 : node381;
							assign node381 = (inp[8]) ? node389 : node382;
								assign node382 = (inp[4]) ? node384 : 3'b100;
									assign node384 = (inp[0]) ? 3'b010 : node385;
										assign node385 = (inp[3]) ? 3'b100 : 3'b000;
								assign node389 = (inp[11]) ? node399 : node390;
									assign node390 = (inp[3]) ? node396 : node391;
										assign node391 = (inp[0]) ? node393 : 3'b010;
											assign node393 = (inp[6]) ? 3'b010 : 3'b000;
										assign node396 = (inp[0]) ? 3'b010 : 3'b000;
									assign node399 = (inp[3]) ? node405 : node400;
										assign node400 = (inp[4]) ? node402 : 3'b000;
											assign node402 = (inp[0]) ? 3'b100 : 3'b000;
										assign node405 = (inp[4]) ? 3'b000 : 3'b010;
							assign node408 = (inp[11]) ? node414 : node409;
								assign node409 = (inp[6]) ? node411 : 3'b010;
									assign node411 = (inp[4]) ? 3'b000 : 3'b100;
								assign node414 = (inp[0]) ? node416 : 3'b010;
									assign node416 = (inp[8]) ? 3'b010 : node417;
										assign node417 = (inp[3]) ? 3'b010 : 3'b110;
						assign node421 = (inp[4]) ? node453 : node422;
							assign node422 = (inp[11]) ? node444 : node423;
								assign node423 = (inp[0]) ? node435 : node424;
									assign node424 = (inp[5]) ? 3'b000 : node425;
										assign node425 = (inp[8]) ? node427 : 3'b000;
											assign node427 = (inp[6]) ? node431 : node428;
												assign node428 = (inp[3]) ? 3'b000 : 3'b010;
												assign node431 = (inp[3]) ? 3'b010 : 3'b000;
									assign node435 = (inp[5]) ? 3'b010 : node436;
										assign node436 = (inp[8]) ? 3'b010 : node437;
											assign node437 = (inp[3]) ? 3'b000 : node438;
												assign node438 = (inp[6]) ? 3'b000 : 3'b010;
								assign node444 = (inp[5]) ? 3'b010 : node445;
									assign node445 = (inp[8]) ? node447 : 3'b000;
										assign node447 = (inp[3]) ? 3'b010 : node448;
											assign node448 = (inp[0]) ? 3'b000 : 3'b010;
							assign node453 = (inp[5]) ? 3'b000 : node454;
								assign node454 = (inp[11]) ? 3'b000 : node455;
									assign node455 = (inp[6]) ? node457 : 3'b000;
										assign node457 = (inp[0]) ? 3'b000 : 3'b010;
		assign node462 = (inp[9]) ? node690 : node463;
			assign node463 = (inp[2]) ? node535 : node464;
				assign node464 = (inp[0]) ? 3'b100 : node465;
					assign node465 = (inp[3]) ? node513 : node466;
						assign node466 = (inp[5]) ? node490 : node467;
							assign node467 = (inp[7]) ? node483 : node468;
								assign node468 = (inp[4]) ? node474 : node469;
									assign node469 = (inp[1]) ? node471 : 3'b101;
										assign node471 = (inp[6]) ? 3'b100 : 3'b110;
									assign node474 = (inp[8]) ? node480 : node475;
										assign node475 = (inp[6]) ? node477 : 3'b010;
											assign node477 = (inp[11]) ? 3'b010 : 3'b000;
										assign node480 = (inp[1]) ? 3'b110 : 3'b101;
								assign node483 = (inp[8]) ? node487 : node484;
									assign node484 = (inp[4]) ? 3'b110 : 3'b010;
									assign node487 = (inp[11]) ? 3'b010 : 3'b000;
							assign node490 = (inp[11]) ? node502 : node491;
								assign node491 = (inp[7]) ? node499 : node492;
									assign node492 = (inp[6]) ? 3'b101 : node493;
										assign node493 = (inp[4]) ? 3'b000 : node494;
											assign node494 = (inp[1]) ? 3'b100 : 3'b101;
									assign node499 = (inp[6]) ? 3'b010 : 3'b000;
								assign node502 = (inp[7]) ? node508 : node503;
									assign node503 = (inp[1]) ? node505 : 3'b000;
										assign node505 = (inp[8]) ? 3'b100 : 3'b000;
									assign node508 = (inp[8]) ? node510 : 3'b100;
										assign node510 = (inp[4]) ? 3'b100 : 3'b000;
						assign node513 = (inp[1]) ? node515 : 3'b101;
							assign node515 = (inp[7]) ? node521 : node516;
								assign node516 = (inp[8]) ? 3'b101 : node517;
									assign node517 = (inp[11]) ? 3'b000 : 3'b010;
								assign node521 = (inp[8]) ? node529 : node522;
									assign node522 = (inp[11]) ? 3'b100 : node523;
										assign node523 = (inp[6]) ? node525 : 3'b100;
											assign node525 = (inp[5]) ? 3'b110 : 3'b100;
									assign node529 = (inp[6]) ? 3'b010 : node530;
										assign node530 = (inp[4]) ? 3'b100 : 3'b000;
				assign node535 = (inp[1]) ? node615 : node536;
					assign node536 = (inp[0]) ? node582 : node537;
						assign node537 = (inp[11]) ? node567 : node538;
							assign node538 = (inp[6]) ? node552 : node539;
								assign node539 = (inp[5]) ? node547 : node540;
									assign node540 = (inp[3]) ? node542 : 3'b000;
										assign node542 = (inp[7]) ? 3'b010 : node543;
											assign node543 = (inp[4]) ? 3'b010 : 3'b110;
									assign node547 = (inp[3]) ? 3'b000 : node548;
										assign node548 = (inp[8]) ? 3'b010 : 3'b110;
								assign node552 = (inp[8]) ? node562 : node553;
									assign node553 = (inp[5]) ? node559 : node554;
										assign node554 = (inp[3]) ? 3'b100 : node555;
											assign node555 = (inp[7]) ? 3'b110 : 3'b010;
										assign node559 = (inp[7]) ? 3'b100 : 3'b110;
									assign node562 = (inp[7]) ? node564 : 3'b100;
										assign node564 = (inp[4]) ? 3'b010 : 3'b000;
							assign node567 = (inp[4]) ? node569 : 3'b000;
								assign node569 = (inp[5]) ? node577 : node570;
									assign node570 = (inp[7]) ? node572 : 3'b100;
										assign node572 = (inp[3]) ? node574 : 3'b010;
											assign node574 = (inp[8]) ? 3'b000 : 3'b100;
									assign node577 = (inp[7]) ? 3'b100 : node578;
										assign node578 = (inp[3]) ? 3'b000 : 3'b100;
						assign node582 = (inp[3]) ? 3'b100 : node583;
							assign node583 = (inp[6]) ? node599 : node584;
								assign node584 = (inp[5]) ? node590 : node585;
									assign node585 = (inp[7]) ? 3'b010 : node586;
										assign node586 = (inp[11]) ? 3'b100 : 3'b010;
									assign node590 = (inp[8]) ? node594 : node591;
										assign node591 = (inp[7]) ? 3'b100 : 3'b000;
										assign node594 = (inp[7]) ? node596 : 3'b100;
											assign node596 = (inp[4]) ? 3'b100 : 3'b000;
								assign node599 = (inp[11]) ? node607 : node600;
									assign node600 = (inp[5]) ? 3'b010 : node601;
										assign node601 = (inp[8]) ? 3'b000 : node602;
											assign node602 = (inp[4]) ? 3'b100 : 3'b000;
									assign node607 = (inp[5]) ? node609 : 3'b010;
										assign node609 = (inp[7]) ? node611 : 3'b000;
											assign node611 = (inp[4]) ? 3'b100 : 3'b000;
					assign node615 = (inp[7]) ? node661 : node616;
						assign node616 = (inp[4]) ? node642 : node617;
							assign node617 = (inp[3]) ? node631 : node618;
								assign node618 = (inp[0]) ? node624 : node619;
									assign node619 = (inp[5]) ? node621 : 3'b000;
										assign node621 = (inp[8]) ? 3'b000 : 3'b100;
									assign node624 = (inp[8]) ? 3'b110 : node625;
										assign node625 = (inp[6]) ? node627 : 3'b010;
											assign node627 = (inp[11]) ? 3'b000 : 3'b100;
								assign node631 = (inp[0]) ? node637 : node632;
									assign node632 = (inp[5]) ? 3'b000 : node633;
										assign node633 = (inp[11]) ? 3'b100 : 3'b110;
									assign node637 = (inp[8]) ? 3'b100 : node638;
										assign node638 = (inp[5]) ? 3'b000 : 3'b100;
							assign node642 = (inp[3]) ? node646 : node643;
								assign node643 = (inp[11]) ? 3'b000 : 3'b010;
								assign node646 = (inp[8]) ? node650 : node647;
									assign node647 = (inp[11]) ? 3'b010 : 3'b000;
									assign node650 = (inp[5]) ? node656 : node651;
										assign node651 = (inp[11]) ? node653 : 3'b100;
											assign node653 = (inp[0]) ? 3'b100 : 3'b000;
										assign node656 = (inp[6]) ? node658 : 3'b000;
											assign node658 = (inp[11]) ? 3'b000 : 3'b100;
						assign node661 = (inp[5]) ? node679 : node662;
							assign node662 = (inp[3]) ? node672 : node663;
								assign node663 = (inp[0]) ? 3'b000 : node664;
									assign node664 = (inp[11]) ? 3'b010 : node665;
										assign node665 = (inp[6]) ? node667 : 3'b000;
											assign node667 = (inp[4]) ? 3'b010 : 3'b000;
								assign node672 = (inp[4]) ? node674 : 3'b010;
									assign node674 = (inp[0]) ? 3'b000 : node675;
										assign node675 = (inp[11]) ? 3'b000 : 3'b010;
							assign node679 = (inp[6]) ? node681 : 3'b000;
								assign node681 = (inp[4]) ? 3'b000 : node682;
									assign node682 = (inp[0]) ? node684 : 3'b000;
										assign node684 = (inp[3]) ? 3'b010 : node685;
											assign node685 = (inp[8]) ? 3'b000 : 3'b010;
			assign node690 = (inp[0]) ? node838 : node691;
				assign node691 = (inp[2]) ? node753 : node692;
					assign node692 = (inp[1]) ? node706 : node693;
						assign node693 = (inp[4]) ? node695 : 3'b001;
							assign node695 = (inp[7]) ? node697 : 3'b001;
								assign node697 = (inp[3]) ? 3'b001 : node698;
									assign node698 = (inp[11]) ? 3'b010 : node699;
										assign node699 = (inp[5]) ? node701 : 3'b000;
											assign node701 = (inp[6]) ? 3'b001 : 3'b000;
						assign node706 = (inp[3]) ? node740 : node707;
							assign node707 = (inp[5]) ? node727 : node708;
								assign node708 = (inp[11]) ? node718 : node709;
									assign node709 = (inp[6]) ? node713 : node710;
										assign node710 = (inp[7]) ? 3'b110 : 3'b010;
										assign node713 = (inp[8]) ? 3'b100 : node714;
											assign node714 = (inp[7]) ? 3'b000 : 3'b100;
									assign node718 = (inp[8]) ? node724 : node719;
										assign node719 = (inp[7]) ? 3'b010 : node720;
											assign node720 = (inp[6]) ? 3'b110 : 3'b010;
										assign node724 = (inp[7]) ? 3'b110 : 3'b010;
								assign node727 = (inp[6]) ? node735 : node728;
									assign node728 = (inp[11]) ? 3'b100 : node729;
										assign node729 = (inp[8]) ? 3'b000 : node730;
											assign node730 = (inp[7]) ? 3'b000 : 3'b100;
									assign node735 = (inp[11]) ? node737 : 3'b110;
										assign node737 = (inp[7]) ? 3'b000 : 3'b100;
							assign node740 = (inp[7]) ? node742 : 3'b001;
								assign node742 = (inp[8]) ? node750 : node743;
									assign node743 = (inp[6]) ? node747 : node744;
										assign node744 = (inp[5]) ? 3'b000 : 3'b010;
										assign node747 = (inp[4]) ? 3'b000 : 3'b001;
									assign node750 = (inp[11]) ? 3'b000 : 3'b001;
					assign node753 = (inp[1]) ? node801 : node754;
						assign node754 = (inp[7]) ? node782 : node755;
							assign node755 = (inp[4]) ? node767 : node756;
								assign node756 = (inp[8]) ? node758 : 3'b010;
									assign node758 = (inp[5]) ? node762 : node759;
										assign node759 = (inp[11]) ? 3'b010 : 3'b000;
										assign node762 = (inp[11]) ? 3'b000 : node763;
											assign node763 = (inp[6]) ? 3'b010 : 3'b000;
								assign node767 = (inp[3]) ? node773 : node768;
									assign node768 = (inp[5]) ? node770 : 3'b100;
										assign node770 = (inp[11]) ? 3'b000 : 3'b010;
									assign node773 = (inp[11]) ? 3'b100 : node774;
										assign node774 = (inp[5]) ? node778 : node775;
											assign node775 = (inp[6]) ? 3'b100 : 3'b110;
											assign node778 = (inp[6]) ? 3'b110 : 3'b100;
							assign node782 = (inp[11]) ? node796 : node783;
								assign node783 = (inp[6]) ? node785 : 3'b110;
									assign node785 = (inp[8]) ? node791 : node786;
										assign node786 = (inp[5]) ? 3'b010 : node787;
											assign node787 = (inp[4]) ? 3'b000 : 3'b010;
										assign node791 = (inp[4]) ? 3'b110 : node792;
											assign node792 = (inp[3]) ? 3'b110 : 3'b010;
								assign node796 = (inp[3]) ? 3'b110 : node797;
									assign node797 = (inp[4]) ? 3'b000 : 3'b100;
						assign node801 = (inp[7]) ? node829 : node802;
							assign node802 = (inp[6]) ? node814 : node803;
								assign node803 = (inp[8]) ? node807 : node804;
									assign node804 = (inp[5]) ? 3'b000 : 3'b100;
									assign node807 = (inp[5]) ? 3'b000 : node808;
										assign node808 = (inp[3]) ? 3'b010 : node809;
											assign node809 = (inp[11]) ? 3'b010 : 3'b000;
								assign node814 = (inp[11]) ? node822 : node815;
									assign node815 = (inp[5]) ? node817 : 3'b010;
										assign node817 = (inp[3]) ? 3'b010 : node818;
											assign node818 = (inp[4]) ? 3'b010 : 3'b100;
									assign node822 = (inp[4]) ? node826 : node823;
										assign node823 = (inp[8]) ? 3'b000 : 3'b100;
										assign node826 = (inp[5]) ? 3'b000 : 3'b010;
							assign node829 = (inp[8]) ? node831 : 3'b000;
								assign node831 = (inp[5]) ? 3'b000 : node832;
									assign node832 = (inp[11]) ? node834 : 3'b000;
										assign node834 = (inp[4]) ? 3'b000 : 3'b010;
				assign node838 = (inp[2]) ? node840 : 3'b000;
					assign node840 = (inp[1]) ? node852 : node841;
						assign node841 = (inp[11]) ? 3'b000 : node842;
							assign node842 = (inp[5]) ? node844 : 3'b000;
								assign node844 = (inp[6]) ? node846 : 3'b000;
									assign node846 = (inp[3]) ? 3'b000 : node847;
										assign node847 = (inp[4]) ? 3'b010 : 3'b000;
						assign node852 = (inp[5]) ? node880 : node853;
							assign node853 = (inp[3]) ? node873 : node854;
								assign node854 = (inp[4]) ? node866 : node855;
									assign node855 = (inp[11]) ? node863 : node856;
										assign node856 = (inp[7]) ? node858 : 3'b000;
											assign node858 = (inp[8]) ? 3'b010 : node859;
												assign node859 = (inp[6]) ? 3'b010 : 3'b000;
										assign node863 = (inp[7]) ? 3'b000 : 3'b010;
									assign node866 = (inp[11]) ? 3'b000 : node867;
										assign node867 = (inp[8]) ? 3'b000 : node868;
											assign node868 = (inp[6]) ? 3'b100 : 3'b110;
								assign node873 = (inp[11]) ? 3'b000 : node874;
									assign node874 = (inp[6]) ? 3'b000 : node875;
										assign node875 = (inp[8]) ? 3'b000 : 3'b010;
							assign node880 = (inp[3]) ? 3'b000 : node881;
								assign node881 = (inp[7]) ? 3'b000 : node882;
									assign node882 = (inp[8]) ? 3'b000 : 3'b100;

endmodule