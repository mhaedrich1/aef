module dtc_split5_bm13 (
	input  wire [11-1:0] inp,
	output wire [1-1:0] outp
);

	wire [1-1:0] node1;
	wire [1-1:0] node2;
	wire [1-1:0] node3;
	wire [1-1:0] node4;
	wire [1-1:0] node6;
	wire [1-1:0] node8;
	wire [1-1:0] node10;
	wire [1-1:0] node12;
	wire [1-1:0] node15;
	wire [1-1:0] node16;
	wire [1-1:0] node18;
	wire [1-1:0] node20;
	wire [1-1:0] node22;
	wire [1-1:0] node25;
	wire [1-1:0] node26;
	wire [1-1:0] node28;
	wire [1-1:0] node30;
	wire [1-1:0] node33;
	wire [1-1:0] node34;
	wire [1-1:0] node36;
	wire [1-1:0] node40;
	wire [1-1:0] node41;
	wire [1-1:0] node42;
	wire [1-1:0] node44;
	wire [1-1:0] node46;
	wire [1-1:0] node48;
	wire [1-1:0] node51;
	wire [1-1:0] node52;
	wire [1-1:0] node54;
	wire [1-1:0] node56;
	wire [1-1:0] node59;
	wire [1-1:0] node60;
	wire [1-1:0] node62;
	wire [1-1:0] node65;
	wire [1-1:0] node66;
	wire [1-1:0] node70;
	wire [1-1:0] node71;
	wire [1-1:0] node72;
	wire [1-1:0] node74;
	wire [1-1:0] node76;
	wire [1-1:0] node79;
	wire [1-1:0] node80;
	wire [1-1:0] node82;
	wire [1-1:0] node85;
	wire [1-1:0] node86;
	wire [1-1:0] node90;
	wire [1-1:0] node91;
	wire [1-1:0] node92;
	wire [1-1:0] node94;
	wire [1-1:0] node97;
	wire [1-1:0] node98;
	wire [1-1:0] node102;
	wire [1-1:0] node103;
	wire [1-1:0] node107;
	wire [1-1:0] node108;
	wire [1-1:0] node109;
	wire [1-1:0] node110;
	wire [1-1:0] node112;
	wire [1-1:0] node114;
	wire [1-1:0] node115;
	wire [1-1:0] node118;
	wire [1-1:0] node121;
	wire [1-1:0] node122;
	wire [1-1:0] node124;
	wire [1-1:0] node126;
	wire [1-1:0] node129;
	wire [1-1:0] node130;
	wire [1-1:0] node132;
	wire [1-1:0] node135;
	wire [1-1:0] node136;
	wire [1-1:0] node140;
	wire [1-1:0] node141;
	wire [1-1:0] node143;
	wire [1-1:0] node144;
	wire [1-1:0] node145;
	wire [1-1:0] node148;
	wire [1-1:0] node151;
	wire [1-1:0] node152;
	wire [1-1:0] node156;
	wire [1-1:0] node157;
	wire [1-1:0] node158;
	wire [1-1:0] node160;
	wire [1-1:0] node163;
	wire [1-1:0] node164;
	wire [1-1:0] node168;
	wire [1-1:0] node169;
	wire [1-1:0] node170;
	wire [1-1:0] node175;
	wire [1-1:0] node176;
	wire [1-1:0] node177;
	wire [1-1:0] node178;
	wire [1-1:0] node180;
	wire [1-1:0] node183;
	wire [1-1:0] node184;
	wire [1-1:0] node186;
	wire [1-1:0] node189;
	wire [1-1:0] node190;
	wire [1-1:0] node194;
	wire [1-1:0] node195;
	wire [1-1:0] node196;
	wire [1-1:0] node197;
	wire [1-1:0] node200;
	wire [1-1:0] node205;
	wire [1-1:0] node206;
	wire [1-1:0] node207;
	wire [1-1:0] node209;
	wire [1-1:0] node211;
	wire [1-1:0] node214;
	wire [1-1:0] node215;
	wire [1-1:0] node216;
	wire [1-1:0] node221;
	wire [1-1:0] node222;
	wire [1-1:0] node223;
	wire [1-1:0] node224;
	wire [1-1:0] node230;
	wire [1-1:0] node231;
	wire [1-1:0] node232;
	wire [1-1:0] node233;
	wire [1-1:0] node235;
	wire [1-1:0] node236;
	wire [1-1:0] node238;
	wire [1-1:0] node240;
	wire [1-1:0] node243;
	wire [1-1:0] node244;
	wire [1-1:0] node246;
	wire [1-1:0] node250;
	wire [1-1:0] node251;
	wire [1-1:0] node252;
	wire [1-1:0] node254;
	wire [1-1:0] node256;
	wire [1-1:0] node259;
	wire [1-1:0] node260;
	wire [1-1:0] node262;
	wire [1-1:0] node265;
	wire [1-1:0] node266;
	wire [1-1:0] node270;
	wire [1-1:0] node271;
	wire [1-1:0] node272;
	wire [1-1:0] node274;
	wire [1-1:0] node277;
	wire [1-1:0] node278;
	wire [1-1:0] node282;
	wire [1-1:0] node283;
	wire [1-1:0] node287;
	wire [1-1:0] node288;
	wire [1-1:0] node289;
	wire [1-1:0] node290;
	wire [1-1:0] node292;
	wire [1-1:0] node294;
	wire [1-1:0] node297;
	wire [1-1:0] node298;
	wire [1-1:0] node300;
	wire [1-1:0] node303;
	wire [1-1:0] node304;
	wire [1-1:0] node308;
	wire [1-1:0] node309;
	wire [1-1:0] node310;
	wire [1-1:0] node312;
	wire [1-1:0] node315;
	wire [1-1:0] node316;
	wire [1-1:0] node320;
	wire [1-1:0] node321;
	wire [1-1:0] node322;
	wire [1-1:0] node327;
	wire [1-1:0] node328;
	wire [1-1:0] node329;
	wire [1-1:0] node330;
	wire [1-1:0] node332;
	wire [1-1:0] node335;
	wire [1-1:0] node336;
	wire [1-1:0] node340;
	wire [1-1:0] node341;
	wire [1-1:0] node342;
	wire [1-1:0] node347;
	wire [1-1:0] node348;
	wire [1-1:0] node349;
	wire [1-1:0] node350;
	wire [1-1:0] node356;
	wire [1-1:0] node357;
	wire [1-1:0] node358;
	wire [1-1:0] node359;
	wire [1-1:0] node360;
	wire [1-1:0] node362;
	wire [1-1:0] node364;
	wire [1-1:0] node367;
	wire [1-1:0] node368;
	wire [1-1:0] node370;
	wire [1-1:0] node373;
	wire [1-1:0] node374;
	wire [1-1:0] node378;
	wire [1-1:0] node379;
	wire [1-1:0] node380;
	wire [1-1:0] node382;
	wire [1-1:0] node385;
	wire [1-1:0] node386;
	wire [1-1:0] node391;
	wire [1-1:0] node392;
	wire [1-1:0] node393;
	wire [1-1:0] node394;
	wire [1-1:0] node396;
	wire [1-1:0] node399;
	wire [1-1:0] node400;
	wire [1-1:0] node404;
	wire [1-1:0] node405;
	wire [1-1:0] node406;
	wire [1-1:0] node411;
	wire [1-1:0] node412;
	wire [1-1:0] node413;
	wire [1-1:0] node414;
	wire [1-1:0] node420;
	wire [1-1:0] node421;
	wire [1-1:0] node422;
	wire [1-1:0] node423;
	wire [1-1:0] node424;
	wire [1-1:0] node426;
	wire [1-1:0] node429;
	wire [1-1:0] node430;
	wire [1-1:0] node434;
	wire [1-1:0] node435;
	wire [1-1:0] node436;
	wire [1-1:0] node439;
	wire [1-1:0] node443;
	wire [1-1:0] node444;
	wire [1-1:0] node445;
	wire [1-1:0] node446;

	assign outp = (inp[7]) ? node230 : node1;
		assign node1 = (inp[5]) ? node107 : node2;
			assign node2 = (inp[6]) ? node40 : node3;
				assign node3 = (inp[4]) ? node15 : node4;
					assign node4 = (inp[0]) ? node6 : 1'b1;
						assign node6 = (inp[8]) ? node8 : 1'b1;
							assign node8 = (inp[10]) ? node10 : 1'b1;
								assign node10 = (inp[3]) ? node12 : 1'b1;
									assign node12 = (inp[9]) ? 1'b0 : 1'b1;
					assign node15 = (inp[3]) ? node25 : node16;
						assign node16 = (inp[1]) ? node18 : 1'b1;
							assign node18 = (inp[2]) ? node20 : 1'b1;
								assign node20 = (inp[10]) ? node22 : 1'b1;
									assign node22 = (inp[8]) ? 1'b0 : 1'b1;
						assign node25 = (inp[0]) ? node33 : node26;
							assign node26 = (inp[2]) ? node28 : 1'b1;
								assign node28 = (inp[10]) ? node30 : 1'b1;
									assign node30 = (inp[8]) ? 1'b0 : 1'b1;
							assign node33 = (inp[1]) ? 1'b0 : node34;
								assign node34 = (inp[10]) ? node36 : 1'b1;
									assign node36 = (inp[8]) ? 1'b0 : 1'b1;
				assign node40 = (inp[2]) ? node70 : node41;
					assign node41 = (inp[8]) ? node51 : node42;
						assign node42 = (inp[3]) ? node44 : 1'b1;
							assign node44 = (inp[9]) ? node46 : 1'b1;
								assign node46 = (inp[1]) ? node48 : 1'b1;
									assign node48 = (inp[0]) ? 1'b0 : 1'b1;
						assign node51 = (inp[4]) ? node59 : node52;
							assign node52 = (inp[9]) ? node54 : 1'b1;
								assign node54 = (inp[3]) ? node56 : 1'b1;
									assign node56 = (inp[1]) ? 1'b0 : 1'b1;
							assign node59 = (inp[1]) ? node65 : node60;
								assign node60 = (inp[9]) ? node62 : 1'b1;
									assign node62 = (inp[0]) ? 1'b0 : 1'b1;
								assign node65 = (inp[0]) ? 1'b0 : node66;
									assign node66 = (inp[9]) ? 1'b0 : 1'b1;
					assign node70 = (inp[0]) ? node90 : node71;
						assign node71 = (inp[4]) ? node79 : node72;
							assign node72 = (inp[3]) ? node74 : 1'b1;
								assign node74 = (inp[10]) ? node76 : 1'b1;
									assign node76 = (inp[1]) ? 1'b0 : 1'b0;
							assign node79 = (inp[1]) ? node85 : node80;
								assign node80 = (inp[10]) ? node82 : 1'b1;
									assign node82 = (inp[9]) ? 1'b0 : 1'b1;
								assign node85 = (inp[3]) ? 1'b0 : node86;
									assign node86 = (inp[10]) ? 1'b0 : 1'b1;
						assign node90 = (inp[10]) ? node102 : node91;
							assign node91 = (inp[4]) ? node97 : node92;
								assign node92 = (inp[8]) ? node94 : 1'b1;
									assign node94 = (inp[3]) ? 1'b0 : 1'b1;
								assign node97 = (inp[1]) ? 1'b0 : node98;
									assign node98 = (inp[3]) ? 1'b0 : 1'b0;
							assign node102 = (inp[8]) ? 1'b0 : node103;
								assign node103 = (inp[9]) ? 1'b0 : 1'b1;
			assign node107 = (inp[1]) ? node175 : node108;
				assign node108 = (inp[2]) ? node140 : node109;
					assign node109 = (inp[0]) ? node121 : node110;
						assign node110 = (inp[3]) ? node112 : 1'b1;
							assign node112 = (inp[6]) ? node114 : 1'b1;
								assign node114 = (inp[4]) ? node118 : node115;
									assign node115 = (inp[10]) ? 1'b1 : 1'b1;
									assign node118 = (inp[9]) ? 1'b0 : 1'b0;
						assign node121 = (inp[4]) ? node129 : node122;
							assign node122 = (inp[10]) ? node124 : 1'b1;
								assign node124 = (inp[9]) ? node126 : 1'b1;
									assign node126 = (inp[8]) ? 1'b0 : 1'b1;
							assign node129 = (inp[8]) ? node135 : node130;
								assign node130 = (inp[10]) ? node132 : 1'b1;
									assign node132 = (inp[3]) ? 1'b0 : 1'b1;
								assign node135 = (inp[9]) ? 1'b0 : node136;
									assign node136 = (inp[10]) ? 1'b0 : 1'b1;
					assign node140 = (inp[10]) ? node156 : node141;
						assign node141 = (inp[4]) ? node143 : 1'b1;
							assign node143 = (inp[9]) ? node151 : node144;
								assign node144 = (inp[6]) ? node148 : node145;
									assign node145 = (inp[3]) ? 1'b1 : 1'b1;
									assign node148 = (inp[8]) ? 1'b0 : 1'b1;
								assign node151 = (inp[0]) ? 1'b0 : node152;
									assign node152 = (inp[8]) ? 1'b0 : 1'b1;
						assign node156 = (inp[0]) ? node168 : node157;
							assign node157 = (inp[8]) ? node163 : node158;
								assign node158 = (inp[6]) ? node160 : 1'b1;
									assign node160 = (inp[9]) ? 1'b0 : 1'b1;
								assign node163 = (inp[9]) ? 1'b0 : node164;
									assign node164 = (inp[6]) ? 1'b1 : 1'b0;
							assign node168 = (inp[3]) ? 1'b0 : node169;
								assign node169 = (inp[9]) ? 1'b0 : node170;
									assign node170 = (inp[6]) ? 1'b0 : 1'b1;
				assign node175 = (inp[8]) ? node205 : node176;
					assign node176 = (inp[2]) ? node194 : node177;
						assign node177 = (inp[0]) ? node183 : node178;
							assign node178 = (inp[3]) ? node180 : 1'b1;
								assign node180 = (inp[10]) ? 1'b0 : 1'b1;
							assign node183 = (inp[9]) ? node189 : node184;
								assign node184 = (inp[10]) ? node186 : 1'b1;
									assign node186 = (inp[3]) ? 1'b0 : 1'b1;
								assign node189 = (inp[6]) ? 1'b0 : node190;
									assign node190 = (inp[10]) ? 1'b0 : 1'b1;
						assign node194 = (inp[6]) ? 1'b0 : node195;
							assign node195 = (inp[10]) ? 1'b0 : node196;
								assign node196 = (inp[9]) ? node200 : node197;
									assign node197 = (inp[3]) ? 1'b1 : 1'b1;
									assign node200 = (inp[4]) ? 1'b0 : 1'b1;
					assign node205 = (inp[6]) ? node221 : node206;
						assign node206 = (inp[3]) ? node214 : node207;
							assign node207 = (inp[4]) ? node209 : 1'b1;
								assign node209 = (inp[0]) ? node211 : 1'b1;
									assign node211 = (inp[9]) ? 1'b0 : 1'b0;
							assign node214 = (inp[0]) ? 1'b0 : node215;
								assign node215 = (inp[9]) ? 1'b0 : node216;
									assign node216 = (inp[2]) ? 1'b0 : 1'b1;
						assign node221 = (inp[4]) ? 1'b0 : node222;
							assign node222 = (inp[2]) ? 1'b0 : node223;
								assign node223 = (inp[9]) ? 1'b0 : node224;
									assign node224 = (inp[3]) ? 1'b0 : 1'b1;
		assign node230 = (inp[9]) ? node356 : node231;
			assign node231 = (inp[3]) ? node287 : node232;
				assign node232 = (inp[8]) ? node250 : node233;
					assign node233 = (inp[4]) ? node235 : 1'b1;
						assign node235 = (inp[2]) ? node243 : node236;
							assign node236 = (inp[0]) ? node238 : 1'b1;
								assign node238 = (inp[5]) ? node240 : 1'b1;
									assign node240 = (inp[1]) ? 1'b0 : 1'b1;
							assign node243 = (inp[10]) ? 1'b0 : node244;
								assign node244 = (inp[6]) ? node246 : 1'b1;
									assign node246 = (inp[5]) ? 1'b0 : 1'b1;
					assign node250 = (inp[10]) ? node270 : node251;
						assign node251 = (inp[0]) ? node259 : node252;
							assign node252 = (inp[5]) ? node254 : 1'b1;
								assign node254 = (inp[6]) ? node256 : 1'b1;
									assign node256 = (inp[4]) ? 1'b0 : 1'b1;
							assign node259 = (inp[6]) ? node265 : node260;
								assign node260 = (inp[4]) ? node262 : 1'b1;
									assign node262 = (inp[1]) ? 1'b0 : 1'b1;
								assign node265 = (inp[2]) ? 1'b0 : node266;
									assign node266 = (inp[5]) ? 1'b0 : 1'b1;
						assign node270 = (inp[5]) ? node282 : node271;
							assign node271 = (inp[4]) ? node277 : node272;
								assign node272 = (inp[2]) ? node274 : 1'b1;
									assign node274 = (inp[6]) ? 1'b0 : 1'b1;
								assign node277 = (inp[6]) ? 1'b0 : node278;
									assign node278 = (inp[0]) ? 1'b0 : 1'b0;
							assign node282 = (inp[6]) ? 1'b0 : node283;
								assign node283 = (inp[2]) ? 1'b0 : 1'b1;
				assign node287 = (inp[2]) ? node327 : node288;
					assign node288 = (inp[4]) ? node308 : node289;
						assign node289 = (inp[1]) ? node297 : node290;
							assign node290 = (inp[10]) ? node292 : 1'b1;
								assign node292 = (inp[0]) ? node294 : 1'b1;
									assign node294 = (inp[5]) ? 1'b0 : 1'b1;
							assign node297 = (inp[8]) ? node303 : node298;
								assign node298 = (inp[5]) ? node300 : 1'b1;
									assign node300 = (inp[10]) ? 1'b0 : 1'b1;
								assign node303 = (inp[0]) ? 1'b0 : node304;
									assign node304 = (inp[5]) ? 1'b0 : 1'b1;
						assign node308 = (inp[8]) ? node320 : node309;
							assign node309 = (inp[5]) ? node315 : node310;
								assign node310 = (inp[0]) ? node312 : 1'b1;
									assign node312 = (inp[1]) ? 1'b0 : 1'b1;
								assign node315 = (inp[6]) ? 1'b0 : node316;
									assign node316 = (inp[1]) ? 1'b0 : 1'b1;
							assign node320 = (inp[10]) ? 1'b0 : node321;
								assign node321 = (inp[0]) ? 1'b0 : node322;
									assign node322 = (inp[1]) ? 1'b0 : 1'b1;
					assign node327 = (inp[6]) ? node347 : node328;
						assign node328 = (inp[8]) ? node340 : node329;
							assign node329 = (inp[10]) ? node335 : node330;
								assign node330 = (inp[5]) ? node332 : 1'b1;
									assign node332 = (inp[4]) ? 1'b0 : 1'b1;
								assign node335 = (inp[4]) ? 1'b0 : node336;
									assign node336 = (inp[1]) ? 1'b0 : 1'b1;
							assign node340 = (inp[5]) ? 1'b0 : node341;
								assign node341 = (inp[0]) ? 1'b0 : node342;
									assign node342 = (inp[10]) ? 1'b0 : 1'b1;
						assign node347 = (inp[4]) ? 1'b0 : node348;
							assign node348 = (inp[0]) ? 1'b0 : node349;
								assign node349 = (inp[5]) ? 1'b0 : node350;
									assign node350 = (inp[8]) ? 1'b0 : 1'b1;
			assign node356 = (inp[0]) ? node420 : node357;
				assign node357 = (inp[1]) ? node391 : node358;
					assign node358 = (inp[6]) ? node378 : node359;
						assign node359 = (inp[5]) ? node367 : node360;
							assign node360 = (inp[2]) ? node362 : 1'b1;
								assign node362 = (inp[10]) ? node364 : 1'b1;
									assign node364 = (inp[3]) ? 1'b0 : 1'b1;
							assign node367 = (inp[10]) ? node373 : node368;
								assign node368 = (inp[8]) ? node370 : 1'b1;
									assign node370 = (inp[4]) ? 1'b0 : 1'b1;
								assign node373 = (inp[3]) ? 1'b0 : node374;
									assign node374 = (inp[4]) ? 1'b0 : 1'b1;
						assign node378 = (inp[2]) ? 1'b0 : node379;
							assign node379 = (inp[3]) ? node385 : node380;
								assign node380 = (inp[8]) ? node382 : 1'b1;
									assign node382 = (inp[10]) ? 1'b0 : 1'b1;
								assign node385 = (inp[4]) ? 1'b0 : node386;
									assign node386 = (inp[5]) ? 1'b0 : 1'b1;
					assign node391 = (inp[10]) ? node411 : node392;
						assign node392 = (inp[4]) ? node404 : node393;
							assign node393 = (inp[8]) ? node399 : node394;
								assign node394 = (inp[5]) ? node396 : 1'b1;
									assign node396 = (inp[6]) ? 1'b0 : 1'b1;
								assign node399 = (inp[3]) ? 1'b0 : node400;
									assign node400 = (inp[5]) ? 1'b0 : 1'b1;
							assign node404 = (inp[5]) ? 1'b0 : node405;
								assign node405 = (inp[3]) ? 1'b0 : node406;
									assign node406 = (inp[6]) ? 1'b0 : 1'b1;
						assign node411 = (inp[4]) ? 1'b0 : node412;
							assign node412 = (inp[6]) ? 1'b0 : node413;
								assign node413 = (inp[2]) ? 1'b0 : node414;
									assign node414 = (inp[5]) ? 1'b0 : 1'b1;
				assign node420 = (inp[8]) ? 1'b0 : node421;
					assign node421 = (inp[2]) ? node443 : node422;
						assign node422 = (inp[4]) ? node434 : node423;
							assign node423 = (inp[6]) ? node429 : node424;
								assign node424 = (inp[5]) ? node426 : 1'b1;
									assign node426 = (inp[1]) ? 1'b0 : 1'b1;
								assign node429 = (inp[5]) ? 1'b0 : node430;
									assign node430 = (inp[3]) ? 1'b0 : 1'b1;
							assign node434 = (inp[1]) ? 1'b0 : node435;
								assign node435 = (inp[5]) ? node439 : node436;
									assign node436 = (inp[10]) ? 1'b0 : 1'b1;
									assign node439 = (inp[6]) ? 1'b0 : 1'b0;
						assign node443 = (inp[5]) ? 1'b0 : node444;
							assign node444 = (inp[4]) ? 1'b0 : node445;
								assign node445 = (inp[10]) ? 1'b0 : node446;
									assign node446 = (inp[3]) ? 1'b0 : 1'b1;

endmodule