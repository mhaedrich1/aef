module dtc_split66_bm83 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node7;
	wire [3-1:0] node8;
	wire [3-1:0] node9;
	wire [3-1:0] node10;
	wire [3-1:0] node13;
	wire [3-1:0] node14;
	wire [3-1:0] node18;
	wire [3-1:0] node20;
	wire [3-1:0] node23;
	wire [3-1:0] node24;
	wire [3-1:0] node25;
	wire [3-1:0] node26;
	wire [3-1:0] node30;
	wire [3-1:0] node31;
	wire [3-1:0] node35;
	wire [3-1:0] node36;
	wire [3-1:0] node37;
	wire [3-1:0] node41;
	wire [3-1:0] node44;
	wire [3-1:0] node45;
	wire [3-1:0] node46;
	wire [3-1:0] node49;
	wire [3-1:0] node52;
	wire [3-1:0] node53;
	wire [3-1:0] node57;
	wire [3-1:0] node58;
	wire [3-1:0] node59;
	wire [3-1:0] node60;
	wire [3-1:0] node63;
	wire [3-1:0] node65;
	wire [3-1:0] node67;
	wire [3-1:0] node70;
	wire [3-1:0] node71;
	wire [3-1:0] node73;
	wire [3-1:0] node76;
	wire [3-1:0] node77;
	wire [3-1:0] node78;
	wire [3-1:0] node83;
	wire [3-1:0] node84;
	wire [3-1:0] node87;
	wire [3-1:0] node89;
	wire [3-1:0] node92;
	wire [3-1:0] node93;
	wire [3-1:0] node94;
	wire [3-1:0] node95;
	wire [3-1:0] node96;
	wire [3-1:0] node97;
	wire [3-1:0] node100;
	wire [3-1:0] node101;
	wire [3-1:0] node105;
	wire [3-1:0] node106;
	wire [3-1:0] node109;
	wire [3-1:0] node112;
	wire [3-1:0] node113;
	wire [3-1:0] node114;
	wire [3-1:0] node117;
	wire [3-1:0] node121;
	wire [3-1:0] node122;
	wire [3-1:0] node123;
	wire [3-1:0] node126;
	wire [3-1:0] node127;
	wire [3-1:0] node129;
	wire [3-1:0] node133;
	wire [3-1:0] node134;
	wire [3-1:0] node136;
	wire [3-1:0] node139;
	wire [3-1:0] node140;
	wire [3-1:0] node142;
	wire [3-1:0] node145;
	wire [3-1:0] node148;
	wire [3-1:0] node149;
	wire [3-1:0] node150;
	wire [3-1:0] node151;
	wire [3-1:0] node152;
	wire [3-1:0] node155;
	wire [3-1:0] node156;
	wire [3-1:0] node160;
	wire [3-1:0] node161;
	wire [3-1:0] node162;
	wire [3-1:0] node167;
	wire [3-1:0] node168;
	wire [3-1:0] node170;
	wire [3-1:0] node173;
	wire [3-1:0] node174;
	wire [3-1:0] node179;
	wire [3-1:0] node180;
	wire [3-1:0] node181;
	wire [3-1:0] node182;
	wire [3-1:0] node184;
	wire [3-1:0] node186;
	wire [3-1:0] node190;
	wire [3-1:0] node191;
	wire [3-1:0] node193;
	wire [3-1:0] node194;
	wire [3-1:0] node196;
	wire [3-1:0] node199;
	wire [3-1:0] node200;
	wire [3-1:0] node205;
	wire [3-1:0] node206;
	wire [3-1:0] node207;
	wire [3-1:0] node209;
	wire [3-1:0] node210;
	wire [3-1:0] node212;
	wire [3-1:0] node216;
	wire [3-1:0] node217;
	wire [3-1:0] node219;
	wire [3-1:0] node221;
	wire [3-1:0] node224;
	wire [3-1:0] node225;
	wire [3-1:0] node229;
	wire [3-1:0] node231;
	wire [3-1:0] node232;
	wire [3-1:0] node233;
	wire [3-1:0] node235;
	wire [3-1:0] node237;
	wire [3-1:0] node242;
	wire [3-1:0] node243;
	wire [3-1:0] node244;
	wire [3-1:0] node245;
	wire [3-1:0] node246;
	wire [3-1:0] node247;
	wire [3-1:0] node248;
	wire [3-1:0] node249;
	wire [3-1:0] node250;
	wire [3-1:0] node255;
	wire [3-1:0] node258;
	wire [3-1:0] node260;
	wire [3-1:0] node261;
	wire [3-1:0] node264;
	wire [3-1:0] node266;
	wire [3-1:0] node269;
	wire [3-1:0] node270;
	wire [3-1:0] node271;
	wire [3-1:0] node275;
	wire [3-1:0] node276;
	wire [3-1:0] node277;
	wire [3-1:0] node279;
	wire [3-1:0] node283;
	wire [3-1:0] node286;
	wire [3-1:0] node287;
	wire [3-1:0] node288;
	wire [3-1:0] node289;
	wire [3-1:0] node290;
	wire [3-1:0] node291;
	wire [3-1:0] node296;
	wire [3-1:0] node297;
	wire [3-1:0] node300;
	wire [3-1:0] node302;
	wire [3-1:0] node305;
	wire [3-1:0] node306;
	wire [3-1:0] node309;
	wire [3-1:0] node311;
	wire [3-1:0] node314;
	wire [3-1:0] node315;
	wire [3-1:0] node316;
	wire [3-1:0] node318;
	wire [3-1:0] node320;
	wire [3-1:0] node324;
	wire [3-1:0] node326;
	wire [3-1:0] node328;
	wire [3-1:0] node331;
	wire [3-1:0] node332;
	wire [3-1:0] node333;
	wire [3-1:0] node334;
	wire [3-1:0] node335;
	wire [3-1:0] node336;
	wire [3-1:0] node339;
	wire [3-1:0] node342;
	wire [3-1:0] node343;
	wire [3-1:0] node346;
	wire [3-1:0] node349;
	wire [3-1:0] node350;
	wire [3-1:0] node352;
	wire [3-1:0] node355;
	wire [3-1:0] node357;
	wire [3-1:0] node359;
	wire [3-1:0] node362;
	wire [3-1:0] node363;
	wire [3-1:0] node364;
	wire [3-1:0] node366;
	wire [3-1:0] node370;
	wire [3-1:0] node372;
	wire [3-1:0] node374;
	wire [3-1:0] node376;
	wire [3-1:0] node379;
	wire [3-1:0] node380;
	wire [3-1:0] node381;
	wire [3-1:0] node383;
	wire [3-1:0] node384;
	wire [3-1:0] node388;
	wire [3-1:0] node389;
	wire [3-1:0] node391;
	wire [3-1:0] node394;
	wire [3-1:0] node396;
	wire [3-1:0] node397;
	wire [3-1:0] node401;
	wire [3-1:0] node402;
	wire [3-1:0] node404;
	wire [3-1:0] node406;
	wire [3-1:0] node408;
	wire [3-1:0] node411;
	wire [3-1:0] node412;
	wire [3-1:0] node415;
	wire [3-1:0] node417;
	wire [3-1:0] node419;
	wire [3-1:0] node422;
	wire [3-1:0] node423;
	wire [3-1:0] node424;
	wire [3-1:0] node425;
	wire [3-1:0] node426;
	wire [3-1:0] node428;
	wire [3-1:0] node429;
	wire [3-1:0] node432;
	wire [3-1:0] node435;
	wire [3-1:0] node437;
	wire [3-1:0] node439;
	wire [3-1:0] node440;
	wire [3-1:0] node444;
	wire [3-1:0] node445;
	wire [3-1:0] node446;
	wire [3-1:0] node448;
	wire [3-1:0] node451;
	wire [3-1:0] node452;
	wire [3-1:0] node455;
	wire [3-1:0] node458;
	wire [3-1:0] node459;
	wire [3-1:0] node460;
	wire [3-1:0] node462;
	wire [3-1:0] node465;
	wire [3-1:0] node468;
	wire [3-1:0] node469;
	wire [3-1:0] node470;
	wire [3-1:0] node474;
	wire [3-1:0] node475;
	wire [3-1:0] node479;
	wire [3-1:0] node480;
	wire [3-1:0] node481;
	wire [3-1:0] node482;
	wire [3-1:0] node483;
	wire [3-1:0] node485;
	wire [3-1:0] node489;
	wire [3-1:0] node490;
	wire [3-1:0] node493;
	wire [3-1:0] node496;
	wire [3-1:0] node497;
	wire [3-1:0] node498;
	wire [3-1:0] node501;
	wire [3-1:0] node503;
	wire [3-1:0] node506;
	wire [3-1:0] node508;
	wire [3-1:0] node509;
	wire [3-1:0] node513;
	wire [3-1:0] node514;
	wire [3-1:0] node515;
	wire [3-1:0] node516;
	wire [3-1:0] node519;
	wire [3-1:0] node520;
	wire [3-1:0] node524;
	wire [3-1:0] node525;
	wire [3-1:0] node529;
	wire [3-1:0] node531;
	wire [3-1:0] node532;
	wire [3-1:0] node536;
	wire [3-1:0] node537;
	wire [3-1:0] node538;
	wire [3-1:0] node539;
	wire [3-1:0] node540;
	wire [3-1:0] node541;
	wire [3-1:0] node543;
	wire [3-1:0] node546;
	wire [3-1:0] node548;
	wire [3-1:0] node553;
	wire [3-1:0] node554;
	wire [3-1:0] node556;
	wire [3-1:0] node558;
	wire [3-1:0] node561;
	wire [3-1:0] node563;
	wire [3-1:0] node566;
	wire [3-1:0] node567;
	wire [3-1:0] node568;
	wire [3-1:0] node569;
	wire [3-1:0] node570;
	wire [3-1:0] node574;
	wire [3-1:0] node575;
	wire [3-1:0] node576;
	wire [3-1:0] node581;
	wire [3-1:0] node583;
	wire [3-1:0] node586;
	wire [3-1:0] node587;
	wire [3-1:0] node588;
	wire [3-1:0] node589;
	wire [3-1:0] node590;
	wire [3-1:0] node594;
	wire [3-1:0] node596;
	wire [3-1:0] node599;
	wire [3-1:0] node600;
	wire [3-1:0] node601;
	wire [3-1:0] node606;
	wire [3-1:0] node607;
	wire [3-1:0] node609;
	wire [3-1:0] node612;
	wire [3-1:0] node614;
	wire [3-1:0] node615;
	wire [3-1:0] node619;
	wire [3-1:0] node620;
	wire [3-1:0] node621;
	wire [3-1:0] node622;
	wire [3-1:0] node623;
	wire [3-1:0] node624;
	wire [3-1:0] node625;
	wire [3-1:0] node626;
	wire [3-1:0] node627;
	wire [3-1:0] node631;
	wire [3-1:0] node634;
	wire [3-1:0] node637;
	wire [3-1:0] node638;
	wire [3-1:0] node639;
	wire [3-1:0] node642;
	wire [3-1:0] node643;
	wire [3-1:0] node644;
	wire [3-1:0] node649;
	wire [3-1:0] node650;
	wire [3-1:0] node651;
	wire [3-1:0] node655;
	wire [3-1:0] node658;
	wire [3-1:0] node659;
	wire [3-1:0] node660;
	wire [3-1:0] node662;
	wire [3-1:0] node663;
	wire [3-1:0] node664;
	wire [3-1:0] node668;
	wire [3-1:0] node671;
	wire [3-1:0] node672;
	wire [3-1:0] node673;
	wire [3-1:0] node676;
	wire [3-1:0] node679;
	wire [3-1:0] node680;
	wire [3-1:0] node682;
	wire [3-1:0] node685;
	wire [3-1:0] node686;
	wire [3-1:0] node690;
	wire [3-1:0] node691;
	wire [3-1:0] node692;
	wire [3-1:0] node693;
	wire [3-1:0] node696;
	wire [3-1:0] node697;
	wire [3-1:0] node701;
	wire [3-1:0] node702;
	wire [3-1:0] node703;
	wire [3-1:0] node707;
	wire [3-1:0] node710;
	wire [3-1:0] node711;
	wire [3-1:0] node712;
	wire [3-1:0] node713;
	wire [3-1:0] node717;
	wire [3-1:0] node718;
	wire [3-1:0] node721;
	wire [3-1:0] node724;
	wire [3-1:0] node727;
	wire [3-1:0] node728;
	wire [3-1:0] node729;
	wire [3-1:0] node730;
	wire [3-1:0] node731;
	wire [3-1:0] node732;
	wire [3-1:0] node733;
	wire [3-1:0] node738;
	wire [3-1:0] node740;
	wire [3-1:0] node741;
	wire [3-1:0] node744;
	wire [3-1:0] node747;
	wire [3-1:0] node749;
	wire [3-1:0] node751;
	wire [3-1:0] node754;
	wire [3-1:0] node755;
	wire [3-1:0] node756;
	wire [3-1:0] node757;
	wire [3-1:0] node761;
	wire [3-1:0] node763;
	wire [3-1:0] node766;
	wire [3-1:0] node767;
	wire [3-1:0] node769;
	wire [3-1:0] node772;
	wire [3-1:0] node774;
	wire [3-1:0] node776;
	wire [3-1:0] node779;
	wire [3-1:0] node780;
	wire [3-1:0] node781;
	wire [3-1:0] node782;
	wire [3-1:0] node784;
	wire [3-1:0] node787;
	wire [3-1:0] node788;
	wire [3-1:0] node792;
	wire [3-1:0] node793;
	wire [3-1:0] node795;
	wire [3-1:0] node797;
	wire [3-1:0] node800;
	wire [3-1:0] node801;
	wire [3-1:0] node805;
	wire [3-1:0] node806;
	wire [3-1:0] node807;
	wire [3-1:0] node808;
	wire [3-1:0] node812;
	wire [3-1:0] node813;
	wire [3-1:0] node817;
	wire [3-1:0] node818;
	wire [3-1:0] node819;
	wire [3-1:0] node821;
	wire [3-1:0] node825;
	wire [3-1:0] node826;
	wire [3-1:0] node830;
	wire [3-1:0] node831;
	wire [3-1:0] node832;
	wire [3-1:0] node833;
	wire [3-1:0] node834;
	wire [3-1:0] node835;
	wire [3-1:0] node836;
	wire [3-1:0] node837;
	wire [3-1:0] node840;
	wire [3-1:0] node843;
	wire [3-1:0] node847;
	wire [3-1:0] node848;
	wire [3-1:0] node849;
	wire [3-1:0] node850;
	wire [3-1:0] node853;
	wire [3-1:0] node857;
	wire [3-1:0] node858;
	wire [3-1:0] node862;
	wire [3-1:0] node863;
	wire [3-1:0] node864;
	wire [3-1:0] node865;
	wire [3-1:0] node867;
	wire [3-1:0] node870;
	wire [3-1:0] node872;
	wire [3-1:0] node875;
	wire [3-1:0] node877;
	wire [3-1:0] node879;
	wire [3-1:0] node882;
	wire [3-1:0] node883;
	wire [3-1:0] node884;
	wire [3-1:0] node886;
	wire [3-1:0] node891;
	wire [3-1:0] node892;
	wire [3-1:0] node893;
	wire [3-1:0] node894;
	wire [3-1:0] node896;
	wire [3-1:0] node897;
	wire [3-1:0] node900;
	wire [3-1:0] node903;
	wire [3-1:0] node904;
	wire [3-1:0] node905;
	wire [3-1:0] node909;
	wire [3-1:0] node911;
	wire [3-1:0] node914;
	wire [3-1:0] node915;
	wire [3-1:0] node916;
	wire [3-1:0] node920;
	wire [3-1:0] node921;
	wire [3-1:0] node924;
	wire [3-1:0] node927;
	wire [3-1:0] node928;
	wire [3-1:0] node929;
	wire [3-1:0] node930;
	wire [3-1:0] node931;
	wire [3-1:0] node934;
	wire [3-1:0] node937;
	wire [3-1:0] node938;
	wire [3-1:0] node942;
	wire [3-1:0] node943;
	wire [3-1:0] node944;
	wire [3-1:0] node949;
	wire [3-1:0] node950;
	wire [3-1:0] node951;
	wire [3-1:0] node952;
	wire [3-1:0] node957;
	wire [3-1:0] node958;
	wire [3-1:0] node961;
	wire [3-1:0] node962;
	wire [3-1:0] node966;
	wire [3-1:0] node967;
	wire [3-1:0] node968;
	wire [3-1:0] node969;
	wire [3-1:0] node970;
	wire [3-1:0] node973;
	wire [3-1:0] node975;
	wire [3-1:0] node976;
	wire [3-1:0] node980;
	wire [3-1:0] node981;
	wire [3-1:0] node982;
	wire [3-1:0] node984;
	wire [3-1:0] node988;
	wire [3-1:0] node991;
	wire [3-1:0] node992;
	wire [3-1:0] node993;
	wire [3-1:0] node994;
	wire [3-1:0] node998;
	wire [3-1:0] node999;
	wire [3-1:0] node1003;
	wire [3-1:0] node1005;
	wire [3-1:0] node1007;
	wire [3-1:0] node1010;
	wire [3-1:0] node1011;
	wire [3-1:0] node1012;
	wire [3-1:0] node1013;
	wire [3-1:0] node1014;
	wire [3-1:0] node1017;
	wire [3-1:0] node1020;
	wire [3-1:0] node1022;
	wire [3-1:0] node1025;
	wire [3-1:0] node1026;
	wire [3-1:0] node1028;
	wire [3-1:0] node1031;
	wire [3-1:0] node1033;
	wire [3-1:0] node1035;
	wire [3-1:0] node1038;
	wire [3-1:0] node1039;
	wire [3-1:0] node1040;
	wire [3-1:0] node1041;
	wire [3-1:0] node1044;
	wire [3-1:0] node1045;
	wire [3-1:0] node1049;
	wire [3-1:0] node1050;
	wire [3-1:0] node1053;
	wire [3-1:0] node1056;
	wire [3-1:0] node1058;
	wire [3-1:0] node1059;
	wire [3-1:0] node1062;
	wire [3-1:0] node1064;
	wire [3-1:0] node1067;
	wire [3-1:0] node1068;
	wire [3-1:0] node1069;
	wire [3-1:0] node1070;
	wire [3-1:0] node1071;
	wire [3-1:0] node1072;
	wire [3-1:0] node1073;
	wire [3-1:0] node1074;
	wire [3-1:0] node1078;
	wire [3-1:0] node1079;
	wire [3-1:0] node1083;
	wire [3-1:0] node1084;
	wire [3-1:0] node1085;
	wire [3-1:0] node1088;
	wire [3-1:0] node1090;
	wire [3-1:0] node1093;
	wire [3-1:0] node1094;
	wire [3-1:0] node1097;
	wire [3-1:0] node1098;
	wire [3-1:0] node1101;
	wire [3-1:0] node1104;
	wire [3-1:0] node1105;
	wire [3-1:0] node1106;
	wire [3-1:0] node1108;
	wire [3-1:0] node1109;
	wire [3-1:0] node1113;
	wire [3-1:0] node1115;
	wire [3-1:0] node1118;
	wire [3-1:0] node1119;
	wire [3-1:0] node1120;
	wire [3-1:0] node1123;
	wire [3-1:0] node1124;
	wire [3-1:0] node1128;
	wire [3-1:0] node1130;
	wire [3-1:0] node1131;
	wire [3-1:0] node1134;
	wire [3-1:0] node1137;
	wire [3-1:0] node1138;
	wire [3-1:0] node1139;
	wire [3-1:0] node1140;
	wire [3-1:0] node1141;
	wire [3-1:0] node1144;
	wire [3-1:0] node1145;
	wire [3-1:0] node1149;
	wire [3-1:0] node1151;
	wire [3-1:0] node1152;
	wire [3-1:0] node1156;
	wire [3-1:0] node1157;
	wire [3-1:0] node1159;
	wire [3-1:0] node1163;
	wire [3-1:0] node1164;
	wire [3-1:0] node1165;
	wire [3-1:0] node1166;
	wire [3-1:0] node1167;
	wire [3-1:0] node1172;
	wire [3-1:0] node1173;
	wire [3-1:0] node1174;
	wire [3-1:0] node1178;
	wire [3-1:0] node1179;
	wire [3-1:0] node1183;
	wire [3-1:0] node1184;
	wire [3-1:0] node1186;
	wire [3-1:0] node1189;
	wire [3-1:0] node1190;
	wire [3-1:0] node1192;
	wire [3-1:0] node1195;
	wire [3-1:0] node1198;
	wire [3-1:0] node1199;
	wire [3-1:0] node1200;
	wire [3-1:0] node1201;
	wire [3-1:0] node1202;
	wire [3-1:0] node1205;
	wire [3-1:0] node1206;
	wire [3-1:0] node1208;
	wire [3-1:0] node1212;
	wire [3-1:0] node1213;
	wire [3-1:0] node1214;
	wire [3-1:0] node1216;
	wire [3-1:0] node1219;
	wire [3-1:0] node1220;
	wire [3-1:0] node1224;
	wire [3-1:0] node1227;
	wire [3-1:0] node1228;
	wire [3-1:0] node1229;
	wire [3-1:0] node1231;
	wire [3-1:0] node1233;
	wire [3-1:0] node1236;
	wire [3-1:0] node1239;
	wire [3-1:0] node1240;
	wire [3-1:0] node1242;
	wire [3-1:0] node1243;
	wire [3-1:0] node1247;
	wire [3-1:0] node1248;
	wire [3-1:0] node1250;
	wire [3-1:0] node1254;
	wire [3-1:0] node1255;
	wire [3-1:0] node1256;
	wire [3-1:0] node1258;
	wire [3-1:0] node1259;
	wire [3-1:0] node1262;
	wire [3-1:0] node1265;
	wire [3-1:0] node1266;
	wire [3-1:0] node1268;
	wire [3-1:0] node1270;
	wire [3-1:0] node1274;
	wire [3-1:0] node1275;
	wire [3-1:0] node1277;
	wire [3-1:0] node1278;
	wire [3-1:0] node1282;
	wire [3-1:0] node1283;
	wire [3-1:0] node1286;
	wire [3-1:0] node1289;
	wire [3-1:0] node1290;
	wire [3-1:0] node1291;
	wire [3-1:0] node1292;
	wire [3-1:0] node1293;
	wire [3-1:0] node1294;
	wire [3-1:0] node1296;
	wire [3-1:0] node1298;
	wire [3-1:0] node1301;
	wire [3-1:0] node1302;
	wire [3-1:0] node1303;
	wire [3-1:0] node1308;
	wire [3-1:0] node1310;
	wire [3-1:0] node1311;
	wire [3-1:0] node1313;
	wire [3-1:0] node1316;
	wire [3-1:0] node1319;
	wire [3-1:0] node1320;
	wire [3-1:0] node1321;
	wire [3-1:0] node1324;
	wire [3-1:0] node1327;
	wire [3-1:0] node1328;
	wire [3-1:0] node1330;
	wire [3-1:0] node1332;
	wire [3-1:0] node1335;
	wire [3-1:0] node1337;
	wire [3-1:0] node1338;
	wire [3-1:0] node1342;
	wire [3-1:0] node1343;
	wire [3-1:0] node1344;
	wire [3-1:0] node1345;
	wire [3-1:0] node1346;
	wire [3-1:0] node1348;
	wire [3-1:0] node1352;
	wire [3-1:0] node1355;
	wire [3-1:0] node1356;
	wire [3-1:0] node1358;
	wire [3-1:0] node1361;
	wire [3-1:0] node1362;
	wire [3-1:0] node1364;
	wire [3-1:0] node1368;
	wire [3-1:0] node1369;
	wire [3-1:0] node1370;
	wire [3-1:0] node1371;
	wire [3-1:0] node1373;
	wire [3-1:0] node1376;
	wire [3-1:0] node1380;
	wire [3-1:0] node1381;
	wire [3-1:0] node1383;
	wire [3-1:0] node1384;
	wire [3-1:0] node1388;
	wire [3-1:0] node1390;
	wire [3-1:0] node1391;
	wire [3-1:0] node1394;
	wire [3-1:0] node1397;
	wire [3-1:0] node1398;
	wire [3-1:0] node1399;
	wire [3-1:0] node1400;
	wire [3-1:0] node1401;
	wire [3-1:0] node1402;
	wire [3-1:0] node1403;
	wire [3-1:0] node1406;
	wire [3-1:0] node1410;
	wire [3-1:0] node1411;
	wire [3-1:0] node1412;
	wire [3-1:0] node1417;
	wire [3-1:0] node1419;
	wire [3-1:0] node1420;
	wire [3-1:0] node1421;
	wire [3-1:0] node1424;
	wire [3-1:0] node1428;
	wire [3-1:0] node1429;
	wire [3-1:0] node1430;
	wire [3-1:0] node1432;
	wire [3-1:0] node1434;
	wire [3-1:0] node1437;
	wire [3-1:0] node1440;
	wire [3-1:0] node1441;
	wire [3-1:0] node1443;
	wire [3-1:0] node1445;
	wire [3-1:0] node1449;
	wire [3-1:0] node1450;
	wire [3-1:0] node1451;
	wire [3-1:0] node1452;
	wire [3-1:0] node1453;
	wire [3-1:0] node1457;
	wire [3-1:0] node1460;
	wire [3-1:0] node1461;
	wire [3-1:0] node1463;
	wire [3-1:0] node1466;
	wire [3-1:0] node1468;
	wire [3-1:0] node1469;
	wire [3-1:0] node1473;
	wire [3-1:0] node1474;
	wire [3-1:0] node1475;
	wire [3-1:0] node1476;
	wire [3-1:0] node1477;
	wire [3-1:0] node1481;
	wire [3-1:0] node1482;
	wire [3-1:0] node1486;
	wire [3-1:0] node1487;
	wire [3-1:0] node1491;
	wire [3-1:0] node1492;
	wire [3-1:0] node1493;
	wire [3-1:0] node1494;
	wire [3-1:0] node1499;
	wire [3-1:0] node1502;
	wire [3-1:0] node1503;
	wire [3-1:0] node1504;
	wire [3-1:0] node1505;
	wire [3-1:0] node1506;
	wire [3-1:0] node1507;
	wire [3-1:0] node1508;
	wire [3-1:0] node1509;
	wire [3-1:0] node1510;
	wire [3-1:0] node1512;
	wire [3-1:0] node1513;
	wire [3-1:0] node1517;
	wire [3-1:0] node1518;
	wire [3-1:0] node1519;
	wire [3-1:0] node1524;
	wire [3-1:0] node1525;
	wire [3-1:0] node1527;
	wire [3-1:0] node1529;
	wire [3-1:0] node1532;
	wire [3-1:0] node1533;
	wire [3-1:0] node1537;
	wire [3-1:0] node1538;
	wire [3-1:0] node1539;
	wire [3-1:0] node1540;
	wire [3-1:0] node1542;
	wire [3-1:0] node1545;
	wire [3-1:0] node1547;
	wire [3-1:0] node1550;
	wire [3-1:0] node1552;
	wire [3-1:0] node1554;
	wire [3-1:0] node1557;
	wire [3-1:0] node1558;
	wire [3-1:0] node1559;
	wire [3-1:0] node1560;
	wire [3-1:0] node1564;
	wire [3-1:0] node1566;
	wire [3-1:0] node1569;
	wire [3-1:0] node1571;
	wire [3-1:0] node1574;
	wire [3-1:0] node1575;
	wire [3-1:0] node1576;
	wire [3-1:0] node1577;
	wire [3-1:0] node1578;
	wire [3-1:0] node1583;
	wire [3-1:0] node1584;
	wire [3-1:0] node1585;
	wire [3-1:0] node1588;
	wire [3-1:0] node1591;
	wire [3-1:0] node1592;
	wire [3-1:0] node1595;
	wire [3-1:0] node1596;
	wire [3-1:0] node1600;
	wire [3-1:0] node1601;
	wire [3-1:0] node1602;
	wire [3-1:0] node1604;
	wire [3-1:0] node1605;
	wire [3-1:0] node1609;
	wire [3-1:0] node1613;
	wire [3-1:0] node1614;
	wire [3-1:0] node1615;
	wire [3-1:0] node1616;
	wire [3-1:0] node1617;
	wire [3-1:0] node1619;
	wire [3-1:0] node1622;
	wire [3-1:0] node1624;
	wire [3-1:0] node1627;
	wire [3-1:0] node1628;
	wire [3-1:0] node1632;
	wire [3-1:0] node1633;
	wire [3-1:0] node1634;
	wire [3-1:0] node1636;
	wire [3-1:0] node1639;
	wire [3-1:0] node1641;
	wire [3-1:0] node1644;
	wire [3-1:0] node1645;
	wire [3-1:0] node1647;
	wire [3-1:0] node1649;
	wire [3-1:0] node1652;
	wire [3-1:0] node1654;
	wire [3-1:0] node1657;
	wire [3-1:0] node1658;
	wire [3-1:0] node1659;
	wire [3-1:0] node1660;
	wire [3-1:0] node1663;
	wire [3-1:0] node1664;
	wire [3-1:0] node1665;
	wire [3-1:0] node1668;
	wire [3-1:0] node1672;
	wire [3-1:0] node1673;
	wire [3-1:0] node1674;
	wire [3-1:0] node1677;
	wire [3-1:0] node1679;
	wire [3-1:0] node1682;
	wire [3-1:0] node1683;
	wire [3-1:0] node1684;
	wire [3-1:0] node1688;
	wire [3-1:0] node1689;
	wire [3-1:0] node1693;
	wire [3-1:0] node1694;
	wire [3-1:0] node1695;
	wire [3-1:0] node1698;
	wire [3-1:0] node1700;
	wire [3-1:0] node1703;
	wire [3-1:0] node1704;
	wire [3-1:0] node1705;
	wire [3-1:0] node1706;
	wire [3-1:0] node1711;
	wire [3-1:0] node1714;
	wire [3-1:0] node1715;
	wire [3-1:0] node1716;
	wire [3-1:0] node1717;
	wire [3-1:0] node1718;
	wire [3-1:0] node1719;
	wire [3-1:0] node1721;
	wire [3-1:0] node1724;
	wire [3-1:0] node1725;
	wire [3-1:0] node1727;
	wire [3-1:0] node1731;
	wire [3-1:0] node1732;
	wire [3-1:0] node1733;
	wire [3-1:0] node1737;
	wire [3-1:0] node1739;
	wire [3-1:0] node1740;
	wire [3-1:0] node1744;
	wire [3-1:0] node1746;
	wire [3-1:0] node1747;
	wire [3-1:0] node1749;
	wire [3-1:0] node1752;
	wire [3-1:0] node1754;
	wire [3-1:0] node1755;
	wire [3-1:0] node1759;
	wire [3-1:0] node1760;
	wire [3-1:0] node1761;
	wire [3-1:0] node1762;
	wire [3-1:0] node1764;
	wire [3-1:0] node1767;
	wire [3-1:0] node1769;
	wire [3-1:0] node1771;
	wire [3-1:0] node1774;
	wire [3-1:0] node1775;
	wire [3-1:0] node1776;
	wire [3-1:0] node1780;
	wire [3-1:0] node1781;
	wire [3-1:0] node1783;
	wire [3-1:0] node1786;
	wire [3-1:0] node1787;
	wire [3-1:0] node1791;
	wire [3-1:0] node1792;
	wire [3-1:0] node1793;
	wire [3-1:0] node1796;
	wire [3-1:0] node1797;
	wire [3-1:0] node1800;
	wire [3-1:0] node1801;
	wire [3-1:0] node1804;
	wire [3-1:0] node1807;
	wire [3-1:0] node1808;
	wire [3-1:0] node1809;
	wire [3-1:0] node1810;
	wire [3-1:0] node1814;
	wire [3-1:0] node1817;
	wire [3-1:0] node1819;
	wire [3-1:0] node1821;
	wire [3-1:0] node1824;
	wire [3-1:0] node1825;
	wire [3-1:0] node1826;
	wire [3-1:0] node1827;
	wire [3-1:0] node1828;
	wire [3-1:0] node1829;
	wire [3-1:0] node1833;
	wire [3-1:0] node1834;
	wire [3-1:0] node1837;
	wire [3-1:0] node1840;
	wire [3-1:0] node1841;
	wire [3-1:0] node1842;
	wire [3-1:0] node1846;
	wire [3-1:0] node1848;
	wire [3-1:0] node1849;
	wire [3-1:0] node1853;
	wire [3-1:0] node1854;
	wire [3-1:0] node1855;
	wire [3-1:0] node1856;
	wire [3-1:0] node1857;
	wire [3-1:0] node1862;
	wire [3-1:0] node1863;
	wire [3-1:0] node1867;
	wire [3-1:0] node1868;
	wire [3-1:0] node1869;
	wire [3-1:0] node1872;
	wire [3-1:0] node1875;
	wire [3-1:0] node1876;
	wire [3-1:0] node1880;
	wire [3-1:0] node1881;
	wire [3-1:0] node1882;
	wire [3-1:0] node1883;
	wire [3-1:0] node1885;
	wire [3-1:0] node1888;
	wire [3-1:0] node1890;
	wire [3-1:0] node1891;
	wire [3-1:0] node1895;
	wire [3-1:0] node1896;
	wire [3-1:0] node1899;
	wire [3-1:0] node1900;
	wire [3-1:0] node1904;
	wire [3-1:0] node1905;
	wire [3-1:0] node1906;
	wire [3-1:0] node1907;
	wire [3-1:0] node1911;
	wire [3-1:0] node1913;
	wire [3-1:0] node1916;
	wire [3-1:0] node1917;
	wire [3-1:0] node1919;
	wire [3-1:0] node1922;
	wire [3-1:0] node1924;
	wire [3-1:0] node1927;
	wire [3-1:0] node1928;
	wire [3-1:0] node1929;
	wire [3-1:0] node1931;
	wire [3-1:0] node1932;
	wire [3-1:0] node1933;
	wire [3-1:0] node1935;
	wire [3-1:0] node1937;
	wire [3-1:0] node1938;
	wire [3-1:0] node1942;
	wire [3-1:0] node1943;
	wire [3-1:0] node1944;
	wire [3-1:0] node1948;
	wire [3-1:0] node1949;
	wire [3-1:0] node1952;
	wire [3-1:0] node1955;
	wire [3-1:0] node1956;
	wire [3-1:0] node1957;
	wire [3-1:0] node1959;
	wire [3-1:0] node1964;
	wire [3-1:0] node1965;
	wire [3-1:0] node1966;
	wire [3-1:0] node1967;
	wire [3-1:0] node1968;
	wire [3-1:0] node1970;
	wire [3-1:0] node1973;
	wire [3-1:0] node1974;
	wire [3-1:0] node1975;
	wire [3-1:0] node1978;
	wire [3-1:0] node1982;
	wire [3-1:0] node1983;
	wire [3-1:0] node1984;
	wire [3-1:0] node1986;
	wire [3-1:0] node1989;
	wire [3-1:0] node1990;
	wire [3-1:0] node1994;
	wire [3-1:0] node1995;
	wire [3-1:0] node1999;
	wire [3-1:0] node2000;
	wire [3-1:0] node2001;
	wire [3-1:0] node2002;
	wire [3-1:0] node2006;
	wire [3-1:0] node2008;
	wire [3-1:0] node2010;
	wire [3-1:0] node2013;
	wire [3-1:0] node2014;
	wire [3-1:0] node2015;
	wire [3-1:0] node2019;
	wire [3-1:0] node2020;
	wire [3-1:0] node2021;
	wire [3-1:0] node2026;
	wire [3-1:0] node2027;
	wire [3-1:0] node2028;
	wire [3-1:0] node2029;
	wire [3-1:0] node2030;
	wire [3-1:0] node2034;
	wire [3-1:0] node2035;
	wire [3-1:0] node2038;
	wire [3-1:0] node2041;
	wire [3-1:0] node2043;
	wire [3-1:0] node2044;
	wire [3-1:0] node2046;
	wire [3-1:0] node2050;
	wire [3-1:0] node2052;
	wire [3-1:0] node2054;
	wire [3-1:0] node2055;
	wire [3-1:0] node2057;
	wire [3-1:0] node2061;
	wire [3-1:0] node2062;
	wire [3-1:0] node2063;
	wire [3-1:0] node2064;
	wire [3-1:0] node2065;
	wire [3-1:0] node2066;
	wire [3-1:0] node2067;
	wire [3-1:0] node2068;
	wire [3-1:0] node2073;
	wire [3-1:0] node2074;
	wire [3-1:0] node2076;
	wire [3-1:0] node2080;
	wire [3-1:0] node2081;
	wire [3-1:0] node2082;
	wire [3-1:0] node2084;
	wire [3-1:0] node2087;
	wire [3-1:0] node2088;
	wire [3-1:0] node2092;
	wire [3-1:0] node2095;
	wire [3-1:0] node2096;
	wire [3-1:0] node2097;
	wire [3-1:0] node2098;
	wire [3-1:0] node2101;
	wire [3-1:0] node2103;
	wire [3-1:0] node2107;
	wire [3-1:0] node2109;
	wire [3-1:0] node2112;
	wire [3-1:0] node2113;
	wire [3-1:0] node2114;
	wire [3-1:0] node2115;
	wire [3-1:0] node2117;
	wire [3-1:0] node2118;
	wire [3-1:0] node2123;
	wire [3-1:0] node2124;
	wire [3-1:0] node2125;
	wire [3-1:0] node2126;
	wire [3-1:0] node2130;
	wire [3-1:0] node2132;
	wire [3-1:0] node2135;
	wire [3-1:0] node2136;
	wire [3-1:0] node2141;
	wire [3-1:0] node2142;
	wire [3-1:0] node2143;
	wire [3-1:0] node2144;
	wire [3-1:0] node2145;
	wire [3-1:0] node2146;
	wire [3-1:0] node2147;
	wire [3-1:0] node2151;
	wire [3-1:0] node2152;
	wire [3-1:0] node2155;
	wire [3-1:0] node2158;
	wire [3-1:0] node2161;
	wire [3-1:0] node2162;
	wire [3-1:0] node2164;
	wire [3-1:0] node2167;
	wire [3-1:0] node2169;
	wire [3-1:0] node2170;
	wire [3-1:0] node2174;
	wire [3-1:0] node2175;
	wire [3-1:0] node2177;
	wire [3-1:0] node2178;
	wire [3-1:0] node2181;
	wire [3-1:0] node2184;
	wire [3-1:0] node2185;
	wire [3-1:0] node2186;
	wire [3-1:0] node2187;
	wire [3-1:0] node2191;
	wire [3-1:0] node2192;
	wire [3-1:0] node2197;
	wire [3-1:0] node2198;
	wire [3-1:0] node2199;
	wire [3-1:0] node2200;
	wire [3-1:0] node2204;
	wire [3-1:0] node2205;
	wire [3-1:0] node2207;
	wire [3-1:0] node2210;
	wire [3-1:0] node2212;
	wire [3-1:0] node2215;
	wire [3-1:0] node2216;
	wire [3-1:0] node2217;
	wire [3-1:0] node2218;
	wire [3-1:0] node2219;
	wire [3-1:0] node2225;
	wire [3-1:0] node2227;
	wire [3-1:0] node2229;
	wire [3-1:0] node2232;
	wire [3-1:0] node2233;
	wire [3-1:0] node2234;
	wire [3-1:0] node2235;
	wire [3-1:0] node2237;
	wire [3-1:0] node2239;
	wire [3-1:0] node2240;
	wire [3-1:0] node2241;
	wire [3-1:0] node2243;
	wire [3-1:0] node2246;
	wire [3-1:0] node2248;
	wire [3-1:0] node2251;
	wire [3-1:0] node2253;
	wire [3-1:0] node2254;
	wire [3-1:0] node2258;
	wire [3-1:0] node2259;
	wire [3-1:0] node2261;
	wire [3-1:0] node2262;
	wire [3-1:0] node2263;
	wire [3-1:0] node2264;
	wire [3-1:0] node2268;
	wire [3-1:0] node2270;
	wire [3-1:0] node2273;
	wire [3-1:0] node2274;
	wire [3-1:0] node2275;
	wire [3-1:0] node2278;
	wire [3-1:0] node2280;
	wire [3-1:0] node2284;
	wire [3-1:0] node2285;
	wire [3-1:0] node2286;
	wire [3-1:0] node2287;
	wire [3-1:0] node2290;
	wire [3-1:0] node2291;
	wire [3-1:0] node2295;
	wire [3-1:0] node2296;
	wire [3-1:0] node2297;
	wire [3-1:0] node2302;
	wire [3-1:0] node2303;
	wire [3-1:0] node2304;
	wire [3-1:0] node2307;
	wire [3-1:0] node2308;
	wire [3-1:0] node2311;
	wire [3-1:0] node2312;
	wire [3-1:0] node2316;
	wire [3-1:0] node2317;
	wire [3-1:0] node2319;
	wire [3-1:0] node2321;
	wire [3-1:0] node2324;
	wire [3-1:0] node2327;
	wire [3-1:0] node2328;
	wire [3-1:0] node2329;
	wire [3-1:0] node2330;
	wire [3-1:0] node2331;
	wire [3-1:0] node2332;
	wire [3-1:0] node2336;
	wire [3-1:0] node2337;
	wire [3-1:0] node2338;
	wire [3-1:0] node2340;
	wire [3-1:0] node2343;
	wire [3-1:0] node2345;
	wire [3-1:0] node2349;
	wire [3-1:0] node2351;
	wire [3-1:0] node2352;
	wire [3-1:0] node2353;
	wire [3-1:0] node2358;
	wire [3-1:0] node2359;
	wire [3-1:0] node2360;
	wire [3-1:0] node2361;
	wire [3-1:0] node2363;
	wire [3-1:0] node2366;
	wire [3-1:0] node2367;
	wire [3-1:0] node2368;
	wire [3-1:0] node2371;
	wire [3-1:0] node2375;
	wire [3-1:0] node2376;
	wire [3-1:0] node2377;
	wire [3-1:0] node2381;
	wire [3-1:0] node2383;
	wire [3-1:0] node2385;
	wire [3-1:0] node2388;
	wire [3-1:0] node2389;
	wire [3-1:0] node2390;
	wire [3-1:0] node2391;
	wire [3-1:0] node2395;
	wire [3-1:0] node2398;
	wire [3-1:0] node2400;
	wire [3-1:0] node2402;
	wire [3-1:0] node2404;
	wire [3-1:0] node2407;
	wire [3-1:0] node2408;
	wire [3-1:0] node2409;
	wire [3-1:0] node2410;
	wire [3-1:0] node2412;
	wire [3-1:0] node2414;
	wire [3-1:0] node2417;
	wire [3-1:0] node2418;
	wire [3-1:0] node2419;
	wire [3-1:0] node2422;
	wire [3-1:0] node2425;
	wire [3-1:0] node2427;
	wire [3-1:0] node2428;
	wire [3-1:0] node2431;
	wire [3-1:0] node2434;
	wire [3-1:0] node2435;
	wire [3-1:0] node2436;
	wire [3-1:0] node2437;
	wire [3-1:0] node2438;
	wire [3-1:0] node2442;
	wire [3-1:0] node2445;
	wire [3-1:0] node2447;
	wire [3-1:0] node2450;
	wire [3-1:0] node2451;
	wire [3-1:0] node2453;
	wire [3-1:0] node2455;
	wire [3-1:0] node2458;
	wire [3-1:0] node2459;
	wire [3-1:0] node2463;
	wire [3-1:0] node2464;
	wire [3-1:0] node2465;
	wire [3-1:0] node2466;
	wire [3-1:0] node2468;
	wire [3-1:0] node2471;
	wire [3-1:0] node2473;
	wire [3-1:0] node2474;
	wire [3-1:0] node2478;
	wire [3-1:0] node2479;
	wire [3-1:0] node2481;
	wire [3-1:0] node2484;
	wire [3-1:0] node2486;
	wire [3-1:0] node2489;
	wire [3-1:0] node2490;
	wire [3-1:0] node2492;
	wire [3-1:0] node2495;
	wire [3-1:0] node2496;
	wire [3-1:0] node2498;
	wire [3-1:0] node2501;
	wire [3-1:0] node2502;
	wire [3-1:0] node2504;
	wire [3-1:0] node2508;
	wire [3-1:0] node2509;
	wire [3-1:0] node2510;
	wire [3-1:0] node2511;
	wire [3-1:0] node2512;
	wire [3-1:0] node2514;
	wire [3-1:0] node2515;
	wire [3-1:0] node2518;
	wire [3-1:0] node2524;
	wire [3-1:0] node2525;
	wire [3-1:0] node2527;
	wire [3-1:0] node2529;
	wire [3-1:0] node2530;
	wire [3-1:0] node2531;
	wire [3-1:0] node2533;
	wire [3-1:0] node2536;
	wire [3-1:0] node2539;
	wire [3-1:0] node2541;
	wire [3-1:0] node2542;
	wire [3-1:0] node2543;
	wire [3-1:0] node2548;
	wire [3-1:0] node2549;
	wire [3-1:0] node2550;
	wire [3-1:0] node2551;
	wire [3-1:0] node2553;
	wire [3-1:0] node2554;
	wire [3-1:0] node2556;
	wire [3-1:0] node2559;
	wire [3-1:0] node2560;
	wire [3-1:0] node2564;
	wire [3-1:0] node2567;
	wire [3-1:0] node2569;
	wire [3-1:0] node2570;
	wire [3-1:0] node2572;
	wire [3-1:0] node2575;
	wire [3-1:0] node2577;
	wire [3-1:0] node2578;
	wire [3-1:0] node2581;
	wire [3-1:0] node2584;
	wire [3-1:0] node2586;
	wire [3-1:0] node2587;
	wire [3-1:0] node2589;
	wire [3-1:0] node2590;
	wire [3-1:0] node2594;
	wire [3-1:0] node2595;
	wire [3-1:0] node2597;
	wire [3-1:0] node2600;
	wire [3-1:0] node2601;

	assign outp = (inp[3]) ? node1502 : node1;
		assign node1 = (inp[4]) ? node619 : node2;
			assign node2 = (inp[9]) ? node242 : node3;
				assign node3 = (inp[7]) ? node179 : node4;
					assign node4 = (inp[1]) ? node92 : node5;
						assign node5 = (inp[5]) ? node57 : node6;
							assign node6 = (inp[0]) ? node44 : node7;
								assign node7 = (inp[6]) ? node23 : node8;
									assign node8 = (inp[2]) ? node18 : node9;
										assign node9 = (inp[8]) ? node13 : node10;
											assign node10 = (inp[10]) ? 3'b001 : 3'b101;
											assign node13 = (inp[11]) ? 3'b001 : node14;
												assign node14 = (inp[10]) ? 3'b101 : 3'b001;
										assign node18 = (inp[11]) ? node20 : 3'b101;
											assign node20 = (inp[10]) ? 3'b001 : 3'b101;
									assign node23 = (inp[11]) ? node35 : node24;
										assign node24 = (inp[10]) ? node30 : node25;
											assign node25 = (inp[8]) ? 3'b001 : node26;
												assign node26 = (inp[2]) ? 3'b101 : 3'b111;
											assign node30 = (inp[8]) ? 3'b111 : node31;
												assign node31 = (inp[2]) ? 3'b111 : 3'b011;
										assign node35 = (inp[2]) ? node41 : node36;
											assign node36 = (inp[8]) ? 3'b011 : node37;
												assign node37 = (inp[10]) ? 3'b011 : 3'b111;
											assign node41 = (inp[8]) ? 3'b001 : 3'b011;
								assign node44 = (inp[11]) ? node52 : node45;
									assign node45 = (inp[2]) ? node49 : node46;
										assign node46 = (inp[8]) ? 3'b111 : 3'b011;
										assign node49 = (inp[8]) ? 3'b011 : 3'b111;
									assign node52 = (inp[8]) ? 3'b111 : node53;
										assign node53 = (inp[2]) ? 3'b111 : 3'b011;
							assign node57 = (inp[0]) ? node83 : node58;
								assign node58 = (inp[6]) ? node70 : node59;
									assign node59 = (inp[11]) ? node63 : node60;
										assign node60 = (inp[10]) ? 3'b001 : 3'b101;
										assign node63 = (inp[10]) ? node65 : 3'b001;
											assign node65 = (inp[2]) ? node67 : 3'b110;
												assign node67 = (inp[8]) ? 3'b101 : 3'b110;
									assign node70 = (inp[10]) ? node76 : node71;
										assign node71 = (inp[11]) ? node73 : 3'b111;
											assign node73 = (inp[8]) ? 3'b111 : 3'b011;
										assign node76 = (inp[11]) ? 3'b101 : node77;
											assign node77 = (inp[8]) ? 3'b011 : node78;
												assign node78 = (inp[2]) ? 3'b011 : 3'b001;
								assign node83 = (inp[8]) ? node87 : node84;
									assign node84 = (inp[2]) ? 3'b101 : 3'b001;
									assign node87 = (inp[2]) ? node89 : 3'b101;
										assign node89 = (inp[11]) ? 3'b101 : 3'b001;
						assign node92 = (inp[0]) ? node148 : node93;
							assign node93 = (inp[2]) ? node121 : node94;
								assign node94 = (inp[11]) ? node112 : node95;
									assign node95 = (inp[5]) ? node105 : node96;
										assign node96 = (inp[10]) ? node100 : node97;
											assign node97 = (inp[6]) ? 3'b001 : 3'b011;
											assign node100 = (inp[8]) ? 3'b011 : node101;
												assign node101 = (inp[6]) ? 3'b011 : 3'b001;
										assign node105 = (inp[8]) ? node109 : node106;
											assign node106 = (inp[6]) ? 3'b011 : 3'b001;
											assign node109 = (inp[10]) ? 3'b101 : 3'b111;
									assign node112 = (inp[5]) ? 3'b001 : node113;
										assign node113 = (inp[10]) ? node117 : node114;
											assign node114 = (inp[6]) ? 3'b101 : 3'b111;
											assign node117 = (inp[6]) ? 3'b111 : 3'b101;
								assign node121 = (inp[6]) ? node133 : node122;
									assign node122 = (inp[5]) ? node126 : node123;
										assign node123 = (inp[10]) ? 3'b011 : 3'b111;
										assign node126 = (inp[10]) ? 3'b001 : node127;
											assign node127 = (inp[11]) ? node129 : 3'b011;
												assign node129 = (inp[8]) ? 3'b011 : 3'b001;
									assign node133 = (inp[8]) ? node139 : node134;
										assign node134 = (inp[11]) ? node136 : 3'b011;
											assign node136 = (inp[5]) ? 3'b011 : 3'b111;
										assign node139 = (inp[11]) ? node145 : node140;
											assign node140 = (inp[5]) ? node142 : 3'b001;
												assign node142 = (inp[10]) ? 3'b111 : 3'b101;
											assign node145 = (inp[5]) ? 3'b011 : 3'b111;
							assign node148 = (inp[6]) ? 3'b111 : node149;
								assign node149 = (inp[5]) ? node167 : node150;
									assign node150 = (inp[10]) ? node160 : node151;
										assign node151 = (inp[11]) ? node155 : node152;
											assign node152 = (inp[8]) ? 3'b011 : 3'b111;
											assign node155 = (inp[8]) ? 3'b111 : node156;
												assign node156 = (inp[2]) ? 3'b111 : 3'b011;
										assign node160 = (inp[2]) ? 3'b111 : node161;
											assign node161 = (inp[8]) ? 3'b111 : node162;
												assign node162 = (inp[11]) ? 3'b011 : 3'b111;
									assign node167 = (inp[11]) ? node173 : node168;
										assign node168 = (inp[2]) ? node170 : 3'b011;
											assign node170 = (inp[8]) ? 3'b111 : 3'b011;
										assign node173 = (inp[2]) ? 3'b011 : node174;
											assign node174 = (inp[8]) ? 3'b011 : 3'b111;
					assign node179 = (inp[5]) ? node205 : node180;
						assign node180 = (inp[2]) ? node190 : node181;
							assign node181 = (inp[6]) ? 3'b111 : node182;
								assign node182 = (inp[1]) ? node184 : 3'b111;
									assign node184 = (inp[11]) ? node186 : 3'b111;
										assign node186 = (inp[8]) ? 3'b111 : 3'b011;
							assign node190 = (inp[11]) ? 3'b111 : node191;
								assign node191 = (inp[8]) ? node193 : 3'b111;
									assign node193 = (inp[0]) ? node199 : node194;
										assign node194 = (inp[1]) ? node196 : 3'b101;
											assign node196 = (inp[6]) ? 3'b101 : 3'b001;
										assign node199 = (inp[6]) ? 3'b111 : node200;
											assign node200 = (inp[1]) ? 3'b011 : 3'b111;
						assign node205 = (inp[0]) ? node229 : node206;
							assign node206 = (inp[11]) ? node216 : node207;
								assign node207 = (inp[1]) ? node209 : 3'b111;
									assign node209 = (inp[6]) ? 3'b111 : node210;
										assign node210 = (inp[2]) ? node212 : 3'b011;
											assign node212 = (inp[8]) ? 3'b111 : 3'b011;
								assign node216 = (inp[2]) ? node224 : node217;
									assign node217 = (inp[8]) ? node219 : 3'b101;
										assign node219 = (inp[1]) ? node221 : 3'b111;
											assign node221 = (inp[6]) ? 3'b111 : 3'b011;
									assign node224 = (inp[6]) ? 3'b111 : node225;
										assign node225 = (inp[1]) ? 3'b011 : 3'b111;
							assign node229 = (inp[1]) ? node231 : 3'b011;
								assign node231 = (inp[6]) ? 3'b111 : node232;
									assign node232 = (inp[10]) ? 3'b011 : node233;
										assign node233 = (inp[2]) ? node235 : 3'b111;
											assign node235 = (inp[8]) ? node237 : 3'b011;
												assign node237 = (inp[11]) ? 3'b011 : 3'b111;
				assign node242 = (inp[6]) ? node422 : node243;
					assign node243 = (inp[0]) ? node331 : node244;
						assign node244 = (inp[10]) ? node286 : node245;
							assign node245 = (inp[1]) ? node269 : node246;
								assign node246 = (inp[7]) ? node258 : node247;
									assign node247 = (inp[5]) ? node255 : node248;
										assign node248 = (inp[8]) ? 3'b001 : node249;
											assign node249 = (inp[11]) ? 3'b110 : node250;
												assign node250 = (inp[2]) ? 3'b001 : 3'b110;
										assign node255 = (inp[11]) ? 3'b010 : 3'b110;
									assign node258 = (inp[11]) ? node260 : 3'b001;
										assign node260 = (inp[5]) ? node264 : node261;
											assign node261 = (inp[8]) ? 3'b101 : 3'b001;
											assign node264 = (inp[2]) ? node266 : 3'b110;
												assign node266 = (inp[8]) ? 3'b001 : 3'b110;
								assign node269 = (inp[11]) ? node275 : node270;
									assign node270 = (inp[5]) ? 3'b001 : node271;
										assign node271 = (inp[8]) ? 3'b101 : 3'b001;
									assign node275 = (inp[5]) ? node283 : node276;
										assign node276 = (inp[7]) ? 3'b101 : node277;
											assign node277 = (inp[2]) ? node279 : 3'b001;
												assign node279 = (inp[8]) ? 3'b101 : 3'b001;
										assign node283 = (inp[7]) ? 3'b001 : 3'b110;
							assign node286 = (inp[5]) ? node314 : node287;
								assign node287 = (inp[11]) ? node305 : node288;
									assign node288 = (inp[2]) ? node296 : node289;
										assign node289 = (inp[8]) ? 3'b001 : node290;
											assign node290 = (inp[7]) ? 3'b110 : node291;
												assign node291 = (inp[1]) ? 3'b110 : 3'b010;
										assign node296 = (inp[7]) ? node300 : node297;
											assign node297 = (inp[1]) ? 3'b001 : 3'b110;
											assign node300 = (inp[1]) ? node302 : 3'b001;
												assign node302 = (inp[8]) ? 3'b101 : 3'b001;
									assign node305 = (inp[1]) ? node309 : node306;
										assign node306 = (inp[7]) ? 3'b110 : 3'b010;
										assign node309 = (inp[7]) ? node311 : 3'b110;
											assign node311 = (inp[2]) ? 3'b001 : 3'b110;
								assign node314 = (inp[7]) ? node324 : node315;
									assign node315 = (inp[1]) ? 3'b010 : node316;
										assign node316 = (inp[8]) ? node318 : 3'b100;
											assign node318 = (inp[11]) ? node320 : 3'b010;
												assign node320 = (inp[2]) ? 3'b010 : 3'b100;
									assign node324 = (inp[11]) ? node326 : 3'b110;
										assign node326 = (inp[1]) ? node328 : 3'b010;
											assign node328 = (inp[2]) ? 3'b110 : 3'b010;
						assign node331 = (inp[10]) ? node379 : node332;
							assign node332 = (inp[5]) ? node362 : node333;
								assign node333 = (inp[1]) ? node349 : node334;
									assign node334 = (inp[2]) ? node342 : node335;
										assign node335 = (inp[7]) ? node339 : node336;
											assign node336 = (inp[8]) ? 3'b101 : 3'b001;
											assign node339 = (inp[8]) ? 3'b011 : 3'b101;
										assign node342 = (inp[7]) ? node346 : node343;
											assign node343 = (inp[11]) ? 3'b101 : 3'b010;
											assign node346 = (inp[11]) ? 3'b011 : 3'b101;
									assign node349 = (inp[7]) ? node355 : node350;
										assign node350 = (inp[11]) ? node352 : 3'b011;
											assign node352 = (inp[2]) ? 3'b011 : 3'b101;
										assign node355 = (inp[11]) ? node357 : 3'b111;
											assign node357 = (inp[2]) ? node359 : 3'b011;
												assign node359 = (inp[8]) ? 3'b111 : 3'b011;
								assign node362 = (inp[8]) ? node370 : node363;
									assign node363 = (inp[7]) ? 3'b101 : node364;
										assign node364 = (inp[1]) ? node366 : 3'b001;
											assign node366 = (inp[2]) ? 3'b101 : 3'b001;
									assign node370 = (inp[11]) ? node372 : 3'b011;
										assign node372 = (inp[1]) ? node374 : 3'b001;
											assign node374 = (inp[2]) ? node376 : 3'b101;
												assign node376 = (inp[7]) ? 3'b011 : 3'b101;
							assign node379 = (inp[5]) ? node401 : node380;
								assign node380 = (inp[1]) ? node388 : node381;
									assign node381 = (inp[7]) ? node383 : 3'b001;
										assign node383 = (inp[2]) ? 3'b011 : node384;
											assign node384 = (inp[8]) ? 3'b101 : 3'b001;
									assign node388 = (inp[8]) ? node394 : node389;
										assign node389 = (inp[11]) ? node391 : 3'b101;
											assign node391 = (inp[7]) ? 3'b101 : 3'b001;
										assign node394 = (inp[7]) ? node396 : 3'b101;
											assign node396 = (inp[2]) ? 3'b011 : node397;
												assign node397 = (inp[11]) ? 3'b101 : 3'b011;
								assign node401 = (inp[7]) ? node411 : node402;
									assign node402 = (inp[1]) ? node404 : 3'b110;
										assign node404 = (inp[11]) ? node406 : 3'b001;
											assign node406 = (inp[8]) ? node408 : 3'b110;
												assign node408 = (inp[2]) ? 3'b001 : 3'b110;
									assign node411 = (inp[1]) ? node415 : node412;
										assign node412 = (inp[8]) ? 3'b001 : 3'b110;
										assign node415 = (inp[11]) ? node417 : 3'b101;
											assign node417 = (inp[2]) ? node419 : 3'b001;
												assign node419 = (inp[8]) ? 3'b101 : 3'b001;
					assign node422 = (inp[0]) ? node536 : node423;
						assign node423 = (inp[7]) ? node479 : node424;
							assign node424 = (inp[10]) ? node444 : node425;
								assign node425 = (inp[5]) ? node435 : node426;
									assign node426 = (inp[1]) ? node428 : 3'b101;
										assign node428 = (inp[8]) ? node432 : node429;
											assign node429 = (inp[2]) ? 3'b011 : 3'b101;
											assign node432 = (inp[11]) ? 3'b011 : 3'b111;
									assign node435 = (inp[1]) ? node437 : 3'b001;
										assign node437 = (inp[8]) ? node439 : 3'b101;
											assign node439 = (inp[11]) ? 3'b101 : node440;
												assign node440 = (inp[2]) ? 3'b001 : 3'b101;
								assign node444 = (inp[5]) ? node458 : node445;
									assign node445 = (inp[1]) ? node451 : node446;
										assign node446 = (inp[2]) ? node448 : 3'b001;
											assign node448 = (inp[8]) ? 3'b101 : 3'b001;
										assign node451 = (inp[2]) ? node455 : node452;
											assign node452 = (inp[8]) ? 3'b101 : 3'b001;
											assign node455 = (inp[8]) ? 3'b011 : 3'b101;
									assign node458 = (inp[1]) ? node468 : node459;
										assign node459 = (inp[11]) ? node465 : node460;
											assign node460 = (inp[8]) ? node462 : 3'b110;
												assign node462 = (inp[2]) ? 3'b010 : 3'b110;
											assign node465 = (inp[2]) ? 3'b110 : 3'b010;
										assign node468 = (inp[8]) ? node474 : node469;
											assign node469 = (inp[2]) ? 3'b001 : node470;
												assign node470 = (inp[11]) ? 3'b110 : 3'b001;
											assign node474 = (inp[11]) ? 3'b001 : node475;
												assign node475 = (inp[2]) ? 3'b101 : 3'b001;
							assign node479 = (inp[1]) ? node513 : node480;
								assign node480 = (inp[5]) ? node496 : node481;
									assign node481 = (inp[10]) ? node489 : node482;
										assign node482 = (inp[2]) ? 3'b011 : node483;
											assign node483 = (inp[11]) ? node485 : 3'b011;
												assign node485 = (inp[8]) ? 3'b011 : 3'b101;
										assign node489 = (inp[2]) ? node493 : node490;
											assign node490 = (inp[8]) ? 3'b101 : 3'b001;
											assign node493 = (inp[8]) ? 3'b011 : 3'b101;
									assign node496 = (inp[10]) ? node506 : node497;
										assign node497 = (inp[2]) ? node501 : node498;
											assign node498 = (inp[11]) ? 3'b001 : 3'b101;
											assign node501 = (inp[8]) ? node503 : 3'b101;
												assign node503 = (inp[11]) ? 3'b101 : 3'b011;
										assign node506 = (inp[11]) ? node508 : 3'b001;
											assign node508 = (inp[8]) ? 3'b001 : node509;
												assign node509 = (inp[2]) ? 3'b001 : 3'b110;
								assign node513 = (inp[10]) ? node529 : node514;
									assign node514 = (inp[5]) ? node524 : node515;
										assign node515 = (inp[8]) ? node519 : node516;
											assign node516 = (inp[2]) ? 3'b111 : 3'b011;
											assign node519 = (inp[11]) ? 3'b111 : node520;
												assign node520 = (inp[2]) ? 3'b001 : 3'b111;
										assign node524 = (inp[11]) ? 3'b011 : node525;
											assign node525 = (inp[2]) ? 3'b111 : 3'b011;
									assign node529 = (inp[11]) ? node531 : 3'b011;
										assign node531 = (inp[5]) ? 3'b001 : node532;
											assign node532 = (inp[8]) ? 3'b011 : 3'b101;
						assign node536 = (inp[5]) ? node566 : node537;
							assign node537 = (inp[11]) ? node553 : node538;
								assign node538 = (inp[8]) ? 3'b111 : node539;
									assign node539 = (inp[2]) ? 3'b111 : node540;
										assign node540 = (inp[1]) ? node546 : node541;
											assign node541 = (inp[10]) ? node543 : 3'b011;
												assign node543 = (inp[7]) ? 3'b011 : 3'b101;
											assign node546 = (inp[10]) ? node548 : 3'b111;
												assign node548 = (inp[7]) ? 3'b111 : 3'b011;
								assign node553 = (inp[7]) ? node561 : node554;
									assign node554 = (inp[8]) ? node556 : 3'b011;
										assign node556 = (inp[1]) ? node558 : 3'b011;
											assign node558 = (inp[2]) ? 3'b111 : 3'b011;
									assign node561 = (inp[10]) ? node563 : 3'b111;
										assign node563 = (inp[1]) ? 3'b111 : 3'b011;
							assign node566 = (inp[10]) ? node586 : node567;
								assign node567 = (inp[1]) ? node581 : node568;
									assign node568 = (inp[7]) ? node574 : node569;
										assign node569 = (inp[2]) ? 3'b011 : node570;
											assign node570 = (inp[11]) ? 3'b101 : 3'b011;
										assign node574 = (inp[2]) ? 3'b111 : node575;
											assign node575 = (inp[11]) ? 3'b011 : node576;
												assign node576 = (inp[8]) ? 3'b111 : 3'b011;
									assign node581 = (inp[11]) ? node583 : 3'b111;
										assign node583 = (inp[7]) ? 3'b111 : 3'b011;
								assign node586 = (inp[7]) ? node606 : node587;
									assign node587 = (inp[1]) ? node599 : node588;
										assign node588 = (inp[11]) ? node594 : node589;
											assign node589 = (inp[2]) ? 3'b101 : node590;
												assign node590 = (inp[8]) ? 3'b101 : 3'b001;
											assign node594 = (inp[8]) ? node596 : 3'b001;
												assign node596 = (inp[2]) ? 3'b101 : 3'b001;
										assign node599 = (inp[11]) ? 3'b101 : node600;
											assign node600 = (inp[2]) ? 3'b011 : node601;
												assign node601 = (inp[8]) ? 3'b011 : 3'b101;
									assign node606 = (inp[11]) ? node612 : node607;
										assign node607 = (inp[8]) ? node609 : 3'b011;
											assign node609 = (inp[1]) ? 3'b111 : 3'b011;
										assign node612 = (inp[8]) ? node614 : 3'b101;
											assign node614 = (inp[2]) ? 3'b011 : node615;
												assign node615 = (inp[1]) ? 3'b011 : 3'b101;
			assign node619 = (inp[0]) ? node1067 : node620;
				assign node620 = (inp[11]) ? node830 : node621;
					assign node621 = (inp[9]) ? node727 : node622;
						assign node622 = (inp[7]) ? node658 : node623;
							assign node623 = (inp[5]) ? node637 : node624;
								assign node624 = (inp[1]) ? node634 : node625;
									assign node625 = (inp[10]) ? node631 : node626;
										assign node626 = (inp[6]) ? 3'b011 : node627;
											assign node627 = (inp[2]) ? 3'b001 : 3'b100;
										assign node631 = (inp[6]) ? 3'b101 : 3'b110;
									assign node634 = (inp[10]) ? 3'b001 : 3'b101;
								assign node637 = (inp[1]) ? node649 : node638;
									assign node638 = (inp[10]) ? node642 : node639;
										assign node639 = (inp[6]) ? 3'b101 : 3'b110;
										assign node642 = (inp[6]) ? 3'b000 : node643;
											assign node643 = (inp[8]) ? 3'b010 : node644;
												assign node644 = (inp[2]) ? 3'b010 : 3'b100;
									assign node649 = (inp[10]) ? node655 : node650;
										assign node650 = (inp[2]) ? 3'b010 : node651;
											assign node651 = (inp[8]) ? 3'b010 : 3'b110;
										assign node655 = (inp[8]) ? 3'b110 : 3'b010;
							assign node658 = (inp[1]) ? node690 : node659;
								assign node659 = (inp[2]) ? node671 : node660;
									assign node660 = (inp[5]) ? node662 : 3'b101;
										assign node662 = (inp[10]) ? node668 : node663;
											assign node663 = (inp[6]) ? 3'b101 : node664;
												assign node664 = (inp[8]) ? 3'b001 : 3'b101;
											assign node668 = (inp[6]) ? 3'b001 : 3'b101;
									assign node671 = (inp[6]) ? node679 : node672;
										assign node672 = (inp[10]) ? node676 : node673;
											assign node673 = (inp[5]) ? 3'b001 : 3'b101;
											assign node676 = (inp[5]) ? 3'b101 : 3'b001;
										assign node679 = (inp[10]) ? node685 : node680;
											assign node680 = (inp[5]) ? node682 : 3'b101;
												assign node682 = (inp[8]) ? 3'b001 : 3'b101;
											assign node685 = (inp[8]) ? 3'b001 : node686;
												assign node686 = (inp[5]) ? 3'b001 : 3'b101;
								assign node690 = (inp[8]) ? node710 : node691;
									assign node691 = (inp[10]) ? node701 : node692;
										assign node692 = (inp[5]) ? node696 : node693;
											assign node693 = (inp[6]) ? 3'b000 : 3'b100;
											assign node696 = (inp[2]) ? 3'b001 : node697;
												assign node697 = (inp[6]) ? 3'b001 : 3'b000;
										assign node701 = (inp[5]) ? node707 : node702;
											assign node702 = (inp[6]) ? 3'b011 : node703;
												assign node703 = (inp[2]) ? 3'b001 : 3'b000;
											assign node707 = (inp[6]) ? 3'b101 : 3'b110;
									assign node710 = (inp[6]) ? node724 : node711;
										assign node711 = (inp[2]) ? node717 : node712;
											assign node712 = (inp[5]) ? 3'b001 : node713;
												assign node713 = (inp[10]) ? 3'b001 : 3'b100;
											assign node717 = (inp[5]) ? node721 : node718;
												assign node718 = (inp[10]) ? 3'b111 : 3'b110;
												assign node721 = (inp[10]) ? 3'b000 : 3'b111;
										assign node724 = (inp[5]) ? 3'b111 : 3'b110;
						assign node727 = (inp[6]) ? node779 : node728;
							assign node728 = (inp[10]) ? node754 : node729;
								assign node729 = (inp[5]) ? node747 : node730;
									assign node730 = (inp[7]) ? node738 : node731;
										assign node731 = (inp[1]) ? 3'b010 : node732;
											assign node732 = (inp[8]) ? 3'b010 : node733;
												assign node733 = (inp[2]) ? 3'b010 : 3'b100;
										assign node738 = (inp[1]) ? node740 : 3'b100;
											assign node740 = (inp[2]) ? node744 : node741;
												assign node741 = (inp[8]) ? 3'b110 : 3'b010;
												assign node744 = (inp[8]) ? 3'b001 : 3'b110;
									assign node747 = (inp[7]) ? node749 : 3'b100;
										assign node749 = (inp[2]) ? node751 : 3'b010;
											assign node751 = (inp[8]) ? 3'b100 : 3'b010;
								assign node754 = (inp[8]) ? node766 : node755;
									assign node755 = (inp[5]) ? node761 : node756;
										assign node756 = (inp[2]) ? 3'b100 : node757;
											assign node757 = (inp[7]) ? 3'b100 : 3'b000;
										assign node761 = (inp[7]) ? node763 : 3'b000;
											assign node763 = (inp[1]) ? 3'b100 : 3'b000;
									assign node766 = (inp[5]) ? node772 : node767;
										assign node767 = (inp[2]) ? node769 : 3'b010;
											assign node769 = (inp[7]) ? 3'b100 : 3'b010;
										assign node772 = (inp[1]) ? node774 : 3'b000;
											assign node774 = (inp[7]) ? node776 : 3'b100;
												assign node776 = (inp[2]) ? 3'b010 : 3'b100;
							assign node779 = (inp[7]) ? node805 : node780;
								assign node780 = (inp[5]) ? node792 : node781;
									assign node781 = (inp[10]) ? node787 : node782;
										assign node782 = (inp[1]) ? node784 : 3'b110;
											assign node784 = (inp[8]) ? 3'b001 : 3'b111;
										assign node787 = (inp[1]) ? 3'b110 : node788;
											assign node788 = (inp[2]) ? 3'b110 : 3'b010;
									assign node792 = (inp[1]) ? node800 : node793;
										assign node793 = (inp[10]) ? node795 : 3'b010;
											assign node795 = (inp[8]) ? node797 : 3'b100;
												assign node797 = (inp[2]) ? 3'b000 : 3'b100;
										assign node800 = (inp[10]) ? 3'b010 : node801;
											assign node801 = (inp[8]) ? 3'b000 : 3'b110;
								assign node805 = (inp[5]) ? node817 : node806;
									assign node806 = (inp[1]) ? node812 : node807;
										assign node807 = (inp[2]) ? 3'b001 : node808;
											assign node808 = (inp[10]) ? 3'b110 : 3'b011;
										assign node812 = (inp[10]) ? 3'b001 : node813;
											assign node813 = (inp[8]) ? 3'b101 : 3'b001;
									assign node817 = (inp[10]) ? node825 : node818;
										assign node818 = (inp[1]) ? 3'b001 : node819;
											assign node819 = (inp[2]) ? node821 : 3'b110;
												assign node821 = (inp[8]) ? 3'b001 : 3'b110;
										assign node825 = (inp[8]) ? 3'b110 : node826;
											assign node826 = (inp[1]) ? 3'b110 : 3'b010;
					assign node830 = (inp[9]) ? node966 : node831;
						assign node831 = (inp[6]) ? node891 : node832;
							assign node832 = (inp[7]) ? node862 : node833;
								assign node833 = (inp[2]) ? node847 : node834;
									assign node834 = (inp[8]) ? 3'b010 : node835;
										assign node835 = (inp[5]) ? node843 : node836;
											assign node836 = (inp[1]) ? node840 : node837;
												assign node837 = (inp[10]) ? 3'b010 : 3'b110;
												assign node840 = (inp[10]) ? 3'b110 : 3'b010;
											assign node843 = (inp[10]) ? 3'b100 : 3'b010;
									assign node847 = (inp[5]) ? node857 : node848;
										assign node848 = (inp[10]) ? 3'b110 : node849;
											assign node849 = (inp[8]) ? node853 : node850;
												assign node850 = (inp[1]) ? 3'b010 : 3'b110;
												assign node853 = (inp[1]) ? 3'b110 : 3'b011;
										assign node857 = (inp[10]) ? 3'b010 : node858;
											assign node858 = (inp[1]) ? 3'b110 : 3'b010;
								assign node862 = (inp[1]) ? node882 : node863;
									assign node863 = (inp[5]) ? node875 : node864;
										assign node864 = (inp[10]) ? node870 : node865;
											assign node865 = (inp[8]) ? node867 : 3'b010;
												assign node867 = (inp[2]) ? 3'b110 : 3'b010;
											assign node870 = (inp[8]) ? node872 : 3'b110;
												assign node872 = (inp[2]) ? 3'b010 : 3'b110;
										assign node875 = (inp[2]) ? node877 : 3'b110;
											assign node877 = (inp[8]) ? node879 : 3'b110;
												assign node879 = (inp[10]) ? 3'b110 : 3'b010;
									assign node882 = (inp[10]) ? 3'b110 : node883;
										assign node883 = (inp[5]) ? 3'b000 : node884;
											assign node884 = (inp[2]) ? node886 : 3'b101;
												assign node886 = (inp[8]) ? 3'b100 : 3'b101;
							assign node891 = (inp[2]) ? node927 : node892;
								assign node892 = (inp[10]) ? node914 : node893;
									assign node893 = (inp[5]) ? node903 : node894;
										assign node894 = (inp[7]) ? node896 : 3'b010;
											assign node896 = (inp[1]) ? node900 : node897;
												assign node897 = (inp[8]) ? 3'b010 : 3'b110;
												assign node900 = (inp[8]) ? 3'b100 : 3'b000;
										assign node903 = (inp[7]) ? node909 : node904;
											assign node904 = (inp[1]) ? 3'b110 : node905;
												assign node905 = (inp[8]) ? 3'b001 : 3'b000;
											assign node909 = (inp[1]) ? node911 : 3'b110;
												assign node911 = (inp[8]) ? 3'b101 : 3'b001;
									assign node914 = (inp[8]) ? node920 : node915;
										assign node915 = (inp[5]) ? 3'b000 : node916;
											assign node916 = (inp[7]) ? 3'b010 : 3'b000;
										assign node920 = (inp[7]) ? node924 : node921;
											assign node921 = (inp[1]) ? 3'b110 : 3'b001;
											assign node924 = (inp[1]) ? 3'b001 : 3'b010;
								assign node927 = (inp[8]) ? node949 : node928;
									assign node928 = (inp[7]) ? node942 : node929;
										assign node929 = (inp[1]) ? node937 : node930;
											assign node930 = (inp[5]) ? node934 : node931;
												assign node931 = (inp[10]) ? 3'b001 : 3'b101;
												assign node934 = (inp[10]) ? 3'b110 : 3'b001;
											assign node937 = (inp[5]) ? 3'b110 : node938;
												assign node938 = (inp[10]) ? 3'b110 : 3'b010;
										assign node942 = (inp[1]) ? 3'b001 : node943;
											assign node943 = (inp[5]) ? 3'b010 : node944;
												assign node944 = (inp[10]) ? 3'b110 : 3'b010;
									assign node949 = (inp[1]) ? node957 : node950;
										assign node950 = (inp[7]) ? 3'b110 : node951;
											assign node951 = (inp[5]) ? 3'b101 : node952;
												assign node952 = (inp[10]) ? 3'b101 : 3'b011;
										assign node957 = (inp[7]) ? node961 : node958;
											assign node958 = (inp[5]) ? 3'b010 : 3'b110;
											assign node961 = (inp[10]) ? 3'b011 : node962;
												assign node962 = (inp[5]) ? 3'b111 : 3'b110;
						assign node966 = (inp[6]) ? node1010 : node967;
							assign node967 = (inp[10]) ? node991 : node968;
								assign node968 = (inp[5]) ? node980 : node969;
									assign node969 = (inp[7]) ? node973 : node970;
										assign node970 = (inp[1]) ? 3'b010 : 3'b100;
										assign node973 = (inp[1]) ? node975 : 3'b010;
											assign node975 = (inp[8]) ? 3'b110 : node976;
												assign node976 = (inp[2]) ? 3'b110 : 3'b010;
									assign node980 = (inp[1]) ? node988 : node981;
										assign node981 = (inp[7]) ? 3'b100 : node982;
											assign node982 = (inp[2]) ? node984 : 3'b000;
												assign node984 = (inp[8]) ? 3'b100 : 3'b000;
										assign node988 = (inp[7]) ? 3'b010 : 3'b100;
								assign node991 = (inp[5]) ? node1003 : node992;
									assign node992 = (inp[1]) ? node998 : node993;
										assign node993 = (inp[7]) ? 3'b100 : node994;
											assign node994 = (inp[2]) ? 3'b100 : 3'b000;
										assign node998 = (inp[7]) ? 3'b010 : node999;
											assign node999 = (inp[8]) ? 3'b100 : 3'b000;
									assign node1003 = (inp[7]) ? node1005 : 3'b000;
										assign node1005 = (inp[1]) ? node1007 : 3'b000;
											assign node1007 = (inp[2]) ? 3'b100 : 3'b000;
							assign node1010 = (inp[5]) ? node1038 : node1011;
								assign node1011 = (inp[10]) ? node1025 : node1012;
									assign node1012 = (inp[7]) ? node1020 : node1013;
										assign node1013 = (inp[1]) ? node1017 : node1014;
											assign node1014 = (inp[8]) ? 3'b110 : 3'b010;
											assign node1017 = (inp[8]) ? 3'b001 : 3'b111;
										assign node1020 = (inp[1]) ? node1022 : 3'b001;
											assign node1022 = (inp[8]) ? 3'b101 : 3'b010;
									assign node1025 = (inp[1]) ? node1031 : node1026;
										assign node1026 = (inp[2]) ? node1028 : 3'b010;
											assign node1028 = (inp[7]) ? 3'b110 : 3'b010;
										assign node1031 = (inp[8]) ? node1033 : 3'b110;
											assign node1033 = (inp[2]) ? node1035 : 3'b110;
												assign node1035 = (inp[7]) ? 3'b001 : 3'b110;
								assign node1038 = (inp[7]) ? node1056 : node1039;
									assign node1039 = (inp[8]) ? node1049 : node1040;
										assign node1040 = (inp[10]) ? node1044 : node1041;
											assign node1041 = (inp[1]) ? 3'b110 : 3'b100;
											assign node1044 = (inp[2]) ? 3'b100 : node1045;
												assign node1045 = (inp[1]) ? 3'b100 : 3'b000;
										assign node1049 = (inp[10]) ? node1053 : node1050;
											assign node1050 = (inp[1]) ? 3'b000 : 3'b010;
											assign node1053 = (inp[1]) ? 3'b010 : 3'b100;
									assign node1056 = (inp[10]) ? node1058 : 3'b110;
										assign node1058 = (inp[1]) ? node1062 : node1059;
											assign node1059 = (inp[8]) ? 3'b010 : 3'b100;
											assign node1062 = (inp[8]) ? node1064 : 3'b010;
												assign node1064 = (inp[2]) ? 3'b110 : 3'b010;
				assign node1067 = (inp[9]) ? node1289 : node1068;
					assign node1068 = (inp[7]) ? node1198 : node1069;
						assign node1069 = (inp[1]) ? node1137 : node1070;
							assign node1070 = (inp[5]) ? node1104 : node1071;
								assign node1071 = (inp[6]) ? node1083 : node1072;
									assign node1072 = (inp[10]) ? node1078 : node1073;
										assign node1073 = (inp[2]) ? 3'b101 : node1074;
											assign node1074 = (inp[8]) ? 3'b101 : 3'b001;
										assign node1078 = (inp[11]) ? 3'b001 : node1079;
											assign node1079 = (inp[2]) ? 3'b111 : 3'b001;
									assign node1083 = (inp[11]) ? node1093 : node1084;
										assign node1084 = (inp[8]) ? node1088 : node1085;
											assign node1085 = (inp[2]) ? 3'b000 : 3'b001;
											assign node1088 = (inp[10]) ? node1090 : 3'b110;
												assign node1090 = (inp[2]) ? 3'b010 : 3'b000;
										assign node1093 = (inp[2]) ? node1097 : node1094;
											assign node1094 = (inp[8]) ? 3'b101 : 3'b111;
											assign node1097 = (inp[8]) ? node1101 : node1098;
												assign node1098 = (inp[10]) ? 3'b101 : 3'b001;
												assign node1101 = (inp[10]) ? 3'b000 : 3'b100;
								assign node1104 = (inp[6]) ? node1118 : node1105;
									assign node1105 = (inp[10]) ? node1113 : node1106;
										assign node1106 = (inp[8]) ? node1108 : 3'b000;
											assign node1108 = (inp[11]) ? 3'b011 : node1109;
												assign node1109 = (inp[2]) ? 3'b101 : 3'b011;
										assign node1113 = (inp[8]) ? node1115 : 3'b110;
											assign node1115 = (inp[2]) ? 3'b000 : 3'b110;
									assign node1118 = (inp[8]) ? node1128 : node1119;
										assign node1119 = (inp[2]) ? node1123 : node1120;
											assign node1120 = (inp[11]) ? 3'b101 : 3'b111;
											assign node1123 = (inp[11]) ? 3'b011 : node1124;
												assign node1124 = (inp[10]) ? 3'b111 : 3'b011;
										assign node1128 = (inp[11]) ? node1130 : 3'b011;
											assign node1130 = (inp[10]) ? node1134 : node1131;
												assign node1131 = (inp[2]) ? 3'b011 : 3'b111;
												assign node1134 = (inp[2]) ? 3'b111 : 3'b011;
							assign node1137 = (inp[10]) ? node1163 : node1138;
								assign node1138 = (inp[5]) ? node1156 : node1139;
									assign node1139 = (inp[6]) ? node1149 : node1140;
										assign node1140 = (inp[2]) ? node1144 : node1141;
											assign node1141 = (inp[11]) ? 3'b001 : 3'b101;
											assign node1144 = (inp[11]) ? 3'b101 : node1145;
												assign node1145 = (inp[8]) ? 3'b001 : 3'b101;
										assign node1149 = (inp[11]) ? node1151 : 3'b101;
											assign node1151 = (inp[8]) ? 3'b011 : node1152;
												assign node1152 = (inp[2]) ? 3'b011 : 3'b101;
									assign node1156 = (inp[6]) ? 3'b101 : node1157;
										assign node1157 = (inp[2]) ? node1159 : 3'b100;
											assign node1159 = (inp[8]) ? 3'b001 : 3'b100;
								assign node1163 = (inp[2]) ? node1183 : node1164;
									assign node1164 = (inp[8]) ? node1172 : node1165;
										assign node1165 = (inp[6]) ? 3'b101 : node1166;
											assign node1166 = (inp[5]) ? 3'b000 : node1167;
												assign node1167 = (inp[11]) ? 3'b001 : 3'b101;
										assign node1172 = (inp[5]) ? node1178 : node1173;
											assign node1173 = (inp[6]) ? 3'b011 : node1174;
												assign node1174 = (inp[11]) ? 3'b101 : 3'b111;
											assign node1178 = (inp[6]) ? 3'b101 : node1179;
												assign node1179 = (inp[11]) ? 3'b110 : 3'b001;
									assign node1183 = (inp[6]) ? node1189 : node1184;
										assign node1184 = (inp[5]) ? node1186 : 3'b101;
											assign node1186 = (inp[11]) ? 3'b011 : 3'b001;
										assign node1189 = (inp[5]) ? node1195 : node1190;
											assign node1190 = (inp[8]) ? node1192 : 3'b011;
												assign node1192 = (inp[11]) ? 3'b011 : 3'b101;
											assign node1195 = (inp[11]) ? 3'b101 : 3'b011;
						assign node1198 = (inp[5]) ? node1254 : node1199;
							assign node1199 = (inp[6]) ? node1227 : node1200;
								assign node1200 = (inp[10]) ? node1212 : node1201;
									assign node1201 = (inp[11]) ? node1205 : node1202;
										assign node1202 = (inp[1]) ? 3'b111 : 3'b011;
										assign node1205 = (inp[2]) ? 3'b011 : node1206;
											assign node1206 = (inp[1]) ? node1208 : 3'b100;
												assign node1208 = (inp[8]) ? 3'b011 : 3'b001;
									assign node1212 = (inp[11]) ? node1224 : node1213;
										assign node1213 = (inp[1]) ? node1219 : node1214;
											assign node1214 = (inp[2]) ? node1216 : 3'b111;
												assign node1216 = (inp[8]) ? 3'b001 : 3'b111;
											assign node1219 = (inp[2]) ? 3'b011 : node1220;
												assign node1220 = (inp[8]) ? 3'b011 : 3'b001;
										assign node1224 = (inp[1]) ? 3'b101 : 3'b111;
								assign node1227 = (inp[10]) ? node1239 : node1228;
									assign node1228 = (inp[1]) ? node1236 : node1229;
										assign node1229 = (inp[8]) ? node1231 : 3'b111;
											assign node1231 = (inp[2]) ? node1233 : 3'b011;
												assign node1233 = (inp[11]) ? 3'b011 : 3'b001;
										assign node1236 = (inp[11]) ? 3'b001 : 3'b101;
									assign node1239 = (inp[1]) ? node1247 : node1240;
										assign node1240 = (inp[11]) ? node1242 : 3'b101;
											assign node1242 = (inp[8]) ? 3'b011 : node1243;
												assign node1243 = (inp[2]) ? 3'b011 : 3'b000;
										assign node1247 = (inp[11]) ? 3'b111 : node1248;
											assign node1248 = (inp[8]) ? node1250 : 3'b011;
												assign node1250 = (inp[2]) ? 3'b001 : 3'b011;
							assign node1254 = (inp[10]) ? node1274 : node1255;
								assign node1255 = (inp[1]) ? node1265 : node1256;
									assign node1256 = (inp[6]) ? node1258 : 3'b101;
										assign node1258 = (inp[11]) ? node1262 : node1259;
											assign node1259 = (inp[8]) ? 3'b111 : 3'b101;
											assign node1262 = (inp[8]) ? 3'b001 : 3'b010;
									assign node1265 = (inp[6]) ? 3'b111 : node1266;
										assign node1266 = (inp[11]) ? node1268 : 3'b011;
											assign node1268 = (inp[8]) ? node1270 : 3'b101;
												assign node1270 = (inp[2]) ? 3'b011 : 3'b111;
								assign node1274 = (inp[1]) ? node1282 : node1275;
									assign node1275 = (inp[2]) ? node1277 : 3'b001;
										assign node1277 = (inp[11]) ? 3'b001 : node1278;
											assign node1278 = (inp[8]) ? 3'b011 : 3'b001;
									assign node1282 = (inp[11]) ? node1286 : node1283;
										assign node1283 = (inp[6]) ? 3'b111 : 3'b101;
										assign node1286 = (inp[8]) ? 3'b101 : 3'b001;
					assign node1289 = (inp[6]) ? node1397 : node1290;
						assign node1290 = (inp[10]) ? node1342 : node1291;
							assign node1291 = (inp[1]) ? node1319 : node1292;
								assign node1292 = (inp[5]) ? node1308 : node1293;
									assign node1293 = (inp[7]) ? node1301 : node1294;
										assign node1294 = (inp[2]) ? node1296 : 3'b110;
											assign node1296 = (inp[8]) ? node1298 : 3'b110;
												assign node1298 = (inp[11]) ? 3'b110 : 3'b001;
										assign node1301 = (inp[8]) ? 3'b110 : node1302;
											assign node1302 = (inp[2]) ? 3'b001 : node1303;
												assign node1303 = (inp[11]) ? 3'b110 : 3'b011;
									assign node1308 = (inp[7]) ? node1310 : 3'b010;
										assign node1310 = (inp[8]) ? node1316 : node1311;
											assign node1311 = (inp[11]) ? node1313 : 3'b110;
												assign node1313 = (inp[2]) ? 3'b110 : 3'b010;
											assign node1316 = (inp[11]) ? 3'b110 : 3'b001;
								assign node1319 = (inp[7]) ? node1327 : node1320;
									assign node1320 = (inp[11]) ? node1324 : node1321;
										assign node1321 = (inp[5]) ? 3'b110 : 3'b001;
										assign node1324 = (inp[5]) ? 3'b010 : 3'b110;
									assign node1327 = (inp[2]) ? node1335 : node1328;
										assign node1328 = (inp[11]) ? node1330 : 3'b001;
											assign node1330 = (inp[8]) ? node1332 : 3'b110;
												assign node1332 = (inp[5]) ? 3'b101 : 3'b001;
										assign node1335 = (inp[5]) ? node1337 : 3'b101;
											assign node1337 = (inp[8]) ? 3'b001 : node1338;
												assign node1338 = (inp[11]) ? 3'b101 : 3'b001;
							assign node1342 = (inp[5]) ? node1368 : node1343;
								assign node1343 = (inp[7]) ? node1355 : node1344;
									assign node1344 = (inp[2]) ? node1352 : node1345;
										assign node1345 = (inp[8]) ? 3'b010 : node1346;
											assign node1346 = (inp[11]) ? node1348 : 3'b010;
												assign node1348 = (inp[1]) ? 3'b010 : 3'b100;
										assign node1352 = (inp[11]) ? 3'b010 : 3'b110;
									assign node1355 = (inp[11]) ? node1361 : node1356;
										assign node1356 = (inp[1]) ? node1358 : 3'b110;
											assign node1358 = (inp[2]) ? 3'b001 : 3'b110;
										assign node1361 = (inp[1]) ? 3'b110 : node1362;
											assign node1362 = (inp[8]) ? node1364 : 3'b010;
												assign node1364 = (inp[2]) ? 3'b110 : 3'b010;
								assign node1368 = (inp[1]) ? node1380 : node1369;
									assign node1369 = (inp[8]) ? 3'b100 : node1370;
										assign node1370 = (inp[11]) ? node1376 : node1371;
											assign node1371 = (inp[2]) ? node1373 : 3'b100;
												assign node1373 = (inp[7]) ? 3'b010 : 3'b100;
											assign node1376 = (inp[7]) ? 3'b100 : 3'b000;
									assign node1380 = (inp[11]) ? node1388 : node1381;
										assign node1381 = (inp[7]) ? node1383 : 3'b010;
											assign node1383 = (inp[2]) ? 3'b110 : node1384;
												assign node1384 = (inp[8]) ? 3'b110 : 3'b010;
										assign node1388 = (inp[2]) ? node1390 : 3'b100;
											assign node1390 = (inp[7]) ? node1394 : node1391;
												assign node1391 = (inp[8]) ? 3'b010 : 3'b100;
												assign node1394 = (inp[8]) ? 3'b110 : 3'b010;
						assign node1397 = (inp[10]) ? node1449 : node1398;
							assign node1398 = (inp[5]) ? node1428 : node1399;
								assign node1399 = (inp[8]) ? node1417 : node1400;
									assign node1400 = (inp[1]) ? node1410 : node1401;
										assign node1401 = (inp[7]) ? 3'b101 : node1402;
											assign node1402 = (inp[11]) ? node1406 : node1403;
												assign node1403 = (inp[2]) ? 3'b101 : 3'b011;
												assign node1406 = (inp[2]) ? 3'b011 : 3'b010;
										assign node1410 = (inp[7]) ? 3'b011 : node1411;
											assign node1411 = (inp[11]) ? 3'b101 : node1412;
												assign node1412 = (inp[2]) ? 3'b011 : 3'b001;
									assign node1417 = (inp[1]) ? node1419 : 3'b011;
										assign node1419 = (inp[2]) ? 3'b111 : node1420;
											assign node1420 = (inp[7]) ? node1424 : node1421;
												assign node1421 = (inp[11]) ? 3'b101 : 3'b011;
												assign node1424 = (inp[11]) ? 3'b011 : 3'b111;
								assign node1428 = (inp[7]) ? node1440 : node1429;
									assign node1429 = (inp[1]) ? node1437 : node1430;
										assign node1430 = (inp[11]) ? node1432 : 3'b011;
											assign node1432 = (inp[2]) ? node1434 : 3'b110;
												assign node1434 = (inp[8]) ? 3'b011 : 3'b111;
										assign node1437 = (inp[11]) ? 3'b001 : 3'b101;
									assign node1440 = (inp[8]) ? 3'b101 : node1441;
										assign node1441 = (inp[1]) ? node1443 : 3'b001;
											assign node1443 = (inp[11]) ? node1445 : 3'b101;
												assign node1445 = (inp[2]) ? 3'b101 : 3'b001;
							assign node1449 = (inp[5]) ? node1473 : node1450;
								assign node1450 = (inp[1]) ? node1460 : node1451;
									assign node1451 = (inp[2]) ? node1457 : node1452;
										assign node1452 = (inp[7]) ? 3'b001 : node1453;
											assign node1453 = (inp[8]) ? 3'b001 : 3'b110;
										assign node1457 = (inp[7]) ? 3'b101 : 3'b001;
									assign node1460 = (inp[11]) ? node1466 : node1461;
										assign node1461 = (inp[8]) ? node1463 : 3'b101;
											assign node1463 = (inp[7]) ? 3'b101 : 3'b100;
										assign node1466 = (inp[7]) ? node1468 : 3'b001;
											assign node1468 = (inp[8]) ? 3'b101 : node1469;
												assign node1469 = (inp[2]) ? 3'b101 : 3'b001;
								assign node1473 = (inp[1]) ? node1491 : node1474;
									assign node1474 = (inp[11]) ? node1486 : node1475;
										assign node1475 = (inp[7]) ? node1481 : node1476;
											assign node1476 = (inp[8]) ? 3'b110 : node1477;
												assign node1477 = (inp[2]) ? 3'b110 : 3'b010;
											assign node1481 = (inp[8]) ? 3'b001 : node1482;
												assign node1482 = (inp[2]) ? 3'b000 : 3'b010;
										assign node1486 = (inp[7]) ? 3'b110 : node1487;
											assign node1487 = (inp[2]) ? 3'b110 : 3'b010;
									assign node1491 = (inp[11]) ? node1499 : node1492;
										assign node1492 = (inp[8]) ? 3'b001 : node1493;
											assign node1493 = (inp[2]) ? 3'b001 : node1494;
												assign node1494 = (inp[7]) ? 3'b001 : 3'b111;
										assign node1499 = (inp[7]) ? 3'b001 : 3'b110;
		assign node1502 = (inp[4]) ? node2232 : node1503;
			assign node1503 = (inp[9]) ? node1927 : node1504;
				assign node1504 = (inp[0]) ? node1714 : node1505;
					assign node1505 = (inp[1]) ? node1613 : node1506;
						assign node1506 = (inp[7]) ? node1574 : node1507;
							assign node1507 = (inp[10]) ? node1537 : node1508;
								assign node1508 = (inp[5]) ? node1524 : node1509;
									assign node1509 = (inp[2]) ? node1517 : node1510;
										assign node1510 = (inp[11]) ? node1512 : 3'b100;
											assign node1512 = (inp[8]) ? 3'b100 : node1513;
												assign node1513 = (inp[6]) ? 3'b000 : 3'b100;
										assign node1517 = (inp[11]) ? 3'b100 : node1518;
											assign node1518 = (inp[8]) ? 3'b000 : node1519;
												assign node1519 = (inp[6]) ? 3'b100 : 3'b000;
									assign node1524 = (inp[6]) ? node1532 : node1525;
										assign node1525 = (inp[11]) ? node1527 : 3'b100;
											assign node1527 = (inp[8]) ? node1529 : 3'b000;
												assign node1529 = (inp[2]) ? 3'b100 : 3'b000;
										assign node1532 = (inp[8]) ? 3'b000 : node1533;
											assign node1533 = (inp[2]) ? 3'b000 : 3'b100;
								assign node1537 = (inp[8]) ? node1557 : node1538;
									assign node1538 = (inp[5]) ? node1550 : node1539;
										assign node1539 = (inp[11]) ? node1545 : node1540;
											assign node1540 = (inp[2]) ? node1542 : 3'b000;
												assign node1542 = (inp[6]) ? 3'b000 : 3'b100;
											assign node1545 = (inp[6]) ? node1547 : 3'b000;
												assign node1547 = (inp[2]) ? 3'b000 : 3'b100;
										assign node1550 = (inp[6]) ? node1552 : 3'b000;
											assign node1552 = (inp[11]) ? node1554 : 3'b100;
												assign node1554 = (inp[2]) ? 3'b100 : 3'b000;
									assign node1557 = (inp[2]) ? node1569 : node1558;
										assign node1558 = (inp[11]) ? node1564 : node1559;
											assign node1559 = (inp[6]) ? 3'b100 : node1560;
												assign node1560 = (inp[5]) ? 3'b000 : 3'b100;
											assign node1564 = (inp[6]) ? node1566 : 3'b000;
												assign node1566 = (inp[5]) ? 3'b100 : 3'b000;
										assign node1569 = (inp[5]) ? node1571 : 3'b100;
											assign node1571 = (inp[6]) ? 3'b100 : 3'b000;
							assign node1574 = (inp[11]) ? node1600 : node1575;
								assign node1575 = (inp[8]) ? node1583 : node1576;
									assign node1576 = (inp[6]) ? 3'b110 : node1577;
										assign node1577 = (inp[10]) ? 3'b100 : node1578;
											assign node1578 = (inp[5]) ? 3'b110 : 3'b100;
									assign node1583 = (inp[6]) ? node1591 : node1584;
										assign node1584 = (inp[10]) ? node1588 : node1585;
											assign node1585 = (inp[5]) ? 3'b010 : 3'b000;
											assign node1588 = (inp[5]) ? 3'b000 : 3'b010;
										assign node1591 = (inp[2]) ? node1595 : node1592;
											assign node1592 = (inp[5]) ? 3'b010 : 3'b011;
											assign node1595 = (inp[10]) ? 3'b001 : node1596;
												assign node1596 = (inp[5]) ? 3'b001 : 3'b010;
								assign node1600 = (inp[10]) ? 3'b100 : node1601;
									assign node1601 = (inp[5]) ? node1609 : node1602;
										assign node1602 = (inp[6]) ? node1604 : 3'b110;
											assign node1604 = (inp[8]) ? 3'b101 : node1605;
												assign node1605 = (inp[2]) ? 3'b101 : 3'b110;
										assign node1609 = (inp[6]) ? 3'b110 : 3'b100;
						assign node1613 = (inp[6]) ? node1657 : node1614;
							assign node1614 = (inp[11]) ? node1632 : node1615;
								assign node1615 = (inp[7]) ? node1627 : node1616;
									assign node1616 = (inp[8]) ? node1622 : node1617;
										assign node1617 = (inp[5]) ? node1619 : 3'b100;
											assign node1619 = (inp[10]) ? 3'b000 : 3'b100;
										assign node1622 = (inp[5]) ? node1624 : 3'b010;
											assign node1624 = (inp[10]) ? 3'b000 : 3'b010;
									assign node1627 = (inp[5]) ? 3'b110 : node1628;
										assign node1628 = (inp[2]) ? 3'b010 : 3'b110;
								assign node1632 = (inp[5]) ? node1644 : node1633;
									assign node1633 = (inp[10]) ? node1639 : node1634;
										assign node1634 = (inp[7]) ? node1636 : 3'b010;
											assign node1636 = (inp[2]) ? 3'b000 : 3'b100;
										assign node1639 = (inp[7]) ? node1641 : 3'b100;
											assign node1641 = (inp[8]) ? 3'b000 : 3'b100;
									assign node1644 = (inp[10]) ? node1652 : node1645;
										assign node1645 = (inp[7]) ? node1647 : 3'b100;
											assign node1647 = (inp[2]) ? node1649 : 3'b000;
												assign node1649 = (inp[8]) ? 3'b100 : 3'b000;
										assign node1652 = (inp[8]) ? node1654 : 3'b000;
											assign node1654 = (inp[7]) ? 3'b100 : 3'b000;
							assign node1657 = (inp[7]) ? node1693 : node1658;
								assign node1658 = (inp[5]) ? node1672 : node1659;
									assign node1659 = (inp[8]) ? node1663 : node1660;
										assign node1660 = (inp[10]) ? 3'b110 : 3'b010;
										assign node1663 = (inp[11]) ? 3'b000 : node1664;
											assign node1664 = (inp[2]) ? node1668 : node1665;
												assign node1665 = (inp[10]) ? 3'b110 : 3'b000;
												assign node1668 = (inp[10]) ? 3'b000 : 3'b110;
									assign node1672 = (inp[10]) ? node1682 : node1673;
										assign node1673 = (inp[2]) ? node1677 : node1674;
											assign node1674 = (inp[8]) ? 3'b110 : 3'b010;
											assign node1677 = (inp[8]) ? node1679 : 3'b110;
												assign node1679 = (inp[11]) ? 3'b110 : 3'b000;
										assign node1682 = (inp[8]) ? node1688 : node1683;
											assign node1683 = (inp[2]) ? 3'b010 : node1684;
												assign node1684 = (inp[11]) ? 3'b100 : 3'b010;
											assign node1688 = (inp[11]) ? 3'b010 : node1689;
												assign node1689 = (inp[2]) ? 3'b110 : 3'b010;
								assign node1693 = (inp[2]) ? node1703 : node1694;
									assign node1694 = (inp[10]) ? node1698 : node1695;
										assign node1695 = (inp[8]) ? 3'b011 : 3'b100;
										assign node1698 = (inp[5]) ? node1700 : 3'b110;
											assign node1700 = (inp[11]) ? 3'b010 : 3'b110;
									assign node1703 = (inp[11]) ? node1711 : node1704;
										assign node1704 = (inp[5]) ? 3'b111 : node1705;
											assign node1705 = (inp[10]) ? 3'b011 : node1706;
												assign node1706 = (inp[8]) ? 3'b011 : 3'b001;
										assign node1711 = (inp[8]) ? 3'b101 : 3'b001;
					assign node1714 = (inp[6]) ? node1824 : node1715;
						assign node1715 = (inp[7]) ? node1759 : node1716;
							assign node1716 = (inp[1]) ? node1744 : node1717;
								assign node1717 = (inp[10]) ? node1731 : node1718;
									assign node1718 = (inp[2]) ? node1724 : node1719;
										assign node1719 = (inp[8]) ? node1721 : 3'b010;
											assign node1721 = (inp[5]) ? 3'b010 : 3'b110;
										assign node1724 = (inp[11]) ? 3'b010 : node1725;
											assign node1725 = (inp[8]) ? node1727 : 3'b110;
												assign node1727 = (inp[5]) ? 3'b100 : 3'b000;
									assign node1731 = (inp[5]) ? node1737 : node1732;
										assign node1732 = (inp[8]) ? 3'b010 : node1733;
											assign node1733 = (inp[2]) ? 3'b010 : 3'b100;
										assign node1737 = (inp[2]) ? node1739 : 3'b100;
											assign node1739 = (inp[11]) ? 3'b100 : node1740;
												assign node1740 = (inp[8]) ? 3'b010 : 3'b100;
								assign node1744 = (inp[10]) ? node1746 : 3'b110;
									assign node1746 = (inp[11]) ? node1752 : node1747;
										assign node1747 = (inp[8]) ? node1749 : 3'b010;
											assign node1749 = (inp[5]) ? 3'b010 : 3'b110;
										assign node1752 = (inp[8]) ? node1754 : 3'b100;
											assign node1754 = (inp[2]) ? 3'b010 : node1755;
												assign node1755 = (inp[5]) ? 3'b100 : 3'b010;
							assign node1759 = (inp[1]) ? node1791 : node1760;
								assign node1760 = (inp[8]) ? node1774 : node1761;
									assign node1761 = (inp[2]) ? node1767 : node1762;
										assign node1762 = (inp[10]) ? node1764 : 3'b010;
											assign node1764 = (inp[5]) ? 3'b000 : 3'b010;
										assign node1767 = (inp[10]) ? node1769 : 3'b100;
											assign node1769 = (inp[5]) ? node1771 : 3'b110;
												assign node1771 = (inp[11]) ? 3'b100 : 3'b110;
									assign node1774 = (inp[2]) ? node1780 : node1775;
										assign node1775 = (inp[10]) ? 3'b110 : node1776;
											assign node1776 = (inp[5]) ? 3'b110 : 3'b100;
										assign node1780 = (inp[11]) ? node1786 : node1781;
											assign node1781 = (inp[5]) ? node1783 : 3'b010;
												assign node1783 = (inp[10]) ? 3'b010 : 3'b000;
											assign node1786 = (inp[5]) ? 3'b110 : node1787;
												assign node1787 = (inp[10]) ? 3'b110 : 3'b100;
								assign node1791 = (inp[10]) ? node1807 : node1792;
									assign node1792 = (inp[2]) ? node1796 : node1793;
										assign node1793 = (inp[5]) ? 3'b001 : 3'b101;
										assign node1796 = (inp[11]) ? node1800 : node1797;
											assign node1797 = (inp[5]) ? 3'b001 : 3'b011;
											assign node1800 = (inp[8]) ? node1804 : node1801;
												assign node1801 = (inp[5]) ? 3'b110 : 3'b101;
												assign node1804 = (inp[5]) ? 3'b001 : 3'b011;
									assign node1807 = (inp[5]) ? node1817 : node1808;
										assign node1808 = (inp[8]) ? node1814 : node1809;
											assign node1809 = (inp[11]) ? 3'b110 : node1810;
												assign node1810 = (inp[2]) ? 3'b101 : 3'b100;
											assign node1814 = (inp[2]) ? 3'b001 : 3'b000;
										assign node1817 = (inp[11]) ? node1819 : 3'b110;
											assign node1819 = (inp[8]) ? node1821 : 3'b010;
												assign node1821 = (inp[2]) ? 3'b110 : 3'b010;
						assign node1824 = (inp[7]) ? node1880 : node1825;
							assign node1825 = (inp[1]) ? node1853 : node1826;
								assign node1826 = (inp[10]) ? node1840 : node1827;
									assign node1827 = (inp[2]) ? node1833 : node1828;
										assign node1828 = (inp[5]) ? 3'b110 : node1829;
											assign node1829 = (inp[8]) ? 3'b111 : 3'b011;
										assign node1833 = (inp[8]) ? node1837 : node1834;
											assign node1834 = (inp[5]) ? 3'b110 : 3'b011;
											assign node1837 = (inp[5]) ? 3'b001 : 3'b100;
									assign node1840 = (inp[5]) ? node1846 : node1841;
										assign node1841 = (inp[11]) ? 3'b110 : node1842;
											assign node1842 = (inp[2]) ? 3'b001 : 3'b000;
										assign node1846 = (inp[2]) ? node1848 : 3'b010;
											assign node1848 = (inp[8]) ? 3'b110 : node1849;
												assign node1849 = (inp[11]) ? 3'b010 : 3'b110;
								assign node1853 = (inp[10]) ? node1867 : node1854;
									assign node1854 = (inp[8]) ? node1862 : node1855;
										assign node1855 = (inp[5]) ? 3'b001 : node1856;
											assign node1856 = (inp[11]) ? 3'b101 : node1857;
												assign node1857 = (inp[2]) ? 3'b111 : 3'b101;
										assign node1862 = (inp[5]) ? 3'b101 : node1863;
											assign node1863 = (inp[2]) ? 3'b011 : 3'b001;
									assign node1867 = (inp[5]) ? node1875 : node1868;
										assign node1868 = (inp[8]) ? node1872 : node1869;
											assign node1869 = (inp[11]) ? 3'b001 : 3'b000;
											assign node1872 = (inp[11]) ? 3'b101 : 3'b100;
										assign node1875 = (inp[11]) ? 3'b110 : node1876;
											assign node1876 = (inp[2]) ? 3'b001 : 3'b110;
							assign node1880 = (inp[1]) ? node1904 : node1881;
								assign node1881 = (inp[10]) ? node1895 : node1882;
									assign node1882 = (inp[5]) ? node1888 : node1883;
										assign node1883 = (inp[8]) ? node1885 : 3'b101;
											assign node1885 = (inp[2]) ? 3'b010 : 3'b101;
										assign node1888 = (inp[2]) ? node1890 : 3'b001;
											assign node1890 = (inp[8]) ? 3'b101 : node1891;
												assign node1891 = (inp[11]) ? 3'b001 : 3'b101;
									assign node1895 = (inp[5]) ? node1899 : node1896;
										assign node1896 = (inp[11]) ? 3'b001 : 3'b101;
										assign node1899 = (inp[11]) ? 3'b110 : node1900;
											assign node1900 = (inp[2]) ? 3'b001 : 3'b110;
								assign node1904 = (inp[10]) ? node1916 : node1905;
									assign node1905 = (inp[2]) ? node1911 : node1906;
										assign node1906 = (inp[5]) ? 3'b011 : node1907;
											assign node1907 = (inp[11]) ? 3'b011 : 3'b111;
										assign node1911 = (inp[5]) ? node1913 : 3'b011;
											assign node1913 = (inp[11]) ? 3'b101 : 3'b011;
									assign node1916 = (inp[11]) ? node1922 : node1917;
										assign node1917 = (inp[5]) ? node1919 : 3'b011;
											assign node1919 = (inp[8]) ? 3'b101 : 3'b001;
										assign node1922 = (inp[5]) ? node1924 : 3'b101;
											assign node1924 = (inp[2]) ? 3'b001 : 3'b101;
				assign node1927 = (inp[0]) ? node2061 : node1928;
					assign node1928 = (inp[6]) ? node1964 : node1929;
						assign node1929 = (inp[1]) ? node1931 : 3'b000;
							assign node1931 = (inp[10]) ? node1955 : node1932;
								assign node1932 = (inp[7]) ? node1942 : node1933;
									assign node1933 = (inp[8]) ? node1935 : 3'b000;
										assign node1935 = (inp[2]) ? node1937 : 3'b000;
											assign node1937 = (inp[5]) ? 3'b000 : node1938;
												assign node1938 = (inp[11]) ? 3'b000 : 3'b100;
									assign node1942 = (inp[5]) ? node1948 : node1943;
										assign node1943 = (inp[11]) ? 3'b100 : node1944;
											assign node1944 = (inp[8]) ? 3'b010 : 3'b100;
										assign node1948 = (inp[2]) ? node1952 : node1949;
											assign node1949 = (inp[8]) ? 3'b000 : 3'b100;
											assign node1952 = (inp[8]) ? 3'b100 : 3'b000;
								assign node1955 = (inp[11]) ? 3'b000 : node1956;
									assign node1956 = (inp[5]) ? 3'b000 : node1957;
										assign node1957 = (inp[2]) ? node1959 : 3'b000;
											assign node1959 = (inp[8]) ? 3'b010 : 3'b000;
						assign node1964 = (inp[10]) ? node2026 : node1965;
							assign node1965 = (inp[5]) ? node1999 : node1966;
								assign node1966 = (inp[8]) ? node1982 : node1967;
									assign node1967 = (inp[7]) ? node1973 : node1968;
										assign node1968 = (inp[1]) ? node1970 : 3'b100;
											assign node1970 = (inp[11]) ? 3'b010 : 3'b110;
										assign node1973 = (inp[2]) ? 3'b010 : node1974;
											assign node1974 = (inp[11]) ? node1978 : node1975;
												assign node1975 = (inp[1]) ? 3'b000 : 3'b010;
												assign node1978 = (inp[1]) ? 3'b010 : 3'b100;
									assign node1982 = (inp[1]) ? node1994 : node1983;
										assign node1983 = (inp[7]) ? node1989 : node1984;
											assign node1984 = (inp[2]) ? node1986 : 3'b100;
												assign node1986 = (inp[11]) ? 3'b100 : 3'b000;
											assign node1989 = (inp[11]) ? 3'b010 : node1990;
												assign node1990 = (inp[2]) ? 3'b100 : 3'b010;
										assign node1994 = (inp[7]) ? 3'b100 : node1995;
											assign node1995 = (inp[11]) ? 3'b010 : 3'b110;
								assign node1999 = (inp[7]) ? node2013 : node2000;
									assign node2000 = (inp[11]) ? node2006 : node2001;
										assign node2001 = (inp[2]) ? 3'b100 : node2002;
											assign node2002 = (inp[8]) ? 3'b100 : 3'b000;
										assign node2006 = (inp[1]) ? node2008 : 3'b000;
											assign node2008 = (inp[2]) ? node2010 : 3'b000;
												assign node2010 = (inp[8]) ? 3'b100 : 3'b000;
									assign node2013 = (inp[11]) ? node2019 : node2014;
										assign node2014 = (inp[2]) ? 3'b010 : node2015;
											assign node2015 = (inp[1]) ? 3'b010 : 3'b100;
										assign node2019 = (inp[1]) ? 3'b100 : node2020;
											assign node2020 = (inp[2]) ? 3'b100 : node2021;
												assign node2021 = (inp[8]) ? 3'b100 : 3'b000;
							assign node2026 = (inp[5]) ? node2050 : node2027;
								assign node2027 = (inp[11]) ? node2041 : node2028;
									assign node2028 = (inp[2]) ? node2034 : node2029;
										assign node2029 = (inp[1]) ? 3'b100 : node2030;
											assign node2030 = (inp[8]) ? 3'b100 : 3'b000;
										assign node2034 = (inp[1]) ? node2038 : node2035;
											assign node2035 = (inp[7]) ? 3'b100 : 3'b000;
											assign node2038 = (inp[7]) ? 3'b010 : 3'b100;
									assign node2041 = (inp[8]) ? node2043 : 3'b000;
										assign node2043 = (inp[7]) ? 3'b100 : node2044;
											assign node2044 = (inp[2]) ? node2046 : 3'b000;
												assign node2046 = (inp[1]) ? 3'b100 : 3'b000;
								assign node2050 = (inp[1]) ? node2052 : 3'b000;
									assign node2052 = (inp[7]) ? node2054 : 3'b000;
										assign node2054 = (inp[8]) ? 3'b100 : node2055;
											assign node2055 = (inp[2]) ? node2057 : 3'b000;
												assign node2057 = (inp[11]) ? 3'b000 : 3'b100;
					assign node2061 = (inp[6]) ? node2141 : node2062;
						assign node2062 = (inp[10]) ? node2112 : node2063;
							assign node2063 = (inp[5]) ? node2095 : node2064;
								assign node2064 = (inp[7]) ? node2080 : node2065;
									assign node2065 = (inp[8]) ? node2073 : node2066;
										assign node2066 = (inp[1]) ? 3'b100 : node2067;
											assign node2067 = (inp[2]) ? 3'b100 : node2068;
												assign node2068 = (inp[11]) ? 3'b000 : 3'b100;
										assign node2073 = (inp[2]) ? 3'b010 : node2074;
											assign node2074 = (inp[1]) ? node2076 : 3'b100;
												assign node2076 = (inp[11]) ? 3'b100 : 3'b010;
									assign node2080 = (inp[1]) ? node2092 : node2081;
										assign node2081 = (inp[8]) ? node2087 : node2082;
											assign node2082 = (inp[2]) ? node2084 : 3'b100;
												assign node2084 = (inp[11]) ? 3'b100 : 3'b010;
											assign node2087 = (inp[2]) ? 3'b010 : node2088;
												assign node2088 = (inp[11]) ? 3'b100 : 3'b010;
										assign node2092 = (inp[8]) ? 3'b110 : 3'b010;
								assign node2095 = (inp[11]) ? node2107 : node2096;
									assign node2096 = (inp[8]) ? 3'b100 : node2097;
										assign node2097 = (inp[2]) ? node2101 : node2098;
											assign node2098 = (inp[7]) ? 3'b100 : 3'b000;
											assign node2101 = (inp[1]) ? node2103 : 3'b100;
												assign node2103 = (inp[7]) ? 3'b010 : 3'b100;
									assign node2107 = (inp[1]) ? node2109 : 3'b000;
										assign node2109 = (inp[8]) ? 3'b100 : 3'b000;
							assign node2112 = (inp[5]) ? 3'b000 : node2113;
								assign node2113 = (inp[7]) ? node2123 : node2114;
									assign node2114 = (inp[11]) ? 3'b000 : node2115;
										assign node2115 = (inp[1]) ? node2117 : 3'b000;
											assign node2117 = (inp[8]) ? 3'b100 : node2118;
												assign node2118 = (inp[2]) ? 3'b100 : 3'b000;
									assign node2123 = (inp[1]) ? node2135 : node2124;
										assign node2124 = (inp[11]) ? node2130 : node2125;
											assign node2125 = (inp[8]) ? 3'b100 : node2126;
												assign node2126 = (inp[2]) ? 3'b100 : 3'b000;
											assign node2130 = (inp[8]) ? node2132 : 3'b000;
												assign node2132 = (inp[2]) ? 3'b100 : 3'b000;
										assign node2135 = (inp[11]) ? 3'b100 : node2136;
											assign node2136 = (inp[8]) ? 3'b010 : 3'b100;
						assign node2141 = (inp[10]) ? node2197 : node2142;
							assign node2142 = (inp[5]) ? node2174 : node2143;
								assign node2143 = (inp[1]) ? node2161 : node2144;
									assign node2144 = (inp[7]) ? node2158 : node2145;
										assign node2145 = (inp[11]) ? node2151 : node2146;
											assign node2146 = (inp[8]) ? 3'b110 : node2147;
												assign node2147 = (inp[2]) ? 3'b110 : 3'b010;
											assign node2151 = (inp[8]) ? node2155 : node2152;
												assign node2152 = (inp[2]) ? 3'b010 : 3'b000;
												assign node2155 = (inp[2]) ? 3'b110 : 3'b010;
										assign node2158 = (inp[2]) ? 3'b001 : 3'b110;
									assign node2161 = (inp[11]) ? node2167 : node2162;
										assign node2162 = (inp[8]) ? node2164 : 3'b001;
											assign node2164 = (inp[7]) ? 3'b111 : 3'b001;
										assign node2167 = (inp[7]) ? node2169 : 3'b110;
											assign node2169 = (inp[8]) ? 3'b001 : node2170;
												assign node2170 = (inp[2]) ? 3'b001 : 3'b110;
								assign node2174 = (inp[7]) ? node2184 : node2175;
									assign node2175 = (inp[8]) ? node2177 : 3'b010;
										assign node2177 = (inp[1]) ? node2181 : node2178;
											assign node2178 = (inp[11]) ? 3'b110 : 3'b010;
											assign node2181 = (inp[11]) ? 3'b010 : 3'b110;
									assign node2184 = (inp[1]) ? 3'b110 : node2185;
										assign node2185 = (inp[8]) ? node2191 : node2186;
											assign node2186 = (inp[11]) ? 3'b010 : node2187;
												assign node2187 = (inp[2]) ? 3'b110 : 3'b010;
											assign node2191 = (inp[2]) ? 3'b110 : node2192;
												assign node2192 = (inp[11]) ? 3'b010 : 3'b110;
							assign node2197 = (inp[5]) ? node2215 : node2198;
								assign node2198 = (inp[11]) ? node2204 : node2199;
									assign node2199 = (inp[7]) ? 3'b110 : node2200;
										assign node2200 = (inp[8]) ? 3'b110 : 3'b010;
									assign node2204 = (inp[2]) ? node2210 : node2205;
										assign node2205 = (inp[7]) ? node2207 : 3'b100;
											assign node2207 = (inp[8]) ? 3'b110 : 3'b010;
										assign node2210 = (inp[1]) ? node2212 : 3'b010;
											assign node2212 = (inp[7]) ? 3'b110 : 3'b010;
								assign node2215 = (inp[7]) ? node2225 : node2216;
									assign node2216 = (inp[8]) ? 3'b100 : node2217;
										assign node2217 = (inp[11]) ? 3'b000 : node2218;
											assign node2218 = (inp[2]) ? 3'b100 : node2219;
												assign node2219 = (inp[1]) ? 3'b100 : 3'b000;
									assign node2225 = (inp[11]) ? node2227 : 3'b010;
										assign node2227 = (inp[2]) ? node2229 : 3'b100;
											assign node2229 = (inp[1]) ? 3'b010 : 3'b100;
			assign node2232 = (inp[9]) ? node2508 : node2233;
				assign node2233 = (inp[6]) ? node2327 : node2234;
					assign node2234 = (inp[0]) ? node2258 : node2235;
						assign node2235 = (inp[1]) ? node2237 : 3'b000;
							assign node2237 = (inp[7]) ? node2239 : 3'b000;
								assign node2239 = (inp[5]) ? node2251 : node2240;
									assign node2240 = (inp[8]) ? node2246 : node2241;
										assign node2241 = (inp[2]) ? node2243 : 3'b000;
											assign node2243 = (inp[10]) ? 3'b000 : 3'b100;
										assign node2246 = (inp[2]) ? node2248 : 3'b100;
											assign node2248 = (inp[10]) ? 3'b100 : 3'b000;
									assign node2251 = (inp[8]) ? node2253 : 3'b000;
										assign node2253 = (inp[11]) ? 3'b000 : node2254;
											assign node2254 = (inp[2]) ? 3'b100 : 3'b000;
						assign node2258 = (inp[7]) ? node2284 : node2259;
							assign node2259 = (inp[1]) ? node2261 : 3'b000;
								assign node2261 = (inp[11]) ? node2273 : node2262;
									assign node2262 = (inp[2]) ? node2268 : node2263;
										assign node2263 = (inp[5]) ? 3'b100 : node2264;
											assign node2264 = (inp[8]) ? 3'b001 : 3'b100;
										assign node2268 = (inp[10]) ? node2270 : 3'b100;
											assign node2270 = (inp[5]) ? 3'b000 : 3'b100;
									assign node2273 = (inp[5]) ? 3'b000 : node2274;
										assign node2274 = (inp[2]) ? node2278 : node2275;
											assign node2275 = (inp[10]) ? 3'b000 : 3'b100;
											assign node2278 = (inp[10]) ? node2280 : 3'b000;
												assign node2280 = (inp[8]) ? 3'b100 : 3'b000;
							assign node2284 = (inp[1]) ? node2302 : node2285;
								assign node2285 = (inp[5]) ? node2295 : node2286;
									assign node2286 = (inp[10]) ? node2290 : node2287;
										assign node2287 = (inp[8]) ? 3'b001 : 3'b100;
										assign node2290 = (inp[8]) ? 3'b100 : node2291;
											assign node2291 = (inp[11]) ? 3'b000 : 3'b100;
									assign node2295 = (inp[10]) ? 3'b000 : node2296;
										assign node2296 = (inp[8]) ? 3'b100 : node2297;
											assign node2297 = (inp[11]) ? 3'b000 : 3'b100;
								assign node2302 = (inp[10]) ? node2316 : node2303;
									assign node2303 = (inp[8]) ? node2307 : node2304;
										assign node2304 = (inp[5]) ? 3'b100 : 3'b110;
										assign node2307 = (inp[11]) ? node2311 : node2308;
											assign node2308 = (inp[5]) ? 3'b010 : 3'b000;
											assign node2311 = (inp[2]) ? 3'b010 : node2312;
												assign node2312 = (inp[5]) ? 3'b100 : 3'b110;
									assign node2316 = (inp[8]) ? node2324 : node2317;
										assign node2317 = (inp[2]) ? node2319 : 3'b000;
											assign node2319 = (inp[5]) ? node2321 : 3'b100;
												assign node2321 = (inp[11]) ? 3'b000 : 3'b100;
										assign node2324 = (inp[2]) ? 3'b010 : 3'b100;
					assign node2327 = (inp[0]) ? node2407 : node2328;
						assign node2328 = (inp[7]) ? node2358 : node2329;
							assign node2329 = (inp[10]) ? node2349 : node2330;
								assign node2330 = (inp[2]) ? node2336 : node2331;
									assign node2331 = (inp[11]) ? 3'b000 : node2332;
										assign node2332 = (inp[8]) ? 3'b100 : 3'b000;
									assign node2336 = (inp[1]) ? 3'b100 : node2337;
										assign node2337 = (inp[5]) ? node2343 : node2338;
											assign node2338 = (inp[8]) ? node2340 : 3'b100;
												assign node2340 = (inp[11]) ? 3'b100 : 3'b000;
											assign node2343 = (inp[8]) ? node2345 : 3'b000;
												assign node2345 = (inp[11]) ? 3'b000 : 3'b100;
								assign node2349 = (inp[8]) ? node2351 : 3'b000;
									assign node2351 = (inp[11]) ? 3'b000 : node2352;
										assign node2352 = (inp[1]) ? 3'b000 : node2353;
											assign node2353 = (inp[5]) ? 3'b000 : 3'b100;
							assign node2358 = (inp[10]) ? node2388 : node2359;
								assign node2359 = (inp[11]) ? node2375 : node2360;
									assign node2360 = (inp[8]) ? node2366 : node2361;
										assign node2361 = (inp[2]) ? node2363 : 3'b100;
											assign node2363 = (inp[5]) ? 3'b010 : 3'b110;
										assign node2366 = (inp[1]) ? 3'b010 : node2367;
											assign node2367 = (inp[5]) ? node2371 : node2368;
												assign node2368 = (inp[2]) ? 3'b000 : 3'b010;
												assign node2371 = (inp[2]) ? 3'b010 : 3'b000;
									assign node2375 = (inp[5]) ? node2381 : node2376;
										assign node2376 = (inp[8]) ? 3'b110 : node2377;
											assign node2377 = (inp[1]) ? 3'b010 : 3'b100;
										assign node2381 = (inp[8]) ? node2383 : 3'b100;
											assign node2383 = (inp[2]) ? node2385 : 3'b100;
												assign node2385 = (inp[1]) ? 3'b010 : 3'b100;
								assign node2388 = (inp[11]) ? node2398 : node2389;
									assign node2389 = (inp[5]) ? node2395 : node2390;
										assign node2390 = (inp[8]) ? 3'b010 : node2391;
											assign node2391 = (inp[1]) ? 3'b010 : 3'b000;
										assign node2395 = (inp[1]) ? 3'b100 : 3'b000;
									assign node2398 = (inp[8]) ? node2400 : 3'b000;
										assign node2400 = (inp[2]) ? node2402 : 3'b000;
											assign node2402 = (inp[5]) ? node2404 : 3'b000;
												assign node2404 = (inp[1]) ? 3'b100 : 3'b000;
						assign node2407 = (inp[1]) ? node2463 : node2408;
							assign node2408 = (inp[10]) ? node2434 : node2409;
								assign node2409 = (inp[2]) ? node2417 : node2410;
									assign node2410 = (inp[5]) ? node2412 : 3'b110;
										assign node2412 = (inp[7]) ? node2414 : 3'b100;
											assign node2414 = (inp[8]) ? 3'b110 : 3'b010;
									assign node2417 = (inp[11]) ? node2425 : node2418;
										assign node2418 = (inp[5]) ? node2422 : node2419;
											assign node2419 = (inp[7]) ? 3'b001 : 3'b000;
											assign node2422 = (inp[7]) ? 3'b110 : 3'b010;
										assign node2425 = (inp[5]) ? node2427 : 3'b110;
											assign node2427 = (inp[7]) ? node2431 : node2428;
												assign node2428 = (inp[8]) ? 3'b010 : 3'b100;
												assign node2431 = (inp[8]) ? 3'b110 : 3'b010;
								assign node2434 = (inp[5]) ? node2450 : node2435;
									assign node2435 = (inp[8]) ? node2445 : node2436;
										assign node2436 = (inp[7]) ? node2442 : node2437;
											assign node2437 = (inp[11]) ? 3'b100 : node2438;
												assign node2438 = (inp[2]) ? 3'b110 : 3'b100;
											assign node2442 = (inp[11]) ? 3'b010 : 3'b110;
										assign node2445 = (inp[7]) ? node2447 : 3'b010;
											assign node2447 = (inp[11]) ? 3'b010 : 3'b110;
									assign node2450 = (inp[7]) ? node2458 : node2451;
										assign node2451 = (inp[11]) ? node2453 : 3'b100;
											assign node2453 = (inp[8]) ? node2455 : 3'b000;
												assign node2455 = (inp[2]) ? 3'b100 : 3'b000;
										assign node2458 = (inp[11]) ? 3'b100 : node2459;
											assign node2459 = (inp[8]) ? 3'b010 : 3'b100;
							assign node2463 = (inp[10]) ? node2489 : node2464;
								assign node2464 = (inp[5]) ? node2478 : node2465;
									assign node2465 = (inp[11]) ? node2471 : node2466;
										assign node2466 = (inp[8]) ? node2468 : 3'b001;
											assign node2468 = (inp[7]) ? 3'b101 : 3'b001;
										assign node2471 = (inp[7]) ? node2473 : 3'b010;
											assign node2473 = (inp[8]) ? 3'b001 : node2474;
												assign node2474 = (inp[2]) ? 3'b001 : 3'b000;
									assign node2478 = (inp[11]) ? node2484 : node2479;
										assign node2479 = (inp[8]) ? node2481 : 3'b110;
											assign node2481 = (inp[2]) ? 3'b001 : 3'b110;
										assign node2484 = (inp[7]) ? node2486 : 3'b010;
											assign node2486 = (inp[2]) ? 3'b110 : 3'b010;
								assign node2489 = (inp[11]) ? node2495 : node2490;
									assign node2490 = (inp[5]) ? node2492 : 3'b110;
										assign node2492 = (inp[7]) ? 3'b110 : 3'b010;
									assign node2495 = (inp[5]) ? node2501 : node2496;
										assign node2496 = (inp[2]) ? node2498 : 3'b010;
											assign node2498 = (inp[7]) ? 3'b110 : 3'b010;
										assign node2501 = (inp[8]) ? 3'b010 : node2502;
											assign node2502 = (inp[7]) ? node2504 : 3'b100;
												assign node2504 = (inp[2]) ? 3'b010 : 3'b100;
				assign node2508 = (inp[6]) ? node2524 : node2509;
					assign node2509 = (inp[10]) ? 3'b000 : node2510;
						assign node2510 = (inp[5]) ? 3'b000 : node2511;
							assign node2511 = (inp[11]) ? 3'b000 : node2512;
								assign node2512 = (inp[0]) ? node2514 : 3'b000;
									assign node2514 = (inp[1]) ? node2518 : node2515;
										assign node2515 = (inp[7]) ? 3'b010 : 3'b000;
										assign node2518 = (inp[7]) ? 3'b100 : 3'b000;
					assign node2524 = (inp[1]) ? node2548 : node2525;
						assign node2525 = (inp[0]) ? node2527 : 3'b000;
							assign node2527 = (inp[7]) ? node2529 : 3'b000;
								assign node2529 = (inp[10]) ? node2539 : node2530;
									assign node2530 = (inp[11]) ? node2536 : node2531;
										assign node2531 = (inp[5]) ? node2533 : 3'b010;
											assign node2533 = (inp[8]) ? 3'b100 : 3'b000;
										assign node2536 = (inp[5]) ? 3'b000 : 3'b100;
									assign node2539 = (inp[2]) ? node2541 : 3'b000;
										assign node2541 = (inp[11]) ? 3'b000 : node2542;
											assign node2542 = (inp[5]) ? 3'b000 : node2543;
												assign node2543 = (inp[8]) ? 3'b100 : 3'b000;
						assign node2548 = (inp[5]) ? node2584 : node2549;
							assign node2549 = (inp[10]) ? node2567 : node2550;
								assign node2550 = (inp[7]) ? node2564 : node2551;
									assign node2551 = (inp[0]) ? node2553 : 3'b000;
										assign node2553 = (inp[11]) ? node2559 : node2554;
											assign node2554 = (inp[2]) ? node2556 : 3'b100;
												assign node2556 = (inp[8]) ? 3'b010 : 3'b100;
											assign node2559 = (inp[8]) ? 3'b100 : node2560;
												assign node2560 = (inp[2]) ? 3'b100 : 3'b000;
									assign node2564 = (inp[0]) ? 3'b010 : 3'b100;
								assign node2567 = (inp[0]) ? node2569 : 3'b000;
									assign node2569 = (inp[8]) ? node2575 : node2570;
										assign node2570 = (inp[2]) ? node2572 : 3'b000;
											assign node2572 = (inp[7]) ? 3'b100 : 3'b000;
										assign node2575 = (inp[2]) ? node2577 : 3'b100;
											assign node2577 = (inp[11]) ? node2581 : node2578;
												assign node2578 = (inp[7]) ? 3'b010 : 3'b100;
												assign node2581 = (inp[7]) ? 3'b100 : 3'b000;
							assign node2584 = (inp[0]) ? node2586 : 3'b000;
								assign node2586 = (inp[8]) ? node2594 : node2587;
									assign node2587 = (inp[7]) ? node2589 : 3'b000;
										assign node2589 = (inp[10]) ? 3'b000 : node2590;
											assign node2590 = (inp[11]) ? 3'b000 : 3'b100;
									assign node2594 = (inp[11]) ? node2600 : node2595;
										assign node2595 = (inp[10]) ? node2597 : 3'b100;
											assign node2597 = (inp[2]) ? 3'b100 : 3'b000;
										assign node2600 = (inp[10]) ? 3'b000 : node2601;
											assign node2601 = (inp[7]) ? 3'b100 : 3'b000;

endmodule