module dtc_split5_bm37 (
	input  wire [8-1:0] inp,
	output wire [63-1:0] outp
);

	wire [63-1:0] node1;
	wire [63-1:0] node2;
	wire [63-1:0] node3;
	wire [63-1:0] node4;
	wire [63-1:0] node5;
	wire [63-1:0] node8;
	wire [63-1:0] node11;
	wire [63-1:0] node12;
	wire [63-1:0] node15;
	wire [63-1:0] node18;
	wire [63-1:0] node19;
	wire [63-1:0] node21;
	wire [63-1:0] node24;
	wire [63-1:0] node25;
	wire [63-1:0] node28;
	wire [63-1:0] node31;
	wire [63-1:0] node32;
	wire [63-1:0] node33;
	wire [63-1:0] node36;
	wire [63-1:0] node38;
	wire [63-1:0] node41;
	wire [63-1:0] node42;
	wire [63-1:0] node43;
	wire [63-1:0] node46;
	wire [63-1:0] node49;
	wire [63-1:0] node50;
	wire [63-1:0] node54;
	wire [63-1:0] node55;
	wire [63-1:0] node56;
	wire [63-1:0] node57;
	wire [63-1:0] node58;
	wire [63-1:0] node61;
	wire [63-1:0] node64;
	wire [63-1:0] node65;
	wire [63-1:0] node69;
	wire [63-1:0] node70;
	wire [63-1:0] node71;
	wire [63-1:0] node74;
	wire [63-1:0] node77;
	wire [63-1:0] node78;
	wire [63-1:0] node82;
	wire [63-1:0] node83;
	wire [63-1:0] node84;
	wire [63-1:0] node85;
	wire [63-1:0] node88;
	wire [63-1:0] node91;
	wire [63-1:0] node92;
	wire [63-1:0] node95;
	wire [63-1:0] node98;
	wire [63-1:0] node99;
	wire [63-1:0] node100;
	wire [63-1:0] node103;
	wire [63-1:0] node106;
	wire [63-1:0] node107;
	wire [63-1:0] node110;

	assign outp = (inp[7]) ? node54 : node1;
		assign node1 = (inp[6]) ? node31 : node2;
			assign node2 = (inp[1]) ? node18 : node3;
				assign node3 = (inp[2]) ? node11 : node4;
					assign node4 = (inp[3]) ? node8 : node5;
						assign node5 = (inp[0]) ? 63'b100111101001100000110001101110110010010101001101001101001010101 : 63'b100111101001100000110001101110110010010101001100001101001010101;
						assign node8 = (inp[4]) ? 63'b100110101001100000110001101110110011010101001100000101001010101 : 63'b100110101001100000110001101110110011010101001100000101001010101;
					assign node11 = (inp[4]) ? node15 : node12;
						assign node12 = (inp[0]) ? 63'b100111101001000000110001101110110011000110001100101001001010101 : 63'b100111101001100000110001101110110011010101001100101101001010101;
						assign node15 = (inp[0]) ? 63'b100110101001100000110001101110110011010101011101000101001010101 : 63'b100101101001110000110001101110110011010101001100101101001010101;
				assign node18 = (inp[2]) ? node24 : node19;
					assign node19 = (inp[3]) ? node21 : 63'b100111101001100000010001101110010010010101001100101101000000101;
						assign node21 = (inp[5]) ? 63'b100001101001100000010001101110010010010101001101101101000010101 : 63'b100001101001100000010001101110010010010101001100101101000010101;
					assign node24 = (inp[4]) ? node28 : node25;
						assign node25 = (inp[3]) ? 63'b100001101001100000110001101110110011010101001100101101001010101 : 63'b100111101001100100110001101110110011010101001100101101001010101;
						assign node28 = (inp[5]) ? 63'b100111101001100000110001101110110011010101001100101101001010101 : 63'b100001101001100000110001101110010010010101011100101101000000101;
			assign node31 = (inp[2]) ? node41 : node32;
				assign node32 = (inp[3]) ? node36 : node33;
					assign node33 = (inp[1]) ? 63'b100110101001100000110001101110110011010101000100001101001010001 : 63'b100110101001100000110001101110110001010101000100101101001010000;
					assign node36 = (inp[1]) ? node38 : 63'b100110101001100000110001101110110011010001001100001101001010101;
						assign node38 = (inp[0]) ? 63'b100110101001100000110001101110100011010101001100100101001010100 : 63'b100110101001100000110001101110100011010101001100100101001010100;
				assign node41 = (inp[5]) ? node49 : node42;
					assign node42 = (inp[4]) ? node46 : node43;
						assign node43 = (inp[0]) ? 63'b100111101001100000110001101110110011010101001100101101001010101 : 63'b100111101001100000110001101110110011010101001100101101011010100;
						assign node46 = (inp[1]) ? 63'b100111101001100000110001101110110011010101001100101101001010101 : 63'b100110101001100000110001101110110001010001010100001101001010000;
					assign node49 = (inp[0]) ? 63'b100111101001000000110001101110110011010100001100101101001110101 : node50;
						assign node50 = (inp[4]) ? 63'b100101101001100000110001101110110011010101001100101101001010101 : 63'b100111101001100100110001101110110011010101001100101101001010101;
		assign node54 = (inp[2]) ? node82 : node55;
			assign node55 = (inp[3]) ? node69 : node56;
				assign node56 = (inp[1]) ? node64 : node57;
					assign node57 = (inp[6]) ? node61 : node58;
						assign node58 = (inp[0]) ? 63'b100111101001100000110001101110110011010101001000101101001000101 : 63'b100111101001100000110001101110110011010101001000101101001000101;
						assign node61 = (inp[4]) ? 63'b100111101001000000110001101000110111010101001100101100001010101 : 63'b100111101000000000110001100000110011010101001100101100001010101;
					assign node64 = (inp[6]) ? 63'b100111101001100000110001001110110011010101001100101101000010101 : node65;
						assign node65 = (inp[0]) ? 63'b100111101001100000110001101110110011010101001100101101000010101 : 63'b100111101001100000110001101110110011010101001100101101000010101;
				assign node69 = (inp[6]) ? node77 : node70;
					assign node70 = (inp[4]) ? node74 : node71;
						assign node71 = (inp[1]) ? 63'b100111101000000000110001100000110011010101001100101100001010101 : 63'b100001101000000000110001100000110011010101001100101100001010101;
						assign node74 = (inp[0]) ? 63'b000111101001001000110001101010110011000101001101101101001010101 : 63'b000111101001001000110001101010110011000101001100101101001010101;
					assign node77 = (inp[1]) ? 63'b100111101000000000110000100100110011010101101100101101001010101 : node78;
						assign node78 = (inp[4]) ? 63'b100111101001100000100001101110110010010101001100101101000010101 : 63'b100111101011100000100001101110110010010101001100101101000010101;
			assign node82 = (inp[0]) ? node98 : node83;
				assign node83 = (inp[4]) ? node91 : node84;
					assign node84 = (inp[5]) ? node88 : node85;
						assign node85 = (inp[6]) ? 63'b100111101001100000010001101110110011010101001100000101001010101 : 63'b100111101001100000110001101110110011010101001100101101001010101;
						assign node88 = (inp[1]) ? 63'b100111101001100100110001101110110011010101001100101101001010101 : 63'b100001101001100100110001101110110011010101001100101101001010101;
					assign node91 = (inp[5]) ? node95 : node92;
						assign node92 = (inp[6]) ? 63'b100111001001100000110001101110110001010101000100101101001000001 : 63'b100111100001000000110001101110110011000100001100101001001010101;
						assign node95 = (inp[1]) ? 63'b100111101001100000110001101110110011010101001100101101001010101 : 63'b100101101001110000110001101110110011010101001100101101001010101;
				assign node98 = (inp[4]) ? node106 : node99;
					assign node99 = (inp[1]) ? node103 : node100;
						assign node100 = (inp[6]) ? 63'b100111101001000000110001101110110011000110001100101001001010101 : 63'b100001101001000000110001101110110011000110001100101001001010101;
						assign node103 = (inp[5]) ? 63'b100111101001000000110001101110110011010100001100101101001110101 : 63'b100111101001100000110001101110110011010101001100101101001010101;
					assign node106 = (inp[6]) ? node110 : node107;
						assign node107 = (inp[5]) ? 63'b100111101000000000110000101100110011010101011101101101001011101 : 63'b100111101000000000110000101100110011010101011100101101001011101;
						assign node110 = (inp[3]) ? 63'b100111101001100000100001101110110010010101011100101101000010101 : 63'b100111101001100000110001001110110010010101011101101101000010101;

endmodule