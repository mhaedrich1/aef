module dtc_split33_bm97 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node7;
	wire [3-1:0] node8;
	wire [3-1:0] node9;
	wire [3-1:0] node11;
	wire [3-1:0] node15;
	wire [3-1:0] node16;
	wire [3-1:0] node17;
	wire [3-1:0] node19;
	wire [3-1:0] node22;
	wire [3-1:0] node23;
	wire [3-1:0] node27;
	wire [3-1:0] node28;
	wire [3-1:0] node34;
	wire [3-1:0] node35;
	wire [3-1:0] node37;
	wire [3-1:0] node39;
	wire [3-1:0] node41;
	wire [3-1:0] node42;
	wire [3-1:0] node43;
	wire [3-1:0] node45;
	wire [3-1:0] node48;
	wire [3-1:0] node50;
	wire [3-1:0] node51;
	wire [3-1:0] node55;
	wire [3-1:0] node57;
	wire [3-1:0] node58;
	wire [3-1:0] node61;
	wire [3-1:0] node62;
	wire [3-1:0] node65;
	wire [3-1:0] node68;
	wire [3-1:0] node69;
	wire [3-1:0] node70;
	wire [3-1:0] node73;
	wire [3-1:0] node75;
	wire [3-1:0] node77;
	wire [3-1:0] node79;
	wire [3-1:0] node80;
	wire [3-1:0] node82;
	wire [3-1:0] node85;
	wire [3-1:0] node86;
	wire [3-1:0] node90;
	wire [3-1:0] node91;
	wire [3-1:0] node92;
	wire [3-1:0] node93;
	wire [3-1:0] node95;
	wire [3-1:0] node98;
	wire [3-1:0] node99;
	wire [3-1:0] node101;
	wire [3-1:0] node104;
	wire [3-1:0] node106;
	wire [3-1:0] node109;
	wire [3-1:0] node111;
	wire [3-1:0] node113;
	wire [3-1:0] node116;
	wire [3-1:0] node118;
	wire [3-1:0] node119;
	wire [3-1:0] node121;
	wire [3-1:0] node122;

	assign outp = (inp[9]) ? node34 : node1;
		assign node1 = (inp[3]) ? node3 : 3'b000;
			assign node3 = (inp[7]) ? 3'b000 : node4;
				assign node4 = (inp[6]) ? 3'b000 : node5;
					assign node5 = (inp[4]) ? node7 : 3'b100;
						assign node7 = (inp[11]) ? node15 : node8;
							assign node8 = (inp[8]) ? 3'b100 : node9;
								assign node9 = (inp[10]) ? node11 : 3'b100;
									assign node11 = (inp[1]) ? 3'b100 : 3'b000;
							assign node15 = (inp[5]) ? node27 : node16;
								assign node16 = (inp[10]) ? node22 : node17;
									assign node17 = (inp[0]) ? node19 : 3'b100;
										assign node19 = (inp[2]) ? 3'b000 : 3'b100;
									assign node22 = (inp[8]) ? 3'b000 : node23;
										assign node23 = (inp[1]) ? 3'b000 : 3'b100;
								assign node27 = (inp[10]) ? 3'b000 : node28;
									assign node28 = (inp[1]) ? 3'b000 : 3'b100;
		assign node34 = (inp[3]) ? node68 : node35;
			assign node35 = (inp[6]) ? node37 : 3'b000;
				assign node37 = (inp[7]) ? node39 : 3'b001;
					assign node39 = (inp[10]) ? node41 : 3'b000;
						assign node41 = (inp[4]) ? node55 : node42;
							assign node42 = (inp[8]) ? node48 : node43;
								assign node43 = (inp[5]) ? node45 : 3'b000;
									assign node45 = (inp[11]) ? 3'b001 : 3'b000;
								assign node48 = (inp[11]) ? node50 : 3'b000;
									assign node50 = (inp[2]) ? 3'b100 : node51;
										assign node51 = (inp[1]) ? 3'b100 : 3'b101;
							assign node55 = (inp[11]) ? node57 : 3'b100;
								assign node57 = (inp[5]) ? node61 : node58;
									assign node58 = (inp[8]) ? 3'b100 : 3'b000;
									assign node61 = (inp[8]) ? node65 : node62;
										assign node62 = (inp[1]) ? 3'b110 : 3'b010;
										assign node65 = (inp[1]) ? 3'b010 : 3'b110;
			assign node68 = (inp[4]) ? node90 : node69;
				assign node69 = (inp[7]) ? node73 : node70;
					assign node70 = (inp[6]) ? 3'b110 : 3'b000;
					assign node73 = (inp[6]) ? node75 : 3'b110;
						assign node75 = (inp[10]) ? node77 : 3'b000;
							assign node77 = (inp[5]) ? node79 : 3'b010;
								assign node79 = (inp[11]) ? node85 : node80;
									assign node80 = (inp[2]) ? node82 : 3'b000;
										assign node82 = (inp[1]) ? 3'b000 : 3'b010;
									assign node85 = (inp[0]) ? 3'b100 : node86;
										assign node86 = (inp[2]) ? 3'b010 : 3'b100;
				assign node90 = (inp[6]) ? node116 : node91;
					assign node91 = (inp[7]) ? node109 : node92;
						assign node92 = (inp[10]) ? node98 : node93;
							assign node93 = (inp[5]) ? node95 : 3'b010;
								assign node95 = (inp[11]) ? 3'b110 : 3'b010;
							assign node98 = (inp[0]) ? node104 : node99;
								assign node99 = (inp[8]) ? node101 : 3'b011;
									assign node101 = (inp[11]) ? 3'b101 : 3'b001;
								assign node104 = (inp[8]) ? node106 : 3'b101;
									assign node106 = (inp[11]) ? 3'b101 : 3'b001;
						assign node109 = (inp[11]) ? node111 : 3'b001;
							assign node111 = (inp[8]) ? node113 : 3'b001;
								assign node113 = (inp[10]) ? 3'b110 : 3'b001;
					assign node116 = (inp[11]) ? node118 : 3'b000;
						assign node118 = (inp[7]) ? 3'b000 : node119;
							assign node119 = (inp[10]) ? node121 : 3'b000;
								assign node121 = (inp[8]) ? 3'b100 : node122;
									assign node122 = (inp[2]) ? 3'b100 : 3'b010;

endmodule