module dtc_split5_bm72 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node9;
	wire [3-1:0] node12;
	wire [3-1:0] node13;
	wire [3-1:0] node16;
	wire [3-1:0] node19;
	wire [3-1:0] node20;
	wire [3-1:0] node21;
	wire [3-1:0] node24;
	wire [3-1:0] node27;
	wire [3-1:0] node28;
	wire [3-1:0] node31;
	wire [3-1:0] node34;
	wire [3-1:0] node35;
	wire [3-1:0] node36;
	wire [3-1:0] node37;
	wire [3-1:0] node40;
	wire [3-1:0] node43;
	wire [3-1:0] node44;
	wire [3-1:0] node47;
	wire [3-1:0] node50;
	wire [3-1:0] node51;
	wire [3-1:0] node52;
	wire [3-1:0] node55;
	wire [3-1:0] node58;
	wire [3-1:0] node59;
	wire [3-1:0] node62;
	wire [3-1:0] node65;
	wire [3-1:0] node66;
	wire [3-1:0] node67;
	wire [3-1:0] node68;
	wire [3-1:0] node70;
	wire [3-1:0] node73;
	wire [3-1:0] node74;
	wire [3-1:0] node77;
	wire [3-1:0] node80;
	wire [3-1:0] node81;
	wire [3-1:0] node82;
	wire [3-1:0] node85;
	wire [3-1:0] node88;
	wire [3-1:0] node89;
	wire [3-1:0] node92;
	wire [3-1:0] node95;
	wire [3-1:0] node96;
	wire [3-1:0] node97;
	wire [3-1:0] node98;
	wire [3-1:0] node101;
	wire [3-1:0] node104;
	wire [3-1:0] node105;
	wire [3-1:0] node108;
	wire [3-1:0] node111;
	wire [3-1:0] node112;
	wire [3-1:0] node113;
	wire [3-1:0] node116;
	wire [3-1:0] node119;
	wire [3-1:0] node120;
	wire [3-1:0] node123;
	wire [3-1:0] node126;
	wire [3-1:0] node127;
	wire [3-1:0] node128;
	wire [3-1:0] node129;
	wire [3-1:0] node130;
	wire [3-1:0] node131;
	wire [3-1:0] node134;
	wire [3-1:0] node137;
	wire [3-1:0] node138;
	wire [3-1:0] node141;
	wire [3-1:0] node144;
	wire [3-1:0] node145;
	wire [3-1:0] node146;
	wire [3-1:0] node149;
	wire [3-1:0] node152;
	wire [3-1:0] node153;
	wire [3-1:0] node157;
	wire [3-1:0] node158;
	wire [3-1:0] node159;
	wire [3-1:0] node160;
	wire [3-1:0] node163;
	wire [3-1:0] node166;
	wire [3-1:0] node167;
	wire [3-1:0] node171;
	wire [3-1:0] node172;
	wire [3-1:0] node174;
	wire [3-1:0] node178;
	wire [3-1:0] node179;
	wire [3-1:0] node180;
	wire [3-1:0] node181;
	wire [3-1:0] node182;
	wire [3-1:0] node185;
	wire [3-1:0] node188;
	wire [3-1:0] node189;
	wire [3-1:0] node192;
	wire [3-1:0] node195;
	wire [3-1:0] node196;
	wire [3-1:0] node197;
	wire [3-1:0] node200;
	wire [3-1:0] node203;
	wire [3-1:0] node204;
	wire [3-1:0] node207;
	wire [3-1:0] node210;
	wire [3-1:0] node211;
	wire [3-1:0] node212;
	wire [3-1:0] node213;
	wire [3-1:0] node216;
	wire [3-1:0] node219;
	wire [3-1:0] node220;
	wire [3-1:0] node223;
	wire [3-1:0] node226;
	wire [3-1:0] node227;
	wire [3-1:0] node228;
	wire [3-1:0] node231;
	wire [3-1:0] node234;
	wire [3-1:0] node235;
	wire [3-1:0] node238;

	assign outp = (inp[3]) ? node126 : node1;
		assign node1 = (inp[6]) ? node65 : node2;
			assign node2 = (inp[9]) ? node34 : node3;
				assign node3 = (inp[0]) ? node19 : node4;
					assign node4 = (inp[7]) ? node12 : node5;
						assign node5 = (inp[4]) ? node9 : node6;
							assign node6 = (inp[8]) ? 3'b001 : 3'b101;
							assign node9 = (inp[10]) ? 3'b010 : 3'b110;
						assign node12 = (inp[4]) ? node16 : node13;
							assign node13 = (inp[10]) ? 3'b001 : 3'b111;
							assign node16 = (inp[1]) ? 3'b001 : 3'b001;
					assign node19 = (inp[4]) ? node27 : node20;
						assign node20 = (inp[10]) ? node24 : node21;
							assign node21 = (inp[7]) ? 3'b101 : 3'b001;
							assign node24 = (inp[7]) ? 3'b010 : 3'b110;
						assign node27 = (inp[7]) ? node31 : node28;
							assign node28 = (inp[1]) ? 3'b000 : 3'b010;
							assign node31 = (inp[5]) ? 3'b110 : 3'b110;
				assign node34 = (inp[0]) ? node50 : node35;
					assign node35 = (inp[4]) ? node43 : node36;
						assign node36 = (inp[7]) ? node40 : node37;
							assign node37 = (inp[2]) ? 3'b110 : 3'b010;
							assign node40 = (inp[1]) ? 3'b110 : 3'b001;
						assign node43 = (inp[5]) ? node47 : node44;
							assign node44 = (inp[10]) ? 3'b010 : 3'b010;
							assign node47 = (inp[7]) ? 3'b110 : 3'b000;
					assign node50 = (inp[4]) ? node58 : node51;
						assign node51 = (inp[7]) ? node55 : node52;
							assign node52 = (inp[5]) ? 3'b000 : 3'b000;
							assign node55 = (inp[10]) ? 3'b010 : 3'b110;
						assign node58 = (inp[7]) ? node62 : node59;
							assign node59 = (inp[2]) ? 3'b000 : 3'b000;
							assign node62 = (inp[5]) ? 3'b000 : 3'b100;
			assign node65 = (inp[9]) ? node95 : node66;
				assign node66 = (inp[0]) ? node80 : node67;
					assign node67 = (inp[4]) ? node73 : node68;
						assign node68 = (inp[1]) ? node70 : 3'b111;
							assign node70 = (inp[10]) ? 3'b111 : 3'b111;
						assign node73 = (inp[7]) ? node77 : node74;
							assign node74 = (inp[1]) ? 3'b001 : 3'b111;
							assign node77 = (inp[10]) ? 3'b111 : 3'b111;
					assign node80 = (inp[7]) ? node88 : node81;
						assign node81 = (inp[4]) ? node85 : node82;
							assign node82 = (inp[8]) ? 3'b011 : 3'b101;
							assign node85 = (inp[11]) ? 3'b101 : 3'b101;
						assign node88 = (inp[4]) ? node92 : node89;
							assign node89 = (inp[10]) ? 3'b111 : 3'b111;
							assign node92 = (inp[1]) ? 3'b101 : 3'b011;
				assign node95 = (inp[0]) ? node111 : node96;
					assign node96 = (inp[4]) ? node104 : node97;
						assign node97 = (inp[7]) ? node101 : node98;
							assign node98 = (inp[5]) ? 3'b101 : 3'b011;
							assign node101 = (inp[1]) ? 3'b011 : 3'b111;
						assign node104 = (inp[11]) ? node108 : node105;
							assign node105 = (inp[7]) ? 3'b001 : 3'b001;
							assign node108 = (inp[7]) ? 3'b101 : 3'b001;
					assign node111 = (inp[4]) ? node119 : node112;
						assign node112 = (inp[10]) ? node116 : node113;
							assign node113 = (inp[7]) ? 3'b001 : 3'b001;
							assign node116 = (inp[1]) ? 3'b110 : 3'b001;
						assign node119 = (inp[7]) ? node123 : node120;
							assign node120 = (inp[10]) ? 3'b110 : 3'b110;
							assign node123 = (inp[8]) ? 3'b001 : 3'b110;
		assign node126 = (inp[6]) ? node178 : node127;
			assign node127 = (inp[9]) ? node157 : node128;
				assign node128 = (inp[0]) ? node144 : node129;
					assign node129 = (inp[4]) ? node137 : node130;
						assign node130 = (inp[10]) ? node134 : node131;
							assign node131 = (inp[7]) ? 3'b000 : 3'b010;
							assign node134 = (inp[7]) ? 3'b010 : 3'b100;
						assign node137 = (inp[7]) ? node141 : node138;
							assign node138 = (inp[5]) ? 3'b000 : 3'b100;
							assign node141 = (inp[1]) ? 3'b100 : 3'b010;
					assign node144 = (inp[4]) ? node152 : node145;
						assign node145 = (inp[10]) ? node149 : node146;
							assign node146 = (inp[7]) ? 3'b110 : 3'b000;
							assign node149 = (inp[7]) ? 3'b000 : 3'b000;
						assign node152 = (inp[10]) ? 3'b000 : node153;
							assign node153 = (inp[7]) ? 3'b000 : 3'b000;
				assign node157 = (inp[4]) ? node171 : node158;
					assign node158 = (inp[0]) ? node166 : node159;
						assign node159 = (inp[7]) ? node163 : node160;
							assign node160 = (inp[8]) ? 3'b000 : 3'b000;
							assign node163 = (inp[8]) ? 3'b010 : 3'b000;
						assign node166 = (inp[1]) ? 3'b000 : node167;
							assign node167 = (inp[2]) ? 3'b000 : 3'b000;
					assign node171 = (inp[10]) ? 3'b000 : node172;
						assign node172 = (inp[8]) ? node174 : 3'b000;
							assign node174 = (inp[0]) ? 3'b000 : 3'b000;
			assign node178 = (inp[9]) ? node210 : node179;
				assign node179 = (inp[0]) ? node195 : node180;
					assign node180 = (inp[7]) ? node188 : node181;
						assign node181 = (inp[4]) ? node185 : node182;
							assign node182 = (inp[10]) ? 3'b101 : 3'b001;
							assign node185 = (inp[8]) ? 3'b110 : 3'b010;
						assign node188 = (inp[4]) ? node192 : node189;
							assign node189 = (inp[10]) ? 3'b001 : 3'b111;
							assign node192 = (inp[8]) ? 3'b001 : 3'b001;
					assign node195 = (inp[7]) ? node203 : node196;
						assign node196 = (inp[4]) ? node200 : node197;
							assign node197 = (inp[10]) ? 3'b010 : 3'b110;
							assign node200 = (inp[10]) ? 3'b000 : 3'b000;
						assign node203 = (inp[4]) ? node207 : node204;
							assign node204 = (inp[10]) ? 3'b010 : 3'b001;
							assign node207 = (inp[10]) ? 3'b010 : 3'b110;
				assign node210 = (inp[0]) ? node226 : node211;
					assign node211 = (inp[4]) ? node219 : node212;
						assign node212 = (inp[7]) ? node216 : node213;
							assign node213 = (inp[1]) ? 3'b010 : 3'b110;
							assign node216 = (inp[10]) ? 3'b010 : 3'b001;
						assign node219 = (inp[7]) ? node223 : node220;
							assign node220 = (inp[10]) ? 3'b000 : 3'b100;
							assign node223 = (inp[1]) ? 3'b110 : 3'b110;
					assign node226 = (inp[7]) ? node234 : node227;
						assign node227 = (inp[4]) ? node231 : node228;
							assign node228 = (inp[10]) ? 3'b000 : 3'b100;
							assign node231 = (inp[5]) ? 3'b000 : 3'b000;
						assign node234 = (inp[4]) ? node238 : node235;
							assign node235 = (inp[5]) ? 3'b000 : 3'b010;
							assign node238 = (inp[10]) ? 3'b000 : 3'b100;

endmodule