module dtc_split66_bm53 (
	input  wire [8-1:0] inp,
	output wire [2-1:0] outp
);

	wire [2-1:0] node1;
	wire [2-1:0] node2;
	wire [2-1:0] node3;
	wire [2-1:0] node4;
	wire [2-1:0] node5;
	wire [2-1:0] node7;
	wire [2-1:0] node10;
	wire [2-1:0] node12;
	wire [2-1:0] node15;
	wire [2-1:0] node17;
	wire [2-1:0] node18;
	wire [2-1:0] node21;
	wire [2-1:0] node23;
	wire [2-1:0] node27;
	wire [2-1:0] node28;
	wire [2-1:0] node29;
	wire [2-1:0] node31;
	wire [2-1:0] node32;
	wire [2-1:0] node36;
	wire [2-1:0] node37;
	wire [2-1:0] node38;
	wire [2-1:0] node41;
	wire [2-1:0] node45;
	wire [2-1:0] node46;
	wire [2-1:0] node47;
	wire [2-1:0] node52;
	wire [2-1:0] node53;
	wire [2-1:0] node54;
	wire [2-1:0] node55;
	wire [2-1:0] node56;
	wire [2-1:0] node59;
	wire [2-1:0] node60;
	wire [2-1:0] node61;
	wire [2-1:0] node66;
	wire [2-1:0] node68;
	wire [2-1:0] node71;
	wire [2-1:0] node72;
	wire [2-1:0] node73;
	wire [2-1:0] node75;
	wire [2-1:0] node78;
	wire [2-1:0] node79;
	wire [2-1:0] node83;
	wire [2-1:0] node85;
	wire [2-1:0] node86;
	wire [2-1:0] node88;

	assign outp = (inp[6]) ? node52 : node1;
		assign node1 = (inp[7]) ? node27 : node2;
			assign node2 = (inp[3]) ? 2'b01 : node3;
				assign node3 = (inp[0]) ? node15 : node4;
					assign node4 = (inp[2]) ? node10 : node5;
						assign node5 = (inp[4]) ? node7 : 2'b00;
							assign node7 = (inp[1]) ? 2'b01 : 2'b00;
						assign node10 = (inp[4]) ? node12 : 2'b01;
							assign node12 = (inp[5]) ? 2'b01 : 2'b00;
					assign node15 = (inp[1]) ? node17 : 2'b11;
						assign node17 = (inp[2]) ? node21 : node18;
							assign node18 = (inp[5]) ? 2'b00 : 2'b11;
							assign node21 = (inp[4]) ? node23 : 2'b01;
								assign node23 = (inp[5]) ? 2'b01 : 2'b00;
			assign node27 = (inp[1]) ? node45 : node28;
				assign node28 = (inp[5]) ? node36 : node29;
					assign node29 = (inp[0]) ? node31 : 2'b00;
						assign node31 = (inp[3]) ? 2'b01 : node32;
							assign node32 = (inp[4]) ? 2'b01 : 2'b00;
					assign node36 = (inp[2]) ? 2'b01 : node37;
						assign node37 = (inp[0]) ? node41 : node38;
							assign node38 = (inp[3]) ? 2'b00 : 2'b01;
							assign node41 = (inp[3]) ? 2'b01 : 2'b00;
				assign node45 = (inp[5]) ? 2'b00 : node46;
					assign node46 = (inp[3]) ? 2'b00 : node47;
						assign node47 = (inp[4]) ? 2'b00 : 2'b01;
		assign node52 = (inp[3]) ? 2'b00 : node53;
			assign node53 = (inp[7]) ? node71 : node54;
				assign node54 = (inp[0]) ? node66 : node55;
					assign node55 = (inp[1]) ? node59 : node56;
						assign node56 = (inp[2]) ? 2'b00 : 2'b10;
						assign node59 = (inp[2]) ? 2'b00 : node60;
							assign node60 = (inp[5]) ? 2'b01 : node61;
								assign node61 = (inp[4]) ? 2'b00 : 2'b01;
					assign node66 = (inp[2]) ? node68 : 2'b10;
						assign node68 = (inp[1]) ? 2'b00 : 2'b10;
				assign node71 = (inp[1]) ? node83 : node72;
					assign node72 = (inp[5]) ? node78 : node73;
						assign node73 = (inp[4]) ? node75 : 2'b01;
							assign node75 = (inp[2]) ? 2'b01 : 2'b00;
						assign node78 = (inp[2]) ? 2'b00 : node79;
							assign node79 = (inp[0]) ? 2'b01 : 2'b00;
					assign node83 = (inp[4]) ? node85 : 2'b00;
						assign node85 = (inp[5]) ? 2'b00 : node86;
							assign node86 = (inp[0]) ? node88 : 2'b00;
								assign node88 = (inp[2]) ? 2'b00 : 2'b01;

endmodule