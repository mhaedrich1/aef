module dtc_split66_bm89 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node7;
	wire [3-1:0] node8;
	wire [3-1:0] node10;
	wire [3-1:0] node12;
	wire [3-1:0] node15;
	wire [3-1:0] node16;
	wire [3-1:0] node18;
	wire [3-1:0] node22;
	wire [3-1:0] node24;
	wire [3-1:0] node25;
	wire [3-1:0] node30;
	wire [3-1:0] node31;
	wire [3-1:0] node32;
	wire [3-1:0] node34;
	wire [3-1:0] node35;
	wire [3-1:0] node39;
	wire [3-1:0] node41;
	wire [3-1:0] node42;
	wire [3-1:0] node43;
	wire [3-1:0] node48;
	wire [3-1:0] node49;
	wire [3-1:0] node50;
	wire [3-1:0] node51;
	wire [3-1:0] node53;
	wire [3-1:0] node56;
	wire [3-1:0] node58;
	wire [3-1:0] node61;
	wire [3-1:0] node62;
	wire [3-1:0] node64;
	wire [3-1:0] node67;
	wire [3-1:0] node69;
	wire [3-1:0] node72;
	wire [3-1:0] node73;
	wire [3-1:0] node74;
	wire [3-1:0] node77;
	wire [3-1:0] node79;
	wire [3-1:0] node82;
	wire [3-1:0] node83;
	wire [3-1:0] node86;
	wire [3-1:0] node88;
	wire [3-1:0] node92;
	wire [3-1:0] node93;
	wire [3-1:0] node94;
	wire [3-1:0] node95;
	wire [3-1:0] node96;
	wire [3-1:0] node97;
	wire [3-1:0] node98;
	wire [3-1:0] node100;
	wire [3-1:0] node103;
	wire [3-1:0] node105;
	wire [3-1:0] node108;
	wire [3-1:0] node110;
	wire [3-1:0] node112;
	wire [3-1:0] node115;
	wire [3-1:0] node116;
	wire [3-1:0] node118;
	wire [3-1:0] node120;
	wire [3-1:0] node124;
	wire [3-1:0] node125;
	wire [3-1:0] node126;
	wire [3-1:0] node127;
	wire [3-1:0] node129;
	wire [3-1:0] node132;
	wire [3-1:0] node135;
	wire [3-1:0] node136;
	wire [3-1:0] node137;
	wire [3-1:0] node139;
	wire [3-1:0] node142;
	wire [3-1:0] node144;
	wire [3-1:0] node147;
	wire [3-1:0] node149;
	wire [3-1:0] node152;
	wire [3-1:0] node153;
	wire [3-1:0] node154;
	wire [3-1:0] node156;
	wire [3-1:0] node159;
	wire [3-1:0] node161;
	wire [3-1:0] node164;
	wire [3-1:0] node165;
	wire [3-1:0] node169;
	wire [3-1:0] node170;
	wire [3-1:0] node171;
	wire [3-1:0] node172;
	wire [3-1:0] node175;
	wire [3-1:0] node177;
	wire [3-1:0] node178;
	wire [3-1:0] node181;
	wire [3-1:0] node184;
	wire [3-1:0] node185;
	wire [3-1:0] node186;
	wire [3-1:0] node187;
	wire [3-1:0] node190;
	wire [3-1:0] node193;
	wire [3-1:0] node195;
	wire [3-1:0] node196;
	wire [3-1:0] node200;
	wire [3-1:0] node202;
	wire [3-1:0] node203;
	wire [3-1:0] node206;
	wire [3-1:0] node209;
	wire [3-1:0] node210;
	wire [3-1:0] node213;
	wire [3-1:0] node214;
	wire [3-1:0] node217;
	wire [3-1:0] node218;
	wire [3-1:0] node219;
	wire [3-1:0] node220;
	wire [3-1:0] node225;
	wire [3-1:0] node228;
	wire [3-1:0] node229;
	wire [3-1:0] node230;
	wire [3-1:0] node231;
	wire [3-1:0] node232;
	wire [3-1:0] node233;
	wire [3-1:0] node234;
	wire [3-1:0] node238;
	wire [3-1:0] node239;
	wire [3-1:0] node243;
	wire [3-1:0] node244;
	wire [3-1:0] node246;
	wire [3-1:0] node250;
	wire [3-1:0] node251;
	wire [3-1:0] node252;
	wire [3-1:0] node254;
	wire [3-1:0] node257;
	wire [3-1:0] node259;
	wire [3-1:0] node262;
	wire [3-1:0] node263;
	wire [3-1:0] node264;
	wire [3-1:0] node267;
	wire [3-1:0] node269;
	wire [3-1:0] node274;
	wire [3-1:0] node275;
	wire [3-1:0] node276;
	wire [3-1:0] node277;
	wire [3-1:0] node279;
	wire [3-1:0] node282;
	wire [3-1:0] node285;
	wire [3-1:0] node286;
	wire [3-1:0] node288;
	wire [3-1:0] node291;
	wire [3-1:0] node292;
	wire [3-1:0] node294;
	wire [3-1:0] node297;
	wire [3-1:0] node299;
	wire [3-1:0] node302;
	wire [3-1:0] node303;
	wire [3-1:0] node304;
	wire [3-1:0] node305;
	wire [3-1:0] node307;
	wire [3-1:0] node310;
	wire [3-1:0] node311;
	wire [3-1:0] node315;
	wire [3-1:0] node317;
	wire [3-1:0] node320;
	wire [3-1:0] node321;
	wire [3-1:0] node323;
	wire [3-1:0] node326;
	wire [3-1:0] node328;
	wire [3-1:0] node331;
	wire [3-1:0] node332;
	wire [3-1:0] node333;
	wire [3-1:0] node334;
	wire [3-1:0] node335;
	wire [3-1:0] node336;
	wire [3-1:0] node337;
	wire [3-1:0] node338;
	wire [3-1:0] node343;
	wire [3-1:0] node344;
	wire [3-1:0] node345;
	wire [3-1:0] node346;
	wire [3-1:0] node350;
	wire [3-1:0] node352;
	wire [3-1:0] node355;
	wire [3-1:0] node356;
	wire [3-1:0] node358;
	wire [3-1:0] node361;
	wire [3-1:0] node366;
	wire [3-1:0] node367;
	wire [3-1:0] node368;
	wire [3-1:0] node369;
	wire [3-1:0] node370;
	wire [3-1:0] node372;
	wire [3-1:0] node373;
	wire [3-1:0] node374;
	wire [3-1:0] node378;
	wire [3-1:0] node381;
	wire [3-1:0] node383;
	wire [3-1:0] node385;
	wire [3-1:0] node387;
	wire [3-1:0] node390;
	wire [3-1:0] node391;
	wire [3-1:0] node393;
	wire [3-1:0] node395;
	wire [3-1:0] node399;
	wire [3-1:0] node400;
	wire [3-1:0] node401;
	wire [3-1:0] node402;
	wire [3-1:0] node404;
	wire [3-1:0] node407;
	wire [3-1:0] node408;
	wire [3-1:0] node410;
	wire [3-1:0] node413;
	wire [3-1:0] node415;
	wire [3-1:0] node418;
	wire [3-1:0] node419;
	wire [3-1:0] node420;
	wire [3-1:0] node424;
	wire [3-1:0] node426;
	wire [3-1:0] node428;
	wire [3-1:0] node431;
	wire [3-1:0] node432;
	wire [3-1:0] node433;
	wire [3-1:0] node434;
	wire [3-1:0] node439;
	wire [3-1:0] node440;
	wire [3-1:0] node441;
	wire [3-1:0] node442;
	wire [3-1:0] node446;
	wire [3-1:0] node449;
	wire [3-1:0] node450;
	wire [3-1:0] node452;
	wire [3-1:0] node456;
	wire [3-1:0] node457;
	wire [3-1:0] node458;
	wire [3-1:0] node459;
	wire [3-1:0] node461;
	wire [3-1:0] node463;
	wire [3-1:0] node464;
	wire [3-1:0] node469;
	wire [3-1:0] node470;
	wire [3-1:0] node471;
	wire [3-1:0] node473;
	wire [3-1:0] node477;
	wire [3-1:0] node478;
	wire [3-1:0] node480;
	wire [3-1:0] node485;
	wire [3-1:0] node486;
	wire [3-1:0] node487;
	wire [3-1:0] node488;
	wire [3-1:0] node489;
	wire [3-1:0] node490;
	wire [3-1:0] node492;
	wire [3-1:0] node494;
	wire [3-1:0] node497;
	wire [3-1:0] node498;
	wire [3-1:0] node500;
	wire [3-1:0] node503;
	wire [3-1:0] node505;
	wire [3-1:0] node508;
	wire [3-1:0] node510;
	wire [3-1:0] node511;
	wire [3-1:0] node516;
	wire [3-1:0] node517;
	wire [3-1:0] node518;
	wire [3-1:0] node519;
	wire [3-1:0] node521;
	wire [3-1:0] node523;
	wire [3-1:0] node526;
	wire [3-1:0] node527;
	wire [3-1:0] node530;
	wire [3-1:0] node533;
	wire [3-1:0] node534;
	wire [3-1:0] node535;
	wire [3-1:0] node536;
	wire [3-1:0] node540;
	wire [3-1:0] node541;
	wire [3-1:0] node544;
	wire [3-1:0] node545;
	wire [3-1:0] node549;
	wire [3-1:0] node550;
	wire [3-1:0] node551;
	wire [3-1:0] node553;
	wire [3-1:0] node556;
	wire [3-1:0] node558;
	wire [3-1:0] node561;
	wire [3-1:0] node563;
	wire [3-1:0] node566;
	wire [3-1:0] node567;
	wire [3-1:0] node569;
	wire [3-1:0] node571;
	wire [3-1:0] node573;
	wire [3-1:0] node576;
	wire [3-1:0] node577;
	wire [3-1:0] node580;
	wire [3-1:0] node582;
	wire [3-1:0] node585;
	wire [3-1:0] node586;
	wire [3-1:0] node587;
	wire [3-1:0] node588;
	wire [3-1:0] node590;
	wire [3-1:0] node593;
	wire [3-1:0] node595;
	wire [3-1:0] node596;
	wire [3-1:0] node598;
	wire [3-1:0] node602;
	wire [3-1:0] node603;
	wire [3-1:0] node604;
	wire [3-1:0] node605;
	wire [3-1:0] node608;
	wire [3-1:0] node610;
	wire [3-1:0] node613;
	wire [3-1:0] node615;
	wire [3-1:0] node618;
	wire [3-1:0] node619;
	wire [3-1:0] node621;
	wire [3-1:0] node623;
	wire [3-1:0] node626;
	wire [3-1:0] node627;
	wire [3-1:0] node630;
	wire [3-1:0] node633;
	wire [3-1:0] node634;
	wire [3-1:0] node635;
	wire [3-1:0] node636;
	wire [3-1:0] node638;
	wire [3-1:0] node639;
	wire [3-1:0] node640;
	wire [3-1:0] node644;
	wire [3-1:0] node645;
	wire [3-1:0] node649;
	wire [3-1:0] node651;
	wire [3-1:0] node654;
	wire [3-1:0] node655;
	wire [3-1:0] node656;
	wire [3-1:0] node658;
	wire [3-1:0] node660;
	wire [3-1:0] node663;
	wire [3-1:0] node664;
	wire [3-1:0] node668;
	wire [3-1:0] node671;
	wire [3-1:0] node672;
	wire [3-1:0] node673;
	wire [3-1:0] node675;
	wire [3-1:0] node678;
	wire [3-1:0] node679;
	wire [3-1:0] node680;
	wire [3-1:0] node684;
	wire [3-1:0] node685;
	wire [3-1:0] node688;
	wire [3-1:0] node691;
	wire [3-1:0] node693;
	wire [3-1:0] node694;
	wire [3-1:0] node696;
	wire [3-1:0] node699;
	wire [3-1:0] node701;
	wire [3-1:0] node703;
	wire [3-1:0] node706;
	wire [3-1:0] node707;
	wire [3-1:0] node708;
	wire [3-1:0] node709;
	wire [3-1:0] node710;
	wire [3-1:0] node711;
	wire [3-1:0] node712;
	wire [3-1:0] node713;
	wire [3-1:0] node715;
	wire [3-1:0] node718;
	wire [3-1:0] node719;
	wire [3-1:0] node721;
	wire [3-1:0] node724;
	wire [3-1:0] node725;
	wire [3-1:0] node729;
	wire [3-1:0] node731;
	wire [3-1:0] node732;
	wire [3-1:0] node736;
	wire [3-1:0] node737;
	wire [3-1:0] node738;
	wire [3-1:0] node739;
	wire [3-1:0] node741;
	wire [3-1:0] node744;
	wire [3-1:0] node746;
	wire [3-1:0] node749;
	wire [3-1:0] node750;
	wire [3-1:0] node752;
	wire [3-1:0] node755;
	wire [3-1:0] node757;
	wire [3-1:0] node760;
	wire [3-1:0] node761;
	wire [3-1:0] node762;
	wire [3-1:0] node765;
	wire [3-1:0] node766;
	wire [3-1:0] node769;
	wire [3-1:0] node772;
	wire [3-1:0] node773;
	wire [3-1:0] node775;
	wire [3-1:0] node777;
	wire [3-1:0] node780;
	wire [3-1:0] node782;
	wire [3-1:0] node785;
	wire [3-1:0] node787;
	wire [3-1:0] node788;
	wire [3-1:0] node789;
	wire [3-1:0] node791;
	wire [3-1:0] node794;
	wire [3-1:0] node796;
	wire [3-1:0] node799;
	wire [3-1:0] node800;
	wire [3-1:0] node801;
	wire [3-1:0] node802;
	wire [3-1:0] node806;
	wire [3-1:0] node808;
	wire [3-1:0] node811;
	wire [3-1:0] node812;
	wire [3-1:0] node815;
	wire [3-1:0] node817;
	wire [3-1:0] node820;
	wire [3-1:0] node822;
	wire [3-1:0] node824;
	wire [3-1:0] node825;
	wire [3-1:0] node827;
	wire [3-1:0] node832;
	wire [3-1:0] node833;
	wire [3-1:0] node834;
	wire [3-1:0] node835;
	wire [3-1:0] node836;
	wire [3-1:0] node837;
	wire [3-1:0] node838;
	wire [3-1:0] node840;
	wire [3-1:0] node842;
	wire [3-1:0] node845;
	wire [3-1:0] node846;
	wire [3-1:0] node848;
	wire [3-1:0] node852;
	wire [3-1:0] node854;
	wire [3-1:0] node855;
	wire [3-1:0] node860;
	wire [3-1:0] node861;
	wire [3-1:0] node862;
	wire [3-1:0] node863;
	wire [3-1:0] node864;
	wire [3-1:0] node867;
	wire [3-1:0] node868;
	wire [3-1:0] node869;
	wire [3-1:0] node872;
	wire [3-1:0] node876;
	wire [3-1:0] node877;
	wire [3-1:0] node881;
	wire [3-1:0] node882;
	wire [3-1:0] node883;
	wire [3-1:0] node885;
	wire [3-1:0] node888;
	wire [3-1:0] node891;
	wire [3-1:0] node892;
	wire [3-1:0] node893;
	wire [3-1:0] node896;
	wire [3-1:0] node898;
	wire [3-1:0] node901;
	wire [3-1:0] node903;
	wire [3-1:0] node905;
	wire [3-1:0] node908;
	wire [3-1:0] node909;
	wire [3-1:0] node910;
	wire [3-1:0] node911;
	wire [3-1:0] node914;
	wire [3-1:0] node916;
	wire [3-1:0] node919;
	wire [3-1:0] node920;
	wire [3-1:0] node924;
	wire [3-1:0] node925;
	wire [3-1:0] node926;
	wire [3-1:0] node927;
	wire [3-1:0] node930;
	wire [3-1:0] node933;
	wire [3-1:0] node936;
	wire [3-1:0] node937;
	wire [3-1:0] node938;
	wire [3-1:0] node941;
	wire [3-1:0] node943;
	wire [3-1:0] node946;
	wire [3-1:0] node947;
	wire [3-1:0] node951;
	wire [3-1:0] node952;
	wire [3-1:0] node953;
	wire [3-1:0] node954;
	wire [3-1:0] node956;
	wire [3-1:0] node957;
	wire [3-1:0] node958;
	wire [3-1:0] node963;
	wire [3-1:0] node965;
	wire [3-1:0] node968;
	wire [3-1:0] node969;
	wire [3-1:0] node970;
	wire [3-1:0] node971;
	wire [3-1:0] node975;
	wire [3-1:0] node976;
	wire [3-1:0] node979;
	wire [3-1:0] node980;
	wire [3-1:0] node984;
	wire [3-1:0] node986;
	wire [3-1:0] node987;
	wire [3-1:0] node988;
	wire [3-1:0] node991;
	wire [3-1:0] node994;
	wire [3-1:0] node995;
	wire [3-1:0] node998;
	wire [3-1:0] node1001;
	wire [3-1:0] node1002;
	wire [3-1:0] node1003;
	wire [3-1:0] node1004;
	wire [3-1:0] node1006;
	wire [3-1:0] node1007;
	wire [3-1:0] node1009;
	wire [3-1:0] node1012;
	wire [3-1:0] node1013;
	wire [3-1:0] node1017;
	wire [3-1:0] node1019;
	wire [3-1:0] node1022;
	wire [3-1:0] node1023;
	wire [3-1:0] node1025;
	wire [3-1:0] node1026;
	wire [3-1:0] node1028;
	wire [3-1:0] node1032;
	wire [3-1:0] node1034;
	wire [3-1:0] node1037;
	wire [3-1:0] node1038;
	wire [3-1:0] node1039;
	wire [3-1:0] node1041;
	wire [3-1:0] node1044;
	wire [3-1:0] node1045;
	wire [3-1:0] node1047;
	wire [3-1:0] node1051;
	wire [3-1:0] node1052;
	wire [3-1:0] node1054;
	wire [3-1:0] node1055;
	wire [3-1:0] node1059;
	wire [3-1:0] node1060;
	wire [3-1:0] node1063;
	wire [3-1:0] node1064;
	wire [3-1:0] node1065;
	wire [3-1:0] node1070;
	wire [3-1:0] node1071;
	wire [3-1:0] node1072;
	wire [3-1:0] node1073;
	wire [3-1:0] node1074;
	wire [3-1:0] node1075;
	wire [3-1:0] node1077;
	wire [3-1:0] node1081;
	wire [3-1:0] node1082;
	wire [3-1:0] node1084;
	wire [3-1:0] node1086;
	wire [3-1:0] node1089;
	wire [3-1:0] node1090;
	wire [3-1:0] node1093;
	wire [3-1:0] node1095;
	wire [3-1:0] node1100;
	wire [3-1:0] node1101;
	wire [3-1:0] node1102;
	wire [3-1:0] node1103;
	wire [3-1:0] node1104;
	wire [3-1:0] node1105;
	wire [3-1:0] node1108;
	wire [3-1:0] node1110;
	wire [3-1:0] node1113;
	wire [3-1:0] node1114;
	wire [3-1:0] node1117;
	wire [3-1:0] node1119;
	wire [3-1:0] node1121;
	wire [3-1:0] node1124;
	wire [3-1:0] node1125;
	wire [3-1:0] node1126;
	wire [3-1:0] node1128;
	wire [3-1:0] node1131;
	wire [3-1:0] node1132;
	wire [3-1:0] node1135;
	wire [3-1:0] node1136;
	wire [3-1:0] node1140;
	wire [3-1:0] node1141;
	wire [3-1:0] node1143;
	wire [3-1:0] node1145;
	wire [3-1:0] node1148;
	wire [3-1:0] node1150;
	wire [3-1:0] node1153;
	wire [3-1:0] node1154;
	wire [3-1:0] node1155;
	wire [3-1:0] node1157;
	wire [3-1:0] node1161;
	wire [3-1:0] node1162;
	wire [3-1:0] node1163;
	wire [3-1:0] node1165;
	wire [3-1:0] node1169;
	wire [3-1:0] node1170;
	wire [3-1:0] node1171;
	wire [3-1:0] node1176;
	wire [3-1:0] node1177;
	wire [3-1:0] node1178;
	wire [3-1:0] node1179;
	wire [3-1:0] node1181;
	wire [3-1:0] node1183;
	wire [3-1:0] node1184;
	wire [3-1:0] node1189;
	wire [3-1:0] node1190;
	wire [3-1:0] node1191;
	wire [3-1:0] node1192;
	wire [3-1:0] node1193;
	wire [3-1:0] node1197;
	wire [3-1:0] node1199;
	wire [3-1:0] node1203;
	wire [3-1:0] node1204;
	wire [3-1:0] node1206;
	wire [3-1:0] node1209;
	wire [3-1:0] node1211;
	wire [3-1:0] node1214;
	wire [3-1:0] node1215;
	wire [3-1:0] node1216;
	wire [3-1:0] node1217;

	assign outp = (inp[3]) ? node706 : node1;
		assign node1 = (inp[6]) ? node331 : node2;
			assign node2 = (inp[7]) ? node92 : node3;
				assign node3 = (inp[9]) ? 3'b111 : node4;
					assign node4 = (inp[4]) ? node30 : node5;
						assign node5 = (inp[10]) ? 3'b111 : node6;
							assign node6 = (inp[5]) ? node22 : node7;
								assign node7 = (inp[8]) ? node15 : node8;
									assign node8 = (inp[0]) ? node10 : 3'b101;
										assign node10 = (inp[2]) ? node12 : 3'b101;
											assign node12 = (inp[11]) ? 3'b011 : 3'b101;
									assign node15 = (inp[11]) ? 3'b011 : node16;
										assign node16 = (inp[0]) ? node18 : 3'b101;
											assign node18 = (inp[1]) ? 3'b011 : 3'b101;
								assign node22 = (inp[11]) ? node24 : 3'b011;
									assign node24 = (inp[2]) ? 3'b101 : node25;
										assign node25 = (inp[8]) ? 3'b101 : 3'b011;
						assign node30 = (inp[10]) ? node48 : node31;
							assign node31 = (inp[8]) ? node39 : node32;
								assign node32 = (inp[11]) ? node34 : 3'b010;
									assign node34 = (inp[0]) ? 3'b110 : node35;
										assign node35 = (inp[1]) ? 3'b110 : 3'b001;
								assign node39 = (inp[11]) ? node41 : 3'b100;
									assign node41 = (inp[1]) ? 3'b010 : node42;
										assign node42 = (inp[0]) ? 3'b110 : node43;
											assign node43 = (inp[2]) ? 3'b110 : 3'b101;
							assign node48 = (inp[2]) ? node72 : node49;
								assign node49 = (inp[8]) ? node61 : node50;
									assign node50 = (inp[11]) ? node56 : node51;
										assign node51 = (inp[5]) ? node53 : 3'b101;
											assign node53 = (inp[0]) ? 3'b001 : 3'b101;
										assign node56 = (inp[5]) ? node58 : 3'b011;
											assign node58 = (inp[0]) ? 3'b101 : 3'b011;
									assign node61 = (inp[11]) ? node67 : node62;
										assign node62 = (inp[5]) ? node64 : 3'b001;
											assign node64 = (inp[0]) ? 3'b110 : 3'b001;
										assign node67 = (inp[0]) ? node69 : 3'b101;
											assign node69 = (inp[5]) ? 3'b001 : 3'b101;
								assign node72 = (inp[8]) ? node82 : node73;
									assign node73 = (inp[11]) ? node77 : node74;
										assign node74 = (inp[1]) ? 3'b001 : 3'b101;
										assign node77 = (inp[0]) ? node79 : 3'b011;
											assign node79 = (inp[5]) ? 3'b101 : 3'b011;
									assign node82 = (inp[11]) ? node86 : node83;
										assign node83 = (inp[1]) ? 3'b110 : 3'b001;
										assign node86 = (inp[0]) ? node88 : 3'b101;
											assign node88 = (inp[5]) ? 3'b001 : 3'b101;
				assign node92 = (inp[10]) ? node228 : node93;
					assign node93 = (inp[4]) ? node169 : node94;
						assign node94 = (inp[11]) ? node124 : node95;
							assign node95 = (inp[5]) ? node115 : node96;
								assign node96 = (inp[9]) ? node108 : node97;
									assign node97 = (inp[0]) ? node103 : node98;
										assign node98 = (inp[8]) ? node100 : 3'b010;
											assign node100 = (inp[2]) ? 3'b010 : 3'b110;
										assign node103 = (inp[8]) ? node105 : 3'b110;
											assign node105 = (inp[2]) ? 3'b010 : 3'b110;
									assign node108 = (inp[8]) ? node110 : 3'b110;
										assign node110 = (inp[1]) ? node112 : 3'b110;
											assign node112 = (inp[0]) ? 3'b000 : 3'b110;
								assign node115 = (inp[9]) ? 3'b000 : node116;
									assign node116 = (inp[8]) ? node118 : 3'b110;
										assign node118 = (inp[1]) ? node120 : 3'b000;
											assign node120 = (inp[2]) ? 3'b100 : 3'b000;
							assign node124 = (inp[9]) ? node152 : node125;
								assign node125 = (inp[5]) ? node135 : node126;
									assign node126 = (inp[8]) ? node132 : node127;
										assign node127 = (inp[0]) ? node129 : 3'b111;
											assign node129 = (inp[2]) ? 3'b001 : 3'b011;
										assign node132 = (inp[2]) ? 3'b101 : 3'b001;
									assign node135 = (inp[8]) ? node147 : node136;
										assign node136 = (inp[2]) ? node142 : node137;
											assign node137 = (inp[0]) ? node139 : 3'b001;
												assign node139 = (inp[1]) ? 3'b100 : 3'b001;
											assign node142 = (inp[1]) ? node144 : 3'b011;
												assign node144 = (inp[0]) ? 3'b110 : 3'b011;
										assign node147 = (inp[1]) ? node149 : 3'b110;
											assign node149 = (inp[0]) ? 3'b010 : 3'b110;
								assign node152 = (inp[5]) ? node164 : node153;
									assign node153 = (inp[8]) ? node159 : node154;
										assign node154 = (inp[2]) ? node156 : 3'b110;
											assign node156 = (inp[0]) ? 3'b000 : 3'b110;
										assign node159 = (inp[2]) ? node161 : 3'b000;
											assign node161 = (inp[1]) ? 3'b110 : 3'b000;
									assign node164 = (inp[8]) ? 3'b110 : node165;
										assign node165 = (inp[2]) ? 3'b110 : 3'b000;
						assign node169 = (inp[9]) ? node209 : node170;
							assign node170 = (inp[8]) ? node184 : node171;
								assign node171 = (inp[11]) ? node175 : node172;
									assign node172 = (inp[5]) ? 3'b000 : 3'b100;
									assign node175 = (inp[5]) ? node177 : 3'b010;
										assign node177 = (inp[0]) ? node181 : node178;
											assign node178 = (inp[2]) ? 3'b100 : 3'b010;
											assign node181 = (inp[2]) ? 3'b010 : 3'b100;
								assign node184 = (inp[5]) ? node200 : node185;
									assign node185 = (inp[2]) ? node193 : node186;
										assign node186 = (inp[1]) ? node190 : node187;
											assign node187 = (inp[11]) ? 3'b000 : 3'b100;
											assign node190 = (inp[11]) ? 3'b100 : 3'b000;
										assign node193 = (inp[1]) ? node195 : 3'b100;
											assign node195 = (inp[11]) ? 3'b100 : node196;
												assign node196 = (inp[0]) ? 3'b000 : 3'b100;
									assign node200 = (inp[11]) ? node202 : 3'b000;
										assign node202 = (inp[2]) ? node206 : node203;
											assign node203 = (inp[1]) ? 3'b100 : 3'b000;
											assign node206 = (inp[1]) ? 3'b000 : 3'b100;
							assign node209 = (inp[8]) ? node213 : node210;
								assign node210 = (inp[11]) ? 3'b101 : 3'b001;
								assign node213 = (inp[11]) ? node217 : node214;
									assign node214 = (inp[5]) ? 3'b110 : 3'b111;
									assign node217 = (inp[1]) ? node225 : node218;
										assign node218 = (inp[5]) ? 3'b111 : node219;
											assign node219 = (inp[2]) ? 3'b100 : node220;
												assign node220 = (inp[0]) ? 3'b100 : 3'b110;
										assign node225 = (inp[5]) ? 3'b001 : 3'b000;
					assign node228 = (inp[4]) ? node274 : node229;
						assign node229 = (inp[9]) ? 3'b100 : node230;
							assign node230 = (inp[11]) ? node250 : node231;
								assign node231 = (inp[5]) ? node243 : node232;
									assign node232 = (inp[2]) ? node238 : node233;
										assign node233 = (inp[0]) ? 3'b101 : node234;
											assign node234 = (inp[8]) ? 3'b101 : 3'b001;
										assign node238 = (inp[8]) ? 3'b001 : node239;
											assign node239 = (inp[0]) ? 3'b101 : 3'b001;
									assign node243 = (inp[8]) ? 3'b010 : node244;
										assign node244 = (inp[1]) ? node246 : 3'b101;
											assign node246 = (inp[0]) ? 3'b001 : 3'b101;
								assign node250 = (inp[5]) ? node262 : node251;
									assign node251 = (inp[8]) ? node257 : node252;
										assign node252 = (inp[0]) ? node254 : 3'b101;
											assign node254 = (inp[1]) ? 3'b011 : 3'b001;
										assign node257 = (inp[2]) ? node259 : 3'b011;
											assign node259 = (inp[1]) ? 3'b101 : 3'b111;
									assign node262 = (inp[8]) ? 3'b101 : node263;
										assign node263 = (inp[2]) ? node267 : node264;
											assign node264 = (inp[0]) ? 3'b111 : 3'b011;
											assign node267 = (inp[1]) ? node269 : 3'b001;
												assign node269 = (inp[0]) ? 3'b101 : 3'b001;
						assign node274 = (inp[9]) ? node302 : node275;
							assign node275 = (inp[11]) ? node285 : node276;
								assign node276 = (inp[8]) ? node282 : node277;
									assign node277 = (inp[0]) ? node279 : 3'b110;
										assign node279 = (inp[5]) ? 3'b010 : 3'b110;
									assign node282 = (inp[0]) ? 3'b100 : 3'b010;
								assign node285 = (inp[8]) ? node291 : node286;
									assign node286 = (inp[0]) ? node288 : 3'b001;
										assign node288 = (inp[5]) ? 3'b110 : 3'b001;
									assign node291 = (inp[5]) ? node297 : node292;
										assign node292 = (inp[2]) ? node294 : 3'b001;
											assign node294 = (inp[0]) ? 3'b110 : 3'b010;
										assign node297 = (inp[1]) ? node299 : 3'b110;
											assign node299 = (inp[0]) ? 3'b010 : 3'b110;
							assign node302 = (inp[8]) ? node320 : node303;
								assign node303 = (inp[11]) ? node315 : node304;
									assign node304 = (inp[5]) ? node310 : node305;
										assign node305 = (inp[2]) ? node307 : 3'b111;
											assign node307 = (inp[0]) ? 3'b011 : 3'b111;
										assign node310 = (inp[0]) ? 3'b011 : node311;
											assign node311 = (inp[2]) ? 3'b011 : 3'b111;
									assign node315 = (inp[0]) ? node317 : 3'b001;
										assign node317 = (inp[5]) ? 3'b111 : 3'b001;
								assign node320 = (inp[11]) ? node326 : node321;
									assign node321 = (inp[1]) ? node323 : 3'b011;
										assign node323 = (inp[2]) ? 3'b101 : 3'b011;
									assign node326 = (inp[5]) ? node328 : 3'b111;
										assign node328 = (inp[0]) ? 3'b011 : 3'b111;
			assign node331 = (inp[9]) ? node485 : node332;
				assign node332 = (inp[10]) ? node366 : node333;
					assign node333 = (inp[7]) ? 3'b000 : node334;
						assign node334 = (inp[4]) ? 3'b000 : node335;
							assign node335 = (inp[11]) ? node343 : node336;
								assign node336 = (inp[8]) ? 3'b000 : node337;
									assign node337 = (inp[2]) ? 3'b100 : node338;
										assign node338 = (inp[0]) ? 3'b000 : 3'b100;
								assign node343 = (inp[5]) ? node355 : node344;
									assign node344 = (inp[2]) ? node350 : node345;
										assign node345 = (inp[0]) ? 3'b010 : node346;
											assign node346 = (inp[8]) ? 3'b010 : 3'b110;
										assign node350 = (inp[0]) ? node352 : 3'b110;
											assign node352 = (inp[1]) ? 3'b100 : 3'b110;
									assign node355 = (inp[8]) ? node361 : node356;
										assign node356 = (inp[1]) ? node358 : 3'b010;
											assign node358 = (inp[0]) ? 3'b100 : 3'b010;
										assign node361 = (inp[2]) ? 3'b000 : 3'b100;
					assign node366 = (inp[4]) ? node456 : node367;
						assign node367 = (inp[11]) ? node399 : node368;
							assign node368 = (inp[7]) ? node390 : node369;
								assign node369 = (inp[2]) ? node381 : node370;
									assign node370 = (inp[1]) ? node372 : 3'b110;
										assign node372 = (inp[5]) ? node378 : node373;
											assign node373 = (inp[8]) ? 3'b110 : node374;
												assign node374 = (inp[0]) ? 3'b110 : 3'b010;
											assign node378 = (inp[8]) ? 3'b000 : 3'b110;
									assign node381 = (inp[5]) ? node383 : 3'b010;
										assign node383 = (inp[8]) ? node385 : 3'b110;
											assign node385 = (inp[0]) ? node387 : 3'b000;
												assign node387 = (inp[1]) ? 3'b100 : 3'b000;
								assign node390 = (inp[8]) ? 3'b000 : node391;
									assign node391 = (inp[0]) ? node393 : 3'b100;
										assign node393 = (inp[2]) ? node395 : 3'b100;
											assign node395 = (inp[5]) ? 3'b000 : 3'b100;
							assign node399 = (inp[7]) ? node431 : node400;
								assign node400 = (inp[8]) ? node418 : node401;
									assign node401 = (inp[1]) ? node407 : node402;
										assign node402 = (inp[2]) ? node404 : 3'b001;
											assign node404 = (inp[0]) ? 3'b001 : 3'b011;
										assign node407 = (inp[5]) ? node413 : node408;
											assign node408 = (inp[0]) ? node410 : 3'b111;
												assign node410 = (inp[2]) ? 3'b001 : 3'b011;
											assign node413 = (inp[0]) ? node415 : 3'b011;
												assign node415 = (inp[2]) ? 3'b110 : 3'b100;
									assign node418 = (inp[5]) ? node424 : node419;
										assign node419 = (inp[1]) ? 3'b110 : node420;
											assign node420 = (inp[2]) ? 3'b101 : 3'b001;
										assign node424 = (inp[2]) ? node426 : 3'b110;
											assign node426 = (inp[0]) ? node428 : 3'b110;
												assign node428 = (inp[1]) ? 3'b010 : 3'b110;
								assign node431 = (inp[2]) ? node439 : node432;
									assign node432 = (inp[0]) ? 3'b010 : node433;
										assign node433 = (inp[8]) ? 3'b010 : node434;
											assign node434 = (inp[5]) ? 3'b010 : 3'b110;
									assign node439 = (inp[8]) ? node449 : node440;
										assign node440 = (inp[1]) ? node446 : node441;
											assign node441 = (inp[5]) ? 3'b010 : node442;
												assign node442 = (inp[0]) ? 3'b010 : 3'b110;
											assign node446 = (inp[5]) ? 3'b100 : 3'b010;
										assign node449 = (inp[5]) ? 3'b100 : node450;
											assign node450 = (inp[1]) ? node452 : 3'b110;
												assign node452 = (inp[0]) ? 3'b100 : 3'b110;
						assign node456 = (inp[7]) ? 3'b000 : node457;
							assign node457 = (inp[11]) ? node469 : node458;
								assign node458 = (inp[8]) ? 3'b000 : node459;
									assign node459 = (inp[0]) ? node461 : 3'b100;
										assign node461 = (inp[5]) ? node463 : 3'b100;
											assign node463 = (inp[2]) ? 3'b000 : node464;
												assign node464 = (inp[1]) ? 3'b000 : 3'b100;
								assign node469 = (inp[5]) ? node477 : node470;
									assign node470 = (inp[0]) ? 3'b010 : node471;
										assign node471 = (inp[8]) ? node473 : 3'b110;
											assign node473 = (inp[2]) ? 3'b110 : 3'b010;
									assign node477 = (inp[8]) ? 3'b100 : node478;
										assign node478 = (inp[0]) ? node480 : 3'b010;
											assign node480 = (inp[1]) ? 3'b100 : 3'b010;
				assign node485 = (inp[4]) ? node585 : node486;
					assign node486 = (inp[7]) ? node516 : node487;
						assign node487 = (inp[10]) ? 3'b011 : node488;
							assign node488 = (inp[5]) ? node508 : node489;
								assign node489 = (inp[8]) ? node497 : node490;
									assign node490 = (inp[0]) ? node492 : 3'b001;
										assign node492 = (inp[2]) ? node494 : 3'b001;
											assign node494 = (inp[11]) ? 3'b011 : 3'b001;
									assign node497 = (inp[11]) ? node503 : node498;
										assign node498 = (inp[1]) ? node500 : 3'b001;
											assign node500 = (inp[0]) ? 3'b011 : 3'b001;
										assign node503 = (inp[1]) ? node505 : 3'b011;
											assign node505 = (inp[0]) ? 3'b001 : 3'b011;
								assign node508 = (inp[11]) ? node510 : 3'b011;
									assign node510 = (inp[2]) ? 3'b001 : node511;
										assign node511 = (inp[8]) ? 3'b001 : 3'b011;
						assign node516 = (inp[10]) ? node566 : node517;
							assign node517 = (inp[11]) ? node533 : node518;
								assign node518 = (inp[5]) ? node526 : node519;
									assign node519 = (inp[0]) ? node521 : 3'b010;
										assign node521 = (inp[2]) ? node523 : 3'b110;
											assign node523 = (inp[8]) ? 3'b010 : 3'b110;
									assign node526 = (inp[8]) ? node530 : node527;
										assign node527 = (inp[1]) ? 3'b010 : 3'b110;
										assign node530 = (inp[1]) ? 3'b100 : 3'b000;
								assign node533 = (inp[5]) ? node549 : node534;
									assign node534 = (inp[2]) ? node540 : node535;
										assign node535 = (inp[8]) ? 3'b001 : node536;
											assign node536 = (inp[0]) ? 3'b011 : 3'b111;
										assign node540 = (inp[1]) ? node544 : node541;
											assign node541 = (inp[8]) ? 3'b101 : 3'b001;
											assign node544 = (inp[0]) ? 3'b110 : node545;
												assign node545 = (inp[8]) ? 3'b101 : 3'b111;
									assign node549 = (inp[8]) ? node561 : node550;
										assign node550 = (inp[2]) ? node556 : node551;
											assign node551 = (inp[0]) ? node553 : 3'b001;
												assign node553 = (inp[1]) ? 3'b100 : 3'b001;
											assign node556 = (inp[1]) ? node558 : 3'b011;
												assign node558 = (inp[0]) ? 3'b110 : 3'b011;
										assign node561 = (inp[0]) ? node563 : 3'b110;
											assign node563 = (inp[1]) ? 3'b010 : 3'b110;
							assign node566 = (inp[5]) ? node576 : node567;
								assign node567 = (inp[11]) ? node569 : 3'b001;
									assign node569 = (inp[1]) ? node571 : 3'b011;
										assign node571 = (inp[8]) ? node573 : 3'b011;
											assign node573 = (inp[0]) ? 3'b101 : 3'b111;
								assign node576 = (inp[11]) ? node580 : node577;
									assign node577 = (inp[8]) ? 3'b110 : 3'b111;
									assign node580 = (inp[8]) ? node582 : 3'b101;
										assign node582 = (inp[1]) ? 3'b001 : 3'b101;
					assign node585 = (inp[10]) ? node633 : node586;
						assign node586 = (inp[11]) ? node602 : node587;
							assign node587 = (inp[8]) ? node593 : node588;
								assign node588 = (inp[7]) ? node590 : 3'b010;
									assign node590 = (inp[5]) ? 3'b000 : 3'b010;
								assign node593 = (inp[7]) ? node595 : 3'b100;
									assign node595 = (inp[5]) ? 3'b000 : node596;
										assign node596 = (inp[0]) ? node598 : 3'b010;
											assign node598 = (inp[1]) ? 3'b000 : 3'b010;
							assign node602 = (inp[7]) ? node618 : node603;
								assign node603 = (inp[0]) ? node613 : node604;
									assign node604 = (inp[2]) ? node608 : node605;
										assign node605 = (inp[8]) ? 3'b101 : 3'b001;
										assign node608 = (inp[8]) ? node610 : 3'b110;
											assign node610 = (inp[1]) ? 3'b010 : 3'b110;
									assign node613 = (inp[8]) ? node615 : 3'b110;
										assign node615 = (inp[1]) ? 3'b010 : 3'b110;
								assign node618 = (inp[5]) ? node626 : node619;
									assign node619 = (inp[8]) ? node621 : 3'b010;
										assign node621 = (inp[0]) ? node623 : 3'b110;
											assign node623 = (inp[1]) ? 3'b100 : 3'b110;
									assign node626 = (inp[8]) ? node630 : node627;
										assign node627 = (inp[0]) ? 3'b100 : 3'b000;
										assign node630 = (inp[0]) ? 3'b000 : 3'b100;
						assign node633 = (inp[7]) ? node671 : node634;
							assign node634 = (inp[8]) ? node654 : node635;
								assign node635 = (inp[11]) ? node649 : node636;
									assign node636 = (inp[5]) ? node638 : 3'b101;
										assign node638 = (inp[1]) ? node644 : node639;
											assign node639 = (inp[2]) ? 3'b101 : node640;
												assign node640 = (inp[0]) ? 3'b001 : 3'b101;
											assign node644 = (inp[2]) ? 3'b001 : node645;
												assign node645 = (inp[0]) ? 3'b001 : 3'b101;
									assign node649 = (inp[0]) ? node651 : 3'b011;
										assign node651 = (inp[5]) ? 3'b101 : 3'b011;
								assign node654 = (inp[11]) ? node668 : node655;
									assign node655 = (inp[1]) ? node663 : node656;
										assign node656 = (inp[5]) ? node658 : 3'b001;
											assign node658 = (inp[0]) ? node660 : 3'b001;
												assign node660 = (inp[2]) ? 3'b001 : 3'b110;
										assign node663 = (inp[5]) ? 3'b110 : node664;
											assign node664 = (inp[2]) ? 3'b110 : 3'b001;
									assign node668 = (inp[5]) ? 3'b001 : 3'b101;
							assign node671 = (inp[11]) ? node691 : node672;
								assign node672 = (inp[8]) ? node678 : node673;
									assign node673 = (inp[2]) ? node675 : 3'b110;
										assign node675 = (inp[0]) ? 3'b010 : 3'b110;
									assign node678 = (inp[1]) ? node684 : node679;
										assign node679 = (inp[5]) ? 3'b010 : node680;
											assign node680 = (inp[0]) ? 3'b010 : 3'b110;
										assign node684 = (inp[5]) ? node688 : node685;
											assign node685 = (inp[0]) ? 3'b010 : 3'b110;
											assign node688 = (inp[0]) ? 3'b100 : 3'b010;
								assign node691 = (inp[5]) ? node693 : 3'b001;
									assign node693 = (inp[8]) ? node699 : node694;
										assign node694 = (inp[0]) ? node696 : 3'b101;
											assign node696 = (inp[1]) ? 3'b110 : 3'b101;
										assign node699 = (inp[1]) ? node701 : 3'b110;
											assign node701 = (inp[2]) ? node703 : 3'b110;
												assign node703 = (inp[0]) ? 3'b010 : 3'b110;
		assign node706 = (inp[9]) ? node832 : node707;
			assign node707 = (inp[6]) ? 3'b000 : node708;
				assign node708 = (inp[4]) ? node820 : node709;
					assign node709 = (inp[7]) ? node785 : node710;
						assign node710 = (inp[11]) ? node736 : node711;
							assign node711 = (inp[8]) ? node729 : node712;
								assign node712 = (inp[10]) ? node718 : node713;
									assign node713 = (inp[5]) ? node715 : 3'b100;
										assign node715 = (inp[0]) ? 3'b000 : 3'b100;
									assign node718 = (inp[2]) ? node724 : node719;
										assign node719 = (inp[5]) ? node721 : 3'b010;
											assign node721 = (inp[0]) ? 3'b010 : 3'b110;
										assign node724 = (inp[0]) ? 3'b110 : node725;
											assign node725 = (inp[5]) ? 3'b110 : 3'b010;
								assign node729 = (inp[10]) ? node731 : 3'b000;
									assign node731 = (inp[5]) ? 3'b000 : node732;
										assign node732 = (inp[2]) ? 3'b010 : 3'b110;
							assign node736 = (inp[10]) ? node760 : node737;
								assign node737 = (inp[5]) ? node749 : node738;
									assign node738 = (inp[0]) ? node744 : node739;
										assign node739 = (inp[8]) ? node741 : 3'b110;
											assign node741 = (inp[2]) ? 3'b110 : 3'b010;
										assign node744 = (inp[2]) ? node746 : 3'b010;
											assign node746 = (inp[1]) ? 3'b010 : 3'b110;
									assign node749 = (inp[8]) ? node755 : node750;
										assign node750 = (inp[0]) ? node752 : 3'b010;
											assign node752 = (inp[1]) ? 3'b100 : 3'b010;
										assign node755 = (inp[2]) ? node757 : 3'b100;
											assign node757 = (inp[1]) ? 3'b000 : 3'b100;
								assign node760 = (inp[5]) ? node772 : node761;
									assign node761 = (inp[2]) ? node765 : node762;
										assign node762 = (inp[8]) ? 3'b001 : 3'b011;
										assign node765 = (inp[8]) ? node769 : node766;
											assign node766 = (inp[0]) ? 3'b001 : 3'b111;
											assign node769 = (inp[1]) ? 3'b110 : 3'b101;
									assign node772 = (inp[8]) ? node780 : node773;
										assign node773 = (inp[0]) ? node775 : 3'b001;
											assign node775 = (inp[1]) ? node777 : 3'b011;
												assign node777 = (inp[2]) ? 3'b110 : 3'b100;
										assign node780 = (inp[0]) ? node782 : 3'b110;
											assign node782 = (inp[2]) ? 3'b010 : 3'b110;
						assign node785 = (inp[10]) ? node787 : 3'b000;
							assign node787 = (inp[11]) ? node799 : node788;
								assign node788 = (inp[8]) ? node794 : node789;
									assign node789 = (inp[0]) ? node791 : 3'b100;
										assign node791 = (inp[5]) ? 3'b000 : 3'b100;
									assign node794 = (inp[0]) ? node796 : 3'b000;
										assign node796 = (inp[5]) ? 3'b100 : 3'b000;
								assign node799 = (inp[8]) ? node811 : node800;
									assign node800 = (inp[5]) ? node806 : node801;
										assign node801 = (inp[1]) ? 3'b010 : node802;
											assign node802 = (inp[2]) ? 3'b010 : 3'b000;
										assign node806 = (inp[1]) ? node808 : 3'b010;
											assign node808 = (inp[2]) ? 3'b100 : 3'b110;
									assign node811 = (inp[0]) ? node815 : node812;
										assign node812 = (inp[5]) ? 3'b100 : 3'b000;
										assign node815 = (inp[1]) ? node817 : 3'b100;
											assign node817 = (inp[5]) ? 3'b000 : 3'b100;
					assign node820 = (inp[10]) ? node822 : 3'b000;
						assign node822 = (inp[11]) ? node824 : 3'b000;
							assign node824 = (inp[7]) ? 3'b000 : node825;
								assign node825 = (inp[5]) ? node827 : 3'b100;
									assign node827 = (inp[8]) ? 3'b000 : 3'b100;
			assign node832 = (inp[6]) ? node1070 : node833;
				assign node833 = (inp[4]) ? node951 : node834;
					assign node834 = (inp[7]) ? node860 : node835;
						assign node835 = (inp[10]) ? 3'b111 : node836;
							assign node836 = (inp[5]) ? node852 : node837;
								assign node837 = (inp[8]) ? node845 : node838;
									assign node838 = (inp[0]) ? node840 : 3'b101;
										assign node840 = (inp[2]) ? node842 : 3'b101;
											assign node842 = (inp[11]) ? 3'b011 : 3'b101;
									assign node845 = (inp[11]) ? 3'b011 : node846;
										assign node846 = (inp[0]) ? node848 : 3'b101;
											assign node848 = (inp[1]) ? 3'b011 : 3'b101;
								assign node852 = (inp[11]) ? node854 : 3'b011;
									assign node854 = (inp[2]) ? 3'b101 : node855;
										assign node855 = (inp[8]) ? 3'b101 : 3'b011;
						assign node860 = (inp[10]) ? node908 : node861;
							assign node861 = (inp[11]) ? node881 : node862;
								assign node862 = (inp[8]) ? node876 : node863;
									assign node863 = (inp[1]) ? node867 : node864;
										assign node864 = (inp[0]) ? 3'b110 : 3'b010;
										assign node867 = (inp[2]) ? 3'b010 : node868;
											assign node868 = (inp[5]) ? node872 : node869;
												assign node869 = (inp[0]) ? 3'b110 : 3'b010;
												assign node872 = (inp[0]) ? 3'b010 : 3'b110;
									assign node876 = (inp[5]) ? 3'b000 : node877;
										assign node877 = (inp[2]) ? 3'b010 : 3'b110;
								assign node881 = (inp[5]) ? node891 : node882;
									assign node882 = (inp[8]) ? node888 : node883;
										assign node883 = (inp[0]) ? node885 : 3'b111;
											assign node885 = (inp[2]) ? 3'b001 : 3'b011;
										assign node888 = (inp[2]) ? 3'b101 : 3'b001;
									assign node891 = (inp[8]) ? node901 : node892;
										assign node892 = (inp[0]) ? node896 : node893;
											assign node893 = (inp[2]) ? 3'b011 : 3'b001;
											assign node896 = (inp[1]) ? node898 : 3'b011;
												assign node898 = (inp[2]) ? 3'b110 : 3'b100;
										assign node901 = (inp[0]) ? node903 : 3'b110;
											assign node903 = (inp[1]) ? node905 : 3'b110;
												assign node905 = (inp[2]) ? 3'b010 : 3'b110;
							assign node908 = (inp[11]) ? node924 : node909;
								assign node909 = (inp[8]) ? node919 : node910;
									assign node910 = (inp[5]) ? node914 : node911;
										assign node911 = (inp[0]) ? 3'b101 : 3'b001;
										assign node914 = (inp[0]) ? node916 : 3'b101;
											assign node916 = (inp[2]) ? 3'b101 : 3'b001;
									assign node919 = (inp[5]) ? 3'b010 : node920;
										assign node920 = (inp[2]) ? 3'b001 : 3'b101;
								assign node924 = (inp[2]) ? node936 : node925;
									assign node925 = (inp[0]) ? node933 : node926;
										assign node926 = (inp[5]) ? node930 : node927;
											assign node927 = (inp[1]) ? 3'b101 : 3'b011;
											assign node930 = (inp[8]) ? 3'b101 : 3'b011;
										assign node933 = (inp[5]) ? 3'b111 : 3'b011;
									assign node936 = (inp[5]) ? node946 : node937;
										assign node937 = (inp[8]) ? node941 : node938;
											assign node938 = (inp[0]) ? 3'b011 : 3'b101;
											assign node941 = (inp[1]) ? node943 : 3'b111;
												assign node943 = (inp[0]) ? 3'b101 : 3'b111;
										assign node946 = (inp[0]) ? 3'b101 : node947;
											assign node947 = (inp[8]) ? 3'b101 : 3'b001;
					assign node951 = (inp[10]) ? node1001 : node952;
						assign node952 = (inp[7]) ? node968 : node953;
							assign node953 = (inp[8]) ? node963 : node954;
								assign node954 = (inp[11]) ? node956 : 3'b010;
									assign node956 = (inp[2]) ? 3'b110 : node957;
										assign node957 = (inp[0]) ? 3'b110 : node958;
											assign node958 = (inp[1]) ? 3'b110 : 3'b001;
								assign node963 = (inp[11]) ? node965 : 3'b100;
									assign node965 = (inp[1]) ? 3'b010 : 3'b110;
							assign node968 = (inp[5]) ? node984 : node969;
								assign node969 = (inp[1]) ? node975 : node970;
									assign node970 = (inp[2]) ? 3'b100 : node971;
										assign node971 = (inp[8]) ? 3'b000 : 3'b100;
									assign node975 = (inp[8]) ? node979 : node976;
										assign node976 = (inp[11]) ? 3'b010 : 3'b100;
										assign node979 = (inp[11]) ? 3'b100 : node980;
											assign node980 = (inp[0]) ? 3'b000 : 3'b100;
								assign node984 = (inp[11]) ? node986 : 3'b000;
									assign node986 = (inp[8]) ? node994 : node987;
										assign node987 = (inp[1]) ? node991 : node988;
											assign node988 = (inp[2]) ? 3'b010 : 3'b100;
											assign node991 = (inp[2]) ? 3'b100 : 3'b010;
										assign node994 = (inp[1]) ? node998 : node995;
											assign node995 = (inp[2]) ? 3'b100 : 3'b000;
											assign node998 = (inp[2]) ? 3'b000 : 3'b100;
						assign node1001 = (inp[7]) ? node1037 : node1002;
							assign node1002 = (inp[8]) ? node1022 : node1003;
								assign node1003 = (inp[11]) ? node1017 : node1004;
									assign node1004 = (inp[5]) ? node1006 : 3'b101;
										assign node1006 = (inp[0]) ? node1012 : node1007;
											assign node1007 = (inp[2]) ? node1009 : 3'b101;
												assign node1009 = (inp[1]) ? 3'b001 : 3'b101;
											assign node1012 = (inp[1]) ? 3'b001 : node1013;
												assign node1013 = (inp[2]) ? 3'b101 : 3'b001;
									assign node1017 = (inp[0]) ? node1019 : 3'b011;
										assign node1019 = (inp[5]) ? 3'b101 : 3'b011;
								assign node1022 = (inp[11]) ? node1032 : node1023;
									assign node1023 = (inp[5]) ? node1025 : 3'b001;
										assign node1025 = (inp[0]) ? 3'b110 : node1026;
											assign node1026 = (inp[2]) ? node1028 : 3'b001;
												assign node1028 = (inp[1]) ? 3'b110 : 3'b001;
									assign node1032 = (inp[0]) ? node1034 : 3'b101;
										assign node1034 = (inp[5]) ? 3'b001 : 3'b101;
							assign node1037 = (inp[11]) ? node1051 : node1038;
								assign node1038 = (inp[8]) ? node1044 : node1039;
									assign node1039 = (inp[0]) ? node1041 : 3'b110;
										assign node1041 = (inp[5]) ? 3'b010 : 3'b110;
									assign node1044 = (inp[1]) ? 3'b100 : node1045;
										assign node1045 = (inp[5]) ? node1047 : 3'b010;
											assign node1047 = (inp[0]) ? 3'b100 : 3'b010;
								assign node1051 = (inp[5]) ? node1059 : node1052;
									assign node1052 = (inp[8]) ? node1054 : 3'b001;
										assign node1054 = (inp[2]) ? 3'b110 : node1055;
											assign node1055 = (inp[0]) ? 3'b101 : 3'b001;
									assign node1059 = (inp[0]) ? node1063 : node1060;
										assign node1060 = (inp[8]) ? 3'b110 : 3'b001;
										assign node1063 = (inp[8]) ? 3'b010 : node1064;
											assign node1064 = (inp[2]) ? 3'b110 : node1065;
												assign node1065 = (inp[1]) ? 3'b110 : 3'b001;
				assign node1070 = (inp[10]) ? node1100 : node1071;
					assign node1071 = (inp[4]) ? 3'b000 : node1072;
						assign node1072 = (inp[7]) ? 3'b000 : node1073;
							assign node1073 = (inp[11]) ? node1081 : node1074;
								assign node1074 = (inp[8]) ? 3'b000 : node1075;
									assign node1075 = (inp[5]) ? node1077 : 3'b100;
										assign node1077 = (inp[0]) ? 3'b000 : 3'b100;
								assign node1081 = (inp[5]) ? node1089 : node1082;
									assign node1082 = (inp[2]) ? node1084 : 3'b010;
										assign node1084 = (inp[0]) ? node1086 : 3'b110;
											assign node1086 = (inp[8]) ? 3'b110 : 3'b010;
									assign node1089 = (inp[8]) ? node1093 : node1090;
										assign node1090 = (inp[0]) ? 3'b100 : 3'b010;
										assign node1093 = (inp[0]) ? node1095 : 3'b100;
											assign node1095 = (inp[1]) ? 3'b000 : 3'b100;
					assign node1100 = (inp[4]) ? node1176 : node1101;
						assign node1101 = (inp[7]) ? node1153 : node1102;
							assign node1102 = (inp[11]) ? node1124 : node1103;
								assign node1103 = (inp[8]) ? node1113 : node1104;
									assign node1104 = (inp[5]) ? node1108 : node1105;
										assign node1105 = (inp[0]) ? 3'b110 : 3'b010;
										assign node1108 = (inp[0]) ? node1110 : 3'b110;
											assign node1110 = (inp[1]) ? 3'b010 : 3'b110;
									assign node1113 = (inp[5]) ? node1117 : node1114;
										assign node1114 = (inp[2]) ? 3'b010 : 3'b110;
										assign node1117 = (inp[2]) ? node1119 : 3'b000;
											assign node1119 = (inp[1]) ? node1121 : 3'b000;
												assign node1121 = (inp[0]) ? 3'b100 : 3'b000;
								assign node1124 = (inp[8]) ? node1140 : node1125;
									assign node1125 = (inp[1]) ? node1131 : node1126;
										assign node1126 = (inp[2]) ? node1128 : 3'b001;
											assign node1128 = (inp[5]) ? 3'b011 : 3'b001;
										assign node1131 = (inp[5]) ? node1135 : node1132;
											assign node1132 = (inp[0]) ? 3'b011 : 3'b111;
											assign node1135 = (inp[0]) ? 3'b100 : node1136;
												assign node1136 = (inp[2]) ? 3'b011 : 3'b001;
									assign node1140 = (inp[5]) ? node1148 : node1141;
										assign node1141 = (inp[2]) ? node1143 : 3'b001;
											assign node1143 = (inp[0]) ? node1145 : 3'b101;
												assign node1145 = (inp[1]) ? 3'b110 : 3'b101;
										assign node1148 = (inp[1]) ? node1150 : 3'b110;
											assign node1150 = (inp[2]) ? 3'b010 : 3'b110;
							assign node1153 = (inp[11]) ? node1161 : node1154;
								assign node1154 = (inp[5]) ? 3'b000 : node1155;
									assign node1155 = (inp[1]) ? node1157 : 3'b100;
										assign node1157 = (inp[0]) ? 3'b000 : 3'b100;
								assign node1161 = (inp[5]) ? node1169 : node1162;
									assign node1162 = (inp[8]) ? 3'b010 : node1163;
										assign node1163 = (inp[0]) ? node1165 : 3'b110;
											assign node1165 = (inp[2]) ? 3'b010 : 3'b110;
									assign node1169 = (inp[8]) ? 3'b100 : node1170;
										assign node1170 = (inp[1]) ? 3'b100 : node1171;
											assign node1171 = (inp[2]) ? 3'b110 : 3'b010;
						assign node1176 = (inp[7]) ? node1214 : node1177;
							assign node1177 = (inp[11]) ? node1189 : node1178;
								assign node1178 = (inp[8]) ? 3'b000 : node1179;
									assign node1179 = (inp[5]) ? node1181 : 3'b100;
										assign node1181 = (inp[0]) ? node1183 : 3'b100;
											assign node1183 = (inp[2]) ? 3'b000 : node1184;
												assign node1184 = (inp[1]) ? 3'b000 : 3'b100;
								assign node1189 = (inp[8]) ? node1203 : node1190;
									assign node1190 = (inp[2]) ? 3'b010 : node1191;
										assign node1191 = (inp[1]) ? node1197 : node1192;
											assign node1192 = (inp[0]) ? 3'b010 : node1193;
												assign node1193 = (inp[5]) ? 3'b010 : 3'b110;
											assign node1197 = (inp[0]) ? node1199 : 3'b010;
												assign node1199 = (inp[5]) ? 3'b100 : 3'b010;
									assign node1203 = (inp[5]) ? node1209 : node1204;
										assign node1204 = (inp[2]) ? node1206 : 3'b010;
											assign node1206 = (inp[1]) ? 3'b100 : 3'b110;
										assign node1209 = (inp[0]) ? node1211 : 3'b100;
											assign node1211 = (inp[1]) ? 3'b000 : 3'b100;
							assign node1214 = (inp[8]) ? 3'b000 : node1215;
								assign node1215 = (inp[5]) ? 3'b000 : node1216;
									assign node1216 = (inp[2]) ? 3'b000 : node1217;
										assign node1217 = (inp[11]) ? 3'b100 : 3'b000;

endmodule