module dtc_split25_bm80 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node7;
	wire [3-1:0] node8;
	wire [3-1:0] node12;
	wire [3-1:0] node14;
	wire [3-1:0] node17;
	wire [3-1:0] node18;
	wire [3-1:0] node19;
	wire [3-1:0] node22;
	wire [3-1:0] node24;
	wire [3-1:0] node27;
	wire [3-1:0] node28;
	wire [3-1:0] node30;
	wire [3-1:0] node33;
	wire [3-1:0] node34;
	wire [3-1:0] node37;
	wire [3-1:0] node40;
	wire [3-1:0] node41;
	wire [3-1:0] node42;
	wire [3-1:0] node43;
	wire [3-1:0] node45;
	wire [3-1:0] node46;
	wire [3-1:0] node51;
	wire [3-1:0] node52;
	wire [3-1:0] node55;
	wire [3-1:0] node56;
	wire [3-1:0] node60;
	wire [3-1:0] node61;
	wire [3-1:0] node62;
	wire [3-1:0] node63;
	wire [3-1:0] node64;
	wire [3-1:0] node69;
	wire [3-1:0] node72;
	wire [3-1:0] node73;
	wire [3-1:0] node74;
	wire [3-1:0] node78;
	wire [3-1:0] node80;
	wire [3-1:0] node83;
	wire [3-1:0] node84;
	wire [3-1:0] node85;
	wire [3-1:0] node86;
	wire [3-1:0] node87;
	wire [3-1:0] node88;
	wire [3-1:0] node93;
	wire [3-1:0] node95;
	wire [3-1:0] node96;
	wire [3-1:0] node100;
	wire [3-1:0] node101;
	wire [3-1:0] node102;
	wire [3-1:0] node103;
	wire [3-1:0] node106;
	wire [3-1:0] node109;
	wire [3-1:0] node112;
	wire [3-1:0] node113;
	wire [3-1:0] node114;
	wire [3-1:0] node117;
	wire [3-1:0] node120;
	wire [3-1:0] node121;
	wire [3-1:0] node125;
	wire [3-1:0] node126;
	wire [3-1:0] node127;
	wire [3-1:0] node128;
	wire [3-1:0] node129;
	wire [3-1:0] node131;
	wire [3-1:0] node135;
	wire [3-1:0] node138;
	wire [3-1:0] node139;
	wire [3-1:0] node142;
	wire [3-1:0] node144;
	wire [3-1:0] node147;
	wire [3-1:0] node148;
	wire [3-1:0] node149;
	wire [3-1:0] node153;
	wire [3-1:0] node154;
	wire [3-1:0] node155;
	wire [3-1:0] node158;
	wire [3-1:0] node159;
	wire [3-1:0] node163;
	wire [3-1:0] node165;
	wire [3-1:0] node167;
	wire [3-1:0] node168;
	wire [3-1:0] node172;
	wire [3-1:0] node173;
	wire [3-1:0] node174;
	wire [3-1:0] node175;
	wire [3-1:0] node176;
	wire [3-1:0] node177;
	wire [3-1:0] node179;
	wire [3-1:0] node181;
	wire [3-1:0] node185;
	wire [3-1:0] node188;
	wire [3-1:0] node189;
	wire [3-1:0] node190;
	wire [3-1:0] node191;
	wire [3-1:0] node193;
	wire [3-1:0] node196;
	wire [3-1:0] node197;
	wire [3-1:0] node201;
	wire [3-1:0] node202;
	wire [3-1:0] node205;
	wire [3-1:0] node208;
	wire [3-1:0] node209;
	wire [3-1:0] node210;
	wire [3-1:0] node211;
	wire [3-1:0] node213;
	wire [3-1:0] node218;
	wire [3-1:0] node220;
	wire [3-1:0] node223;
	wire [3-1:0] node224;
	wire [3-1:0] node225;
	wire [3-1:0] node226;
	wire [3-1:0] node229;
	wire [3-1:0] node231;
	wire [3-1:0] node232;
	wire [3-1:0] node235;
	wire [3-1:0] node238;
	wire [3-1:0] node239;
	wire [3-1:0] node240;
	wire [3-1:0] node244;
	wire [3-1:0] node245;
	wire [3-1:0] node248;
	wire [3-1:0] node251;
	wire [3-1:0] node252;
	wire [3-1:0] node254;
	wire [3-1:0] node255;
	wire [3-1:0] node259;
	wire [3-1:0] node260;
	wire [3-1:0] node262;
	wire [3-1:0] node265;
	wire [3-1:0] node267;
	wire [3-1:0] node270;
	wire [3-1:0] node271;
	wire [3-1:0] node272;
	wire [3-1:0] node273;
	wire [3-1:0] node275;
	wire [3-1:0] node276;
	wire [3-1:0] node280;
	wire [3-1:0] node281;
	wire [3-1:0] node282;
	wire [3-1:0] node283;
	wire [3-1:0] node285;
	wire [3-1:0] node289;
	wire [3-1:0] node291;
	wire [3-1:0] node293;
	wire [3-1:0] node297;
	wire [3-1:0] node298;
	wire [3-1:0] node299;
	wire [3-1:0] node300;
	wire [3-1:0] node302;
	wire [3-1:0] node306;
	wire [3-1:0] node307;
	wire [3-1:0] node309;
	wire [3-1:0] node311;
	wire [3-1:0] node315;
	wire [3-1:0] node316;
	wire [3-1:0] node318;
	wire [3-1:0] node319;
	wire [3-1:0] node322;
	wire [3-1:0] node325;
	wire [3-1:0] node328;
	wire [3-1:0] node330;
	wire [3-1:0] node331;
	wire [3-1:0] node334;
	wire [3-1:0] node335;
	wire [3-1:0] node339;
	wire [3-1:0] node340;
	wire [3-1:0] node341;
	wire [3-1:0] node342;
	wire [3-1:0] node343;
	wire [3-1:0] node344;
	wire [3-1:0] node345;
	wire [3-1:0] node347;
	wire [3-1:0] node349;
	wire [3-1:0] node352;
	wire [3-1:0] node355;
	wire [3-1:0] node356;
	wire [3-1:0] node358;
	wire [3-1:0] node362;
	wire [3-1:0] node364;
	wire [3-1:0] node365;
	wire [3-1:0] node370;
	wire [3-1:0] node371;
	wire [3-1:0] node372;
	wire [3-1:0] node373;
	wire [3-1:0] node374;
	wire [3-1:0] node377;
	wire [3-1:0] node379;
	wire [3-1:0] node381;
	wire [3-1:0] node384;
	wire [3-1:0] node385;
	wire [3-1:0] node386;
	wire [3-1:0] node388;
	wire [3-1:0] node392;
	wire [3-1:0] node393;
	wire [3-1:0] node396;
	wire [3-1:0] node398;
	wire [3-1:0] node399;
	wire [3-1:0] node403;
	wire [3-1:0] node404;
	wire [3-1:0] node406;
	wire [3-1:0] node409;
	wire [3-1:0] node410;
	wire [3-1:0] node414;
	wire [3-1:0] node415;
	wire [3-1:0] node416;
	wire [3-1:0] node417;
	wire [3-1:0] node421;
	wire [3-1:0] node422;
	wire [3-1:0] node423;
	wire [3-1:0] node424;
	wire [3-1:0] node429;
	wire [3-1:0] node431;
	wire [3-1:0] node435;
	wire [3-1:0] node437;
	wire [3-1:0] node438;
	wire [3-1:0] node439;
	wire [3-1:0] node440;
	wire [3-1:0] node441;
	wire [3-1:0] node442;
	wire [3-1:0] node444;
	wire [3-1:0] node449;
	wire [3-1:0] node450;
	wire [3-1:0] node454;
	wire [3-1:0] node455;
	wire [3-1:0] node456;
	wire [3-1:0] node462;
	wire [3-1:0] node463;
	wire [3-1:0] node464;
	wire [3-1:0] node465;
	wire [3-1:0] node466;
	wire [3-1:0] node468;
	wire [3-1:0] node470;
	wire [3-1:0] node471;
	wire [3-1:0] node472;
	wire [3-1:0] node477;
	wire [3-1:0] node478;
	wire [3-1:0] node479;
	wire [3-1:0] node480;
	wire [3-1:0] node482;
	wire [3-1:0] node483;
	wire [3-1:0] node486;
	wire [3-1:0] node489;
	wire [3-1:0] node490;
	wire [3-1:0] node494;
	wire [3-1:0] node495;
	wire [3-1:0] node497;
	wire [3-1:0] node500;
	wire [3-1:0] node501;
	wire [3-1:0] node503;
	wire [3-1:0] node507;
	wire [3-1:0] node509;
	wire [3-1:0] node511;
	wire [3-1:0] node514;
	wire [3-1:0] node515;
	wire [3-1:0] node516;
	wire [3-1:0] node517;
	wire [3-1:0] node518;
	wire [3-1:0] node520;
	wire [3-1:0] node522;
	wire [3-1:0] node526;
	wire [3-1:0] node527;
	wire [3-1:0] node530;
	wire [3-1:0] node532;
	wire [3-1:0] node535;
	wire [3-1:0] node536;
	wire [3-1:0] node538;
	wire [3-1:0] node541;
	wire [3-1:0] node542;
	wire [3-1:0] node543;
	wire [3-1:0] node546;
	wire [3-1:0] node550;
	wire [3-1:0] node551;
	wire [3-1:0] node552;
	wire [3-1:0] node553;
	wire [3-1:0] node556;
	wire [3-1:0] node558;
	wire [3-1:0] node561;
	wire [3-1:0] node562;
	wire [3-1:0] node563;
	wire [3-1:0] node564;
	wire [3-1:0] node567;
	wire [3-1:0] node571;
	wire [3-1:0] node573;
	wire [3-1:0] node574;
	wire [3-1:0] node578;
	wire [3-1:0] node579;
	wire [3-1:0] node580;
	wire [3-1:0] node582;
	wire [3-1:0] node583;
	wire [3-1:0] node585;
	wire [3-1:0] node589;
	wire [3-1:0] node591;
	wire [3-1:0] node594;
	wire [3-1:0] node595;
	wire [3-1:0] node597;
	wire [3-1:0] node600;
	wire [3-1:0] node603;
	wire [3-1:0] node604;
	wire [3-1:0] node605;
	wire [3-1:0] node606;
	wire [3-1:0] node607;
	wire [3-1:0] node608;
	wire [3-1:0] node612;
	wire [3-1:0] node613;
	wire [3-1:0] node614;
	wire [3-1:0] node618;
	wire [3-1:0] node619;
	wire [3-1:0] node622;
	wire [3-1:0] node624;
	wire [3-1:0] node627;
	wire [3-1:0] node629;
	wire [3-1:0] node630;
	wire [3-1:0] node633;
	wire [3-1:0] node634;
	wire [3-1:0] node638;
	wire [3-1:0] node639;
	wire [3-1:0] node640;
	wire [3-1:0] node641;
	wire [3-1:0] node645;
	wire [3-1:0] node646;
	wire [3-1:0] node648;
	wire [3-1:0] node650;
	wire [3-1:0] node654;
	wire [3-1:0] node655;
	wire [3-1:0] node656;
	wire [3-1:0] node657;
	wire [3-1:0] node660;
	wire [3-1:0] node661;
	wire [3-1:0] node665;
	wire [3-1:0] node666;
	wire [3-1:0] node667;
	wire [3-1:0] node669;
	wire [3-1:0] node673;
	wire [3-1:0] node676;
	wire [3-1:0] node677;
	wire [3-1:0] node679;
	wire [3-1:0] node682;
	wire [3-1:0] node683;
	wire [3-1:0] node687;
	wire [3-1:0] node688;
	wire [3-1:0] node689;
	wire [3-1:0] node690;
	wire [3-1:0] node691;
	wire [3-1:0] node692;
	wire [3-1:0] node693;
	wire [3-1:0] node698;
	wire [3-1:0] node702;
	wire [3-1:0] node703;
	wire [3-1:0] node704;
	wire [3-1:0] node706;
	wire [3-1:0] node708;
	wire [3-1:0] node711;
	wire [3-1:0] node713;
	wire [3-1:0] node716;
	wire [3-1:0] node717;
	wire [3-1:0] node718;
	wire [3-1:0] node721;
	wire [3-1:0] node725;
	wire [3-1:0] node726;
	wire [3-1:0] node727;
	wire [3-1:0] node728;
	wire [3-1:0] node729;
	wire [3-1:0] node731;
	wire [3-1:0] node732;
	wire [3-1:0] node736;
	wire [3-1:0] node737;
	wire [3-1:0] node742;
	wire [3-1:0] node743;
	wire [3-1:0] node744;
	wire [3-1:0] node747;
	wire [3-1:0] node750;
	wire [3-1:0] node752;
	wire [3-1:0] node755;
	wire [3-1:0] node756;
	wire [3-1:0] node757;
	wire [3-1:0] node758;
	wire [3-1:0] node761;
	wire [3-1:0] node764;
	wire [3-1:0] node767;
	wire [3-1:0] node768;
	wire [3-1:0] node772;
	wire [3-1:0] node773;
	wire [3-1:0] node774;
	wire [3-1:0] node775;
	wire [3-1:0] node776;
	wire [3-1:0] node777;
	wire [3-1:0] node778;
	wire [3-1:0] node779;
	wire [3-1:0] node782;
	wire [3-1:0] node785;
	wire [3-1:0] node786;
	wire [3-1:0] node787;
	wire [3-1:0] node792;
	wire [3-1:0] node793;
	wire [3-1:0] node794;
	wire [3-1:0] node798;
	wire [3-1:0] node800;
	wire [3-1:0] node802;
	wire [3-1:0] node805;
	wire [3-1:0] node806;
	wire [3-1:0] node808;
	wire [3-1:0] node809;
	wire [3-1:0] node813;
	wire [3-1:0] node815;
	wire [3-1:0] node817;
	wire [3-1:0] node820;
	wire [3-1:0] node821;
	wire [3-1:0] node822;
	wire [3-1:0] node823;
	wire [3-1:0] node826;
	wire [3-1:0] node827;
	wire [3-1:0] node830;
	wire [3-1:0] node833;
	wire [3-1:0] node834;
	wire [3-1:0] node836;
	wire [3-1:0] node839;
	wire [3-1:0] node840;
	wire [3-1:0] node842;
	wire [3-1:0] node844;
	wire [3-1:0] node848;
	wire [3-1:0] node849;
	wire [3-1:0] node850;
	wire [3-1:0] node852;
	wire [3-1:0] node855;
	wire [3-1:0] node858;
	wire [3-1:0] node859;
	wire [3-1:0] node860;
	wire [3-1:0] node865;
	wire [3-1:0] node866;
	wire [3-1:0] node867;
	wire [3-1:0] node868;
	wire [3-1:0] node869;
	wire [3-1:0] node872;
	wire [3-1:0] node874;
	wire [3-1:0] node877;
	wire [3-1:0] node879;
	wire [3-1:0] node882;
	wire [3-1:0] node883;
	wire [3-1:0] node885;
	wire [3-1:0] node887;
	wire [3-1:0] node889;
	wire [3-1:0] node890;
	wire [3-1:0] node894;
	wire [3-1:0] node895;
	wire [3-1:0] node896;
	wire [3-1:0] node897;
	wire [3-1:0] node901;
	wire [3-1:0] node904;
	wire [3-1:0] node905;
	wire [3-1:0] node906;
	wire [3-1:0] node911;
	wire [3-1:0] node912;
	wire [3-1:0] node913;
	wire [3-1:0] node914;
	wire [3-1:0] node916;
	wire [3-1:0] node919;
	wire [3-1:0] node922;
	wire [3-1:0] node923;
	wire [3-1:0] node924;
	wire [3-1:0] node928;
	wire [3-1:0] node931;
	wire [3-1:0] node932;
	wire [3-1:0] node933;
	wire [3-1:0] node936;
	wire [3-1:0] node939;
	wire [3-1:0] node942;
	wire [3-1:0] node943;
	wire [3-1:0] node944;
	wire [3-1:0] node945;
	wire [3-1:0] node946;
	wire [3-1:0] node947;
	wire [3-1:0] node948;
	wire [3-1:0] node950;
	wire [3-1:0] node954;
	wire [3-1:0] node956;
	wire [3-1:0] node959;
	wire [3-1:0] node961;
	wire [3-1:0] node962;
	wire [3-1:0] node966;
	wire [3-1:0] node967;
	wire [3-1:0] node969;
	wire [3-1:0] node972;
	wire [3-1:0] node974;
	wire [3-1:0] node976;
	wire [3-1:0] node977;
	wire [3-1:0] node978;
	wire [3-1:0] node981;
	wire [3-1:0] node985;
	wire [3-1:0] node986;
	wire [3-1:0] node987;
	wire [3-1:0] node990;
	wire [3-1:0] node991;
	wire [3-1:0] node992;
	wire [3-1:0] node994;
	wire [3-1:0] node997;
	wire [3-1:0] node1000;
	wire [3-1:0] node1001;
	wire [3-1:0] node1004;
	wire [3-1:0] node1007;
	wire [3-1:0] node1008;
	wire [3-1:0] node1009;
	wire [3-1:0] node1010;
	wire [3-1:0] node1014;
	wire [3-1:0] node1016;
	wire [3-1:0] node1019;
	wire [3-1:0] node1020;
	wire [3-1:0] node1023;
	wire [3-1:0] node1026;
	wire [3-1:0] node1027;
	wire [3-1:0] node1028;
	wire [3-1:0] node1029;
	wire [3-1:0] node1030;
	wire [3-1:0] node1033;
	wire [3-1:0] node1037;
	wire [3-1:0] node1038;
	wire [3-1:0] node1039;
	wire [3-1:0] node1040;
	wire [3-1:0] node1045;
	wire [3-1:0] node1046;
	wire [3-1:0] node1047;
	wire [3-1:0] node1050;
	wire [3-1:0] node1054;
	wire [3-1:0] node1055;
	wire [3-1:0] node1057;
	wire [3-1:0] node1058;
	wire [3-1:0] node1061;
	wire [3-1:0] node1062;
	wire [3-1:0] node1063;

	assign outp = (inp[6]) ? node462 : node1;
		assign node1 = (inp[3]) ? node339 : node2;
			assign node2 = (inp[9]) ? node172 : node3;
				assign node3 = (inp[10]) ? node83 : node4;
					assign node4 = (inp[7]) ? node40 : node5;
						assign node5 = (inp[4]) ? node17 : node6;
							assign node6 = (inp[0]) ? node12 : node7;
								assign node7 = (inp[1]) ? 3'b001 : node8;
									assign node8 = (inp[2]) ? 3'b101 : 3'b111;
								assign node12 = (inp[8]) ? node14 : 3'b110;
									assign node14 = (inp[11]) ? 3'b010 : 3'b001;
							assign node17 = (inp[5]) ? node27 : node18;
								assign node18 = (inp[1]) ? node22 : node19;
									assign node19 = (inp[0]) ? 3'b110 : 3'b100;
									assign node22 = (inp[8]) ? node24 : 3'b100;
										assign node24 = (inp[11]) ? 3'b000 : 3'b001;
								assign node27 = (inp[0]) ? node33 : node28;
									assign node28 = (inp[1]) ? node30 : 3'b000;
										assign node30 = (inp[8]) ? 3'b110 : 3'b010;
									assign node33 = (inp[8]) ? node37 : node34;
										assign node34 = (inp[11]) ? 3'b000 : 3'b100;
										assign node37 = (inp[1]) ? 3'b100 : 3'b010;
						assign node40 = (inp[0]) ? node60 : node41;
							assign node41 = (inp[8]) ? node51 : node42;
								assign node42 = (inp[2]) ? 3'b101 : node43;
									assign node43 = (inp[5]) ? node45 : 3'b001;
										assign node45 = (inp[11]) ? 3'b001 : node46;
											assign node46 = (inp[1]) ? 3'b101 : 3'b111;
								assign node51 = (inp[11]) ? node55 : node52;
									assign node52 = (inp[4]) ? 3'b011 : 3'b001;
									assign node55 = (inp[5]) ? 3'b001 : node56;
										assign node56 = (inp[4]) ? 3'b101 : 3'b011;
							assign node60 = (inp[1]) ? node72 : node61;
								assign node61 = (inp[4]) ? node69 : node62;
									assign node62 = (inp[11]) ? 3'b101 : node63;
										assign node63 = (inp[5]) ? 3'b101 : node64;
											assign node64 = (inp[8]) ? 3'b011 : 3'b101;
									assign node69 = (inp[8]) ? 3'b001 : 3'b010;
								assign node72 = (inp[2]) ? node78 : node73;
									assign node73 = (inp[8]) ? 3'b110 : node74;
										assign node74 = (inp[4]) ? 3'b010 : 3'b110;
									assign node78 = (inp[4]) ? node80 : 3'b001;
										assign node80 = (inp[5]) ? 3'b100 : 3'b010;
					assign node83 = (inp[0]) ? node125 : node84;
						assign node84 = (inp[4]) ? node100 : node85;
							assign node85 = (inp[7]) ? node93 : node86;
								assign node86 = (inp[11]) ? 3'b001 : node87;
									assign node87 = (inp[5]) ? 3'b101 : node88;
										assign node88 = (inp[8]) ? 3'b001 : 3'b101;
								assign node93 = (inp[11]) ? node95 : 3'b011;
									assign node95 = (inp[8]) ? 3'b001 : node96;
										assign node96 = (inp[1]) ? 3'b001 : 3'b000;
							assign node100 = (inp[1]) ? node112 : node101;
								assign node101 = (inp[7]) ? node109 : node102;
									assign node102 = (inp[11]) ? node106 : node103;
										assign node103 = (inp[2]) ? 3'b000 : 3'b100;
										assign node106 = (inp[8]) ? 3'b110 : 3'b010;
									assign node109 = (inp[2]) ? 3'b101 : 3'b001;
								assign node112 = (inp[11]) ? node120 : node113;
									assign node113 = (inp[8]) ? node117 : node114;
										assign node114 = (inp[7]) ? 3'b110 : 3'b010;
										assign node117 = (inp[7]) ? 3'b001 : 3'b110;
									assign node120 = (inp[7]) ? 3'b110 : node121;
										assign node121 = (inp[8]) ? 3'b110 : 3'b100;
						assign node125 = (inp[4]) ? node147 : node126;
							assign node126 = (inp[2]) ? node138 : node127;
								assign node127 = (inp[8]) ? node135 : node128;
									assign node128 = (inp[11]) ? 3'b110 : node129;
										assign node129 = (inp[1]) ? node131 : 3'b010;
											assign node131 = (inp[5]) ? 3'b100 : 3'b010;
									assign node135 = (inp[5]) ? 3'b110 : 3'b101;
								assign node138 = (inp[11]) ? node142 : node139;
									assign node139 = (inp[5]) ? 3'b010 : 3'b110;
									assign node142 = (inp[7]) ? node144 : 3'b010;
										assign node144 = (inp[1]) ? 3'b010 : 3'b110;
							assign node147 = (inp[7]) ? node153 : node148;
								assign node148 = (inp[5]) ? 3'b000 : node149;
									assign node149 = (inp[2]) ? 3'b100 : 3'b000;
								assign node153 = (inp[2]) ? node163 : node154;
									assign node154 = (inp[5]) ? node158 : node155;
										assign node155 = (inp[11]) ? 3'b010 : 3'b110;
										assign node158 = (inp[1]) ? 3'b100 : node159;
											assign node159 = (inp[8]) ? 3'b010 : 3'b000;
									assign node163 = (inp[5]) ? node165 : 3'b010;
										assign node165 = (inp[8]) ? node167 : 3'b010;
											assign node167 = (inp[1]) ? 3'b010 : node168;
												assign node168 = (inp[11]) ? 3'b010 : 3'b110;
				assign node172 = (inp[10]) ? node270 : node173;
					assign node173 = (inp[11]) ? node223 : node174;
						assign node174 = (inp[7]) ? node188 : node175;
							assign node175 = (inp[0]) ? node185 : node176;
								assign node176 = (inp[4]) ? 3'b010 : node177;
									assign node177 = (inp[1]) ? node179 : 3'b010;
										assign node179 = (inp[8]) ? node181 : 3'b010;
											assign node181 = (inp[2]) ? 3'b110 : 3'b111;
								assign node185 = (inp[4]) ? 3'b000 : 3'b010;
							assign node188 = (inp[4]) ? node208 : node189;
								assign node189 = (inp[0]) ? node201 : node190;
									assign node190 = (inp[2]) ? node196 : node191;
										assign node191 = (inp[8]) ? node193 : 3'b110;
											assign node193 = (inp[1]) ? 3'b001 : 3'b000;
										assign node196 = (inp[8]) ? 3'b101 : node197;
											assign node197 = (inp[5]) ? 3'b000 : 3'b101;
									assign node201 = (inp[8]) ? node205 : node202;
										assign node202 = (inp[2]) ? 3'b110 : 3'b100;
										assign node205 = (inp[5]) ? 3'b010 : 3'b110;
								assign node208 = (inp[0]) ? node218 : node209;
									assign node209 = (inp[8]) ? 3'b110 : node210;
										assign node210 = (inp[2]) ? 3'b010 : node211;
											assign node211 = (inp[1]) ? node213 : 3'b010;
												assign node213 = (inp[5]) ? 3'b010 : 3'b011;
									assign node218 = (inp[1]) ? node220 : 3'b010;
										assign node220 = (inp[2]) ? 3'b000 : 3'b100;
						assign node223 = (inp[0]) ? node251 : node224;
							assign node224 = (inp[1]) ? node238 : node225;
								assign node225 = (inp[4]) ? node229 : node226;
									assign node226 = (inp[5]) ? 3'b000 : 3'b100;
									assign node229 = (inp[7]) ? node231 : 3'b010;
										assign node231 = (inp[5]) ? node235 : node232;
											assign node232 = (inp[2]) ? 3'b010 : 3'b000;
											assign node235 = (inp[8]) ? 3'b100 : 3'b000;
								assign node238 = (inp[4]) ? node244 : node239;
									assign node239 = (inp[7]) ? 3'b101 : node240;
										assign node240 = (inp[2]) ? 3'b100 : 3'b110;
									assign node244 = (inp[7]) ? node248 : node245;
										assign node245 = (inp[5]) ? 3'b100 : 3'b000;
										assign node248 = (inp[2]) ? 3'b110 : 3'b010;
							assign node251 = (inp[7]) ? node259 : node252;
								assign node252 = (inp[5]) ? node254 : 3'b000;
									assign node254 = (inp[4]) ? 3'b000 : node255;
										assign node255 = (inp[8]) ? 3'b000 : 3'b100;
								assign node259 = (inp[8]) ? node265 : node260;
									assign node260 = (inp[5]) ? node262 : 3'b100;
										assign node262 = (inp[1]) ? 3'b100 : 3'b010;
									assign node265 = (inp[5]) ? node267 : 3'b000;
										assign node267 = (inp[4]) ? 3'b000 : 3'b010;
					assign node270 = (inp[4]) ? node328 : node271;
						assign node271 = (inp[7]) ? node297 : node272;
							assign node272 = (inp[2]) ? node280 : node273;
								assign node273 = (inp[1]) ? node275 : 3'b100;
									assign node275 = (inp[5]) ? 3'b100 : node276;
										assign node276 = (inp[0]) ? 3'b000 : 3'b010;
								assign node280 = (inp[0]) ? 3'b000 : node281;
									assign node281 = (inp[11]) ? node289 : node282;
										assign node282 = (inp[1]) ? 3'b010 : node283;
											assign node283 = (inp[8]) ? node285 : 3'b000;
												assign node285 = (inp[5]) ? 3'b100 : 3'b000;
										assign node289 = (inp[1]) ? node291 : 3'b000;
											assign node291 = (inp[5]) ? node293 : 3'b100;
												assign node293 = (inp[8]) ? 3'b100 : 3'b000;
							assign node297 = (inp[11]) ? node315 : node298;
								assign node298 = (inp[1]) ? node306 : node299;
									assign node299 = (inp[8]) ? 3'b110 : node300;
										assign node300 = (inp[2]) ? node302 : 3'b000;
											assign node302 = (inp[5]) ? 3'b100 : 3'b000;
									assign node306 = (inp[2]) ? 3'b110 : node307;
										assign node307 = (inp[5]) ? node309 : 3'b001;
											assign node309 = (inp[8]) ? node311 : 3'b101;
												assign node311 = (inp[0]) ? 3'b100 : 3'b110;
								assign node315 = (inp[8]) ? node325 : node316;
									assign node316 = (inp[0]) ? node318 : 3'b010;
										assign node318 = (inp[5]) ? node322 : node319;
											assign node319 = (inp[1]) ? 3'b100 : 3'b010;
											assign node322 = (inp[1]) ? 3'b000 : 3'b100;
									assign node325 = (inp[0]) ? 3'b010 : 3'b001;
						assign node328 = (inp[7]) ? node330 : 3'b000;
							assign node330 = (inp[11]) ? node334 : node331;
								assign node331 = (inp[8]) ? 3'b100 : 3'b000;
								assign node334 = (inp[0]) ? 3'b000 : node335;
									assign node335 = (inp[1]) ? 3'b010 : 3'b000;
			assign node339 = (inp[4]) ? node435 : node340;
				assign node340 = (inp[7]) ? node370 : node341;
					assign node341 = (inp[9]) ? 3'b000 : node342;
						assign node342 = (inp[5]) ? node362 : node343;
							assign node343 = (inp[11]) ? node355 : node344;
								assign node344 = (inp[10]) ? node352 : node345;
									assign node345 = (inp[1]) ? node347 : 3'b100;
										assign node347 = (inp[0]) ? node349 : 3'b010;
											assign node349 = (inp[8]) ? 3'b100 : 3'b000;
									assign node352 = (inp[1]) ? 3'b100 : 3'b000;
								assign node355 = (inp[10]) ? 3'b000 : node356;
									assign node356 = (inp[2]) ? node358 : 3'b000;
										assign node358 = (inp[0]) ? 3'b000 : 3'b010;
							assign node362 = (inp[1]) ? node364 : 3'b000;
								assign node364 = (inp[0]) ? 3'b000 : node365;
									assign node365 = (inp[8]) ? 3'b100 : 3'b000;
					assign node370 = (inp[0]) ? node414 : node371;
						assign node371 = (inp[9]) ? node403 : node372;
							assign node372 = (inp[10]) ? node384 : node373;
								assign node373 = (inp[11]) ? node377 : node374;
									assign node374 = (inp[1]) ? 3'b010 : 3'b000;
									assign node377 = (inp[2]) ? node379 : 3'b110;
										assign node379 = (inp[8]) ? node381 : 3'b010;
											assign node381 = (inp[5]) ? 3'b010 : 3'b000;
								assign node384 = (inp[8]) ? node392 : node385;
									assign node385 = (inp[1]) ? 3'b100 : node386;
										assign node386 = (inp[5]) ? node388 : 3'b110;
											assign node388 = (inp[11]) ? 3'b010 : 3'b000;
									assign node392 = (inp[1]) ? node396 : node393;
										assign node393 = (inp[5]) ? 3'b110 : 3'b000;
										assign node396 = (inp[2]) ? node398 : 3'b010;
											assign node398 = (inp[5]) ? 3'b010 : node399;
												assign node399 = (inp[11]) ? 3'b010 : 3'b110;
							assign node403 = (inp[1]) ? node409 : node404;
								assign node404 = (inp[5]) ? node406 : 3'b010;
									assign node406 = (inp[10]) ? 3'b000 : 3'b010;
								assign node409 = (inp[5]) ? 3'b000 : node410;
									assign node410 = (inp[10]) ? 3'b000 : 3'b100;
						assign node414 = (inp[9]) ? 3'b000 : node415;
							assign node415 = (inp[5]) ? node421 : node416;
								assign node416 = (inp[2]) ? 3'b010 : node417;
									assign node417 = (inp[8]) ? 3'b100 : 3'b110;
								assign node421 = (inp[8]) ? node429 : node422;
									assign node422 = (inp[11]) ? 3'b000 : node423;
										assign node423 = (inp[1]) ? 3'b000 : node424;
											assign node424 = (inp[10]) ? 3'b000 : 3'b100;
									assign node429 = (inp[10]) ? node431 : 3'b100;
										assign node431 = (inp[2]) ? 3'b000 : 3'b100;
				assign node435 = (inp[7]) ? node437 : 3'b000;
					assign node437 = (inp[9]) ? 3'b000 : node438;
						assign node438 = (inp[11]) ? node454 : node439;
							assign node439 = (inp[0]) ? node449 : node440;
								assign node440 = (inp[10]) ? 3'b100 : node441;
									assign node441 = (inp[8]) ? 3'b010 : node442;
										assign node442 = (inp[2]) ? node444 : 3'b100;
											assign node444 = (inp[1]) ? 3'b010 : 3'b100;
								assign node449 = (inp[5]) ? 3'b000 : node450;
									assign node450 = (inp[1]) ? 3'b000 : 3'b100;
							assign node454 = (inp[5]) ? 3'b000 : node455;
								assign node455 = (inp[0]) ? 3'b000 : node456;
									assign node456 = (inp[2]) ? 3'b100 : 3'b000;
		assign node462 = (inp[3]) ? node772 : node463;
			assign node463 = (inp[9]) ? node603 : node464;
				assign node464 = (inp[0]) ? node514 : node465;
					assign node465 = (inp[1]) ? node477 : node466;
						assign node466 = (inp[4]) ? node468 : 3'b111;
							assign node468 = (inp[10]) ? node470 : 3'b111;
								assign node470 = (inp[7]) ? 3'b111 : node471;
									assign node471 = (inp[11]) ? 3'b011 : node472;
										assign node472 = (inp[5]) ? 3'b011 : 3'b111;
						assign node477 = (inp[7]) ? node507 : node478;
							assign node478 = (inp[11]) ? node494 : node479;
								assign node479 = (inp[4]) ? node489 : node480;
									assign node480 = (inp[10]) ? node482 : 3'b111;
										assign node482 = (inp[2]) ? node486 : node483;
											assign node483 = (inp[5]) ? 3'b111 : 3'b011;
											assign node486 = (inp[5]) ? 3'b011 : 3'b111;
									assign node489 = (inp[5]) ? 3'b011 : node490;
										assign node490 = (inp[8]) ? 3'b111 : 3'b011;
								assign node494 = (inp[4]) ? node500 : node495;
									assign node495 = (inp[8]) ? node497 : 3'b011;
										assign node497 = (inp[10]) ? 3'b011 : 3'b111;
									assign node500 = (inp[2]) ? 3'b101 : node501;
										assign node501 = (inp[8]) ? node503 : 3'b101;
											assign node503 = (inp[10]) ? 3'b101 : 3'b011;
							assign node507 = (inp[4]) ? node509 : 3'b111;
								assign node509 = (inp[2]) ? node511 : 3'b011;
									assign node511 = (inp[8]) ? 3'b111 : 3'b011;
					assign node514 = (inp[4]) ? node550 : node515;
						assign node515 = (inp[7]) ? node535 : node516;
							assign node516 = (inp[5]) ? node526 : node517;
								assign node517 = (inp[10]) ? 3'b101 : node518;
									assign node518 = (inp[1]) ? node520 : 3'b111;
										assign node520 = (inp[11]) ? node522 : 3'b011;
											assign node522 = (inp[8]) ? 3'b011 : 3'b101;
								assign node526 = (inp[11]) ? node530 : node527;
									assign node527 = (inp[1]) ? 3'b101 : 3'b011;
									assign node530 = (inp[2]) ? node532 : 3'b001;
										assign node532 = (inp[10]) ? 3'b001 : 3'b101;
							assign node535 = (inp[1]) ? node541 : node536;
								assign node536 = (inp[11]) ? node538 : 3'b111;
									assign node538 = (inp[10]) ? 3'b011 : 3'b111;
								assign node541 = (inp[2]) ? 3'b111 : node542;
									assign node542 = (inp[10]) ? node546 : node543;
										assign node543 = (inp[5]) ? 3'b111 : 3'b011;
										assign node546 = (inp[5]) ? 3'b001 : 3'b011;
						assign node550 = (inp[10]) ? node578 : node551;
							assign node551 = (inp[1]) ? node561 : node552;
								assign node552 = (inp[7]) ? node556 : node553;
									assign node553 = (inp[8]) ? 3'b101 : 3'b001;
									assign node556 = (inp[8]) ? node558 : 3'b011;
										assign node558 = (inp[5]) ? 3'b011 : 3'b111;
								assign node561 = (inp[5]) ? node571 : node562;
									assign node562 = (inp[11]) ? 3'b001 : node563;
										assign node563 = (inp[7]) ? node567 : node564;
											assign node564 = (inp[8]) ? 3'b101 : 3'b001;
											assign node567 = (inp[2]) ? 3'b101 : 3'b001;
									assign node571 = (inp[7]) ? node573 : 3'b110;
										assign node573 = (inp[8]) ? 3'b101 : node574;
											assign node574 = (inp[11]) ? 3'b001 : 3'b101;
							assign node578 = (inp[1]) ? node594 : node579;
								assign node579 = (inp[8]) ? node589 : node580;
									assign node580 = (inp[7]) ? node582 : 3'b110;
										assign node582 = (inp[11]) ? 3'b101 : node583;
											assign node583 = (inp[2]) ? node585 : 3'b111;
												assign node585 = (inp[5]) ? 3'b101 : 3'b111;
									assign node589 = (inp[7]) ? node591 : 3'b001;
										assign node591 = (inp[11]) ? 3'b011 : 3'b111;
								assign node594 = (inp[7]) ? node600 : node595;
									assign node595 = (inp[5]) ? node597 : 3'b110;
										assign node597 = (inp[8]) ? 3'b110 : 3'b010;
									assign node600 = (inp[5]) ? 3'b010 : 3'b001;
				assign node603 = (inp[4]) ? node687 : node604;
					assign node604 = (inp[0]) ? node638 : node605;
						assign node605 = (inp[7]) ? node627 : node606;
							assign node606 = (inp[5]) ? node612 : node607;
								assign node607 = (inp[11]) ? 3'b011 : node608;
									assign node608 = (inp[1]) ? 3'b001 : 3'b011;
								assign node612 = (inp[1]) ? node618 : node613;
									assign node613 = (inp[8]) ? 3'b011 : node614;
										assign node614 = (inp[10]) ? 3'b111 : 3'b101;
									assign node618 = (inp[8]) ? node622 : node619;
										assign node619 = (inp[10]) ? 3'b111 : 3'b001;
										assign node622 = (inp[10]) ? node624 : 3'b101;
											assign node624 = (inp[11]) ? 3'b001 : 3'b101;
							assign node627 = (inp[10]) ? node629 : 3'b111;
								assign node629 = (inp[2]) ? node633 : node630;
									assign node630 = (inp[1]) ? 3'b101 : 3'b111;
									assign node633 = (inp[5]) ? 3'b011 : node634;
										assign node634 = (inp[1]) ? 3'b011 : 3'b111;
						assign node638 = (inp[8]) ? node654 : node639;
							assign node639 = (inp[10]) ? node645 : node640;
								assign node640 = (inp[5]) ? 3'b101 : node641;
									assign node641 = (inp[1]) ? 3'b001 : 3'b011;
								assign node645 = (inp[2]) ? 3'b110 : node646;
									assign node646 = (inp[11]) ? node648 : 3'b110;
										assign node648 = (inp[1]) ? node650 : 3'b101;
											assign node650 = (inp[7]) ? 3'b110 : 3'b000;
							assign node654 = (inp[2]) ? node676 : node655;
								assign node655 = (inp[10]) ? node665 : node656;
									assign node656 = (inp[5]) ? node660 : node657;
										assign node657 = (inp[7]) ? 3'b111 : 3'b101;
										assign node660 = (inp[1]) ? 3'b010 : node661;
											assign node661 = (inp[7]) ? 3'b011 : 3'b101;
									assign node665 = (inp[11]) ? node673 : node666;
										assign node666 = (inp[5]) ? 3'b101 : node667;
											assign node667 = (inp[7]) ? node669 : 3'b101;
												assign node669 = (inp[1]) ? 3'b101 : 3'b011;
										assign node673 = (inp[7]) ? 3'b001 : 3'b010;
								assign node676 = (inp[11]) ? node682 : node677;
									assign node677 = (inp[5]) ? node679 : 3'b101;
										assign node679 = (inp[7]) ? 3'b101 : 3'b001;
									assign node682 = (inp[1]) ? 3'b001 : node683;
										assign node683 = (inp[5]) ? 3'b001 : 3'b101;
					assign node687 = (inp[0]) ? node725 : node688;
						assign node688 = (inp[10]) ? node702 : node689;
							assign node689 = (inp[2]) ? 3'b101 : node690;
								assign node690 = (inp[1]) ? node698 : node691;
									assign node691 = (inp[7]) ? 3'b111 : node692;
										assign node692 = (inp[8]) ? 3'b101 : node693;
											assign node693 = (inp[11]) ? 3'b101 : 3'b001;
									assign node698 = (inp[11]) ? 3'b001 : 3'b011;
							assign node702 = (inp[7]) ? node716 : node703;
								assign node703 = (inp[1]) ? node711 : node704;
									assign node704 = (inp[11]) ? node706 : 3'b110;
										assign node706 = (inp[8]) ? node708 : 3'b000;
											assign node708 = (inp[5]) ? 3'b000 : 3'b001;
									assign node711 = (inp[5]) ? node713 : 3'b110;
										assign node713 = (inp[8]) ? 3'b110 : 3'b101;
								assign node716 = (inp[1]) ? 3'b101 : node717;
									assign node717 = (inp[11]) ? node721 : node718;
										assign node718 = (inp[8]) ? 3'b011 : 3'b111;
										assign node721 = (inp[5]) ? 3'b001 : 3'b101;
						assign node725 = (inp[8]) ? node755 : node726;
							assign node726 = (inp[2]) ? node742 : node727;
								assign node727 = (inp[7]) ? 3'b110 : node728;
									assign node728 = (inp[1]) ? node736 : node729;
										assign node729 = (inp[11]) ? node731 : 3'b010;
											assign node731 = (inp[10]) ? 3'b010 : node732;
												assign node732 = (inp[5]) ? 3'b010 : 3'b101;
										assign node736 = (inp[11]) ? 3'b010 : node737;
											assign node737 = (inp[10]) ? 3'b100 : 3'b110;
								assign node742 = (inp[10]) ? node750 : node743;
									assign node743 = (inp[7]) ? node747 : node744;
										assign node744 = (inp[5]) ? 3'b100 : 3'b010;
										assign node747 = (inp[11]) ? 3'b010 : 3'b001;
									assign node750 = (inp[5]) ? node752 : 3'b110;
										assign node752 = (inp[7]) ? 3'b010 : 3'b000;
							assign node755 = (inp[7]) ? node767 : node756;
								assign node756 = (inp[5]) ? node764 : node757;
									assign node757 = (inp[11]) ? node761 : node758;
										assign node758 = (inp[10]) ? 3'b010 : 3'b001;
										assign node761 = (inp[1]) ? 3'b000 : 3'b110;
									assign node764 = (inp[10]) ? 3'b100 : 3'b110;
								assign node767 = (inp[2]) ? 3'b001 : node768;
									assign node768 = (inp[1]) ? 3'b000 : 3'b101;
			assign node772 = (inp[0]) ? node942 : node773;
				assign node773 = (inp[7]) ? node865 : node774;
					assign node774 = (inp[4]) ? node820 : node775;
						assign node775 = (inp[10]) ? node805 : node776;
							assign node776 = (inp[5]) ? node792 : node777;
								assign node777 = (inp[11]) ? node785 : node778;
									assign node778 = (inp[2]) ? node782 : node779;
										assign node779 = (inp[9]) ? 3'b101 : 3'b011;
										assign node782 = (inp[9]) ? 3'b100 : 3'b101;
									assign node785 = (inp[1]) ? 3'b110 : node786;
										assign node786 = (inp[8]) ? 3'b111 : node787;
											assign node787 = (inp[2]) ? 3'b111 : 3'b101;
								assign node792 = (inp[1]) ? node798 : node793;
									assign node793 = (inp[2]) ? 3'b110 : node794;
										assign node794 = (inp[11]) ? 3'b110 : 3'b100;
									assign node798 = (inp[9]) ? node800 : 3'b001;
										assign node800 = (inp[11]) ? node802 : 3'b010;
											assign node802 = (inp[2]) ? 3'b100 : 3'b010;
							assign node805 = (inp[1]) ? node813 : node806;
								assign node806 = (inp[8]) ? node808 : 3'b010;
									assign node808 = (inp[5]) ? 3'b110 : node809;
										assign node809 = (inp[11]) ? 3'b110 : 3'b100;
								assign node813 = (inp[9]) ? node815 : 3'b110;
									assign node815 = (inp[8]) ? node817 : 3'b100;
										assign node817 = (inp[5]) ? 3'b100 : 3'b010;
						assign node820 = (inp[11]) ? node848 : node821;
							assign node821 = (inp[9]) ? node833 : node822;
								assign node822 = (inp[8]) ? node826 : node823;
									assign node823 = (inp[2]) ? 3'b110 : 3'b010;
									assign node826 = (inp[2]) ? node830 : node827;
										assign node827 = (inp[5]) ? 3'b110 : 3'b100;
										assign node830 = (inp[1]) ? 3'b001 : 3'b000;
								assign node833 = (inp[1]) ? node839 : node834;
									assign node834 = (inp[10]) ? node836 : 3'b110;
										assign node836 = (inp[5]) ? 3'b100 : 3'b110;
									assign node839 = (inp[5]) ? 3'b000 : node840;
										assign node840 = (inp[2]) ? node842 : 3'b100;
											assign node842 = (inp[10]) ? node844 : 3'b100;
												assign node844 = (inp[8]) ? 3'b100 : 3'b000;
							assign node848 = (inp[1]) ? node858 : node849;
								assign node849 = (inp[8]) ? node855 : node850;
									assign node850 = (inp[5]) ? node852 : 3'b010;
										assign node852 = (inp[9]) ? 3'b000 : 3'b010;
									assign node855 = (inp[10]) ? 3'b110 : 3'b000;
								assign node858 = (inp[9]) ? 3'b000 : node859;
									assign node859 = (inp[8]) ? 3'b110 : node860;
										assign node860 = (inp[10]) ? 3'b100 : 3'b000;
					assign node865 = (inp[9]) ? node911 : node866;
						assign node866 = (inp[4]) ? node882 : node867;
							assign node867 = (inp[10]) ? node877 : node868;
								assign node868 = (inp[8]) ? node872 : node869;
									assign node869 = (inp[1]) ? 3'b101 : 3'b011;
									assign node872 = (inp[5]) ? node874 : 3'b111;
										assign node874 = (inp[1]) ? 3'b011 : 3'b111;
								assign node877 = (inp[2]) ? node879 : 3'b011;
									assign node879 = (inp[5]) ? 3'b111 : 3'b011;
							assign node882 = (inp[5]) ? node894 : node883;
								assign node883 = (inp[1]) ? node885 : 3'b101;
									assign node885 = (inp[11]) ? node887 : 3'b001;
										assign node887 = (inp[2]) ? node889 : 3'b101;
											assign node889 = (inp[10]) ? 3'b001 : node890;
												assign node890 = (inp[8]) ? 3'b101 : 3'b001;
								assign node894 = (inp[2]) ? node904 : node895;
									assign node895 = (inp[10]) ? node901 : node896;
										assign node896 = (inp[11]) ? 3'b001 : node897;
											assign node897 = (inp[8]) ? 3'b011 : 3'b111;
										assign node901 = (inp[1]) ? 3'b001 : 3'b101;
									assign node904 = (inp[10]) ? 3'b110 : node905;
										assign node905 = (inp[8]) ? 3'b001 : node906;
											assign node906 = (inp[1]) ? 3'b110 : 3'b001;
						assign node911 = (inp[5]) ? node931 : node912;
							assign node912 = (inp[8]) ? node922 : node913;
								assign node913 = (inp[1]) ? node919 : node914;
									assign node914 = (inp[11]) ? node916 : 3'b001;
										assign node916 = (inp[4]) ? 3'b110 : 3'b101;
									assign node919 = (inp[4]) ? 3'b100 : 3'b110;
								assign node922 = (inp[4]) ? node928 : node923;
									assign node923 = (inp[10]) ? 3'b001 : node924;
										assign node924 = (inp[2]) ? 3'b001 : 3'b101;
									assign node928 = (inp[10]) ? 3'b110 : 3'b001;
							assign node931 = (inp[1]) ? node939 : node932;
								assign node932 = (inp[10]) ? node936 : node933;
									assign node933 = (inp[4]) ? 3'b110 : 3'b001;
									assign node936 = (inp[4]) ? 3'b010 : 3'b110;
								assign node939 = (inp[10]) ? 3'b100 : 3'b010;
				assign node942 = (inp[9]) ? node1026 : node943;
					assign node943 = (inp[7]) ? node985 : node944;
						assign node944 = (inp[2]) ? node966 : node945;
							assign node945 = (inp[8]) ? node959 : node946;
								assign node946 = (inp[4]) ? node954 : node947;
									assign node947 = (inp[5]) ? 3'b010 : node948;
										assign node948 = (inp[10]) ? node950 : 3'b100;
											assign node950 = (inp[11]) ? 3'b010 : 3'b110;
									assign node954 = (inp[1]) ? node956 : 3'b110;
										assign node956 = (inp[5]) ? 3'b100 : 3'b000;
								assign node959 = (inp[5]) ? node961 : 3'b110;
									assign node961 = (inp[11]) ? 3'b100 : node962;
										assign node962 = (inp[1]) ? 3'b010 : 3'b100;
							assign node966 = (inp[1]) ? node972 : node967;
								assign node967 = (inp[8]) ? node969 : 3'b110;
									assign node969 = (inp[4]) ? 3'b010 : 3'b001;
								assign node972 = (inp[5]) ? node974 : 3'b010;
									assign node974 = (inp[10]) ? node976 : 3'b100;
										assign node976 = (inp[4]) ? 3'b000 : node977;
											assign node977 = (inp[11]) ? node981 : node978;
												assign node978 = (inp[8]) ? 3'b010 : 3'b100;
												assign node981 = (inp[8]) ? 3'b100 : 3'b000;
						assign node985 = (inp[4]) ? node1007 : node986;
							assign node986 = (inp[1]) ? node990 : node987;
								assign node987 = (inp[5]) ? 3'b001 : 3'b101;
								assign node990 = (inp[10]) ? node1000 : node991;
									assign node991 = (inp[2]) ? node997 : node992;
										assign node992 = (inp[8]) ? node994 : 3'b001;
											assign node994 = (inp[5]) ? 3'b001 : 3'b101;
										assign node997 = (inp[8]) ? 3'b001 : 3'b110;
									assign node1000 = (inp[11]) ? node1004 : node1001;
										assign node1001 = (inp[8]) ? 3'b001 : 3'b110;
										assign node1004 = (inp[8]) ? 3'b110 : 3'b010;
							assign node1007 = (inp[10]) ? node1019 : node1008;
								assign node1008 = (inp[8]) ? node1014 : node1009;
									assign node1009 = (inp[1]) ? 3'b010 : node1010;
										assign node1010 = (inp[5]) ? 3'b010 : 3'b110;
									assign node1014 = (inp[2]) ? node1016 : 3'b001;
										assign node1016 = (inp[5]) ? 3'b110 : 3'b001;
								assign node1019 = (inp[11]) ? node1023 : node1020;
									assign node1020 = (inp[2]) ? 3'b110 : 3'b010;
									assign node1023 = (inp[5]) ? 3'b100 : 3'b000;
					assign node1026 = (inp[4]) ? node1054 : node1027;
						assign node1027 = (inp[7]) ? node1037 : node1028;
							assign node1028 = (inp[11]) ? 3'b000 : node1029;
								assign node1029 = (inp[1]) ? node1033 : node1030;
									assign node1030 = (inp[5]) ? 3'b110 : 3'b010;
									assign node1033 = (inp[5]) ? 3'b000 : 3'b100;
							assign node1037 = (inp[10]) ? node1045 : node1038;
								assign node1038 = (inp[2]) ? 3'b010 : node1039;
									assign node1039 = (inp[11]) ? 3'b010 : node1040;
										assign node1040 = (inp[5]) ? 3'b010 : 3'b110;
								assign node1045 = (inp[5]) ? 3'b100 : node1046;
									assign node1046 = (inp[8]) ? node1050 : node1047;
										assign node1047 = (inp[2]) ? 3'b100 : 3'b010;
										assign node1050 = (inp[2]) ? 3'b010 : 3'b110;
						assign node1054 = (inp[1]) ? 3'b000 : node1055;
							assign node1055 = (inp[7]) ? node1057 : 3'b000;
								assign node1057 = (inp[8]) ? node1061 : node1058;
									assign node1058 = (inp[11]) ? 3'b000 : 3'b100;
									assign node1061 = (inp[5]) ? 3'b100 : node1062;
										assign node1062 = (inp[10]) ? 3'b100 : node1063;
											assign node1063 = (inp[2]) ? 3'b010 : 3'b110;

endmodule