module dtc_split5_bm68 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node6;
	wire [3-1:0] node8;
	wire [3-1:0] node10;
	wire [3-1:0] node11;
	wire [3-1:0] node15;
	wire [3-1:0] node16;
	wire [3-1:0] node17;
	wire [3-1:0] node19;
	wire [3-1:0] node21;
	wire [3-1:0] node23;
	wire [3-1:0] node24;
	wire [3-1:0] node28;
	wire [3-1:0] node29;
	wire [3-1:0] node31;
	wire [3-1:0] node32;
	wire [3-1:0] node33;
	wire [3-1:0] node35;
	wire [3-1:0] node38;
	wire [3-1:0] node39;
	wire [3-1:0] node45;
	wire [3-1:0] node46;
	wire [3-1:0] node47;
	wire [3-1:0] node48;
	wire [3-1:0] node49;
	wire [3-1:0] node50;
	wire [3-1:0] node52;
	wire [3-1:0] node56;
	wire [3-1:0] node57;
	wire [3-1:0] node59;
	wire [3-1:0] node64;
	wire [3-1:0] node66;
	wire [3-1:0] node67;
	wire [3-1:0] node71;
	wire [3-1:0] node72;
	wire [3-1:0] node74;
	wire [3-1:0] node75;
	wire [3-1:0] node80;
	wire [3-1:0] node81;
	wire [3-1:0] node82;
	wire [3-1:0] node83;
	wire [3-1:0] node85;
	wire [3-1:0] node86;
	wire [3-1:0] node87;
	wire [3-1:0] node92;
	wire [3-1:0] node94;
	wire [3-1:0] node95;
	wire [3-1:0] node96;
	wire [3-1:0] node98;
	wire [3-1:0] node103;
	wire [3-1:0] node104;
	wire [3-1:0] node105;
	wire [3-1:0] node107;
	wire [3-1:0] node109;
	wire [3-1:0] node113;
	wire [3-1:0] node115;
	wire [3-1:0] node116;
	wire [3-1:0] node117;
	wire [3-1:0] node122;
	wire [3-1:0] node123;
	wire [3-1:0] node124;
	wire [3-1:0] node125;
	wire [3-1:0] node126;
	wire [3-1:0] node128;
	wire [3-1:0] node129;
	wire [3-1:0] node134;
	wire [3-1:0] node135;
	wire [3-1:0] node137;
	wire [3-1:0] node139;
	wire [3-1:0] node142;
	wire [3-1:0] node143;
	wire [3-1:0] node145;
	wire [3-1:0] node149;
	wire [3-1:0] node150;
	wire [3-1:0] node152;
	wire [3-1:0] node154;
	wire [3-1:0] node155;
	wire [3-1:0] node160;
	wire [3-1:0] node161;
	wire [3-1:0] node162;
	wire [3-1:0] node163;
	wire [3-1:0] node164;
	wire [3-1:0] node169;
	wire [3-1:0] node172;
	wire [3-1:0] node173;
	wire [3-1:0] node174;
	wire [3-1:0] node176;
	wire [3-1:0] node179;
	wire [3-1:0] node180;
	wire [3-1:0] node184;
	wire [3-1:0] node186;
	wire [3-1:0] node188;
	wire [3-1:0] node191;
	wire [3-1:0] node192;
	wire [3-1:0] node193;
	wire [3-1:0] node194;
	wire [3-1:0] node195;
	wire [3-1:0] node197;
	wire [3-1:0] node198;
	wire [3-1:0] node199;
	wire [3-1:0] node204;
	wire [3-1:0] node205;
	wire [3-1:0] node206;
	wire [3-1:0] node207;
	wire [3-1:0] node208;
	wire [3-1:0] node214;
	wire [3-1:0] node215;
	wire [3-1:0] node217;
	wire [3-1:0] node221;
	wire [3-1:0] node222;
	wire [3-1:0] node225;
	wire [3-1:0] node227;
	wire [3-1:0] node228;
	wire [3-1:0] node230;
	wire [3-1:0] node231;
	wire [3-1:0] node236;
	wire [3-1:0] node237;
	wire [3-1:0] node238;
	wire [3-1:0] node239;
	wire [3-1:0] node240;
	wire [3-1:0] node241;
	wire [3-1:0] node243;
	wire [3-1:0] node246;
	wire [3-1:0] node247;
	wire [3-1:0] node252;
	wire [3-1:0] node254;
	wire [3-1:0] node257;
	wire [3-1:0] node258;
	wire [3-1:0] node261;
	wire [3-1:0] node262;
	wire [3-1:0] node263;
	wire [3-1:0] node267;
	wire [3-1:0] node269;
	wire [3-1:0] node272;
	wire [3-1:0] node273;
	wire [3-1:0] node274;
	wire [3-1:0] node275;
	wire [3-1:0] node279;
	wire [3-1:0] node281;
	wire [3-1:0] node282;
	wire [3-1:0] node286;
	wire [3-1:0] node287;
	wire [3-1:0] node288;
	wire [3-1:0] node290;
	wire [3-1:0] node294;
	wire [3-1:0] node296;
	wire [3-1:0] node298;
	wire [3-1:0] node300;
	wire [3-1:0] node303;
	wire [3-1:0] node304;
	wire [3-1:0] node305;
	wire [3-1:0] node306;
	wire [3-1:0] node307;
	wire [3-1:0] node309;
	wire [3-1:0] node311;
	wire [3-1:0] node315;
	wire [3-1:0] node317;
	wire [3-1:0] node318;
	wire [3-1:0] node322;
	wire [3-1:0] node323;
	wire [3-1:0] node324;
	wire [3-1:0] node326;
	wire [3-1:0] node328;
	wire [3-1:0] node329;
	wire [3-1:0] node334;
	wire [3-1:0] node336;
	wire [3-1:0] node337;
	wire [3-1:0] node338;
	wire [3-1:0] node343;
	wire [3-1:0] node344;
	wire [3-1:0] node345;
	wire [3-1:0] node346;
	wire [3-1:0] node347;
	wire [3-1:0] node351;
	wire [3-1:0] node352;
	wire [3-1:0] node354;
	wire [3-1:0] node358;
	wire [3-1:0] node359;
	wire [3-1:0] node360;
	wire [3-1:0] node362;
	wire [3-1:0] node366;
	wire [3-1:0] node368;
	wire [3-1:0] node370;
	wire [3-1:0] node373;
	wire [3-1:0] node374;
	wire [3-1:0] node375;
	wire [3-1:0] node376;
	wire [3-1:0] node377;
	wire [3-1:0] node379;
	wire [3-1:0] node380;
	wire [3-1:0] node386;
	wire [3-1:0] node387;
	wire [3-1:0] node389;
	wire [3-1:0] node391;
	wire [3-1:0] node395;
	wire [3-1:0] node396;
	wire [3-1:0] node397;
	wire [3-1:0] node398;
	wire [3-1:0] node404;
	wire [3-1:0] node405;
	wire [3-1:0] node406;
	wire [3-1:0] node407;
	wire [3-1:0] node408;
	wire [3-1:0] node409;
	wire [3-1:0] node410;
	wire [3-1:0] node412;
	wire [3-1:0] node414;
	wire [3-1:0] node418;
	wire [3-1:0] node420;
	wire [3-1:0] node421;
	wire [3-1:0] node422;
	wire [3-1:0] node424;
	wire [3-1:0] node429;
	wire [3-1:0] node430;
	wire [3-1:0] node431;
	wire [3-1:0] node433;
	wire [3-1:0] node437;
	wire [3-1:0] node440;
	wire [3-1:0] node441;
	wire [3-1:0] node442;
	wire [3-1:0] node444;
	wire [3-1:0] node445;
	wire [3-1:0] node447;
	wire [3-1:0] node449;
	wire [3-1:0] node452;
	wire [3-1:0] node453;
	wire [3-1:0] node457;
	wire [3-1:0] node458;
	wire [3-1:0] node461;
	wire [3-1:0] node463;
	wire [3-1:0] node464;
	wire [3-1:0] node466;
	wire [3-1:0] node469;
	wire [3-1:0] node470;
	wire [3-1:0] node474;
	wire [3-1:0] node475;
	wire [3-1:0] node476;
	wire [3-1:0] node477;
	wire [3-1:0] node481;
	wire [3-1:0] node482;
	wire [3-1:0] node484;
	wire [3-1:0] node485;
	wire [3-1:0] node490;
	wire [3-1:0] node491;
	wire [3-1:0] node492;
	wire [3-1:0] node494;
	wire [3-1:0] node496;
	wire [3-1:0] node500;
	wire [3-1:0] node502;
	wire [3-1:0] node503;
	wire [3-1:0] node505;
	wire [3-1:0] node509;
	wire [3-1:0] node510;
	wire [3-1:0] node511;
	wire [3-1:0] node512;
	wire [3-1:0] node513;
	wire [3-1:0] node515;
	wire [3-1:0] node516;
	wire [3-1:0] node518;
	wire [3-1:0] node521;
	wire [3-1:0] node522;
	wire [3-1:0] node523;
	wire [3-1:0] node529;
	wire [3-1:0] node530;
	wire [3-1:0] node532;
	wire [3-1:0] node534;
	wire [3-1:0] node538;
	wire [3-1:0] node539;
	wire [3-1:0] node540;
	wire [3-1:0] node542;
	wire [3-1:0] node543;
	wire [3-1:0] node548;
	wire [3-1:0] node549;
	wire [3-1:0] node551;
	wire [3-1:0] node553;
	wire [3-1:0] node555;
	wire [3-1:0] node557;
	wire [3-1:0] node561;
	wire [3-1:0] node562;
	wire [3-1:0] node563;
	wire [3-1:0] node564;
	wire [3-1:0] node565;
	wire [3-1:0] node569;
	wire [3-1:0] node570;
	wire [3-1:0] node574;
	wire [3-1:0] node575;
	wire [3-1:0] node576;
	wire [3-1:0] node577;
	wire [3-1:0] node579;
	wire [3-1:0] node582;
	wire [3-1:0] node583;
	wire [3-1:0] node590;
	wire [3-1:0] node591;
	wire [3-1:0] node592;
	wire [3-1:0] node593;
	wire [3-1:0] node594;
	wire [3-1:0] node595;
	wire [3-1:0] node597;
	wire [3-1:0] node598;
	wire [3-1:0] node600;
	wire [3-1:0] node603;
	wire [3-1:0] node604;
	wire [3-1:0] node609;
	wire [3-1:0] node611;
	wire [3-1:0] node613;
	wire [3-1:0] node614;
	wire [3-1:0] node615;
	wire [3-1:0] node620;
	wire [3-1:0] node621;
	wire [3-1:0] node622;
	wire [3-1:0] node624;
	wire [3-1:0] node625;
	wire [3-1:0] node631;
	wire [3-1:0] node632;
	wire [3-1:0] node633;
	wire [3-1:0] node634;
	wire [3-1:0] node635;

	assign outp = (inp[9]) ? node404 : node1;
		assign node1 = (inp[6]) ? node191 : node2;
			assign node2 = (inp[10]) ? node80 : node3;
				assign node3 = (inp[7]) ? node15 : node4;
					assign node4 = (inp[8]) ? node6 : 3'b111;
						assign node6 = (inp[11]) ? node8 : 3'b111;
							assign node8 = (inp[3]) ? node10 : 3'b111;
								assign node10 = (inp[0]) ? 3'b011 : node11;
									assign node11 = (inp[4]) ? 3'b011 : 3'b111;
					assign node15 = (inp[11]) ? node45 : node16;
						assign node16 = (inp[8]) ? node28 : node17;
							assign node17 = (inp[0]) ? node19 : 3'b111;
								assign node19 = (inp[4]) ? node21 : 3'b111;
									assign node21 = (inp[3]) ? node23 : 3'b111;
										assign node23 = (inp[5]) ? 3'b011 : node24;
											assign node24 = (inp[1]) ? 3'b011 : 3'b111;
							assign node28 = (inp[3]) ? 3'b011 : node29;
								assign node29 = (inp[4]) ? node31 : 3'b111;
									assign node31 = (inp[2]) ? 3'b011 : node32;
										assign node32 = (inp[1]) ? node38 : node33;
											assign node33 = (inp[0]) ? node35 : 3'b111;
												assign node35 = (inp[5]) ? 3'b011 : 3'b111;
											assign node38 = (inp[0]) ? 3'b011 : node39;
												assign node39 = (inp[5]) ? 3'b011 : 3'b111;
						assign node45 = (inp[8]) ? node71 : node46;
							assign node46 = (inp[3]) ? node64 : node47;
								assign node47 = (inp[4]) ? 3'b011 : node48;
									assign node48 = (inp[2]) ? node56 : node49;
										assign node49 = (inp[1]) ? 3'b111 : node50;
											assign node50 = (inp[5]) ? node52 : 3'b111;
												assign node52 = (inp[0]) ? 3'b011 : 3'b111;
										assign node56 = (inp[5]) ? 3'b011 : node57;
											assign node57 = (inp[1]) ? node59 : 3'b111;
												assign node59 = (inp[0]) ? 3'b011 : 3'b111;
								assign node64 = (inp[4]) ? node66 : 3'b011;
									assign node66 = (inp[5]) ? 3'b101 : node67;
										assign node67 = (inp[0]) ? 3'b101 : 3'b011;
							assign node71 = (inp[3]) ? 3'b101 : node72;
								assign node72 = (inp[4]) ? node74 : 3'b011;
									assign node74 = (inp[0]) ? 3'b101 : node75;
										assign node75 = (inp[5]) ? 3'b101 : 3'b011;
				assign node80 = (inp[7]) ? node122 : node81;
					assign node81 = (inp[11]) ? node103 : node82;
						assign node82 = (inp[8]) ? node92 : node83;
							assign node83 = (inp[3]) ? node85 : 3'b111;
								assign node85 = (inp[0]) ? 3'b011 : node86;
									assign node86 = (inp[5]) ? 3'b011 : node87;
										assign node87 = (inp[1]) ? 3'b011 : 3'b111;
							assign node92 = (inp[3]) ? node94 : 3'b011;
								assign node94 = (inp[0]) ? 3'b101 : node95;
									assign node95 = (inp[4]) ? 3'b101 : node96;
										assign node96 = (inp[5]) ? node98 : 3'b011;
											assign node98 = (inp[2]) ? 3'b101 : 3'b011;
						assign node103 = (inp[3]) ? node113 : node104;
							assign node104 = (inp[8]) ? 3'b101 : node105;
								assign node105 = (inp[5]) ? node107 : 3'b011;
									assign node107 = (inp[0]) ? node109 : 3'b011;
										assign node109 = (inp[4]) ? 3'b101 : 3'b011;
							assign node113 = (inp[8]) ? node115 : 3'b101;
								assign node115 = (inp[4]) ? 3'b001 : node116;
									assign node116 = (inp[5]) ? 3'b001 : node117;
										assign node117 = (inp[1]) ? 3'b001 : 3'b101;
					assign node122 = (inp[11]) ? node160 : node123;
						assign node123 = (inp[3]) ? node149 : node124;
							assign node124 = (inp[8]) ? node134 : node125;
								assign node125 = (inp[4]) ? 3'b101 : node126;
									assign node126 = (inp[1]) ? node128 : 3'b011;
										assign node128 = (inp[0]) ? 3'b101 : node129;
											assign node129 = (inp[5]) ? 3'b101 : 3'b011;
								assign node134 = (inp[4]) ? node142 : node135;
									assign node135 = (inp[2]) ? node137 : 3'b101;
										assign node137 = (inp[5]) ? node139 : 3'b101;
											assign node139 = (inp[1]) ? 3'b001 : 3'b101;
									assign node142 = (inp[0]) ? 3'b001 : node143;
										assign node143 = (inp[2]) ? node145 : 3'b001;
											assign node145 = (inp[1]) ? 3'b001 : 3'b101;
							assign node149 = (inp[8]) ? 3'b001 : node150;
								assign node150 = (inp[4]) ? node152 : 3'b101;
									assign node152 = (inp[2]) ? node154 : 3'b001;
										assign node154 = (inp[5]) ? 3'b001 : node155;
											assign node155 = (inp[0]) ? 3'b001 : 3'b101;
						assign node160 = (inp[8]) ? node172 : node161;
							assign node161 = (inp[3]) ? node169 : node162;
								assign node162 = (inp[4]) ? 3'b001 : node163;
									assign node163 = (inp[0]) ? 3'b001 : node164;
										assign node164 = (inp[5]) ? 3'b001 : 3'b101;
								assign node169 = (inp[4]) ? 3'b110 : 3'b001;
							assign node172 = (inp[3]) ? node184 : node173;
								assign node173 = (inp[4]) ? node179 : node174;
									assign node174 = (inp[1]) ? node176 : 3'b001;
										assign node176 = (inp[5]) ? 3'b110 : 3'b001;
									assign node179 = (inp[5]) ? 3'b110 : node180;
										assign node180 = (inp[2]) ? 3'b110 : 3'b001;
								assign node184 = (inp[0]) ? node186 : 3'b110;
									assign node186 = (inp[4]) ? node188 : 3'b110;
										assign node188 = (inp[2]) ? 3'b010 : 3'b110;
			assign node191 = (inp[10]) ? node303 : node192;
				assign node192 = (inp[7]) ? node236 : node193;
					assign node193 = (inp[11]) ? node221 : node194;
						assign node194 = (inp[3]) ? node204 : node195;
							assign node195 = (inp[8]) ? node197 : 3'b011;
								assign node197 = (inp[0]) ? 3'b101 : node198;
									assign node198 = (inp[1]) ? 3'b101 : node199;
										assign node199 = (inp[4]) ? 3'b101 : 3'b011;
							assign node204 = (inp[8]) ? node214 : node205;
								assign node205 = (inp[0]) ? 3'b101 : node206;
									assign node206 = (inp[5]) ? 3'b101 : node207;
										assign node207 = (inp[4]) ? 3'b101 : node208;
											assign node208 = (inp[1]) ? 3'b101 : 3'b011;
								assign node214 = (inp[4]) ? 3'b001 : node215;
									assign node215 = (inp[0]) ? node217 : 3'b101;
										assign node217 = (inp[5]) ? 3'b001 : 3'b101;
						assign node221 = (inp[8]) ? node225 : node222;
							assign node222 = (inp[3]) ? 3'b001 : 3'b101;
							assign node225 = (inp[3]) ? node227 : 3'b001;
								assign node227 = (inp[4]) ? 3'b110 : node228;
									assign node228 = (inp[5]) ? node230 : 3'b001;
										assign node230 = (inp[1]) ? 3'b110 : node231;
											assign node231 = (inp[0]) ? 3'b110 : 3'b001;
					assign node236 = (inp[11]) ? node272 : node237;
						assign node237 = (inp[8]) ? node257 : node238;
							assign node238 = (inp[3]) ? node252 : node239;
								assign node239 = (inp[4]) ? 3'b001 : node240;
									assign node240 = (inp[1]) ? node246 : node241;
										assign node241 = (inp[5]) ? node243 : 3'b101;
											assign node243 = (inp[0]) ? 3'b001 : 3'b101;
										assign node246 = (inp[5]) ? 3'b001 : node247;
											assign node247 = (inp[0]) ? 3'b001 : 3'b101;
								assign node252 = (inp[4]) ? node254 : 3'b001;
									assign node254 = (inp[5]) ? 3'b110 : 3'b001;
							assign node257 = (inp[4]) ? node261 : node258;
								assign node258 = (inp[3]) ? 3'b110 : 3'b001;
								assign node261 = (inp[5]) ? node267 : node262;
									assign node262 = (inp[0]) ? 3'b110 : node263;
										assign node263 = (inp[3]) ? 3'b110 : 3'b001;
									assign node267 = (inp[0]) ? node269 : 3'b110;
										assign node269 = (inp[3]) ? 3'b010 : 3'b110;
						assign node272 = (inp[8]) ? node286 : node273;
							assign node273 = (inp[3]) ? node279 : node274;
								assign node274 = (inp[4]) ? 3'b110 : node275;
									assign node275 = (inp[5]) ? 3'b110 : 3'b001;
								assign node279 = (inp[4]) ? node281 : 3'b110;
									assign node281 = (inp[0]) ? 3'b010 : node282;
										assign node282 = (inp[5]) ? 3'b010 : 3'b110;
							assign node286 = (inp[4]) ? node294 : node287;
								assign node287 = (inp[3]) ? 3'b010 : node288;
									assign node288 = (inp[5]) ? node290 : 3'b110;
										assign node290 = (inp[1]) ? 3'b010 : 3'b110;
								assign node294 = (inp[3]) ? node296 : 3'b010;
									assign node296 = (inp[5]) ? node298 : 3'b010;
										assign node298 = (inp[0]) ? node300 : 3'b010;
											assign node300 = (inp[1]) ? 3'b100 : 3'b010;
				assign node303 = (inp[7]) ? node343 : node304;
					assign node304 = (inp[11]) ? node322 : node305;
						assign node305 = (inp[3]) ? node315 : node306;
							assign node306 = (inp[8]) ? 3'b110 : node307;
								assign node307 = (inp[5]) ? node309 : 3'b001;
									assign node309 = (inp[4]) ? node311 : 3'b001;
										assign node311 = (inp[0]) ? 3'b110 : 3'b001;
							assign node315 = (inp[8]) ? node317 : 3'b110;
								assign node317 = (inp[4]) ? 3'b010 : node318;
									assign node318 = (inp[5]) ? 3'b010 : 3'b110;
						assign node322 = (inp[3]) ? node334 : node323;
							assign node323 = (inp[8]) ? 3'b010 : node324;
								assign node324 = (inp[4]) ? node326 : 3'b110;
									assign node326 = (inp[2]) ? node328 : 3'b110;
										assign node328 = (inp[5]) ? 3'b010 : node329;
											assign node329 = (inp[0]) ? 3'b010 : 3'b110;
							assign node334 = (inp[8]) ? node336 : 3'b010;
								assign node336 = (inp[4]) ? 3'b100 : node337;
									assign node337 = (inp[5]) ? 3'b100 : node338;
										assign node338 = (inp[0]) ? 3'b100 : 3'b010;
					assign node343 = (inp[11]) ? node373 : node344;
						assign node344 = (inp[8]) ? node358 : node345;
							assign node345 = (inp[3]) ? node351 : node346;
								assign node346 = (inp[4]) ? 3'b010 : node347;
									assign node347 = (inp[0]) ? 3'b010 : 3'b110;
								assign node351 = (inp[4]) ? 3'b100 : node352;
									assign node352 = (inp[2]) ? node354 : 3'b010;
										assign node354 = (inp[0]) ? 3'b100 : 3'b010;
							assign node358 = (inp[4]) ? node366 : node359;
								assign node359 = (inp[3]) ? 3'b100 : node360;
									assign node360 = (inp[1]) ? node362 : 3'b010;
										assign node362 = (inp[5]) ? 3'b100 : 3'b010;
								assign node366 = (inp[3]) ? node368 : 3'b100;
									assign node368 = (inp[5]) ? node370 : 3'b100;
										assign node370 = (inp[0]) ? 3'b000 : 3'b100;
						assign node373 = (inp[8]) ? node395 : node374;
							assign node374 = (inp[3]) ? node386 : node375;
								assign node375 = (inp[0]) ? 3'b100 : node376;
									assign node376 = (inp[4]) ? 3'b100 : node377;
										assign node377 = (inp[2]) ? node379 : 3'b010;
											assign node379 = (inp[1]) ? 3'b100 : node380;
												assign node380 = (inp[5]) ? 3'b100 : 3'b010;
								assign node386 = (inp[4]) ? 3'b000 : node387;
									assign node387 = (inp[5]) ? node389 : 3'b100;
										assign node389 = (inp[1]) ? node391 : 3'b100;
											assign node391 = (inp[0]) ? 3'b000 : 3'b100;
							assign node395 = (inp[4]) ? 3'b000 : node396;
								assign node396 = (inp[3]) ? 3'b000 : node397;
									assign node397 = (inp[1]) ? 3'b100 : node398;
										assign node398 = (inp[5]) ? 3'b000 : 3'b100;
		assign node404 = (inp[6]) ? node590 : node405;
			assign node405 = (inp[10]) ? node509 : node406;
				assign node406 = (inp[7]) ? node440 : node407;
					assign node407 = (inp[11]) ? node429 : node408;
						assign node408 = (inp[8]) ? node418 : node409;
							assign node409 = (inp[3]) ? 3'b001 : node410;
								assign node410 = (inp[0]) ? node412 : 3'b101;
									assign node412 = (inp[5]) ? node414 : 3'b101;
										assign node414 = (inp[2]) ? 3'b101 : 3'b001;
							assign node418 = (inp[3]) ? node420 : 3'b001;
								assign node420 = (inp[4]) ? 3'b110 : node421;
									assign node421 = (inp[5]) ? 3'b110 : node422;
										assign node422 = (inp[0]) ? node424 : 3'b001;
											assign node424 = (inp[1]) ? 3'b110 : 3'b001;
						assign node429 = (inp[3]) ? node437 : node430;
							assign node430 = (inp[8]) ? 3'b110 : node431;
								assign node431 = (inp[4]) ? node433 : 3'b001;
									assign node433 = (inp[1]) ? 3'b110 : 3'b001;
							assign node437 = (inp[8]) ? 3'b010 : 3'b110;
					assign node440 = (inp[11]) ? node474 : node441;
						assign node441 = (inp[8]) ? node457 : node442;
							assign node442 = (inp[3]) ? node444 : 3'b110;
								assign node444 = (inp[4]) ? node452 : node445;
									assign node445 = (inp[0]) ? node447 : 3'b110;
										assign node447 = (inp[1]) ? node449 : 3'b110;
											assign node449 = (inp[5]) ? 3'b010 : 3'b110;
									assign node452 = (inp[0]) ? 3'b010 : node453;
										assign node453 = (inp[5]) ? 3'b010 : 3'b110;
							assign node457 = (inp[4]) ? node461 : node458;
								assign node458 = (inp[3]) ? 3'b010 : 3'b110;
								assign node461 = (inp[3]) ? node463 : 3'b010;
									assign node463 = (inp[5]) ? node469 : node464;
										assign node464 = (inp[2]) ? node466 : 3'b010;
											assign node466 = (inp[1]) ? 3'b100 : 3'b010;
										assign node469 = (inp[0]) ? 3'b100 : node470;
											assign node470 = (inp[2]) ? 3'b100 : 3'b010;
						assign node474 = (inp[3]) ? node490 : node475;
							assign node475 = (inp[8]) ? node481 : node476;
								assign node476 = (inp[5]) ? 3'b010 : node477;
									assign node477 = (inp[1]) ? 3'b010 : 3'b110;
								assign node481 = (inp[4]) ? 3'b100 : node482;
									assign node482 = (inp[5]) ? node484 : 3'b010;
										assign node484 = (inp[0]) ? 3'b100 : node485;
											assign node485 = (inp[1]) ? 3'b100 : 3'b010;
							assign node490 = (inp[8]) ? node500 : node491;
								assign node491 = (inp[4]) ? 3'b100 : node492;
									assign node492 = (inp[5]) ? node494 : 3'b010;
										assign node494 = (inp[2]) ? node496 : 3'b010;
											assign node496 = (inp[0]) ? 3'b100 : 3'b010;
								assign node500 = (inp[4]) ? node502 : 3'b100;
									assign node502 = (inp[5]) ? 3'b000 : node503;
										assign node503 = (inp[1]) ? node505 : 3'b100;
											assign node505 = (inp[0]) ? 3'b000 : 3'b100;
				assign node509 = (inp[7]) ? node561 : node510;
					assign node510 = (inp[11]) ? node538 : node511;
						assign node511 = (inp[8]) ? node529 : node512;
							assign node512 = (inp[3]) ? 3'b010 : node513;
								assign node513 = (inp[4]) ? node515 : 3'b110;
									assign node515 = (inp[5]) ? node521 : node516;
										assign node516 = (inp[2]) ? node518 : 3'b110;
											assign node518 = (inp[0]) ? 3'b010 : 3'b110;
										assign node521 = (inp[1]) ? 3'b010 : node522;
											assign node522 = (inp[2]) ? 3'b010 : node523;
												assign node523 = (inp[0]) ? 3'b010 : 3'b110;
							assign node529 = (inp[3]) ? 3'b100 : node530;
								assign node530 = (inp[1]) ? node532 : 3'b010;
									assign node532 = (inp[5]) ? node534 : 3'b010;
										assign node534 = (inp[0]) ? 3'b100 : 3'b010;
						assign node538 = (inp[3]) ? node548 : node539;
							assign node539 = (inp[8]) ? 3'b100 : node540;
								assign node540 = (inp[4]) ? node542 : 3'b010;
									assign node542 = (inp[5]) ? 3'b100 : node543;
										assign node543 = (inp[0]) ? 3'b100 : 3'b010;
							assign node548 = (inp[8]) ? 3'b000 : node549;
								assign node549 = (inp[0]) ? node551 : 3'b100;
									assign node551 = (inp[2]) ? node553 : 3'b100;
										assign node553 = (inp[5]) ? node555 : 3'b100;
											assign node555 = (inp[4]) ? node557 : 3'b100;
												assign node557 = (inp[1]) ? 3'b000 : 3'b100;
					assign node561 = (inp[11]) ? 3'b000 : node562;
						assign node562 = (inp[8]) ? node574 : node563;
							assign node563 = (inp[3]) ? node569 : node564;
								assign node564 = (inp[2]) ? 3'b100 : node565;
									assign node565 = (inp[4]) ? 3'b100 : 3'b010;
								assign node569 = (inp[4]) ? 3'b000 : node570;
									assign node570 = (inp[5]) ? 3'b000 : 3'b100;
							assign node574 = (inp[4]) ? 3'b000 : node575;
								assign node575 = (inp[3]) ? 3'b000 : node576;
									assign node576 = (inp[5]) ? node582 : node577;
										assign node577 = (inp[1]) ? node579 : 3'b100;
											assign node579 = (inp[0]) ? 3'b000 : 3'b100;
										assign node582 = (inp[0]) ? 3'b000 : node583;
											assign node583 = (inp[1]) ? 3'b000 : 3'b100;
			assign node590 = (inp[10]) ? 3'b000 : node591;
				assign node591 = (inp[7]) ? node631 : node592;
					assign node592 = (inp[11]) ? node620 : node593;
						assign node593 = (inp[8]) ? node609 : node594;
							assign node594 = (inp[3]) ? 3'b100 : node595;
								assign node595 = (inp[4]) ? node597 : 3'b010;
									assign node597 = (inp[0]) ? node603 : node598;
										assign node598 = (inp[1]) ? node600 : 3'b010;
											assign node600 = (inp[5]) ? 3'b100 : 3'b010;
										assign node603 = (inp[1]) ? 3'b100 : node604;
											assign node604 = (inp[5]) ? 3'b100 : 3'b010;
							assign node609 = (inp[3]) ? node611 : 3'b100;
								assign node611 = (inp[1]) ? node613 : 3'b000;
									assign node613 = (inp[2]) ? 3'b000 : node614;
										assign node614 = (inp[5]) ? 3'b000 : node615;
											assign node615 = (inp[0]) ? 3'b000 : 3'b100;
						assign node620 = (inp[3]) ? 3'b000 : node621;
							assign node621 = (inp[8]) ? 3'b000 : node622;
								assign node622 = (inp[4]) ? node624 : 3'b100;
									assign node624 = (inp[0]) ? 3'b000 : node625;
										assign node625 = (inp[5]) ? 3'b000 : 3'b100;
					assign node631 = (inp[5]) ? 3'b000 : node632;
						assign node632 = (inp[11]) ? 3'b000 : node633;
							assign node633 = (inp[3]) ? 3'b000 : node634;
								assign node634 = (inp[8]) ? 3'b000 : node635;
									assign node635 = (inp[1]) ? 3'b000 : 3'b100;

endmodule