module dtc_split75_bm32 (
	input  wire [15-1:0] inp,
	output wire [9-1:0] outp
);

	wire [9-1:0] node1;
	wire [9-1:0] node2;
	wire [9-1:0] node5;
	wire [9-1:0] node6;
	wire [9-1:0] node7;
	wire [9-1:0] node9;
	wire [9-1:0] node11;
	wire [9-1:0] node12;
	wire [9-1:0] node14;
	wire [9-1:0] node18;
	wire [9-1:0] node21;
	wire [9-1:0] node22;
	wire [9-1:0] node24;
	wire [9-1:0] node26;
	wire [9-1:0] node29;
	wire [9-1:0] node30;
	wire [9-1:0] node32;
	wire [9-1:0] node34;
	wire [9-1:0] node35;
	wire [9-1:0] node39;
	wire [9-1:0] node41;
	wire [9-1:0] node42;
	wire [9-1:0] node45;
	wire [9-1:0] node48;
	wire [9-1:0] node49;
	wire [9-1:0] node50;
	wire [9-1:0] node51;
	wire [9-1:0] node52;
	wire [9-1:0] node53;
	wire [9-1:0] node54;
	wire [9-1:0] node55;
	wire [9-1:0] node60;
	wire [9-1:0] node61;
	wire [9-1:0] node62;
	wire [9-1:0] node63;
	wire [9-1:0] node68;
	wire [9-1:0] node71;
	wire [9-1:0] node72;
	wire [9-1:0] node73;
	wire [9-1:0] node74;
	wire [9-1:0] node79;
	wire [9-1:0] node80;
	wire [9-1:0] node81;
	wire [9-1:0] node82;
	wire [9-1:0] node87;
	wire [9-1:0] node90;
	wire [9-1:0] node91;
	wire [9-1:0] node92;
	wire [9-1:0] node93;
	wire [9-1:0] node94;
	wire [9-1:0] node99;
	wire [9-1:0] node100;
	wire [9-1:0] node101;
	wire [9-1:0] node102;
	wire [9-1:0] node107;
	wire [9-1:0] node110;
	wire [9-1:0] node111;
	wire [9-1:0] node112;
	wire [9-1:0] node113;
	wire [9-1:0] node114;
	wire [9-1:0] node116;
	wire [9-1:0] node118;
	wire [9-1:0] node121;
	wire [9-1:0] node123;
	wire [9-1:0] node126;
	wire [9-1:0] node127;
	wire [9-1:0] node128;
	wire [9-1:0] node132;
	wire [9-1:0] node133;
	wire [9-1:0] node134;
	wire [9-1:0] node139;
	wire [9-1:0] node140;
	wire [9-1:0] node143;
	wire [9-1:0] node146;
	wire [9-1:0] node147;
	wire [9-1:0] node148;
	wire [9-1:0] node149;
	wire [9-1:0] node150;
	wire [9-1:0] node154;
	wire [9-1:0] node155;
	wire [9-1:0] node156;
	wire [9-1:0] node161;
	wire [9-1:0] node162;
	wire [9-1:0] node164;
	wire [9-1:0] node166;
	wire [9-1:0] node169;
	wire [9-1:0] node171;
	wire [9-1:0] node174;
	wire [9-1:0] node175;
	wire [9-1:0] node178;
	wire [9-1:0] node181;
	wire [9-1:0] node182;
	wire [9-1:0] node183;
	wire [9-1:0] node184;
	wire [9-1:0] node185;
	wire [9-1:0] node186;
	wire [9-1:0] node191;
	wire [9-1:0] node192;
	wire [9-1:0] node193;
	wire [9-1:0] node194;
	wire [9-1:0] node199;
	wire [9-1:0] node202;
	wire [9-1:0] node203;
	wire [9-1:0] node204;
	wire [9-1:0] node205;
	wire [9-1:0] node210;
	wire [9-1:0] node211;
	wire [9-1:0] node212;
	wire [9-1:0] node213;
	wire [9-1:0] node218;
	wire [9-1:0] node221;
	wire [9-1:0] node222;
	wire [9-1:0] node223;
	wire [9-1:0] node224;
	wire [9-1:0] node225;
	wire [9-1:0] node230;
	wire [9-1:0] node231;
	wire [9-1:0] node232;
	wire [9-1:0] node233;
	wire [9-1:0] node238;
	wire [9-1:0] node241;
	wire [9-1:0] node242;
	wire [9-1:0] node243;
	wire [9-1:0] node244;
	wire [9-1:0] node245;
	wire [9-1:0] node246;
	wire [9-1:0] node248;
	wire [9-1:0] node250;
	wire [9-1:0] node253;
	wire [9-1:0] node255;
	wire [9-1:0] node258;
	wire [9-1:0] node259;
	wire [9-1:0] node260;
	wire [9-1:0] node264;
	wire [9-1:0] node265;
	wire [9-1:0] node266;
	wire [9-1:0] node271;
	wire [9-1:0] node272;
	wire [9-1:0] node275;
	wire [9-1:0] node278;
	wire [9-1:0] node279;
	wire [9-1:0] node280;
	wire [9-1:0] node281;
	wire [9-1:0] node282;
	wire [9-1:0] node286;
	wire [9-1:0] node287;
	wire [9-1:0] node288;
	wire [9-1:0] node293;
	wire [9-1:0] node294;
	wire [9-1:0] node296;
	wire [9-1:0] node298;
	wire [9-1:0] node301;
	wire [9-1:0] node303;
	wire [9-1:0] node306;
	wire [9-1:0] node308;
	wire [9-1:0] node311;
	wire [9-1:0] node312;
	wire [9-1:0] node313;
	wire [9-1:0] node314;
	wire [9-1:0] node315;
	wire [9-1:0] node317;
	wire [9-1:0] node319;
	wire [9-1:0] node322;
	wire [9-1:0] node323;
	wire [9-1:0] node326;
	wire [9-1:0] node329;
	wire [9-1:0] node330;
	wire [9-1:0] node332;
	wire [9-1:0] node334;
	wire [9-1:0] node337;
	wire [9-1:0] node339;
	wire [9-1:0] node342;
	wire [9-1:0] node343;
	wire [9-1:0] node346;
	wire [9-1:0] node349;
	wire [9-1:0] node350;
	wire [9-1:0] node351;
	wire [9-1:0] node352;
	wire [9-1:0] node353;
	wire [9-1:0] node357;
	wire [9-1:0] node358;
	wire [9-1:0] node359;
	wire [9-1:0] node364;
	wire [9-1:0] node365;
	wire [9-1:0] node367;
	wire [9-1:0] node369;
	wire [9-1:0] node372;
	wire [9-1:0] node374;
	wire [9-1:0] node377;
	wire [9-1:0] node378;
	wire [9-1:0] node381;
	wire [9-1:0] node384;
	wire [9-1:0] node385;
	wire [9-1:0] node386;
	wire [9-1:0] node387;
	wire [9-1:0] node389;
	wire [9-1:0] node392;
	wire [9-1:0] node393;
	wire [9-1:0] node396;
	wire [9-1:0] node397;
	wire [9-1:0] node400;
	wire [9-1:0] node401;
	wire [9-1:0] node404;
	wire [9-1:0] node407;
	wire [9-1:0] node408;
	wire [9-1:0] node410;
	wire [9-1:0] node413;
	wire [9-1:0] node414;
	wire [9-1:0] node417;
	wire [9-1:0] node418;
	wire [9-1:0] node421;
	wire [9-1:0] node422;
	wire [9-1:0] node425;
	wire [9-1:0] node428;
	wire [9-1:0] node429;
	wire [9-1:0] node430;
	wire [9-1:0] node431;
	wire [9-1:0] node434;
	wire [9-1:0] node435;
	wire [9-1:0] node438;
	wire [9-1:0] node441;
	wire [9-1:0] node442;
	wire [9-1:0] node445;
	wire [9-1:0] node447;
	wire [9-1:0] node448;
	wire [9-1:0] node451;
	wire [9-1:0] node454;
	wire [9-1:0] node455;
	wire [9-1:0] node456;
	wire [9-1:0] node459;
	wire [9-1:0] node462;
	wire [9-1:0] node463;
	wire [9-1:0] node466;
	wire [9-1:0] node467;
	wire [9-1:0] node468;
	wire [9-1:0] node471;
	wire [9-1:0] node472;
	wire [9-1:0] node475;
	wire [9-1:0] node478;
	wire [9-1:0] node479;
	wire [9-1:0] node482;
	wire [9-1:0] node483;
	wire [9-1:0] node486;

	assign outp = (inp[12]) ? node48 : node1;
		assign node1 = (inp[13]) ? node5 : node2;
			assign node2 = (inp[11]) ? 9'b101010101 : 9'b101010000;
			assign node5 = (inp[14]) ? node21 : node6;
				assign node6 = (inp[0]) ? node18 : node7;
					assign node7 = (inp[3]) ? node9 : 9'b101010001;
						assign node9 = (inp[9]) ? node11 : 9'b100010001;
							assign node11 = (inp[4]) ? 9'b100010001 : node12;
								assign node12 = (inp[8]) ? node14 : 9'b100010001;
									assign node14 = (inp[6]) ? 9'b001010001 : 9'b101010001;
					assign node18 = (inp[3]) ? 9'b000010101 : 9'b101010101;
				assign node21 = (inp[3]) ? node29 : node22;
					assign node22 = (inp[8]) ? node24 : 9'b111010101;
						assign node24 = (inp[4]) ? node26 : 9'b101010101;
							assign node26 = (inp[9]) ? 9'b111010101 : 9'b101010101;
					assign node29 = (inp[0]) ? node39 : node30;
						assign node30 = (inp[8]) ? node32 : 9'b111010111;
							assign node32 = (inp[9]) ? node34 : 9'b101010111;
								assign node34 = (inp[4]) ? 9'b111010111 : node35;
									assign node35 = (inp[6]) ? 9'b011010101 : 9'b111010101;
						assign node39 = (inp[8]) ? node41 : 9'b011010111;
							assign node41 = (inp[4]) ? node45 : node42;
								assign node42 = (inp[9]) ? 9'b000010111 : 9'b001010111;
								assign node45 = (inp[9]) ? 9'b001010101 : 9'b001010111;
		assign node48 = (inp[8]) ? node384 : node49;
			assign node49 = (inp[6]) ? node181 : node50;
				assign node50 = (inp[13]) ? node90 : node51;
					assign node51 = (inp[11]) ? node71 : node52;
						assign node52 = (inp[7]) ? node60 : node53;
							assign node53 = (inp[1]) ? 9'b111011000 : node54;
								assign node54 = (inp[9]) ? 9'b111011000 : node55;
									assign node55 = (inp[2]) ? 9'b111111000 : 9'b111110000;
							assign node60 = (inp[4]) ? node68 : node61;
								assign node61 = (inp[1]) ? 9'b111111000 : node62;
									assign node62 = (inp[2]) ? 9'b111111000 : node63;
										assign node63 = (inp[9]) ? 9'b111111000 : 9'b111110000;
								assign node68 = (inp[9]) ? 9'b111010000 : 9'b111110000;
						assign node71 = (inp[7]) ? node79 : node72;
							assign node72 = (inp[9]) ? 9'b111011100 : node73;
								assign node73 = (inp[1]) ? 9'b111011100 : node74;
									assign node74 = (inp[2]) ? 9'b111111100 : 9'b111110100;
							assign node79 = (inp[4]) ? node87 : node80;
								assign node80 = (inp[1]) ? 9'b111111100 : node81;
									assign node81 = (inp[2]) ? 9'b111111100 : node82;
										assign node82 = (inp[9]) ? 9'b111111100 : 9'b111110100;
								assign node87 = (inp[9]) ? 9'b111010100 : 9'b111110100;
					assign node90 = (inp[3]) ? node110 : node91;
						assign node91 = (inp[7]) ? node99 : node92;
							assign node92 = (inp[1]) ? 9'b111011100 : node93;
								assign node93 = (inp[9]) ? 9'b111011100 : node94;
									assign node94 = (inp[2]) ? 9'b111111100 : 9'b111110100;
							assign node99 = (inp[4]) ? node107 : node100;
								assign node100 = (inp[9]) ? 9'b111111100 : node101;
									assign node101 = (inp[2]) ? 9'b111111100 : node102;
										assign node102 = (inp[1]) ? 9'b111111100 : 9'b111110100;
								assign node107 = (inp[9]) ? 9'b111010100 : 9'b111110100;
						assign node110 = (inp[14]) ? node146 : node111;
							assign node111 = (inp[9]) ? node139 : node112;
								assign node112 = (inp[10]) ? node126 : node113;
									assign node113 = (inp[1]) ? node121 : node114;
										assign node114 = (inp[2]) ? node116 : 9'b110110100;
											assign node116 = (inp[7]) ? node118 : 9'b110111100;
												assign node118 = (inp[4]) ? 9'b110110100 : 9'b110111100;
										assign node121 = (inp[7]) ? node123 : 9'b110011100;
											assign node123 = (inp[4]) ? 9'b110110100 : 9'b110111100;
									assign node126 = (inp[7]) ? node132 : node127;
										assign node127 = (inp[1]) ? 9'b110011110 : node128;
											assign node128 = (inp[2]) ? 9'b110111110 : 9'b110110110;
										assign node132 = (inp[4]) ? 9'b110110110 : node133;
											assign node133 = (inp[1]) ? 9'b110111110 : node134;
												assign node134 = (inp[2]) ? 9'b110111110 : 9'b110110110;
								assign node139 = (inp[4]) ? node143 : node140;
									assign node140 = (inp[7]) ? 9'b110111110 : 9'b110011110;
									assign node143 = (inp[7]) ? 9'b110010110 : 9'b110011110;
							assign node146 = (inp[9]) ? node174 : node147;
								assign node147 = (inp[10]) ? node161 : node148;
									assign node148 = (inp[7]) ? node154 : node149;
										assign node149 = (inp[1]) ? 9'b111011100 : node150;
											assign node150 = (inp[2]) ? 9'b111111100 : 9'b111110100;
										assign node154 = (inp[4]) ? 9'b111110100 : node155;
											assign node155 = (inp[2]) ? 9'b111111100 : node156;
												assign node156 = (inp[1]) ? 9'b111111100 : 9'b111110100;
									assign node161 = (inp[1]) ? node169 : node162;
										assign node162 = (inp[2]) ? node164 : 9'b111110110;
											assign node164 = (inp[4]) ? node166 : 9'b111111110;
												assign node166 = (inp[7]) ? 9'b111110110 : 9'b111111110;
										assign node169 = (inp[7]) ? node171 : 9'b111011110;
											assign node171 = (inp[4]) ? 9'b111110110 : 9'b111111110;
								assign node174 = (inp[4]) ? node178 : node175;
									assign node175 = (inp[7]) ? 9'b111111110 : 9'b111011110;
									assign node178 = (inp[7]) ? 9'b111010110 : 9'b111011110;
				assign node181 = (inp[13]) ? node221 : node182;
					assign node182 = (inp[11]) ? node202 : node183;
						assign node183 = (inp[7]) ? node191 : node184;
							assign node184 = (inp[1]) ? 9'b111011000 : node185;
								assign node185 = (inp[9]) ? 9'b111011000 : node186;
									assign node186 = (inp[2]) ? 9'b111111000 : 9'b111110000;
							assign node191 = (inp[4]) ? node199 : node192;
								assign node192 = (inp[1]) ? 9'b111111000 : node193;
									assign node193 = (inp[9]) ? 9'b111111000 : node194;
										assign node194 = (inp[2]) ? 9'b111111000 : 9'b111110000;
								assign node199 = (inp[9]) ? 9'b111010000 : 9'b111110000;
						assign node202 = (inp[7]) ? node210 : node203;
							assign node203 = (inp[9]) ? 9'b111011101 : node204;
								assign node204 = (inp[1]) ? 9'b111011101 : node205;
									assign node205 = (inp[2]) ? 9'b111111101 : 9'b111110101;
							assign node210 = (inp[4]) ? node218 : node211;
								assign node211 = (inp[1]) ? 9'b111111101 : node212;
									assign node212 = (inp[9]) ? 9'b111111101 : node213;
										assign node213 = (inp[2]) ? 9'b111111101 : 9'b111110101;
								assign node218 = (inp[9]) ? 9'b111010101 : 9'b111110101;
					assign node221 = (inp[3]) ? node241 : node222;
						assign node222 = (inp[7]) ? node230 : node223;
							assign node223 = (inp[9]) ? 9'b111011101 : node224;
								assign node224 = (inp[1]) ? 9'b111011101 : node225;
									assign node225 = (inp[2]) ? 9'b111111101 : 9'b111110101;
							assign node230 = (inp[4]) ? node238 : node231;
								assign node231 = (inp[9]) ? 9'b111111101 : node232;
									assign node232 = (inp[2]) ? 9'b111111101 : node233;
										assign node233 = (inp[1]) ? 9'b111111101 : 9'b111110101;
								assign node238 = (inp[9]) ? 9'b111010101 : 9'b111110101;
						assign node241 = (inp[5]) ? node311 : node242;
							assign node242 = (inp[14]) ? node278 : node243;
								assign node243 = (inp[9]) ? node271 : node244;
									assign node244 = (inp[10]) ? node258 : node245;
										assign node245 = (inp[1]) ? node253 : node246;
											assign node246 = (inp[2]) ? node248 : 9'b110100101;
												assign node248 = (inp[7]) ? node250 : 9'b110101101;
													assign node250 = (inp[4]) ? 9'b110100101 : 9'b110101101;
											assign node253 = (inp[7]) ? node255 : 9'b110001101;
												assign node255 = (inp[4]) ? 9'b110100101 : 9'b110101101;
										assign node258 = (inp[7]) ? node264 : node259;
											assign node259 = (inp[1]) ? 9'b110001111 : node260;
												assign node260 = (inp[2]) ? 9'b110101111 : 9'b110100111;
											assign node264 = (inp[4]) ? 9'b110100111 : node265;
												assign node265 = (inp[2]) ? 9'b110101111 : node266;
													assign node266 = (inp[1]) ? 9'b110101111 : 9'b110100111;
									assign node271 = (inp[4]) ? node275 : node272;
										assign node272 = (inp[7]) ? 9'b110101111 : 9'b110001111;
										assign node275 = (inp[7]) ? 9'b110000111 : 9'b110001111;
								assign node278 = (inp[9]) ? node306 : node279;
									assign node279 = (inp[10]) ? node293 : node280;
										assign node280 = (inp[7]) ? node286 : node281;
											assign node281 = (inp[1]) ? 9'b111001101 : node282;
												assign node282 = (inp[2]) ? 9'b111101101 : 9'b111100101;
											assign node286 = (inp[4]) ? 9'b111100101 : node287;
												assign node287 = (inp[1]) ? 9'b111101101 : node288;
													assign node288 = (inp[2]) ? 9'b111101101 : 9'b111100101;
										assign node293 = (inp[1]) ? node301 : node294;
											assign node294 = (inp[2]) ? node296 : 9'b111100111;
												assign node296 = (inp[7]) ? node298 : 9'b111101111;
													assign node298 = (inp[4]) ? 9'b111100111 : 9'b111101111;
											assign node301 = (inp[7]) ? node303 : 9'b111001111;
												assign node303 = (inp[4]) ? 9'b111100111 : 9'b111101111;
									assign node306 = (inp[7]) ? node308 : 9'b111001111;
										assign node308 = (inp[4]) ? 9'b111000111 : 9'b111101111;
							assign node311 = (inp[14]) ? node349 : node312;
								assign node312 = (inp[9]) ? node342 : node313;
									assign node313 = (inp[10]) ? node329 : node314;
										assign node314 = (inp[2]) ? node322 : node315;
											assign node315 = (inp[1]) ? node317 : 9'b110110101;
												assign node317 = (inp[7]) ? node319 : 9'b110011101;
													assign node319 = (inp[4]) ? 9'b110110101 : 9'b110111101;
											assign node322 = (inp[7]) ? node326 : node323;
												assign node323 = (inp[1]) ? 9'b110011101 : 9'b110111101;
												assign node326 = (inp[4]) ? 9'b110110101 : 9'b110111101;
										assign node329 = (inp[1]) ? node337 : node330;
											assign node330 = (inp[2]) ? node332 : 9'b110110111;
												assign node332 = (inp[7]) ? node334 : 9'b110111111;
													assign node334 = (inp[4]) ? 9'b110110111 : 9'b110111111;
											assign node337 = (inp[7]) ? node339 : 9'b110011111;
												assign node339 = (inp[4]) ? 9'b110110111 : 9'b110111111;
									assign node342 = (inp[4]) ? node346 : node343;
										assign node343 = (inp[7]) ? 9'b110111111 : 9'b110011111;
										assign node346 = (inp[7]) ? 9'b110010111 : 9'b110011111;
								assign node349 = (inp[9]) ? node377 : node350;
									assign node350 = (inp[10]) ? node364 : node351;
										assign node351 = (inp[7]) ? node357 : node352;
											assign node352 = (inp[1]) ? 9'b111011101 : node353;
												assign node353 = (inp[2]) ? 9'b111111101 : 9'b111110101;
											assign node357 = (inp[4]) ? 9'b111110101 : node358;
												assign node358 = (inp[2]) ? 9'b111111101 : node359;
													assign node359 = (inp[1]) ? 9'b111111101 : 9'b111110101;
										assign node364 = (inp[1]) ? node372 : node365;
											assign node365 = (inp[2]) ? node367 : 9'b111110111;
												assign node367 = (inp[7]) ? node369 : 9'b111111111;
													assign node369 = (inp[4]) ? 9'b111110111 : 9'b111111111;
											assign node372 = (inp[7]) ? node374 : 9'b111011111;
												assign node374 = (inp[4]) ? 9'b111110111 : 9'b111111111;
									assign node377 = (inp[4]) ? node381 : node378;
										assign node378 = (inp[7]) ? 9'b111111111 : 9'b111011111;
										assign node381 = (inp[7]) ? 9'b111010111 : 9'b111011111;
			assign node384 = (inp[9]) ? node428 : node385;
				assign node385 = (inp[4]) ? node407 : node386;
					assign node386 = (inp[13]) ? node392 : node387;
						assign node387 = (inp[11]) ? node389 : 9'b101111000;
							assign node389 = (inp[6]) ? 9'b101111101 : 9'b101111100;
						assign node392 = (inp[3]) ? node396 : node393;
							assign node393 = (inp[6]) ? 9'b101111101 : 9'b101111100;
							assign node396 = (inp[6]) ? node400 : node397;
								assign node397 = (inp[14]) ? 9'b101111110 : 9'b100111110;
								assign node400 = (inp[14]) ? node404 : node401;
									assign node401 = (inp[5]) ? 9'b100111111 : 9'b100101111;
									assign node404 = (inp[5]) ? 9'b101111111 : 9'b101101111;
					assign node407 = (inp[13]) ? node413 : node408;
						assign node408 = (inp[11]) ? node410 : 9'b101010000;
							assign node410 = (inp[6]) ? 9'b101010101 : 9'b101010100;
						assign node413 = (inp[3]) ? node417 : node414;
							assign node414 = (inp[6]) ? 9'b101010101 : 9'b101010100;
							assign node417 = (inp[6]) ? node421 : node418;
								assign node418 = (inp[14]) ? 9'b101010110 : 9'b100010110;
								assign node421 = (inp[14]) ? node425 : node422;
									assign node422 = (inp[5]) ? 9'b100010111 : 9'b100000111;
									assign node425 = (inp[5]) ? 9'b101010111 : 9'b101000111;
				assign node428 = (inp[6]) ? node454 : node429;
					assign node429 = (inp[4]) ? node441 : node430;
						assign node430 = (inp[13]) ? node434 : node431;
							assign node431 = (inp[11]) ? 9'b101010100 : 9'b101010000;
							assign node434 = (inp[0]) ? node438 : node435;
								assign node435 = (inp[3]) ? 9'b111010100 : 9'b101010100;
								assign node438 = (inp[3]) ? 9'b100010110 : 9'b101010100;
						assign node441 = (inp[13]) ? node445 : node442;
							assign node442 = (inp[11]) ? 9'b111010100 : 9'b111010000;
							assign node445 = (inp[3]) ? node447 : 9'b111010100;
								assign node447 = (inp[0]) ? node451 : node448;
									assign node448 = (inp[14]) ? 9'b111010110 : 9'b110010110;
									assign node451 = (inp[14]) ? 9'b101010100 : 9'b100010100;
					assign node454 = (inp[13]) ? node462 : node455;
						assign node455 = (inp[11]) ? node459 : node456;
							assign node456 = (inp[4]) ? 9'b111010000 : 9'b101010000;
							assign node459 = (inp[4]) ? 9'b111010101 : 9'b101010101;
						assign node462 = (inp[3]) ? node466 : node463;
							assign node463 = (inp[4]) ? 9'b111010101 : 9'b101010101;
							assign node466 = (inp[0]) ? node478 : node467;
								assign node467 = (inp[4]) ? node471 : node468;
									assign node468 = (inp[5]) ? 9'b011010101 : 9'b011000101;
									assign node471 = (inp[14]) ? node475 : node472;
										assign node472 = (inp[5]) ? 9'b110010111 : 9'b110000111;
										assign node475 = (inp[5]) ? 9'b111010111 : 9'b111000111;
								assign node478 = (inp[4]) ? node482 : node479;
									assign node479 = (inp[5]) ? 9'b100010111 : 9'b100000111;
									assign node482 = (inp[14]) ? node486 : node483;
										assign node483 = (inp[5]) ? 9'b100010101 : 9'b100000101;
										assign node486 = (inp[5]) ? 9'b101010101 : 9'b101000101;

endmodule