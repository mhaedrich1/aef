module dtc_split33_bm19 (
	input  wire [8-1:0] inp,
	output wire [8-1:0] outp
);

	wire [8-1:0] node1;
	wire [8-1:0] node2;
	wire [8-1:0] node3;
	wire [8-1:0] node4;
	wire [8-1:0] node5;
	wire [8-1:0] node6;
	wire [8-1:0] node9;
	wire [8-1:0] node12;
	wire [8-1:0] node15;
	wire [8-1:0] node17;
	wire [8-1:0] node20;
	wire [8-1:0] node21;
	wire [8-1:0] node22;
	wire [8-1:0] node25;
	wire [8-1:0] node26;
	wire [8-1:0] node30;
	wire [8-1:0] node31;
	wire [8-1:0] node35;
	wire [8-1:0] node36;
	wire [8-1:0] node37;
	wire [8-1:0] node40;
	wire [8-1:0] node41;
	wire [8-1:0] node42;
	wire [8-1:0] node46;
	wire [8-1:0] node48;
	wire [8-1:0] node51;
	wire [8-1:0] node52;
	wire [8-1:0] node54;
	wire [8-1:0] node55;
	wire [8-1:0] node59;
	wire [8-1:0] node61;
	wire [8-1:0] node62;
	wire [8-1:0] node65;
	wire [8-1:0] node68;
	wire [8-1:0] node69;
	wire [8-1:0] node70;
	wire [8-1:0] node71;
	wire [8-1:0] node72;
	wire [8-1:0] node75;
	wire [8-1:0] node76;
	wire [8-1:0] node80;
	wire [8-1:0] node82;
	wire [8-1:0] node85;
	wire [8-1:0] node86;
	wire [8-1:0] node87;
	wire [8-1:0] node90;
	wire [8-1:0] node91;
	wire [8-1:0] node94;
	wire [8-1:0] node98;
	wire [8-1:0] node99;
	wire [8-1:0] node100;
	wire [8-1:0] node101;
	wire [8-1:0] node104;
	wire [8-1:0] node107;
	wire [8-1:0] node109;
	wire [8-1:0] node111;
	wire [8-1:0] node114;
	wire [8-1:0] node115;
	wire [8-1:0] node117;
	wire [8-1:0] node120;
	wire [8-1:0] node122;

	assign outp = (inp[5]) ? node68 : node1;
		assign node1 = (inp[3]) ? node35 : node2;
			assign node2 = (inp[7]) ? node20 : node3;
				assign node3 = (inp[2]) ? node15 : node4;
					assign node4 = (inp[1]) ? node12 : node5;
						assign node5 = (inp[0]) ? node9 : node6;
							assign node6 = (inp[4]) ? 8'b00111111 : 8'b01111111;
							assign node9 = (inp[6]) ? 8'b00011111 : 8'b00111111;
						assign node12 = (inp[4]) ? 8'b00011111 : 8'b00111111;
					assign node15 = (inp[1]) ? node17 : 8'b00011111;
						assign node17 = (inp[4]) ? 8'b00001111 : 8'b00011111;
				assign node20 = (inp[1]) ? node30 : node21;
					assign node21 = (inp[4]) ? node25 : node22;
						assign node22 = (inp[2]) ? 8'b00011111 : 8'b00111111;
						assign node25 = (inp[2]) ? 8'b00001111 : node26;
							assign node26 = (inp[0]) ? 8'b00001111 : 8'b00011111;
					assign node30 = (inp[6]) ? 8'b00001111 : node31;
						assign node31 = (inp[0]) ? 8'b00001111 : 8'b00011111;
			assign node35 = (inp[0]) ? node51 : node36;
				assign node36 = (inp[1]) ? node40 : node37;
					assign node37 = (inp[4]) ? 8'b00011111 : 8'b00111111;
					assign node40 = (inp[4]) ? node46 : node41;
						assign node41 = (inp[2]) ? 8'b00001111 : node42;
							assign node42 = (inp[6]) ? 8'b00011111 : 8'b00111111;
						assign node46 = (inp[7]) ? node48 : 8'b00001111;
							assign node48 = (inp[6]) ? 8'b00000111 : 8'b00001111;
				assign node51 = (inp[6]) ? node59 : node52;
					assign node52 = (inp[7]) ? node54 : 8'b00001111;
						assign node54 = (inp[1]) ? 8'b00000111 : node55;
							assign node55 = (inp[2]) ? 8'b00000111 : 8'b00001111;
					assign node59 = (inp[4]) ? node61 : 8'b00011111;
						assign node61 = (inp[7]) ? node65 : node62;
							assign node62 = (inp[2]) ? 8'b00000011 : 8'b00000111;
							assign node65 = (inp[2]) ? 8'b00000001 : 8'b00000011;
		assign node68 = (inp[1]) ? node98 : node69;
			assign node69 = (inp[0]) ? node85 : node70;
				assign node70 = (inp[7]) ? node80 : node71;
					assign node71 = (inp[6]) ? node75 : node72;
						assign node72 = (inp[3]) ? 8'b00011111 : 8'b00111111;
						assign node75 = (inp[4]) ? 8'b00001111 : node76;
							assign node76 = (inp[2]) ? 8'b00001111 : 8'b00011111;
					assign node80 = (inp[4]) ? node82 : 8'b00001111;
						assign node82 = (inp[3]) ? 8'b00000011 : 8'b00001111;
				assign node85 = (inp[2]) ? 8'b00000111 : node86;
					assign node86 = (inp[4]) ? node90 : node87;
						assign node87 = (inp[3]) ? 8'b00001111 : 8'b00011111;
						assign node90 = (inp[6]) ? node94 : node91;
							assign node91 = (inp[3]) ? 8'b00000111 : 8'b00001111;
							assign node94 = (inp[3]) ? 8'b00000011 : 8'b00000111;
			assign node98 = (inp[2]) ? node114 : node99;
				assign node99 = (inp[6]) ? node107 : node100;
					assign node100 = (inp[7]) ? node104 : node101;
						assign node101 = (inp[0]) ? 8'b00001111 : 8'b00011111;
						assign node104 = (inp[0]) ? 8'b00000111 : 8'b00001111;
					assign node107 = (inp[3]) ? node109 : 8'b00000111;
						assign node109 = (inp[4]) ? node111 : 8'b00000111;
							assign node111 = (inp[7]) ? 8'b00000011 : 8'b00000111;
				assign node114 = (inp[4]) ? node120 : node115;
					assign node115 = (inp[3]) ? node117 : 8'b00001111;
						assign node117 = (inp[0]) ? 8'b00000011 : 8'b00000111;
					assign node120 = (inp[6]) ? node122 : 8'b00000011;
						assign node122 = (inp[7]) ? 8'b00000000 : 8'b00000001;

endmodule