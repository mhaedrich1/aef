module dtc_split5_bm55 (
	input  wire [8-1:0] inp,
	output wire [7-1:0] outp
);

	wire [7-1:0] node1;
	wire [7-1:0] node2;
	wire [7-1:0] node3;
	wire [7-1:0] node4;
	wire [7-1:0] node6;
	wire [7-1:0] node7;
	wire [7-1:0] node10;
	wire [7-1:0] node13;
	wire [7-1:0] node16;
	wire [7-1:0] node17;
	wire [7-1:0] node18;
	wire [7-1:0] node19;
	wire [7-1:0] node22;
	wire [7-1:0] node25;
	wire [7-1:0] node28;
	wire [7-1:0] node29;
	wire [7-1:0] node30;
	wire [7-1:0] node33;
	wire [7-1:0] node34;
	wire [7-1:0] node37;
	wire [7-1:0] node40;
	wire [7-1:0] node42;
	wire [7-1:0] node43;
	wire [7-1:0] node47;
	wire [7-1:0] node48;
	wire [7-1:0] node49;
	wire [7-1:0] node50;
	wire [7-1:0] node52;
	wire [7-1:0] node53;
	wire [7-1:0] node57;
	wire [7-1:0] node59;
	wire [7-1:0] node62;
	wire [7-1:0] node63;
	wire [7-1:0] node64;
	wire [7-1:0] node66;
	wire [7-1:0] node69;
	wire [7-1:0] node71;
	wire [7-1:0] node74;
	wire [7-1:0] node76;
	wire [7-1:0] node79;
	wire [7-1:0] node80;
	wire [7-1:0] node81;
	wire [7-1:0] node82;
	wire [7-1:0] node83;
	wire [7-1:0] node87;
	wire [7-1:0] node90;
	wire [7-1:0] node91;
	wire [7-1:0] node95;
	wire [7-1:0] node96;
	wire [7-1:0] node97;
	wire [7-1:0] node100;
	wire [7-1:0] node102;
	wire [7-1:0] node105;
	wire [7-1:0] node106;
	wire [7-1:0] node110;
	wire [7-1:0] node111;
	wire [7-1:0] node112;
	wire [7-1:0] node113;
	wire [7-1:0] node114;
	wire [7-1:0] node117;
	wire [7-1:0] node118;
	wire [7-1:0] node119;
	wire [7-1:0] node123;
	wire [7-1:0] node126;
	wire [7-1:0] node127;
	wire [7-1:0] node128;
	wire [7-1:0] node129;
	wire [7-1:0] node133;
	wire [7-1:0] node136;
	wire [7-1:0] node137;
	wire [7-1:0] node140;
	wire [7-1:0] node143;
	wire [7-1:0] node144;
	wire [7-1:0] node145;
	wire [7-1:0] node147;
	wire [7-1:0] node148;
	wire [7-1:0] node152;
	wire [7-1:0] node153;
	wire [7-1:0] node157;
	wire [7-1:0] node158;
	wire [7-1:0] node159;
	wire [7-1:0] node162;
	wire [7-1:0] node164;
	wire [7-1:0] node167;
	wire [7-1:0] node169;
	wire [7-1:0] node172;
	wire [7-1:0] node173;
	wire [7-1:0] node174;
	wire [7-1:0] node175;
	wire [7-1:0] node177;
	wire [7-1:0] node180;
	wire [7-1:0] node181;
	wire [7-1:0] node182;
	wire [7-1:0] node186;
	wire [7-1:0] node187;
	wire [7-1:0] node191;
	wire [7-1:0] node192;
	wire [7-1:0] node193;
	wire [7-1:0] node194;
	wire [7-1:0] node198;
	wire [7-1:0] node199;
	wire [7-1:0] node202;
	wire [7-1:0] node205;
	wire [7-1:0] node206;
	wire [7-1:0] node210;
	wire [7-1:0] node211;
	wire [7-1:0] node212;
	wire [7-1:0] node213;
	wire [7-1:0] node215;
	wire [7-1:0] node218;
	wire [7-1:0] node221;
	wire [7-1:0] node223;
	wire [7-1:0] node226;
	wire [7-1:0] node227;
	wire [7-1:0] node228;
	wire [7-1:0] node230;
	wire [7-1:0] node234;
	wire [7-1:0] node235;

	assign outp = (inp[6]) ? node110 : node1;
		assign node1 = (inp[2]) ? node47 : node2;
			assign node2 = (inp[4]) ? node16 : node3;
				assign node3 = (inp[3]) ? node13 : node4;
					assign node4 = (inp[5]) ? node6 : 7'b0110101;
						assign node6 = (inp[7]) ? node10 : node7;
							assign node7 = (inp[1]) ? 7'b0101101 : 7'b0100101;
							assign node10 = (inp[1]) ? 7'b1100101 : 7'b0100101;
					assign node13 = (inp[5]) ? 7'b1100100 : 7'b1111100;
				assign node16 = (inp[7]) ? node28 : node17;
					assign node17 = (inp[1]) ? node25 : node18;
						assign node18 = (inp[5]) ? node22 : node19;
							assign node19 = (inp[3]) ? 7'b1101110 : 7'b0111100;
							assign node22 = (inp[0]) ? 7'b1100100 : 7'b1001100;
						assign node25 = (inp[5]) ? 7'b0001101 : 7'b0000111;
					assign node28 = (inp[3]) ? node40 : node29;
						assign node29 = (inp[0]) ? node33 : node30;
							assign node30 = (inp[1]) ? 7'b1000111 : 7'b1000101;
							assign node33 = (inp[5]) ? node37 : node34;
								assign node34 = (inp[1]) ? 7'b1010110 : 7'b0101110;
								assign node37 = (inp[1]) ? 7'b0010100 : 7'b1110100;
						assign node40 = (inp[0]) ? node42 : 7'b0000100;
							assign node42 = (inp[5]) ? 7'b0000101 : node43;
								assign node43 = (inp[1]) ? 7'b1000100 : 7'b1000101;
			assign node47 = (inp[0]) ? node79 : node48;
				assign node48 = (inp[1]) ? node62 : node49;
					assign node49 = (inp[4]) ? node57 : node50;
						assign node50 = (inp[7]) ? node52 : 7'b0110011;
							assign node52 = (inp[5]) ? 7'b0100001 : node53;
								assign node53 = (inp[3]) ? 7'b0101001 : 7'b0100011;
						assign node57 = (inp[3]) ? node59 : 7'b0101000;
							assign node59 = (inp[7]) ? 7'b0110001 : 7'b1111001;
					assign node62 = (inp[5]) ? node74 : node63;
						assign node63 = (inp[7]) ? node69 : node64;
							assign node64 = (inp[3]) ? node66 : 7'b0110000;
								assign node66 = (inp[4]) ? 7'b0110010 : 7'b1111010;
							assign node69 = (inp[3]) ? node71 : 7'b1110010;
								assign node71 = (inp[4]) ? 7'b1100000 : 7'b1101000;
						assign node74 = (inp[3]) ? node76 : 7'b0110000;
							assign node76 = (inp[7]) ? 7'b0100000 : 7'b1100000;
				assign node79 = (inp[4]) ? node95 : node80;
					assign node80 = (inp[1]) ? node90 : node81;
						assign node81 = (inp[5]) ? node87 : node82;
							assign node82 = (inp[7]) ? 7'b1100010 : node83;
								assign node83 = (inp[3]) ? 7'b0100010 : 7'b0110000;
							assign node87 = (inp[3]) ? 7'b0010001 : 7'b0100000;
						assign node90 = (inp[3]) ? 7'b1001001 : node91;
							assign node91 = (inp[7]) ? 7'b0001011 : 7'b1001001;
					assign node95 = (inp[3]) ? node105 : node96;
						assign node96 = (inp[5]) ? node100 : node97;
							assign node97 = (inp[7]) ? 7'b0011010 : 7'b0001001;
							assign node100 = (inp[1]) ? node102 : 7'b1010000;
								assign node102 = (inp[7]) ? 7'b0010000 : 7'b0011000;
						assign node105 = (inp[5]) ? 7'b0001000 : node106;
							assign node106 = (inp[7]) ? 7'b1000000 : 7'b1000010;
		assign node110 = (inp[5]) ? node172 : node111;
			assign node111 = (inp[0]) ? node143 : node112;
				assign node112 = (inp[4]) ? node126 : node113;
					assign node113 = (inp[3]) ? node117 : node114;
						assign node114 = (inp[1]) ? 7'b1010100 : 7'b1010111;
						assign node117 = (inp[1]) ? node123 : node118;
							assign node118 = (inp[7]) ? 7'b1001100 : node119;
								assign node119 = (inp[2]) ? 7'b1000011 : 7'b1000111;
							assign node123 = (inp[2]) ? 7'b0011011 : 7'b0101011;
					assign node126 = (inp[2]) ? node136 : node127;
						assign node127 = (inp[7]) ? node133 : node128;
							assign node128 = (inp[1]) ? 7'b1101001 : node129;
								assign node129 = (inp[3]) ? 7'b0111010 : 7'b1111000;
							assign node133 = (inp[3]) ? 7'b1110001 : 7'b0110011;
						assign node136 = (inp[3]) ? node140 : node137;
							assign node137 = (inp[1]) ? 7'b1001000 : 7'b1001001;
							assign node140 = (inp[1]) ? 7'b1000010 : 7'b1010000;
				assign node143 = (inp[1]) ? node157 : node144;
					assign node144 = (inp[2]) ? node152 : node145;
						assign node145 = (inp[4]) ? node147 : 7'b1000011;
							assign node147 = (inp[7]) ? 7'b0000001 : node148;
								assign node148 = (inp[3]) ? 7'b0011011 : 7'b1011001;
						assign node152 = (inp[4]) ? 7'b1001000 : node153;
							assign node153 = (inp[3]) ? 7'b1010010 : 7'b1010000;
					assign node157 = (inp[4]) ? node167 : node158;
						assign node158 = (inp[3]) ? node162 : node159;
							assign node159 = (inp[7]) ? 7'b1001010 : 7'b0000001;
							assign node162 = (inp[7]) ? node164 : 7'b0001010;
								assign node164 = (inp[2]) ? 7'b0001000 : 7'b0011000;
						assign node167 = (inp[7]) ? node169 : 7'b0011000;
							assign node169 = (inp[3]) ? 7'b0000000 : 7'b0000010;
			assign node172 = (inp[7]) ? node210 : node173;
				assign node173 = (inp[2]) ? node191 : node174;
					assign node174 = (inp[0]) ? node180 : node175;
						assign node175 = (inp[1]) ? node177 : 7'b0110000;
							assign node177 = (inp[3]) ? 7'b1110000 : 7'b1111001;
						assign node180 = (inp[4]) ? node186 : node181;
							assign node181 = (inp[3]) ? 7'b1001001 : node182;
								assign node182 = (inp[1]) ? 7'b1011000 : 7'b1100000;
							assign node186 = (inp[1]) ? 7'b0011000 : node187;
								assign node187 = (inp[3]) ? 7'b0011001 : 7'b1010001;
					assign node191 = (inp[0]) ? node205 : node192;
						assign node192 = (inp[3]) ? node198 : node193;
							assign node193 = (inp[4]) ? 7'b0000001 : node194;
								assign node194 = (inp[1]) ? 7'b0011001 : 7'b0010001;
							assign node198 = (inp[1]) ? node202 : node199;
								assign node199 = (inp[4]) ? 7'b1011000 : 7'b0001001;
								assign node202 = (inp[4]) ? 7'b1000000 : 7'b1000001;
						assign node205 = (inp[1]) ? 7'b1001000 : node206;
							assign node206 = (inp[4]) ? 7'b1000000 : 7'b1010000;
				assign node210 = (inp[0]) ? node226 : node211;
					assign node211 = (inp[4]) ? node221 : node212;
						assign node212 = (inp[1]) ? node218 : node213;
							assign node213 = (inp[2]) ? node215 : 7'b0010101;
								assign node215 = (inp[3]) ? 7'b0000001 : 7'b0010001;
							assign node218 = (inp[2]) ? 7'b1010001 : 7'b1110001;
						assign node221 = (inp[3]) ? node223 : 7'b1110000;
							assign node223 = (inp[2]) ? 7'b0010000 : 7'b0100000;
					assign node226 = (inp[1]) ? node234 : node227;
						assign node227 = (inp[2]) ? 7'b0000000 : node228;
							assign node228 = (inp[4]) ? node230 : 7'b0010001;
								assign node230 = (inp[3]) ? 7'b0000001 : 7'b1000001;
						assign node234 = (inp[2]) ? 7'b0000000 : node235;
							assign node235 = (inp[4]) ? 7'b0000000 : 7'b1000000;

endmodule