module dtc_split75_bm51 (
	input  wire [8-1:0] inp,
	output wire [2-1:0] outp
);

	wire [2-1:0] node1;
	wire [2-1:0] node2;
	wire [2-1:0] node3;
	wire [2-1:0] node4;
	wire [2-1:0] node5;
	wire [2-1:0] node6;
	wire [2-1:0] node8;
	wire [2-1:0] node11;
	wire [2-1:0] node13;
	wire [2-1:0] node16;
	wire [2-1:0] node17;
	wire [2-1:0] node19;
	wire [2-1:0] node22;
	wire [2-1:0] node25;
	wire [2-1:0] node26;
	wire [2-1:0] node29;
	wire [2-1:0] node32;
	wire [2-1:0] node33;
	wire [2-1:0] node34;
	wire [2-1:0] node35;
	wire [2-1:0] node36;
	wire [2-1:0] node39;
	wire [2-1:0] node43;
	wire [2-1:0] node45;
	wire [2-1:0] node46;
	wire [2-1:0] node50;
	wire [2-1:0] node51;
	wire [2-1:0] node52;
	wire [2-1:0] node56;
	wire [2-1:0] node57;
	wire [2-1:0] node61;
	wire [2-1:0] node62;
	wire [2-1:0] node63;
	wire [2-1:0] node64;
	wire [2-1:0] node65;
	wire [2-1:0] node68;
	wire [2-1:0] node71;
	wire [2-1:0] node72;
	wire [2-1:0] node75;
	wire [2-1:0] node78;
	wire [2-1:0] node79;
	wire [2-1:0] node82;
	wire [2-1:0] node85;
	wire [2-1:0] node86;
	wire [2-1:0] node87;
	wire [2-1:0] node91;
	wire [2-1:0] node92;
	wire [2-1:0] node96;
	wire [2-1:0] node97;
	wire [2-1:0] node98;
	wire [2-1:0] node99;
	wire [2-1:0] node100;
	wire [2-1:0] node103;
	wire [2-1:0] node105;
	wire [2-1:0] node106;
	wire [2-1:0] node110;
	wire [2-1:0] node111;
	wire [2-1:0] node114;
	wire [2-1:0] node117;
	wire [2-1:0] node118;
	wire [2-1:0] node119;
	wire [2-1:0] node123;
	wire [2-1:0] node124;
	wire [2-1:0] node128;
	wire [2-1:0] node129;
	wire [2-1:0] node130;
	wire [2-1:0] node131;
	wire [2-1:0] node132;
	wire [2-1:0] node133;
	wire [2-1:0] node137;
	wire [2-1:0] node141;
	wire [2-1:0] node142;
	wire [2-1:0] node144;
	wire [2-1:0] node148;
	wire [2-1:0] node149;

	assign outp = (inp[6]) ? node96 : node1;
		assign node1 = (inp[2]) ? node61 : node2;
			assign node2 = (inp[7]) ? node32 : node3;
				assign node3 = (inp[0]) ? node25 : node4;
					assign node4 = (inp[5]) ? node16 : node5;
						assign node5 = (inp[4]) ? node11 : node6;
							assign node6 = (inp[3]) ? node8 : 2'b00;
								assign node8 = (inp[1]) ? 2'b01 : 2'b00;
							assign node11 = (inp[3]) ? node13 : 2'b01;
								assign node13 = (inp[1]) ? 2'b00 : 2'b01;
						assign node16 = (inp[4]) ? node22 : node17;
							assign node17 = (inp[1]) ? node19 : 2'b01;
								assign node19 = (inp[3]) ? 2'b00 : 2'b01;
							assign node22 = (inp[1]) ? 2'b01 : 2'b00;
					assign node25 = (inp[3]) ? node29 : node26;
						assign node26 = (inp[5]) ? 2'b11 : 2'b10;
						assign node29 = (inp[5]) ? 2'b10 : 2'b11;
				assign node32 = (inp[3]) ? node50 : node33;
					assign node33 = (inp[5]) ? node43 : node34;
						assign node34 = (inp[0]) ? 2'b10 : node35;
							assign node35 = (inp[1]) ? node39 : node36;
								assign node36 = (inp[4]) ? 2'b11 : 2'b10;
								assign node39 = (inp[4]) ? 2'b10 : 2'b11;
						assign node43 = (inp[4]) ? node45 : 2'b10;
							assign node45 = (inp[1]) ? 2'b11 : node46;
								assign node46 = (inp[0]) ? 2'b11 : 2'b10;
					assign node50 = (inp[5]) ? node56 : node51;
						assign node51 = (inp[4]) ? 2'b11 : node52;
							assign node52 = (inp[0]) ? 2'b11 : 2'b10;
						assign node56 = (inp[0]) ? 2'b10 : node57;
							assign node57 = (inp[4]) ? 2'b10 : 2'b11;
			assign node61 = (inp[0]) ? node85 : node62;
				assign node62 = (inp[7]) ? node78 : node63;
					assign node63 = (inp[3]) ? node71 : node64;
						assign node64 = (inp[1]) ? node68 : node65;
							assign node65 = (inp[4]) ? 2'b11 : 2'b10;
							assign node68 = (inp[4]) ? 2'b10 : 2'b11;
						assign node71 = (inp[1]) ? node75 : node72;
							assign node72 = (inp[4]) ? 2'b11 : 2'b10;
							assign node75 = (inp[5]) ? 2'b11 : 2'b10;
					assign node78 = (inp[3]) ? node82 : node79;
						assign node79 = (inp[4]) ? 2'b01 : 2'b00;
						assign node82 = (inp[4]) ? 2'b00 : 2'b01;
				assign node85 = (inp[3]) ? node91 : node86;
					assign node86 = (inp[1]) ? 2'b01 : node87;
						assign node87 = (inp[7]) ? 2'b01 : 2'b00;
					assign node91 = (inp[7]) ? 2'b00 : node92;
						assign node92 = (inp[1]) ? 2'b00 : 2'b01;
		assign node96 = (inp[7]) ? node128 : node97;
			assign node97 = (inp[0]) ? node117 : node98;
				assign node98 = (inp[2]) ? node110 : node99;
					assign node99 = (inp[4]) ? node103 : node100;
						assign node100 = (inp[3]) ? 2'b11 : 2'b10;
						assign node103 = (inp[3]) ? node105 : 2'b11;
							assign node105 = (inp[1]) ? 2'b10 : node106;
								assign node106 = (inp[5]) ? 2'b11 : 2'b10;
					assign node110 = (inp[4]) ? node114 : node111;
						assign node111 = (inp[1]) ? 2'b11 : 2'b10;
						assign node114 = (inp[1]) ? 2'b10 : 2'b11;
				assign node117 = (inp[1]) ? node123 : node118;
					assign node118 = (inp[2]) ? 2'b01 : node119;
						assign node119 = (inp[5]) ? 2'b01 : 2'b00;
					assign node123 = (inp[2]) ? 2'b00 : node124;
						assign node124 = (inp[5]) ? 2'b00 : 2'b01;
			assign node128 = (inp[2]) ? node148 : node129;
				assign node129 = (inp[5]) ? node141 : node130;
					assign node130 = (inp[0]) ? 2'b01 : node131;
						assign node131 = (inp[3]) ? node137 : node132;
							assign node132 = (inp[1]) ? 2'b01 : node133;
								assign node133 = (inp[4]) ? 2'b00 : 2'b01;
							assign node137 = (inp[4]) ? 2'b01 : 2'b00;
					assign node141 = (inp[0]) ? 2'b00 : node142;
						assign node142 = (inp[1]) ? node144 : 2'b00;
							assign node144 = (inp[4]) ? 2'b00 : 2'b01;
				assign node148 = (inp[0]) ? 2'b00 : node149;
					assign node149 = (inp[4]) ? 2'b00 : 2'b01;

endmodule