module dtc_split125_bm60 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node6;
	wire [3-1:0] node8;
	wire [3-1:0] node10;
	wire [3-1:0] node13;
	wire [3-1:0] node14;
	wire [3-1:0] node16;
	wire [3-1:0] node20;
	wire [3-1:0] node21;
	wire [3-1:0] node22;
	wire [3-1:0] node23;
	wire [3-1:0] node25;
	wire [3-1:0] node30;
	wire [3-1:0] node32;
	wire [3-1:0] node33;
	wire [3-1:0] node37;
	wire [3-1:0] node38;
	wire [3-1:0] node39;
	wire [3-1:0] node41;
	wire [3-1:0] node43;
	wire [3-1:0] node46;
	wire [3-1:0] node48;
	wire [3-1:0] node51;
	wire [3-1:0] node52;
	wire [3-1:0] node54;
	wire [3-1:0] node56;
	wire [3-1:0] node58;
	wire [3-1:0] node62;
	wire [3-1:0] node63;
	wire [3-1:0] node64;
	wire [3-1:0] node65;
	wire [3-1:0] node67;
	wire [3-1:0] node70;
	wire [3-1:0] node71;
	wire [3-1:0] node72;
	wire [3-1:0] node77;
	wire [3-1:0] node78;
	wire [3-1:0] node79;
	wire [3-1:0] node81;
	wire [3-1:0] node85;
	wire [3-1:0] node87;
	wire [3-1:0] node88;
	wire [3-1:0] node90;
	wire [3-1:0] node94;
	wire [3-1:0] node95;
	wire [3-1:0] node96;
	wire [3-1:0] node98;
	wire [3-1:0] node100;
	wire [3-1:0] node103;
	wire [3-1:0] node105;
	wire [3-1:0] node106;
	wire [3-1:0] node108;
	wire [3-1:0] node109;
	wire [3-1:0] node114;
	wire [3-1:0] node115;
	wire [3-1:0] node116;
	wire [3-1:0] node118;
	wire [3-1:0] node120;
	wire [3-1:0] node123;
	wire [3-1:0] node125;
	wire [3-1:0] node128;
	wire [3-1:0] node129;
	wire [3-1:0] node132;
	wire [3-1:0] node133;
	wire [3-1:0] node136;
	wire [3-1:0] node137;
	wire [3-1:0] node138;
	wire [3-1:0] node142;
	wire [3-1:0] node144;

	assign outp = (inp[2]) ? node62 : node1;
		assign node1 = (inp[3]) ? node37 : node2;
			assign node2 = (inp[5]) ? node20 : node3;
				assign node3 = (inp[10]) ? node13 : node4;
					assign node4 = (inp[4]) ? node6 : 3'b111;
						assign node6 = (inp[9]) ? node8 : 3'b110;
							assign node8 = (inp[8]) ? node10 : 3'b110;
								assign node10 = (inp[7]) ? 3'b111 : 3'b110;
					assign node13 = (inp[9]) ? 3'b110 : node14;
						assign node14 = (inp[4]) ? node16 : 3'b110;
							assign node16 = (inp[7]) ? 3'b110 : 3'b111;
				assign node20 = (inp[10]) ? node30 : node21;
					assign node21 = (inp[4]) ? 3'b111 : node22;
						assign node22 = (inp[0]) ? 3'b111 : node23;
							assign node23 = (inp[7]) ? node25 : 3'b111;
								assign node25 = (inp[6]) ? 3'b110 : 3'b111;
					assign node30 = (inp[9]) ? node32 : 3'b110;
						assign node32 = (inp[4]) ? 3'b011 : node33;
							assign node33 = (inp[0]) ? 3'b110 : 3'b111;
			assign node37 = (inp[4]) ? node51 : node38;
				assign node38 = (inp[10]) ? node46 : node39;
					assign node39 = (inp[9]) ? node41 : 3'b111;
						assign node41 = (inp[5]) ? node43 : 3'b111;
							assign node43 = (inp[7]) ? 3'b110 : 3'b111;
					assign node46 = (inp[5]) ? node48 : 3'b110;
						assign node48 = (inp[9]) ? 3'b011 : 3'b110;
				assign node51 = (inp[5]) ? 3'b010 : node52;
					assign node52 = (inp[7]) ? node54 : 3'b011;
						assign node54 = (inp[9]) ? node56 : 3'b011;
							assign node56 = (inp[0]) ? node58 : 3'b010;
								assign node58 = (inp[10]) ? 3'b011 : 3'b010;
		assign node62 = (inp[4]) ? node94 : node63;
			assign node63 = (inp[10]) ? node77 : node64;
				assign node64 = (inp[5]) ? node70 : node65;
					assign node65 = (inp[9]) ? node67 : 3'b011;
						assign node67 = (inp[3]) ? 3'b010 : 3'b011;
					assign node70 = (inp[7]) ? 3'b010 : node71;
						assign node71 = (inp[3]) ? 3'b010 : node72;
							assign node72 = (inp[9]) ? 3'b010 : 3'b011;
				assign node77 = (inp[3]) ? node85 : node78;
					assign node78 = (inp[5]) ? 3'b011 : node79;
						assign node79 = (inp[9]) ? node81 : 3'b010;
							assign node81 = (inp[11]) ? 3'b011 : 3'b010;
					assign node85 = (inp[5]) ? node87 : 3'b111;
						assign node87 = (inp[9]) ? 3'b110 : node88;
							assign node88 = (inp[0]) ? node90 : 3'b111;
								assign node90 = (inp[1]) ? 3'b111 : 3'b110;
			assign node94 = (inp[3]) ? node114 : node95;
				assign node95 = (inp[5]) ? node103 : node96;
					assign node96 = (inp[9]) ? node98 : 3'b101;
						assign node98 = (inp[10]) ? node100 : 3'b101;
							assign node100 = (inp[7]) ? 3'b100 : 3'b101;
					assign node103 = (inp[9]) ? node105 : 3'b100;
						assign node105 = (inp[10]) ? 3'b001 : node106;
							assign node106 = (inp[1]) ? node108 : 3'b101;
								assign node108 = (inp[0]) ? 3'b100 : node109;
									assign node109 = (inp[8]) ? 3'b100 : 3'b100;
				assign node114 = (inp[10]) ? node128 : node115;
					assign node115 = (inp[9]) ? node123 : node116;
						assign node116 = (inp[6]) ? node118 : 3'b001;
							assign node118 = (inp[7]) ? node120 : 3'b001;
								assign node120 = (inp[0]) ? 3'b001 : 3'b000;
						assign node123 = (inp[8]) ? node125 : 3'b000;
							assign node125 = (inp[5]) ? 3'b000 : 3'b001;
					assign node128 = (inp[5]) ? node132 : node129;
						assign node129 = (inp[9]) ? 3'b100 : 3'b101;
						assign node132 = (inp[9]) ? node136 : node133;
							assign node133 = (inp[7]) ? 3'b100 : 3'b101;
							assign node136 = (inp[7]) ? node142 : node137;
								assign node137 = (inp[0]) ? 3'b001 : node138;
									assign node138 = (inp[8]) ? 3'b000 : 3'b001;
								assign node142 = (inp[8]) ? node144 : 3'b000;
									assign node144 = (inp[6]) ? 3'b000 : 3'b001;

endmodule