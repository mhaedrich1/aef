module dtc_split25_bm50 (
	input  wire [8-1:0] inp,
	output wire [2-1:0] outp
);

	wire [2-1:0] node1;
	wire [2-1:0] node2;
	wire [2-1:0] node3;
	wire [2-1:0] node4;
	wire [2-1:0] node6;
	wire [2-1:0] node8;
	wire [2-1:0] node11;
	wire [2-1:0] node14;
	wire [2-1:0] node15;
	wire [2-1:0] node16;
	wire [2-1:0] node21;
	wire [2-1:0] node22;
	wire [2-1:0] node23;
	wire [2-1:0] node26;
	wire [2-1:0] node29;
	wire [2-1:0] node32;
	wire [2-1:0] node33;
	wire [2-1:0] node34;
	wire [2-1:0] node35;
	wire [2-1:0] node38;
	wire [2-1:0] node39;
	wire [2-1:0] node43;
	wire [2-1:0] node44;
	wire [2-1:0] node45;
	wire [2-1:0] node46;
	wire [2-1:0] node51;
	wire [2-1:0] node52;
	wire [2-1:0] node55;
	wire [2-1:0] node56;
	wire [2-1:0] node60;
	wire [2-1:0] node61;
	wire [2-1:0] node62;
	wire [2-1:0] node63;
	wire [2-1:0] node64;
	wire [2-1:0] node65;
	wire [2-1:0] node70;
	wire [2-1:0] node72;
	wire [2-1:0] node75;
	wire [2-1:0] node77;
	wire [2-1:0] node80;
	wire [2-1:0] node81;

	assign outp = (inp[5]) ? node32 : node1;
		assign node1 = (inp[0]) ? node21 : node2;
			assign node2 = (inp[7]) ? node14 : node3;
				assign node3 = (inp[2]) ? node11 : node4;
					assign node4 = (inp[3]) ? node6 : 2'b10;
						assign node6 = (inp[4]) ? node8 : 2'b11;
							assign node8 = (inp[1]) ? 2'b11 : 2'b01;
					assign node11 = (inp[1]) ? 2'b00 : 2'b10;
				assign node14 = (inp[1]) ? 2'b11 : node15;
					assign node15 = (inp[6]) ? 2'b01 : node16;
						assign node16 = (inp[2]) ? 2'b01 : 2'b10;
			assign node21 = (inp[7]) ? node29 : node22;
				assign node22 = (inp[6]) ? node26 : node23;
					assign node23 = (inp[3]) ? 2'b01 : 2'b10;
					assign node26 = (inp[4]) ? 2'b01 : 2'b11;
				assign node29 = (inp[6]) ? 2'b00 : 2'b01;
		assign node32 = (inp[1]) ? node60 : node33;
			assign node33 = (inp[4]) ? node43 : node34;
				assign node34 = (inp[3]) ? node38 : node35;
					assign node35 = (inp[6]) ? 2'b00 : 2'b01;
					assign node38 = (inp[0]) ? 2'b11 : node39;
						assign node39 = (inp[7]) ? 2'b11 : 2'b00;
				assign node43 = (inp[3]) ? node51 : node44;
					assign node44 = (inp[2]) ? 2'b11 : node45;
						assign node45 = (inp[6]) ? 2'b11 : node46;
							assign node46 = (inp[0]) ? 2'b11 : 2'b00;
					assign node51 = (inp[2]) ? node55 : node52;
						assign node52 = (inp[6]) ? 2'b11 : 2'b10;
						assign node55 = (inp[7]) ? 2'b10 : node56;
							assign node56 = (inp[0]) ? 2'b11 : 2'b10;
			assign node60 = (inp[3]) ? node80 : node61;
				assign node61 = (inp[4]) ? node75 : node62;
					assign node62 = (inp[2]) ? node70 : node63;
						assign node63 = (inp[7]) ? 2'b11 : node64;
							assign node64 = (inp[0]) ? 2'b11 : node65;
								assign node65 = (inp[6]) ? 2'b10 : 2'b11;
						assign node70 = (inp[7]) ? node72 : 2'b10;
							assign node72 = (inp[0]) ? 2'b10 : 2'b11;
					assign node75 = (inp[0]) ? node77 : 2'b10;
						assign node77 = (inp[2]) ? 2'b01 : 2'b00;
				assign node80 = (inp[0]) ? 2'b00 : node81;
					assign node81 = (inp[7]) ? 2'b01 : 2'b11;

endmodule