module dtc_split875_bm63 (
	input  wire [16-1:0] inp,
	output wire [4-1:0] outp
);

	wire [4-1:0] node1;
	wire [4-1:0] node2;
	wire [4-1:0] node3;
	wire [4-1:0] node4;
	wire [4-1:0] node5;
	wire [4-1:0] node6;
	wire [4-1:0] node7;
	wire [4-1:0] node8;
	wire [4-1:0] node9;
	wire [4-1:0] node10;
	wire [4-1:0] node11;
	wire [4-1:0] node12;
	wire [4-1:0] node13;
	wire [4-1:0] node15;
	wire [4-1:0] node17;
	wire [4-1:0] node20;
	wire [4-1:0] node21;
	wire [4-1:0] node25;
	wire [4-1:0] node26;
	wire [4-1:0] node27;
	wire [4-1:0] node30;
	wire [4-1:0] node32;
	wire [4-1:0] node35;
	wire [4-1:0] node36;
	wire [4-1:0] node37;
	wire [4-1:0] node41;
	wire [4-1:0] node42;
	wire [4-1:0] node45;
	wire [4-1:0] node48;
	wire [4-1:0] node49;
	wire [4-1:0] node50;
	wire [4-1:0] node53;
	wire [4-1:0] node54;
	wire [4-1:0] node55;
	wire [4-1:0] node58;
	wire [4-1:0] node61;
	wire [4-1:0] node62;
	wire [4-1:0] node65;
	wire [4-1:0] node68;
	wire [4-1:0] node69;
	wire [4-1:0] node70;
	wire [4-1:0] node71;
	wire [4-1:0] node74;
	wire [4-1:0] node77;
	wire [4-1:0] node78;
	wire [4-1:0] node81;
	wire [4-1:0] node84;
	wire [4-1:0] node85;
	wire [4-1:0] node86;
	wire [4-1:0] node90;
	wire [4-1:0] node91;
	wire [4-1:0] node95;
	wire [4-1:0] node96;
	wire [4-1:0] node97;
	wire [4-1:0] node98;
	wire [4-1:0] node101;
	wire [4-1:0] node102;
	wire [4-1:0] node104;
	wire [4-1:0] node107;
	wire [4-1:0] node108;
	wire [4-1:0] node111;
	wire [4-1:0] node114;
	wire [4-1:0] node115;
	wire [4-1:0] node116;
	wire [4-1:0] node119;
	wire [4-1:0] node121;
	wire [4-1:0] node124;
	wire [4-1:0] node125;
	wire [4-1:0] node126;
	wire [4-1:0] node129;
	wire [4-1:0] node132;
	wire [4-1:0] node133;
	wire [4-1:0] node136;
	wire [4-1:0] node139;
	wire [4-1:0] node140;
	wire [4-1:0] node141;
	wire [4-1:0] node142;
	wire [4-1:0] node144;
	wire [4-1:0] node147;
	wire [4-1:0] node148;
	wire [4-1:0] node152;
	wire [4-1:0] node154;
	wire [4-1:0] node156;
	wire [4-1:0] node159;
	wire [4-1:0] node160;
	wire [4-1:0] node161;
	wire [4-1:0] node163;
	wire [4-1:0] node166;
	wire [4-1:0] node167;
	wire [4-1:0] node171;
	wire [4-1:0] node172;
	wire [4-1:0] node174;
	wire [4-1:0] node177;
	wire [4-1:0] node179;
	wire [4-1:0] node182;
	wire [4-1:0] node183;
	wire [4-1:0] node184;
	wire [4-1:0] node185;
	wire [4-1:0] node188;
	wire [4-1:0] node189;
	wire [4-1:0] node190;
	wire [4-1:0] node193;
	wire [4-1:0] node195;
	wire [4-1:0] node198;
	wire [4-1:0] node199;
	wire [4-1:0] node200;
	wire [4-1:0] node204;
	wire [4-1:0] node207;
	wire [4-1:0] node208;
	wire [4-1:0] node209;
	wire [4-1:0] node210;
	wire [4-1:0] node213;
	wire [4-1:0] node214;
	wire [4-1:0] node217;
	wire [4-1:0] node220;
	wire [4-1:0] node221;
	wire [4-1:0] node222;
	wire [4-1:0] node226;
	wire [4-1:0] node227;
	wire [4-1:0] node231;
	wire [4-1:0] node232;
	wire [4-1:0] node233;
	wire [4-1:0] node234;
	wire [4-1:0] node238;
	wire [4-1:0] node241;
	wire [4-1:0] node242;
	wire [4-1:0] node245;
	wire [4-1:0] node248;
	wire [4-1:0] node249;
	wire [4-1:0] node250;
	wire [4-1:0] node251;
	wire [4-1:0] node252;
	wire [4-1:0] node255;
	wire [4-1:0] node258;
	wire [4-1:0] node259;
	wire [4-1:0] node261;
	wire [4-1:0] node264;
	wire [4-1:0] node267;
	wire [4-1:0] node268;
	wire [4-1:0] node269;
	wire [4-1:0] node270;
	wire [4-1:0] node274;
	wire [4-1:0] node276;
	wire [4-1:0] node279;
	wire [4-1:0] node280;
	wire [4-1:0] node283;
	wire [4-1:0] node286;
	wire [4-1:0] node287;
	wire [4-1:0] node288;
	wire [4-1:0] node289;
	wire [4-1:0] node292;
	wire [4-1:0] node295;
	wire [4-1:0] node296;
	wire [4-1:0] node299;
	wire [4-1:0] node300;
	wire [4-1:0] node303;
	wire [4-1:0] node306;
	wire [4-1:0] node307;
	wire [4-1:0] node308;
	wire [4-1:0] node309;
	wire [4-1:0] node313;
	wire [4-1:0] node316;
	wire [4-1:0] node317;
	wire [4-1:0] node319;
	wire [4-1:0] node322;
	wire [4-1:0] node324;
	wire [4-1:0] node327;
	wire [4-1:0] node328;
	wire [4-1:0] node329;
	wire [4-1:0] node330;
	wire [4-1:0] node331;
	wire [4-1:0] node334;
	wire [4-1:0] node335;
	wire [4-1:0] node336;
	wire [4-1:0] node339;
	wire [4-1:0] node340;
	wire [4-1:0] node343;
	wire [4-1:0] node346;
	wire [4-1:0] node347;
	wire [4-1:0] node350;
	wire [4-1:0] node353;
	wire [4-1:0] node354;
	wire [4-1:0] node355;
	wire [4-1:0] node356;
	wire [4-1:0] node359;
	wire [4-1:0] node360;
	wire [4-1:0] node363;
	wire [4-1:0] node366;
	wire [4-1:0] node368;
	wire [4-1:0] node370;
	wire [4-1:0] node373;
	wire [4-1:0] node374;
	wire [4-1:0] node375;
	wire [4-1:0] node378;
	wire [4-1:0] node381;
	wire [4-1:0] node382;
	wire [4-1:0] node385;
	wire [4-1:0] node386;
	wire [4-1:0] node390;
	wire [4-1:0] node391;
	wire [4-1:0] node392;
	wire [4-1:0] node393;
	wire [4-1:0] node394;
	wire [4-1:0] node397;
	wire [4-1:0] node400;
	wire [4-1:0] node401;
	wire [4-1:0] node404;
	wire [4-1:0] node405;
	wire [4-1:0] node408;
	wire [4-1:0] node411;
	wire [4-1:0] node412;
	wire [4-1:0] node413;
	wire [4-1:0] node414;
	wire [4-1:0] node417;
	wire [4-1:0] node420;
	wire [4-1:0] node421;
	wire [4-1:0] node424;
	wire [4-1:0] node427;
	wire [4-1:0] node428;
	wire [4-1:0] node430;
	wire [4-1:0] node433;
	wire [4-1:0] node434;
	wire [4-1:0] node437;
	wire [4-1:0] node440;
	wire [4-1:0] node441;
	wire [4-1:0] node442;
	wire [4-1:0] node443;
	wire [4-1:0] node445;
	wire [4-1:0] node448;
	wire [4-1:0] node450;
	wire [4-1:0] node453;
	wire [4-1:0] node454;
	wire [4-1:0] node456;
	wire [4-1:0] node459;
	wire [4-1:0] node462;
	wire [4-1:0] node463;
	wire [4-1:0] node464;
	wire [4-1:0] node465;
	wire [4-1:0] node470;
	wire [4-1:0] node471;
	wire [4-1:0] node473;
	wire [4-1:0] node476;
	wire [4-1:0] node477;
	wire [4-1:0] node480;
	wire [4-1:0] node483;
	wire [4-1:0] node484;
	wire [4-1:0] node485;
	wire [4-1:0] node486;
	wire [4-1:0] node487;
	wire [4-1:0] node488;
	wire [4-1:0] node492;
	wire [4-1:0] node493;
	wire [4-1:0] node496;
	wire [4-1:0] node499;
	wire [4-1:0] node500;
	wire [4-1:0] node501;
	wire [4-1:0] node502;
	wire [4-1:0] node505;
	wire [4-1:0] node508;
	wire [4-1:0] node509;
	wire [4-1:0] node512;
	wire [4-1:0] node515;
	wire [4-1:0] node516;
	wire [4-1:0] node519;
	wire [4-1:0] node521;
	wire [4-1:0] node524;
	wire [4-1:0] node525;
	wire [4-1:0] node526;
	wire [4-1:0] node527;
	wire [4-1:0] node528;
	wire [4-1:0] node531;
	wire [4-1:0] node534;
	wire [4-1:0] node535;
	wire [4-1:0] node538;
	wire [4-1:0] node541;
	wire [4-1:0] node543;
	wire [4-1:0] node546;
	wire [4-1:0] node547;
	wire [4-1:0] node548;
	wire [4-1:0] node550;
	wire [4-1:0] node553;
	wire [4-1:0] node556;
	wire [4-1:0] node557;
	wire [4-1:0] node559;
	wire [4-1:0] node562;
	wire [4-1:0] node565;
	wire [4-1:0] node566;
	wire [4-1:0] node567;
	wire [4-1:0] node568;
	wire [4-1:0] node569;
	wire [4-1:0] node570;
	wire [4-1:0] node575;
	wire [4-1:0] node576;
	wire [4-1:0] node577;
	wire [4-1:0] node581;
	wire [4-1:0] node584;
	wire [4-1:0] node585;
	wire [4-1:0] node586;
	wire [4-1:0] node588;
	wire [4-1:0] node591;
	wire [4-1:0] node593;
	wire [4-1:0] node596;
	wire [4-1:0] node597;
	wire [4-1:0] node598;
	wire [4-1:0] node601;
	wire [4-1:0] node604;
	wire [4-1:0] node606;
	wire [4-1:0] node609;
	wire [4-1:0] node610;
	wire [4-1:0] node611;
	wire [4-1:0] node612;
	wire [4-1:0] node613;
	wire [4-1:0] node617;
	wire [4-1:0] node619;
	wire [4-1:0] node622;
	wire [4-1:0] node623;
	wire [4-1:0] node624;
	wire [4-1:0] node627;
	wire [4-1:0] node630;
	wire [4-1:0] node633;
	wire [4-1:0] node634;
	wire [4-1:0] node635;
	wire [4-1:0] node636;
	wire [4-1:0] node639;
	wire [4-1:0] node642;
	wire [4-1:0] node645;
	wire [4-1:0] node646;
	wire [4-1:0] node649;
	wire [4-1:0] node652;
	wire [4-1:0] node653;
	wire [4-1:0] node654;
	wire [4-1:0] node655;
	wire [4-1:0] node656;
	wire [4-1:0] node657;
	wire [4-1:0] node659;
	wire [4-1:0] node660;
	wire [4-1:0] node662;
	wire [4-1:0] node665;
	wire [4-1:0] node667;
	wire [4-1:0] node670;
	wire [4-1:0] node672;
	wire [4-1:0] node673;
	wire [4-1:0] node675;
	wire [4-1:0] node678;
	wire [4-1:0] node679;
	wire [4-1:0] node683;
	wire [4-1:0] node684;
	wire [4-1:0] node685;
	wire [4-1:0] node686;
	wire [4-1:0] node689;
	wire [4-1:0] node692;
	wire [4-1:0] node693;
	wire [4-1:0] node696;
	wire [4-1:0] node697;
	wire [4-1:0] node701;
	wire [4-1:0] node702;
	wire [4-1:0] node703;
	wire [4-1:0] node704;
	wire [4-1:0] node707;
	wire [4-1:0] node710;
	wire [4-1:0] node711;
	wire [4-1:0] node715;
	wire [4-1:0] node716;
	wire [4-1:0] node717;
	wire [4-1:0] node720;
	wire [4-1:0] node723;
	wire [4-1:0] node724;
	wire [4-1:0] node728;
	wire [4-1:0] node729;
	wire [4-1:0] node730;
	wire [4-1:0] node731;
	wire [4-1:0] node732;
	wire [4-1:0] node735;
	wire [4-1:0] node737;
	wire [4-1:0] node740;
	wire [4-1:0] node741;
	wire [4-1:0] node744;
	wire [4-1:0] node745;
	wire [4-1:0] node749;
	wire [4-1:0] node750;
	wire [4-1:0] node752;
	wire [4-1:0] node753;
	wire [4-1:0] node757;
	wire [4-1:0] node758;
	wire [4-1:0] node759;
	wire [4-1:0] node762;
	wire [4-1:0] node765;
	wire [4-1:0] node766;
	wire [4-1:0] node769;
	wire [4-1:0] node772;
	wire [4-1:0] node773;
	wire [4-1:0] node774;
	wire [4-1:0] node775;
	wire [4-1:0] node777;
	wire [4-1:0] node780;
	wire [4-1:0] node781;
	wire [4-1:0] node785;
	wire [4-1:0] node786;
	wire [4-1:0] node788;
	wire [4-1:0] node791;
	wire [4-1:0] node793;
	wire [4-1:0] node796;
	wire [4-1:0] node797;
	wire [4-1:0] node799;
	wire [4-1:0] node800;
	wire [4-1:0] node804;
	wire [4-1:0] node805;
	wire [4-1:0] node807;
	wire [4-1:0] node810;
	wire [4-1:0] node811;
	wire [4-1:0] node815;
	wire [4-1:0] node816;
	wire [4-1:0] node817;
	wire [4-1:0] node818;
	wire [4-1:0] node819;
	wire [4-1:0] node821;
	wire [4-1:0] node823;
	wire [4-1:0] node826;
	wire [4-1:0] node828;
	wire [4-1:0] node831;
	wire [4-1:0] node832;
	wire [4-1:0] node834;
	wire [4-1:0] node835;
	wire [4-1:0] node839;
	wire [4-1:0] node841;
	wire [4-1:0] node842;
	wire [4-1:0] node846;
	wire [4-1:0] node847;
	wire [4-1:0] node848;
	wire [4-1:0] node850;
	wire [4-1:0] node852;
	wire [4-1:0] node855;
	wire [4-1:0] node856;
	wire [4-1:0] node857;
	wire [4-1:0] node860;
	wire [4-1:0] node863;
	wire [4-1:0] node866;
	wire [4-1:0] node867;
	wire [4-1:0] node868;
	wire [4-1:0] node871;
	wire [4-1:0] node874;
	wire [4-1:0] node875;
	wire [4-1:0] node878;
	wire [4-1:0] node879;
	wire [4-1:0] node883;
	wire [4-1:0] node884;
	wire [4-1:0] node885;
	wire [4-1:0] node886;
	wire [4-1:0] node887;
	wire [4-1:0] node888;
	wire [4-1:0] node892;
	wire [4-1:0] node895;
	wire [4-1:0] node896;
	wire [4-1:0] node897;
	wire [4-1:0] node901;
	wire [4-1:0] node902;
	wire [4-1:0] node906;
	wire [4-1:0] node907;
	wire [4-1:0] node908;
	wire [4-1:0] node911;
	wire [4-1:0] node914;
	wire [4-1:0] node915;
	wire [4-1:0] node918;
	wire [4-1:0] node919;
	wire [4-1:0] node923;
	wire [4-1:0] node924;
	wire [4-1:0] node925;
	wire [4-1:0] node926;
	wire [4-1:0] node928;
	wire [4-1:0] node931;
	wire [4-1:0] node932;
	wire [4-1:0] node936;
	wire [4-1:0] node937;
	wire [4-1:0] node938;
	wire [4-1:0] node942;
	wire [4-1:0] node945;
	wire [4-1:0] node946;
	wire [4-1:0] node948;
	wire [4-1:0] node951;
	wire [4-1:0] node952;
	wire [4-1:0] node955;
	wire [4-1:0] node957;
	wire [4-1:0] node960;
	wire [4-1:0] node961;
	wire [4-1:0] node962;
	wire [4-1:0] node963;
	wire [4-1:0] node964;
	wire [4-1:0] node966;
	wire [4-1:0] node968;
	wire [4-1:0] node971;
	wire [4-1:0] node972;
	wire [4-1:0] node973;
	wire [4-1:0] node974;
	wire [4-1:0] node977;
	wire [4-1:0] node981;
	wire [4-1:0] node982;
	wire [4-1:0] node983;
	wire [4-1:0] node987;
	wire [4-1:0] node988;
	wire [4-1:0] node992;
	wire [4-1:0] node993;
	wire [4-1:0] node995;
	wire [4-1:0] node996;
	wire [4-1:0] node997;
	wire [4-1:0] node1001;
	wire [4-1:0] node1004;
	wire [4-1:0] node1005;
	wire [4-1:0] node1006;
	wire [4-1:0] node1007;
	wire [4-1:0] node1011;
	wire [4-1:0] node1013;
	wire [4-1:0] node1016;
	wire [4-1:0] node1017;
	wire [4-1:0] node1020;
	wire [4-1:0] node1022;
	wire [4-1:0] node1025;
	wire [4-1:0] node1026;
	wire [4-1:0] node1027;
	wire [4-1:0] node1028;
	wire [4-1:0] node1029;
	wire [4-1:0] node1031;
	wire [4-1:0] node1034;
	wire [4-1:0] node1037;
	wire [4-1:0] node1038;
	wire [4-1:0] node1040;
	wire [4-1:0] node1043;
	wire [4-1:0] node1046;
	wire [4-1:0] node1047;
	wire [4-1:0] node1048;
	wire [4-1:0] node1051;
	wire [4-1:0] node1054;
	wire [4-1:0] node1055;
	wire [4-1:0] node1058;
	wire [4-1:0] node1061;
	wire [4-1:0] node1062;
	wire [4-1:0] node1063;
	wire [4-1:0] node1064;
	wire [4-1:0] node1065;
	wire [4-1:0] node1069;
	wire [4-1:0] node1071;
	wire [4-1:0] node1074;
	wire [4-1:0] node1075;
	wire [4-1:0] node1076;
	wire [4-1:0] node1080;
	wire [4-1:0] node1083;
	wire [4-1:0] node1084;
	wire [4-1:0] node1085;
	wire [4-1:0] node1087;
	wire [4-1:0] node1090;
	wire [4-1:0] node1093;
	wire [4-1:0] node1094;
	wire [4-1:0] node1096;
	wire [4-1:0] node1099;
	wire [4-1:0] node1100;
	wire [4-1:0] node1104;
	wire [4-1:0] node1105;
	wire [4-1:0] node1106;
	wire [4-1:0] node1107;
	wire [4-1:0] node1108;
	wire [4-1:0] node1109;
	wire [4-1:0] node1111;
	wire [4-1:0] node1114;
	wire [4-1:0] node1117;
	wire [4-1:0] node1118;
	wire [4-1:0] node1121;
	wire [4-1:0] node1123;
	wire [4-1:0] node1126;
	wire [4-1:0] node1127;
	wire [4-1:0] node1128;
	wire [4-1:0] node1129;
	wire [4-1:0] node1132;
	wire [4-1:0] node1135;
	wire [4-1:0] node1136;
	wire [4-1:0] node1140;
	wire [4-1:0] node1141;
	wire [4-1:0] node1142;
	wire [4-1:0] node1146;
	wire [4-1:0] node1148;
	wire [4-1:0] node1151;
	wire [4-1:0] node1152;
	wire [4-1:0] node1153;
	wire [4-1:0] node1154;
	wire [4-1:0] node1157;
	wire [4-1:0] node1158;
	wire [4-1:0] node1162;
	wire [4-1:0] node1163;
	wire [4-1:0] node1166;
	wire [4-1:0] node1168;
	wire [4-1:0] node1171;
	wire [4-1:0] node1172;
	wire [4-1:0] node1173;
	wire [4-1:0] node1176;
	wire [4-1:0] node1179;
	wire [4-1:0] node1180;
	wire [4-1:0] node1182;
	wire [4-1:0] node1185;
	wire [4-1:0] node1186;
	wire [4-1:0] node1190;
	wire [4-1:0] node1191;
	wire [4-1:0] node1192;
	wire [4-1:0] node1193;
	wire [4-1:0] node1194;
	wire [4-1:0] node1195;
	wire [4-1:0] node1199;
	wire [4-1:0] node1200;
	wire [4-1:0] node1204;
	wire [4-1:0] node1205;
	wire [4-1:0] node1206;
	wire [4-1:0] node1210;
	wire [4-1:0] node1213;
	wire [4-1:0] node1214;
	wire [4-1:0] node1215;
	wire [4-1:0] node1217;
	wire [4-1:0] node1220;
	wire [4-1:0] node1221;
	wire [4-1:0] node1224;
	wire [4-1:0] node1227;
	wire [4-1:0] node1228;
	wire [4-1:0] node1229;
	wire [4-1:0] node1232;
	wire [4-1:0] node1235;
	wire [4-1:0] node1238;
	wire [4-1:0] node1239;
	wire [4-1:0] node1240;
	wire [4-1:0] node1241;
	wire [4-1:0] node1243;
	wire [4-1:0] node1246;
	wire [4-1:0] node1248;
	wire [4-1:0] node1251;
	wire [4-1:0] node1252;
	wire [4-1:0] node1254;
	wire [4-1:0] node1257;
	wire [4-1:0] node1260;
	wire [4-1:0] node1261;
	wire [4-1:0] node1262;
	wire [4-1:0] node1263;
	wire [4-1:0] node1266;
	wire [4-1:0] node1269;
	wire [4-1:0] node1272;
	wire [4-1:0] node1273;
	wire [4-1:0] node1276;
	wire [4-1:0] node1279;
	wire [4-1:0] node1280;
	wire [4-1:0] node1281;
	wire [4-1:0] node1282;
	wire [4-1:0] node1283;
	wire [4-1:0] node1284;
	wire [4-1:0] node1285;
	wire [4-1:0] node1288;
	wire [4-1:0] node1289;
	wire [4-1:0] node1290;
	wire [4-1:0] node1293;
	wire [4-1:0] node1296;
	wire [4-1:0] node1297;
	wire [4-1:0] node1298;
	wire [4-1:0] node1302;
	wire [4-1:0] node1303;
	wire [4-1:0] node1306;
	wire [4-1:0] node1309;
	wire [4-1:0] node1310;
	wire [4-1:0] node1311;
	wire [4-1:0] node1312;
	wire [4-1:0] node1313;
	wire [4-1:0] node1316;
	wire [4-1:0] node1320;
	wire [4-1:0] node1321;
	wire [4-1:0] node1323;
	wire [4-1:0] node1326;
	wire [4-1:0] node1327;
	wire [4-1:0] node1331;
	wire [4-1:0] node1332;
	wire [4-1:0] node1333;
	wire [4-1:0] node1335;
	wire [4-1:0] node1338;
	wire [4-1:0] node1339;
	wire [4-1:0] node1343;
	wire [4-1:0] node1344;
	wire [4-1:0] node1347;
	wire [4-1:0] node1348;
	wire [4-1:0] node1352;
	wire [4-1:0] node1353;
	wire [4-1:0] node1354;
	wire [4-1:0] node1355;
	wire [4-1:0] node1358;
	wire [4-1:0] node1359;
	wire [4-1:0] node1360;
	wire [4-1:0] node1363;
	wire [4-1:0] node1366;
	wire [4-1:0] node1368;
	wire [4-1:0] node1371;
	wire [4-1:0] node1372;
	wire [4-1:0] node1373;
	wire [4-1:0] node1376;
	wire [4-1:0] node1377;
	wire [4-1:0] node1381;
	wire [4-1:0] node1382;
	wire [4-1:0] node1383;
	wire [4-1:0] node1387;
	wire [4-1:0] node1388;
	wire [4-1:0] node1392;
	wire [4-1:0] node1393;
	wire [4-1:0] node1394;
	wire [4-1:0] node1395;
	wire [4-1:0] node1397;
	wire [4-1:0] node1401;
	wire [4-1:0] node1402;
	wire [4-1:0] node1404;
	wire [4-1:0] node1407;
	wire [4-1:0] node1409;
	wire [4-1:0] node1412;
	wire [4-1:0] node1413;
	wire [4-1:0] node1414;
	wire [4-1:0] node1416;
	wire [4-1:0] node1419;
	wire [4-1:0] node1421;
	wire [4-1:0] node1424;
	wire [4-1:0] node1425;
	wire [4-1:0] node1428;
	wire [4-1:0] node1429;
	wire [4-1:0] node1432;
	wire [4-1:0] node1435;
	wire [4-1:0] node1436;
	wire [4-1:0] node1437;
	wire [4-1:0] node1438;
	wire [4-1:0] node1440;
	wire [4-1:0] node1441;
	wire [4-1:0] node1443;
	wire [4-1:0] node1446;
	wire [4-1:0] node1449;
	wire [4-1:0] node1450;
	wire [4-1:0] node1451;
	wire [4-1:0] node1452;
	wire [4-1:0] node1455;
	wire [4-1:0] node1458;
	wire [4-1:0] node1459;
	wire [4-1:0] node1463;
	wire [4-1:0] node1464;
	wire [4-1:0] node1466;
	wire [4-1:0] node1469;
	wire [4-1:0] node1472;
	wire [4-1:0] node1473;
	wire [4-1:0] node1474;
	wire [4-1:0] node1476;
	wire [4-1:0] node1477;
	wire [4-1:0] node1481;
	wire [4-1:0] node1483;
	wire [4-1:0] node1484;
	wire [4-1:0] node1488;
	wire [4-1:0] node1489;
	wire [4-1:0] node1490;
	wire [4-1:0] node1491;
	wire [4-1:0] node1495;
	wire [4-1:0] node1498;
	wire [4-1:0] node1499;
	wire [4-1:0] node1501;
	wire [4-1:0] node1504;
	wire [4-1:0] node1506;
	wire [4-1:0] node1509;
	wire [4-1:0] node1510;
	wire [4-1:0] node1511;
	wire [4-1:0] node1512;
	wire [4-1:0] node1513;
	wire [4-1:0] node1516;
	wire [4-1:0] node1519;
	wire [4-1:0] node1520;
	wire [4-1:0] node1523;
	wire [4-1:0] node1524;
	wire [4-1:0] node1528;
	wire [4-1:0] node1529;
	wire [4-1:0] node1530;
	wire [4-1:0] node1531;
	wire [4-1:0] node1535;
	wire [4-1:0] node1538;
	wire [4-1:0] node1539;
	wire [4-1:0] node1542;
	wire [4-1:0] node1545;
	wire [4-1:0] node1546;
	wire [4-1:0] node1547;
	wire [4-1:0] node1548;
	wire [4-1:0] node1549;
	wire [4-1:0] node1553;
	wire [4-1:0] node1556;
	wire [4-1:0] node1557;
	wire [4-1:0] node1558;
	wire [4-1:0] node1562;
	wire [4-1:0] node1565;
	wire [4-1:0] node1566;
	wire [4-1:0] node1567;
	wire [4-1:0] node1569;
	wire [4-1:0] node1572;
	wire [4-1:0] node1575;
	wire [4-1:0] node1576;
	wire [4-1:0] node1578;
	wire [4-1:0] node1581;
	wire [4-1:0] node1582;
	wire [4-1:0] node1585;
	wire [4-1:0] node1588;
	wire [4-1:0] node1589;
	wire [4-1:0] node1590;
	wire [4-1:0] node1591;
	wire [4-1:0] node1592;
	wire [4-1:0] node1595;
	wire [4-1:0] node1596;
	wire [4-1:0] node1597;
	wire [4-1:0] node1601;
	wire [4-1:0] node1602;
	wire [4-1:0] node1603;
	wire [4-1:0] node1607;
	wire [4-1:0] node1610;
	wire [4-1:0] node1611;
	wire [4-1:0] node1612;
	wire [4-1:0] node1613;
	wire [4-1:0] node1615;
	wire [4-1:0] node1619;
	wire [4-1:0] node1620;
	wire [4-1:0] node1623;
	wire [4-1:0] node1626;
	wire [4-1:0] node1627;
	wire [4-1:0] node1628;
	wire [4-1:0] node1629;
	wire [4-1:0] node1634;
	wire [4-1:0] node1635;
	wire [4-1:0] node1636;
	wire [4-1:0] node1640;
	wire [4-1:0] node1642;
	wire [4-1:0] node1645;
	wire [4-1:0] node1646;
	wire [4-1:0] node1647;
	wire [4-1:0] node1648;
	wire [4-1:0] node1650;
	wire [4-1:0] node1653;
	wire [4-1:0] node1655;
	wire [4-1:0] node1656;
	wire [4-1:0] node1660;
	wire [4-1:0] node1661;
	wire [4-1:0] node1662;
	wire [4-1:0] node1663;
	wire [4-1:0] node1667;
	wire [4-1:0] node1668;
	wire [4-1:0] node1672;
	wire [4-1:0] node1673;
	wire [4-1:0] node1675;
	wire [4-1:0] node1678;
	wire [4-1:0] node1679;
	wire [4-1:0] node1683;
	wire [4-1:0] node1684;
	wire [4-1:0] node1685;
	wire [4-1:0] node1686;
	wire [4-1:0] node1690;
	wire [4-1:0] node1691;
	wire [4-1:0] node1692;
	wire [4-1:0] node1696;
	wire [4-1:0] node1698;
	wire [4-1:0] node1701;
	wire [4-1:0] node1702;
	wire [4-1:0] node1703;
	wire [4-1:0] node1705;
	wire [4-1:0] node1708;
	wire [4-1:0] node1709;
	wire [4-1:0] node1712;
	wire [4-1:0] node1715;
	wire [4-1:0] node1717;
	wire [4-1:0] node1718;
	wire [4-1:0] node1721;
	wire [4-1:0] node1724;
	wire [4-1:0] node1725;
	wire [4-1:0] node1726;
	wire [4-1:0] node1727;
	wire [4-1:0] node1728;
	wire [4-1:0] node1729;
	wire [4-1:0] node1732;
	wire [4-1:0] node1733;
	wire [4-1:0] node1737;
	wire [4-1:0] node1738;
	wire [4-1:0] node1741;
	wire [4-1:0] node1742;
	wire [4-1:0] node1746;
	wire [4-1:0] node1747;
	wire [4-1:0] node1748;
	wire [4-1:0] node1749;
	wire [4-1:0] node1752;
	wire [4-1:0] node1755;
	wire [4-1:0] node1756;
	wire [4-1:0] node1760;
	wire [4-1:0] node1762;
	wire [4-1:0] node1763;
	wire [4-1:0] node1767;
	wire [4-1:0] node1768;
	wire [4-1:0] node1769;
	wire [4-1:0] node1770;
	wire [4-1:0] node1773;
	wire [4-1:0] node1774;
	wire [4-1:0] node1778;
	wire [4-1:0] node1779;
	wire [4-1:0] node1782;
	wire [4-1:0] node1784;
	wire [4-1:0] node1787;
	wire [4-1:0] node1788;
	wire [4-1:0] node1789;
	wire [4-1:0] node1792;
	wire [4-1:0] node1795;
	wire [4-1:0] node1796;
	wire [4-1:0] node1798;
	wire [4-1:0] node1801;
	wire [4-1:0] node1802;
	wire [4-1:0] node1806;
	wire [4-1:0] node1807;
	wire [4-1:0] node1808;
	wire [4-1:0] node1809;
	wire [4-1:0] node1810;
	wire [4-1:0] node1814;
	wire [4-1:0] node1815;
	wire [4-1:0] node1816;
	wire [4-1:0] node1820;
	wire [4-1:0] node1821;
	wire [4-1:0] node1824;
	wire [4-1:0] node1827;
	wire [4-1:0] node1828;
	wire [4-1:0] node1829;
	wire [4-1:0] node1830;
	wire [4-1:0] node1834;
	wire [4-1:0] node1837;
	wire [4-1:0] node1838;
	wire [4-1:0] node1839;
	wire [4-1:0] node1842;
	wire [4-1:0] node1845;
	wire [4-1:0] node1846;
	wire [4-1:0] node1849;
	wire [4-1:0] node1852;
	wire [4-1:0] node1853;
	wire [4-1:0] node1854;
	wire [4-1:0] node1856;
	wire [4-1:0] node1858;
	wire [4-1:0] node1861;
	wire [4-1:0] node1862;
	wire [4-1:0] node1863;
	wire [4-1:0] node1866;
	wire [4-1:0] node1869;
	wire [4-1:0] node1872;
	wire [4-1:0] node1873;
	wire [4-1:0] node1874;
	wire [4-1:0] node1875;
	wire [4-1:0] node1878;
	wire [4-1:0] node1881;
	wire [4-1:0] node1884;
	wire [4-1:0] node1885;
	wire [4-1:0] node1888;
	wire [4-1:0] node1891;
	wire [4-1:0] node1892;
	wire [4-1:0] node1893;
	wire [4-1:0] node1894;
	wire [4-1:0] node1895;
	wire [4-1:0] node1896;
	wire [4-1:0] node1899;
	wire [4-1:0] node1900;
	wire [4-1:0] node1902;
	wire [4-1:0] node1905;
	wire [4-1:0] node1906;
	wire [4-1:0] node1909;
	wire [4-1:0] node1910;
	wire [4-1:0] node1914;
	wire [4-1:0] node1915;
	wire [4-1:0] node1916;
	wire [4-1:0] node1919;
	wire [4-1:0] node1921;
	wire [4-1:0] node1924;
	wire [4-1:0] node1925;
	wire [4-1:0] node1926;
	wire [4-1:0] node1928;
	wire [4-1:0] node1931;
	wire [4-1:0] node1932;
	wire [4-1:0] node1936;
	wire [4-1:0] node1937;
	wire [4-1:0] node1938;
	wire [4-1:0] node1942;
	wire [4-1:0] node1943;
	wire [4-1:0] node1947;
	wire [4-1:0] node1948;
	wire [4-1:0] node1949;
	wire [4-1:0] node1950;
	wire [4-1:0] node1953;
	wire [4-1:0] node1954;
	wire [4-1:0] node1957;
	wire [4-1:0] node1958;
	wire [4-1:0] node1961;
	wire [4-1:0] node1964;
	wire [4-1:0] node1965;
	wire [4-1:0] node1966;
	wire [4-1:0] node1969;
	wire [4-1:0] node1972;
	wire [4-1:0] node1973;
	wire [4-1:0] node1974;
	wire [4-1:0] node1977;
	wire [4-1:0] node1980;
	wire [4-1:0] node1981;
	wire [4-1:0] node1985;
	wire [4-1:0] node1986;
	wire [4-1:0] node1987;
	wire [4-1:0] node1988;
	wire [4-1:0] node1989;
	wire [4-1:0] node1992;
	wire [4-1:0] node1995;
	wire [4-1:0] node1996;
	wire [4-1:0] node1999;
	wire [4-1:0] node2002;
	wire [4-1:0] node2003;
	wire [4-1:0] node2004;
	wire [4-1:0] node2008;
	wire [4-1:0] node2009;
	wire [4-1:0] node2013;
	wire [4-1:0] node2014;
	wire [4-1:0] node2015;
	wire [4-1:0] node2016;
	wire [4-1:0] node2020;
	wire [4-1:0] node2023;
	wire [4-1:0] node2024;
	wire [4-1:0] node2026;
	wire [4-1:0] node2029;
	wire [4-1:0] node2032;
	wire [4-1:0] node2033;
	wire [4-1:0] node2034;
	wire [4-1:0] node2035;
	wire [4-1:0] node2036;
	wire [4-1:0] node2039;
	wire [4-1:0] node2040;
	wire [4-1:0] node2043;
	wire [4-1:0] node2045;
	wire [4-1:0] node2048;
	wire [4-1:0] node2049;
	wire [4-1:0] node2052;
	wire [4-1:0] node2053;
	wire [4-1:0] node2056;
	wire [4-1:0] node2057;
	wire [4-1:0] node2060;
	wire [4-1:0] node2063;
	wire [4-1:0] node2064;
	wire [4-1:0] node2065;
	wire [4-1:0] node2066;
	wire [4-1:0] node2069;
	wire [4-1:0] node2071;
	wire [4-1:0] node2074;
	wire [4-1:0] node2075;
	wire [4-1:0] node2078;
	wire [4-1:0] node2079;
	wire [4-1:0] node2082;
	wire [4-1:0] node2085;
	wire [4-1:0] node2086;
	wire [4-1:0] node2087;
	wire [4-1:0] node2088;
	wire [4-1:0] node2091;
	wire [4-1:0] node2094;
	wire [4-1:0] node2095;
	wire [4-1:0] node2098;
	wire [4-1:0] node2101;
	wire [4-1:0] node2102;
	wire [4-1:0] node2105;
	wire [4-1:0] node2107;
	wire [4-1:0] node2110;
	wire [4-1:0] node2111;
	wire [4-1:0] node2112;
	wire [4-1:0] node2113;
	wire [4-1:0] node2114;
	wire [4-1:0] node2115;
	wire [4-1:0] node2118;
	wire [4-1:0] node2121;
	wire [4-1:0] node2122;
	wire [4-1:0] node2125;
	wire [4-1:0] node2128;
	wire [4-1:0] node2129;
	wire [4-1:0] node2132;
	wire [4-1:0] node2133;
	wire [4-1:0] node2136;
	wire [4-1:0] node2139;
	wire [4-1:0] node2140;
	wire [4-1:0] node2141;
	wire [4-1:0] node2142;
	wire [4-1:0] node2145;
	wire [4-1:0] node2148;
	wire [4-1:0] node2149;
	wire [4-1:0] node2152;
	wire [4-1:0] node2155;
	wire [4-1:0] node2156;
	wire [4-1:0] node2158;
	wire [4-1:0] node2161;
	wire [4-1:0] node2162;
	wire [4-1:0] node2165;
	wire [4-1:0] node2168;
	wire [4-1:0] node2169;
	wire [4-1:0] node2170;
	wire [4-1:0] node2171;
	wire [4-1:0] node2174;
	wire [4-1:0] node2175;
	wire [4-1:0] node2179;
	wire [4-1:0] node2180;
	wire [4-1:0] node2181;
	wire [4-1:0] node2185;
	wire [4-1:0] node2186;
	wire [4-1:0] node2189;
	wire [4-1:0] node2192;
	wire [4-1:0] node2193;
	wire [4-1:0] node2194;
	wire [4-1:0] node2195;
	wire [4-1:0] node2199;
	wire [4-1:0] node2202;
	wire [4-1:0] node2203;
	wire [4-1:0] node2206;
	wire [4-1:0] node2207;
	wire [4-1:0] node2211;
	wire [4-1:0] node2212;
	wire [4-1:0] node2213;
	wire [4-1:0] node2214;
	wire [4-1:0] node2215;
	wire [4-1:0] node2216;
	wire [4-1:0] node2217;
	wire [4-1:0] node2218;
	wire [4-1:0] node2221;
	wire [4-1:0] node2224;
	wire [4-1:0] node2225;
	wire [4-1:0] node2229;
	wire [4-1:0] node2230;
	wire [4-1:0] node2231;
	wire [4-1:0] node2234;
	wire [4-1:0] node2238;
	wire [4-1:0] node2239;
	wire [4-1:0] node2240;
	wire [4-1:0] node2242;
	wire [4-1:0] node2245;
	wire [4-1:0] node2246;
	wire [4-1:0] node2250;
	wire [4-1:0] node2251;
	wire [4-1:0] node2252;
	wire [4-1:0] node2255;
	wire [4-1:0] node2258;
	wire [4-1:0] node2259;
	wire [4-1:0] node2262;
	wire [4-1:0] node2265;
	wire [4-1:0] node2266;
	wire [4-1:0] node2267;
	wire [4-1:0] node2268;
	wire [4-1:0] node2271;
	wire [4-1:0] node2274;
	wire [4-1:0] node2275;
	wire [4-1:0] node2277;
	wire [4-1:0] node2280;
	wire [4-1:0] node2282;
	wire [4-1:0] node2285;
	wire [4-1:0] node2286;
	wire [4-1:0] node2287;
	wire [4-1:0] node2288;
	wire [4-1:0] node2292;
	wire [4-1:0] node2293;
	wire [4-1:0] node2297;
	wire [4-1:0] node2298;
	wire [4-1:0] node2301;
	wire [4-1:0] node2302;
	wire [4-1:0] node2305;
	wire [4-1:0] node2308;
	wire [4-1:0] node2309;
	wire [4-1:0] node2310;
	wire [4-1:0] node2311;
	wire [4-1:0] node2312;
	wire [4-1:0] node2314;
	wire [4-1:0] node2317;
	wire [4-1:0] node2318;
	wire [4-1:0] node2321;
	wire [4-1:0] node2324;
	wire [4-1:0] node2325;
	wire [4-1:0] node2327;
	wire [4-1:0] node2330;
	wire [4-1:0] node2331;
	wire [4-1:0] node2335;
	wire [4-1:0] node2336;
	wire [4-1:0] node2337;
	wire [4-1:0] node2338;
	wire [4-1:0] node2341;
	wire [4-1:0] node2344;
	wire [4-1:0] node2347;
	wire [4-1:0] node2348;
	wire [4-1:0] node2350;
	wire [4-1:0] node2353;
	wire [4-1:0] node2354;
	wire [4-1:0] node2357;
	wire [4-1:0] node2360;
	wire [4-1:0] node2361;
	wire [4-1:0] node2362;
	wire [4-1:0] node2363;
	wire [4-1:0] node2364;
	wire [4-1:0] node2367;
	wire [4-1:0] node2370;
	wire [4-1:0] node2372;
	wire [4-1:0] node2375;
	wire [4-1:0] node2376;
	wire [4-1:0] node2378;
	wire [4-1:0] node2381;
	wire [4-1:0] node2383;
	wire [4-1:0] node2386;
	wire [4-1:0] node2387;
	wire [4-1:0] node2388;
	wire [4-1:0] node2389;
	wire [4-1:0] node2393;
	wire [4-1:0] node2396;
	wire [4-1:0] node2397;
	wire [4-1:0] node2398;
	wire [4-1:0] node2401;
	wire [4-1:0] node2404;
	wire [4-1:0] node2405;
	wire [4-1:0] node2408;
	wire [4-1:0] node2411;
	wire [4-1:0] node2412;
	wire [4-1:0] node2413;
	wire [4-1:0] node2414;
	wire [4-1:0] node2415;
	wire [4-1:0] node2417;
	wire [4-1:0] node2418;
	wire [4-1:0] node2422;
	wire [4-1:0] node2423;
	wire [4-1:0] node2424;
	wire [4-1:0] node2427;
	wire [4-1:0] node2430;
	wire [4-1:0] node2433;
	wire [4-1:0] node2434;
	wire [4-1:0] node2436;
	wire [4-1:0] node2437;
	wire [4-1:0] node2441;
	wire [4-1:0] node2442;
	wire [4-1:0] node2444;
	wire [4-1:0] node2447;
	wire [4-1:0] node2448;
	wire [4-1:0] node2452;
	wire [4-1:0] node2453;
	wire [4-1:0] node2454;
	wire [4-1:0] node2455;
	wire [4-1:0] node2458;
	wire [4-1:0] node2459;
	wire [4-1:0] node2463;
	wire [4-1:0] node2464;
	wire [4-1:0] node2465;
	wire [4-1:0] node2469;
	wire [4-1:0] node2470;
	wire [4-1:0] node2474;
	wire [4-1:0] node2475;
	wire [4-1:0] node2476;
	wire [4-1:0] node2478;
	wire [4-1:0] node2481;
	wire [4-1:0] node2484;
	wire [4-1:0] node2485;
	wire [4-1:0] node2488;
	wire [4-1:0] node2490;
	wire [4-1:0] node2493;
	wire [4-1:0] node2494;
	wire [4-1:0] node2495;
	wire [4-1:0] node2496;
	wire [4-1:0] node2497;
	wire [4-1:0] node2499;
	wire [4-1:0] node2502;
	wire [4-1:0] node2503;
	wire [4-1:0] node2507;
	wire [4-1:0] node2508;
	wire [4-1:0] node2510;
	wire [4-1:0] node2513;
	wire [4-1:0] node2514;
	wire [4-1:0] node2518;
	wire [4-1:0] node2519;
	wire [4-1:0] node2520;
	wire [4-1:0] node2522;
	wire [4-1:0] node2525;
	wire [4-1:0] node2527;
	wire [4-1:0] node2530;
	wire [4-1:0] node2531;
	wire [4-1:0] node2533;
	wire [4-1:0] node2536;
	wire [4-1:0] node2537;
	wire [4-1:0] node2540;
	wire [4-1:0] node2543;
	wire [4-1:0] node2544;
	wire [4-1:0] node2545;
	wire [4-1:0] node2546;
	wire [4-1:0] node2547;
	wire [4-1:0] node2550;
	wire [4-1:0] node2553;
	wire [4-1:0] node2556;
	wire [4-1:0] node2557;
	wire [4-1:0] node2558;
	wire [4-1:0] node2562;
	wire [4-1:0] node2564;
	wire [4-1:0] node2567;
	wire [4-1:0] node2568;
	wire [4-1:0] node2569;
	wire [4-1:0] node2571;
	wire [4-1:0] node2574;
	wire [4-1:0] node2575;
	wire [4-1:0] node2579;
	wire [4-1:0] node2580;
	wire [4-1:0] node2581;
	wire [4-1:0] node2585;
	wire [4-1:0] node2588;
	wire [4-1:0] node2589;
	wire [4-1:0] node2590;
	wire [4-1:0] node2591;
	wire [4-1:0] node2592;
	wire [4-1:0] node2593;
	wire [4-1:0] node2594;
	wire [4-1:0] node2595;
	wire [4-1:0] node2596;
	wire [4-1:0] node2598;
	wire [4-1:0] node2599;
	wire [4-1:0] node2603;
	wire [4-1:0] node2605;
	wire [4-1:0] node2606;
	wire [4-1:0] node2609;
	wire [4-1:0] node2612;
	wire [4-1:0] node2613;
	wire [4-1:0] node2614;
	wire [4-1:0] node2616;
	wire [4-1:0] node2619;
	wire [4-1:0] node2620;
	wire [4-1:0] node2623;
	wire [4-1:0] node2626;
	wire [4-1:0] node2627;
	wire [4-1:0] node2628;
	wire [4-1:0] node2631;
	wire [4-1:0] node2634;
	wire [4-1:0] node2635;
	wire [4-1:0] node2639;
	wire [4-1:0] node2640;
	wire [4-1:0] node2641;
	wire [4-1:0] node2642;
	wire [4-1:0] node2645;
	wire [4-1:0] node2647;
	wire [4-1:0] node2650;
	wire [4-1:0] node2651;
	wire [4-1:0] node2654;
	wire [4-1:0] node2655;
	wire [4-1:0] node2658;
	wire [4-1:0] node2661;
	wire [4-1:0] node2662;
	wire [4-1:0] node2663;
	wire [4-1:0] node2666;
	wire [4-1:0] node2667;
	wire [4-1:0] node2671;
	wire [4-1:0] node2672;
	wire [4-1:0] node2675;
	wire [4-1:0] node2677;
	wire [4-1:0] node2680;
	wire [4-1:0] node2681;
	wire [4-1:0] node2682;
	wire [4-1:0] node2683;
	wire [4-1:0] node2684;
	wire [4-1:0] node2686;
	wire [4-1:0] node2689;
	wire [4-1:0] node2690;
	wire [4-1:0] node2694;
	wire [4-1:0] node2695;
	wire [4-1:0] node2698;
	wire [4-1:0] node2701;
	wire [4-1:0] node2702;
	wire [4-1:0] node2703;
	wire [4-1:0] node2704;
	wire [4-1:0] node2708;
	wire [4-1:0] node2709;
	wire [4-1:0] node2713;
	wire [4-1:0] node2714;
	wire [4-1:0] node2715;
	wire [4-1:0] node2718;
	wire [4-1:0] node2721;
	wire [4-1:0] node2723;
	wire [4-1:0] node2726;
	wire [4-1:0] node2727;
	wire [4-1:0] node2728;
	wire [4-1:0] node2729;
	wire [4-1:0] node2732;
	wire [4-1:0] node2733;
	wire [4-1:0] node2736;
	wire [4-1:0] node2739;
	wire [4-1:0] node2740;
	wire [4-1:0] node2741;
	wire [4-1:0] node2744;
	wire [4-1:0] node2747;
	wire [4-1:0] node2748;
	wire [4-1:0] node2751;
	wire [4-1:0] node2754;
	wire [4-1:0] node2755;
	wire [4-1:0] node2756;
	wire [4-1:0] node2758;
	wire [4-1:0] node2761;
	wire [4-1:0] node2763;
	wire [4-1:0] node2766;
	wire [4-1:0] node2767;
	wire [4-1:0] node2769;
	wire [4-1:0] node2772;
	wire [4-1:0] node2773;
	wire [4-1:0] node2776;
	wire [4-1:0] node2779;
	wire [4-1:0] node2780;
	wire [4-1:0] node2781;
	wire [4-1:0] node2782;
	wire [4-1:0] node2783;
	wire [4-1:0] node2785;
	wire [4-1:0] node2786;
	wire [4-1:0] node2790;
	wire [4-1:0] node2792;
	wire [4-1:0] node2795;
	wire [4-1:0] node2796;
	wire [4-1:0] node2797;
	wire [4-1:0] node2800;
	wire [4-1:0] node2801;
	wire [4-1:0] node2804;
	wire [4-1:0] node2807;
	wire [4-1:0] node2808;
	wire [4-1:0] node2810;
	wire [4-1:0] node2814;
	wire [4-1:0] node2815;
	wire [4-1:0] node2816;
	wire [4-1:0] node2818;
	wire [4-1:0] node2821;
	wire [4-1:0] node2823;
	wire [4-1:0] node2824;
	wire [4-1:0] node2828;
	wire [4-1:0] node2829;
	wire [4-1:0] node2830;
	wire [4-1:0] node2831;
	wire [4-1:0] node2834;
	wire [4-1:0] node2837;
	wire [4-1:0] node2839;
	wire [4-1:0] node2842;
	wire [4-1:0] node2843;
	wire [4-1:0] node2845;
	wire [4-1:0] node2848;
	wire [4-1:0] node2851;
	wire [4-1:0] node2852;
	wire [4-1:0] node2853;
	wire [4-1:0] node2854;
	wire [4-1:0] node2855;
	wire [4-1:0] node2857;
	wire [4-1:0] node2860;
	wire [4-1:0] node2861;
	wire [4-1:0] node2865;
	wire [4-1:0] node2866;
	wire [4-1:0] node2869;
	wire [4-1:0] node2870;
	wire [4-1:0] node2873;
	wire [4-1:0] node2876;
	wire [4-1:0] node2877;
	wire [4-1:0] node2878;
	wire [4-1:0] node2879;
	wire [4-1:0] node2882;
	wire [4-1:0] node2885;
	wire [4-1:0] node2886;
	wire [4-1:0] node2889;
	wire [4-1:0] node2892;
	wire [4-1:0] node2893;
	wire [4-1:0] node2896;
	wire [4-1:0] node2897;
	wire [4-1:0] node2901;
	wire [4-1:0] node2902;
	wire [4-1:0] node2903;
	wire [4-1:0] node2904;
	wire [4-1:0] node2907;
	wire [4-1:0] node2908;
	wire [4-1:0] node2911;
	wire [4-1:0] node2914;
	wire [4-1:0] node2915;
	wire [4-1:0] node2918;
	wire [4-1:0] node2919;
	wire [4-1:0] node2923;
	wire [4-1:0] node2924;
	wire [4-1:0] node2925;
	wire [4-1:0] node2927;
	wire [4-1:0] node2930;
	wire [4-1:0] node2933;
	wire [4-1:0] node2934;
	wire [4-1:0] node2935;
	wire [4-1:0] node2938;
	wire [4-1:0] node2941;
	wire [4-1:0] node2942;
	wire [4-1:0] node2946;
	wire [4-1:0] node2947;
	wire [4-1:0] node2948;
	wire [4-1:0] node2949;
	wire [4-1:0] node2950;
	wire [4-1:0] node2951;
	wire [4-1:0] node2952;
	wire [4-1:0] node2955;
	wire [4-1:0] node2958;
	wire [4-1:0] node2959;
	wire [4-1:0] node2962;
	wire [4-1:0] node2965;
	wire [4-1:0] node2966;
	wire [4-1:0] node2967;
	wire [4-1:0] node2970;
	wire [4-1:0] node2973;
	wire [4-1:0] node2974;
	wire [4-1:0] node2976;
	wire [4-1:0] node2979;
	wire [4-1:0] node2980;
	wire [4-1:0] node2983;
	wire [4-1:0] node2986;
	wire [4-1:0] node2987;
	wire [4-1:0] node2988;
	wire [4-1:0] node2989;
	wire [4-1:0] node2990;
	wire [4-1:0] node2993;
	wire [4-1:0] node2996;
	wire [4-1:0] node2997;
	wire [4-1:0] node3000;
	wire [4-1:0] node3003;
	wire [4-1:0] node3004;
	wire [4-1:0] node3005;
	wire [4-1:0] node3008;
	wire [4-1:0] node3011;
	wire [4-1:0] node3012;
	wire [4-1:0] node3015;
	wire [4-1:0] node3018;
	wire [4-1:0] node3019;
	wire [4-1:0] node3020;
	wire [4-1:0] node3023;
	wire [4-1:0] node3024;
	wire [4-1:0] node3027;
	wire [4-1:0] node3030;
	wire [4-1:0] node3031;
	wire [4-1:0] node3032;
	wire [4-1:0] node3036;
	wire [4-1:0] node3037;
	wire [4-1:0] node3040;
	wire [4-1:0] node3043;
	wire [4-1:0] node3044;
	wire [4-1:0] node3045;
	wire [4-1:0] node3046;
	wire [4-1:0] node3047;
	wire [4-1:0] node3049;
	wire [4-1:0] node3052;
	wire [4-1:0] node3054;
	wire [4-1:0] node3057;
	wire [4-1:0] node3058;
	wire [4-1:0] node3059;
	wire [4-1:0] node3062;
	wire [4-1:0] node3065;
	wire [4-1:0] node3066;
	wire [4-1:0] node3069;
	wire [4-1:0] node3072;
	wire [4-1:0] node3073;
	wire [4-1:0] node3074;
	wire [4-1:0] node3075;
	wire [4-1:0] node3078;
	wire [4-1:0] node3081;
	wire [4-1:0] node3082;
	wire [4-1:0] node3085;
	wire [4-1:0] node3088;
	wire [4-1:0] node3089;
	wire [4-1:0] node3092;
	wire [4-1:0] node3093;
	wire [4-1:0] node3097;
	wire [4-1:0] node3098;
	wire [4-1:0] node3099;
	wire [4-1:0] node3100;
	wire [4-1:0] node3101;
	wire [4-1:0] node3105;
	wire [4-1:0] node3106;
	wire [4-1:0] node3110;
	wire [4-1:0] node3111;
	wire [4-1:0] node3114;
	wire [4-1:0] node3115;
	wire [4-1:0] node3118;
	wire [4-1:0] node3121;
	wire [4-1:0] node3122;
	wire [4-1:0] node3123;
	wire [4-1:0] node3124;
	wire [4-1:0] node3127;
	wire [4-1:0] node3130;
	wire [4-1:0] node3131;
	wire [4-1:0] node3134;
	wire [4-1:0] node3137;
	wire [4-1:0] node3138;
	wire [4-1:0] node3139;
	wire [4-1:0] node3142;
	wire [4-1:0] node3145;
	wire [4-1:0] node3146;
	wire [4-1:0] node3149;
	wire [4-1:0] node3152;
	wire [4-1:0] node3153;
	wire [4-1:0] node3154;
	wire [4-1:0] node3155;
	wire [4-1:0] node3156;
	wire [4-1:0] node3157;
	wire [4-1:0] node3158;
	wire [4-1:0] node3161;
	wire [4-1:0] node3164;
	wire [4-1:0] node3165;
	wire [4-1:0] node3168;
	wire [4-1:0] node3171;
	wire [4-1:0] node3172;
	wire [4-1:0] node3176;
	wire [4-1:0] node3177;
	wire [4-1:0] node3178;
	wire [4-1:0] node3179;
	wire [4-1:0] node3182;
	wire [4-1:0] node3185;
	wire [4-1:0] node3186;
	wire [4-1:0] node3189;
	wire [4-1:0] node3192;
	wire [4-1:0] node3193;
	wire [4-1:0] node3194;
	wire [4-1:0] node3197;
	wire [4-1:0] node3200;
	wire [4-1:0] node3201;
	wire [4-1:0] node3204;
	wire [4-1:0] node3207;
	wire [4-1:0] node3208;
	wire [4-1:0] node3209;
	wire [4-1:0] node3210;
	wire [4-1:0] node3212;
	wire [4-1:0] node3215;
	wire [4-1:0] node3216;
	wire [4-1:0] node3220;
	wire [4-1:0] node3221;
	wire [4-1:0] node3223;
	wire [4-1:0] node3226;
	wire [4-1:0] node3228;
	wire [4-1:0] node3231;
	wire [4-1:0] node3232;
	wire [4-1:0] node3233;
	wire [4-1:0] node3235;
	wire [4-1:0] node3238;
	wire [4-1:0] node3241;
	wire [4-1:0] node3242;
	wire [4-1:0] node3243;
	wire [4-1:0] node3246;
	wire [4-1:0] node3249;
	wire [4-1:0] node3250;
	wire [4-1:0] node3253;
	wire [4-1:0] node3256;
	wire [4-1:0] node3257;
	wire [4-1:0] node3258;
	wire [4-1:0] node3259;
	wire [4-1:0] node3260;
	wire [4-1:0] node3262;
	wire [4-1:0] node3265;
	wire [4-1:0] node3266;
	wire [4-1:0] node3269;
	wire [4-1:0] node3272;
	wire [4-1:0] node3273;
	wire [4-1:0] node3276;
	wire [4-1:0] node3277;
	wire [4-1:0] node3280;
	wire [4-1:0] node3283;
	wire [4-1:0] node3284;
	wire [4-1:0] node3285;
	wire [4-1:0] node3288;
	wire [4-1:0] node3289;
	wire [4-1:0] node3292;
	wire [4-1:0] node3295;
	wire [4-1:0] node3296;
	wire [4-1:0] node3299;
	wire [4-1:0] node3300;
	wire [4-1:0] node3304;
	wire [4-1:0] node3305;
	wire [4-1:0] node3306;
	wire [4-1:0] node3307;
	wire [4-1:0] node3308;
	wire [4-1:0] node3311;
	wire [4-1:0] node3314;
	wire [4-1:0] node3315;
	wire [4-1:0] node3318;
	wire [4-1:0] node3321;
	wire [4-1:0] node3322;
	wire [4-1:0] node3323;
	wire [4-1:0] node3326;
	wire [4-1:0] node3329;
	wire [4-1:0] node3330;
	wire [4-1:0] node3334;
	wire [4-1:0] node3335;
	wire [4-1:0] node3336;
	wire [4-1:0] node3338;
	wire [4-1:0] node3341;
	wire [4-1:0] node3342;
	wire [4-1:0] node3345;
	wire [4-1:0] node3348;
	wire [4-1:0] node3349;
	wire [4-1:0] node3350;
	wire [4-1:0] node3354;
	wire [4-1:0] node3355;
	wire [4-1:0] node3358;
	wire [4-1:0] node3361;
	wire [4-1:0] node3362;
	wire [4-1:0] node3363;
	wire [4-1:0] node3364;
	wire [4-1:0] node3365;
	wire [4-1:0] node3366;
	wire [4-1:0] node3367;
	wire [4-1:0] node3368;
	wire [4-1:0] node3370;
	wire [4-1:0] node3373;
	wire [4-1:0] node3375;
	wire [4-1:0] node3378;
	wire [4-1:0] node3379;
	wire [4-1:0] node3380;
	wire [4-1:0] node3383;
	wire [4-1:0] node3386;
	wire [4-1:0] node3387;
	wire [4-1:0] node3391;
	wire [4-1:0] node3392;
	wire [4-1:0] node3393;
	wire [4-1:0] node3394;
	wire [4-1:0] node3397;
	wire [4-1:0] node3400;
	wire [4-1:0] node3403;
	wire [4-1:0] node3404;
	wire [4-1:0] node3406;
	wire [4-1:0] node3409;
	wire [4-1:0] node3410;
	wire [4-1:0] node3413;
	wire [4-1:0] node3416;
	wire [4-1:0] node3417;
	wire [4-1:0] node3418;
	wire [4-1:0] node3419;
	wire [4-1:0] node3422;
	wire [4-1:0] node3424;
	wire [4-1:0] node3427;
	wire [4-1:0] node3428;
	wire [4-1:0] node3429;
	wire [4-1:0] node3432;
	wire [4-1:0] node3435;
	wire [4-1:0] node3436;
	wire [4-1:0] node3439;
	wire [4-1:0] node3442;
	wire [4-1:0] node3443;
	wire [4-1:0] node3445;
	wire [4-1:0] node3446;
	wire [4-1:0] node3450;
	wire [4-1:0] node3451;
	wire [4-1:0] node3454;
	wire [4-1:0] node3455;
	wire [4-1:0] node3459;
	wire [4-1:0] node3460;
	wire [4-1:0] node3461;
	wire [4-1:0] node3462;
	wire [4-1:0] node3463;
	wire [4-1:0] node3465;
	wire [4-1:0] node3468;
	wire [4-1:0] node3469;
	wire [4-1:0] node3472;
	wire [4-1:0] node3475;
	wire [4-1:0] node3476;
	wire [4-1:0] node3478;
	wire [4-1:0] node3481;
	wire [4-1:0] node3482;
	wire [4-1:0] node3485;
	wire [4-1:0] node3488;
	wire [4-1:0] node3489;
	wire [4-1:0] node3490;
	wire [4-1:0] node3491;
	wire [4-1:0] node3495;
	wire [4-1:0] node3496;
	wire [4-1:0] node3499;
	wire [4-1:0] node3502;
	wire [4-1:0] node3503;
	wire [4-1:0] node3504;
	wire [4-1:0] node3508;
	wire [4-1:0] node3509;
	wire [4-1:0] node3512;
	wire [4-1:0] node3515;
	wire [4-1:0] node3516;
	wire [4-1:0] node3517;
	wire [4-1:0] node3518;
	wire [4-1:0] node3520;
	wire [4-1:0] node3523;
	wire [4-1:0] node3524;
	wire [4-1:0] node3528;
	wire [4-1:0] node3529;
	wire [4-1:0] node3532;
	wire [4-1:0] node3533;
	wire [4-1:0] node3537;
	wire [4-1:0] node3538;
	wire [4-1:0] node3539;
	wire [4-1:0] node3540;
	wire [4-1:0] node3543;
	wire [4-1:0] node3546;
	wire [4-1:0] node3547;
	wire [4-1:0] node3550;
	wire [4-1:0] node3553;
	wire [4-1:0] node3554;
	wire [4-1:0] node3555;
	wire [4-1:0] node3558;
	wire [4-1:0] node3561;
	wire [4-1:0] node3562;
	wire [4-1:0] node3565;
	wire [4-1:0] node3568;
	wire [4-1:0] node3569;
	wire [4-1:0] node3570;
	wire [4-1:0] node3571;
	wire [4-1:0] node3572;
	wire [4-1:0] node3573;
	wire [4-1:0] node3574;
	wire [4-1:0] node3578;
	wire [4-1:0] node3580;
	wire [4-1:0] node3583;
	wire [4-1:0] node3584;
	wire [4-1:0] node3587;
	wire [4-1:0] node3589;
	wire [4-1:0] node3592;
	wire [4-1:0] node3593;
	wire [4-1:0] node3594;
	wire [4-1:0] node3597;
	wire [4-1:0] node3598;
	wire [4-1:0] node3602;
	wire [4-1:0] node3603;
	wire [4-1:0] node3605;
	wire [4-1:0] node3608;
	wire [4-1:0] node3609;
	wire [4-1:0] node3613;
	wire [4-1:0] node3614;
	wire [4-1:0] node3615;
	wire [4-1:0] node3616;
	wire [4-1:0] node3617;
	wire [4-1:0] node3621;
	wire [4-1:0] node3622;
	wire [4-1:0] node3625;
	wire [4-1:0] node3628;
	wire [4-1:0] node3629;
	wire [4-1:0] node3631;
	wire [4-1:0] node3634;
	wire [4-1:0] node3636;
	wire [4-1:0] node3639;
	wire [4-1:0] node3640;
	wire [4-1:0] node3641;
	wire [4-1:0] node3643;
	wire [4-1:0] node3646;
	wire [4-1:0] node3648;
	wire [4-1:0] node3651;
	wire [4-1:0] node3652;
	wire [4-1:0] node3653;
	wire [4-1:0] node3657;
	wire [4-1:0] node3658;
	wire [4-1:0] node3662;
	wire [4-1:0] node3663;
	wire [4-1:0] node3664;
	wire [4-1:0] node3665;
	wire [4-1:0] node3666;
	wire [4-1:0] node3669;
	wire [4-1:0] node3671;
	wire [4-1:0] node3674;
	wire [4-1:0] node3675;
	wire [4-1:0] node3677;
	wire [4-1:0] node3680;
	wire [4-1:0] node3681;
	wire [4-1:0] node3685;
	wire [4-1:0] node3686;
	wire [4-1:0] node3688;
	wire [4-1:0] node3689;
	wire [4-1:0] node3692;
	wire [4-1:0] node3695;
	wire [4-1:0] node3696;
	wire [4-1:0] node3697;
	wire [4-1:0] node3700;
	wire [4-1:0] node3703;
	wire [4-1:0] node3704;
	wire [4-1:0] node3707;
	wire [4-1:0] node3710;
	wire [4-1:0] node3711;
	wire [4-1:0] node3712;
	wire [4-1:0] node3713;
	wire [4-1:0] node3714;
	wire [4-1:0] node3717;
	wire [4-1:0] node3720;
	wire [4-1:0] node3721;
	wire [4-1:0] node3724;
	wire [4-1:0] node3727;
	wire [4-1:0] node3728;
	wire [4-1:0] node3729;
	wire [4-1:0] node3732;
	wire [4-1:0] node3735;
	wire [4-1:0] node3738;
	wire [4-1:0] node3739;
	wire [4-1:0] node3740;
	wire [4-1:0] node3741;
	wire [4-1:0] node3745;
	wire [4-1:0] node3746;
	wire [4-1:0] node3749;
	wire [4-1:0] node3752;
	wire [4-1:0] node3753;
	wire [4-1:0] node3754;
	wire [4-1:0] node3758;
	wire [4-1:0] node3759;
	wire [4-1:0] node3762;
	wire [4-1:0] node3765;
	wire [4-1:0] node3766;
	wire [4-1:0] node3767;
	wire [4-1:0] node3768;
	wire [4-1:0] node3769;
	wire [4-1:0] node3770;
	wire [4-1:0] node3771;
	wire [4-1:0] node3773;
	wire [4-1:0] node3776;
	wire [4-1:0] node3778;
	wire [4-1:0] node3781;
	wire [4-1:0] node3782;
	wire [4-1:0] node3784;
	wire [4-1:0] node3787;
	wire [4-1:0] node3788;
	wire [4-1:0] node3792;
	wire [4-1:0] node3793;
	wire [4-1:0] node3794;
	wire [4-1:0] node3797;
	wire [4-1:0] node3799;
	wire [4-1:0] node3802;
	wire [4-1:0] node3803;
	wire [4-1:0] node3805;
	wire [4-1:0] node3808;
	wire [4-1:0] node3809;
	wire [4-1:0] node3813;
	wire [4-1:0] node3814;
	wire [4-1:0] node3815;
	wire [4-1:0] node3816;
	wire [4-1:0] node3819;
	wire [4-1:0] node3822;
	wire [4-1:0] node3823;
	wire [4-1:0] node3826;
	wire [4-1:0] node3827;
	wire [4-1:0] node3831;
	wire [4-1:0] node3832;
	wire [4-1:0] node3833;
	wire [4-1:0] node3834;
	wire [4-1:0] node3838;
	wire [4-1:0] node3839;
	wire [4-1:0] node3843;
	wire [4-1:0] node3846;
	wire [4-1:0] node3847;
	wire [4-1:0] node3848;
	wire [4-1:0] node3849;
	wire [4-1:0] node3850;
	wire [4-1:0] node3853;
	wire [4-1:0] node3855;
	wire [4-1:0] node3858;
	wire [4-1:0] node3859;
	wire [4-1:0] node3860;
	wire [4-1:0] node3863;
	wire [4-1:0] node3866;
	wire [4-1:0] node3867;
	wire [4-1:0] node3870;
	wire [4-1:0] node3873;
	wire [4-1:0] node3874;
	wire [4-1:0] node3875;
	wire [4-1:0] node3877;
	wire [4-1:0] node3880;
	wire [4-1:0] node3882;
	wire [4-1:0] node3885;
	wire [4-1:0] node3886;
	wire [4-1:0] node3889;
	wire [4-1:0] node3890;
	wire [4-1:0] node3894;
	wire [4-1:0] node3895;
	wire [4-1:0] node3896;
	wire [4-1:0] node3897;
	wire [4-1:0] node3898;
	wire [4-1:0] node3901;
	wire [4-1:0] node3904;
	wire [4-1:0] node3907;
	wire [4-1:0] node3909;
	wire [4-1:0] node3912;
	wire [4-1:0] node3913;
	wire [4-1:0] node3914;
	wire [4-1:0] node3916;
	wire [4-1:0] node3919;
	wire [4-1:0] node3920;
	wire [4-1:0] node3923;
	wire [4-1:0] node3926;
	wire [4-1:0] node3927;
	wire [4-1:0] node3928;
	wire [4-1:0] node3932;
	wire [4-1:0] node3935;
	wire [4-1:0] node3936;
	wire [4-1:0] node3937;
	wire [4-1:0] node3938;
	wire [4-1:0] node3939;
	wire [4-1:0] node3940;
	wire [4-1:0] node3941;
	wire [4-1:0] node3945;
	wire [4-1:0] node3946;
	wire [4-1:0] node3949;
	wire [4-1:0] node3952;
	wire [4-1:0] node3953;
	wire [4-1:0] node3955;
	wire [4-1:0] node3958;
	wire [4-1:0] node3960;
	wire [4-1:0] node3963;
	wire [4-1:0] node3964;
	wire [4-1:0] node3965;
	wire [4-1:0] node3966;
	wire [4-1:0] node3969;
	wire [4-1:0] node3972;
	wire [4-1:0] node3973;
	wire [4-1:0] node3976;
	wire [4-1:0] node3979;
	wire [4-1:0] node3980;
	wire [4-1:0] node3983;
	wire [4-1:0] node3984;
	wire [4-1:0] node3987;
	wire [4-1:0] node3990;
	wire [4-1:0] node3991;
	wire [4-1:0] node3992;
	wire [4-1:0] node3993;
	wire [4-1:0] node3995;
	wire [4-1:0] node3998;
	wire [4-1:0] node4001;
	wire [4-1:0] node4002;
	wire [4-1:0] node4003;
	wire [4-1:0] node4006;
	wire [4-1:0] node4009;
	wire [4-1:0] node4012;
	wire [4-1:0] node4013;
	wire [4-1:0] node4014;
	wire [4-1:0] node4015;
	wire [4-1:0] node4019;
	wire [4-1:0] node4020;
	wire [4-1:0] node4023;
	wire [4-1:0] node4026;
	wire [4-1:0] node4027;
	wire [4-1:0] node4028;
	wire [4-1:0] node4031;
	wire [4-1:0] node4034;
	wire [4-1:0] node4035;
	wire [4-1:0] node4038;
	wire [4-1:0] node4041;
	wire [4-1:0] node4042;
	wire [4-1:0] node4043;
	wire [4-1:0] node4044;
	wire [4-1:0] node4045;
	wire [4-1:0] node4047;
	wire [4-1:0] node4050;
	wire [4-1:0] node4052;
	wire [4-1:0] node4055;
	wire [4-1:0] node4056;
	wire [4-1:0] node4057;
	wire [4-1:0] node4061;
	wire [4-1:0] node4062;
	wire [4-1:0] node4065;
	wire [4-1:0] node4068;
	wire [4-1:0] node4069;
	wire [4-1:0] node4070;
	wire [4-1:0] node4071;
	wire [4-1:0] node4075;
	wire [4-1:0] node4077;
	wire [4-1:0] node4080;
	wire [4-1:0] node4081;
	wire [4-1:0] node4082;
	wire [4-1:0] node4085;
	wire [4-1:0] node4088;
	wire [4-1:0] node4089;
	wire [4-1:0] node4092;
	wire [4-1:0] node4095;
	wire [4-1:0] node4096;
	wire [4-1:0] node4097;
	wire [4-1:0] node4098;
	wire [4-1:0] node4100;
	wire [4-1:0] node4103;
	wire [4-1:0] node4105;
	wire [4-1:0] node4108;
	wire [4-1:0] node4109;
	wire [4-1:0] node4110;
	wire [4-1:0] node4113;
	wire [4-1:0] node4116;
	wire [4-1:0] node4119;
	wire [4-1:0] node4120;
	wire [4-1:0] node4121;
	wire [4-1:0] node4123;
	wire [4-1:0] node4126;
	wire [4-1:0] node4127;
	wire [4-1:0] node4131;
	wire [4-1:0] node4132;
	wire [4-1:0] node4134;
	wire [4-1:0] node4138;
	wire [4-1:0] node4139;
	wire [4-1:0] node4140;
	wire [4-1:0] node4141;
	wire [4-1:0] node4142;
	wire [4-1:0] node4143;
	wire [4-1:0] node4144;
	wire [4-1:0] node4145;
	wire [4-1:0] node4146;
	wire [4-1:0] node4149;
	wire [4-1:0] node4150;
	wire [4-1:0] node4153;
	wire [4-1:0] node4156;
	wire [4-1:0] node4157;
	wire [4-1:0] node4158;
	wire [4-1:0] node4161;
	wire [4-1:0] node4164;
	wire [4-1:0] node4165;
	wire [4-1:0] node4168;
	wire [4-1:0] node4171;
	wire [4-1:0] node4172;
	wire [4-1:0] node4173;
	wire [4-1:0] node4176;
	wire [4-1:0] node4177;
	wire [4-1:0] node4181;
	wire [4-1:0] node4182;
	wire [4-1:0] node4183;
	wire [4-1:0] node4186;
	wire [4-1:0] node4189;
	wire [4-1:0] node4190;
	wire [4-1:0] node4193;
	wire [4-1:0] node4196;
	wire [4-1:0] node4197;
	wire [4-1:0] node4198;
	wire [4-1:0] node4199;
	wire [4-1:0] node4202;
	wire [4-1:0] node4203;
	wire [4-1:0] node4206;
	wire [4-1:0] node4209;
	wire [4-1:0] node4210;
	wire [4-1:0] node4213;
	wire [4-1:0] node4214;
	wire [4-1:0] node4218;
	wire [4-1:0] node4219;
	wire [4-1:0] node4220;
	wire [4-1:0] node4221;
	wire [4-1:0] node4225;
	wire [4-1:0] node4226;
	wire [4-1:0] node4229;
	wire [4-1:0] node4232;
	wire [4-1:0] node4233;
	wire [4-1:0] node4235;
	wire [4-1:0] node4238;
	wire [4-1:0] node4239;
	wire [4-1:0] node4242;
	wire [4-1:0] node4245;
	wire [4-1:0] node4246;
	wire [4-1:0] node4247;
	wire [4-1:0] node4248;
	wire [4-1:0] node4249;
	wire [4-1:0] node4252;
	wire [4-1:0] node4253;
	wire [4-1:0] node4256;
	wire [4-1:0] node4259;
	wire [4-1:0] node4260;
	wire [4-1:0] node4261;
	wire [4-1:0] node4264;
	wire [4-1:0] node4267;
	wire [4-1:0] node4268;
	wire [4-1:0] node4271;
	wire [4-1:0] node4274;
	wire [4-1:0] node4275;
	wire [4-1:0] node4276;
	wire [4-1:0] node4279;
	wire [4-1:0] node4280;
	wire [4-1:0] node4283;
	wire [4-1:0] node4286;
	wire [4-1:0] node4287;
	wire [4-1:0] node4288;
	wire [4-1:0] node4291;
	wire [4-1:0] node4294;
	wire [4-1:0] node4296;
	wire [4-1:0] node4299;
	wire [4-1:0] node4300;
	wire [4-1:0] node4301;
	wire [4-1:0] node4302;
	wire [4-1:0] node4303;
	wire [4-1:0] node4306;
	wire [4-1:0] node4309;
	wire [4-1:0] node4310;
	wire [4-1:0] node4313;
	wire [4-1:0] node4316;
	wire [4-1:0] node4317;
	wire [4-1:0] node4318;
	wire [4-1:0] node4321;
	wire [4-1:0] node4324;
	wire [4-1:0] node4325;
	wire [4-1:0] node4328;
	wire [4-1:0] node4331;
	wire [4-1:0] node4332;
	wire [4-1:0] node4333;
	wire [4-1:0] node4335;
	wire [4-1:0] node4338;
	wire [4-1:0] node4340;
	wire [4-1:0] node4343;
	wire [4-1:0] node4344;
	wire [4-1:0] node4347;
	wire [4-1:0] node4348;
	wire [4-1:0] node4351;
	wire [4-1:0] node4354;
	wire [4-1:0] node4355;
	wire [4-1:0] node4356;
	wire [4-1:0] node4357;
	wire [4-1:0] node4358;
	wire [4-1:0] node4359;
	wire [4-1:0] node4362;
	wire [4-1:0] node4363;
	wire [4-1:0] node4366;
	wire [4-1:0] node4369;
	wire [4-1:0] node4370;
	wire [4-1:0] node4371;
	wire [4-1:0] node4374;
	wire [4-1:0] node4377;
	wire [4-1:0] node4379;
	wire [4-1:0] node4382;
	wire [4-1:0] node4383;
	wire [4-1:0] node4384;
	wire [4-1:0] node4387;
	wire [4-1:0] node4389;
	wire [4-1:0] node4392;
	wire [4-1:0] node4393;
	wire [4-1:0] node4394;
	wire [4-1:0] node4397;
	wire [4-1:0] node4400;
	wire [4-1:0] node4401;
	wire [4-1:0] node4405;
	wire [4-1:0] node4406;
	wire [4-1:0] node4407;
	wire [4-1:0] node4408;
	wire [4-1:0] node4411;
	wire [4-1:0] node4412;
	wire [4-1:0] node4415;
	wire [4-1:0] node4418;
	wire [4-1:0] node4419;
	wire [4-1:0] node4421;
	wire [4-1:0] node4424;
	wire [4-1:0] node4425;
	wire [4-1:0] node4428;
	wire [4-1:0] node4431;
	wire [4-1:0] node4432;
	wire [4-1:0] node4433;
	wire [4-1:0] node4434;
	wire [4-1:0] node4437;
	wire [4-1:0] node4440;
	wire [4-1:0] node4441;
	wire [4-1:0] node4444;
	wire [4-1:0] node4447;
	wire [4-1:0] node4448;
	wire [4-1:0] node4450;
	wire [4-1:0] node4453;
	wire [4-1:0] node4455;
	wire [4-1:0] node4458;
	wire [4-1:0] node4459;
	wire [4-1:0] node4460;
	wire [4-1:0] node4461;
	wire [4-1:0] node4462;
	wire [4-1:0] node4465;
	wire [4-1:0] node4467;
	wire [4-1:0] node4470;
	wire [4-1:0] node4471;
	wire [4-1:0] node4474;
	wire [4-1:0] node4477;
	wire [4-1:0] node4478;
	wire [4-1:0] node4479;
	wire [4-1:0] node4480;
	wire [4-1:0] node4484;
	wire [4-1:0] node4485;
	wire [4-1:0] node4488;
	wire [4-1:0] node4491;
	wire [4-1:0] node4492;
	wire [4-1:0] node4493;
	wire [4-1:0] node4496;
	wire [4-1:0] node4499;
	wire [4-1:0] node4501;
	wire [4-1:0] node4504;
	wire [4-1:0] node4505;
	wire [4-1:0] node4506;
	wire [4-1:0] node4507;
	wire [4-1:0] node4510;
	wire [4-1:0] node4511;
	wire [4-1:0] node4514;
	wire [4-1:0] node4517;
	wire [4-1:0] node4518;
	wire [4-1:0] node4521;
	wire [4-1:0] node4523;
	wire [4-1:0] node4526;
	wire [4-1:0] node4527;
	wire [4-1:0] node4528;
	wire [4-1:0] node4530;
	wire [4-1:0] node4533;
	wire [4-1:0] node4534;
	wire [4-1:0] node4537;
	wire [4-1:0] node4540;
	wire [4-1:0] node4541;
	wire [4-1:0] node4542;
	wire [4-1:0] node4545;
	wire [4-1:0] node4548;
	wire [4-1:0] node4550;
	wire [4-1:0] node4553;
	wire [4-1:0] node4554;
	wire [4-1:0] node4555;
	wire [4-1:0] node4556;
	wire [4-1:0] node4557;
	wire [4-1:0] node4558;
	wire [4-1:0] node4559;
	wire [4-1:0] node4560;
	wire [4-1:0] node4564;
	wire [4-1:0] node4567;
	wire [4-1:0] node4568;
	wire [4-1:0] node4570;
	wire [4-1:0] node4573;
	wire [4-1:0] node4575;
	wire [4-1:0] node4578;
	wire [4-1:0] node4579;
	wire [4-1:0] node4580;
	wire [4-1:0] node4581;
	wire [4-1:0] node4585;
	wire [4-1:0] node4586;
	wire [4-1:0] node4589;
	wire [4-1:0] node4592;
	wire [4-1:0] node4593;
	wire [4-1:0] node4595;
	wire [4-1:0] node4598;
	wire [4-1:0] node4601;
	wire [4-1:0] node4602;
	wire [4-1:0] node4603;
	wire [4-1:0] node4605;
	wire [4-1:0] node4608;
	wire [4-1:0] node4609;
	wire [4-1:0] node4611;
	wire [4-1:0] node4614;
	wire [4-1:0] node4615;
	wire [4-1:0] node4619;
	wire [4-1:0] node4620;
	wire [4-1:0] node4621;
	wire [4-1:0] node4624;
	wire [4-1:0] node4625;
	wire [4-1:0] node4629;
	wire [4-1:0] node4630;
	wire [4-1:0] node4631;
	wire [4-1:0] node4635;
	wire [4-1:0] node4637;
	wire [4-1:0] node4640;
	wire [4-1:0] node4641;
	wire [4-1:0] node4642;
	wire [4-1:0] node4643;
	wire [4-1:0] node4644;
	wire [4-1:0] node4645;
	wire [4-1:0] node4648;
	wire [4-1:0] node4651;
	wire [4-1:0] node4652;
	wire [4-1:0] node4655;
	wire [4-1:0] node4658;
	wire [4-1:0] node4659;
	wire [4-1:0] node4661;
	wire [4-1:0] node4664;
	wire [4-1:0] node4667;
	wire [4-1:0] node4668;
	wire [4-1:0] node4670;
	wire [4-1:0] node4671;
	wire [4-1:0] node4675;
	wire [4-1:0] node4676;
	wire [4-1:0] node4678;
	wire [4-1:0] node4682;
	wire [4-1:0] node4683;
	wire [4-1:0] node4684;
	wire [4-1:0] node4685;
	wire [4-1:0] node4687;
	wire [4-1:0] node4690;
	wire [4-1:0] node4692;
	wire [4-1:0] node4695;
	wire [4-1:0] node4697;
	wire [4-1:0] node4698;
	wire [4-1:0] node4702;
	wire [4-1:0] node4703;
	wire [4-1:0] node4704;
	wire [4-1:0] node4706;
	wire [4-1:0] node4709;
	wire [4-1:0] node4710;
	wire [4-1:0] node4713;
	wire [4-1:0] node4716;
	wire [4-1:0] node4717;
	wire [4-1:0] node4720;
	wire [4-1:0] node4723;
	wire [4-1:0] node4724;
	wire [4-1:0] node4725;
	wire [4-1:0] node4726;
	wire [4-1:0] node4727;
	wire [4-1:0] node4728;
	wire [4-1:0] node4729;
	wire [4-1:0] node4732;
	wire [4-1:0] node4735;
	wire [4-1:0] node4736;
	wire [4-1:0] node4739;
	wire [4-1:0] node4742;
	wire [4-1:0] node4743;
	wire [4-1:0] node4745;
	wire [4-1:0] node4748;
	wire [4-1:0] node4751;
	wire [4-1:0] node4752;
	wire [4-1:0] node4753;
	wire [4-1:0] node4754;
	wire [4-1:0] node4758;
	wire [4-1:0] node4760;
	wire [4-1:0] node4763;
	wire [4-1:0] node4765;
	wire [4-1:0] node4768;
	wire [4-1:0] node4769;
	wire [4-1:0] node4770;
	wire [4-1:0] node4771;
	wire [4-1:0] node4772;
	wire [4-1:0] node4776;
	wire [4-1:0] node4777;
	wire [4-1:0] node4780;
	wire [4-1:0] node4783;
	wire [4-1:0] node4784;
	wire [4-1:0] node4786;
	wire [4-1:0] node4789;
	wire [4-1:0] node4790;
	wire [4-1:0] node4794;
	wire [4-1:0] node4795;
	wire [4-1:0] node4796;
	wire [4-1:0] node4798;
	wire [4-1:0] node4801;
	wire [4-1:0] node4804;
	wire [4-1:0] node4805;
	wire [4-1:0] node4807;
	wire [4-1:0] node4810;
	wire [4-1:0] node4811;
	wire [4-1:0] node4815;
	wire [4-1:0] node4816;
	wire [4-1:0] node4817;
	wire [4-1:0] node4818;
	wire [4-1:0] node4819;
	wire [4-1:0] node4820;
	wire [4-1:0] node4824;
	wire [4-1:0] node4827;
	wire [4-1:0] node4828;
	wire [4-1:0] node4829;
	wire [4-1:0] node4832;
	wire [4-1:0] node4835;
	wire [4-1:0] node4837;
	wire [4-1:0] node4840;
	wire [4-1:0] node4841;
	wire [4-1:0] node4842;
	wire [4-1:0] node4844;
	wire [4-1:0] node4847;
	wire [4-1:0] node4850;
	wire [4-1:0] node4851;
	wire [4-1:0] node4852;
	wire [4-1:0] node4856;
	wire [4-1:0] node4859;
	wire [4-1:0] node4860;
	wire [4-1:0] node4861;
	wire [4-1:0] node4862;
	wire [4-1:0] node4864;
	wire [4-1:0] node4867;
	wire [4-1:0] node4868;
	wire [4-1:0] node4872;
	wire [4-1:0] node4873;
	wire [4-1:0] node4874;
	wire [4-1:0] node4878;
	wire [4-1:0] node4879;
	wire [4-1:0] node4883;
	wire [4-1:0] node4884;
	wire [4-1:0] node4885;
	wire [4-1:0] node4887;
	wire [4-1:0] node4890;
	wire [4-1:0] node4891;
	wire [4-1:0] node4895;
	wire [4-1:0] node4896;
	wire [4-1:0] node4897;
	wire [4-1:0] node4900;
	wire [4-1:0] node4903;
	wire [4-1:0] node4904;
	wire [4-1:0] node4907;
	wire [4-1:0] node4910;
	wire [4-1:0] node4911;
	wire [4-1:0] node4912;
	wire [4-1:0] node4913;
	wire [4-1:0] node4914;
	wire [4-1:0] node4915;
	wire [4-1:0] node4916;
	wire [4-1:0] node4917;
	wire [4-1:0] node4920;
	wire [4-1:0] node4921;
	wire [4-1:0] node4924;
	wire [4-1:0] node4927;
	wire [4-1:0] node4928;
	wire [4-1:0] node4931;
	wire [4-1:0] node4932;
	wire [4-1:0] node4936;
	wire [4-1:0] node4937;
	wire [4-1:0] node4938;
	wire [4-1:0] node4940;
	wire [4-1:0] node4943;
	wire [4-1:0] node4944;
	wire [4-1:0] node4947;
	wire [4-1:0] node4950;
	wire [4-1:0] node4951;
	wire [4-1:0] node4952;
	wire [4-1:0] node4955;
	wire [4-1:0] node4958;
	wire [4-1:0] node4959;
	wire [4-1:0] node4962;
	wire [4-1:0] node4965;
	wire [4-1:0] node4966;
	wire [4-1:0] node4967;
	wire [4-1:0] node4968;
	wire [4-1:0] node4971;
	wire [4-1:0] node4972;
	wire [4-1:0] node4975;
	wire [4-1:0] node4978;
	wire [4-1:0] node4979;
	wire [4-1:0] node4980;
	wire [4-1:0] node4984;
	wire [4-1:0] node4985;
	wire [4-1:0] node4989;
	wire [4-1:0] node4990;
	wire [4-1:0] node4991;
	wire [4-1:0] node4994;
	wire [4-1:0] node4995;
	wire [4-1:0] node4999;
	wire [4-1:0] node5000;
	wire [4-1:0] node5002;
	wire [4-1:0] node5005;
	wire [4-1:0] node5006;
	wire [4-1:0] node5010;
	wire [4-1:0] node5011;
	wire [4-1:0] node5012;
	wire [4-1:0] node5013;
	wire [4-1:0] node5014;
	wire [4-1:0] node5017;
	wire [4-1:0] node5019;
	wire [4-1:0] node5022;
	wire [4-1:0] node5023;
	wire [4-1:0] node5026;
	wire [4-1:0] node5028;
	wire [4-1:0] node5031;
	wire [4-1:0] node5032;
	wire [4-1:0] node5033;
	wire [4-1:0] node5034;
	wire [4-1:0] node5037;
	wire [4-1:0] node5040;
	wire [4-1:0] node5041;
	wire [4-1:0] node5044;
	wire [4-1:0] node5047;
	wire [4-1:0] node5048;
	wire [4-1:0] node5050;
	wire [4-1:0] node5053;
	wire [4-1:0] node5054;
	wire [4-1:0] node5058;
	wire [4-1:0] node5059;
	wire [4-1:0] node5060;
	wire [4-1:0] node5061;
	wire [4-1:0] node5063;
	wire [4-1:0] node5066;
	wire [4-1:0] node5067;
	wire [4-1:0] node5070;
	wire [4-1:0] node5073;
	wire [4-1:0] node5074;
	wire [4-1:0] node5077;
	wire [4-1:0] node5078;
	wire [4-1:0] node5082;
	wire [4-1:0] node5083;
	wire [4-1:0] node5084;
	wire [4-1:0] node5085;
	wire [4-1:0] node5088;
	wire [4-1:0] node5091;
	wire [4-1:0] node5092;
	wire [4-1:0] node5095;
	wire [4-1:0] node5098;
	wire [4-1:0] node5099;
	wire [4-1:0] node5100;
	wire [4-1:0] node5104;
	wire [4-1:0] node5105;
	wire [4-1:0] node5108;
	wire [4-1:0] node5111;
	wire [4-1:0] node5112;
	wire [4-1:0] node5113;
	wire [4-1:0] node5114;
	wire [4-1:0] node5115;
	wire [4-1:0] node5116;
	wire [4-1:0] node5118;
	wire [4-1:0] node5122;
	wire [4-1:0] node5123;
	wire [4-1:0] node5127;
	wire [4-1:0] node5128;
	wire [4-1:0] node5129;
	wire [4-1:0] node5131;
	wire [4-1:0] node5134;
	wire [4-1:0] node5137;
	wire [4-1:0] node5138;
	wire [4-1:0] node5140;
	wire [4-1:0] node5143;
	wire [4-1:0] node5144;
	wire [4-1:0] node5147;
	wire [4-1:0] node5150;
	wire [4-1:0] node5151;
	wire [4-1:0] node5152;
	wire [4-1:0] node5153;
	wire [4-1:0] node5156;
	wire [4-1:0] node5157;
	wire [4-1:0] node5160;
	wire [4-1:0] node5163;
	wire [4-1:0] node5164;
	wire [4-1:0] node5167;
	wire [4-1:0] node5168;
	wire [4-1:0] node5171;
	wire [4-1:0] node5174;
	wire [4-1:0] node5175;
	wire [4-1:0] node5176;
	wire [4-1:0] node5179;
	wire [4-1:0] node5182;
	wire [4-1:0] node5183;
	wire [4-1:0] node5185;
	wire [4-1:0] node5188;
	wire [4-1:0] node5189;
	wire [4-1:0] node5192;
	wire [4-1:0] node5195;
	wire [4-1:0] node5196;
	wire [4-1:0] node5197;
	wire [4-1:0] node5198;
	wire [4-1:0] node5199;
	wire [4-1:0] node5200;
	wire [4-1:0] node5204;
	wire [4-1:0] node5206;
	wire [4-1:0] node5209;
	wire [4-1:0] node5210;
	wire [4-1:0] node5211;
	wire [4-1:0] node5214;
	wire [4-1:0] node5217;
	wire [4-1:0] node5218;
	wire [4-1:0] node5221;
	wire [4-1:0] node5224;
	wire [4-1:0] node5225;
	wire [4-1:0] node5226;
	wire [4-1:0] node5228;
	wire [4-1:0] node5231;
	wire [4-1:0] node5232;
	wire [4-1:0] node5235;
	wire [4-1:0] node5238;
	wire [4-1:0] node5239;
	wire [4-1:0] node5240;
	wire [4-1:0] node5244;
	wire [4-1:0] node5245;
	wire [4-1:0] node5248;
	wire [4-1:0] node5251;
	wire [4-1:0] node5252;
	wire [4-1:0] node5253;
	wire [4-1:0] node5254;
	wire [4-1:0] node5255;
	wire [4-1:0] node5258;
	wire [4-1:0] node5261;
	wire [4-1:0] node5262;
	wire [4-1:0] node5266;
	wire [4-1:0] node5267;
	wire [4-1:0] node5268;
	wire [4-1:0] node5271;
	wire [4-1:0] node5274;
	wire [4-1:0] node5276;
	wire [4-1:0] node5279;
	wire [4-1:0] node5280;
	wire [4-1:0] node5281;
	wire [4-1:0] node5282;
	wire [4-1:0] node5285;
	wire [4-1:0] node5288;
	wire [4-1:0] node5289;
	wire [4-1:0] node5292;
	wire [4-1:0] node5295;
	wire [4-1:0] node5296;
	wire [4-1:0] node5297;
	wire [4-1:0] node5300;
	wire [4-1:0] node5303;
	wire [4-1:0] node5304;
	wire [4-1:0] node5307;
	wire [4-1:0] node5310;
	wire [4-1:0] node5311;
	wire [4-1:0] node5312;
	wire [4-1:0] node5313;
	wire [4-1:0] node5314;
	wire [4-1:0] node5315;
	wire [4-1:0] node5316;
	wire [4-1:0] node5319;
	wire [4-1:0] node5321;
	wire [4-1:0] node5324;
	wire [4-1:0] node5325;
	wire [4-1:0] node5327;
	wire [4-1:0] node5330;
	wire [4-1:0] node5331;
	wire [4-1:0] node5335;
	wire [4-1:0] node5336;
	wire [4-1:0] node5337;
	wire [4-1:0] node5340;
	wire [4-1:0] node5341;
	wire [4-1:0] node5344;
	wire [4-1:0] node5347;
	wire [4-1:0] node5349;
	wire [4-1:0] node5350;
	wire [4-1:0] node5354;
	wire [4-1:0] node5355;
	wire [4-1:0] node5356;
	wire [4-1:0] node5357;
	wire [4-1:0] node5360;
	wire [4-1:0] node5363;
	wire [4-1:0] node5364;
	wire [4-1:0] node5367;
	wire [4-1:0] node5370;
	wire [4-1:0] node5371;
	wire [4-1:0] node5372;
	wire [4-1:0] node5374;
	wire [4-1:0] node5377;
	wire [4-1:0] node5380;
	wire [4-1:0] node5381;
	wire [4-1:0] node5382;
	wire [4-1:0] node5385;
	wire [4-1:0] node5388;
	wire [4-1:0] node5389;
	wire [4-1:0] node5393;
	wire [4-1:0] node5394;
	wire [4-1:0] node5395;
	wire [4-1:0] node5396;
	wire [4-1:0] node5397;
	wire [4-1:0] node5399;
	wire [4-1:0] node5402;
	wire [4-1:0] node5403;
	wire [4-1:0] node5406;
	wire [4-1:0] node5409;
	wire [4-1:0] node5411;
	wire [4-1:0] node5414;
	wire [4-1:0] node5415;
	wire [4-1:0] node5416;
	wire [4-1:0] node5418;
	wire [4-1:0] node5421;
	wire [4-1:0] node5423;
	wire [4-1:0] node5426;
	wire [4-1:0] node5427;
	wire [4-1:0] node5428;
	wire [4-1:0] node5432;
	wire [4-1:0] node5435;
	wire [4-1:0] node5436;
	wire [4-1:0] node5437;
	wire [4-1:0] node5438;
	wire [4-1:0] node5440;
	wire [4-1:0] node5443;
	wire [4-1:0] node5444;
	wire [4-1:0] node5447;
	wire [4-1:0] node5450;
	wire [4-1:0] node5451;
	wire [4-1:0] node5452;
	wire [4-1:0] node5456;
	wire [4-1:0] node5458;
	wire [4-1:0] node5461;
	wire [4-1:0] node5462;
	wire [4-1:0] node5463;
	wire [4-1:0] node5464;
	wire [4-1:0] node5468;
	wire [4-1:0] node5469;
	wire [4-1:0] node5472;
	wire [4-1:0] node5475;
	wire [4-1:0] node5476;
	wire [4-1:0] node5477;
	wire [4-1:0] node5480;
	wire [4-1:0] node5483;
	wire [4-1:0] node5484;
	wire [4-1:0] node5487;
	wire [4-1:0] node5490;
	wire [4-1:0] node5491;
	wire [4-1:0] node5492;
	wire [4-1:0] node5493;
	wire [4-1:0] node5494;
	wire [4-1:0] node5495;
	wire [4-1:0] node5498;
	wire [4-1:0] node5500;
	wire [4-1:0] node5503;
	wire [4-1:0] node5504;
	wire [4-1:0] node5507;
	wire [4-1:0] node5510;
	wire [4-1:0] node5511;
	wire [4-1:0] node5512;
	wire [4-1:0] node5515;
	wire [4-1:0] node5518;
	wire [4-1:0] node5519;
	wire [4-1:0] node5520;
	wire [4-1:0] node5523;
	wire [4-1:0] node5526;
	wire [4-1:0] node5527;
	wire [4-1:0] node5531;
	wire [4-1:0] node5532;
	wire [4-1:0] node5533;
	wire [4-1:0] node5534;
	wire [4-1:0] node5536;
	wire [4-1:0] node5539;
	wire [4-1:0] node5542;
	wire [4-1:0] node5543;
	wire [4-1:0] node5544;
	wire [4-1:0] node5548;
	wire [4-1:0] node5551;
	wire [4-1:0] node5552;
	wire [4-1:0] node5553;
	wire [4-1:0] node5554;
	wire [4-1:0] node5557;
	wire [4-1:0] node5560;
	wire [4-1:0] node5561;
	wire [4-1:0] node5564;
	wire [4-1:0] node5567;
	wire [4-1:0] node5568;
	wire [4-1:0] node5571;
	wire [4-1:0] node5572;
	wire [4-1:0] node5575;
	wire [4-1:0] node5578;
	wire [4-1:0] node5579;
	wire [4-1:0] node5580;
	wire [4-1:0] node5581;
	wire [4-1:0] node5582;
	wire [4-1:0] node5583;
	wire [4-1:0] node5586;
	wire [4-1:0] node5589;
	wire [4-1:0] node5590;
	wire [4-1:0] node5593;
	wire [4-1:0] node5596;
	wire [4-1:0] node5597;
	wire [4-1:0] node5598;
	wire [4-1:0] node5601;
	wire [4-1:0] node5604;
	wire [4-1:0] node5606;
	wire [4-1:0] node5609;
	wire [4-1:0] node5610;
	wire [4-1:0] node5611;
	wire [4-1:0] node5614;
	wire [4-1:0] node5617;
	wire [4-1:0] node5618;
	wire [4-1:0] node5619;
	wire [4-1:0] node5622;
	wire [4-1:0] node5625;
	wire [4-1:0] node5628;
	wire [4-1:0] node5629;
	wire [4-1:0] node5630;
	wire [4-1:0] node5631;
	wire [4-1:0] node5633;
	wire [4-1:0] node5636;
	wire [4-1:0] node5637;
	wire [4-1:0] node5640;
	wire [4-1:0] node5643;
	wire [4-1:0] node5644;
	wire [4-1:0] node5645;
	wire [4-1:0] node5648;
	wire [4-1:0] node5651;
	wire [4-1:0] node5652;
	wire [4-1:0] node5655;
	wire [4-1:0] node5658;
	wire [4-1:0] node5659;
	wire [4-1:0] node5660;
	wire [4-1:0] node5661;
	wire [4-1:0] node5665;
	wire [4-1:0] node5667;
	wire [4-1:0] node5670;
	wire [4-1:0] node5671;
	wire [4-1:0] node5672;
	wire [4-1:0] node5675;
	wire [4-1:0] node5678;
	wire [4-1:0] node5680;
	wire [4-1:0] node5683;
	wire [4-1:0] node5684;
	wire [4-1:0] node5685;
	wire [4-1:0] node5686;
	wire [4-1:0] node5687;
	wire [4-1:0] node5688;
	wire [4-1:0] node5689;
	wire [4-1:0] node5690;
	wire [4-1:0] node5693;
	wire [4-1:0] node5694;
	wire [4-1:0] node5696;
	wire [4-1:0] node5697;
	wire [4-1:0] node5700;
	wire [4-1:0] node5703;
	wire [4-1:0] node5704;
	wire [4-1:0] node5706;
	wire [4-1:0] node5710;
	wire [4-1:0] node5711;
	wire [4-1:0] node5714;
	wire [4-1:0] node5715;
	wire [4-1:0] node5717;
	wire [4-1:0] node5718;
	wire [4-1:0] node5722;
	wire [4-1:0] node5723;
	wire [4-1:0] node5724;
	wire [4-1:0] node5727;
	wire [4-1:0] node5731;
	wire [4-1:0] node5732;
	wire [4-1:0] node5733;
	wire [4-1:0] node5734;
	wire [4-1:0] node5736;
	wire [4-1:0] node5739;
	wire [4-1:0] node5741;
	wire [4-1:0] node5744;
	wire [4-1:0] node5745;
	wire [4-1:0] node5747;
	wire [4-1:0] node5748;
	wire [4-1:0] node5751;
	wire [4-1:0] node5754;
	wire [4-1:0] node5755;
	wire [4-1:0] node5756;
	wire [4-1:0] node5760;
	wire [4-1:0] node5762;
	wire [4-1:0] node5765;
	wire [4-1:0] node5766;
	wire [4-1:0] node5767;
	wire [4-1:0] node5768;
	wire [4-1:0] node5772;
	wire [4-1:0] node5773;
	wire [4-1:0] node5777;
	wire [4-1:0] node5778;
	wire [4-1:0] node5779;
	wire [4-1:0] node5780;
	wire [4-1:0] node5784;
	wire [4-1:0] node5786;
	wire [4-1:0] node5789;
	wire [4-1:0] node5790;
	wire [4-1:0] node5791;
	wire [4-1:0] node5794;
	wire [4-1:0] node5797;
	wire [4-1:0] node5798;
	wire [4-1:0] node5802;
	wire [4-1:0] node5803;
	wire [4-1:0] node5804;
	wire [4-1:0] node5805;
	wire [4-1:0] node5806;
	wire [4-1:0] node5807;
	wire [4-1:0] node5810;
	wire [4-1:0] node5813;
	wire [4-1:0] node5814;
	wire [4-1:0] node5817;
	wire [4-1:0] node5820;
	wire [4-1:0] node5821;
	wire [4-1:0] node5822;
	wire [4-1:0] node5825;
	wire [4-1:0] node5828;
	wire [4-1:0] node5829;
	wire [4-1:0] node5832;
	wire [4-1:0] node5835;
	wire [4-1:0] node5836;
	wire [4-1:0] node5837;
	wire [4-1:0] node5838;
	wire [4-1:0] node5841;
	wire [4-1:0] node5844;
	wire [4-1:0] node5845;
	wire [4-1:0] node5849;
	wire [4-1:0] node5850;
	wire [4-1:0] node5851;
	wire [4-1:0] node5852;
	wire [4-1:0] node5855;
	wire [4-1:0] node5858;
	wire [4-1:0] node5859;
	wire [4-1:0] node5862;
	wire [4-1:0] node5865;
	wire [4-1:0] node5866;
	wire [4-1:0] node5870;
	wire [4-1:0] node5871;
	wire [4-1:0] node5872;
	wire [4-1:0] node5873;
	wire [4-1:0] node5874;
	wire [4-1:0] node5875;
	wire [4-1:0] node5879;
	wire [4-1:0] node5880;
	wire [4-1:0] node5884;
	wire [4-1:0] node5885;
	wire [4-1:0] node5886;
	wire [4-1:0] node5890;
	wire [4-1:0] node5893;
	wire [4-1:0] node5894;
	wire [4-1:0] node5895;
	wire [4-1:0] node5896;
	wire [4-1:0] node5897;
	wire [4-1:0] node5900;
	wire [4-1:0] node5903;
	wire [4-1:0] node5905;
	wire [4-1:0] node5908;
	wire [4-1:0] node5910;
	wire [4-1:0] node5913;
	wire [4-1:0] node5914;
	wire [4-1:0] node5916;
	wire [4-1:0] node5919;
	wire [4-1:0] node5922;
	wire [4-1:0] node5923;
	wire [4-1:0] node5924;
	wire [4-1:0] node5925;
	wire [4-1:0] node5926;
	wire [4-1:0] node5930;
	wire [4-1:0] node5931;
	wire [4-1:0] node5934;
	wire [4-1:0] node5937;
	wire [4-1:0] node5938;
	wire [4-1:0] node5940;
	wire [4-1:0] node5943;
	wire [4-1:0] node5944;
	wire [4-1:0] node5948;
	wire [4-1:0] node5949;
	wire [4-1:0] node5950;
	wire [4-1:0] node5953;
	wire [4-1:0] node5956;
	wire [4-1:0] node5957;
	wire [4-1:0] node5958;
	wire [4-1:0] node5961;
	wire [4-1:0] node5965;
	wire [4-1:0] node5966;
	wire [4-1:0] node5967;
	wire [4-1:0] node5968;
	wire [4-1:0] node5969;
	wire [4-1:0] node5970;
	wire [4-1:0] node5971;
	wire [4-1:0] node5974;
	wire [4-1:0] node5976;
	wire [4-1:0] node5979;
	wire [4-1:0] node5980;
	wire [4-1:0] node5982;
	wire [4-1:0] node5985;
	wire [4-1:0] node5988;
	wire [4-1:0] node5989;
	wire [4-1:0] node5990;
	wire [4-1:0] node5991;
	wire [4-1:0] node5994;
	wire [4-1:0] node5997;
	wire [4-1:0] node5998;
	wire [4-1:0] node6001;
	wire [4-1:0] node6004;
	wire [4-1:0] node6005;
	wire [4-1:0] node6006;
	wire [4-1:0] node6009;
	wire [4-1:0] node6012;
	wire [4-1:0] node6013;
	wire [4-1:0] node6016;
	wire [4-1:0] node6019;
	wire [4-1:0] node6020;
	wire [4-1:0] node6021;
	wire [4-1:0] node6022;
	wire [4-1:0] node6024;
	wire [4-1:0] node6027;
	wire [4-1:0] node6028;
	wire [4-1:0] node6032;
	wire [4-1:0] node6033;
	wire [4-1:0] node6036;
	wire [4-1:0] node6038;
	wire [4-1:0] node6041;
	wire [4-1:0] node6042;
	wire [4-1:0] node6043;
	wire [4-1:0] node6046;
	wire [4-1:0] node6047;
	wire [4-1:0] node6051;
	wire [4-1:0] node6052;
	wire [4-1:0] node6053;
	wire [4-1:0] node6057;
	wire [4-1:0] node6059;
	wire [4-1:0] node6062;
	wire [4-1:0] node6063;
	wire [4-1:0] node6064;
	wire [4-1:0] node6065;
	wire [4-1:0] node6066;
	wire [4-1:0] node6067;
	wire [4-1:0] node6070;
	wire [4-1:0] node6073;
	wire [4-1:0] node6074;
	wire [4-1:0] node6077;
	wire [4-1:0] node6080;
	wire [4-1:0] node6081;
	wire [4-1:0] node6082;
	wire [4-1:0] node6085;
	wire [4-1:0] node6088;
	wire [4-1:0] node6089;
	wire [4-1:0] node6092;
	wire [4-1:0] node6095;
	wire [4-1:0] node6096;
	wire [4-1:0] node6097;
	wire [4-1:0] node6098;
	wire [4-1:0] node6101;
	wire [4-1:0] node6104;
	wire [4-1:0] node6105;
	wire [4-1:0] node6108;
	wire [4-1:0] node6111;
	wire [4-1:0] node6112;
	wire [4-1:0] node6113;
	wire [4-1:0] node6116;
	wire [4-1:0] node6119;
	wire [4-1:0] node6120;
	wire [4-1:0] node6123;
	wire [4-1:0] node6126;
	wire [4-1:0] node6127;
	wire [4-1:0] node6128;
	wire [4-1:0] node6129;
	wire [4-1:0] node6131;
	wire [4-1:0] node6134;
	wire [4-1:0] node6137;
	wire [4-1:0] node6138;
	wire [4-1:0] node6140;
	wire [4-1:0] node6143;
	wire [4-1:0] node6145;
	wire [4-1:0] node6148;
	wire [4-1:0] node6149;
	wire [4-1:0] node6150;
	wire [4-1:0] node6152;
	wire [4-1:0] node6155;
	wire [4-1:0] node6156;
	wire [4-1:0] node6160;
	wire [4-1:0] node6161;
	wire [4-1:0] node6163;
	wire [4-1:0] node6166;
	wire [4-1:0] node6169;
	wire [4-1:0] node6170;
	wire [4-1:0] node6171;
	wire [4-1:0] node6172;
	wire [4-1:0] node6173;
	wire [4-1:0] node6174;
	wire [4-1:0] node6175;
	wire [4-1:0] node6178;
	wire [4-1:0] node6181;
	wire [4-1:0] node6182;
	wire [4-1:0] node6186;
	wire [4-1:0] node6187;
	wire [4-1:0] node6190;
	wire [4-1:0] node6192;
	wire [4-1:0] node6195;
	wire [4-1:0] node6196;
	wire [4-1:0] node6197;
	wire [4-1:0] node6198;
	wire [4-1:0] node6202;
	wire [4-1:0] node6204;
	wire [4-1:0] node6207;
	wire [4-1:0] node6208;
	wire [4-1:0] node6209;
	wire [4-1:0] node6212;
	wire [4-1:0] node6215;
	wire [4-1:0] node6216;
	wire [4-1:0] node6220;
	wire [4-1:0] node6221;
	wire [4-1:0] node6222;
	wire [4-1:0] node6223;
	wire [4-1:0] node6224;
	wire [4-1:0] node6227;
	wire [4-1:0] node6230;
	wire [4-1:0] node6231;
	wire [4-1:0] node6234;
	wire [4-1:0] node6237;
	wire [4-1:0] node6238;
	wire [4-1:0] node6239;
	wire [4-1:0] node6242;
	wire [4-1:0] node6245;
	wire [4-1:0] node6246;
	wire [4-1:0] node6249;
	wire [4-1:0] node6252;
	wire [4-1:0] node6253;
	wire [4-1:0] node6254;
	wire [4-1:0] node6256;
	wire [4-1:0] node6259;
	wire [4-1:0] node6260;
	wire [4-1:0] node6263;
	wire [4-1:0] node6266;
	wire [4-1:0] node6267;
	wire [4-1:0] node6270;
	wire [4-1:0] node6271;
	wire [4-1:0] node6275;
	wire [4-1:0] node6276;
	wire [4-1:0] node6277;
	wire [4-1:0] node6278;
	wire [4-1:0] node6279;
	wire [4-1:0] node6280;
	wire [4-1:0] node6283;
	wire [4-1:0] node6286;
	wire [4-1:0] node6287;
	wire [4-1:0] node6290;
	wire [4-1:0] node6293;
	wire [4-1:0] node6294;
	wire [4-1:0] node6295;
	wire [4-1:0] node6298;
	wire [4-1:0] node6301;
	wire [4-1:0] node6302;
	wire [4-1:0] node6306;
	wire [4-1:0] node6307;
	wire [4-1:0] node6308;
	wire [4-1:0] node6309;
	wire [4-1:0] node6312;
	wire [4-1:0] node6315;
	wire [4-1:0] node6316;
	wire [4-1:0] node6319;
	wire [4-1:0] node6322;
	wire [4-1:0] node6323;
	wire [4-1:0] node6324;
	wire [4-1:0] node6327;
	wire [4-1:0] node6330;
	wire [4-1:0] node6331;
	wire [4-1:0] node6334;
	wire [4-1:0] node6337;
	wire [4-1:0] node6338;
	wire [4-1:0] node6339;
	wire [4-1:0] node6340;
	wire [4-1:0] node6342;
	wire [4-1:0] node6345;
	wire [4-1:0] node6346;
	wire [4-1:0] node6349;
	wire [4-1:0] node6352;
	wire [4-1:0] node6353;
	wire [4-1:0] node6354;
	wire [4-1:0] node6357;
	wire [4-1:0] node6360;
	wire [4-1:0] node6361;
	wire [4-1:0] node6364;
	wire [4-1:0] node6367;
	wire [4-1:0] node6368;
	wire [4-1:0] node6369;
	wire [4-1:0] node6370;
	wire [4-1:0] node6373;
	wire [4-1:0] node6376;
	wire [4-1:0] node6377;
	wire [4-1:0] node6380;
	wire [4-1:0] node6383;
	wire [4-1:0] node6384;
	wire [4-1:0] node6386;
	wire [4-1:0] node6389;
	wire [4-1:0] node6390;
	wire [4-1:0] node6394;
	wire [4-1:0] node6395;
	wire [4-1:0] node6396;
	wire [4-1:0] node6397;
	wire [4-1:0] node6398;
	wire [4-1:0] node6399;
	wire [4-1:0] node6402;
	wire [4-1:0] node6403;
	wire [4-1:0] node6405;
	wire [4-1:0] node6406;
	wire [4-1:0] node6409;
	wire [4-1:0] node6412;
	wire [4-1:0] node6413;
	wire [4-1:0] node6417;
	wire [4-1:0] node6418;
	wire [4-1:0] node6421;
	wire [4-1:0] node6422;
	wire [4-1:0] node6424;
	wire [4-1:0] node6425;
	wire [4-1:0] node6429;
	wire [4-1:0] node6430;
	wire [4-1:0] node6431;
	wire [4-1:0] node6434;
	wire [4-1:0] node6438;
	wire [4-1:0] node6439;
	wire [4-1:0] node6440;
	wire [4-1:0] node6441;
	wire [4-1:0] node6443;
	wire [4-1:0] node6446;
	wire [4-1:0] node6448;
	wire [4-1:0] node6451;
	wire [4-1:0] node6452;
	wire [4-1:0] node6453;
	wire [4-1:0] node6455;
	wire [4-1:0] node6458;
	wire [4-1:0] node6459;
	wire [4-1:0] node6462;
	wire [4-1:0] node6465;
	wire [4-1:0] node6466;
	wire [4-1:0] node6467;
	wire [4-1:0] node6471;
	wire [4-1:0] node6473;
	wire [4-1:0] node6476;
	wire [4-1:0] node6477;
	wire [4-1:0] node6478;
	wire [4-1:0] node6479;
	wire [4-1:0] node6483;
	wire [4-1:0] node6484;
	wire [4-1:0] node6488;
	wire [4-1:0] node6489;
	wire [4-1:0] node6490;
	wire [4-1:0] node6491;
	wire [4-1:0] node6495;
	wire [4-1:0] node6497;
	wire [4-1:0] node6500;
	wire [4-1:0] node6501;
	wire [4-1:0] node6502;
	wire [4-1:0] node6505;
	wire [4-1:0] node6508;
	wire [4-1:0] node6509;
	wire [4-1:0] node6513;
	wire [4-1:0] node6514;
	wire [4-1:0] node6515;
	wire [4-1:0] node6516;
	wire [4-1:0] node6517;
	wire [4-1:0] node6518;
	wire [4-1:0] node6521;
	wire [4-1:0] node6524;
	wire [4-1:0] node6525;
	wire [4-1:0] node6526;
	wire [4-1:0] node6527;
	wire [4-1:0] node6530;
	wire [4-1:0] node6533;
	wire [4-1:0] node6534;
	wire [4-1:0] node6538;
	wire [4-1:0] node6539;
	wire [4-1:0] node6542;
	wire [4-1:0] node6545;
	wire [4-1:0] node6546;
	wire [4-1:0] node6547;
	wire [4-1:0] node6550;
	wire [4-1:0] node6553;
	wire [4-1:0] node6554;
	wire [4-1:0] node6557;
	wire [4-1:0] node6560;
	wire [4-1:0] node6561;
	wire [4-1:0] node6562;
	wire [4-1:0] node6563;
	wire [4-1:0] node6566;
	wire [4-1:0] node6569;
	wire [4-1:0] node6570;
	wire [4-1:0] node6573;
	wire [4-1:0] node6576;
	wire [4-1:0] node6577;
	wire [4-1:0] node6578;
	wire [4-1:0] node6581;
	wire [4-1:0] node6584;
	wire [4-1:0] node6585;
	wire [4-1:0] node6589;
	wire [4-1:0] node6590;
	wire [4-1:0] node6591;
	wire [4-1:0] node6592;
	wire [4-1:0] node6593;
	wire [4-1:0] node6594;
	wire [4-1:0] node6598;
	wire [4-1:0] node6599;
	wire [4-1:0] node6603;
	wire [4-1:0] node6604;
	wire [4-1:0] node6606;
	wire [4-1:0] node6609;
	wire [4-1:0] node6612;
	wire [4-1:0] node6613;
	wire [4-1:0] node6614;
	wire [4-1:0] node6615;
	wire [4-1:0] node6619;
	wire [4-1:0] node6620;
	wire [4-1:0] node6623;
	wire [4-1:0] node6626;
	wire [4-1:0] node6628;
	wire [4-1:0] node6629;
	wire [4-1:0] node6633;
	wire [4-1:0] node6634;
	wire [4-1:0] node6635;
	wire [4-1:0] node6636;
	wire [4-1:0] node6637;
	wire [4-1:0] node6641;
	wire [4-1:0] node6642;
	wire [4-1:0] node6645;
	wire [4-1:0] node6648;
	wire [4-1:0] node6649;
	wire [4-1:0] node6651;
	wire [4-1:0] node6654;
	wire [4-1:0] node6655;
	wire [4-1:0] node6659;
	wire [4-1:0] node6660;
	wire [4-1:0] node6661;
	wire [4-1:0] node6663;
	wire [4-1:0] node6666;
	wire [4-1:0] node6668;
	wire [4-1:0] node6671;
	wire [4-1:0] node6672;
	wire [4-1:0] node6675;
	wire [4-1:0] node6677;
	wire [4-1:0] node6680;
	wire [4-1:0] node6681;
	wire [4-1:0] node6682;
	wire [4-1:0] node6683;
	wire [4-1:0] node6684;
	wire [4-1:0] node6685;
	wire [4-1:0] node6686;
	wire [4-1:0] node6687;
	wire [4-1:0] node6690;
	wire [4-1:0] node6693;
	wire [4-1:0] node6694;
	wire [4-1:0] node6697;
	wire [4-1:0] node6700;
	wire [4-1:0] node6701;
	wire [4-1:0] node6702;
	wire [4-1:0] node6703;
	wire [4-1:0] node6706;
	wire [4-1:0] node6709;
	wire [4-1:0] node6710;
	wire [4-1:0] node6713;
	wire [4-1:0] node6716;
	wire [4-1:0] node6717;
	wire [4-1:0] node6720;
	wire [4-1:0] node6723;
	wire [4-1:0] node6724;
	wire [4-1:0] node6725;
	wire [4-1:0] node6726;
	wire [4-1:0] node6729;
	wire [4-1:0] node6732;
	wire [4-1:0] node6733;
	wire [4-1:0] node6736;
	wire [4-1:0] node6739;
	wire [4-1:0] node6740;
	wire [4-1:0] node6741;
	wire [4-1:0] node6742;
	wire [4-1:0] node6745;
	wire [4-1:0] node6748;
	wire [4-1:0] node6749;
	wire [4-1:0] node6753;
	wire [4-1:0] node6754;
	wire [4-1:0] node6755;
	wire [4-1:0] node6758;
	wire [4-1:0] node6761;
	wire [4-1:0] node6762;
	wire [4-1:0] node6765;
	wire [4-1:0] node6768;
	wire [4-1:0] node6769;
	wire [4-1:0] node6770;
	wire [4-1:0] node6771;
	wire [4-1:0] node6772;
	wire [4-1:0] node6775;
	wire [4-1:0] node6778;
	wire [4-1:0] node6779;
	wire [4-1:0] node6782;
	wire [4-1:0] node6785;
	wire [4-1:0] node6786;
	wire [4-1:0] node6787;
	wire [4-1:0] node6791;
	wire [4-1:0] node6794;
	wire [4-1:0] node6795;
	wire [4-1:0] node6796;
	wire [4-1:0] node6797;
	wire [4-1:0] node6800;
	wire [4-1:0] node6803;
	wire [4-1:0] node6804;
	wire [4-1:0] node6807;
	wire [4-1:0] node6810;
	wire [4-1:0] node6811;
	wire [4-1:0] node6814;
	wire [4-1:0] node6816;
	wire [4-1:0] node6819;
	wire [4-1:0] node6820;
	wire [4-1:0] node6821;
	wire [4-1:0] node6822;
	wire [4-1:0] node6823;
	wire [4-1:0] node6825;
	wire [4-1:0] node6828;
	wire [4-1:0] node6829;
	wire [4-1:0] node6833;
	wire [4-1:0] node6834;
	wire [4-1:0] node6837;
	wire [4-1:0] node6839;
	wire [4-1:0] node6842;
	wire [4-1:0] node6843;
	wire [4-1:0] node6844;
	wire [4-1:0] node6846;
	wire [4-1:0] node6849;
	wire [4-1:0] node6852;
	wire [4-1:0] node6853;
	wire [4-1:0] node6854;
	wire [4-1:0] node6858;
	wire [4-1:0] node6859;
	wire [4-1:0] node6863;
	wire [4-1:0] node6864;
	wire [4-1:0] node6865;
	wire [4-1:0] node6866;
	wire [4-1:0] node6867;
	wire [4-1:0] node6871;
	wire [4-1:0] node6874;
	wire [4-1:0] node6875;
	wire [4-1:0] node6877;
	wire [4-1:0] node6880;
	wire [4-1:0] node6882;
	wire [4-1:0] node6885;
	wire [4-1:0] node6886;
	wire [4-1:0] node6887;
	wire [4-1:0] node6888;
	wire [4-1:0] node6892;
	wire [4-1:0] node6893;
	wire [4-1:0] node6897;
	wire [4-1:0] node6898;
	wire [4-1:0] node6899;
	wire [4-1:0] node6903;
	wire [4-1:0] node6906;
	wire [4-1:0] node6907;
	wire [4-1:0] node6908;
	wire [4-1:0] node6909;
	wire [4-1:0] node6910;
	wire [4-1:0] node6911;
	wire [4-1:0] node6912;
	wire [4-1:0] node6915;
	wire [4-1:0] node6918;
	wire [4-1:0] node6919;
	wire [4-1:0] node6923;
	wire [4-1:0] node6924;
	wire [4-1:0] node6926;
	wire [4-1:0] node6927;
	wire [4-1:0] node6930;
	wire [4-1:0] node6933;
	wire [4-1:0] node6934;
	wire [4-1:0] node6937;
	wire [4-1:0] node6940;
	wire [4-1:0] node6941;
	wire [4-1:0] node6942;
	wire [4-1:0] node6943;
	wire [4-1:0] node6947;
	wire [4-1:0] node6949;
	wire [4-1:0] node6952;
	wire [4-1:0] node6953;
	wire [4-1:0] node6954;
	wire [4-1:0] node6957;
	wire [4-1:0] node6960;
	wire [4-1:0] node6961;
	wire [4-1:0] node6965;
	wire [4-1:0] node6966;
	wire [4-1:0] node6967;
	wire [4-1:0] node6968;
	wire [4-1:0] node6969;
	wire [4-1:0] node6973;
	wire [4-1:0] node6976;
	wire [4-1:0] node6977;
	wire [4-1:0] node6979;
	wire [4-1:0] node6982;
	wire [4-1:0] node6983;
	wire [4-1:0] node6986;
	wire [4-1:0] node6989;
	wire [4-1:0] node6990;
	wire [4-1:0] node6991;
	wire [4-1:0] node6992;
	wire [4-1:0] node6995;
	wire [4-1:0] node6998;
	wire [4-1:0] node7000;
	wire [4-1:0] node7003;
	wire [4-1:0] node7004;
	wire [4-1:0] node7005;
	wire [4-1:0] node7009;
	wire [4-1:0] node7011;
	wire [4-1:0] node7014;
	wire [4-1:0] node7015;
	wire [4-1:0] node7016;
	wire [4-1:0] node7017;
	wire [4-1:0] node7018;
	wire [4-1:0] node7019;
	wire [4-1:0] node7022;
	wire [4-1:0] node7025;
	wire [4-1:0] node7026;
	wire [4-1:0] node7029;
	wire [4-1:0] node7032;
	wire [4-1:0] node7033;
	wire [4-1:0] node7034;
	wire [4-1:0] node7037;
	wire [4-1:0] node7040;
	wire [4-1:0] node7041;
	wire [4-1:0] node7045;
	wire [4-1:0] node7046;
	wire [4-1:0] node7047;
	wire [4-1:0] node7048;
	wire [4-1:0] node7051;
	wire [4-1:0] node7054;
	wire [4-1:0] node7055;
	wire [4-1:0] node7058;
	wire [4-1:0] node7061;
	wire [4-1:0] node7062;
	wire [4-1:0] node7063;
	wire [4-1:0] node7066;
	wire [4-1:0] node7069;
	wire [4-1:0] node7070;
	wire [4-1:0] node7073;
	wire [4-1:0] node7076;
	wire [4-1:0] node7077;
	wire [4-1:0] node7078;
	wire [4-1:0] node7079;
	wire [4-1:0] node7080;
	wire [4-1:0] node7084;
	wire [4-1:0] node7085;
	wire [4-1:0] node7088;
	wire [4-1:0] node7091;
	wire [4-1:0] node7092;
	wire [4-1:0] node7093;
	wire [4-1:0] node7096;
	wire [4-1:0] node7099;
	wire [4-1:0] node7100;
	wire [4-1:0] node7103;
	wire [4-1:0] node7106;
	wire [4-1:0] node7107;
	wire [4-1:0] node7108;
	wire [4-1:0] node7109;
	wire [4-1:0] node7112;
	wire [4-1:0] node7115;
	wire [4-1:0] node7116;
	wire [4-1:0] node7119;
	wire [4-1:0] node7122;
	wire [4-1:0] node7123;
	wire [4-1:0] node7124;
	wire [4-1:0] node7128;
	wire [4-1:0] node7129;
	wire [4-1:0] node7133;
	wire [4-1:0] node7134;
	wire [4-1:0] node7135;
	wire [4-1:0] node7136;
	wire [4-1:0] node7137;
	wire [4-1:0] node7138;
	wire [4-1:0] node7139;
	wire [4-1:0] node7142;
	wire [4-1:0] node7143;
	wire [4-1:0] node7145;
	wire [4-1:0] node7146;
	wire [4-1:0] node7149;
	wire [4-1:0] node7152;
	wire [4-1:0] node7153;
	wire [4-1:0] node7155;
	wire [4-1:0] node7159;
	wire [4-1:0] node7160;
	wire [4-1:0] node7163;
	wire [4-1:0] node7164;
	wire [4-1:0] node7166;
	wire [4-1:0] node7167;
	wire [4-1:0] node7171;
	wire [4-1:0] node7172;
	wire [4-1:0] node7173;
	wire [4-1:0] node7176;
	wire [4-1:0] node7180;
	wire [4-1:0] node7181;
	wire [4-1:0] node7182;
	wire [4-1:0] node7183;
	wire [4-1:0] node7185;
	wire [4-1:0] node7188;
	wire [4-1:0] node7190;
	wire [4-1:0] node7193;
	wire [4-1:0] node7194;
	wire [4-1:0] node7195;
	wire [4-1:0] node7197;
	wire [4-1:0] node7200;
	wire [4-1:0] node7201;
	wire [4-1:0] node7204;
	wire [4-1:0] node7207;
	wire [4-1:0] node7208;
	wire [4-1:0] node7209;
	wire [4-1:0] node7213;
	wire [4-1:0] node7215;
	wire [4-1:0] node7218;
	wire [4-1:0] node7219;
	wire [4-1:0] node7220;
	wire [4-1:0] node7221;
	wire [4-1:0] node7225;
	wire [4-1:0] node7226;
	wire [4-1:0] node7230;
	wire [4-1:0] node7231;
	wire [4-1:0] node7232;
	wire [4-1:0] node7233;
	wire [4-1:0] node7237;
	wire [4-1:0] node7239;
	wire [4-1:0] node7242;
	wire [4-1:0] node7243;
	wire [4-1:0] node7244;
	wire [4-1:0] node7247;
	wire [4-1:0] node7250;
	wire [4-1:0] node7251;
	wire [4-1:0] node7255;
	wire [4-1:0] node7256;
	wire [4-1:0] node7257;
	wire [4-1:0] node7258;
	wire [4-1:0] node7259;
	wire [4-1:0] node7260;
	wire [4-1:0] node7261;
	wire [4-1:0] node7264;
	wire [4-1:0] node7267;
	wire [4-1:0] node7268;
	wire [4-1:0] node7269;
	wire [4-1:0] node7272;
	wire [4-1:0] node7275;
	wire [4-1:0] node7277;
	wire [4-1:0] node7280;
	wire [4-1:0] node7282;
	wire [4-1:0] node7285;
	wire [4-1:0] node7286;
	wire [4-1:0] node7287;
	wire [4-1:0] node7288;
	wire [4-1:0] node7291;
	wire [4-1:0] node7294;
	wire [4-1:0] node7295;
	wire [4-1:0] node7296;
	wire [4-1:0] node7299;
	wire [4-1:0] node7302;
	wire [4-1:0] node7303;
	wire [4-1:0] node7306;
	wire [4-1:0] node7309;
	wire [4-1:0] node7311;
	wire [4-1:0] node7314;
	wire [4-1:0] node7315;
	wire [4-1:0] node7316;
	wire [4-1:0] node7317;
	wire [4-1:0] node7320;
	wire [4-1:0] node7323;
	wire [4-1:0] node7324;
	wire [4-1:0] node7327;
	wire [4-1:0] node7330;
	wire [4-1:0] node7331;
	wire [4-1:0] node7332;
	wire [4-1:0] node7335;
	wire [4-1:0] node7338;
	wire [4-1:0] node7339;
	wire [4-1:0] node7342;
	wire [4-1:0] node7345;
	wire [4-1:0] node7346;
	wire [4-1:0] node7347;
	wire [4-1:0] node7348;
	wire [4-1:0] node7349;
	wire [4-1:0] node7350;
	wire [4-1:0] node7354;
	wire [4-1:0] node7355;
	wire [4-1:0] node7359;
	wire [4-1:0] node7360;
	wire [4-1:0] node7361;
	wire [4-1:0] node7365;
	wire [4-1:0] node7368;
	wire [4-1:0] node7369;
	wire [4-1:0] node7370;
	wire [4-1:0] node7371;
	wire [4-1:0] node7375;
	wire [4-1:0] node7377;
	wire [4-1:0] node7380;
	wire [4-1:0] node7381;
	wire [4-1:0] node7383;
	wire [4-1:0] node7386;
	wire [4-1:0] node7387;
	wire [4-1:0] node7391;
	wire [4-1:0] node7392;
	wire [4-1:0] node7393;
	wire [4-1:0] node7394;
	wire [4-1:0] node7395;
	wire [4-1:0] node7398;
	wire [4-1:0] node7401;
	wire [4-1:0] node7403;
	wire [4-1:0] node7406;
	wire [4-1:0] node7407;
	wire [4-1:0] node7409;
	wire [4-1:0] node7412;
	wire [4-1:0] node7414;
	wire [4-1:0] node7417;
	wire [4-1:0] node7418;
	wire [4-1:0] node7419;
	wire [4-1:0] node7422;
	wire [4-1:0] node7424;
	wire [4-1:0] node7427;
	wire [4-1:0] node7428;
	wire [4-1:0] node7431;
	wire [4-1:0] node7432;
	wire [4-1:0] node7436;
	wire [4-1:0] node7437;
	wire [4-1:0] node7438;
	wire [4-1:0] node7439;
	wire [4-1:0] node7440;
	wire [4-1:0] node7441;
	wire [4-1:0] node7442;
	wire [4-1:0] node7444;
	wire [4-1:0] node7447;
	wire [4-1:0] node7449;
	wire [4-1:0] node7452;
	wire [4-1:0] node7453;
	wire [4-1:0] node7455;
	wire [4-1:0] node7458;
	wire [4-1:0] node7460;
	wire [4-1:0] node7463;
	wire [4-1:0] node7464;
	wire [4-1:0] node7465;
	wire [4-1:0] node7466;
	wire [4-1:0] node7470;
	wire [4-1:0] node7472;
	wire [4-1:0] node7475;
	wire [4-1:0] node7476;
	wire [4-1:0] node7477;
	wire [4-1:0] node7481;
	wire [4-1:0] node7483;
	wire [4-1:0] node7486;
	wire [4-1:0] node7487;
	wire [4-1:0] node7488;
	wire [4-1:0] node7490;
	wire [4-1:0] node7491;
	wire [4-1:0] node7492;
	wire [4-1:0] node7495;
	wire [4-1:0] node7498;
	wire [4-1:0] node7499;
	wire [4-1:0] node7502;
	wire [4-1:0] node7505;
	wire [4-1:0] node7506;
	wire [4-1:0] node7507;
	wire [4-1:0] node7511;
	wire [4-1:0] node7512;
	wire [4-1:0] node7516;
	wire [4-1:0] node7517;
	wire [4-1:0] node7518;
	wire [4-1:0] node7520;
	wire [4-1:0] node7523;
	wire [4-1:0] node7524;
	wire [4-1:0] node7528;
	wire [4-1:0] node7529;
	wire [4-1:0] node7530;
	wire [4-1:0] node7534;
	wire [4-1:0] node7535;
	wire [4-1:0] node7539;
	wire [4-1:0] node7540;
	wire [4-1:0] node7541;
	wire [4-1:0] node7542;
	wire [4-1:0] node7543;
	wire [4-1:0] node7545;
	wire [4-1:0] node7548;
	wire [4-1:0] node7550;
	wire [4-1:0] node7553;
	wire [4-1:0] node7554;
	wire [4-1:0] node7555;
	wire [4-1:0] node7559;
	wire [4-1:0] node7560;
	wire [4-1:0] node7564;
	wire [4-1:0] node7565;
	wire [4-1:0] node7566;
	wire [4-1:0] node7567;
	wire [4-1:0] node7571;
	wire [4-1:0] node7573;
	wire [4-1:0] node7576;
	wire [4-1:0] node7577;
	wire [4-1:0] node7579;
	wire [4-1:0] node7582;
	wire [4-1:0] node7583;
	wire [4-1:0] node7587;
	wire [4-1:0] node7588;
	wire [4-1:0] node7589;
	wire [4-1:0] node7591;
	wire [4-1:0] node7592;
	wire [4-1:0] node7595;
	wire [4-1:0] node7598;
	wire [4-1:0] node7599;
	wire [4-1:0] node7601;
	wire [4-1:0] node7604;
	wire [4-1:0] node7606;
	wire [4-1:0] node7609;
	wire [4-1:0] node7610;
	wire [4-1:0] node7611;
	wire [4-1:0] node7612;
	wire [4-1:0] node7614;
	wire [4-1:0] node7617;
	wire [4-1:0] node7618;
	wire [4-1:0] node7623;
	wire [4-1:0] node7624;
	wire [4-1:0] node7626;
	wire [4-1:0] node7629;
	wire [4-1:0] node7631;
	wire [4-1:0] node7634;
	wire [4-1:0] node7635;
	wire [4-1:0] node7636;
	wire [4-1:0] node7637;
	wire [4-1:0] node7638;
	wire [4-1:0] node7639;
	wire [4-1:0] node7641;
	wire [4-1:0] node7644;
	wire [4-1:0] node7645;
	wire [4-1:0] node7649;
	wire [4-1:0] node7650;
	wire [4-1:0] node7651;
	wire [4-1:0] node7655;
	wire [4-1:0] node7657;
	wire [4-1:0] node7660;
	wire [4-1:0] node7661;
	wire [4-1:0] node7662;
	wire [4-1:0] node7663;
	wire [4-1:0] node7667;
	wire [4-1:0] node7668;
	wire [4-1:0] node7672;
	wire [4-1:0] node7673;
	wire [4-1:0] node7675;
	wire [4-1:0] node7678;
	wire [4-1:0] node7680;
	wire [4-1:0] node7683;
	wire [4-1:0] node7684;
	wire [4-1:0] node7685;
	wire [4-1:0] node7686;
	wire [4-1:0] node7688;
	wire [4-1:0] node7691;
	wire [4-1:0] node7693;
	wire [4-1:0] node7696;
	wire [4-1:0] node7697;
	wire [4-1:0] node7698;
	wire [4-1:0] node7702;
	wire [4-1:0] node7704;
	wire [4-1:0] node7707;
	wire [4-1:0] node7708;
	wire [4-1:0] node7709;
	wire [4-1:0] node7711;
	wire [4-1:0] node7714;
	wire [4-1:0] node7716;
	wire [4-1:0] node7719;
	wire [4-1:0] node7720;
	wire [4-1:0] node7722;
	wire [4-1:0] node7725;
	wire [4-1:0] node7727;
	wire [4-1:0] node7730;
	wire [4-1:0] node7731;
	wire [4-1:0] node7732;
	wire [4-1:0] node7733;
	wire [4-1:0] node7734;
	wire [4-1:0] node7735;
	wire [4-1:0] node7739;
	wire [4-1:0] node7740;
	wire [4-1:0] node7744;
	wire [4-1:0] node7745;
	wire [4-1:0] node7746;
	wire [4-1:0] node7750;
	wire [4-1:0] node7752;
	wire [4-1:0] node7755;
	wire [4-1:0] node7756;
	wire [4-1:0] node7757;
	wire [4-1:0] node7759;
	wire [4-1:0] node7762;
	wire [4-1:0] node7763;
	wire [4-1:0] node7767;
	wire [4-1:0] node7768;
	wire [4-1:0] node7770;
	wire [4-1:0] node7773;
	wire [4-1:0] node7774;
	wire [4-1:0] node7778;
	wire [4-1:0] node7779;
	wire [4-1:0] node7780;
	wire [4-1:0] node7781;
	wire [4-1:0] node7782;
	wire [4-1:0] node7785;
	wire [4-1:0] node7789;
	wire [4-1:0] node7790;
	wire [4-1:0] node7792;
	wire [4-1:0] node7795;
	wire [4-1:0] node7797;
	wire [4-1:0] node7800;
	wire [4-1:0] node7801;
	wire [4-1:0] node7802;
	wire [4-1:0] node7803;
	wire [4-1:0] node7807;
	wire [4-1:0] node7808;
	wire [4-1:0] node7812;
	wire [4-1:0] node7814;
	wire [4-1:0] node7816;
	wire [4-1:0] node7819;
	wire [4-1:0] node7820;
	wire [4-1:0] node7821;
	wire [4-1:0] node7822;
	wire [4-1:0] node7823;
	wire [4-1:0] node7824;
	wire [4-1:0] node7826;
	wire [4-1:0] node7827;
	wire [4-1:0] node7828;
	wire [4-1:0] node7829;
	wire [4-1:0] node7832;
	wire [4-1:0] node7835;
	wire [4-1:0] node7837;
	wire [4-1:0] node7840;
	wire [4-1:0] node7841;
	wire [4-1:0] node7844;
	wire [4-1:0] node7847;
	wire [4-1:0] node7849;
	wire [4-1:0] node7850;
	wire [4-1:0] node7853;
	wire [4-1:0] node7856;
	wire [4-1:0] node7857;
	wire [4-1:0] node7858;
	wire [4-1:0] node7859;
	wire [4-1:0] node7861;
	wire [4-1:0] node7864;
	wire [4-1:0] node7865;
	wire [4-1:0] node7869;
	wire [4-1:0] node7870;
	wire [4-1:0] node7871;
	wire [4-1:0] node7875;
	wire [4-1:0] node7876;
	wire [4-1:0] node7880;
	wire [4-1:0] node7881;
	wire [4-1:0] node7882;
	wire [4-1:0] node7884;
	wire [4-1:0] node7887;
	wire [4-1:0] node7889;
	wire [4-1:0] node7892;
	wire [4-1:0] node7894;
	wire [4-1:0] node7895;
	wire [4-1:0] node7897;
	wire [4-1:0] node7900;
	wire [4-1:0] node7901;
	wire [4-1:0] node7904;
	wire [4-1:0] node7907;
	wire [4-1:0] node7908;
	wire [4-1:0] node7909;
	wire [4-1:0] node7910;
	wire [4-1:0] node7911;
	wire [4-1:0] node7913;
	wire [4-1:0] node7916;
	wire [4-1:0] node7917;
	wire [4-1:0] node7921;
	wire [4-1:0] node7922;
	wire [4-1:0] node7925;
	wire [4-1:0] node7927;
	wire [4-1:0] node7930;
	wire [4-1:0] node7931;
	wire [4-1:0] node7932;
	wire [4-1:0] node7933;
	wire [4-1:0] node7937;
	wire [4-1:0] node7938;
	wire [4-1:0] node7942;
	wire [4-1:0] node7943;
	wire [4-1:0] node7944;
	wire [4-1:0] node7948;
	wire [4-1:0] node7949;
	wire [4-1:0] node7953;
	wire [4-1:0] node7954;
	wire [4-1:0] node7955;
	wire [4-1:0] node7957;
	wire [4-1:0] node7958;
	wire [4-1:0] node7961;
	wire [4-1:0] node7964;
	wire [4-1:0] node7965;
	wire [4-1:0] node7966;
	wire [4-1:0] node7970;
	wire [4-1:0] node7971;
	wire [4-1:0] node7975;
	wire [4-1:0] node7976;
	wire [4-1:0] node7977;
	wire [4-1:0] node7979;
	wire [4-1:0] node7982;
	wire [4-1:0] node7983;
	wire [4-1:0] node7987;
	wire [4-1:0] node7988;
	wire [4-1:0] node7989;
	wire [4-1:0] node7991;
	wire [4-1:0] node7994;
	wire [4-1:0] node7995;
	wire [4-1:0] node7998;
	wire [4-1:0] node8002;
	wire [4-1:0] node8003;
	wire [4-1:0] node8004;
	wire [4-1:0] node8005;
	wire [4-1:0] node8007;
	wire [4-1:0] node8008;
	wire [4-1:0] node8009;
	wire [4-1:0] node8011;
	wire [4-1:0] node8014;
	wire [4-1:0] node8015;
	wire [4-1:0] node8019;
	wire [4-1:0] node8020;
	wire [4-1:0] node8023;
	wire [4-1:0] node8026;
	wire [4-1:0] node8028;
	wire [4-1:0] node8029;
	wire [4-1:0] node8032;
	wire [4-1:0] node8035;
	wire [4-1:0] node8036;
	wire [4-1:0] node8037;
	wire [4-1:0] node8039;
	wire [4-1:0] node8040;
	wire [4-1:0] node8043;
	wire [4-1:0] node8046;
	wire [4-1:0] node8047;
	wire [4-1:0] node8050;
	wire [4-1:0] node8052;
	wire [4-1:0] node8055;
	wire [4-1:0] node8056;
	wire [4-1:0] node8057;
	wire [4-1:0] node8058;
	wire [4-1:0] node8062;
	wire [4-1:0] node8065;
	wire [4-1:0] node8067;
	wire [4-1:0] node8068;
	wire [4-1:0] node8069;
	wire [4-1:0] node8072;
	wire [4-1:0] node8075;
	wire [4-1:0] node8076;
	wire [4-1:0] node8080;
	wire [4-1:0] node8081;
	wire [4-1:0] node8082;
	wire [4-1:0] node8083;
	wire [4-1:0] node8084;
	wire [4-1:0] node8086;
	wire [4-1:0] node8089;
	wire [4-1:0] node8091;
	wire [4-1:0] node8094;
	wire [4-1:0] node8095;
	wire [4-1:0] node8096;
	wire [4-1:0] node8101;
	wire [4-1:0] node8102;
	wire [4-1:0] node8103;
	wire [4-1:0] node8104;
	wire [4-1:0] node8108;
	wire [4-1:0] node8110;
	wire [4-1:0] node8113;
	wire [4-1:0] node8114;
	wire [4-1:0] node8116;
	wire [4-1:0] node8119;
	wire [4-1:0] node8120;
	wire [4-1:0] node8124;
	wire [4-1:0] node8125;
	wire [4-1:0] node8126;
	wire [4-1:0] node8127;
	wire [4-1:0] node8129;
	wire [4-1:0] node8132;
	wire [4-1:0] node8134;
	wire [4-1:0] node8137;
	wire [4-1:0] node8138;
	wire [4-1:0] node8139;
	wire [4-1:0] node8143;
	wire [4-1:0] node8144;
	wire [4-1:0] node8148;
	wire [4-1:0] node8149;
	wire [4-1:0] node8150;
	wire [4-1:0] node8152;
	wire [4-1:0] node8155;
	wire [4-1:0] node8157;
	wire [4-1:0] node8160;
	wire [4-1:0] node8161;
	wire [4-1:0] node8162;
	wire [4-1:0] node8165;
	wire [4-1:0] node8169;
	wire [4-1:0] node8170;
	wire [4-1:0] node8171;
	wire [4-1:0] node8172;
	wire [4-1:0] node8173;
	wire [4-1:0] node8175;
	wire [4-1:0] node8176;
	wire [4-1:0] node8179;
	wire [4-1:0] node8182;
	wire [4-1:0] node8184;
	wire [4-1:0] node8185;
	wire [4-1:0] node8186;
	wire [4-1:0] node8187;
	wire [4-1:0] node8190;
	wire [4-1:0] node8193;
	wire [4-1:0] node8194;
	wire [4-1:0] node8197;
	wire [4-1:0] node8200;
	wire [4-1:0] node8201;
	wire [4-1:0] node8204;
	wire [4-1:0] node8207;
	wire [4-1:0] node8208;
	wire [4-1:0] node8209;
	wire [4-1:0] node8211;
	wire [4-1:0] node8212;
	wire [4-1:0] node8214;
	wire [4-1:0] node8217;
	wire [4-1:0] node8220;
	wire [4-1:0] node8221;
	wire [4-1:0] node8222;
	wire [4-1:0] node8226;
	wire [4-1:0] node8227;
	wire [4-1:0] node8231;
	wire [4-1:0] node8232;
	wire [4-1:0] node8233;
	wire [4-1:0] node8234;
	wire [4-1:0] node8238;
	wire [4-1:0] node8239;
	wire [4-1:0] node8243;
	wire [4-1:0] node8245;
	wire [4-1:0] node8246;
	wire [4-1:0] node8249;
	wire [4-1:0] node8252;
	wire [4-1:0] node8253;
	wire [4-1:0] node8254;
	wire [4-1:0] node8255;
	wire [4-1:0] node8256;
	wire [4-1:0] node8258;
	wire [4-1:0] node8261;
	wire [4-1:0] node8262;
	wire [4-1:0] node8266;
	wire [4-1:0] node8267;
	wire [4-1:0] node8268;
	wire [4-1:0] node8272;
	wire [4-1:0] node8274;
	wire [4-1:0] node8277;
	wire [4-1:0] node8278;
	wire [4-1:0] node8279;
	wire [4-1:0] node8280;
	wire [4-1:0] node8284;
	wire [4-1:0] node8286;
	wire [4-1:0] node8289;
	wire [4-1:0] node8290;
	wire [4-1:0] node8292;
	wire [4-1:0] node8295;
	wire [4-1:0] node8296;
	wire [4-1:0] node8300;
	wire [4-1:0] node8301;
	wire [4-1:0] node8302;
	wire [4-1:0] node8303;
	wire [4-1:0] node8304;
	wire [4-1:0] node8308;
	wire [4-1:0] node8309;
	wire [4-1:0] node8313;
	wire [4-1:0] node8314;
	wire [4-1:0] node8316;
	wire [4-1:0] node8319;
	wire [4-1:0] node8321;
	wire [4-1:0] node8324;
	wire [4-1:0] node8325;
	wire [4-1:0] node8326;
	wire [4-1:0] node8328;
	wire [4-1:0] node8331;
	wire [4-1:0] node8333;
	wire [4-1:0] node8336;
	wire [4-1:0] node8337;
	wire [4-1:0] node8339;
	wire [4-1:0] node8342;
	wire [4-1:0] node8345;
	wire [4-1:0] node8346;
	wire [4-1:0] node8347;
	wire [4-1:0] node8348;
	wire [4-1:0] node8349;
	wire [4-1:0] node8350;
	wire [4-1:0] node8353;
	wire [4-1:0] node8357;
	wire [4-1:0] node8358;
	wire [4-1:0] node8359;
	wire [4-1:0] node8360;
	wire [4-1:0] node8361;
	wire [4-1:0] node8364;
	wire [4-1:0] node8367;
	wire [4-1:0] node8368;
	wire [4-1:0] node8371;
	wire [4-1:0] node8374;
	wire [4-1:0] node8375;
	wire [4-1:0] node8378;
	wire [4-1:0] node8382;
	wire [4-1:0] node8383;
	wire [4-1:0] node8384;
	wire [4-1:0] node8385;
	wire [4-1:0] node8387;
	wire [4-1:0] node8391;
	wire [4-1:0] node8392;
	wire [4-1:0] node8394;
	wire [4-1:0] node8397;
	wire [4-1:0] node8399;
	wire [4-1:0] node8402;
	wire [4-1:0] node8403;
	wire [4-1:0] node8404;
	wire [4-1:0] node8405;
	wire [4-1:0] node8409;
	wire [4-1:0] node8411;
	wire [4-1:0] node8414;
	wire [4-1:0] node8415;
	wire [4-1:0] node8416;
	wire [4-1:0] node8417;
	wire [4-1:0] node8420;
	wire [4-1:0] node8423;
	wire [4-1:0] node8424;
	wire [4-1:0] node8429;
	wire [4-1:0] node8430;
	wire [4-1:0] node8431;
	wire [4-1:0] node8432;
	wire [4-1:0] node8433;
	wire [4-1:0] node8434;
	wire [4-1:0] node8438;
	wire [4-1:0] node8439;
	wire [4-1:0] node8443;
	wire [4-1:0] node8444;
	wire [4-1:0] node8445;
	wire [4-1:0] node8449;
	wire [4-1:0] node8450;
	wire [4-1:0] node8454;
	wire [4-1:0] node8455;
	wire [4-1:0] node8456;
	wire [4-1:0] node8458;
	wire [4-1:0] node8461;
	wire [4-1:0] node8463;
	wire [4-1:0] node8466;
	wire [4-1:0] node8467;
	wire [4-1:0] node8468;
	wire [4-1:0] node8472;
	wire [4-1:0] node8474;
	wire [4-1:0] node8477;
	wire [4-1:0] node8478;
	wire [4-1:0] node8479;
	wire [4-1:0] node8480;
	wire [4-1:0] node8481;
	wire [4-1:0] node8482;
	wire [4-1:0] node8485;
	wire [4-1:0] node8488;
	wire [4-1:0] node8489;
	wire [4-1:0] node8492;
	wire [4-1:0] node8496;
	wire [4-1:0] node8497;
	wire [4-1:0] node8499;
	wire [4-1:0] node8502;
	wire [4-1:0] node8504;
	wire [4-1:0] node8507;
	wire [4-1:0] node8508;
	wire [4-1:0] node8509;
	wire [4-1:0] node8510;
	wire [4-1:0] node8514;
	wire [4-1:0] node8516;
	wire [4-1:0] node8519;
	wire [4-1:0] node8520;
	wire [4-1:0] node8521;
	wire [4-1:0] node8525;
	wire [4-1:0] node8527;
	wire [4-1:0] node8530;
	wire [4-1:0] node8531;
	wire [4-1:0] node8532;
	wire [4-1:0] node8533;
	wire [4-1:0] node8534;
	wire [4-1:0] node8535;
	wire [4-1:0] node8536;
	wire [4-1:0] node8537;
	wire [4-1:0] node8538;
	wire [4-1:0] node8539;
	wire [4-1:0] node8540;
	wire [4-1:0] node8542;
	wire [4-1:0] node8545;
	wire [4-1:0] node8547;
	wire [4-1:0] node8550;
	wire [4-1:0] node8551;
	wire [4-1:0] node8552;
	wire [4-1:0] node8556;
	wire [4-1:0] node8557;
	wire [4-1:0] node8561;
	wire [4-1:0] node8562;
	wire [4-1:0] node8563;
	wire [4-1:0] node8564;
	wire [4-1:0] node8566;
	wire [4-1:0] node8570;
	wire [4-1:0] node8571;
	wire [4-1:0] node8572;
	wire [4-1:0] node8575;
	wire [4-1:0] node8578;
	wire [4-1:0] node8580;
	wire [4-1:0] node8583;
	wire [4-1:0] node8584;
	wire [4-1:0] node8585;
	wire [4-1:0] node8588;
	wire [4-1:0] node8591;
	wire [4-1:0] node8592;
	wire [4-1:0] node8596;
	wire [4-1:0] node8597;
	wire [4-1:0] node8598;
	wire [4-1:0] node8599;
	wire [4-1:0] node8600;
	wire [4-1:0] node8602;
	wire [4-1:0] node8605;
	wire [4-1:0] node8606;
	wire [4-1:0] node8610;
	wire [4-1:0] node8611;
	wire [4-1:0] node8614;
	wire [4-1:0] node8616;
	wire [4-1:0] node8619;
	wire [4-1:0] node8620;
	wire [4-1:0] node8621;
	wire [4-1:0] node8622;
	wire [4-1:0] node8626;
	wire [4-1:0] node8627;
	wire [4-1:0] node8631;
	wire [4-1:0] node8632;
	wire [4-1:0] node8633;
	wire [4-1:0] node8638;
	wire [4-1:0] node8639;
	wire [4-1:0] node8640;
	wire [4-1:0] node8641;
	wire [4-1:0] node8642;
	wire [4-1:0] node8646;
	wire [4-1:0] node8647;
	wire [4-1:0] node8651;
	wire [4-1:0] node8654;
	wire [4-1:0] node8655;
	wire [4-1:0] node8656;
	wire [4-1:0] node8657;
	wire [4-1:0] node8660;
	wire [4-1:0] node8663;
	wire [4-1:0] node8665;
	wire [4-1:0] node8668;
	wire [4-1:0] node8669;
	wire [4-1:0] node8670;
	wire [4-1:0] node8673;
	wire [4-1:0] node8676;
	wire [4-1:0] node8677;
	wire [4-1:0] node8680;
	wire [4-1:0] node8683;
	wire [4-1:0] node8684;
	wire [4-1:0] node8685;
	wire [4-1:0] node8686;
	wire [4-1:0] node8687;
	wire [4-1:0] node8688;
	wire [4-1:0] node8690;
	wire [4-1:0] node8693;
	wire [4-1:0] node8694;
	wire [4-1:0] node8698;
	wire [4-1:0] node8699;
	wire [4-1:0] node8700;
	wire [4-1:0] node8704;
	wire [4-1:0] node8705;
	wire [4-1:0] node8708;
	wire [4-1:0] node8711;
	wire [4-1:0] node8712;
	wire [4-1:0] node8713;
	wire [4-1:0] node8716;
	wire [4-1:0] node8718;
	wire [4-1:0] node8721;
	wire [4-1:0] node8722;
	wire [4-1:0] node8725;
	wire [4-1:0] node8727;
	wire [4-1:0] node8730;
	wire [4-1:0] node8731;
	wire [4-1:0] node8732;
	wire [4-1:0] node8733;
	wire [4-1:0] node8734;
	wire [4-1:0] node8737;
	wire [4-1:0] node8740;
	wire [4-1:0] node8742;
	wire [4-1:0] node8745;
	wire [4-1:0] node8747;
	wire [4-1:0] node8748;
	wire [4-1:0] node8752;
	wire [4-1:0] node8753;
	wire [4-1:0] node8754;
	wire [4-1:0] node8756;
	wire [4-1:0] node8759;
	wire [4-1:0] node8761;
	wire [4-1:0] node8764;
	wire [4-1:0] node8765;
	wire [4-1:0] node8766;
	wire [4-1:0] node8769;
	wire [4-1:0] node8772;
	wire [4-1:0] node8773;
	wire [4-1:0] node8776;
	wire [4-1:0] node8779;
	wire [4-1:0] node8780;
	wire [4-1:0] node8781;
	wire [4-1:0] node8782;
	wire [4-1:0] node8783;
	wire [4-1:0] node8785;
	wire [4-1:0] node8788;
	wire [4-1:0] node8791;
	wire [4-1:0] node8792;
	wire [4-1:0] node8794;
	wire [4-1:0] node8797;
	wire [4-1:0] node8799;
	wire [4-1:0] node8802;
	wire [4-1:0] node8803;
	wire [4-1:0] node8804;
	wire [4-1:0] node8806;
	wire [4-1:0] node8809;
	wire [4-1:0] node8811;
	wire [4-1:0] node8814;
	wire [4-1:0] node8815;
	wire [4-1:0] node8816;
	wire [4-1:0] node8820;
	wire [4-1:0] node8823;
	wire [4-1:0] node8824;
	wire [4-1:0] node8825;
	wire [4-1:0] node8826;
	wire [4-1:0] node8827;
	wire [4-1:0] node8830;
	wire [4-1:0] node8833;
	wire [4-1:0] node8834;
	wire [4-1:0] node8837;
	wire [4-1:0] node8840;
	wire [4-1:0] node8841;
	wire [4-1:0] node8845;
	wire [4-1:0] node8846;
	wire [4-1:0] node8848;
	wire [4-1:0] node8849;
	wire [4-1:0] node8852;
	wire [4-1:0] node8855;
	wire [4-1:0] node8856;
	wire [4-1:0] node8858;
	wire [4-1:0] node8861;
	wire [4-1:0] node8863;
	wire [4-1:0] node8866;
	wire [4-1:0] node8867;
	wire [4-1:0] node8868;
	wire [4-1:0] node8869;
	wire [4-1:0] node8870;
	wire [4-1:0] node8871;
	wire [4-1:0] node8874;
	wire [4-1:0] node8875;
	wire [4-1:0] node8877;
	wire [4-1:0] node8881;
	wire [4-1:0] node8882;
	wire [4-1:0] node8885;
	wire [4-1:0] node8886;
	wire [4-1:0] node8889;
	wire [4-1:0] node8892;
	wire [4-1:0] node8893;
	wire [4-1:0] node8894;
	wire [4-1:0] node8897;
	wire [4-1:0] node8898;
	wire [4-1:0] node8901;
	wire [4-1:0] node8902;
	wire [4-1:0] node8906;
	wire [4-1:0] node8907;
	wire [4-1:0] node8910;
	wire [4-1:0] node8911;
	wire [4-1:0] node8913;
	wire [4-1:0] node8916;
	wire [4-1:0] node8917;
	wire [4-1:0] node8921;
	wire [4-1:0] node8922;
	wire [4-1:0] node8923;
	wire [4-1:0] node8924;
	wire [4-1:0] node8925;
	wire [4-1:0] node8926;
	wire [4-1:0] node8930;
	wire [4-1:0] node8931;
	wire [4-1:0] node8934;
	wire [4-1:0] node8937;
	wire [4-1:0] node8938;
	wire [4-1:0] node8939;
	wire [4-1:0] node8942;
	wire [4-1:0] node8945;
	wire [4-1:0] node8946;
	wire [4-1:0] node8949;
	wire [4-1:0] node8952;
	wire [4-1:0] node8953;
	wire [4-1:0] node8954;
	wire [4-1:0] node8957;
	wire [4-1:0] node8958;
	wire [4-1:0] node8961;
	wire [4-1:0] node8964;
	wire [4-1:0] node8965;
	wire [4-1:0] node8966;
	wire [4-1:0] node8969;
	wire [4-1:0] node8972;
	wire [4-1:0] node8973;
	wire [4-1:0] node8976;
	wire [4-1:0] node8979;
	wire [4-1:0] node8980;
	wire [4-1:0] node8981;
	wire [4-1:0] node8982;
	wire [4-1:0] node8983;
	wire [4-1:0] node8987;
	wire [4-1:0] node8988;
	wire [4-1:0] node8991;
	wire [4-1:0] node8994;
	wire [4-1:0] node8995;
	wire [4-1:0] node8996;
	wire [4-1:0] node8999;
	wire [4-1:0] node9002;
	wire [4-1:0] node9003;
	wire [4-1:0] node9006;
	wire [4-1:0] node9009;
	wire [4-1:0] node9010;
	wire [4-1:0] node9011;
	wire [4-1:0] node9012;
	wire [4-1:0] node9015;
	wire [4-1:0] node9018;
	wire [4-1:0] node9019;
	wire [4-1:0] node9022;
	wire [4-1:0] node9025;
	wire [4-1:0] node9026;
	wire [4-1:0] node9028;
	wire [4-1:0] node9032;
	wire [4-1:0] node9033;
	wire [4-1:0] node9034;
	wire [4-1:0] node9035;
	wire [4-1:0] node9036;
	wire [4-1:0] node9037;
	wire [4-1:0] node9040;
	wire [4-1:0] node9041;
	wire [4-1:0] node9045;
	wire [4-1:0] node9046;
	wire [4-1:0] node9047;
	wire [4-1:0] node9051;
	wire [4-1:0] node9054;
	wire [4-1:0] node9055;
	wire [4-1:0] node9056;
	wire [4-1:0] node9057;
	wire [4-1:0] node9060;
	wire [4-1:0] node9064;
	wire [4-1:0] node9065;
	wire [4-1:0] node9068;
	wire [4-1:0] node9071;
	wire [4-1:0] node9072;
	wire [4-1:0] node9073;
	wire [4-1:0] node9074;
	wire [4-1:0] node9077;
	wire [4-1:0] node9080;
	wire [4-1:0] node9081;
	wire [4-1:0] node9082;
	wire [4-1:0] node9085;
	wire [4-1:0] node9088;
	wire [4-1:0] node9089;
	wire [4-1:0] node9092;
	wire [4-1:0] node9095;
	wire [4-1:0] node9096;
	wire [4-1:0] node9098;
	wire [4-1:0] node9099;
	wire [4-1:0] node9103;
	wire [4-1:0] node9104;
	wire [4-1:0] node9106;
	wire [4-1:0] node9109;
	wire [4-1:0] node9111;
	wire [4-1:0] node9114;
	wire [4-1:0] node9115;
	wire [4-1:0] node9116;
	wire [4-1:0] node9117;
	wire [4-1:0] node9118;
	wire [4-1:0] node9121;
	wire [4-1:0] node9124;
	wire [4-1:0] node9125;
	wire [4-1:0] node9126;
	wire [4-1:0] node9131;
	wire [4-1:0] node9132;
	wire [4-1:0] node9133;
	wire [4-1:0] node9136;
	wire [4-1:0] node9139;
	wire [4-1:0] node9140;
	wire [4-1:0] node9143;
	wire [4-1:0] node9146;
	wire [4-1:0] node9147;
	wire [4-1:0] node9148;
	wire [4-1:0] node9150;
	wire [4-1:0] node9151;
	wire [4-1:0] node9154;
	wire [4-1:0] node9157;
	wire [4-1:0] node9158;
	wire [4-1:0] node9159;
	wire [4-1:0] node9162;
	wire [4-1:0] node9165;
	wire [4-1:0] node9167;
	wire [4-1:0] node9170;
	wire [4-1:0] node9171;
	wire [4-1:0] node9172;
	wire [4-1:0] node9175;
	wire [4-1:0] node9178;
	wire [4-1:0] node9179;
	wire [4-1:0] node9180;
	wire [4-1:0] node9184;
	wire [4-1:0] node9185;
	wire [4-1:0] node9188;
	wire [4-1:0] node9191;
	wire [4-1:0] node9192;
	wire [4-1:0] node9193;
	wire [4-1:0] node9194;
	wire [4-1:0] node9195;
	wire [4-1:0] node9196;
	wire [4-1:0] node9197;
	wire [4-1:0] node9198;
	wire [4-1:0] node9202;
	wire [4-1:0] node9203;
	wire [4-1:0] node9204;
	wire [4-1:0] node9208;
	wire [4-1:0] node9211;
	wire [4-1:0] node9212;
	wire [4-1:0] node9213;
	wire [4-1:0] node9215;
	wire [4-1:0] node9218;
	wire [4-1:0] node9219;
	wire [4-1:0] node9223;
	wire [4-1:0] node9224;
	wire [4-1:0] node9227;
	wire [4-1:0] node9229;
	wire [4-1:0] node9232;
	wire [4-1:0] node9233;
	wire [4-1:0] node9234;
	wire [4-1:0] node9235;
	wire [4-1:0] node9237;
	wire [4-1:0] node9240;
	wire [4-1:0] node9242;
	wire [4-1:0] node9245;
	wire [4-1:0] node9246;
	wire [4-1:0] node9247;
	wire [4-1:0] node9250;
	wire [4-1:0] node9253;
	wire [4-1:0] node9254;
	wire [4-1:0] node9257;
	wire [4-1:0] node9260;
	wire [4-1:0] node9261;
	wire [4-1:0] node9262;
	wire [4-1:0] node9263;
	wire [4-1:0] node9267;
	wire [4-1:0] node9268;
	wire [4-1:0] node9272;
	wire [4-1:0] node9273;
	wire [4-1:0] node9274;
	wire [4-1:0] node9278;
	wire [4-1:0] node9279;
	wire [4-1:0] node9283;
	wire [4-1:0] node9284;
	wire [4-1:0] node9285;
	wire [4-1:0] node9286;
	wire [4-1:0] node9287;
	wire [4-1:0] node9288;
	wire [4-1:0] node9292;
	wire [4-1:0] node9295;
	wire [4-1:0] node9296;
	wire [4-1:0] node9297;
	wire [4-1:0] node9301;
	wire [4-1:0] node9304;
	wire [4-1:0] node9305;
	wire [4-1:0] node9306;
	wire [4-1:0] node9309;
	wire [4-1:0] node9312;
	wire [4-1:0] node9313;
	wire [4-1:0] node9314;
	wire [4-1:0] node9318;
	wire [4-1:0] node9321;
	wire [4-1:0] node9322;
	wire [4-1:0] node9323;
	wire [4-1:0] node9324;
	wire [4-1:0] node9325;
	wire [4-1:0] node9328;
	wire [4-1:0] node9332;
	wire [4-1:0] node9333;
	wire [4-1:0] node9335;
	wire [4-1:0] node9338;
	wire [4-1:0] node9339;
	wire [4-1:0] node9342;
	wire [4-1:0] node9345;
	wire [4-1:0] node9346;
	wire [4-1:0] node9347;
	wire [4-1:0] node9348;
	wire [4-1:0] node9351;
	wire [4-1:0] node9354;
	wire [4-1:0] node9355;
	wire [4-1:0] node9358;
	wire [4-1:0] node9361;
	wire [4-1:0] node9362;
	wire [4-1:0] node9363;
	wire [4-1:0] node9367;
	wire [4-1:0] node9368;
	wire [4-1:0] node9371;
	wire [4-1:0] node9374;
	wire [4-1:0] node9375;
	wire [4-1:0] node9376;
	wire [4-1:0] node9377;
	wire [4-1:0] node9378;
	wire [4-1:0] node9379;
	wire [4-1:0] node9381;
	wire [4-1:0] node9384;
	wire [4-1:0] node9385;
	wire [4-1:0] node9389;
	wire [4-1:0] node9391;
	wire [4-1:0] node9392;
	wire [4-1:0] node9396;
	wire [4-1:0] node9397;
	wire [4-1:0] node9398;
	wire [4-1:0] node9400;
	wire [4-1:0] node9403;
	wire [4-1:0] node9405;
	wire [4-1:0] node9408;
	wire [4-1:0] node9409;
	wire [4-1:0] node9410;
	wire [4-1:0] node9414;
	wire [4-1:0] node9416;
	wire [4-1:0] node9419;
	wire [4-1:0] node9420;
	wire [4-1:0] node9421;
	wire [4-1:0] node9422;
	wire [4-1:0] node9424;
	wire [4-1:0] node9427;
	wire [4-1:0] node9428;
	wire [4-1:0] node9431;
	wire [4-1:0] node9434;
	wire [4-1:0] node9435;
	wire [4-1:0] node9438;
	wire [4-1:0] node9441;
	wire [4-1:0] node9442;
	wire [4-1:0] node9443;
	wire [4-1:0] node9444;
	wire [4-1:0] node9447;
	wire [4-1:0] node9450;
	wire [4-1:0] node9451;
	wire [4-1:0] node9454;
	wire [4-1:0] node9457;
	wire [4-1:0] node9458;
	wire [4-1:0] node9460;
	wire [4-1:0] node9463;
	wire [4-1:0] node9464;
	wire [4-1:0] node9467;
	wire [4-1:0] node9470;
	wire [4-1:0] node9471;
	wire [4-1:0] node9472;
	wire [4-1:0] node9473;
	wire [4-1:0] node9474;
	wire [4-1:0] node9475;
	wire [4-1:0] node9478;
	wire [4-1:0] node9481;
	wire [4-1:0] node9482;
	wire [4-1:0] node9485;
	wire [4-1:0] node9488;
	wire [4-1:0] node9489;
	wire [4-1:0] node9491;
	wire [4-1:0] node9494;
	wire [4-1:0] node9495;
	wire [4-1:0] node9498;
	wire [4-1:0] node9501;
	wire [4-1:0] node9502;
	wire [4-1:0] node9503;
	wire [4-1:0] node9504;
	wire [4-1:0] node9507;
	wire [4-1:0] node9510;
	wire [4-1:0] node9511;
	wire [4-1:0] node9514;
	wire [4-1:0] node9517;
	wire [4-1:0] node9518;
	wire [4-1:0] node9519;
	wire [4-1:0] node9522;
	wire [4-1:0] node9525;
	wire [4-1:0] node9526;
	wire [4-1:0] node9530;
	wire [4-1:0] node9531;
	wire [4-1:0] node9532;
	wire [4-1:0] node9533;
	wire [4-1:0] node9534;
	wire [4-1:0] node9537;
	wire [4-1:0] node9540;
	wire [4-1:0] node9541;
	wire [4-1:0] node9544;
	wire [4-1:0] node9547;
	wire [4-1:0] node9548;
	wire [4-1:0] node9551;
	wire [4-1:0] node9554;
	wire [4-1:0] node9555;
	wire [4-1:0] node9556;
	wire [4-1:0] node9559;
	wire [4-1:0] node9562;
	wire [4-1:0] node9563;
	wire [4-1:0] node9566;
	wire [4-1:0] node9569;
	wire [4-1:0] node9570;
	wire [4-1:0] node9571;
	wire [4-1:0] node9572;
	wire [4-1:0] node9573;
	wire [4-1:0] node9574;
	wire [4-1:0] node9575;
	wire [4-1:0] node9576;
	wire [4-1:0] node9580;
	wire [4-1:0] node9583;
	wire [4-1:0] node9584;
	wire [4-1:0] node9587;
	wire [4-1:0] node9590;
	wire [4-1:0] node9591;
	wire [4-1:0] node9592;
	wire [4-1:0] node9593;
	wire [4-1:0] node9597;
	wire [4-1:0] node9598;
	wire [4-1:0] node9602;
	wire [4-1:0] node9603;
	wire [4-1:0] node9606;
	wire [4-1:0] node9609;
	wire [4-1:0] node9610;
	wire [4-1:0] node9611;
	wire [4-1:0] node9612;
	wire [4-1:0] node9613;
	wire [4-1:0] node9617;
	wire [4-1:0] node9620;
	wire [4-1:0] node9621;
	wire [4-1:0] node9623;
	wire [4-1:0] node9626;
	wire [4-1:0] node9627;
	wire [4-1:0] node9630;
	wire [4-1:0] node9633;
	wire [4-1:0] node9634;
	wire [4-1:0] node9635;
	wire [4-1:0] node9638;
	wire [4-1:0] node9641;
	wire [4-1:0] node9642;
	wire [4-1:0] node9645;
	wire [4-1:0] node9648;
	wire [4-1:0] node9649;
	wire [4-1:0] node9650;
	wire [4-1:0] node9651;
	wire [4-1:0] node9652;
	wire [4-1:0] node9656;
	wire [4-1:0] node9658;
	wire [4-1:0] node9659;
	wire [4-1:0] node9662;
	wire [4-1:0] node9665;
	wire [4-1:0] node9666;
	wire [4-1:0] node9667;
	wire [4-1:0] node9669;
	wire [4-1:0] node9672;
	wire [4-1:0] node9673;
	wire [4-1:0] node9676;
	wire [4-1:0] node9679;
	wire [4-1:0] node9680;
	wire [4-1:0] node9683;
	wire [4-1:0] node9684;
	wire [4-1:0] node9687;
	wire [4-1:0] node9690;
	wire [4-1:0] node9691;
	wire [4-1:0] node9692;
	wire [4-1:0] node9693;
	wire [4-1:0] node9694;
	wire [4-1:0] node9697;
	wire [4-1:0] node9700;
	wire [4-1:0] node9701;
	wire [4-1:0] node9704;
	wire [4-1:0] node9707;
	wire [4-1:0] node9709;
	wire [4-1:0] node9710;
	wire [4-1:0] node9713;
	wire [4-1:0] node9716;
	wire [4-1:0] node9717;
	wire [4-1:0] node9718;
	wire [4-1:0] node9719;
	wire [4-1:0] node9722;
	wire [4-1:0] node9726;
	wire [4-1:0] node9727;
	wire [4-1:0] node9728;
	wire [4-1:0] node9731;
	wire [4-1:0] node9734;
	wire [4-1:0] node9736;
	wire [4-1:0] node9739;
	wire [4-1:0] node9740;
	wire [4-1:0] node9741;
	wire [4-1:0] node9742;
	wire [4-1:0] node9743;
	wire [4-1:0] node9744;
	wire [4-1:0] node9746;
	wire [4-1:0] node9749;
	wire [4-1:0] node9750;
	wire [4-1:0] node9753;
	wire [4-1:0] node9756;
	wire [4-1:0] node9758;
	wire [4-1:0] node9760;
	wire [4-1:0] node9763;
	wire [4-1:0] node9764;
	wire [4-1:0] node9765;
	wire [4-1:0] node9766;
	wire [4-1:0] node9769;
	wire [4-1:0] node9772;
	wire [4-1:0] node9773;
	wire [4-1:0] node9776;
	wire [4-1:0] node9779;
	wire [4-1:0] node9780;
	wire [4-1:0] node9781;
	wire [4-1:0] node9784;
	wire [4-1:0] node9787;
	wire [4-1:0] node9788;
	wire [4-1:0] node9791;
	wire [4-1:0] node9794;
	wire [4-1:0] node9795;
	wire [4-1:0] node9796;
	wire [4-1:0] node9797;
	wire [4-1:0] node9798;
	wire [4-1:0] node9802;
	wire [4-1:0] node9804;
	wire [4-1:0] node9807;
	wire [4-1:0] node9808;
	wire [4-1:0] node9809;
	wire [4-1:0] node9812;
	wire [4-1:0] node9815;
	wire [4-1:0] node9817;
	wire [4-1:0] node9820;
	wire [4-1:0] node9821;
	wire [4-1:0] node9822;
	wire [4-1:0] node9823;
	wire [4-1:0] node9826;
	wire [4-1:0] node9829;
	wire [4-1:0] node9830;
	wire [4-1:0] node9833;
	wire [4-1:0] node9836;
	wire [4-1:0] node9837;
	wire [4-1:0] node9838;
	wire [4-1:0] node9841;
	wire [4-1:0] node9844;
	wire [4-1:0] node9845;
	wire [4-1:0] node9848;
	wire [4-1:0] node9851;
	wire [4-1:0] node9852;
	wire [4-1:0] node9853;
	wire [4-1:0] node9854;
	wire [4-1:0] node9855;
	wire [4-1:0] node9857;
	wire [4-1:0] node9860;
	wire [4-1:0] node9863;
	wire [4-1:0] node9864;
	wire [4-1:0] node9865;
	wire [4-1:0] node9868;
	wire [4-1:0] node9871;
	wire [4-1:0] node9872;
	wire [4-1:0] node9875;
	wire [4-1:0] node9878;
	wire [4-1:0] node9879;
	wire [4-1:0] node9880;
	wire [4-1:0] node9882;
	wire [4-1:0] node9885;
	wire [4-1:0] node9887;
	wire [4-1:0] node9890;
	wire [4-1:0] node9891;
	wire [4-1:0] node9892;
	wire [4-1:0] node9896;
	wire [4-1:0] node9898;
	wire [4-1:0] node9901;
	wire [4-1:0] node9902;
	wire [4-1:0] node9903;
	wire [4-1:0] node9905;
	wire [4-1:0] node9908;
	wire [4-1:0] node9909;
	wire [4-1:0] node9910;
	wire [4-1:0] node9913;
	wire [4-1:0] node9916;
	wire [4-1:0] node9918;
	wire [4-1:0] node9921;
	wire [4-1:0] node9922;
	wire [4-1:0] node9923;
	wire [4-1:0] node9925;
	wire [4-1:0] node9928;
	wire [4-1:0] node9931;
	wire [4-1:0] node9932;
	wire [4-1:0] node9934;
	wire [4-1:0] node9937;
	wire [4-1:0] node9940;
	wire [4-1:0] node9941;
	wire [4-1:0] node9942;
	wire [4-1:0] node9943;
	wire [4-1:0] node9944;
	wire [4-1:0] node9945;
	wire [4-1:0] node9946;
	wire [4-1:0] node9947;
	wire [4-1:0] node9948;
	wire [4-1:0] node9951;
	wire [4-1:0] node9954;
	wire [4-1:0] node9955;
	wire [4-1:0] node9958;
	wire [4-1:0] node9961;
	wire [4-1:0] node9962;
	wire [4-1:0] node9963;
	wire [4-1:0] node9966;
	wire [4-1:0] node9969;
	wire [4-1:0] node9970;
	wire [4-1:0] node9973;
	wire [4-1:0] node9976;
	wire [4-1:0] node9977;
	wire [4-1:0] node9978;
	wire [4-1:0] node9979;
	wire [4-1:0] node9980;
	wire [4-1:0] node9983;
	wire [4-1:0] node9986;
	wire [4-1:0] node9987;
	wire [4-1:0] node9991;
	wire [4-1:0] node9993;
	wire [4-1:0] node9994;
	wire [4-1:0] node9997;
	wire [4-1:0] node10000;
	wire [4-1:0] node10001;
	wire [4-1:0] node10003;
	wire [4-1:0] node10004;
	wire [4-1:0] node10008;
	wire [4-1:0] node10009;
	wire [4-1:0] node10010;
	wire [4-1:0] node10013;
	wire [4-1:0] node10016;
	wire [4-1:0] node10017;
	wire [4-1:0] node10021;
	wire [4-1:0] node10022;
	wire [4-1:0] node10023;
	wire [4-1:0] node10024;
	wire [4-1:0] node10025;
	wire [4-1:0] node10027;
	wire [4-1:0] node10030;
	wire [4-1:0] node10031;
	wire [4-1:0] node10035;
	wire [4-1:0] node10036;
	wire [4-1:0] node10038;
	wire [4-1:0] node10041;
	wire [4-1:0] node10043;
	wire [4-1:0] node10046;
	wire [4-1:0] node10047;
	wire [4-1:0] node10048;
	wire [4-1:0] node10049;
	wire [4-1:0] node10052;
	wire [4-1:0] node10056;
	wire [4-1:0] node10057;
	wire [4-1:0] node10059;
	wire [4-1:0] node10062;
	wire [4-1:0] node10063;
	wire [4-1:0] node10067;
	wire [4-1:0] node10068;
	wire [4-1:0] node10069;
	wire [4-1:0] node10072;
	wire [4-1:0] node10075;
	wire [4-1:0] node10076;
	wire [4-1:0] node10077;
	wire [4-1:0] node10078;
	wire [4-1:0] node10082;
	wire [4-1:0] node10083;
	wire [4-1:0] node10086;
	wire [4-1:0] node10089;
	wire [4-1:0] node10090;
	wire [4-1:0] node10093;
	wire [4-1:0] node10096;
	wire [4-1:0] node10097;
	wire [4-1:0] node10098;
	wire [4-1:0] node10099;
	wire [4-1:0] node10100;
	wire [4-1:0] node10102;
	wire [4-1:0] node10105;
	wire [4-1:0] node10106;
	wire [4-1:0] node10110;
	wire [4-1:0] node10111;
	wire [4-1:0] node10112;
	wire [4-1:0] node10116;
	wire [4-1:0] node10118;
	wire [4-1:0] node10121;
	wire [4-1:0] node10122;
	wire [4-1:0] node10123;
	wire [4-1:0] node10124;
	wire [4-1:0] node10128;
	wire [4-1:0] node10129;
	wire [4-1:0] node10133;
	wire [4-1:0] node10134;
	wire [4-1:0] node10135;
	wire [4-1:0] node10136;
	wire [4-1:0] node10140;
	wire [4-1:0] node10142;
	wire [4-1:0] node10146;
	wire [4-1:0] node10147;
	wire [4-1:0] node10148;
	wire [4-1:0] node10149;
	wire [4-1:0] node10150;
	wire [4-1:0] node10153;
	wire [4-1:0] node10156;
	wire [4-1:0] node10157;
	wire [4-1:0] node10160;
	wire [4-1:0] node10163;
	wire [4-1:0] node10164;
	wire [4-1:0] node10167;
	wire [4-1:0] node10170;
	wire [4-1:0] node10171;
	wire [4-1:0] node10172;
	wire [4-1:0] node10173;
	wire [4-1:0] node10174;
	wire [4-1:0] node10177;
	wire [4-1:0] node10180;
	wire [4-1:0] node10181;
	wire [4-1:0] node10185;
	wire [4-1:0] node10186;
	wire [4-1:0] node10187;
	wire [4-1:0] node10191;
	wire [4-1:0] node10193;
	wire [4-1:0] node10196;
	wire [4-1:0] node10197;
	wire [4-1:0] node10198;
	wire [4-1:0] node10199;
	wire [4-1:0] node10202;
	wire [4-1:0] node10206;
	wire [4-1:0] node10207;
	wire [4-1:0] node10208;
	wire [4-1:0] node10211;
	wire [4-1:0] node10214;
	wire [4-1:0] node10216;
	wire [4-1:0] node10219;
	wire [4-1:0] node10220;
	wire [4-1:0] node10221;
	wire [4-1:0] node10222;
	wire [4-1:0] node10223;
	wire [4-1:0] node10224;
	wire [4-1:0] node10225;
	wire [4-1:0] node10229;
	wire [4-1:0] node10230;
	wire [4-1:0] node10234;
	wire [4-1:0] node10235;
	wire [4-1:0] node10236;
	wire [4-1:0] node10240;
	wire [4-1:0] node10241;
	wire [4-1:0] node10245;
	wire [4-1:0] node10246;
	wire [4-1:0] node10247;
	wire [4-1:0] node10248;
	wire [4-1:0] node10252;
	wire [4-1:0] node10253;
	wire [4-1:0] node10257;
	wire [4-1:0] node10258;
	wire [4-1:0] node10259;
	wire [4-1:0] node10263;
	wire [4-1:0] node10264;
	wire [4-1:0] node10268;
	wire [4-1:0] node10269;
	wire [4-1:0] node10270;
	wire [4-1:0] node10271;
	wire [4-1:0] node10273;
	wire [4-1:0] node10276;
	wire [4-1:0] node10278;
	wire [4-1:0] node10281;
	wire [4-1:0] node10282;
	wire [4-1:0] node10283;
	wire [4-1:0] node10287;
	wire [4-1:0] node10288;
	wire [4-1:0] node10292;
	wire [4-1:0] node10293;
	wire [4-1:0] node10294;
	wire [4-1:0] node10295;
	wire [4-1:0] node10299;
	wire [4-1:0] node10301;
	wire [4-1:0] node10304;
	wire [4-1:0] node10305;
	wire [4-1:0] node10306;
	wire [4-1:0] node10310;
	wire [4-1:0] node10311;
	wire [4-1:0] node10315;
	wire [4-1:0] node10316;
	wire [4-1:0] node10317;
	wire [4-1:0] node10318;
	wire [4-1:0] node10319;
	wire [4-1:0] node10322;
	wire [4-1:0] node10323;
	wire [4-1:0] node10327;
	wire [4-1:0] node10328;
	wire [4-1:0] node10331;
	wire [4-1:0] node10332;
	wire [4-1:0] node10336;
	wire [4-1:0] node10337;
	wire [4-1:0] node10338;
	wire [4-1:0] node10339;
	wire [4-1:0] node10342;
	wire [4-1:0] node10345;
	wire [4-1:0] node10346;
	wire [4-1:0] node10349;
	wire [4-1:0] node10352;
	wire [4-1:0] node10353;
	wire [4-1:0] node10354;
	wire [4-1:0] node10357;
	wire [4-1:0] node10360;
	wire [4-1:0] node10362;
	wire [4-1:0] node10365;
	wire [4-1:0] node10366;
	wire [4-1:0] node10367;
	wire [4-1:0] node10368;
	wire [4-1:0] node10370;
	wire [4-1:0] node10373;
	wire [4-1:0] node10374;
	wire [4-1:0] node10378;
	wire [4-1:0] node10379;
	wire [4-1:0] node10381;
	wire [4-1:0] node10384;
	wire [4-1:0] node10386;
	wire [4-1:0] node10389;
	wire [4-1:0] node10390;
	wire [4-1:0] node10391;
	wire [4-1:0] node10392;
	wire [4-1:0] node10396;
	wire [4-1:0] node10397;
	wire [4-1:0] node10401;
	wire [4-1:0] node10402;
	wire [4-1:0] node10404;
	wire [4-1:0] node10407;
	wire [4-1:0] node10409;
	wire [4-1:0] node10412;
	wire [4-1:0] node10413;
	wire [4-1:0] node10414;
	wire [4-1:0] node10415;
	wire [4-1:0] node10416;
	wire [4-1:0] node10417;
	wire [4-1:0] node10418;
	wire [4-1:0] node10420;
	wire [4-1:0] node10423;
	wire [4-1:0] node10425;
	wire [4-1:0] node10428;
	wire [4-1:0] node10429;
	wire [4-1:0] node10430;
	wire [4-1:0] node10434;
	wire [4-1:0] node10436;
	wire [4-1:0] node10439;
	wire [4-1:0] node10440;
	wire [4-1:0] node10441;
	wire [4-1:0] node10442;
	wire [4-1:0] node10446;
	wire [4-1:0] node10448;
	wire [4-1:0] node10451;
	wire [4-1:0] node10452;
	wire [4-1:0] node10453;
	wire [4-1:0] node10457;
	wire [4-1:0] node10459;
	wire [4-1:0] node10462;
	wire [4-1:0] node10463;
	wire [4-1:0] node10464;
	wire [4-1:0] node10465;
	wire [4-1:0] node10467;
	wire [4-1:0] node10470;
	wire [4-1:0] node10472;
	wire [4-1:0] node10475;
	wire [4-1:0] node10476;
	wire [4-1:0] node10478;
	wire [4-1:0] node10482;
	wire [4-1:0] node10483;
	wire [4-1:0] node10484;
	wire [4-1:0] node10487;
	wire [4-1:0] node10490;
	wire [4-1:0] node10491;
	wire [4-1:0] node10492;
	wire [4-1:0] node10493;
	wire [4-1:0] node10497;
	wire [4-1:0] node10498;
	wire [4-1:0] node10501;
	wire [4-1:0] node10504;
	wire [4-1:0] node10505;
	wire [4-1:0] node10506;
	wire [4-1:0] node10509;
	wire [4-1:0] node10512;
	wire [4-1:0] node10513;
	wire [4-1:0] node10516;
	wire [4-1:0] node10519;
	wire [4-1:0] node10520;
	wire [4-1:0] node10521;
	wire [4-1:0] node10522;
	wire [4-1:0] node10523;
	wire [4-1:0] node10524;
	wire [4-1:0] node10528;
	wire [4-1:0] node10529;
	wire [4-1:0] node10533;
	wire [4-1:0] node10534;
	wire [4-1:0] node10535;
	wire [4-1:0] node10539;
	wire [4-1:0] node10541;
	wire [4-1:0] node10544;
	wire [4-1:0] node10545;
	wire [4-1:0] node10547;
	wire [4-1:0] node10548;
	wire [4-1:0] node10552;
	wire [4-1:0] node10553;
	wire [4-1:0] node10554;
	wire [4-1:0] node10558;
	wire [4-1:0] node10559;
	wire [4-1:0] node10563;
	wire [4-1:0] node10564;
	wire [4-1:0] node10565;
	wire [4-1:0] node10567;
	wire [4-1:0] node10568;
	wire [4-1:0] node10569;
	wire [4-1:0] node10572;
	wire [4-1:0] node10575;
	wire [4-1:0] node10576;
	wire [4-1:0] node10580;
	wire [4-1:0] node10582;
	wire [4-1:0] node10583;
	wire [4-1:0] node10586;
	wire [4-1:0] node10589;
	wire [4-1:0] node10590;
	wire [4-1:0] node10592;
	wire [4-1:0] node10593;
	wire [4-1:0] node10596;
	wire [4-1:0] node10599;
	wire [4-1:0] node10601;
	wire [4-1:0] node10602;
	wire [4-1:0] node10603;
	wire [4-1:0] node10606;
	wire [4-1:0] node10609;
	wire [4-1:0] node10610;
	wire [4-1:0] node10613;
	wire [4-1:0] node10616;
	wire [4-1:0] node10617;
	wire [4-1:0] node10618;
	wire [4-1:0] node10619;
	wire [4-1:0] node10620;
	wire [4-1:0] node10621;
	wire [4-1:0] node10622;
	wire [4-1:0] node10623;
	wire [4-1:0] node10626;
	wire [4-1:0] node10629;
	wire [4-1:0] node10630;
	wire [4-1:0] node10633;
	wire [4-1:0] node10636;
	wire [4-1:0] node10637;
	wire [4-1:0] node10639;
	wire [4-1:0] node10642;
	wire [4-1:0] node10643;
	wire [4-1:0] node10646;
	wire [4-1:0] node10649;
	wire [4-1:0] node10650;
	wire [4-1:0] node10651;
	wire [4-1:0] node10653;
	wire [4-1:0] node10656;
	wire [4-1:0] node10657;
	wire [4-1:0] node10661;
	wire [4-1:0] node10662;
	wire [4-1:0] node10663;
	wire [4-1:0] node10666;
	wire [4-1:0] node10669;
	wire [4-1:0] node10670;
	wire [4-1:0] node10673;
	wire [4-1:0] node10676;
	wire [4-1:0] node10677;
	wire [4-1:0] node10678;
	wire [4-1:0] node10680;
	wire [4-1:0] node10683;
	wire [4-1:0] node10685;
	wire [4-1:0] node10688;
	wire [4-1:0] node10689;
	wire [4-1:0] node10690;
	wire [4-1:0] node10694;
	wire [4-1:0] node10696;
	wire [4-1:0] node10699;
	wire [4-1:0] node10700;
	wire [4-1:0] node10701;
	wire [4-1:0] node10704;
	wire [4-1:0] node10707;
	wire [4-1:0] node10708;
	wire [4-1:0] node10709;
	wire [4-1:0] node10710;
	wire [4-1:0] node10712;
	wire [4-1:0] node10715;
	wire [4-1:0] node10717;
	wire [4-1:0] node10720;
	wire [4-1:0] node10722;
	wire [4-1:0] node10723;
	wire [4-1:0] node10726;
	wire [4-1:0] node10729;
	wire [4-1:0] node10730;
	wire [4-1:0] node10731;
	wire [4-1:0] node10732;
	wire [4-1:0] node10736;
	wire [4-1:0] node10737;
	wire [4-1:0] node10740;
	wire [4-1:0] node10743;
	wire [4-1:0] node10744;
	wire [4-1:0] node10745;
	wire [4-1:0] node10748;
	wire [4-1:0] node10751;
	wire [4-1:0] node10752;
	wire [4-1:0] node10755;
	wire [4-1:0] node10758;
	wire [4-1:0] node10759;
	wire [4-1:0] node10760;
	wire [4-1:0] node10761;
	wire [4-1:0] node10763;
	wire [4-1:0] node10766;
	wire [4-1:0] node10768;
	wire [4-1:0] node10771;
	wire [4-1:0] node10772;
	wire [4-1:0] node10773;
	wire [4-1:0] node10777;
	wire [4-1:0] node10778;
	wire [4-1:0] node10782;
	wire [4-1:0] node10783;
	wire [4-1:0] node10784;
	wire [4-1:0] node10787;
	wire [4-1:0] node10790;
	wire [4-1:0] node10791;
	wire [4-1:0] node10792;
	wire [4-1:0] node10793;
	wire [4-1:0] node10796;
	wire [4-1:0] node10800;
	wire [4-1:0] node10801;
	wire [4-1:0] node10802;
	wire [4-1:0] node10804;
	wire [4-1:0] node10807;
	wire [4-1:0] node10808;
	wire [4-1:0] node10812;
	wire [4-1:0] node10813;
	wire [4-1:0] node10816;
	wire [4-1:0] node10819;
	wire [4-1:0] node10820;
	wire [4-1:0] node10821;
	wire [4-1:0] node10822;
	wire [4-1:0] node10823;
	wire [4-1:0] node10824;
	wire [4-1:0] node10825;
	wire [4-1:0] node10826;
	wire [4-1:0] node10827;
	wire [4-1:0] node10828;
	wire [4-1:0] node10829;
	wire [4-1:0] node10832;
	wire [4-1:0] node10835;
	wire [4-1:0] node10836;
	wire [4-1:0] node10839;
	wire [4-1:0] node10843;
	wire [4-1:0] node10844;
	wire [4-1:0] node10846;
	wire [4-1:0] node10847;
	wire [4-1:0] node10850;
	wire [4-1:0] node10853;
	wire [4-1:0] node10854;
	wire [4-1:0] node10855;
	wire [4-1:0] node10859;
	wire [4-1:0] node10861;
	wire [4-1:0] node10864;
	wire [4-1:0] node10865;
	wire [4-1:0] node10866;
	wire [4-1:0] node10867;
	wire [4-1:0] node10868;
	wire [4-1:0] node10871;
	wire [4-1:0] node10874;
	wire [4-1:0] node10875;
	wire [4-1:0] node10879;
	wire [4-1:0] node10880;
	wire [4-1:0] node10882;
	wire [4-1:0] node10885;
	wire [4-1:0] node10886;
	wire [4-1:0] node10889;
	wire [4-1:0] node10892;
	wire [4-1:0] node10893;
	wire [4-1:0] node10894;
	wire [4-1:0] node10896;
	wire [4-1:0] node10899;
	wire [4-1:0] node10901;
	wire [4-1:0] node10904;
	wire [4-1:0] node10905;
	wire [4-1:0] node10908;
	wire [4-1:0] node10910;
	wire [4-1:0] node10913;
	wire [4-1:0] node10914;
	wire [4-1:0] node10915;
	wire [4-1:0] node10916;
	wire [4-1:0] node10918;
	wire [4-1:0] node10921;
	wire [4-1:0] node10922;
	wire [4-1:0] node10923;
	wire [4-1:0] node10927;
	wire [4-1:0] node10929;
	wire [4-1:0] node10932;
	wire [4-1:0] node10933;
	wire [4-1:0] node10934;
	wire [4-1:0] node10937;
	wire [4-1:0] node10940;
	wire [4-1:0] node10941;
	wire [4-1:0] node10945;
	wire [4-1:0] node10946;
	wire [4-1:0] node10947;
	wire [4-1:0] node10948;
	wire [4-1:0] node10951;
	wire [4-1:0] node10954;
	wire [4-1:0] node10956;
	wire [4-1:0] node10957;
	wire [4-1:0] node10960;
	wire [4-1:0] node10963;
	wire [4-1:0] node10964;
	wire [4-1:0] node10965;
	wire [4-1:0] node10967;
	wire [4-1:0] node10970;
	wire [4-1:0] node10972;
	wire [4-1:0] node10975;
	wire [4-1:0] node10976;
	wire [4-1:0] node10978;
	wire [4-1:0] node10981;
	wire [4-1:0] node10983;
	wire [4-1:0] node10986;
	wire [4-1:0] node10987;
	wire [4-1:0] node10988;
	wire [4-1:0] node10989;
	wire [4-1:0] node10990;
	wire [4-1:0] node10991;
	wire [4-1:0] node10992;
	wire [4-1:0] node10996;
	wire [4-1:0] node10999;
	wire [4-1:0] node11000;
	wire [4-1:0] node11003;
	wire [4-1:0] node11004;
	wire [4-1:0] node11008;
	wire [4-1:0] node11009;
	wire [4-1:0] node11010;
	wire [4-1:0] node11013;
	wire [4-1:0] node11014;
	wire [4-1:0] node11018;
	wire [4-1:0] node11020;
	wire [4-1:0] node11023;
	wire [4-1:0] node11024;
	wire [4-1:0] node11025;
	wire [4-1:0] node11026;
	wire [4-1:0] node11028;
	wire [4-1:0] node11031;
	wire [4-1:0] node11033;
	wire [4-1:0] node11036;
	wire [4-1:0] node11037;
	wire [4-1:0] node11040;
	wire [4-1:0] node11042;
	wire [4-1:0] node11045;
	wire [4-1:0] node11046;
	wire [4-1:0] node11047;
	wire [4-1:0] node11048;
	wire [4-1:0] node11051;
	wire [4-1:0] node11054;
	wire [4-1:0] node11055;
	wire [4-1:0] node11058;
	wire [4-1:0] node11061;
	wire [4-1:0] node11062;
	wire [4-1:0] node11063;
	wire [4-1:0] node11066;
	wire [4-1:0] node11069;
	wire [4-1:0] node11070;
	wire [4-1:0] node11073;
	wire [4-1:0] node11076;
	wire [4-1:0] node11077;
	wire [4-1:0] node11078;
	wire [4-1:0] node11079;
	wire [4-1:0] node11080;
	wire [4-1:0] node11081;
	wire [4-1:0] node11085;
	wire [4-1:0] node11087;
	wire [4-1:0] node11090;
	wire [4-1:0] node11091;
	wire [4-1:0] node11092;
	wire [4-1:0] node11096;
	wire [4-1:0] node11097;
	wire [4-1:0] node11101;
	wire [4-1:0] node11102;
	wire [4-1:0] node11103;
	wire [4-1:0] node11105;
	wire [4-1:0] node11108;
	wire [4-1:0] node11111;
	wire [4-1:0] node11112;
	wire [4-1:0] node11115;
	wire [4-1:0] node11117;
	wire [4-1:0] node11120;
	wire [4-1:0] node11121;
	wire [4-1:0] node11122;
	wire [4-1:0] node11123;
	wire [4-1:0] node11125;
	wire [4-1:0] node11128;
	wire [4-1:0] node11129;
	wire [4-1:0] node11132;
	wire [4-1:0] node11135;
	wire [4-1:0] node11136;
	wire [4-1:0] node11139;
	wire [4-1:0] node11140;
	wire [4-1:0] node11143;
	wire [4-1:0] node11146;
	wire [4-1:0] node11147;
	wire [4-1:0] node11150;
	wire [4-1:0] node11151;
	wire [4-1:0] node11154;
	wire [4-1:0] node11157;
	wire [4-1:0] node11158;
	wire [4-1:0] node11159;
	wire [4-1:0] node11160;
	wire [4-1:0] node11161;
	wire [4-1:0] node11162;
	wire [4-1:0] node11163;
	wire [4-1:0] node11164;
	wire [4-1:0] node11167;
	wire [4-1:0] node11170;
	wire [4-1:0] node11171;
	wire [4-1:0] node11174;
	wire [4-1:0] node11177;
	wire [4-1:0] node11178;
	wire [4-1:0] node11181;
	wire [4-1:0] node11184;
	wire [4-1:0] node11185;
	wire [4-1:0] node11186;
	wire [4-1:0] node11187;
	wire [4-1:0] node11192;
	wire [4-1:0] node11193;
	wire [4-1:0] node11197;
	wire [4-1:0] node11198;
	wire [4-1:0] node11199;
	wire [4-1:0] node11200;
	wire [4-1:0] node11201;
	wire [4-1:0] node11205;
	wire [4-1:0] node11207;
	wire [4-1:0] node11210;
	wire [4-1:0] node11211;
	wire [4-1:0] node11213;
	wire [4-1:0] node11216;
	wire [4-1:0] node11217;
	wire [4-1:0] node11221;
	wire [4-1:0] node11222;
	wire [4-1:0] node11223;
	wire [4-1:0] node11224;
	wire [4-1:0] node11228;
	wire [4-1:0] node11230;
	wire [4-1:0] node11233;
	wire [4-1:0] node11234;
	wire [4-1:0] node11235;
	wire [4-1:0] node11240;
	wire [4-1:0] node11241;
	wire [4-1:0] node11242;
	wire [4-1:0] node11243;
	wire [4-1:0] node11244;
	wire [4-1:0] node11248;
	wire [4-1:0] node11249;
	wire [4-1:0] node11253;
	wire [4-1:0] node11254;
	wire [4-1:0] node11256;
	wire [4-1:0] node11259;
	wire [4-1:0] node11261;
	wire [4-1:0] node11264;
	wire [4-1:0] node11265;
	wire [4-1:0] node11266;
	wire [4-1:0] node11269;
	wire [4-1:0] node11272;
	wire [4-1:0] node11273;
	wire [4-1:0] node11274;
	wire [4-1:0] node11277;
	wire [4-1:0] node11280;
	wire [4-1:0] node11281;
	wire [4-1:0] node11282;
	wire [4-1:0] node11285;
	wire [4-1:0] node11288;
	wire [4-1:0] node11289;
	wire [4-1:0] node11293;
	wire [4-1:0] node11294;
	wire [4-1:0] node11295;
	wire [4-1:0] node11296;
	wire [4-1:0] node11297;
	wire [4-1:0] node11298;
	wire [4-1:0] node11301;
	wire [4-1:0] node11304;
	wire [4-1:0] node11305;
	wire [4-1:0] node11306;
	wire [4-1:0] node11309;
	wire [4-1:0] node11312;
	wire [4-1:0] node11314;
	wire [4-1:0] node11317;
	wire [4-1:0] node11318;
	wire [4-1:0] node11319;
	wire [4-1:0] node11321;
	wire [4-1:0] node11324;
	wire [4-1:0] node11327;
	wire [4-1:0] node11328;
	wire [4-1:0] node11329;
	wire [4-1:0] node11333;
	wire [4-1:0] node11336;
	wire [4-1:0] node11337;
	wire [4-1:0] node11338;
	wire [4-1:0] node11340;
	wire [4-1:0] node11341;
	wire [4-1:0] node11345;
	wire [4-1:0] node11346;
	wire [4-1:0] node11348;
	wire [4-1:0] node11351;
	wire [4-1:0] node11352;
	wire [4-1:0] node11356;
	wire [4-1:0] node11358;
	wire [4-1:0] node11359;
	wire [4-1:0] node11361;
	wire [4-1:0] node11364;
	wire [4-1:0] node11367;
	wire [4-1:0] node11368;
	wire [4-1:0] node11369;
	wire [4-1:0] node11370;
	wire [4-1:0] node11373;
	wire [4-1:0] node11376;
	wire [4-1:0] node11377;
	wire [4-1:0] node11378;
	wire [4-1:0] node11381;
	wire [4-1:0] node11384;
	wire [4-1:0] node11385;
	wire [4-1:0] node11386;
	wire [4-1:0] node11389;
	wire [4-1:0] node11392;
	wire [4-1:0] node11393;
	wire [4-1:0] node11396;
	wire [4-1:0] node11399;
	wire [4-1:0] node11400;
	wire [4-1:0] node11401;
	wire [4-1:0] node11402;
	wire [4-1:0] node11405;
	wire [4-1:0] node11408;
	wire [4-1:0] node11410;
	wire [4-1:0] node11411;
	wire [4-1:0] node11414;
	wire [4-1:0] node11417;
	wire [4-1:0] node11418;
	wire [4-1:0] node11419;
	wire [4-1:0] node11420;
	wire [4-1:0] node11423;
	wire [4-1:0] node11426;
	wire [4-1:0] node11427;
	wire [4-1:0] node11431;
	wire [4-1:0] node11432;
	wire [4-1:0] node11435;
	wire [4-1:0] node11438;
	wire [4-1:0] node11439;
	wire [4-1:0] node11440;
	wire [4-1:0] node11441;
	wire [4-1:0] node11442;
	wire [4-1:0] node11443;
	wire [4-1:0] node11444;
	wire [4-1:0] node11445;
	wire [4-1:0] node11447;
	wire [4-1:0] node11450;
	wire [4-1:0] node11451;
	wire [4-1:0] node11455;
	wire [4-1:0] node11456;
	wire [4-1:0] node11458;
	wire [4-1:0] node11461;
	wire [4-1:0] node11463;
	wire [4-1:0] node11466;
	wire [4-1:0] node11467;
	wire [4-1:0] node11468;
	wire [4-1:0] node11470;
	wire [4-1:0] node11473;
	wire [4-1:0] node11474;
	wire [4-1:0] node11478;
	wire [4-1:0] node11479;
	wire [4-1:0] node11481;
	wire [4-1:0] node11484;
	wire [4-1:0] node11486;
	wire [4-1:0] node11489;
	wire [4-1:0] node11490;
	wire [4-1:0] node11491;
	wire [4-1:0] node11492;
	wire [4-1:0] node11493;
	wire [4-1:0] node11497;
	wire [4-1:0] node11498;
	wire [4-1:0] node11502;
	wire [4-1:0] node11503;
	wire [4-1:0] node11506;
	wire [4-1:0] node11507;
	wire [4-1:0] node11511;
	wire [4-1:0] node11512;
	wire [4-1:0] node11513;
	wire [4-1:0] node11516;
	wire [4-1:0] node11519;
	wire [4-1:0] node11520;
	wire [4-1:0] node11521;
	wire [4-1:0] node11524;
	wire [4-1:0] node11527;
	wire [4-1:0] node11528;
	wire [4-1:0] node11531;
	wire [4-1:0] node11534;
	wire [4-1:0] node11535;
	wire [4-1:0] node11536;
	wire [4-1:0] node11537;
	wire [4-1:0] node11538;
	wire [4-1:0] node11541;
	wire [4-1:0] node11544;
	wire [4-1:0] node11545;
	wire [4-1:0] node11546;
	wire [4-1:0] node11549;
	wire [4-1:0] node11552;
	wire [4-1:0] node11553;
	wire [4-1:0] node11557;
	wire [4-1:0] node11558;
	wire [4-1:0] node11559;
	wire [4-1:0] node11560;
	wire [4-1:0] node11564;
	wire [4-1:0] node11565;
	wire [4-1:0] node11568;
	wire [4-1:0] node11571;
	wire [4-1:0] node11572;
	wire [4-1:0] node11575;
	wire [4-1:0] node11578;
	wire [4-1:0] node11579;
	wire [4-1:0] node11580;
	wire [4-1:0] node11581;
	wire [4-1:0] node11584;
	wire [4-1:0] node11587;
	wire [4-1:0] node11588;
	wire [4-1:0] node11589;
	wire [4-1:0] node11592;
	wire [4-1:0] node11595;
	wire [4-1:0] node11597;
	wire [4-1:0] node11600;
	wire [4-1:0] node11601;
	wire [4-1:0] node11603;
	wire [4-1:0] node11605;
	wire [4-1:0] node11608;
	wire [4-1:0] node11609;
	wire [4-1:0] node11612;
	wire [4-1:0] node11615;
	wire [4-1:0] node11616;
	wire [4-1:0] node11617;
	wire [4-1:0] node11618;
	wire [4-1:0] node11619;
	wire [4-1:0] node11620;
	wire [4-1:0] node11622;
	wire [4-1:0] node11625;
	wire [4-1:0] node11626;
	wire [4-1:0] node11629;
	wire [4-1:0] node11632;
	wire [4-1:0] node11633;
	wire [4-1:0] node11635;
	wire [4-1:0] node11638;
	wire [4-1:0] node11639;
	wire [4-1:0] node11642;
	wire [4-1:0] node11645;
	wire [4-1:0] node11646;
	wire [4-1:0] node11647;
	wire [4-1:0] node11650;
	wire [4-1:0] node11653;
	wire [4-1:0] node11654;
	wire [4-1:0] node11655;
	wire [4-1:0] node11659;
	wire [4-1:0] node11660;
	wire [4-1:0] node11663;
	wire [4-1:0] node11666;
	wire [4-1:0] node11667;
	wire [4-1:0] node11668;
	wire [4-1:0] node11669;
	wire [4-1:0] node11670;
	wire [4-1:0] node11673;
	wire [4-1:0] node11676;
	wire [4-1:0] node11677;
	wire [4-1:0] node11680;
	wire [4-1:0] node11683;
	wire [4-1:0] node11684;
	wire [4-1:0] node11687;
	wire [4-1:0] node11690;
	wire [4-1:0] node11691;
	wire [4-1:0] node11692;
	wire [4-1:0] node11693;
	wire [4-1:0] node11697;
	wire [4-1:0] node11698;
	wire [4-1:0] node11702;
	wire [4-1:0] node11704;
	wire [4-1:0] node11707;
	wire [4-1:0] node11708;
	wire [4-1:0] node11709;
	wire [4-1:0] node11710;
	wire [4-1:0] node11711;
	wire [4-1:0] node11712;
	wire [4-1:0] node11715;
	wire [4-1:0] node11718;
	wire [4-1:0] node11719;
	wire [4-1:0] node11722;
	wire [4-1:0] node11725;
	wire [4-1:0] node11726;
	wire [4-1:0] node11729;
	wire [4-1:0] node11732;
	wire [4-1:0] node11733;
	wire [4-1:0] node11734;
	wire [4-1:0] node11735;
	wire [4-1:0] node11738;
	wire [4-1:0] node11741;
	wire [4-1:0] node11742;
	wire [4-1:0] node11745;
	wire [4-1:0] node11748;
	wire [4-1:0] node11749;
	wire [4-1:0] node11752;
	wire [4-1:0] node11755;
	wire [4-1:0] node11756;
	wire [4-1:0] node11757;
	wire [4-1:0] node11758;
	wire [4-1:0] node11762;
	wire [4-1:0] node11765;
	wire [4-1:0] node11766;
	wire [4-1:0] node11768;
	wire [4-1:0] node11771;
	wire [4-1:0] node11773;
	wire [4-1:0] node11776;
	wire [4-1:0] node11777;
	wire [4-1:0] node11778;
	wire [4-1:0] node11779;
	wire [4-1:0] node11780;
	wire [4-1:0] node11781;
	wire [4-1:0] node11782;
	wire [4-1:0] node11784;
	wire [4-1:0] node11787;
	wire [4-1:0] node11788;
	wire [4-1:0] node11791;
	wire [4-1:0] node11794;
	wire [4-1:0] node11795;
	wire [4-1:0] node11798;
	wire [4-1:0] node11801;
	wire [4-1:0] node11802;
	wire [4-1:0] node11803;
	wire [4-1:0] node11804;
	wire [4-1:0] node11809;
	wire [4-1:0] node11810;
	wire [4-1:0] node11814;
	wire [4-1:0] node11815;
	wire [4-1:0] node11816;
	wire [4-1:0] node11817;
	wire [4-1:0] node11818;
	wire [4-1:0] node11822;
	wire [4-1:0] node11824;
	wire [4-1:0] node11827;
	wire [4-1:0] node11828;
	wire [4-1:0] node11830;
	wire [4-1:0] node11833;
	wire [4-1:0] node11834;
	wire [4-1:0] node11838;
	wire [4-1:0] node11839;
	wire [4-1:0] node11840;
	wire [4-1:0] node11842;
	wire [4-1:0] node11845;
	wire [4-1:0] node11846;
	wire [4-1:0] node11850;
	wire [4-1:0] node11851;
	wire [4-1:0] node11852;
	wire [4-1:0] node11856;
	wire [4-1:0] node11857;
	wire [4-1:0] node11861;
	wire [4-1:0] node11862;
	wire [4-1:0] node11863;
	wire [4-1:0] node11864;
	wire [4-1:0] node11865;
	wire [4-1:0] node11867;
	wire [4-1:0] node11870;
	wire [4-1:0] node11871;
	wire [4-1:0] node11874;
	wire [4-1:0] node11877;
	wire [4-1:0] node11878;
	wire [4-1:0] node11879;
	wire [4-1:0] node11882;
	wire [4-1:0] node11885;
	wire [4-1:0] node11886;
	wire [4-1:0] node11890;
	wire [4-1:0] node11891;
	wire [4-1:0] node11892;
	wire [4-1:0] node11893;
	wire [4-1:0] node11896;
	wire [4-1:0] node11899;
	wire [4-1:0] node11900;
	wire [4-1:0] node11903;
	wire [4-1:0] node11906;
	wire [4-1:0] node11907;
	wire [4-1:0] node11908;
	wire [4-1:0] node11911;
	wire [4-1:0] node11914;
	wire [4-1:0] node11915;
	wire [4-1:0] node11918;
	wire [4-1:0] node11921;
	wire [4-1:0] node11922;
	wire [4-1:0] node11923;
	wire [4-1:0] node11924;
	wire [4-1:0] node11925;
	wire [4-1:0] node11928;
	wire [4-1:0] node11931;
	wire [4-1:0] node11932;
	wire [4-1:0] node11935;
	wire [4-1:0] node11938;
	wire [4-1:0] node11940;
	wire [4-1:0] node11942;
	wire [4-1:0] node11945;
	wire [4-1:0] node11946;
	wire [4-1:0] node11947;
	wire [4-1:0] node11948;
	wire [4-1:0] node11952;
	wire [4-1:0] node11953;
	wire [4-1:0] node11957;
	wire [4-1:0] node11958;
	wire [4-1:0] node11960;
	wire [4-1:0] node11963;
	wire [4-1:0] node11964;
	wire [4-1:0] node11967;
	wire [4-1:0] node11970;
	wire [4-1:0] node11971;
	wire [4-1:0] node11972;
	wire [4-1:0] node11973;
	wire [4-1:0] node11974;
	wire [4-1:0] node11975;
	wire [4-1:0] node11976;
	wire [4-1:0] node11980;
	wire [4-1:0] node11983;
	wire [4-1:0] node11984;
	wire [4-1:0] node11985;
	wire [4-1:0] node11990;
	wire [4-1:0] node11991;
	wire [4-1:0] node11993;
	wire [4-1:0] node11994;
	wire [4-1:0] node11998;
	wire [4-1:0] node11999;
	wire [4-1:0] node12000;
	wire [4-1:0] node12004;
	wire [4-1:0] node12006;
	wire [4-1:0] node12009;
	wire [4-1:0] node12010;
	wire [4-1:0] node12011;
	wire [4-1:0] node12013;
	wire [4-1:0] node12016;
	wire [4-1:0] node12017;
	wire [4-1:0] node12019;
	wire [4-1:0] node12022;
	wire [4-1:0] node12023;
	wire [4-1:0] node12027;
	wire [4-1:0] node12028;
	wire [4-1:0] node12029;
	wire [4-1:0] node12032;
	wire [4-1:0] node12035;
	wire [4-1:0] node12036;
	wire [4-1:0] node12037;
	wire [4-1:0] node12042;
	wire [4-1:0] node12043;
	wire [4-1:0] node12044;
	wire [4-1:0] node12045;
	wire [4-1:0] node12049;
	wire [4-1:0] node12051;
	wire [4-1:0] node12054;
	wire [4-1:0] node12055;
	wire [4-1:0] node12057;
	wire [4-1:0] node12060;
	wire [4-1:0] node12061;
	wire [4-1:0] node12065;
	wire [4-1:0] node12066;
	wire [4-1:0] node12067;
	wire [4-1:0] node12068;
	wire [4-1:0] node12069;
	wire [4-1:0] node12070;
	wire [4-1:0] node12071;
	wire [4-1:0] node12072;
	wire [4-1:0] node12074;
	wire [4-1:0] node12075;
	wire [4-1:0] node12078;
	wire [4-1:0] node12081;
	wire [4-1:0] node12082;
	wire [4-1:0] node12084;
	wire [4-1:0] node12087;
	wire [4-1:0] node12088;
	wire [4-1:0] node12091;
	wire [4-1:0] node12094;
	wire [4-1:0] node12095;
	wire [4-1:0] node12098;
	wire [4-1:0] node12101;
	wire [4-1:0] node12102;
	wire [4-1:0] node12103;
	wire [4-1:0] node12104;
	wire [4-1:0] node12108;
	wire [4-1:0] node12111;
	wire [4-1:0] node12112;
	wire [4-1:0] node12113;
	wire [4-1:0] node12117;
	wire [4-1:0] node12118;
	wire [4-1:0] node12122;
	wire [4-1:0] node12123;
	wire [4-1:0] node12124;
	wire [4-1:0] node12125;
	wire [4-1:0] node12126;
	wire [4-1:0] node12130;
	wire [4-1:0] node12132;
	wire [4-1:0] node12135;
	wire [4-1:0] node12136;
	wire [4-1:0] node12138;
	wire [4-1:0] node12141;
	wire [4-1:0] node12143;
	wire [4-1:0] node12146;
	wire [4-1:0] node12147;
	wire [4-1:0] node12148;
	wire [4-1:0] node12149;
	wire [4-1:0] node12151;
	wire [4-1:0] node12154;
	wire [4-1:0] node12155;
	wire [4-1:0] node12159;
	wire [4-1:0] node12160;
	wire [4-1:0] node12164;
	wire [4-1:0] node12165;
	wire [4-1:0] node12166;
	wire [4-1:0] node12167;
	wire [4-1:0] node12171;
	wire [4-1:0] node12173;
	wire [4-1:0] node12176;
	wire [4-1:0] node12177;
	wire [4-1:0] node12179;
	wire [4-1:0] node12182;
	wire [4-1:0] node12183;
	wire [4-1:0] node12187;
	wire [4-1:0] node12188;
	wire [4-1:0] node12189;
	wire [4-1:0] node12190;
	wire [4-1:0] node12191;
	wire [4-1:0] node12193;
	wire [4-1:0] node12196;
	wire [4-1:0] node12198;
	wire [4-1:0] node12201;
	wire [4-1:0] node12202;
	wire [4-1:0] node12204;
	wire [4-1:0] node12207;
	wire [4-1:0] node12209;
	wire [4-1:0] node12212;
	wire [4-1:0] node12213;
	wire [4-1:0] node12214;
	wire [4-1:0] node12215;
	wire [4-1:0] node12219;
	wire [4-1:0] node12220;
	wire [4-1:0] node12224;
	wire [4-1:0] node12225;
	wire [4-1:0] node12226;
	wire [4-1:0] node12230;
	wire [4-1:0] node12231;
	wire [4-1:0] node12235;
	wire [4-1:0] node12236;
	wire [4-1:0] node12237;
	wire [4-1:0] node12238;
	wire [4-1:0] node12239;
	wire [4-1:0] node12243;
	wire [4-1:0] node12244;
	wire [4-1:0] node12248;
	wire [4-1:0] node12249;
	wire [4-1:0] node12250;
	wire [4-1:0] node12254;
	wire [4-1:0] node12255;
	wire [4-1:0] node12259;
	wire [4-1:0] node12260;
	wire [4-1:0] node12261;
	wire [4-1:0] node12262;
	wire [4-1:0] node12264;
	wire [4-1:0] node12268;
	wire [4-1:0] node12269;
	wire [4-1:0] node12272;
	wire [4-1:0] node12275;
	wire [4-1:0] node12276;
	wire [4-1:0] node12279;
	wire [4-1:0] node12282;
	wire [4-1:0] node12283;
	wire [4-1:0] node12284;
	wire [4-1:0] node12285;
	wire [4-1:0] node12286;
	wire [4-1:0] node12287;
	wire [4-1:0] node12288;
	wire [4-1:0] node12289;
	wire [4-1:0] node12293;
	wire [4-1:0] node12294;
	wire [4-1:0] node12298;
	wire [4-1:0] node12299;
	wire [4-1:0] node12300;
	wire [4-1:0] node12303;
	wire [4-1:0] node12307;
	wire [4-1:0] node12308;
	wire [4-1:0] node12309;
	wire [4-1:0] node12311;
	wire [4-1:0] node12314;
	wire [4-1:0] node12315;
	wire [4-1:0] node12318;
	wire [4-1:0] node12321;
	wire [4-1:0] node12322;
	wire [4-1:0] node12325;
	wire [4-1:0] node12326;
	wire [4-1:0] node12329;
	wire [4-1:0] node12332;
	wire [4-1:0] node12333;
	wire [4-1:0] node12334;
	wire [4-1:0] node12335;
	wire [4-1:0] node12337;
	wire [4-1:0] node12340;
	wire [4-1:0] node12341;
	wire [4-1:0] node12344;
	wire [4-1:0] node12347;
	wire [4-1:0] node12348;
	wire [4-1:0] node12349;
	wire [4-1:0] node12352;
	wire [4-1:0] node12355;
	wire [4-1:0] node12356;
	wire [4-1:0] node12359;
	wire [4-1:0] node12362;
	wire [4-1:0] node12363;
	wire [4-1:0] node12364;
	wire [4-1:0] node12365;
	wire [4-1:0] node12368;
	wire [4-1:0] node12371;
	wire [4-1:0] node12372;
	wire [4-1:0] node12376;
	wire [4-1:0] node12377;
	wire [4-1:0] node12381;
	wire [4-1:0] node12382;
	wire [4-1:0] node12383;
	wire [4-1:0] node12384;
	wire [4-1:0] node12385;
	wire [4-1:0] node12386;
	wire [4-1:0] node12390;
	wire [4-1:0] node12391;
	wire [4-1:0] node12394;
	wire [4-1:0] node12397;
	wire [4-1:0] node12399;
	wire [4-1:0] node12401;
	wire [4-1:0] node12404;
	wire [4-1:0] node12405;
	wire [4-1:0] node12406;
	wire [4-1:0] node12407;
	wire [4-1:0] node12411;
	wire [4-1:0] node12412;
	wire [4-1:0] node12415;
	wire [4-1:0] node12418;
	wire [4-1:0] node12419;
	wire [4-1:0] node12420;
	wire [4-1:0] node12424;
	wire [4-1:0] node12426;
	wire [4-1:0] node12429;
	wire [4-1:0] node12430;
	wire [4-1:0] node12431;
	wire [4-1:0] node12432;
	wire [4-1:0] node12433;
	wire [4-1:0] node12436;
	wire [4-1:0] node12439;
	wire [4-1:0] node12440;
	wire [4-1:0] node12443;
	wire [4-1:0] node12446;
	wire [4-1:0] node12447;
	wire [4-1:0] node12450;
	wire [4-1:0] node12453;
	wire [4-1:0] node12454;
	wire [4-1:0] node12455;
	wire [4-1:0] node12456;
	wire [4-1:0] node12459;
	wire [4-1:0] node12462;
	wire [4-1:0] node12463;
	wire [4-1:0] node12466;
	wire [4-1:0] node12469;
	wire [4-1:0] node12470;
	wire [4-1:0] node12471;
	wire [4-1:0] node12474;
	wire [4-1:0] node12477;
	wire [4-1:0] node12478;
	wire [4-1:0] node12481;
	wire [4-1:0] node12484;
	wire [4-1:0] node12485;
	wire [4-1:0] node12486;
	wire [4-1:0] node12487;
	wire [4-1:0] node12488;
	wire [4-1:0] node12489;
	wire [4-1:0] node12493;
	wire [4-1:0] node12494;
	wire [4-1:0] node12497;
	wire [4-1:0] node12500;
	wire [4-1:0] node12501;
	wire [4-1:0] node12502;
	wire [4-1:0] node12506;
	wire [4-1:0] node12508;
	wire [4-1:0] node12511;
	wire [4-1:0] node12512;
	wire [4-1:0] node12513;
	wire [4-1:0] node12514;
	wire [4-1:0] node12518;
	wire [4-1:0] node12519;
	wire [4-1:0] node12522;
	wire [4-1:0] node12525;
	wire [4-1:0] node12526;
	wire [4-1:0] node12527;
	wire [4-1:0] node12530;
	wire [4-1:0] node12533;
	wire [4-1:0] node12535;
	wire [4-1:0] node12538;
	wire [4-1:0] node12539;
	wire [4-1:0] node12540;
	wire [4-1:0] node12541;
	wire [4-1:0] node12543;
	wire [4-1:0] node12546;
	wire [4-1:0] node12549;
	wire [4-1:0] node12550;
	wire [4-1:0] node12553;
	wire [4-1:0] node12556;
	wire [4-1:0] node12557;
	wire [4-1:0] node12558;
	wire [4-1:0] node12560;
	wire [4-1:0] node12563;
	wire [4-1:0] node12566;
	wire [4-1:0] node12567;
	wire [4-1:0] node12569;
	wire [4-1:0] node12572;
	wire [4-1:0] node12575;
	wire [4-1:0] node12576;
	wire [4-1:0] node12577;
	wire [4-1:0] node12578;
	wire [4-1:0] node12579;
	wire [4-1:0] node12580;
	wire [4-1:0] node12581;
	wire [4-1:0] node12582;
	wire [4-1:0] node12583;
	wire [4-1:0] node12586;
	wire [4-1:0] node12589;
	wire [4-1:0] node12590;
	wire [4-1:0] node12593;
	wire [4-1:0] node12597;
	wire [4-1:0] node12598;
	wire [4-1:0] node12599;
	wire [4-1:0] node12600;
	wire [4-1:0] node12603;
	wire [4-1:0] node12606;
	wire [4-1:0] node12607;
	wire [4-1:0] node12610;
	wire [4-1:0] node12614;
	wire [4-1:0] node12615;
	wire [4-1:0] node12616;
	wire [4-1:0] node12617;
	wire [4-1:0] node12620;
	wire [4-1:0] node12624;
	wire [4-1:0] node12625;
	wire [4-1:0] node12626;
	wire [4-1:0] node12629;
	wire [4-1:0] node12633;
	wire [4-1:0] node12634;
	wire [4-1:0] node12635;
	wire [4-1:0] node12636;
	wire [4-1:0] node12638;
	wire [4-1:0] node12641;
	wire [4-1:0] node12643;
	wire [4-1:0] node12646;
	wire [4-1:0] node12647;
	wire [4-1:0] node12649;
	wire [4-1:0] node12652;
	wire [4-1:0] node12653;
	wire [4-1:0] node12657;
	wire [4-1:0] node12658;
	wire [4-1:0] node12659;
	wire [4-1:0] node12660;
	wire [4-1:0] node12661;
	wire [4-1:0] node12665;
	wire [4-1:0] node12666;
	wire [4-1:0] node12669;
	wire [4-1:0] node12672;
	wire [4-1:0] node12673;
	wire [4-1:0] node12674;
	wire [4-1:0] node12677;
	wire [4-1:0] node12680;
	wire [4-1:0] node12681;
	wire [4-1:0] node12684;
	wire [4-1:0] node12687;
	wire [4-1:0] node12688;
	wire [4-1:0] node12690;
	wire [4-1:0] node12691;
	wire [4-1:0] node12694;
	wire [4-1:0] node12697;
	wire [4-1:0] node12698;
	wire [4-1:0] node12700;
	wire [4-1:0] node12703;
	wire [4-1:0] node12705;
	wire [4-1:0] node12708;
	wire [4-1:0] node12709;
	wire [4-1:0] node12710;
	wire [4-1:0] node12711;
	wire [4-1:0] node12712;
	wire [4-1:0] node12713;
	wire [4-1:0] node12714;
	wire [4-1:0] node12717;
	wire [4-1:0] node12720;
	wire [4-1:0] node12721;
	wire [4-1:0] node12724;
	wire [4-1:0] node12727;
	wire [4-1:0] node12728;
	wire [4-1:0] node12730;
	wire [4-1:0] node12733;
	wire [4-1:0] node12734;
	wire [4-1:0] node12738;
	wire [4-1:0] node12739;
	wire [4-1:0] node12742;
	wire [4-1:0] node12745;
	wire [4-1:0] node12746;
	wire [4-1:0] node12747;
	wire [4-1:0] node12750;
	wire [4-1:0] node12753;
	wire [4-1:0] node12754;
	wire [4-1:0] node12755;
	wire [4-1:0] node12756;
	wire [4-1:0] node12759;
	wire [4-1:0] node12762;
	wire [4-1:0] node12763;
	wire [4-1:0] node12766;
	wire [4-1:0] node12769;
	wire [4-1:0] node12770;
	wire [4-1:0] node12771;
	wire [4-1:0] node12774;
	wire [4-1:0] node12777;
	wire [4-1:0] node12778;
	wire [4-1:0] node12782;
	wire [4-1:0] node12783;
	wire [4-1:0] node12784;
	wire [4-1:0] node12785;
	wire [4-1:0] node12786;
	wire [4-1:0] node12787;
	wire [4-1:0] node12790;
	wire [4-1:0] node12794;
	wire [4-1:0] node12795;
	wire [4-1:0] node12797;
	wire [4-1:0] node12800;
	wire [4-1:0] node12803;
	wire [4-1:0] node12804;
	wire [4-1:0] node12805;
	wire [4-1:0] node12808;
	wire [4-1:0] node12811;
	wire [4-1:0] node12813;
	wire [4-1:0] node12815;
	wire [4-1:0] node12818;
	wire [4-1:0] node12819;
	wire [4-1:0] node12820;
	wire [4-1:0] node12821;
	wire [4-1:0] node12825;
	wire [4-1:0] node12826;
	wire [4-1:0] node12830;
	wire [4-1:0] node12831;
	wire [4-1:0] node12834;
	wire [4-1:0] node12835;
	wire [4-1:0] node12839;
	wire [4-1:0] node12840;
	wire [4-1:0] node12841;
	wire [4-1:0] node12842;
	wire [4-1:0] node12843;
	wire [4-1:0] node12844;
	wire [4-1:0] node12845;
	wire [4-1:0] node12848;
	wire [4-1:0] node12851;
	wire [4-1:0] node12852;
	wire [4-1:0] node12853;
	wire [4-1:0] node12856;
	wire [4-1:0] node12859;
	wire [4-1:0] node12860;
	wire [4-1:0] node12863;
	wire [4-1:0] node12866;
	wire [4-1:0] node12867;
	wire [4-1:0] node12869;
	wire [4-1:0] node12870;
	wire [4-1:0] node12873;
	wire [4-1:0] node12876;
	wire [4-1:0] node12877;
	wire [4-1:0] node12879;
	wire [4-1:0] node12882;
	wire [4-1:0] node12884;
	wire [4-1:0] node12887;
	wire [4-1:0] node12888;
	wire [4-1:0] node12891;
	wire [4-1:0] node12894;
	wire [4-1:0] node12895;
	wire [4-1:0] node12896;
	wire [4-1:0] node12897;
	wire [4-1:0] node12898;
	wire [4-1:0] node12899;
	wire [4-1:0] node12902;
	wire [4-1:0] node12905;
	wire [4-1:0] node12906;
	wire [4-1:0] node12909;
	wire [4-1:0] node12912;
	wire [4-1:0] node12913;
	wire [4-1:0] node12914;
	wire [4-1:0] node12917;
	wire [4-1:0] node12920;
	wire [4-1:0] node12921;
	wire [4-1:0] node12924;
	wire [4-1:0] node12927;
	wire [4-1:0] node12928;
	wire [4-1:0] node12929;
	wire [4-1:0] node12932;
	wire [4-1:0] node12935;
	wire [4-1:0] node12936;
	wire [4-1:0] node12939;
	wire [4-1:0] node12942;
	wire [4-1:0] node12943;
	wire [4-1:0] node12944;
	wire [4-1:0] node12945;
	wire [4-1:0] node12948;
	wire [4-1:0] node12951;
	wire [4-1:0] node12952;
	wire [4-1:0] node12955;
	wire [4-1:0] node12958;
	wire [4-1:0] node12959;
	wire [4-1:0] node12960;
	wire [4-1:0] node12961;
	wire [4-1:0] node12965;
	wire [4-1:0] node12966;
	wire [4-1:0] node12969;
	wire [4-1:0] node12972;
	wire [4-1:0] node12973;
	wire [4-1:0] node12974;
	wire [4-1:0] node12977;
	wire [4-1:0] node12981;
	wire [4-1:0] node12982;
	wire [4-1:0] node12983;
	wire [4-1:0] node12984;
	wire [4-1:0] node12985;
	wire [4-1:0] node12986;
	wire [4-1:0] node12987;
	wire [4-1:0] node12990;
	wire [4-1:0] node12993;
	wire [4-1:0] node12994;
	wire [4-1:0] node12997;
	wire [4-1:0] node13000;
	wire [4-1:0] node13001;
	wire [4-1:0] node13002;
	wire [4-1:0] node13005;
	wire [4-1:0] node13008;
	wire [4-1:0] node13009;
	wire [4-1:0] node13012;
	wire [4-1:0] node13015;
	wire [4-1:0] node13016;
	wire [4-1:0] node13017;
	wire [4-1:0] node13018;
	wire [4-1:0] node13021;
	wire [4-1:0] node13024;
	wire [4-1:0] node13025;
	wire [4-1:0] node13028;
	wire [4-1:0] node13031;
	wire [4-1:0] node13032;
	wire [4-1:0] node13033;
	wire [4-1:0] node13036;
	wire [4-1:0] node13039;
	wire [4-1:0] node13040;
	wire [4-1:0] node13044;
	wire [4-1:0] node13045;
	wire [4-1:0] node13048;
	wire [4-1:0] node13051;
	wire [4-1:0] node13052;
	wire [4-1:0] node13053;
	wire [4-1:0] node13054;
	wire [4-1:0] node13055;
	wire [4-1:0] node13058;
	wire [4-1:0] node13061;
	wire [4-1:0] node13062;
	wire [4-1:0] node13063;
	wire [4-1:0] node13066;
	wire [4-1:0] node13069;
	wire [4-1:0] node13070;
	wire [4-1:0] node13073;
	wire [4-1:0] node13076;
	wire [4-1:0] node13077;
	wire [4-1:0] node13078;
	wire [4-1:0] node13079;
	wire [4-1:0] node13083;
	wire [4-1:0] node13085;
	wire [4-1:0] node13088;
	wire [4-1:0] node13089;
	wire [4-1:0] node13090;
	wire [4-1:0] node13093;
	wire [4-1:0] node13096;
	wire [4-1:0] node13097;
	wire [4-1:0] node13100;
	wire [4-1:0] node13103;
	wire [4-1:0] node13104;
	wire [4-1:0] node13105;
	wire [4-1:0] node13108;
	wire [4-1:0] node13111;
	wire [4-1:0] node13112;
	wire [4-1:0] node13113;
	wire [4-1:0] node13114;
	wire [4-1:0] node13117;
	wire [4-1:0] node13121;
	wire [4-1:0] node13122;
	wire [4-1:0] node13124;
	wire [4-1:0] node13127;
	wire [4-1:0] node13128;
	wire [4-1:0] node13131;
	wire [4-1:0] node13134;
	wire [4-1:0] node13135;
	wire [4-1:0] node13136;
	wire [4-1:0] node13137;
	wire [4-1:0] node13138;
	wire [4-1:0] node13139;
	wire [4-1:0] node13140;
	wire [4-1:0] node13141;
	wire [4-1:0] node13142;
	wire [4-1:0] node13143;
	wire [4-1:0] node13144;
	wire [4-1:0] node13145;
	wire [4-1:0] node13149;
	wire [4-1:0] node13150;
	wire [4-1:0] node13154;
	wire [4-1:0] node13155;
	wire [4-1:0] node13156;
	wire [4-1:0] node13159;
	wire [4-1:0] node13162;
	wire [4-1:0] node13163;
	wire [4-1:0] node13166;
	wire [4-1:0] node13169;
	wire [4-1:0] node13170;
	wire [4-1:0] node13171;
	wire [4-1:0] node13173;
	wire [4-1:0] node13176;
	wire [4-1:0] node13177;
	wire [4-1:0] node13180;
	wire [4-1:0] node13183;
	wire [4-1:0] node13184;
	wire [4-1:0] node13185;
	wire [4-1:0] node13189;
	wire [4-1:0] node13192;
	wire [4-1:0] node13193;
	wire [4-1:0] node13194;
	wire [4-1:0] node13195;
	wire [4-1:0] node13196;
	wire [4-1:0] node13201;
	wire [4-1:0] node13202;
	wire [4-1:0] node13203;
	wire [4-1:0] node13207;
	wire [4-1:0] node13210;
	wire [4-1:0] node13211;
	wire [4-1:0] node13212;
	wire [4-1:0] node13214;
	wire [4-1:0] node13217;
	wire [4-1:0] node13220;
	wire [4-1:0] node13221;
	wire [4-1:0] node13224;
	wire [4-1:0] node13227;
	wire [4-1:0] node13228;
	wire [4-1:0] node13229;
	wire [4-1:0] node13230;
	wire [4-1:0] node13231;
	wire [4-1:0] node13232;
	wire [4-1:0] node13235;
	wire [4-1:0] node13238;
	wire [4-1:0] node13239;
	wire [4-1:0] node13242;
	wire [4-1:0] node13245;
	wire [4-1:0] node13246;
	wire [4-1:0] node13249;
	wire [4-1:0] node13252;
	wire [4-1:0] node13253;
	wire [4-1:0] node13254;
	wire [4-1:0] node13255;
	wire [4-1:0] node13258;
	wire [4-1:0] node13261;
	wire [4-1:0] node13262;
	wire [4-1:0] node13265;
	wire [4-1:0] node13268;
	wire [4-1:0] node13269;
	wire [4-1:0] node13272;
	wire [4-1:0] node13275;
	wire [4-1:0] node13276;
	wire [4-1:0] node13277;
	wire [4-1:0] node13278;
	wire [4-1:0] node13279;
	wire [4-1:0] node13282;
	wire [4-1:0] node13285;
	wire [4-1:0] node13286;
	wire [4-1:0] node13289;
	wire [4-1:0] node13292;
	wire [4-1:0] node13293;
	wire [4-1:0] node13294;
	wire [4-1:0] node13297;
	wire [4-1:0] node13300;
	wire [4-1:0] node13301;
	wire [4-1:0] node13304;
	wire [4-1:0] node13307;
	wire [4-1:0] node13308;
	wire [4-1:0] node13309;
	wire [4-1:0] node13310;
	wire [4-1:0] node13313;
	wire [4-1:0] node13316;
	wire [4-1:0] node13317;
	wire [4-1:0] node13320;
	wire [4-1:0] node13323;
	wire [4-1:0] node13324;
	wire [4-1:0] node13325;
	wire [4-1:0] node13328;
	wire [4-1:0] node13331;
	wire [4-1:0] node13333;
	wire [4-1:0] node13336;
	wire [4-1:0] node13337;
	wire [4-1:0] node13338;
	wire [4-1:0] node13339;
	wire [4-1:0] node13340;
	wire [4-1:0] node13341;
	wire [4-1:0] node13342;
	wire [4-1:0] node13345;
	wire [4-1:0] node13349;
	wire [4-1:0] node13350;
	wire [4-1:0] node13353;
	wire [4-1:0] node13356;
	wire [4-1:0] node13357;
	wire [4-1:0] node13358;
	wire [4-1:0] node13362;
	wire [4-1:0] node13363;
	wire [4-1:0] node13366;
	wire [4-1:0] node13369;
	wire [4-1:0] node13370;
	wire [4-1:0] node13371;
	wire [4-1:0] node13372;
	wire [4-1:0] node13373;
	wire [4-1:0] node13376;
	wire [4-1:0] node13379;
	wire [4-1:0] node13380;
	wire [4-1:0] node13383;
	wire [4-1:0] node13386;
	wire [4-1:0] node13387;
	wire [4-1:0] node13390;
	wire [4-1:0] node13393;
	wire [4-1:0] node13394;
	wire [4-1:0] node13395;
	wire [4-1:0] node13398;
	wire [4-1:0] node13400;
	wire [4-1:0] node13403;
	wire [4-1:0] node13404;
	wire [4-1:0] node13407;
	wire [4-1:0] node13408;
	wire [4-1:0] node13412;
	wire [4-1:0] node13413;
	wire [4-1:0] node13414;
	wire [4-1:0] node13415;
	wire [4-1:0] node13416;
	wire [4-1:0] node13417;
	wire [4-1:0] node13421;
	wire [4-1:0] node13422;
	wire [4-1:0] node13426;
	wire [4-1:0] node13427;
	wire [4-1:0] node13430;
	wire [4-1:0] node13432;
	wire [4-1:0] node13435;
	wire [4-1:0] node13436;
	wire [4-1:0] node13437;
	wire [4-1:0] node13438;
	wire [4-1:0] node13441;
	wire [4-1:0] node13444;
	wire [4-1:0] node13445;
	wire [4-1:0] node13448;
	wire [4-1:0] node13451;
	wire [4-1:0] node13452;
	wire [4-1:0] node13455;
	wire [4-1:0] node13457;
	wire [4-1:0] node13460;
	wire [4-1:0] node13461;
	wire [4-1:0] node13462;
	wire [4-1:0] node13464;
	wire [4-1:0] node13467;
	wire [4-1:0] node13468;
	wire [4-1:0] node13469;
	wire [4-1:0] node13472;
	wire [4-1:0] node13475;
	wire [4-1:0] node13476;
	wire [4-1:0] node13479;
	wire [4-1:0] node13482;
	wire [4-1:0] node13483;
	wire [4-1:0] node13484;
	wire [4-1:0] node13485;
	wire [4-1:0] node13488;
	wire [4-1:0] node13492;
	wire [4-1:0] node13493;
	wire [4-1:0] node13496;
	wire [4-1:0] node13498;
	wire [4-1:0] node13501;
	wire [4-1:0] node13502;
	wire [4-1:0] node13503;
	wire [4-1:0] node13504;
	wire [4-1:0] node13505;
	wire [4-1:0] node13506;
	wire [4-1:0] node13507;
	wire [4-1:0] node13508;
	wire [4-1:0] node13512;
	wire [4-1:0] node13515;
	wire [4-1:0] node13516;
	wire [4-1:0] node13519;
	wire [4-1:0] node13520;
	wire [4-1:0] node13524;
	wire [4-1:0] node13525;
	wire [4-1:0] node13526;
	wire [4-1:0] node13527;
	wire [4-1:0] node13531;
	wire [4-1:0] node13534;
	wire [4-1:0] node13535;
	wire [4-1:0] node13538;
	wire [4-1:0] node13541;
	wire [4-1:0] node13542;
	wire [4-1:0] node13543;
	wire [4-1:0] node13544;
	wire [4-1:0] node13545;
	wire [4-1:0] node13549;
	wire [4-1:0] node13552;
	wire [4-1:0] node13553;
	wire [4-1:0] node13554;
	wire [4-1:0] node13557;
	wire [4-1:0] node13560;
	wire [4-1:0] node13561;
	wire [4-1:0] node13564;
	wire [4-1:0] node13567;
	wire [4-1:0] node13568;
	wire [4-1:0] node13569;
	wire [4-1:0] node13570;
	wire [4-1:0] node13574;
	wire [4-1:0] node13577;
	wire [4-1:0] node13578;
	wire [4-1:0] node13581;
	wire [4-1:0] node13582;
	wire [4-1:0] node13586;
	wire [4-1:0] node13587;
	wire [4-1:0] node13588;
	wire [4-1:0] node13589;
	wire [4-1:0] node13590;
	wire [4-1:0] node13593;
	wire [4-1:0] node13596;
	wire [4-1:0] node13597;
	wire [4-1:0] node13600;
	wire [4-1:0] node13603;
	wire [4-1:0] node13604;
	wire [4-1:0] node13605;
	wire [4-1:0] node13608;
	wire [4-1:0] node13611;
	wire [4-1:0] node13612;
	wire [4-1:0] node13613;
	wire [4-1:0] node13616;
	wire [4-1:0] node13619;
	wire [4-1:0] node13620;
	wire [4-1:0] node13623;
	wire [4-1:0] node13626;
	wire [4-1:0] node13627;
	wire [4-1:0] node13628;
	wire [4-1:0] node13629;
	wire [4-1:0] node13632;
	wire [4-1:0] node13635;
	wire [4-1:0] node13636;
	wire [4-1:0] node13637;
	wire [4-1:0] node13640;
	wire [4-1:0] node13643;
	wire [4-1:0] node13644;
	wire [4-1:0] node13648;
	wire [4-1:0] node13649;
	wire [4-1:0] node13650;
	wire [4-1:0] node13651;
	wire [4-1:0] node13654;
	wire [4-1:0] node13657;
	wire [4-1:0] node13658;
	wire [4-1:0] node13661;
	wire [4-1:0] node13664;
	wire [4-1:0] node13665;
	wire [4-1:0] node13666;
	wire [4-1:0] node13669;
	wire [4-1:0] node13672;
	wire [4-1:0] node13673;
	wire [4-1:0] node13676;
	wire [4-1:0] node13679;
	wire [4-1:0] node13680;
	wire [4-1:0] node13681;
	wire [4-1:0] node13682;
	wire [4-1:0] node13683;
	wire [4-1:0] node13684;
	wire [4-1:0] node13685;
	wire [4-1:0] node13688;
	wire [4-1:0] node13691;
	wire [4-1:0] node13692;
	wire [4-1:0] node13696;
	wire [4-1:0] node13697;
	wire [4-1:0] node13699;
	wire [4-1:0] node13702;
	wire [4-1:0] node13703;
	wire [4-1:0] node13707;
	wire [4-1:0] node13708;
	wire [4-1:0] node13709;
	wire [4-1:0] node13710;
	wire [4-1:0] node13713;
	wire [4-1:0] node13716;
	wire [4-1:0] node13717;
	wire [4-1:0] node13721;
	wire [4-1:0] node13722;
	wire [4-1:0] node13723;
	wire [4-1:0] node13726;
	wire [4-1:0] node13729;
	wire [4-1:0] node13732;
	wire [4-1:0] node13733;
	wire [4-1:0] node13734;
	wire [4-1:0] node13735;
	wire [4-1:0] node13736;
	wire [4-1:0] node13739;
	wire [4-1:0] node13742;
	wire [4-1:0] node13744;
	wire [4-1:0] node13747;
	wire [4-1:0] node13748;
	wire [4-1:0] node13749;
	wire [4-1:0] node13753;
	wire [4-1:0] node13754;
	wire [4-1:0] node13757;
	wire [4-1:0] node13760;
	wire [4-1:0] node13761;
	wire [4-1:0] node13762;
	wire [4-1:0] node13763;
	wire [4-1:0] node13766;
	wire [4-1:0] node13769;
	wire [4-1:0] node13770;
	wire [4-1:0] node13773;
	wire [4-1:0] node13776;
	wire [4-1:0] node13777;
	wire [4-1:0] node13779;
	wire [4-1:0] node13782;
	wire [4-1:0] node13783;
	wire [4-1:0] node13786;
	wire [4-1:0] node13789;
	wire [4-1:0] node13790;
	wire [4-1:0] node13791;
	wire [4-1:0] node13792;
	wire [4-1:0] node13793;
	wire [4-1:0] node13794;
	wire [4-1:0] node13798;
	wire [4-1:0] node13801;
	wire [4-1:0] node13802;
	wire [4-1:0] node13803;
	wire [4-1:0] node13807;
	wire [4-1:0] node13810;
	wire [4-1:0] node13811;
	wire [4-1:0] node13812;
	wire [4-1:0] node13813;
	wire [4-1:0] node13816;
	wire [4-1:0] node13819;
	wire [4-1:0] node13820;
	wire [4-1:0] node13823;
	wire [4-1:0] node13826;
	wire [4-1:0] node13827;
	wire [4-1:0] node13828;
	wire [4-1:0] node13832;
	wire [4-1:0] node13835;
	wire [4-1:0] node13836;
	wire [4-1:0] node13837;
	wire [4-1:0] node13838;
	wire [4-1:0] node13839;
	wire [4-1:0] node13842;
	wire [4-1:0] node13845;
	wire [4-1:0] node13846;
	wire [4-1:0] node13849;
	wire [4-1:0] node13852;
	wire [4-1:0] node13853;
	wire [4-1:0] node13854;
	wire [4-1:0] node13858;
	wire [4-1:0] node13859;
	wire [4-1:0] node13862;
	wire [4-1:0] node13865;
	wire [4-1:0] node13866;
	wire [4-1:0] node13867;
	wire [4-1:0] node13868;
	wire [4-1:0] node13872;
	wire [4-1:0] node13873;
	wire [4-1:0] node13876;
	wire [4-1:0] node13879;
	wire [4-1:0] node13880;
	wire [4-1:0] node13881;
	wire [4-1:0] node13884;
	wire [4-1:0] node13887;
	wire [4-1:0] node13890;
	wire [4-1:0] node13891;
	wire [4-1:0] node13892;
	wire [4-1:0] node13893;
	wire [4-1:0] node13894;
	wire [4-1:0] node13895;
	wire [4-1:0] node13896;
	wire [4-1:0] node13897;
	wire [4-1:0] node13898;
	wire [4-1:0] node13901;
	wire [4-1:0] node13904;
	wire [4-1:0] node13905;
	wire [4-1:0] node13908;
	wire [4-1:0] node13911;
	wire [4-1:0] node13912;
	wire [4-1:0] node13913;
	wire [4-1:0] node13916;
	wire [4-1:0] node13919;
	wire [4-1:0] node13920;
	wire [4-1:0] node13924;
	wire [4-1:0] node13925;
	wire [4-1:0] node13926;
	wire [4-1:0] node13927;
	wire [4-1:0] node13930;
	wire [4-1:0] node13933;
	wire [4-1:0] node13934;
	wire [4-1:0] node13937;
	wire [4-1:0] node13940;
	wire [4-1:0] node13941;
	wire [4-1:0] node13943;
	wire [4-1:0] node13946;
	wire [4-1:0] node13947;
	wire [4-1:0] node13951;
	wire [4-1:0] node13952;
	wire [4-1:0] node13953;
	wire [4-1:0] node13955;
	wire [4-1:0] node13957;
	wire [4-1:0] node13960;
	wire [4-1:0] node13961;
	wire [4-1:0] node13964;
	wire [4-1:0] node13967;
	wire [4-1:0] node13968;
	wire [4-1:0] node13969;
	wire [4-1:0] node13970;
	wire [4-1:0] node13973;
	wire [4-1:0] node13976;
	wire [4-1:0] node13977;
	wire [4-1:0] node13980;
	wire [4-1:0] node13983;
	wire [4-1:0] node13984;
	wire [4-1:0] node13985;
	wire [4-1:0] node13989;
	wire [4-1:0] node13990;
	wire [4-1:0] node13993;
	wire [4-1:0] node13996;
	wire [4-1:0] node13997;
	wire [4-1:0] node13998;
	wire [4-1:0] node13999;
	wire [4-1:0] node14000;
	wire [4-1:0] node14001;
	wire [4-1:0] node14004;
	wire [4-1:0] node14007;
	wire [4-1:0] node14008;
	wire [4-1:0] node14012;
	wire [4-1:0] node14013;
	wire [4-1:0] node14016;
	wire [4-1:0] node14018;
	wire [4-1:0] node14021;
	wire [4-1:0] node14022;
	wire [4-1:0] node14023;
	wire [4-1:0] node14024;
	wire [4-1:0] node14027;
	wire [4-1:0] node14030;
	wire [4-1:0] node14031;
	wire [4-1:0] node14034;
	wire [4-1:0] node14037;
	wire [4-1:0] node14038;
	wire [4-1:0] node14039;
	wire [4-1:0] node14043;
	wire [4-1:0] node14044;
	wire [4-1:0] node14047;
	wire [4-1:0] node14050;
	wire [4-1:0] node14051;
	wire [4-1:0] node14052;
	wire [4-1:0] node14053;
	wire [4-1:0] node14054;
	wire [4-1:0] node14058;
	wire [4-1:0] node14059;
	wire [4-1:0] node14062;
	wire [4-1:0] node14065;
	wire [4-1:0] node14067;
	wire [4-1:0] node14068;
	wire [4-1:0] node14071;
	wire [4-1:0] node14074;
	wire [4-1:0] node14075;
	wire [4-1:0] node14076;
	wire [4-1:0] node14079;
	wire [4-1:0] node14080;
	wire [4-1:0] node14083;
	wire [4-1:0] node14086;
	wire [4-1:0] node14087;
	wire [4-1:0] node14088;
	wire [4-1:0] node14091;
	wire [4-1:0] node14095;
	wire [4-1:0] node14096;
	wire [4-1:0] node14097;
	wire [4-1:0] node14098;
	wire [4-1:0] node14099;
	wire [4-1:0] node14100;
	wire [4-1:0] node14101;
	wire [4-1:0] node14104;
	wire [4-1:0] node14107;
	wire [4-1:0] node14108;
	wire [4-1:0] node14111;
	wire [4-1:0] node14114;
	wire [4-1:0] node14115;
	wire [4-1:0] node14116;
	wire [4-1:0] node14119;
	wire [4-1:0] node14122;
	wire [4-1:0] node14123;
	wire [4-1:0] node14126;
	wire [4-1:0] node14129;
	wire [4-1:0] node14130;
	wire [4-1:0] node14131;
	wire [4-1:0] node14133;
	wire [4-1:0] node14136;
	wire [4-1:0] node14137;
	wire [4-1:0] node14140;
	wire [4-1:0] node14143;
	wire [4-1:0] node14144;
	wire [4-1:0] node14145;
	wire [4-1:0] node14148;
	wire [4-1:0] node14151;
	wire [4-1:0] node14152;
	wire [4-1:0] node14155;
	wire [4-1:0] node14158;
	wire [4-1:0] node14159;
	wire [4-1:0] node14160;
	wire [4-1:0] node14161;
	wire [4-1:0] node14162;
	wire [4-1:0] node14165;
	wire [4-1:0] node14168;
	wire [4-1:0] node14169;
	wire [4-1:0] node14172;
	wire [4-1:0] node14175;
	wire [4-1:0] node14176;
	wire [4-1:0] node14177;
	wire [4-1:0] node14180;
	wire [4-1:0] node14184;
	wire [4-1:0] node14185;
	wire [4-1:0] node14186;
	wire [4-1:0] node14187;
	wire [4-1:0] node14190;
	wire [4-1:0] node14193;
	wire [4-1:0] node14194;
	wire [4-1:0] node14198;
	wire [4-1:0] node14199;
	wire [4-1:0] node14200;
	wire [4-1:0] node14203;
	wire [4-1:0] node14206;
	wire [4-1:0] node14207;
	wire [4-1:0] node14211;
	wire [4-1:0] node14212;
	wire [4-1:0] node14213;
	wire [4-1:0] node14214;
	wire [4-1:0] node14216;
	wire [4-1:0] node14217;
	wire [4-1:0] node14220;
	wire [4-1:0] node14223;
	wire [4-1:0] node14224;
	wire [4-1:0] node14226;
	wire [4-1:0] node14229;
	wire [4-1:0] node14230;
	wire [4-1:0] node14233;
	wire [4-1:0] node14236;
	wire [4-1:0] node14237;
	wire [4-1:0] node14238;
	wire [4-1:0] node14239;
	wire [4-1:0] node14242;
	wire [4-1:0] node14245;
	wire [4-1:0] node14246;
	wire [4-1:0] node14249;
	wire [4-1:0] node14252;
	wire [4-1:0] node14253;
	wire [4-1:0] node14254;
	wire [4-1:0] node14257;
	wire [4-1:0] node14260;
	wire [4-1:0] node14261;
	wire [4-1:0] node14265;
	wire [4-1:0] node14266;
	wire [4-1:0] node14267;
	wire [4-1:0] node14268;
	wire [4-1:0] node14269;
	wire [4-1:0] node14272;
	wire [4-1:0] node14275;
	wire [4-1:0] node14276;
	wire [4-1:0] node14279;
	wire [4-1:0] node14282;
	wire [4-1:0] node14283;
	wire [4-1:0] node14284;
	wire [4-1:0] node14287;
	wire [4-1:0] node14290;
	wire [4-1:0] node14291;
	wire [4-1:0] node14294;
	wire [4-1:0] node14297;
	wire [4-1:0] node14298;
	wire [4-1:0] node14299;
	wire [4-1:0] node14300;
	wire [4-1:0] node14303;
	wire [4-1:0] node14306;
	wire [4-1:0] node14307;
	wire [4-1:0] node14310;
	wire [4-1:0] node14313;
	wire [4-1:0] node14314;
	wire [4-1:0] node14315;
	wire [4-1:0] node14318;
	wire [4-1:0] node14321;
	wire [4-1:0] node14322;
	wire [4-1:0] node14325;
	wire [4-1:0] node14328;
	wire [4-1:0] node14329;
	wire [4-1:0] node14330;
	wire [4-1:0] node14331;
	wire [4-1:0] node14332;
	wire [4-1:0] node14333;
	wire [4-1:0] node14334;
	wire [4-1:0] node14337;
	wire [4-1:0] node14338;
	wire [4-1:0] node14341;
	wire [4-1:0] node14344;
	wire [4-1:0] node14345;
	wire [4-1:0] node14348;
	wire [4-1:0] node14351;
	wire [4-1:0] node14352;
	wire [4-1:0] node14354;
	wire [4-1:0] node14355;
	wire [4-1:0] node14359;
	wire [4-1:0] node14360;
	wire [4-1:0] node14363;
	wire [4-1:0] node14364;
	wire [4-1:0] node14368;
	wire [4-1:0] node14369;
	wire [4-1:0] node14370;
	wire [4-1:0] node14371;
	wire [4-1:0] node14373;
	wire [4-1:0] node14376;
	wire [4-1:0] node14377;
	wire [4-1:0] node14380;
	wire [4-1:0] node14383;
	wire [4-1:0] node14384;
	wire [4-1:0] node14385;
	wire [4-1:0] node14388;
	wire [4-1:0] node14391;
	wire [4-1:0] node14392;
	wire [4-1:0] node14395;
	wire [4-1:0] node14398;
	wire [4-1:0] node14399;
	wire [4-1:0] node14401;
	wire [4-1:0] node14402;
	wire [4-1:0] node14405;
	wire [4-1:0] node14408;
	wire [4-1:0] node14409;
	wire [4-1:0] node14412;
	wire [4-1:0] node14414;
	wire [4-1:0] node14417;
	wire [4-1:0] node14418;
	wire [4-1:0] node14419;
	wire [4-1:0] node14420;
	wire [4-1:0] node14421;
	wire [4-1:0] node14422;
	wire [4-1:0] node14425;
	wire [4-1:0] node14429;
	wire [4-1:0] node14431;
	wire [4-1:0] node14432;
	wire [4-1:0] node14435;
	wire [4-1:0] node14438;
	wire [4-1:0] node14439;
	wire [4-1:0] node14442;
	wire [4-1:0] node14443;
	wire [4-1:0] node14446;
	wire [4-1:0] node14449;
	wire [4-1:0] node14450;
	wire [4-1:0] node14451;
	wire [4-1:0] node14453;
	wire [4-1:0] node14454;
	wire [4-1:0] node14457;
	wire [4-1:0] node14460;
	wire [4-1:0] node14461;
	wire [4-1:0] node14462;
	wire [4-1:0] node14465;
	wire [4-1:0] node14468;
	wire [4-1:0] node14469;
	wire [4-1:0] node14472;
	wire [4-1:0] node14475;
	wire [4-1:0] node14476;
	wire [4-1:0] node14477;
	wire [4-1:0] node14478;
	wire [4-1:0] node14481;
	wire [4-1:0] node14484;
	wire [4-1:0] node14485;
	wire [4-1:0] node14488;
	wire [4-1:0] node14491;
	wire [4-1:0] node14492;
	wire [4-1:0] node14493;
	wire [4-1:0] node14496;
	wire [4-1:0] node14499;
	wire [4-1:0] node14501;
	wire [4-1:0] node14504;
	wire [4-1:0] node14505;
	wire [4-1:0] node14506;
	wire [4-1:0] node14507;
	wire [4-1:0] node14508;
	wire [4-1:0] node14509;
	wire [4-1:0] node14510;
	wire [4-1:0] node14513;
	wire [4-1:0] node14516;
	wire [4-1:0] node14517;
	wire [4-1:0] node14520;
	wire [4-1:0] node14523;
	wire [4-1:0] node14524;
	wire [4-1:0] node14527;
	wire [4-1:0] node14530;
	wire [4-1:0] node14531;
	wire [4-1:0] node14532;
	wire [4-1:0] node14533;
	wire [4-1:0] node14536;
	wire [4-1:0] node14539;
	wire [4-1:0] node14540;
	wire [4-1:0] node14543;
	wire [4-1:0] node14546;
	wire [4-1:0] node14547;
	wire [4-1:0] node14548;
	wire [4-1:0] node14551;
	wire [4-1:0] node14554;
	wire [4-1:0] node14555;
	wire [4-1:0] node14558;
	wire [4-1:0] node14561;
	wire [4-1:0] node14562;
	wire [4-1:0] node14563;
	wire [4-1:0] node14564;
	wire [4-1:0] node14565;
	wire [4-1:0] node14569;
	wire [4-1:0] node14570;
	wire [4-1:0] node14574;
	wire [4-1:0] node14575;
	wire [4-1:0] node14576;
	wire [4-1:0] node14579;
	wire [4-1:0] node14582;
	wire [4-1:0] node14583;
	wire [4-1:0] node14587;
	wire [4-1:0] node14588;
	wire [4-1:0] node14589;
	wire [4-1:0] node14590;
	wire [4-1:0] node14593;
	wire [4-1:0] node14596;
	wire [4-1:0] node14599;
	wire [4-1:0] node14600;
	wire [4-1:0] node14601;
	wire [4-1:0] node14605;
	wire [4-1:0] node14606;
	wire [4-1:0] node14610;
	wire [4-1:0] node14611;
	wire [4-1:0] node14612;
	wire [4-1:0] node14613;
	wire [4-1:0] node14614;
	wire [4-1:0] node14617;
	wire [4-1:0] node14620;
	wire [4-1:0] node14621;
	wire [4-1:0] node14624;
	wire [4-1:0] node14627;
	wire [4-1:0] node14628;
	wire [4-1:0] node14629;
	wire [4-1:0] node14630;
	wire [4-1:0] node14634;
	wire [4-1:0] node14635;
	wire [4-1:0] node14639;
	wire [4-1:0] node14640;
	wire [4-1:0] node14641;
	wire [4-1:0] node14644;
	wire [4-1:0] node14647;
	wire [4-1:0] node14648;
	wire [4-1:0] node14652;
	wire [4-1:0] node14653;
	wire [4-1:0] node14654;
	wire [4-1:0] node14655;
	wire [4-1:0] node14657;
	wire [4-1:0] node14660;
	wire [4-1:0] node14661;
	wire [4-1:0] node14664;
	wire [4-1:0] node14667;
	wire [4-1:0] node14668;
	wire [4-1:0] node14671;
	wire [4-1:0] node14672;
	wire [4-1:0] node14675;
	wire [4-1:0] node14678;
	wire [4-1:0] node14679;
	wire [4-1:0] node14681;
	wire [4-1:0] node14683;
	wire [4-1:0] node14686;
	wire [4-1:0] node14687;
	wire [4-1:0] node14688;
	wire [4-1:0] node14692;
	wire [4-1:0] node14695;
	wire [4-1:0] node14696;
	wire [4-1:0] node14697;
	wire [4-1:0] node14698;
	wire [4-1:0] node14699;
	wire [4-1:0] node14700;
	wire [4-1:0] node14701;
	wire [4-1:0] node14702;
	wire [4-1:0] node14703;
	wire [4-1:0] node14705;
	wire [4-1:0] node14708;
	wire [4-1:0] node14709;
	wire [4-1:0] node14713;
	wire [4-1:0] node14715;
	wire [4-1:0] node14717;
	wire [4-1:0] node14720;
	wire [4-1:0] node14721;
	wire [4-1:0] node14722;
	wire [4-1:0] node14723;
	wire [4-1:0] node14728;
	wire [4-1:0] node14729;
	wire [4-1:0] node14730;
	wire [4-1:0] node14734;
	wire [4-1:0] node14735;
	wire [4-1:0] node14739;
	wire [4-1:0] node14740;
	wire [4-1:0] node14741;
	wire [4-1:0] node14742;
	wire [4-1:0] node14744;
	wire [4-1:0] node14747;
	wire [4-1:0] node14749;
	wire [4-1:0] node14752;
	wire [4-1:0] node14753;
	wire [4-1:0] node14755;
	wire [4-1:0] node14758;
	wire [4-1:0] node14760;
	wire [4-1:0] node14763;
	wire [4-1:0] node14764;
	wire [4-1:0] node14766;
	wire [4-1:0] node14769;
	wire [4-1:0] node14771;
	wire [4-1:0] node14773;
	wire [4-1:0] node14776;
	wire [4-1:0] node14777;
	wire [4-1:0] node14778;
	wire [4-1:0] node14779;
	wire [4-1:0] node14780;
	wire [4-1:0] node14784;
	wire [4-1:0] node14785;
	wire [4-1:0] node14789;
	wire [4-1:0] node14790;
	wire [4-1:0] node14791;
	wire [4-1:0] node14795;
	wire [4-1:0] node14796;
	wire [4-1:0] node14800;
	wire [4-1:0] node14801;
	wire [4-1:0] node14802;
	wire [4-1:0] node14804;
	wire [4-1:0] node14805;
	wire [4-1:0] node14808;
	wire [4-1:0] node14811;
	wire [4-1:0] node14812;
	wire [4-1:0] node14815;
	wire [4-1:0] node14818;
	wire [4-1:0] node14819;
	wire [4-1:0] node14820;
	wire [4-1:0] node14821;
	wire [4-1:0] node14824;
	wire [4-1:0] node14827;
	wire [4-1:0] node14828;
	wire [4-1:0] node14831;
	wire [4-1:0] node14834;
	wire [4-1:0] node14835;
	wire [4-1:0] node14839;
	wire [4-1:0] node14840;
	wire [4-1:0] node14841;
	wire [4-1:0] node14842;
	wire [4-1:0] node14843;
	wire [4-1:0] node14844;
	wire [4-1:0] node14848;
	wire [4-1:0] node14851;
	wire [4-1:0] node14852;
	wire [4-1:0] node14853;
	wire [4-1:0] node14857;
	wire [4-1:0] node14858;
	wire [4-1:0] node14862;
	wire [4-1:0] node14863;
	wire [4-1:0] node14864;
	wire [4-1:0] node14865;
	wire [4-1:0] node14866;
	wire [4-1:0] node14869;
	wire [4-1:0] node14872;
	wire [4-1:0] node14873;
	wire [4-1:0] node14876;
	wire [4-1:0] node14879;
	wire [4-1:0] node14880;
	wire [4-1:0] node14883;
	wire [4-1:0] node14886;
	wire [4-1:0] node14887;
	wire [4-1:0] node14890;
	wire [4-1:0] node14893;
	wire [4-1:0] node14894;
	wire [4-1:0] node14895;
	wire [4-1:0] node14896;
	wire [4-1:0] node14898;
	wire [4-1:0] node14901;
	wire [4-1:0] node14903;
	wire [4-1:0] node14906;
	wire [4-1:0] node14907;
	wire [4-1:0] node14909;
	wire [4-1:0] node14912;
	wire [4-1:0] node14914;
	wire [4-1:0] node14917;
	wire [4-1:0] node14918;
	wire [4-1:0] node14919;
	wire [4-1:0] node14922;
	wire [4-1:0] node14925;
	wire [4-1:0] node14926;
	wire [4-1:0] node14927;
	wire [4-1:0] node14930;
	wire [4-1:0] node14933;
	wire [4-1:0] node14934;
	wire [4-1:0] node14937;
	wire [4-1:0] node14940;
	wire [4-1:0] node14941;
	wire [4-1:0] node14942;
	wire [4-1:0] node14943;
	wire [4-1:0] node14944;
	wire [4-1:0] node14945;
	wire [4-1:0] node14946;
	wire [4-1:0] node14950;
	wire [4-1:0] node14951;
	wire [4-1:0] node14955;
	wire [4-1:0] node14956;
	wire [4-1:0] node14957;
	wire [4-1:0] node14961;
	wire [4-1:0] node14962;
	wire [4-1:0] node14966;
	wire [4-1:0] node14967;
	wire [4-1:0] node14968;
	wire [4-1:0] node14969;
	wire [4-1:0] node14973;
	wire [4-1:0] node14974;
	wire [4-1:0] node14978;
	wire [4-1:0] node14979;
	wire [4-1:0] node14980;
	wire [4-1:0] node14984;
	wire [4-1:0] node14985;
	wire [4-1:0] node14989;
	wire [4-1:0] node14990;
	wire [4-1:0] node14991;
	wire [4-1:0] node14992;
	wire [4-1:0] node14993;
	wire [4-1:0] node14994;
	wire [4-1:0] node14997;
	wire [4-1:0] node15000;
	wire [4-1:0] node15001;
	wire [4-1:0] node15004;
	wire [4-1:0] node15007;
	wire [4-1:0] node15008;
	wire [4-1:0] node15011;
	wire [4-1:0] node15014;
	wire [4-1:0] node15015;
	wire [4-1:0] node15016;
	wire [4-1:0] node15019;
	wire [4-1:0] node15022;
	wire [4-1:0] node15023;
	wire [4-1:0] node15026;
	wire [4-1:0] node15029;
	wire [4-1:0] node15030;
	wire [4-1:0] node15031;
	wire [4-1:0] node15032;
	wire [4-1:0] node15035;
	wire [4-1:0] node15038;
	wire [4-1:0] node15039;
	wire [4-1:0] node15040;
	wire [4-1:0] node15043;
	wire [4-1:0] node15046;
	wire [4-1:0] node15047;
	wire [4-1:0] node15050;
	wire [4-1:0] node15053;
	wire [4-1:0] node15054;
	wire [4-1:0] node15055;
	wire [4-1:0] node15057;
	wire [4-1:0] node15060;
	wire [4-1:0] node15061;
	wire [4-1:0] node15064;
	wire [4-1:0] node15067;
	wire [4-1:0] node15068;
	wire [4-1:0] node15071;
	wire [4-1:0] node15074;
	wire [4-1:0] node15075;
	wire [4-1:0] node15076;
	wire [4-1:0] node15077;
	wire [4-1:0] node15078;
	wire [4-1:0] node15079;
	wire [4-1:0] node15080;
	wire [4-1:0] node15083;
	wire [4-1:0] node15087;
	wire [4-1:0] node15088;
	wire [4-1:0] node15091;
	wire [4-1:0] node15094;
	wire [4-1:0] node15095;
	wire [4-1:0] node15098;
	wire [4-1:0] node15101;
	wire [4-1:0] node15102;
	wire [4-1:0] node15103;
	wire [4-1:0] node15104;
	wire [4-1:0] node15108;
	wire [4-1:0] node15109;
	wire [4-1:0] node15113;
	wire [4-1:0] node15114;
	wire [4-1:0] node15117;
	wire [4-1:0] node15119;
	wire [4-1:0] node15122;
	wire [4-1:0] node15123;
	wire [4-1:0] node15124;
	wire [4-1:0] node15125;
	wire [4-1:0] node15126;
	wire [4-1:0] node15128;
	wire [4-1:0] node15131;
	wire [4-1:0] node15134;
	wire [4-1:0] node15135;
	wire [4-1:0] node15137;
	wire [4-1:0] node15140;
	wire [4-1:0] node15142;
	wire [4-1:0] node15145;
	wire [4-1:0] node15146;
	wire [4-1:0] node15147;
	wire [4-1:0] node15150;
	wire [4-1:0] node15153;
	wire [4-1:0] node15154;
	wire [4-1:0] node15155;
	wire [4-1:0] node15158;
	wire [4-1:0] node15161;
	wire [4-1:0] node15162;
	wire [4-1:0] node15165;
	wire [4-1:0] node15168;
	wire [4-1:0] node15169;
	wire [4-1:0] node15170;
	wire [4-1:0] node15171;
	wire [4-1:0] node15175;
	wire [4-1:0] node15176;
	wire [4-1:0] node15180;
	wire [4-1:0] node15181;
	wire [4-1:0] node15182;
	wire [4-1:0] node15186;
	wire [4-1:0] node15187;
	wire [4-1:0] node15191;
	wire [4-1:0] node15192;
	wire [4-1:0] node15193;
	wire [4-1:0] node15194;
	wire [4-1:0] node15195;
	wire [4-1:0] node15196;
	wire [4-1:0] node15197;
	wire [4-1:0] node15198;
	wire [4-1:0] node15202;
	wire [4-1:0] node15203;
	wire [4-1:0] node15207;
	wire [4-1:0] node15208;
	wire [4-1:0] node15210;
	wire [4-1:0] node15213;
	wire [4-1:0] node15214;
	wire [4-1:0] node15218;
	wire [4-1:0] node15219;
	wire [4-1:0] node15220;
	wire [4-1:0] node15222;
	wire [4-1:0] node15225;
	wire [4-1:0] node15226;
	wire [4-1:0] node15230;
	wire [4-1:0] node15231;
	wire [4-1:0] node15232;
	wire [4-1:0] node15236;
	wire [4-1:0] node15238;
	wire [4-1:0] node15241;
	wire [4-1:0] node15242;
	wire [4-1:0] node15243;
	wire [4-1:0] node15244;
	wire [4-1:0] node15247;
	wire [4-1:0] node15248;
	wire [4-1:0] node15252;
	wire [4-1:0] node15253;
	wire [4-1:0] node15254;
	wire [4-1:0] node15258;
	wire [4-1:0] node15259;
	wire [4-1:0] node15263;
	wire [4-1:0] node15264;
	wire [4-1:0] node15265;
	wire [4-1:0] node15268;
	wire [4-1:0] node15271;
	wire [4-1:0] node15272;
	wire [4-1:0] node15273;
	wire [4-1:0] node15274;
	wire [4-1:0] node15277;
	wire [4-1:0] node15280;
	wire [4-1:0] node15282;
	wire [4-1:0] node15285;
	wire [4-1:0] node15286;
	wire [4-1:0] node15287;
	wire [4-1:0] node15290;
	wire [4-1:0] node15293;
	wire [4-1:0] node15294;
	wire [4-1:0] node15297;
	wire [4-1:0] node15300;
	wire [4-1:0] node15301;
	wire [4-1:0] node15302;
	wire [4-1:0] node15303;
	wire [4-1:0] node15304;
	wire [4-1:0] node15305;
	wire [4-1:0] node15306;
	wire [4-1:0] node15311;
	wire [4-1:0] node15313;
	wire [4-1:0] node15314;
	wire [4-1:0] node15317;
	wire [4-1:0] node15320;
	wire [4-1:0] node15321;
	wire [4-1:0] node15322;
	wire [4-1:0] node15323;
	wire [4-1:0] node15326;
	wire [4-1:0] node15330;
	wire [4-1:0] node15331;
	wire [4-1:0] node15332;
	wire [4-1:0] node15335;
	wire [4-1:0] node15338;
	wire [4-1:0] node15340;
	wire [4-1:0] node15343;
	wire [4-1:0] node15344;
	wire [4-1:0] node15345;
	wire [4-1:0] node15347;
	wire [4-1:0] node15350;
	wire [4-1:0] node15351;
	wire [4-1:0] node15355;
	wire [4-1:0] node15356;
	wire [4-1:0] node15357;
	wire [4-1:0] node15361;
	wire [4-1:0] node15362;
	wire [4-1:0] node15366;
	wire [4-1:0] node15367;
	wire [4-1:0] node15368;
	wire [4-1:0] node15369;
	wire [4-1:0] node15370;
	wire [4-1:0] node15373;
	wire [4-1:0] node15376;
	wire [4-1:0] node15377;
	wire [4-1:0] node15378;
	wire [4-1:0] node15381;
	wire [4-1:0] node15384;
	wire [4-1:0] node15385;
	wire [4-1:0] node15388;
	wire [4-1:0] node15391;
	wire [4-1:0] node15392;
	wire [4-1:0] node15393;
	wire [4-1:0] node15394;
	wire [4-1:0] node15398;
	wire [4-1:0] node15399;
	wire [4-1:0] node15403;
	wire [4-1:0] node15404;
	wire [4-1:0] node15405;
	wire [4-1:0] node15410;
	wire [4-1:0] node15411;
	wire [4-1:0] node15412;
	wire [4-1:0] node15413;
	wire [4-1:0] node15416;
	wire [4-1:0] node15419;
	wire [4-1:0] node15420;
	wire [4-1:0] node15421;
	wire [4-1:0] node15424;
	wire [4-1:0] node15427;
	wire [4-1:0] node15428;
	wire [4-1:0] node15431;
	wire [4-1:0] node15434;
	wire [4-1:0] node15435;
	wire [4-1:0] node15437;
	wire [4-1:0] node15438;
	wire [4-1:0] node15442;
	wire [4-1:0] node15443;
	wire [4-1:0] node15444;
	wire [4-1:0] node15448;
	wire [4-1:0] node15449;
	wire [4-1:0] node15453;
	wire [4-1:0] node15454;
	wire [4-1:0] node15455;
	wire [4-1:0] node15456;
	wire [4-1:0] node15457;
	wire [4-1:0] node15458;
	wire [4-1:0] node15459;
	wire [4-1:0] node15460;
	wire [4-1:0] node15463;
	wire [4-1:0] node15466;
	wire [4-1:0] node15467;
	wire [4-1:0] node15470;
	wire [4-1:0] node15473;
	wire [4-1:0] node15474;
	wire [4-1:0] node15476;
	wire [4-1:0] node15479;
	wire [4-1:0] node15480;
	wire [4-1:0] node15483;
	wire [4-1:0] node15486;
	wire [4-1:0] node15487;
	wire [4-1:0] node15488;
	wire [4-1:0] node15491;
	wire [4-1:0] node15494;
	wire [4-1:0] node15496;
	wire [4-1:0] node15497;
	wire [4-1:0] node15500;
	wire [4-1:0] node15503;
	wire [4-1:0] node15504;
	wire [4-1:0] node15505;
	wire [4-1:0] node15507;
	wire [4-1:0] node15508;
	wire [4-1:0] node15511;
	wire [4-1:0] node15514;
	wire [4-1:0] node15515;
	wire [4-1:0] node15516;
	wire [4-1:0] node15519;
	wire [4-1:0] node15522;
	wire [4-1:0] node15523;
	wire [4-1:0] node15526;
	wire [4-1:0] node15529;
	wire [4-1:0] node15530;
	wire [4-1:0] node15531;
	wire [4-1:0] node15532;
	wire [4-1:0] node15535;
	wire [4-1:0] node15538;
	wire [4-1:0] node15540;
	wire [4-1:0] node15543;
	wire [4-1:0] node15544;
	wire [4-1:0] node15546;
	wire [4-1:0] node15549;
	wire [4-1:0] node15550;
	wire [4-1:0] node15553;
	wire [4-1:0] node15556;
	wire [4-1:0] node15557;
	wire [4-1:0] node15558;
	wire [4-1:0] node15559;
	wire [4-1:0] node15562;
	wire [4-1:0] node15565;
	wire [4-1:0] node15566;
	wire [4-1:0] node15567;
	wire [4-1:0] node15570;
	wire [4-1:0] node15573;
	wire [4-1:0] node15574;
	wire [4-1:0] node15575;
	wire [4-1:0] node15580;
	wire [4-1:0] node15581;
	wire [4-1:0] node15583;
	wire [4-1:0] node15584;
	wire [4-1:0] node15587;
	wire [4-1:0] node15590;
	wire [4-1:0] node15591;
	wire [4-1:0] node15592;
	wire [4-1:0] node15593;
	wire [4-1:0] node15596;
	wire [4-1:0] node15599;
	wire [4-1:0] node15600;
	wire [4-1:0] node15603;
	wire [4-1:0] node15606;
	wire [4-1:0] node15607;
	wire [4-1:0] node15610;
	wire [4-1:0] node15613;
	wire [4-1:0] node15614;
	wire [4-1:0] node15615;
	wire [4-1:0] node15616;
	wire [4-1:0] node15617;
	wire [4-1:0] node15620;
	wire [4-1:0] node15624;
	wire [4-1:0] node15625;
	wire [4-1:0] node15626;
	wire [4-1:0] node15627;
	wire [4-1:0] node15630;
	wire [4-1:0] node15633;
	wire [4-1:0] node15634;
	wire [4-1:0] node15639;
	wire [4-1:0] node15640;
	wire [4-1:0] node15641;
	wire [4-1:0] node15642;
	wire [4-1:0] node15643;
	wire [4-1:0] node15646;
	wire [4-1:0] node15649;
	wire [4-1:0] node15650;
	wire [4-1:0] node15653;
	wire [4-1:0] node15657;
	wire [4-1:0] node15658;
	wire [4-1:0] node15659;
	wire [4-1:0] node15660;
	wire [4-1:0] node15662;
	wire [4-1:0] node15665;
	wire [4-1:0] node15666;
	wire [4-1:0] node15669;
	wire [4-1:0] node15672;
	wire [4-1:0] node15673;
	wire [4-1:0] node15674;
	wire [4-1:0] node15677;
	wire [4-1:0] node15680;
	wire [4-1:0] node15681;
	wire [4-1:0] node15684;
	wire [4-1:0] node15688;
	wire [4-1:0] node15689;
	wire [4-1:0] node15690;
	wire [4-1:0] node15691;
	wire [4-1:0] node15692;
	wire [4-1:0] node15693;
	wire [4-1:0] node15694;
	wire [4-1:0] node15695;
	wire [4-1:0] node15696;
	wire [4-1:0] node15697;
	wire [4-1:0] node15698;
	wire [4-1:0] node15702;
	wire [4-1:0] node15703;
	wire [4-1:0] node15707;
	wire [4-1:0] node15708;
	wire [4-1:0] node15709;
	wire [4-1:0] node15713;
	wire [4-1:0] node15715;
	wire [4-1:0] node15718;
	wire [4-1:0] node15719;
	wire [4-1:0] node15720;
	wire [4-1:0] node15721;
	wire [4-1:0] node15724;
	wire [4-1:0] node15728;
	wire [4-1:0] node15729;
	wire [4-1:0] node15732;
	wire [4-1:0] node15734;
	wire [4-1:0] node15737;
	wire [4-1:0] node15738;
	wire [4-1:0] node15739;
	wire [4-1:0] node15740;
	wire [4-1:0] node15742;
	wire [4-1:0] node15745;
	wire [4-1:0] node15747;
	wire [4-1:0] node15750;
	wire [4-1:0] node15751;
	wire [4-1:0] node15753;
	wire [4-1:0] node15756;
	wire [4-1:0] node15757;
	wire [4-1:0] node15761;
	wire [4-1:0] node15762;
	wire [4-1:0] node15763;
	wire [4-1:0] node15764;
	wire [4-1:0] node15768;
	wire [4-1:0] node15769;
	wire [4-1:0] node15773;
	wire [4-1:0] node15774;
	wire [4-1:0] node15776;
	wire [4-1:0] node15779;
	wire [4-1:0] node15780;
	wire [4-1:0] node15784;
	wire [4-1:0] node15785;
	wire [4-1:0] node15786;
	wire [4-1:0] node15787;
	wire [4-1:0] node15788;
	wire [4-1:0] node15791;
	wire [4-1:0] node15794;
	wire [4-1:0] node15795;
	wire [4-1:0] node15798;
	wire [4-1:0] node15801;
	wire [4-1:0] node15802;
	wire [4-1:0] node15803;
	wire [4-1:0] node15804;
	wire [4-1:0] node15807;
	wire [4-1:0] node15810;
	wire [4-1:0] node15811;
	wire [4-1:0] node15814;
	wire [4-1:0] node15817;
	wire [4-1:0] node15819;
	wire [4-1:0] node15820;
	wire [4-1:0] node15823;
	wire [4-1:0] node15826;
	wire [4-1:0] node15827;
	wire [4-1:0] node15828;
	wire [4-1:0] node15829;
	wire [4-1:0] node15830;
	wire [4-1:0] node15834;
	wire [4-1:0] node15835;
	wire [4-1:0] node15839;
	wire [4-1:0] node15840;
	wire [4-1:0] node15842;
	wire [4-1:0] node15845;
	wire [4-1:0] node15848;
	wire [4-1:0] node15849;
	wire [4-1:0] node15850;
	wire [4-1:0] node15851;
	wire [4-1:0] node15854;
	wire [4-1:0] node15857;
	wire [4-1:0] node15858;
	wire [4-1:0] node15862;
	wire [4-1:0] node15863;
	wire [4-1:0] node15866;
	wire [4-1:0] node15869;
	wire [4-1:0] node15870;
	wire [4-1:0] node15871;
	wire [4-1:0] node15872;
	wire [4-1:0] node15873;
	wire [4-1:0] node15874;
	wire [4-1:0] node15877;
	wire [4-1:0] node15880;
	wire [4-1:0] node15882;
	wire [4-1:0] node15884;
	wire [4-1:0] node15887;
	wire [4-1:0] node15888;
	wire [4-1:0] node15889;
	wire [4-1:0] node15891;
	wire [4-1:0] node15894;
	wire [4-1:0] node15895;
	wire [4-1:0] node15898;
	wire [4-1:0] node15901;
	wire [4-1:0] node15902;
	wire [4-1:0] node15905;
	wire [4-1:0] node15908;
	wire [4-1:0] node15909;
	wire [4-1:0] node15910;
	wire [4-1:0] node15911;
	wire [4-1:0] node15912;
	wire [4-1:0] node15915;
	wire [4-1:0] node15918;
	wire [4-1:0] node15919;
	wire [4-1:0] node15922;
	wire [4-1:0] node15925;
	wire [4-1:0] node15926;
	wire [4-1:0] node15927;
	wire [4-1:0] node15930;
	wire [4-1:0] node15933;
	wire [4-1:0] node15934;
	wire [4-1:0] node15937;
	wire [4-1:0] node15940;
	wire [4-1:0] node15941;
	wire [4-1:0] node15942;
	wire [4-1:0] node15943;
	wire [4-1:0] node15946;
	wire [4-1:0] node15949;
	wire [4-1:0] node15950;
	wire [4-1:0] node15953;
	wire [4-1:0] node15956;
	wire [4-1:0] node15957;
	wire [4-1:0] node15960;
	wire [4-1:0] node15963;
	wire [4-1:0] node15964;
	wire [4-1:0] node15965;
	wire [4-1:0] node15966;
	wire [4-1:0] node15967;
	wire [4-1:0] node15968;
	wire [4-1:0] node15971;
	wire [4-1:0] node15974;
	wire [4-1:0] node15975;
	wire [4-1:0] node15978;
	wire [4-1:0] node15981;
	wire [4-1:0] node15982;
	wire [4-1:0] node15983;
	wire [4-1:0] node15986;
	wire [4-1:0] node15989;
	wire [4-1:0] node15991;
	wire [4-1:0] node15994;
	wire [4-1:0] node15995;
	wire [4-1:0] node15996;
	wire [4-1:0] node15997;
	wire [4-1:0] node16000;
	wire [4-1:0] node16003;
	wire [4-1:0] node16004;
	wire [4-1:0] node16007;
	wire [4-1:0] node16010;
	wire [4-1:0] node16011;
	wire [4-1:0] node16014;
	wire [4-1:0] node16017;
	wire [4-1:0] node16018;
	wire [4-1:0] node16019;
	wire [4-1:0] node16022;
	wire [4-1:0] node16025;
	wire [4-1:0] node16026;
	wire [4-1:0] node16027;
	wire [4-1:0] node16029;
	wire [4-1:0] node16032;
	wire [4-1:0] node16035;
	wire [4-1:0] node16036;
	wire [4-1:0] node16039;
	wire [4-1:0] node16042;
	wire [4-1:0] node16043;
	wire [4-1:0] node16044;
	wire [4-1:0] node16045;
	wire [4-1:0] node16046;
	wire [4-1:0] node16047;
	wire [4-1:0] node16048;
	wire [4-1:0] node16051;
	wire [4-1:0] node16054;
	wire [4-1:0] node16055;
	wire [4-1:0] node16058;
	wire [4-1:0] node16061;
	wire [4-1:0] node16062;
	wire [4-1:0] node16063;
	wire [4-1:0] node16066;
	wire [4-1:0] node16069;
	wire [4-1:0] node16070;
	wire [4-1:0] node16073;
	wire [4-1:0] node16076;
	wire [4-1:0] node16077;
	wire [4-1:0] node16078;
	wire [4-1:0] node16079;
	wire [4-1:0] node16080;
	wire [4-1:0] node16083;
	wire [4-1:0] node16086;
	wire [4-1:0] node16088;
	wire [4-1:0] node16091;
	wire [4-1:0] node16092;
	wire [4-1:0] node16093;
	wire [4-1:0] node16096;
	wire [4-1:0] node16099;
	wire [4-1:0] node16100;
	wire [4-1:0] node16103;
	wire [4-1:0] node16106;
	wire [4-1:0] node16107;
	wire [4-1:0] node16108;
	wire [4-1:0] node16109;
	wire [4-1:0] node16112;
	wire [4-1:0] node16115;
	wire [4-1:0] node16116;
	wire [4-1:0] node16119;
	wire [4-1:0] node16122;
	wire [4-1:0] node16124;
	wire [4-1:0] node16125;
	wire [4-1:0] node16128;
	wire [4-1:0] node16131;
	wire [4-1:0] node16132;
	wire [4-1:0] node16133;
	wire [4-1:0] node16134;
	wire [4-1:0] node16135;
	wire [4-1:0] node16136;
	wire [4-1:0] node16140;
	wire [4-1:0] node16141;
	wire [4-1:0] node16145;
	wire [4-1:0] node16147;
	wire [4-1:0] node16150;
	wire [4-1:0] node16151;
	wire [4-1:0] node16153;
	wire [4-1:0] node16154;
	wire [4-1:0] node16158;
	wire [4-1:0] node16159;
	wire [4-1:0] node16161;
	wire [4-1:0] node16164;
	wire [4-1:0] node16166;
	wire [4-1:0] node16169;
	wire [4-1:0] node16170;
	wire [4-1:0] node16171;
	wire [4-1:0] node16172;
	wire [4-1:0] node16173;
	wire [4-1:0] node16178;
	wire [4-1:0] node16179;
	wire [4-1:0] node16182;
	wire [4-1:0] node16185;
	wire [4-1:0] node16186;
	wire [4-1:0] node16187;
	wire [4-1:0] node16190;
	wire [4-1:0] node16191;
	wire [4-1:0] node16195;
	wire [4-1:0] node16196;
	wire [4-1:0] node16198;
	wire [4-1:0] node16202;
	wire [4-1:0] node16203;
	wire [4-1:0] node16204;
	wire [4-1:0] node16205;
	wire [4-1:0] node16206;
	wire [4-1:0] node16207;
	wire [4-1:0] node16208;
	wire [4-1:0] node16212;
	wire [4-1:0] node16213;
	wire [4-1:0] node16217;
	wire [4-1:0] node16219;
	wire [4-1:0] node16222;
	wire [4-1:0] node16223;
	wire [4-1:0] node16224;
	wire [4-1:0] node16225;
	wire [4-1:0] node16230;
	wire [4-1:0] node16231;
	wire [4-1:0] node16233;
	wire [4-1:0] node16236;
	wire [4-1:0] node16237;
	wire [4-1:0] node16241;
	wire [4-1:0] node16242;
	wire [4-1:0] node16243;
	wire [4-1:0] node16244;
	wire [4-1:0] node16247;
	wire [4-1:0] node16250;
	wire [4-1:0] node16251;
	wire [4-1:0] node16252;
	wire [4-1:0] node16255;
	wire [4-1:0] node16258;
	wire [4-1:0] node16260;
	wire [4-1:0] node16263;
	wire [4-1:0] node16264;
	wire [4-1:0] node16267;
	wire [4-1:0] node16270;
	wire [4-1:0] node16271;
	wire [4-1:0] node16272;
	wire [4-1:0] node16273;
	wire [4-1:0] node16275;
	wire [4-1:0] node16276;
	wire [4-1:0] node16280;
	wire [4-1:0] node16281;
	wire [4-1:0] node16282;
	wire [4-1:0] node16286;
	wire [4-1:0] node16288;
	wire [4-1:0] node16291;
	wire [4-1:0] node16292;
	wire [4-1:0] node16293;
	wire [4-1:0] node16294;
	wire [4-1:0] node16298;
	wire [4-1:0] node16299;
	wire [4-1:0] node16303;
	wire [4-1:0] node16305;
	wire [4-1:0] node16307;
	wire [4-1:0] node16310;
	wire [4-1:0] node16311;
	wire [4-1:0] node16312;
	wire [4-1:0] node16313;
	wire [4-1:0] node16317;
	wire [4-1:0] node16319;
	wire [4-1:0] node16322;
	wire [4-1:0] node16323;
	wire [4-1:0] node16325;
	wire [4-1:0] node16328;
	wire [4-1:0] node16329;
	wire [4-1:0] node16333;
	wire [4-1:0] node16334;
	wire [4-1:0] node16335;
	wire [4-1:0] node16336;
	wire [4-1:0] node16337;
	wire [4-1:0] node16338;
	wire [4-1:0] node16339;
	wire [4-1:0] node16340;
	wire [4-1:0] node16343;
	wire [4-1:0] node16346;
	wire [4-1:0] node16347;
	wire [4-1:0] node16348;
	wire [4-1:0] node16351;
	wire [4-1:0] node16354;
	wire [4-1:0] node16355;
	wire [4-1:0] node16358;
	wire [4-1:0] node16361;
	wire [4-1:0] node16362;
	wire [4-1:0] node16363;
	wire [4-1:0] node16364;
	wire [4-1:0] node16368;
	wire [4-1:0] node16369;
	wire [4-1:0] node16373;
	wire [4-1:0] node16374;
	wire [4-1:0] node16375;
	wire [4-1:0] node16379;
	wire [4-1:0] node16380;
	wire [4-1:0] node16384;
	wire [4-1:0] node16385;
	wire [4-1:0] node16386;
	wire [4-1:0] node16387;
	wire [4-1:0] node16388;
	wire [4-1:0] node16391;
	wire [4-1:0] node16394;
	wire [4-1:0] node16395;
	wire [4-1:0] node16398;
	wire [4-1:0] node16401;
	wire [4-1:0] node16402;
	wire [4-1:0] node16403;
	wire [4-1:0] node16406;
	wire [4-1:0] node16410;
	wire [4-1:0] node16411;
	wire [4-1:0] node16412;
	wire [4-1:0] node16414;
	wire [4-1:0] node16417;
	wire [4-1:0] node16419;
	wire [4-1:0] node16422;
	wire [4-1:0] node16423;
	wire [4-1:0] node16425;
	wire [4-1:0] node16428;
	wire [4-1:0] node16431;
	wire [4-1:0] node16432;
	wire [4-1:0] node16433;
	wire [4-1:0] node16434;
	wire [4-1:0] node16435;
	wire [4-1:0] node16439;
	wire [4-1:0] node16440;
	wire [4-1:0] node16441;
	wire [4-1:0] node16444;
	wire [4-1:0] node16447;
	wire [4-1:0] node16448;
	wire [4-1:0] node16452;
	wire [4-1:0] node16453;
	wire [4-1:0] node16454;
	wire [4-1:0] node16456;
	wire [4-1:0] node16459;
	wire [4-1:0] node16460;
	wire [4-1:0] node16464;
	wire [4-1:0] node16465;
	wire [4-1:0] node16468;
	wire [4-1:0] node16469;
	wire [4-1:0] node16473;
	wire [4-1:0] node16474;
	wire [4-1:0] node16475;
	wire [4-1:0] node16476;
	wire [4-1:0] node16479;
	wire [4-1:0] node16482;
	wire [4-1:0] node16483;
	wire [4-1:0] node16485;
	wire [4-1:0] node16488;
	wire [4-1:0] node16489;
	wire [4-1:0] node16492;
	wire [4-1:0] node16495;
	wire [4-1:0] node16496;
	wire [4-1:0] node16498;
	wire [4-1:0] node16499;
	wire [4-1:0] node16502;
	wire [4-1:0] node16505;
	wire [4-1:0] node16506;
	wire [4-1:0] node16507;
	wire [4-1:0] node16510;
	wire [4-1:0] node16513;
	wire [4-1:0] node16514;
	wire [4-1:0] node16517;
	wire [4-1:0] node16520;
	wire [4-1:0] node16521;
	wire [4-1:0] node16522;
	wire [4-1:0] node16523;
	wire [4-1:0] node16524;
	wire [4-1:0] node16525;
	wire [4-1:0] node16528;
	wire [4-1:0] node16529;
	wire [4-1:0] node16533;
	wire [4-1:0] node16534;
	wire [4-1:0] node16535;
	wire [4-1:0] node16539;
	wire [4-1:0] node16542;
	wire [4-1:0] node16543;
	wire [4-1:0] node16544;
	wire [4-1:0] node16547;
	wire [4-1:0] node16549;
	wire [4-1:0] node16552;
	wire [4-1:0] node16554;
	wire [4-1:0] node16556;
	wire [4-1:0] node16559;
	wire [4-1:0] node16560;
	wire [4-1:0] node16561;
	wire [4-1:0] node16562;
	wire [4-1:0] node16563;
	wire [4-1:0] node16567;
	wire [4-1:0] node16569;
	wire [4-1:0] node16572;
	wire [4-1:0] node16573;
	wire [4-1:0] node16575;
	wire [4-1:0] node16578;
	wire [4-1:0] node16579;
	wire [4-1:0] node16583;
	wire [4-1:0] node16584;
	wire [4-1:0] node16585;
	wire [4-1:0] node16586;
	wire [4-1:0] node16590;
	wire [4-1:0] node16593;
	wire [4-1:0] node16594;
	wire [4-1:0] node16595;
	wire [4-1:0] node16600;
	wire [4-1:0] node16601;
	wire [4-1:0] node16602;
	wire [4-1:0] node16603;
	wire [4-1:0] node16604;
	wire [4-1:0] node16605;
	wire [4-1:0] node16610;
	wire [4-1:0] node16611;
	wire [4-1:0] node16613;
	wire [4-1:0] node16616;
	wire [4-1:0] node16617;
	wire [4-1:0] node16621;
	wire [4-1:0] node16622;
	wire [4-1:0] node16623;
	wire [4-1:0] node16625;
	wire [4-1:0] node16629;
	wire [4-1:0] node16630;
	wire [4-1:0] node16631;
	wire [4-1:0] node16635;
	wire [4-1:0] node16637;
	wire [4-1:0] node16640;
	wire [4-1:0] node16641;
	wire [4-1:0] node16642;
	wire [4-1:0] node16643;
	wire [4-1:0] node16644;
	wire [4-1:0] node16648;
	wire [4-1:0] node16651;
	wire [4-1:0] node16653;
	wire [4-1:0] node16654;
	wire [4-1:0] node16658;
	wire [4-1:0] node16659;
	wire [4-1:0] node16660;
	wire [4-1:0] node16661;
	wire [4-1:0] node16664;
	wire [4-1:0] node16667;
	wire [4-1:0] node16668;
	wire [4-1:0] node16671;
	wire [4-1:0] node16674;
	wire [4-1:0] node16676;
	wire [4-1:0] node16677;
	wire [4-1:0] node16680;
	wire [4-1:0] node16683;
	wire [4-1:0] node16684;
	wire [4-1:0] node16685;
	wire [4-1:0] node16686;
	wire [4-1:0] node16687;
	wire [4-1:0] node16688;
	wire [4-1:0] node16689;
	wire [4-1:0] node16690;
	wire [4-1:0] node16693;
	wire [4-1:0] node16696;
	wire [4-1:0] node16697;
	wire [4-1:0] node16701;
	wire [4-1:0] node16702;
	wire [4-1:0] node16703;
	wire [4-1:0] node16706;
	wire [4-1:0] node16709;
	wire [4-1:0] node16710;
	wire [4-1:0] node16713;
	wire [4-1:0] node16716;
	wire [4-1:0] node16717;
	wire [4-1:0] node16718;
	wire [4-1:0] node16720;
	wire [4-1:0] node16723;
	wire [4-1:0] node16725;
	wire [4-1:0] node16728;
	wire [4-1:0] node16730;
	wire [4-1:0] node16733;
	wire [4-1:0] node16734;
	wire [4-1:0] node16735;
	wire [4-1:0] node16736;
	wire [4-1:0] node16737;
	wire [4-1:0] node16740;
	wire [4-1:0] node16743;
	wire [4-1:0] node16744;
	wire [4-1:0] node16747;
	wire [4-1:0] node16750;
	wire [4-1:0] node16751;
	wire [4-1:0] node16752;
	wire [4-1:0] node16756;
	wire [4-1:0] node16757;
	wire [4-1:0] node16760;
	wire [4-1:0] node16763;
	wire [4-1:0] node16764;
	wire [4-1:0] node16765;
	wire [4-1:0] node16768;
	wire [4-1:0] node16771;
	wire [4-1:0] node16772;
	wire [4-1:0] node16775;
	wire [4-1:0] node16778;
	wire [4-1:0] node16779;
	wire [4-1:0] node16780;
	wire [4-1:0] node16781;
	wire [4-1:0] node16782;
	wire [4-1:0] node16784;
	wire [4-1:0] node16787;
	wire [4-1:0] node16789;
	wire [4-1:0] node16792;
	wire [4-1:0] node16793;
	wire [4-1:0] node16796;
	wire [4-1:0] node16798;
	wire [4-1:0] node16801;
	wire [4-1:0] node16802;
	wire [4-1:0] node16803;
	wire [4-1:0] node16804;
	wire [4-1:0] node16807;
	wire [4-1:0] node16810;
	wire [4-1:0] node16811;
	wire [4-1:0] node16814;
	wire [4-1:0] node16817;
	wire [4-1:0] node16819;
	wire [4-1:0] node16820;
	wire [4-1:0] node16823;
	wire [4-1:0] node16826;
	wire [4-1:0] node16827;
	wire [4-1:0] node16828;
	wire [4-1:0] node16830;
	wire [4-1:0] node16833;
	wire [4-1:0] node16835;
	wire [4-1:0] node16838;
	wire [4-1:0] node16839;
	wire [4-1:0] node16841;
	wire [4-1:0] node16844;
	wire [4-1:0] node16845;
	wire [4-1:0] node16849;
	wire [4-1:0] node16850;
	wire [4-1:0] node16851;
	wire [4-1:0] node16852;
	wire [4-1:0] node16853;
	wire [4-1:0] node16854;
	wire [4-1:0] node16856;
	wire [4-1:0] node16859;
	wire [4-1:0] node16860;
	wire [4-1:0] node16864;
	wire [4-1:0] node16865;
	wire [4-1:0] node16868;
	wire [4-1:0] node16869;
	wire [4-1:0] node16873;
	wire [4-1:0] node16874;
	wire [4-1:0] node16876;
	wire [4-1:0] node16877;
	wire [4-1:0] node16881;
	wire [4-1:0] node16882;
	wire [4-1:0] node16885;
	wire [4-1:0] node16886;
	wire [4-1:0] node16890;
	wire [4-1:0] node16891;
	wire [4-1:0] node16892;
	wire [4-1:0] node16893;
	wire [4-1:0] node16894;
	wire [4-1:0] node16897;
	wire [4-1:0] node16900;
	wire [4-1:0] node16902;
	wire [4-1:0] node16905;
	wire [4-1:0] node16906;
	wire [4-1:0] node16907;
	wire [4-1:0] node16910;
	wire [4-1:0] node16913;
	wire [4-1:0] node16915;
	wire [4-1:0] node16918;
	wire [4-1:0] node16919;
	wire [4-1:0] node16920;
	wire [4-1:0] node16921;
	wire [4-1:0] node16925;
	wire [4-1:0] node16926;
	wire [4-1:0] node16930;
	wire [4-1:0] node16931;
	wire [4-1:0] node16932;
	wire [4-1:0] node16936;
	wire [4-1:0] node16937;
	wire [4-1:0] node16941;
	wire [4-1:0] node16942;
	wire [4-1:0] node16943;
	wire [4-1:0] node16944;
	wire [4-1:0] node16945;
	wire [4-1:0] node16948;
	wire [4-1:0] node16951;
	wire [4-1:0] node16952;
	wire [4-1:0] node16955;
	wire [4-1:0] node16958;
	wire [4-1:0] node16959;
	wire [4-1:0] node16960;
	wire [4-1:0] node16963;
	wire [4-1:0] node16966;
	wire [4-1:0] node16967;
	wire [4-1:0] node16970;
	wire [4-1:0] node16973;
	wire [4-1:0] node16974;
	wire [4-1:0] node16975;
	wire [4-1:0] node16978;
	wire [4-1:0] node16981;
	wire [4-1:0] node16982;
	wire [4-1:0] node16983;
	wire [4-1:0] node16984;
	wire [4-1:0] node16987;
	wire [4-1:0] node16990;
	wire [4-1:0] node16991;
	wire [4-1:0] node16994;
	wire [4-1:0] node16997;
	wire [4-1:0] node16998;
	wire [4-1:0] node17001;
	wire [4-1:0] node17004;
	wire [4-1:0] node17005;
	wire [4-1:0] node17006;
	wire [4-1:0] node17007;
	wire [4-1:0] node17008;
	wire [4-1:0] node17009;
	wire [4-1:0] node17010;
	wire [4-1:0] node17011;
	wire [4-1:0] node17012;
	wire [4-1:0] node17013;
	wire [4-1:0] node17017;
	wire [4-1:0] node17018;
	wire [4-1:0] node17021;
	wire [4-1:0] node17024;
	wire [4-1:0] node17025;
	wire [4-1:0] node17026;
	wire [4-1:0] node17029;
	wire [4-1:0] node17032;
	wire [4-1:0] node17033;
	wire [4-1:0] node17036;
	wire [4-1:0] node17039;
	wire [4-1:0] node17040;
	wire [4-1:0] node17041;
	wire [4-1:0] node17044;
	wire [4-1:0] node17047;
	wire [4-1:0] node17049;
	wire [4-1:0] node17052;
	wire [4-1:0] node17053;
	wire [4-1:0] node17054;
	wire [4-1:0] node17055;
	wire [4-1:0] node17056;
	wire [4-1:0] node17060;
	wire [4-1:0] node17063;
	wire [4-1:0] node17064;
	wire [4-1:0] node17065;
	wire [4-1:0] node17069;
	wire [4-1:0] node17071;
	wire [4-1:0] node17074;
	wire [4-1:0] node17075;
	wire [4-1:0] node17076;
	wire [4-1:0] node17077;
	wire [4-1:0] node17080;
	wire [4-1:0] node17083;
	wire [4-1:0] node17084;
	wire [4-1:0] node17087;
	wire [4-1:0] node17090;
	wire [4-1:0] node17091;
	wire [4-1:0] node17092;
	wire [4-1:0] node17095;
	wire [4-1:0] node17099;
	wire [4-1:0] node17100;
	wire [4-1:0] node17101;
	wire [4-1:0] node17102;
	wire [4-1:0] node17104;
	wire [4-1:0] node17107;
	wire [4-1:0] node17108;
	wire [4-1:0] node17112;
	wire [4-1:0] node17113;
	wire [4-1:0] node17114;
	wire [4-1:0] node17118;
	wire [4-1:0] node17119;
	wire [4-1:0] node17123;
	wire [4-1:0] node17124;
	wire [4-1:0] node17125;
	wire [4-1:0] node17126;
	wire [4-1:0] node17129;
	wire [4-1:0] node17132;
	wire [4-1:0] node17133;
	wire [4-1:0] node17134;
	wire [4-1:0] node17137;
	wire [4-1:0] node17141;
	wire [4-1:0] node17142;
	wire [4-1:0] node17143;
	wire [4-1:0] node17146;
	wire [4-1:0] node17149;
	wire [4-1:0] node17150;
	wire [4-1:0] node17151;
	wire [4-1:0] node17154;
	wire [4-1:0] node17157;
	wire [4-1:0] node17158;
	wire [4-1:0] node17161;
	wire [4-1:0] node17164;
	wire [4-1:0] node17165;
	wire [4-1:0] node17166;
	wire [4-1:0] node17167;
	wire [4-1:0] node17168;
	wire [4-1:0] node17171;
	wire [4-1:0] node17174;
	wire [4-1:0] node17175;
	wire [4-1:0] node17176;
	wire [4-1:0] node17179;
	wire [4-1:0] node17182;
	wire [4-1:0] node17184;
	wire [4-1:0] node17185;
	wire [4-1:0] node17188;
	wire [4-1:0] node17191;
	wire [4-1:0] node17192;
	wire [4-1:0] node17193;
	wire [4-1:0] node17195;
	wire [4-1:0] node17198;
	wire [4-1:0] node17199;
	wire [4-1:0] node17203;
	wire [4-1:0] node17204;
	wire [4-1:0] node17205;
	wire [4-1:0] node17209;
	wire [4-1:0] node17211;
	wire [4-1:0] node17214;
	wire [4-1:0] node17215;
	wire [4-1:0] node17216;
	wire [4-1:0] node17217;
	wire [4-1:0] node17218;
	wire [4-1:0] node17219;
	wire [4-1:0] node17222;
	wire [4-1:0] node17225;
	wire [4-1:0] node17226;
	wire [4-1:0] node17230;
	wire [4-1:0] node17231;
	wire [4-1:0] node17234;
	wire [4-1:0] node17237;
	wire [4-1:0] node17238;
	wire [4-1:0] node17239;
	wire [4-1:0] node17241;
	wire [4-1:0] node17245;
	wire [4-1:0] node17246;
	wire [4-1:0] node17247;
	wire [4-1:0] node17251;
	wire [4-1:0] node17252;
	wire [4-1:0] node17255;
	wire [4-1:0] node17258;
	wire [4-1:0] node17259;
	wire [4-1:0] node17260;
	wire [4-1:0] node17261;
	wire [4-1:0] node17265;
	wire [4-1:0] node17266;
	wire [4-1:0] node17270;
	wire [4-1:0] node17271;
	wire [4-1:0] node17272;
	wire [4-1:0] node17276;
	wire [4-1:0] node17277;
	wire [4-1:0] node17281;
	wire [4-1:0] node17282;
	wire [4-1:0] node17283;
	wire [4-1:0] node17284;
	wire [4-1:0] node17285;
	wire [4-1:0] node17286;
	wire [4-1:0] node17287;
	wire [4-1:0] node17289;
	wire [4-1:0] node17292;
	wire [4-1:0] node17293;
	wire [4-1:0] node17296;
	wire [4-1:0] node17299;
	wire [4-1:0] node17300;
	wire [4-1:0] node17302;
	wire [4-1:0] node17305;
	wire [4-1:0] node17306;
	wire [4-1:0] node17309;
	wire [4-1:0] node17312;
	wire [4-1:0] node17313;
	wire [4-1:0] node17314;
	wire [4-1:0] node17317;
	wire [4-1:0] node17320;
	wire [4-1:0] node17321;
	wire [4-1:0] node17324;
	wire [4-1:0] node17327;
	wire [4-1:0] node17328;
	wire [4-1:0] node17329;
	wire [4-1:0] node17330;
	wire [4-1:0] node17331;
	wire [4-1:0] node17334;
	wire [4-1:0] node17337;
	wire [4-1:0] node17338;
	wire [4-1:0] node17341;
	wire [4-1:0] node17344;
	wire [4-1:0] node17345;
	wire [4-1:0] node17346;
	wire [4-1:0] node17350;
	wire [4-1:0] node17351;
	wire [4-1:0] node17355;
	wire [4-1:0] node17356;
	wire [4-1:0] node17357;
	wire [4-1:0] node17358;
	wire [4-1:0] node17363;
	wire [4-1:0] node17364;
	wire [4-1:0] node17365;
	wire [4-1:0] node17368;
	wire [4-1:0] node17371;
	wire [4-1:0] node17372;
	wire [4-1:0] node17375;
	wire [4-1:0] node17378;
	wire [4-1:0] node17379;
	wire [4-1:0] node17380;
	wire [4-1:0] node17381;
	wire [4-1:0] node17383;
	wire [4-1:0] node17386;
	wire [4-1:0] node17387;
	wire [4-1:0] node17390;
	wire [4-1:0] node17393;
	wire [4-1:0] node17394;
	wire [4-1:0] node17395;
	wire [4-1:0] node17398;
	wire [4-1:0] node17401;
	wire [4-1:0] node17402;
	wire [4-1:0] node17405;
	wire [4-1:0] node17408;
	wire [4-1:0] node17409;
	wire [4-1:0] node17410;
	wire [4-1:0] node17411;
	wire [4-1:0] node17414;
	wire [4-1:0] node17417;
	wire [4-1:0] node17418;
	wire [4-1:0] node17421;
	wire [4-1:0] node17424;
	wire [4-1:0] node17425;
	wire [4-1:0] node17427;
	wire [4-1:0] node17430;
	wire [4-1:0] node17431;
	wire [4-1:0] node17434;
	wire [4-1:0] node17437;
	wire [4-1:0] node17438;
	wire [4-1:0] node17439;
	wire [4-1:0] node17440;
	wire [4-1:0] node17441;
	wire [4-1:0] node17442;
	wire [4-1:0] node17443;
	wire [4-1:0] node17446;
	wire [4-1:0] node17450;
	wire [4-1:0] node17451;
	wire [4-1:0] node17454;
	wire [4-1:0] node17457;
	wire [4-1:0] node17458;
	wire [4-1:0] node17459;
	wire [4-1:0] node17462;
	wire [4-1:0] node17465;
	wire [4-1:0] node17466;
	wire [4-1:0] node17469;
	wire [4-1:0] node17472;
	wire [4-1:0] node17473;
	wire [4-1:0] node17474;
	wire [4-1:0] node17475;
	wire [4-1:0] node17476;
	wire [4-1:0] node17480;
	wire [4-1:0] node17481;
	wire [4-1:0] node17484;
	wire [4-1:0] node17487;
	wire [4-1:0] node17488;
	wire [4-1:0] node17489;
	wire [4-1:0] node17492;
	wire [4-1:0] node17495;
	wire [4-1:0] node17496;
	wire [4-1:0] node17499;
	wire [4-1:0] node17502;
	wire [4-1:0] node17503;
	wire [4-1:0] node17504;
	wire [4-1:0] node17507;
	wire [4-1:0] node17510;
	wire [4-1:0] node17512;
	wire [4-1:0] node17515;
	wire [4-1:0] node17516;
	wire [4-1:0] node17517;
	wire [4-1:0] node17518;
	wire [4-1:0] node17520;
	wire [4-1:0] node17523;
	wire [4-1:0] node17526;
	wire [4-1:0] node17527;
	wire [4-1:0] node17528;
	wire [4-1:0] node17532;
	wire [4-1:0] node17535;
	wire [4-1:0] node17536;
	wire [4-1:0] node17537;
	wire [4-1:0] node17538;
	wire [4-1:0] node17539;
	wire [4-1:0] node17544;
	wire [4-1:0] node17545;
	wire [4-1:0] node17546;
	wire [4-1:0] node17550;
	wire [4-1:0] node17551;
	wire [4-1:0] node17555;
	wire [4-1:0] node17556;
	wire [4-1:0] node17557;
	wire [4-1:0] node17558;
	wire [4-1:0] node17561;
	wire [4-1:0] node17564;
	wire [4-1:0] node17565;
	wire [4-1:0] node17569;
	wire [4-1:0] node17570;
	wire [4-1:0] node17573;
	wire [4-1:0] node17576;
	wire [4-1:0] node17577;
	wire [4-1:0] node17578;
	wire [4-1:0] node17579;
	wire [4-1:0] node17580;
	wire [4-1:0] node17581;
	wire [4-1:0] node17582;
	wire [4-1:0] node17583;
	wire [4-1:0] node17584;
	wire [4-1:0] node17587;
	wire [4-1:0] node17590;
	wire [4-1:0] node17591;
	wire [4-1:0] node17594;
	wire [4-1:0] node17597;
	wire [4-1:0] node17598;
	wire [4-1:0] node17599;
	wire [4-1:0] node17602;
	wire [4-1:0] node17605;
	wire [4-1:0] node17607;
	wire [4-1:0] node17610;
	wire [4-1:0] node17611;
	wire [4-1:0] node17612;
	wire [4-1:0] node17614;
	wire [4-1:0] node17617;
	wire [4-1:0] node17618;
	wire [4-1:0] node17622;
	wire [4-1:0] node17623;
	wire [4-1:0] node17624;
	wire [4-1:0] node17629;
	wire [4-1:0] node17630;
	wire [4-1:0] node17631;
	wire [4-1:0] node17632;
	wire [4-1:0] node17633;
	wire [4-1:0] node17637;
	wire [4-1:0] node17640;
	wire [4-1:0] node17641;
	wire [4-1:0] node17642;
	wire [4-1:0] node17646;
	wire [4-1:0] node17648;
	wire [4-1:0] node17651;
	wire [4-1:0] node17652;
	wire [4-1:0] node17653;
	wire [4-1:0] node17654;
	wire [4-1:0] node17658;
	wire [4-1:0] node17659;
	wire [4-1:0] node17663;
	wire [4-1:0] node17664;
	wire [4-1:0] node17665;
	wire [4-1:0] node17669;
	wire [4-1:0] node17670;
	wire [4-1:0] node17674;
	wire [4-1:0] node17675;
	wire [4-1:0] node17676;
	wire [4-1:0] node17677;
	wire [4-1:0] node17678;
	wire [4-1:0] node17681;
	wire [4-1:0] node17684;
	wire [4-1:0] node17685;
	wire [4-1:0] node17688;
	wire [4-1:0] node17691;
	wire [4-1:0] node17692;
	wire [4-1:0] node17695;
	wire [4-1:0] node17698;
	wire [4-1:0] node17699;
	wire [4-1:0] node17700;
	wire [4-1:0] node17701;
	wire [4-1:0] node17705;
	wire [4-1:0] node17706;
	wire [4-1:0] node17710;
	wire [4-1:0] node17711;
	wire [4-1:0] node17712;
	wire [4-1:0] node17716;
	wire [4-1:0] node17717;
	wire [4-1:0] node17721;
	wire [4-1:0] node17722;
	wire [4-1:0] node17723;
	wire [4-1:0] node17724;
	wire [4-1:0] node17725;
	wire [4-1:0] node17726;
	wire [4-1:0] node17729;
	wire [4-1:0] node17732;
	wire [4-1:0] node17733;
	wire [4-1:0] node17734;
	wire [4-1:0] node17737;
	wire [4-1:0] node17740;
	wire [4-1:0] node17741;
	wire [4-1:0] node17744;
	wire [4-1:0] node17747;
	wire [4-1:0] node17748;
	wire [4-1:0] node17749;
	wire [4-1:0] node17752;
	wire [4-1:0] node17755;
	wire [4-1:0] node17756;
	wire [4-1:0] node17759;
	wire [4-1:0] node17762;
	wire [4-1:0] node17763;
	wire [4-1:0] node17764;
	wire [4-1:0] node17765;
	wire [4-1:0] node17766;
	wire [4-1:0] node17769;
	wire [4-1:0] node17772;
	wire [4-1:0] node17774;
	wire [4-1:0] node17777;
	wire [4-1:0] node17778;
	wire [4-1:0] node17779;
	wire [4-1:0] node17782;
	wire [4-1:0] node17785;
	wire [4-1:0] node17786;
	wire [4-1:0] node17790;
	wire [4-1:0] node17791;
	wire [4-1:0] node17792;
	wire [4-1:0] node17795;
	wire [4-1:0] node17798;
	wire [4-1:0] node17799;
	wire [4-1:0] node17800;
	wire [4-1:0] node17804;
	wire [4-1:0] node17805;
	wire [4-1:0] node17808;
	wire [4-1:0] node17811;
	wire [4-1:0] node17812;
	wire [4-1:0] node17813;
	wire [4-1:0] node17814;
	wire [4-1:0] node17815;
	wire [4-1:0] node17816;
	wire [4-1:0] node17819;
	wire [4-1:0] node17822;
	wire [4-1:0] node17823;
	wire [4-1:0] node17827;
	wire [4-1:0] node17828;
	wire [4-1:0] node17829;
	wire [4-1:0] node17833;
	wire [4-1:0] node17834;
	wire [4-1:0] node17838;
	wire [4-1:0] node17839;
	wire [4-1:0] node17840;
	wire [4-1:0] node17843;
	wire [4-1:0] node17844;
	wire [4-1:0] node17848;
	wire [4-1:0] node17849;
	wire [4-1:0] node17850;
	wire [4-1:0] node17854;
	wire [4-1:0] node17855;
	wire [4-1:0] node17859;
	wire [4-1:0] node17860;
	wire [4-1:0] node17861;
	wire [4-1:0] node17862;
	wire [4-1:0] node17865;
	wire [4-1:0] node17867;
	wire [4-1:0] node17870;
	wire [4-1:0] node17871;
	wire [4-1:0] node17873;
	wire [4-1:0] node17876;
	wire [4-1:0] node17879;
	wire [4-1:0] node17880;
	wire [4-1:0] node17881;
	wire [4-1:0] node17882;
	wire [4-1:0] node17886;
	wire [4-1:0] node17887;
	wire [4-1:0] node17891;
	wire [4-1:0] node17892;
	wire [4-1:0] node17893;
	wire [4-1:0] node17897;
	wire [4-1:0] node17898;
	wire [4-1:0] node17902;
	wire [4-1:0] node17903;
	wire [4-1:0] node17904;
	wire [4-1:0] node17905;
	wire [4-1:0] node17906;
	wire [4-1:0] node17907;
	wire [4-1:0] node17908;
	wire [4-1:0] node17909;
	wire [4-1:0] node17912;
	wire [4-1:0] node17915;
	wire [4-1:0] node17916;
	wire [4-1:0] node17919;
	wire [4-1:0] node17922;
	wire [4-1:0] node17923;
	wire [4-1:0] node17925;
	wire [4-1:0] node17928;
	wire [4-1:0] node17929;
	wire [4-1:0] node17932;
	wire [4-1:0] node17935;
	wire [4-1:0] node17936;
	wire [4-1:0] node17939;
	wire [4-1:0] node17942;
	wire [4-1:0] node17943;
	wire [4-1:0] node17944;
	wire [4-1:0] node17945;
	wire [4-1:0] node17946;
	wire [4-1:0] node17949;
	wire [4-1:0] node17952;
	wire [4-1:0] node17953;
	wire [4-1:0] node17956;
	wire [4-1:0] node17959;
	wire [4-1:0] node17960;
	wire [4-1:0] node17963;
	wire [4-1:0] node17966;
	wire [4-1:0] node17967;
	wire [4-1:0] node17970;
	wire [4-1:0] node17973;
	wire [4-1:0] node17974;
	wire [4-1:0] node17975;
	wire [4-1:0] node17976;
	wire [4-1:0] node17977;
	wire [4-1:0] node17979;
	wire [4-1:0] node17983;
	wire [4-1:0] node17984;
	wire [4-1:0] node17987;
	wire [4-1:0] node17990;
	wire [4-1:0] node17991;
	wire [4-1:0] node17992;
	wire [4-1:0] node17993;
	wire [4-1:0] node17996;
	wire [4-1:0] node17999;
	wire [4-1:0] node18000;
	wire [4-1:0] node18003;
	wire [4-1:0] node18006;
	wire [4-1:0] node18007;
	wire [4-1:0] node18010;
	wire [4-1:0] node18013;
	wire [4-1:0] node18014;
	wire [4-1:0] node18015;
	wire [4-1:0] node18016;
	wire [4-1:0] node18020;
	wire [4-1:0] node18021;
	wire [4-1:0] node18025;
	wire [4-1:0] node18026;
	wire [4-1:0] node18027;
	wire [4-1:0] node18031;
	wire [4-1:0] node18032;
	wire [4-1:0] node18036;
	wire [4-1:0] node18037;
	wire [4-1:0] node18038;
	wire [4-1:0] node18039;
	wire [4-1:0] node18040;
	wire [4-1:0] node18041;
	wire [4-1:0] node18044;
	wire [4-1:0] node18047;
	wire [4-1:0] node18048;
	wire [4-1:0] node18051;
	wire [4-1:0] node18055;
	wire [4-1:0] node18056;
	wire [4-1:0] node18057;
	wire [4-1:0] node18060;
	wire [4-1:0] node18064;
	wire [4-1:0] node18065;
	wire [4-1:0] node18066;
	wire [4-1:0] node18067;
	wire [4-1:0] node18069;
	wire [4-1:0] node18072;
	wire [4-1:0] node18073;
	wire [4-1:0] node18076;
	wire [4-1:0] node18080;
	wire [4-1:0] node18081;
	wire [4-1:0] node18082;
	wire [4-1:0] node18083;
	wire [4-1:0] node18086;
	wire [4-1:0] node18089;
	wire [4-1:0] node18090;
	wire [4-1:0] node18091;
	wire [4-1:0] node18094;
	wire [4-1:0] node18097;
	wire [4-1:0] node18099;
	wire [4-1:0] node18103;
	wire [4-1:0] node18104;
	wire [4-1:0] node18105;
	wire [4-1:0] node18106;
	wire [4-1:0] node18107;
	wire [4-1:0] node18108;
	wire [4-1:0] node18109;
	wire [4-1:0] node18110;
	wire [4-1:0] node18111;
	wire [4-1:0] node18112;
	wire [4-1:0] node18115;
	wire [4-1:0] node18116;
	wire [4-1:0] node18118;
	wire [4-1:0] node18119;
	wire [4-1:0] node18122;
	wire [4-1:0] node18125;
	wire [4-1:0] node18126;
	wire [4-1:0] node18128;
	wire [4-1:0] node18132;
	wire [4-1:0] node18133;
	wire [4-1:0] node18136;
	wire [4-1:0] node18137;
	wire [4-1:0] node18139;
	wire [4-1:0] node18140;
	wire [4-1:0] node18144;
	wire [4-1:0] node18145;
	wire [4-1:0] node18146;
	wire [4-1:0] node18149;
	wire [4-1:0] node18153;
	wire [4-1:0] node18154;
	wire [4-1:0] node18155;
	wire [4-1:0] node18156;
	wire [4-1:0] node18158;
	wire [4-1:0] node18161;
	wire [4-1:0] node18163;
	wire [4-1:0] node18166;
	wire [4-1:0] node18167;
	wire [4-1:0] node18168;
	wire [4-1:0] node18169;
	wire [4-1:0] node18171;
	wire [4-1:0] node18175;
	wire [4-1:0] node18176;
	wire [4-1:0] node18179;
	wire [4-1:0] node18182;
	wire [4-1:0] node18183;
	wire [4-1:0] node18184;
	wire [4-1:0] node18188;
	wire [4-1:0] node18190;
	wire [4-1:0] node18193;
	wire [4-1:0] node18194;
	wire [4-1:0] node18195;
	wire [4-1:0] node18196;
	wire [4-1:0] node18200;
	wire [4-1:0] node18201;
	wire [4-1:0] node18205;
	wire [4-1:0] node18206;
	wire [4-1:0] node18207;
	wire [4-1:0] node18208;
	wire [4-1:0] node18212;
	wire [4-1:0] node18214;
	wire [4-1:0] node18217;
	wire [4-1:0] node18218;
	wire [4-1:0] node18219;
	wire [4-1:0] node18222;
	wire [4-1:0] node18225;
	wire [4-1:0] node18226;
	wire [4-1:0] node18230;
	wire [4-1:0] node18231;
	wire [4-1:0] node18232;
	wire [4-1:0] node18233;
	wire [4-1:0] node18234;
	wire [4-1:0] node18235;
	wire [4-1:0] node18236;
	wire [4-1:0] node18239;
	wire [4-1:0] node18242;
	wire [4-1:0] node18243;
	wire [4-1:0] node18246;
	wire [4-1:0] node18249;
	wire [4-1:0] node18250;
	wire [4-1:0] node18251;
	wire [4-1:0] node18254;
	wire [4-1:0] node18257;
	wire [4-1:0] node18258;
	wire [4-1:0] node18261;
	wire [4-1:0] node18264;
	wire [4-1:0] node18265;
	wire [4-1:0] node18266;
	wire [4-1:0] node18268;
	wire [4-1:0] node18271;
	wire [4-1:0] node18273;
	wire [4-1:0] node18276;
	wire [4-1:0] node18277;
	wire [4-1:0] node18278;
	wire [4-1:0] node18282;
	wire [4-1:0] node18284;
	wire [4-1:0] node18287;
	wire [4-1:0] node18288;
	wire [4-1:0] node18289;
	wire [4-1:0] node18290;
	wire [4-1:0] node18291;
	wire [4-1:0] node18294;
	wire [4-1:0] node18297;
	wire [4-1:0] node18298;
	wire [4-1:0] node18302;
	wire [4-1:0] node18303;
	wire [4-1:0] node18304;
	wire [4-1:0] node18307;
	wire [4-1:0] node18310;
	wire [4-1:0] node18312;
	wire [4-1:0] node18315;
	wire [4-1:0] node18316;
	wire [4-1:0] node18317;
	wire [4-1:0] node18320;
	wire [4-1:0] node18323;
	wire [4-1:0] node18324;
	wire [4-1:0] node18325;
	wire [4-1:0] node18328;
	wire [4-1:0] node18331;
	wire [4-1:0] node18332;
	wire [4-1:0] node18336;
	wire [4-1:0] node18337;
	wire [4-1:0] node18338;
	wire [4-1:0] node18339;
	wire [4-1:0] node18340;
	wire [4-1:0] node18341;
	wire [4-1:0] node18344;
	wire [4-1:0] node18347;
	wire [4-1:0] node18349;
	wire [4-1:0] node18352;
	wire [4-1:0] node18353;
	wire [4-1:0] node18354;
	wire [4-1:0] node18357;
	wire [4-1:0] node18360;
	wire [4-1:0] node18362;
	wire [4-1:0] node18365;
	wire [4-1:0] node18366;
	wire [4-1:0] node18367;
	wire [4-1:0] node18368;
	wire [4-1:0] node18372;
	wire [4-1:0] node18373;
	wire [4-1:0] node18376;
	wire [4-1:0] node18379;
	wire [4-1:0] node18380;
	wire [4-1:0] node18383;
	wire [4-1:0] node18386;
	wire [4-1:0] node18387;
	wire [4-1:0] node18388;
	wire [4-1:0] node18389;
	wire [4-1:0] node18390;
	wire [4-1:0] node18393;
	wire [4-1:0] node18396;
	wire [4-1:0] node18397;
	wire [4-1:0] node18400;
	wire [4-1:0] node18403;
	wire [4-1:0] node18404;
	wire [4-1:0] node18405;
	wire [4-1:0] node18408;
	wire [4-1:0] node18411;
	wire [4-1:0] node18412;
	wire [4-1:0] node18415;
	wire [4-1:0] node18418;
	wire [4-1:0] node18419;
	wire [4-1:0] node18420;
	wire [4-1:0] node18422;
	wire [4-1:0] node18425;
	wire [4-1:0] node18426;
	wire [4-1:0] node18430;
	wire [4-1:0] node18431;
	wire [4-1:0] node18433;
	wire [4-1:0] node18436;
	wire [4-1:0] node18438;
	wire [4-1:0] node18441;
	wire [4-1:0] node18442;
	wire [4-1:0] node18443;
	wire [4-1:0] node18444;
	wire [4-1:0] node18445;
	wire [4-1:0] node18446;
	wire [4-1:0] node18447;
	wire [4-1:0] node18448;
	wire [4-1:0] node18451;
	wire [4-1:0] node18454;
	wire [4-1:0] node18455;
	wire [4-1:0] node18458;
	wire [4-1:0] node18461;
	wire [4-1:0] node18462;
	wire [4-1:0] node18465;
	wire [4-1:0] node18467;
	wire [4-1:0] node18470;
	wire [4-1:0] node18471;
	wire [4-1:0] node18472;
	wire [4-1:0] node18473;
	wire [4-1:0] node18476;
	wire [4-1:0] node18479;
	wire [4-1:0] node18480;
	wire [4-1:0] node18484;
	wire [4-1:0] node18485;
	wire [4-1:0] node18488;
	wire [4-1:0] node18490;
	wire [4-1:0] node18493;
	wire [4-1:0] node18494;
	wire [4-1:0] node18495;
	wire [4-1:0] node18496;
	wire [4-1:0] node18497;
	wire [4-1:0] node18498;
	wire [4-1:0] node18501;
	wire [4-1:0] node18504;
	wire [4-1:0] node18505;
	wire [4-1:0] node18508;
	wire [4-1:0] node18511;
	wire [4-1:0] node18512;
	wire [4-1:0] node18515;
	wire [4-1:0] node18518;
	wire [4-1:0] node18519;
	wire [4-1:0] node18520;
	wire [4-1:0] node18523;
	wire [4-1:0] node18526;
	wire [4-1:0] node18527;
	wire [4-1:0] node18530;
	wire [4-1:0] node18533;
	wire [4-1:0] node18534;
	wire [4-1:0] node18535;
	wire [4-1:0] node18536;
	wire [4-1:0] node18539;
	wire [4-1:0] node18542;
	wire [4-1:0] node18543;
	wire [4-1:0] node18546;
	wire [4-1:0] node18549;
	wire [4-1:0] node18550;
	wire [4-1:0] node18551;
	wire [4-1:0] node18554;
	wire [4-1:0] node18557;
	wire [4-1:0] node18558;
	wire [4-1:0] node18559;
	wire [4-1:0] node18562;
	wire [4-1:0] node18565;
	wire [4-1:0] node18566;
	wire [4-1:0] node18570;
	wire [4-1:0] node18571;
	wire [4-1:0] node18572;
	wire [4-1:0] node18573;
	wire [4-1:0] node18574;
	wire [4-1:0] node18575;
	wire [4-1:0] node18578;
	wire [4-1:0] node18581;
	wire [4-1:0] node18582;
	wire [4-1:0] node18585;
	wire [4-1:0] node18588;
	wire [4-1:0] node18589;
	wire [4-1:0] node18590;
	wire [4-1:0] node18593;
	wire [4-1:0] node18596;
	wire [4-1:0] node18597;
	wire [4-1:0] node18600;
	wire [4-1:0] node18603;
	wire [4-1:0] node18604;
	wire [4-1:0] node18605;
	wire [4-1:0] node18606;
	wire [4-1:0] node18609;
	wire [4-1:0] node18612;
	wire [4-1:0] node18613;
	wire [4-1:0] node18616;
	wire [4-1:0] node18619;
	wire [4-1:0] node18620;
	wire [4-1:0] node18621;
	wire [4-1:0] node18622;
	wire [4-1:0] node18625;
	wire [4-1:0] node18628;
	wire [4-1:0] node18629;
	wire [4-1:0] node18632;
	wire [4-1:0] node18635;
	wire [4-1:0] node18636;
	wire [4-1:0] node18639;
	wire [4-1:0] node18642;
	wire [4-1:0] node18643;
	wire [4-1:0] node18644;
	wire [4-1:0] node18645;
	wire [4-1:0] node18646;
	wire [4-1:0] node18649;
	wire [4-1:0] node18652;
	wire [4-1:0] node18653;
	wire [4-1:0] node18656;
	wire [4-1:0] node18659;
	wire [4-1:0] node18660;
	wire [4-1:0] node18661;
	wire [4-1:0] node18664;
	wire [4-1:0] node18667;
	wire [4-1:0] node18668;
	wire [4-1:0] node18671;
	wire [4-1:0] node18674;
	wire [4-1:0] node18675;
	wire [4-1:0] node18676;
	wire [4-1:0] node18677;
	wire [4-1:0] node18681;
	wire [4-1:0] node18684;
	wire [4-1:0] node18685;
	wire [4-1:0] node18686;
	wire [4-1:0] node18690;
	wire [4-1:0] node18693;
	wire [4-1:0] node18694;
	wire [4-1:0] node18695;
	wire [4-1:0] node18696;
	wire [4-1:0] node18697;
	wire [4-1:0] node18698;
	wire [4-1:0] node18699;
	wire [4-1:0] node18702;
	wire [4-1:0] node18705;
	wire [4-1:0] node18706;
	wire [4-1:0] node18710;
	wire [4-1:0] node18711;
	wire [4-1:0] node18714;
	wire [4-1:0] node18716;
	wire [4-1:0] node18719;
	wire [4-1:0] node18720;
	wire [4-1:0] node18721;
	wire [4-1:0] node18722;
	wire [4-1:0] node18726;
	wire [4-1:0] node18728;
	wire [4-1:0] node18731;
	wire [4-1:0] node18732;
	wire [4-1:0] node18734;
	wire [4-1:0] node18737;
	wire [4-1:0] node18738;
	wire [4-1:0] node18741;
	wire [4-1:0] node18744;
	wire [4-1:0] node18745;
	wire [4-1:0] node18746;
	wire [4-1:0] node18747;
	wire [4-1:0] node18748;
	wire [4-1:0] node18751;
	wire [4-1:0] node18754;
	wire [4-1:0] node18755;
	wire [4-1:0] node18756;
	wire [4-1:0] node18759;
	wire [4-1:0] node18762;
	wire [4-1:0] node18763;
	wire [4-1:0] node18766;
	wire [4-1:0] node18769;
	wire [4-1:0] node18770;
	wire [4-1:0] node18772;
	wire [4-1:0] node18775;
	wire [4-1:0] node18776;
	wire [4-1:0] node18779;
	wire [4-1:0] node18782;
	wire [4-1:0] node18783;
	wire [4-1:0] node18784;
	wire [4-1:0] node18785;
	wire [4-1:0] node18789;
	wire [4-1:0] node18790;
	wire [4-1:0] node18793;
	wire [4-1:0] node18796;
	wire [4-1:0] node18797;
	wire [4-1:0] node18799;
	wire [4-1:0] node18802;
	wire [4-1:0] node18804;
	wire [4-1:0] node18807;
	wire [4-1:0] node18808;
	wire [4-1:0] node18809;
	wire [4-1:0] node18810;
	wire [4-1:0] node18811;
	wire [4-1:0] node18812;
	wire [4-1:0] node18815;
	wire [4-1:0] node18818;
	wire [4-1:0] node18819;
	wire [4-1:0] node18822;
	wire [4-1:0] node18825;
	wire [4-1:0] node18826;
	wire [4-1:0] node18828;
	wire [4-1:0] node18831;
	wire [4-1:0] node18832;
	wire [4-1:0] node18836;
	wire [4-1:0] node18837;
	wire [4-1:0] node18838;
	wire [4-1:0] node18839;
	wire [4-1:0] node18842;
	wire [4-1:0] node18845;
	wire [4-1:0] node18846;
	wire [4-1:0] node18849;
	wire [4-1:0] node18852;
	wire [4-1:0] node18853;
	wire [4-1:0] node18854;
	wire [4-1:0] node18857;
	wire [4-1:0] node18860;
	wire [4-1:0] node18861;
	wire [4-1:0] node18864;
	wire [4-1:0] node18867;
	wire [4-1:0] node18868;
	wire [4-1:0] node18869;
	wire [4-1:0] node18870;
	wire [4-1:0] node18871;
	wire [4-1:0] node18874;
	wire [4-1:0] node18877;
	wire [4-1:0] node18878;
	wire [4-1:0] node18881;
	wire [4-1:0] node18884;
	wire [4-1:0] node18885;
	wire [4-1:0] node18886;
	wire [4-1:0] node18889;
	wire [4-1:0] node18892;
	wire [4-1:0] node18893;
	wire [4-1:0] node18896;
	wire [4-1:0] node18899;
	wire [4-1:0] node18900;
	wire [4-1:0] node18901;
	wire [4-1:0] node18902;
	wire [4-1:0] node18905;
	wire [4-1:0] node18908;
	wire [4-1:0] node18909;
	wire [4-1:0] node18912;
	wire [4-1:0] node18915;
	wire [4-1:0] node18916;
	wire [4-1:0] node18917;
	wire [4-1:0] node18921;
	wire [4-1:0] node18923;
	wire [4-1:0] node18926;
	wire [4-1:0] node18927;
	wire [4-1:0] node18928;
	wire [4-1:0] node18929;
	wire [4-1:0] node18930;
	wire [4-1:0] node18931;
	wire [4-1:0] node18934;
	wire [4-1:0] node18935;
	wire [4-1:0] node18937;
	wire [4-1:0] node18938;
	wire [4-1:0] node18941;
	wire [4-1:0] node18944;
	wire [4-1:0] node18945;
	wire [4-1:0] node18947;
	wire [4-1:0] node18951;
	wire [4-1:0] node18952;
	wire [4-1:0] node18955;
	wire [4-1:0] node18956;
	wire [4-1:0] node18958;
	wire [4-1:0] node18959;
	wire [4-1:0] node18963;
	wire [4-1:0] node18964;
	wire [4-1:0] node18965;
	wire [4-1:0] node18968;
	wire [4-1:0] node18972;
	wire [4-1:0] node18973;
	wire [4-1:0] node18974;
	wire [4-1:0] node18975;
	wire [4-1:0] node18977;
	wire [4-1:0] node18980;
	wire [4-1:0] node18982;
	wire [4-1:0] node18985;
	wire [4-1:0] node18986;
	wire [4-1:0] node18987;
	wire [4-1:0] node18989;
	wire [4-1:0] node18992;
	wire [4-1:0] node18993;
	wire [4-1:0] node18996;
	wire [4-1:0] node18999;
	wire [4-1:0] node19000;
	wire [4-1:0] node19001;
	wire [4-1:0] node19005;
	wire [4-1:0] node19007;
	wire [4-1:0] node19010;
	wire [4-1:0] node19011;
	wire [4-1:0] node19012;
	wire [4-1:0] node19013;
	wire [4-1:0] node19017;
	wire [4-1:0] node19018;
	wire [4-1:0] node19022;
	wire [4-1:0] node19023;
	wire [4-1:0] node19024;
	wire [4-1:0] node19025;
	wire [4-1:0] node19029;
	wire [4-1:0] node19031;
	wire [4-1:0] node19034;
	wire [4-1:0] node19035;
	wire [4-1:0] node19036;
	wire [4-1:0] node19039;
	wire [4-1:0] node19042;
	wire [4-1:0] node19043;
	wire [4-1:0] node19047;
	wire [4-1:0] node19048;
	wire [4-1:0] node19049;
	wire [4-1:0] node19050;
	wire [4-1:0] node19051;
	wire [4-1:0] node19052;
	wire [4-1:0] node19055;
	wire [4-1:0] node19058;
	wire [4-1:0] node19059;
	wire [4-1:0] node19060;
	wire [4-1:0] node19063;
	wire [4-1:0] node19066;
	wire [4-1:0] node19067;
	wire [4-1:0] node19070;
	wire [4-1:0] node19073;
	wire [4-1:0] node19074;
	wire [4-1:0] node19075;
	wire [4-1:0] node19078;
	wire [4-1:0] node19081;
	wire [4-1:0] node19082;
	wire [4-1:0] node19085;
	wire [4-1:0] node19088;
	wire [4-1:0] node19089;
	wire [4-1:0] node19090;
	wire [4-1:0] node19091;
	wire [4-1:0] node19094;
	wire [4-1:0] node19097;
	wire [4-1:0] node19098;
	wire [4-1:0] node19102;
	wire [4-1:0] node19103;
	wire [4-1:0] node19104;
	wire [4-1:0] node19107;
	wire [4-1:0] node19110;
	wire [4-1:0] node19111;
	wire [4-1:0] node19114;
	wire [4-1:0] node19117;
	wire [4-1:0] node19118;
	wire [4-1:0] node19119;
	wire [4-1:0] node19120;
	wire [4-1:0] node19121;
	wire [4-1:0] node19122;
	wire [4-1:0] node19126;
	wire [4-1:0] node19127;
	wire [4-1:0] node19131;
	wire [4-1:0] node19132;
	wire [4-1:0] node19135;
	wire [4-1:0] node19138;
	wire [4-1:0] node19139;
	wire [4-1:0] node19141;
	wire [4-1:0] node19142;
	wire [4-1:0] node19145;
	wire [4-1:0] node19148;
	wire [4-1:0] node19149;
	wire [4-1:0] node19150;
	wire [4-1:0] node19154;
	wire [4-1:0] node19155;
	wire [4-1:0] node19159;
	wire [4-1:0] node19160;
	wire [4-1:0] node19161;
	wire [4-1:0] node19162;
	wire [4-1:0] node19163;
	wire [4-1:0] node19167;
	wire [4-1:0] node19168;
	wire [4-1:0] node19169;
	wire [4-1:0] node19172;
	wire [4-1:0] node19175;
	wire [4-1:0] node19176;
	wire [4-1:0] node19179;
	wire [4-1:0] node19182;
	wire [4-1:0] node19183;
	wire [4-1:0] node19186;
	wire [4-1:0] node19187;
	wire [4-1:0] node19191;
	wire [4-1:0] node19192;
	wire [4-1:0] node19193;
	wire [4-1:0] node19195;
	wire [4-1:0] node19198;
	wire [4-1:0] node19200;
	wire [4-1:0] node19203;
	wire [4-1:0] node19204;
	wire [4-1:0] node19207;
	wire [4-1:0] node19209;
	wire [4-1:0] node19212;
	wire [4-1:0] node19213;
	wire [4-1:0] node19214;
	wire [4-1:0] node19215;
	wire [4-1:0] node19216;
	wire [4-1:0] node19217;
	wire [4-1:0] node19218;
	wire [4-1:0] node19220;
	wire [4-1:0] node19223;
	wire [4-1:0] node19224;
	wire [4-1:0] node19228;
	wire [4-1:0] node19230;
	wire [4-1:0] node19232;
	wire [4-1:0] node19235;
	wire [4-1:0] node19236;
	wire [4-1:0] node19237;
	wire [4-1:0] node19238;
	wire [4-1:0] node19242;
	wire [4-1:0] node19244;
	wire [4-1:0] node19247;
	wire [4-1:0] node19248;
	wire [4-1:0] node19249;
	wire [4-1:0] node19253;
	wire [4-1:0] node19255;
	wire [4-1:0] node19258;
	wire [4-1:0] node19259;
	wire [4-1:0] node19260;
	wire [4-1:0] node19262;
	wire [4-1:0] node19263;
	wire [4-1:0] node19264;
	wire [4-1:0] node19267;
	wire [4-1:0] node19270;
	wire [4-1:0] node19271;
	wire [4-1:0] node19274;
	wire [4-1:0] node19277;
	wire [4-1:0] node19278;
	wire [4-1:0] node19279;
	wire [4-1:0] node19283;
	wire [4-1:0] node19285;
	wire [4-1:0] node19288;
	wire [4-1:0] node19289;
	wire [4-1:0] node19290;
	wire [4-1:0] node19292;
	wire [4-1:0] node19295;
	wire [4-1:0] node19296;
	wire [4-1:0] node19300;
	wire [4-1:0] node19301;
	wire [4-1:0] node19302;
	wire [4-1:0] node19305;
	wire [4-1:0] node19309;
	wire [4-1:0] node19310;
	wire [4-1:0] node19311;
	wire [4-1:0] node19312;
	wire [4-1:0] node19313;
	wire [4-1:0] node19315;
	wire [4-1:0] node19318;
	wire [4-1:0] node19319;
	wire [4-1:0] node19323;
	wire [4-1:0] node19324;
	wire [4-1:0] node19325;
	wire [4-1:0] node19329;
	wire [4-1:0] node19330;
	wire [4-1:0] node19334;
	wire [4-1:0] node19335;
	wire [4-1:0] node19336;
	wire [4-1:0] node19337;
	wire [4-1:0] node19341;
	wire [4-1:0] node19343;
	wire [4-1:0] node19346;
	wire [4-1:0] node19347;
	wire [4-1:0] node19349;
	wire [4-1:0] node19352;
	wire [4-1:0] node19354;
	wire [4-1:0] node19357;
	wire [4-1:0] node19358;
	wire [4-1:0] node19359;
	wire [4-1:0] node19361;
	wire [4-1:0] node19362;
	wire [4-1:0] node19363;
	wire [4-1:0] node19366;
	wire [4-1:0] node19369;
	wire [4-1:0] node19370;
	wire [4-1:0] node19374;
	wire [4-1:0] node19375;
	wire [4-1:0] node19377;
	wire [4-1:0] node19380;
	wire [4-1:0] node19382;
	wire [4-1:0] node19385;
	wire [4-1:0] node19386;
	wire [4-1:0] node19388;
	wire [4-1:0] node19390;
	wire [4-1:0] node19393;
	wire [4-1:0] node19394;
	wire [4-1:0] node19395;
	wire [4-1:0] node19399;
	wire [4-1:0] node19401;
	wire [4-1:0] node19404;
	wire [4-1:0] node19405;
	wire [4-1:0] node19406;
	wire [4-1:0] node19407;
	wire [4-1:0] node19408;
	wire [4-1:0] node19409;
	wire [4-1:0] node19411;
	wire [4-1:0] node19414;
	wire [4-1:0] node19415;
	wire [4-1:0] node19419;
	wire [4-1:0] node19420;
	wire [4-1:0] node19421;
	wire [4-1:0] node19425;
	wire [4-1:0] node19427;
	wire [4-1:0] node19430;
	wire [4-1:0] node19431;
	wire [4-1:0] node19432;
	wire [4-1:0] node19433;
	wire [4-1:0] node19437;
	wire [4-1:0] node19439;
	wire [4-1:0] node19442;
	wire [4-1:0] node19443;
	wire [4-1:0] node19446;
	wire [4-1:0] node19447;
	wire [4-1:0] node19451;
	wire [4-1:0] node19452;
	wire [4-1:0] node19453;
	wire [4-1:0] node19454;
	wire [4-1:0] node19457;
	wire [4-1:0] node19458;
	wire [4-1:0] node19462;
	wire [4-1:0] node19463;
	wire [4-1:0] node19464;
	wire [4-1:0] node19467;
	wire [4-1:0] node19470;
	wire [4-1:0] node19472;
	wire [4-1:0] node19475;
	wire [4-1:0] node19476;
	wire [4-1:0] node19477;
	wire [4-1:0] node19479;
	wire [4-1:0] node19482;
	wire [4-1:0] node19483;
	wire [4-1:0] node19487;
	wire [4-1:0] node19488;
	wire [4-1:0] node19489;
	wire [4-1:0] node19493;
	wire [4-1:0] node19494;
	wire [4-1:0] node19498;
	wire [4-1:0] node19499;
	wire [4-1:0] node19500;
	wire [4-1:0] node19501;
	wire [4-1:0] node19502;
	wire [4-1:0] node19503;
	wire [4-1:0] node19507;
	wire [4-1:0] node19510;
	wire [4-1:0] node19511;
	wire [4-1:0] node19513;
	wire [4-1:0] node19516;
	wire [4-1:0] node19517;
	wire [4-1:0] node19521;
	wire [4-1:0] node19522;
	wire [4-1:0] node19523;
	wire [4-1:0] node19524;
	wire [4-1:0] node19528;
	wire [4-1:0] node19530;
	wire [4-1:0] node19533;
	wire [4-1:0] node19534;
	wire [4-1:0] node19536;
	wire [4-1:0] node19540;
	wire [4-1:0] node19541;
	wire [4-1:0] node19542;
	wire [4-1:0] node19543;
	wire [4-1:0] node19544;
	wire [4-1:0] node19548;
	wire [4-1:0] node19549;
	wire [4-1:0] node19553;
	wire [4-1:0] node19554;
	wire [4-1:0] node19555;
	wire [4-1:0] node19559;
	wire [4-1:0] node19561;
	wire [4-1:0] node19564;
	wire [4-1:0] node19565;
	wire [4-1:0] node19566;
	wire [4-1:0] node19567;
	wire [4-1:0] node19571;
	wire [4-1:0] node19572;
	wire [4-1:0] node19575;
	wire [4-1:0] node19578;
	wire [4-1:0] node19579;
	wire [4-1:0] node19580;
	wire [4-1:0] node19583;
	wire [4-1:0] node19586;
	wire [4-1:0] node19587;
	wire [4-1:0] node19590;
	wire [4-1:0] node19593;
	wire [4-1:0] node19594;
	wire [4-1:0] node19595;
	wire [4-1:0] node19596;
	wire [4-1:0] node19597;
	wire [4-1:0] node19598;
	wire [4-1:0] node19599;
	wire [4-1:0] node19602;
	wire [4-1:0] node19603;
	wire [4-1:0] node19605;
	wire [4-1:0] node19606;
	wire [4-1:0] node19609;
	wire [4-1:0] node19612;
	wire [4-1:0] node19613;
	wire [4-1:0] node19615;
	wire [4-1:0] node19619;
	wire [4-1:0] node19620;
	wire [4-1:0] node19623;
	wire [4-1:0] node19624;
	wire [4-1:0] node19626;
	wire [4-1:0] node19627;
	wire [4-1:0] node19631;
	wire [4-1:0] node19632;
	wire [4-1:0] node19633;
	wire [4-1:0] node19638;
	wire [4-1:0] node19639;
	wire [4-1:0] node19640;
	wire [4-1:0] node19641;
	wire [4-1:0] node19643;
	wire [4-1:0] node19646;
	wire [4-1:0] node19648;
	wire [4-1:0] node19651;
	wire [4-1:0] node19652;
	wire [4-1:0] node19653;
	wire [4-1:0] node19655;
	wire [4-1:0] node19658;
	wire [4-1:0] node19659;
	wire [4-1:0] node19662;
	wire [4-1:0] node19665;
	wire [4-1:0] node19666;
	wire [4-1:0] node19667;
	wire [4-1:0] node19671;
	wire [4-1:0] node19673;
	wire [4-1:0] node19676;
	wire [4-1:0] node19677;
	wire [4-1:0] node19678;
	wire [4-1:0] node19679;
	wire [4-1:0] node19683;
	wire [4-1:0] node19684;
	wire [4-1:0] node19688;
	wire [4-1:0] node19689;
	wire [4-1:0] node19690;
	wire [4-1:0] node19691;
	wire [4-1:0] node19695;
	wire [4-1:0] node19698;
	wire [4-1:0] node19699;
	wire [4-1:0] node19700;
	wire [4-1:0] node19703;
	wire [4-1:0] node19706;
	wire [4-1:0] node19707;
	wire [4-1:0] node19711;
	wire [4-1:0] node19712;
	wire [4-1:0] node19713;
	wire [4-1:0] node19714;
	wire [4-1:0] node19715;
	wire [4-1:0] node19716;
	wire [4-1:0] node19719;
	wire [4-1:0] node19721;
	wire [4-1:0] node19724;
	wire [4-1:0] node19725;
	wire [4-1:0] node19726;
	wire [4-1:0] node19727;
	wire [4-1:0] node19731;
	wire [4-1:0] node19732;
	wire [4-1:0] node19735;
	wire [4-1:0] node19738;
	wire [4-1:0] node19739;
	wire [4-1:0] node19742;
	wire [4-1:0] node19745;
	wire [4-1:0] node19746;
	wire [4-1:0] node19747;
	wire [4-1:0] node19749;
	wire [4-1:0] node19752;
	wire [4-1:0] node19755;
	wire [4-1:0] node19756;
	wire [4-1:0] node19757;
	wire [4-1:0] node19758;
	wire [4-1:0] node19761;
	wire [4-1:0] node19764;
	wire [4-1:0] node19765;
	wire [4-1:0] node19768;
	wire [4-1:0] node19771;
	wire [4-1:0] node19772;
	wire [4-1:0] node19775;
	wire [4-1:0] node19778;
	wire [4-1:0] node19779;
	wire [4-1:0] node19780;
	wire [4-1:0] node19781;
	wire [4-1:0] node19782;
	wire [4-1:0] node19785;
	wire [4-1:0] node19788;
	wire [4-1:0] node19789;
	wire [4-1:0] node19793;
	wire [4-1:0] node19794;
	wire [4-1:0] node19795;
	wire [4-1:0] node19799;
	wire [4-1:0] node19802;
	wire [4-1:0] node19803;
	wire [4-1:0] node19804;
	wire [4-1:0] node19805;
	wire [4-1:0] node19808;
	wire [4-1:0] node19811;
	wire [4-1:0] node19812;
	wire [4-1:0] node19816;
	wire [4-1:0] node19817;
	wire [4-1:0] node19818;
	wire [4-1:0] node19821;
	wire [4-1:0] node19824;
	wire [4-1:0] node19825;
	wire [4-1:0] node19828;
	wire [4-1:0] node19831;
	wire [4-1:0] node19832;
	wire [4-1:0] node19833;
	wire [4-1:0] node19834;
	wire [4-1:0] node19835;
	wire [4-1:0] node19837;
	wire [4-1:0] node19840;
	wire [4-1:0] node19842;
	wire [4-1:0] node19845;
	wire [4-1:0] node19846;
	wire [4-1:0] node19849;
	wire [4-1:0] node19850;
	wire [4-1:0] node19854;
	wire [4-1:0] node19855;
	wire [4-1:0] node19856;
	wire [4-1:0] node19858;
	wire [4-1:0] node19861;
	wire [4-1:0] node19864;
	wire [4-1:0] node19865;
	wire [4-1:0] node19866;
	wire [4-1:0] node19870;
	wire [4-1:0] node19871;
	wire [4-1:0] node19875;
	wire [4-1:0] node19876;
	wire [4-1:0] node19877;
	wire [4-1:0] node19878;
	wire [4-1:0] node19879;
	wire [4-1:0] node19883;
	wire [4-1:0] node19886;
	wire [4-1:0] node19887;
	wire [4-1:0] node19889;
	wire [4-1:0] node19892;
	wire [4-1:0] node19894;
	wire [4-1:0] node19897;
	wire [4-1:0] node19898;
	wire [4-1:0] node19899;
	wire [4-1:0] node19901;
	wire [4-1:0] node19904;
	wire [4-1:0] node19905;
	wire [4-1:0] node19909;
	wire [4-1:0] node19910;
	wire [4-1:0] node19911;
	wire [4-1:0] node19915;
	wire [4-1:0] node19918;
	wire [4-1:0] node19919;
	wire [4-1:0] node19920;
	wire [4-1:0] node19921;
	wire [4-1:0] node19922;
	wire [4-1:0] node19923;
	wire [4-1:0] node19924;
	wire [4-1:0] node19927;
	wire [4-1:0] node19930;
	wire [4-1:0] node19931;
	wire [4-1:0] node19932;
	wire [4-1:0] node19935;
	wire [4-1:0] node19938;
	wire [4-1:0] node19939;
	wire [4-1:0] node19942;
	wire [4-1:0] node19945;
	wire [4-1:0] node19946;
	wire [4-1:0] node19947;
	wire [4-1:0] node19948;
	wire [4-1:0] node19952;
	wire [4-1:0] node19953;
	wire [4-1:0] node19957;
	wire [4-1:0] node19958;
	wire [4-1:0] node19959;
	wire [4-1:0] node19963;
	wire [4-1:0] node19964;
	wire [4-1:0] node19967;
	wire [4-1:0] node19970;
	wire [4-1:0] node19971;
	wire [4-1:0] node19972;
	wire [4-1:0] node19973;
	wire [4-1:0] node19974;
	wire [4-1:0] node19977;
	wire [4-1:0] node19980;
	wire [4-1:0] node19981;
	wire [4-1:0] node19985;
	wire [4-1:0] node19986;
	wire [4-1:0] node19989;
	wire [4-1:0] node19991;
	wire [4-1:0] node19994;
	wire [4-1:0] node19995;
	wire [4-1:0] node19996;
	wire [4-1:0] node19997;
	wire [4-1:0] node20001;
	wire [4-1:0] node20002;
	wire [4-1:0] node20006;
	wire [4-1:0] node20007;
	wire [4-1:0] node20008;
	wire [4-1:0] node20011;
	wire [4-1:0] node20014;
	wire [4-1:0] node20015;
	wire [4-1:0] node20019;
	wire [4-1:0] node20020;
	wire [4-1:0] node20021;
	wire [4-1:0] node20022;
	wire [4-1:0] node20023;
	wire [4-1:0] node20024;
	wire [4-1:0] node20025;
	wire [4-1:0] node20028;
	wire [4-1:0] node20031;
	wire [4-1:0] node20032;
	wire [4-1:0] node20036;
	wire [4-1:0] node20037;
	wire [4-1:0] node20040;
	wire [4-1:0] node20043;
	wire [4-1:0] node20044;
	wire [4-1:0] node20045;
	wire [4-1:0] node20046;
	wire [4-1:0] node20049;
	wire [4-1:0] node20052;
	wire [4-1:0] node20053;
	wire [4-1:0] node20056;
	wire [4-1:0] node20059;
	wire [4-1:0] node20060;
	wire [4-1:0] node20061;
	wire [4-1:0] node20064;
	wire [4-1:0] node20067;
	wire [4-1:0] node20068;
	wire [4-1:0] node20071;
	wire [4-1:0] node20074;
	wire [4-1:0] node20075;
	wire [4-1:0] node20076;
	wire [4-1:0] node20077;
	wire [4-1:0] node20081;
	wire [4-1:0] node20082;
	wire [4-1:0] node20085;
	wire [4-1:0] node20088;
	wire [4-1:0] node20089;
	wire [4-1:0] node20091;
	wire [4-1:0] node20094;
	wire [4-1:0] node20096;
	wire [4-1:0] node20099;
	wire [4-1:0] node20100;
	wire [4-1:0] node20101;
	wire [4-1:0] node20102;
	wire [4-1:0] node20103;
	wire [4-1:0] node20106;
	wire [4-1:0] node20109;
	wire [4-1:0] node20110;
	wire [4-1:0] node20113;
	wire [4-1:0] node20116;
	wire [4-1:0] node20117;
	wire [4-1:0] node20119;
	wire [4-1:0] node20122;
	wire [4-1:0] node20123;
	wire [4-1:0] node20126;
	wire [4-1:0] node20129;
	wire [4-1:0] node20130;
	wire [4-1:0] node20131;
	wire [4-1:0] node20132;
	wire [4-1:0] node20135;
	wire [4-1:0] node20138;
	wire [4-1:0] node20140;
	wire [4-1:0] node20143;
	wire [4-1:0] node20144;
	wire [4-1:0] node20145;
	wire [4-1:0] node20149;
	wire [4-1:0] node20151;
	wire [4-1:0] node20154;
	wire [4-1:0] node20155;
	wire [4-1:0] node20156;
	wire [4-1:0] node20157;
	wire [4-1:0] node20158;
	wire [4-1:0] node20160;
	wire [4-1:0] node20162;
	wire [4-1:0] node20165;
	wire [4-1:0] node20167;
	wire [4-1:0] node20168;
	wire [4-1:0] node20172;
	wire [4-1:0] node20173;
	wire [4-1:0] node20174;
	wire [4-1:0] node20175;
	wire [4-1:0] node20178;
	wire [4-1:0] node20181;
	wire [4-1:0] node20182;
	wire [4-1:0] node20185;
	wire [4-1:0] node20188;
	wire [4-1:0] node20189;
	wire [4-1:0] node20191;
	wire [4-1:0] node20194;
	wire [4-1:0] node20195;
	wire [4-1:0] node20199;
	wire [4-1:0] node20200;
	wire [4-1:0] node20201;
	wire [4-1:0] node20202;
	wire [4-1:0] node20204;
	wire [4-1:0] node20207;
	wire [4-1:0] node20208;
	wire [4-1:0] node20212;
	wire [4-1:0] node20213;
	wire [4-1:0] node20215;
	wire [4-1:0] node20218;
	wire [4-1:0] node20219;
	wire [4-1:0] node20222;
	wire [4-1:0] node20225;
	wire [4-1:0] node20226;
	wire [4-1:0] node20227;
	wire [4-1:0] node20229;
	wire [4-1:0] node20232;
	wire [4-1:0] node20233;
	wire [4-1:0] node20237;
	wire [4-1:0] node20238;
	wire [4-1:0] node20239;
	wire [4-1:0] node20242;
	wire [4-1:0] node20245;
	wire [4-1:0] node20246;
	wire [4-1:0] node20250;
	wire [4-1:0] node20251;
	wire [4-1:0] node20252;
	wire [4-1:0] node20253;
	wire [4-1:0] node20255;
	wire [4-1:0] node20258;
	wire [4-1:0] node20259;
	wire [4-1:0] node20263;
	wire [4-1:0] node20264;
	wire [4-1:0] node20265;
	wire [4-1:0] node20267;
	wire [4-1:0] node20270;
	wire [4-1:0] node20271;
	wire [4-1:0] node20275;
	wire [4-1:0] node20276;
	wire [4-1:0] node20279;
	wire [4-1:0] node20281;
	wire [4-1:0] node20284;
	wire [4-1:0] node20285;
	wire [4-1:0] node20286;
	wire [4-1:0] node20287;
	wire [4-1:0] node20288;
	wire [4-1:0] node20291;
	wire [4-1:0] node20294;
	wire [4-1:0] node20295;
	wire [4-1:0] node20298;
	wire [4-1:0] node20301;
	wire [4-1:0] node20302;
	wire [4-1:0] node20303;
	wire [4-1:0] node20306;
	wire [4-1:0] node20309;
	wire [4-1:0] node20310;
	wire [4-1:0] node20313;
	wire [4-1:0] node20316;
	wire [4-1:0] node20317;
	wire [4-1:0] node20318;
	wire [4-1:0] node20319;
	wire [4-1:0] node20322;
	wire [4-1:0] node20325;
	wire [4-1:0] node20326;
	wire [4-1:0] node20329;
	wire [4-1:0] node20332;
	wire [4-1:0] node20333;
	wire [4-1:0] node20334;
	wire [4-1:0] node20338;
	wire [4-1:0] node20339;
	wire [4-1:0] node20343;
	wire [4-1:0] node20344;
	wire [4-1:0] node20345;
	wire [4-1:0] node20346;
	wire [4-1:0] node20347;
	wire [4-1:0] node20348;
	wire [4-1:0] node20351;
	wire [4-1:0] node20352;
	wire [4-1:0] node20354;
	wire [4-1:0] node20355;
	wire [4-1:0] node20358;
	wire [4-1:0] node20361;
	wire [4-1:0] node20362;
	wire [4-1:0] node20364;
	wire [4-1:0] node20368;
	wire [4-1:0] node20369;
	wire [4-1:0] node20372;
	wire [4-1:0] node20373;
	wire [4-1:0] node20375;
	wire [4-1:0] node20376;
	wire [4-1:0] node20380;
	wire [4-1:0] node20381;
	wire [4-1:0] node20382;
	wire [4-1:0] node20385;
	wire [4-1:0] node20389;
	wire [4-1:0] node20390;
	wire [4-1:0] node20391;
	wire [4-1:0] node20392;
	wire [4-1:0] node20394;
	wire [4-1:0] node20397;
	wire [4-1:0] node20399;
	wire [4-1:0] node20402;
	wire [4-1:0] node20403;
	wire [4-1:0] node20404;
	wire [4-1:0] node20406;
	wire [4-1:0] node20409;
	wire [4-1:0] node20410;
	wire [4-1:0] node20413;
	wire [4-1:0] node20416;
	wire [4-1:0] node20417;
	wire [4-1:0] node20418;
	wire [4-1:0] node20422;
	wire [4-1:0] node20424;
	wire [4-1:0] node20427;
	wire [4-1:0] node20428;
	wire [4-1:0] node20429;
	wire [4-1:0] node20430;
	wire [4-1:0] node20434;
	wire [4-1:0] node20435;
	wire [4-1:0] node20439;
	wire [4-1:0] node20440;
	wire [4-1:0] node20441;
	wire [4-1:0] node20442;
	wire [4-1:0] node20446;
	wire [4-1:0] node20448;
	wire [4-1:0] node20451;
	wire [4-1:0] node20452;
	wire [4-1:0] node20453;
	wire [4-1:0] node20456;
	wire [4-1:0] node20459;
	wire [4-1:0] node20460;
	wire [4-1:0] node20464;
	wire [4-1:0] node20465;
	wire [4-1:0] node20466;
	wire [4-1:0] node20467;
	wire [4-1:0] node20468;
	wire [4-1:0] node20469;
	wire [4-1:0] node20472;
	wire [4-1:0] node20474;
	wire [4-1:0] node20477;
	wire [4-1:0] node20478;
	wire [4-1:0] node20479;
	wire [4-1:0] node20481;
	wire [4-1:0] node20484;
	wire [4-1:0] node20485;
	wire [4-1:0] node20489;
	wire [4-1:0] node20490;
	wire [4-1:0] node20493;
	wire [4-1:0] node20496;
	wire [4-1:0] node20497;
	wire [4-1:0] node20498;
	wire [4-1:0] node20500;
	wire [4-1:0] node20503;
	wire [4-1:0] node20506;
	wire [4-1:0] node20507;
	wire [4-1:0] node20508;
	wire [4-1:0] node20511;
	wire [4-1:0] node20514;
	wire [4-1:0] node20515;
	wire [4-1:0] node20518;
	wire [4-1:0] node20521;
	wire [4-1:0] node20522;
	wire [4-1:0] node20523;
	wire [4-1:0] node20524;
	wire [4-1:0] node20525;
	wire [4-1:0] node20528;
	wire [4-1:0] node20531;
	wire [4-1:0] node20532;
	wire [4-1:0] node20536;
	wire [4-1:0] node20537;
	wire [4-1:0] node20538;
	wire [4-1:0] node20542;
	wire [4-1:0] node20545;
	wire [4-1:0] node20546;
	wire [4-1:0] node20547;
	wire [4-1:0] node20548;
	wire [4-1:0] node20549;
	wire [4-1:0] node20554;
	wire [4-1:0] node20555;
	wire [4-1:0] node20558;
	wire [4-1:0] node20561;
	wire [4-1:0] node20562;
	wire [4-1:0] node20564;
	wire [4-1:0] node20567;
	wire [4-1:0] node20570;
	wire [4-1:0] node20571;
	wire [4-1:0] node20572;
	wire [4-1:0] node20573;
	wire [4-1:0] node20574;
	wire [4-1:0] node20576;
	wire [4-1:0] node20579;
	wire [4-1:0] node20581;
	wire [4-1:0] node20584;
	wire [4-1:0] node20585;
	wire [4-1:0] node20588;
	wire [4-1:0] node20590;
	wire [4-1:0] node20593;
	wire [4-1:0] node20594;
	wire [4-1:0] node20595;
	wire [4-1:0] node20598;
	wire [4-1:0] node20599;
	wire [4-1:0] node20603;
	wire [4-1:0] node20604;
	wire [4-1:0] node20605;
	wire [4-1:0] node20609;
	wire [4-1:0] node20610;
	wire [4-1:0] node20614;
	wire [4-1:0] node20615;
	wire [4-1:0] node20616;
	wire [4-1:0] node20617;
	wire [4-1:0] node20620;
	wire [4-1:0] node20621;
	wire [4-1:0] node20625;
	wire [4-1:0] node20626;
	wire [4-1:0] node20628;
	wire [4-1:0] node20631;
	wire [4-1:0] node20633;
	wire [4-1:0] node20636;
	wire [4-1:0] node20637;
	wire [4-1:0] node20638;
	wire [4-1:0] node20640;
	wire [4-1:0] node20643;
	wire [4-1:0] node20644;
	wire [4-1:0] node20648;
	wire [4-1:0] node20649;
	wire [4-1:0] node20650;
	wire [4-1:0] node20654;
	wire [4-1:0] node20657;
	wire [4-1:0] node20658;
	wire [4-1:0] node20659;
	wire [4-1:0] node20660;
	wire [4-1:0] node20661;
	wire [4-1:0] node20662;
	wire [4-1:0] node20663;
	wire [4-1:0] node20664;
	wire [4-1:0] node20668;
	wire [4-1:0] node20669;
	wire [4-1:0] node20671;
	wire [4-1:0] node20674;
	wire [4-1:0] node20676;
	wire [4-1:0] node20679;
	wire [4-1:0] node20680;
	wire [4-1:0] node20683;
	wire [4-1:0] node20686;
	wire [4-1:0] node20687;
	wire [4-1:0] node20688;
	wire [4-1:0] node20689;
	wire [4-1:0] node20693;
	wire [4-1:0] node20694;
	wire [4-1:0] node20698;
	wire [4-1:0] node20699;
	wire [4-1:0] node20700;
	wire [4-1:0] node20704;
	wire [4-1:0] node20705;
	wire [4-1:0] node20708;
	wire [4-1:0] node20711;
	wire [4-1:0] node20712;
	wire [4-1:0] node20713;
	wire [4-1:0] node20714;
	wire [4-1:0] node20715;
	wire [4-1:0] node20717;
	wire [4-1:0] node20721;
	wire [4-1:0] node20722;
	wire [4-1:0] node20725;
	wire [4-1:0] node20728;
	wire [4-1:0] node20729;
	wire [4-1:0] node20732;
	wire [4-1:0] node20734;
	wire [4-1:0] node20737;
	wire [4-1:0] node20738;
	wire [4-1:0] node20739;
	wire [4-1:0] node20740;
	wire [4-1:0] node20744;
	wire [4-1:0] node20746;
	wire [4-1:0] node20749;
	wire [4-1:0] node20750;
	wire [4-1:0] node20752;
	wire [4-1:0] node20755;
	wire [4-1:0] node20756;
	wire [4-1:0] node20759;
	wire [4-1:0] node20762;
	wire [4-1:0] node20763;
	wire [4-1:0] node20764;
	wire [4-1:0] node20765;
	wire [4-1:0] node20766;
	wire [4-1:0] node20769;
	wire [4-1:0] node20772;
	wire [4-1:0] node20773;
	wire [4-1:0] node20776;
	wire [4-1:0] node20779;
	wire [4-1:0] node20780;
	wire [4-1:0] node20781;
	wire [4-1:0] node20782;
	wire [4-1:0] node20785;
	wire [4-1:0] node20788;
	wire [4-1:0] node20790;
	wire [4-1:0] node20793;
	wire [4-1:0] node20794;
	wire [4-1:0] node20796;
	wire [4-1:0] node20799;
	wire [4-1:0] node20801;
	wire [4-1:0] node20804;
	wire [4-1:0] node20805;
	wire [4-1:0] node20806;
	wire [4-1:0] node20807;
	wire [4-1:0] node20808;
	wire [4-1:0] node20811;
	wire [4-1:0] node20814;
	wire [4-1:0] node20815;
	wire [4-1:0] node20818;
	wire [4-1:0] node20821;
	wire [4-1:0] node20822;
	wire [4-1:0] node20823;
	wire [4-1:0] node20824;
	wire [4-1:0] node20827;
	wire [4-1:0] node20830;
	wire [4-1:0] node20831;
	wire [4-1:0] node20834;
	wire [4-1:0] node20837;
	wire [4-1:0] node20838;
	wire [4-1:0] node20841;
	wire [4-1:0] node20844;
	wire [4-1:0] node20845;
	wire [4-1:0] node20846;
	wire [4-1:0] node20848;
	wire [4-1:0] node20851;
	wire [4-1:0] node20852;
	wire [4-1:0] node20855;
	wire [4-1:0] node20858;
	wire [4-1:0] node20859;
	wire [4-1:0] node20860;
	wire [4-1:0] node20864;
	wire [4-1:0] node20865;
	wire [4-1:0] node20869;
	wire [4-1:0] node20870;
	wire [4-1:0] node20871;
	wire [4-1:0] node20872;
	wire [4-1:0] node20873;
	wire [4-1:0] node20874;
	wire [4-1:0] node20878;
	wire [4-1:0] node20880;
	wire [4-1:0] node20883;
	wire [4-1:0] node20884;
	wire [4-1:0] node20885;
	wire [4-1:0] node20886;
	wire [4-1:0] node20890;
	wire [4-1:0] node20893;
	wire [4-1:0] node20894;
	wire [4-1:0] node20896;
	wire [4-1:0] node20899;
	wire [4-1:0] node20900;
	wire [4-1:0] node20904;
	wire [4-1:0] node20905;
	wire [4-1:0] node20906;
	wire [4-1:0] node20907;
	wire [4-1:0] node20908;
	wire [4-1:0] node20911;
	wire [4-1:0] node20914;
	wire [4-1:0] node20915;
	wire [4-1:0] node20918;
	wire [4-1:0] node20921;
	wire [4-1:0] node20922;
	wire [4-1:0] node20923;
	wire [4-1:0] node20927;
	wire [4-1:0] node20928;
	wire [4-1:0] node20932;
	wire [4-1:0] node20933;
	wire [4-1:0] node20934;
	wire [4-1:0] node20935;
	wire [4-1:0] node20938;
	wire [4-1:0] node20941;
	wire [4-1:0] node20942;
	wire [4-1:0] node20945;
	wire [4-1:0] node20948;
	wire [4-1:0] node20949;
	wire [4-1:0] node20950;
	wire [4-1:0] node20953;
	wire [4-1:0] node20956;
	wire [4-1:0] node20957;
	wire [4-1:0] node20960;
	wire [4-1:0] node20963;
	wire [4-1:0] node20964;
	wire [4-1:0] node20965;
	wire [4-1:0] node20966;
	wire [4-1:0] node20968;
	wire [4-1:0] node20971;
	wire [4-1:0] node20973;
	wire [4-1:0] node20976;
	wire [4-1:0] node20977;
	wire [4-1:0] node20978;
	wire [4-1:0] node20980;
	wire [4-1:0] node20983;
	wire [4-1:0] node20984;
	wire [4-1:0] node20988;
	wire [4-1:0] node20989;
	wire [4-1:0] node20992;
	wire [4-1:0] node20993;
	wire [4-1:0] node20997;
	wire [4-1:0] node20998;
	wire [4-1:0] node20999;
	wire [4-1:0] node21000;
	wire [4-1:0] node21001;
	wire [4-1:0] node21004;
	wire [4-1:0] node21007;
	wire [4-1:0] node21008;
	wire [4-1:0] node21011;
	wire [4-1:0] node21014;
	wire [4-1:0] node21015;
	wire [4-1:0] node21016;
	wire [4-1:0] node21019;
	wire [4-1:0] node21022;
	wire [4-1:0] node21023;
	wire [4-1:0] node21026;
	wire [4-1:0] node21029;
	wire [4-1:0] node21030;
	wire [4-1:0] node21031;
	wire [4-1:0] node21032;
	wire [4-1:0] node21035;
	wire [4-1:0] node21038;
	wire [4-1:0] node21039;
	wire [4-1:0] node21042;
	wire [4-1:0] node21045;
	wire [4-1:0] node21046;
	wire [4-1:0] node21047;
	wire [4-1:0] node21051;
	wire [4-1:0] node21052;
	wire [4-1:0] node21056;
	wire [4-1:0] node21057;
	wire [4-1:0] node21058;
	wire [4-1:0] node21059;
	wire [4-1:0] node21060;
	wire [4-1:0] node21061;
	wire [4-1:0] node21062;
	wire [4-1:0] node21063;
	wire [4-1:0] node21064;
	wire [4-1:0] node21066;
	wire [4-1:0] node21068;
	wire [4-1:0] node21071;
	wire [4-1:0] node21073;
	wire [4-1:0] node21076;
	wire [4-1:0] node21077;
	wire [4-1:0] node21078;
	wire [4-1:0] node21081;
	wire [4-1:0] node21084;
	wire [4-1:0] node21085;
	wire [4-1:0] node21087;
	wire [4-1:0] node21088;
	wire [4-1:0] node21091;
	wire [4-1:0] node21094;
	wire [4-1:0] node21095;
	wire [4-1:0] node21099;
	wire [4-1:0] node21100;
	wire [4-1:0] node21101;
	wire [4-1:0] node21102;
	wire [4-1:0] node21105;
	wire [4-1:0] node21108;
	wire [4-1:0] node21109;
	wire [4-1:0] node21110;
	wire [4-1:0] node21113;
	wire [4-1:0] node21116;
	wire [4-1:0] node21118;
	wire [4-1:0] node21121;
	wire [4-1:0] node21122;
	wire [4-1:0] node21123;
	wire [4-1:0] node21125;
	wire [4-1:0] node21129;
	wire [4-1:0] node21130;
	wire [4-1:0] node21133;
	wire [4-1:0] node21136;
	wire [4-1:0] node21137;
	wire [4-1:0] node21138;
	wire [4-1:0] node21139;
	wire [4-1:0] node21140;
	wire [4-1:0] node21143;
	wire [4-1:0] node21144;
	wire [4-1:0] node21145;
	wire [4-1:0] node21148;
	wire [4-1:0] node21151;
	wire [4-1:0] node21152;
	wire [4-1:0] node21155;
	wire [4-1:0] node21158;
	wire [4-1:0] node21159;
	wire [4-1:0] node21160;
	wire [4-1:0] node21163;
	wire [4-1:0] node21166;
	wire [4-1:0] node21167;
	wire [4-1:0] node21171;
	wire [4-1:0] node21172;
	wire [4-1:0] node21173;
	wire [4-1:0] node21176;
	wire [4-1:0] node21177;
	wire [4-1:0] node21181;
	wire [4-1:0] node21182;
	wire [4-1:0] node21183;
	wire [4-1:0] node21186;
	wire [4-1:0] node21189;
	wire [4-1:0] node21190;
	wire [4-1:0] node21194;
	wire [4-1:0] node21195;
	wire [4-1:0] node21196;
	wire [4-1:0] node21197;
	wire [4-1:0] node21198;
	wire [4-1:0] node21201;
	wire [4-1:0] node21204;
	wire [4-1:0] node21206;
	wire [4-1:0] node21209;
	wire [4-1:0] node21210;
	wire [4-1:0] node21211;
	wire [4-1:0] node21215;
	wire [4-1:0] node21216;
	wire [4-1:0] node21220;
	wire [4-1:0] node21221;
	wire [4-1:0] node21222;
	wire [4-1:0] node21223;
	wire [4-1:0] node21226;
	wire [4-1:0] node21229;
	wire [4-1:0] node21230;
	wire [4-1:0] node21233;
	wire [4-1:0] node21236;
	wire [4-1:0] node21237;
	wire [4-1:0] node21238;
	wire [4-1:0] node21242;
	wire [4-1:0] node21243;
	wire [4-1:0] node21247;
	wire [4-1:0] node21248;
	wire [4-1:0] node21249;
	wire [4-1:0] node21250;
	wire [4-1:0] node21251;
	wire [4-1:0] node21252;
	wire [4-1:0] node21255;
	wire [4-1:0] node21256;
	wire [4-1:0] node21259;
	wire [4-1:0] node21262;
	wire [4-1:0] node21263;
	wire [4-1:0] node21264;
	wire [4-1:0] node21267;
	wire [4-1:0] node21270;
	wire [4-1:0] node21271;
	wire [4-1:0] node21274;
	wire [4-1:0] node21277;
	wire [4-1:0] node21278;
	wire [4-1:0] node21279;
	wire [4-1:0] node21281;
	wire [4-1:0] node21284;
	wire [4-1:0] node21286;
	wire [4-1:0] node21289;
	wire [4-1:0] node21290;
	wire [4-1:0] node21291;
	wire [4-1:0] node21294;
	wire [4-1:0] node21297;
	wire [4-1:0] node21298;
	wire [4-1:0] node21301;
	wire [4-1:0] node21304;
	wire [4-1:0] node21305;
	wire [4-1:0] node21306;
	wire [4-1:0] node21307;
	wire [4-1:0] node21308;
	wire [4-1:0] node21311;
	wire [4-1:0] node21314;
	wire [4-1:0] node21316;
	wire [4-1:0] node21319;
	wire [4-1:0] node21320;
	wire [4-1:0] node21321;
	wire [4-1:0] node21324;
	wire [4-1:0] node21327;
	wire [4-1:0] node21328;
	wire [4-1:0] node21332;
	wire [4-1:0] node21333;
	wire [4-1:0] node21334;
	wire [4-1:0] node21335;
	wire [4-1:0] node21338;
	wire [4-1:0] node21341;
	wire [4-1:0] node21342;
	wire [4-1:0] node21346;
	wire [4-1:0] node21347;
	wire [4-1:0] node21348;
	wire [4-1:0] node21351;
	wire [4-1:0] node21354;
	wire [4-1:0] node21357;
	wire [4-1:0] node21358;
	wire [4-1:0] node21359;
	wire [4-1:0] node21360;
	wire [4-1:0] node21361;
	wire [4-1:0] node21364;
	wire [4-1:0] node21367;
	wire [4-1:0] node21368;
	wire [4-1:0] node21369;
	wire [4-1:0] node21373;
	wire [4-1:0] node21374;
	wire [4-1:0] node21375;
	wire [4-1:0] node21378;
	wire [4-1:0] node21381;
	wire [4-1:0] node21382;
	wire [4-1:0] node21385;
	wire [4-1:0] node21388;
	wire [4-1:0] node21389;
	wire [4-1:0] node21390;
	wire [4-1:0] node21392;
	wire [4-1:0] node21396;
	wire [4-1:0] node21397;
	wire [4-1:0] node21400;
	wire [4-1:0] node21403;
	wire [4-1:0] node21404;
	wire [4-1:0] node21405;
	wire [4-1:0] node21406;
	wire [4-1:0] node21407;
	wire [4-1:0] node21410;
	wire [4-1:0] node21413;
	wire [4-1:0] node21414;
	wire [4-1:0] node21417;
	wire [4-1:0] node21420;
	wire [4-1:0] node21421;
	wire [4-1:0] node21424;
	wire [4-1:0] node21425;
	wire [4-1:0] node21429;
	wire [4-1:0] node21430;
	wire [4-1:0] node21431;
	wire [4-1:0] node21432;
	wire [4-1:0] node21436;
	wire [4-1:0] node21439;
	wire [4-1:0] node21442;
	wire [4-1:0] node21443;
	wire [4-1:0] node21444;
	wire [4-1:0] node21445;
	wire [4-1:0] node21446;
	wire [4-1:0] node21447;
	wire [4-1:0] node21449;
	wire [4-1:0] node21452;
	wire [4-1:0] node21454;
	wire [4-1:0] node21457;
	wire [4-1:0] node21458;
	wire [4-1:0] node21459;
	wire [4-1:0] node21460;
	wire [4-1:0] node21464;
	wire [4-1:0] node21465;
	wire [4-1:0] node21469;
	wire [4-1:0] node21470;
	wire [4-1:0] node21471;
	wire [4-1:0] node21475;
	wire [4-1:0] node21478;
	wire [4-1:0] node21479;
	wire [4-1:0] node21480;
	wire [4-1:0] node21482;
	wire [4-1:0] node21485;
	wire [4-1:0] node21487;
	wire [4-1:0] node21490;
	wire [4-1:0] node21491;
	wire [4-1:0] node21492;
	wire [4-1:0] node21494;
	wire [4-1:0] node21497;
	wire [4-1:0] node21498;
	wire [4-1:0] node21502;
	wire [4-1:0] node21503;
	wire [4-1:0] node21504;
	wire [4-1:0] node21508;
	wire [4-1:0] node21509;
	wire [4-1:0] node21513;
	wire [4-1:0] node21514;
	wire [4-1:0] node21515;
	wire [4-1:0] node21516;
	wire [4-1:0] node21517;
	wire [4-1:0] node21519;
	wire [4-1:0] node21522;
	wire [4-1:0] node21523;
	wire [4-1:0] node21527;
	wire [4-1:0] node21528;
	wire [4-1:0] node21529;
	wire [4-1:0] node21533;
	wire [4-1:0] node21534;
	wire [4-1:0] node21538;
	wire [4-1:0] node21539;
	wire [4-1:0] node21540;
	wire [4-1:0] node21542;
	wire [4-1:0] node21545;
	wire [4-1:0] node21547;
	wire [4-1:0] node21550;
	wire [4-1:0] node21551;
	wire [4-1:0] node21553;
	wire [4-1:0] node21556;
	wire [4-1:0] node21557;
	wire [4-1:0] node21561;
	wire [4-1:0] node21562;
	wire [4-1:0] node21563;
	wire [4-1:0] node21564;
	wire [4-1:0] node21565;
	wire [4-1:0] node21569;
	wire [4-1:0] node21570;
	wire [4-1:0] node21574;
	wire [4-1:0] node21575;
	wire [4-1:0] node21576;
	wire [4-1:0] node21580;
	wire [4-1:0] node21581;
	wire [4-1:0] node21585;
	wire [4-1:0] node21586;
	wire [4-1:0] node21587;
	wire [4-1:0] node21588;
	wire [4-1:0] node21592;
	wire [4-1:0] node21594;
	wire [4-1:0] node21597;
	wire [4-1:0] node21598;
	wire [4-1:0] node21600;
	wire [4-1:0] node21603;
	wire [4-1:0] node21604;
	wire [4-1:0] node21608;
	wire [4-1:0] node21609;
	wire [4-1:0] node21610;
	wire [4-1:0] node21611;
	wire [4-1:0] node21612;
	wire [4-1:0] node21613;
	wire [4-1:0] node21615;
	wire [4-1:0] node21618;
	wire [4-1:0] node21619;
	wire [4-1:0] node21623;
	wire [4-1:0] node21624;
	wire [4-1:0] node21625;
	wire [4-1:0] node21629;
	wire [4-1:0] node21631;
	wire [4-1:0] node21634;
	wire [4-1:0] node21635;
	wire [4-1:0] node21636;
	wire [4-1:0] node21637;
	wire [4-1:0] node21641;
	wire [4-1:0] node21644;
	wire [4-1:0] node21645;
	wire [4-1:0] node21647;
	wire [4-1:0] node21650;
	wire [4-1:0] node21652;
	wire [4-1:0] node21655;
	wire [4-1:0] node21656;
	wire [4-1:0] node21657;
	wire [4-1:0] node21658;
	wire [4-1:0] node21660;
	wire [4-1:0] node21663;
	wire [4-1:0] node21665;
	wire [4-1:0] node21668;
	wire [4-1:0] node21669;
	wire [4-1:0] node21670;
	wire [4-1:0] node21674;
	wire [4-1:0] node21676;
	wire [4-1:0] node21679;
	wire [4-1:0] node21680;
	wire [4-1:0] node21681;
	wire [4-1:0] node21682;
	wire [4-1:0] node21686;
	wire [4-1:0] node21687;
	wire [4-1:0] node21691;
	wire [4-1:0] node21692;
	wire [4-1:0] node21696;
	wire [4-1:0] node21697;
	wire [4-1:0] node21698;
	wire [4-1:0] node21699;
	wire [4-1:0] node21700;
	wire [4-1:0] node21702;
	wire [4-1:0] node21705;
	wire [4-1:0] node21707;
	wire [4-1:0] node21710;
	wire [4-1:0] node21711;
	wire [4-1:0] node21712;
	wire [4-1:0] node21716;
	wire [4-1:0] node21717;
	wire [4-1:0] node21721;
	wire [4-1:0] node21722;
	wire [4-1:0] node21724;
	wire [4-1:0] node21727;
	wire [4-1:0] node21728;
	wire [4-1:0] node21732;
	wire [4-1:0] node21733;
	wire [4-1:0] node21734;
	wire [4-1:0] node21735;
	wire [4-1:0] node21736;
	wire [4-1:0] node21740;
	wire [4-1:0] node21742;
	wire [4-1:0] node21745;
	wire [4-1:0] node21746;
	wire [4-1:0] node21748;
	wire [4-1:0] node21751;
	wire [4-1:0] node21753;
	wire [4-1:0] node21756;
	wire [4-1:0] node21757;
	wire [4-1:0] node21759;
	wire [4-1:0] node21762;
	wire [4-1:0] node21763;
	wire [4-1:0] node21767;
	wire [4-1:0] node21768;
	wire [4-1:0] node21769;
	wire [4-1:0] node21770;
	wire [4-1:0] node21771;
	wire [4-1:0] node21772;
	wire [4-1:0] node21773;
	wire [4-1:0] node21775;
	wire [4-1:0] node21777;
	wire [4-1:0] node21780;
	wire [4-1:0] node21782;
	wire [4-1:0] node21785;
	wire [4-1:0] node21786;
	wire [4-1:0] node21788;
	wire [4-1:0] node21791;
	wire [4-1:0] node21792;
	wire [4-1:0] node21793;
	wire [4-1:0] node21796;
	wire [4-1:0] node21799;
	wire [4-1:0] node21800;
	wire [4-1:0] node21804;
	wire [4-1:0] node21805;
	wire [4-1:0] node21806;
	wire [4-1:0] node21808;
	wire [4-1:0] node21811;
	wire [4-1:0] node21812;
	wire [4-1:0] node21814;
	wire [4-1:0] node21815;
	wire [4-1:0] node21818;
	wire [4-1:0] node21821;
	wire [4-1:0] node21823;
	wire [4-1:0] node21826;
	wire [4-1:0] node21827;
	wire [4-1:0] node21828;
	wire [4-1:0] node21830;
	wire [4-1:0] node21834;
	wire [4-1:0] node21835;
	wire [4-1:0] node21839;
	wire [4-1:0] node21840;
	wire [4-1:0] node21841;
	wire [4-1:0] node21842;
	wire [4-1:0] node21843;
	wire [4-1:0] node21846;
	wire [4-1:0] node21847;
	wire [4-1:0] node21850;
	wire [4-1:0] node21853;
	wire [4-1:0] node21854;
	wire [4-1:0] node21855;
	wire [4-1:0] node21858;
	wire [4-1:0] node21861;
	wire [4-1:0] node21862;
	wire [4-1:0] node21865;
	wire [4-1:0] node21868;
	wire [4-1:0] node21869;
	wire [4-1:0] node21870;
	wire [4-1:0] node21873;
	wire [4-1:0] node21874;
	wire [4-1:0] node21877;
	wire [4-1:0] node21880;
	wire [4-1:0] node21881;
	wire [4-1:0] node21883;
	wire [4-1:0] node21886;
	wire [4-1:0] node21887;
	wire [4-1:0] node21891;
	wire [4-1:0] node21892;
	wire [4-1:0] node21893;
	wire [4-1:0] node21894;
	wire [4-1:0] node21895;
	wire [4-1:0] node21898;
	wire [4-1:0] node21901;
	wire [4-1:0] node21902;
	wire [4-1:0] node21905;
	wire [4-1:0] node21908;
	wire [4-1:0] node21909;
	wire [4-1:0] node21910;
	wire [4-1:0] node21913;
	wire [4-1:0] node21916;
	wire [4-1:0] node21917;
	wire [4-1:0] node21921;
	wire [4-1:0] node21922;
	wire [4-1:0] node21923;
	wire [4-1:0] node21924;
	wire [4-1:0] node21927;
	wire [4-1:0] node21930;
	wire [4-1:0] node21931;
	wire [4-1:0] node21934;
	wire [4-1:0] node21937;
	wire [4-1:0] node21938;
	wire [4-1:0] node21939;
	wire [4-1:0] node21940;
	wire [4-1:0] node21943;
	wire [4-1:0] node21946;
	wire [4-1:0] node21947;
	wire [4-1:0] node21950;
	wire [4-1:0] node21953;
	wire [4-1:0] node21956;
	wire [4-1:0] node21957;
	wire [4-1:0] node21958;
	wire [4-1:0] node21959;
	wire [4-1:0] node21960;
	wire [4-1:0] node21961;
	wire [4-1:0] node21963;
	wire [4-1:0] node21966;
	wire [4-1:0] node21967;
	wire [4-1:0] node21970;
	wire [4-1:0] node21973;
	wire [4-1:0] node21974;
	wire [4-1:0] node21976;
	wire [4-1:0] node21979;
	wire [4-1:0] node21980;
	wire [4-1:0] node21983;
	wire [4-1:0] node21986;
	wire [4-1:0] node21987;
	wire [4-1:0] node21988;
	wire [4-1:0] node21990;
	wire [4-1:0] node21993;
	wire [4-1:0] node21995;
	wire [4-1:0] node21998;
	wire [4-1:0] node21999;
	wire [4-1:0] node22001;
	wire [4-1:0] node22004;
	wire [4-1:0] node22005;
	wire [4-1:0] node22008;
	wire [4-1:0] node22011;
	wire [4-1:0] node22012;
	wire [4-1:0] node22013;
	wire [4-1:0] node22014;
	wire [4-1:0] node22015;
	wire [4-1:0] node22018;
	wire [4-1:0] node22021;
	wire [4-1:0] node22023;
	wire [4-1:0] node22026;
	wire [4-1:0] node22027;
	wire [4-1:0] node22028;
	wire [4-1:0] node22031;
	wire [4-1:0] node22034;
	wire [4-1:0] node22035;
	wire [4-1:0] node22038;
	wire [4-1:0] node22041;
	wire [4-1:0] node22042;
	wire [4-1:0] node22043;
	wire [4-1:0] node22045;
	wire [4-1:0] node22048;
	wire [4-1:0] node22049;
	wire [4-1:0] node22053;
	wire [4-1:0] node22054;
	wire [4-1:0] node22055;
	wire [4-1:0] node22058;
	wire [4-1:0] node22061;
	wire [4-1:0] node22062;
	wire [4-1:0] node22066;
	wire [4-1:0] node22067;
	wire [4-1:0] node22068;
	wire [4-1:0] node22069;
	wire [4-1:0] node22070;
	wire [4-1:0] node22073;
	wire [4-1:0] node22076;
	wire [4-1:0] node22077;
	wire [4-1:0] node22078;
	wire [4-1:0] node22081;
	wire [4-1:0] node22084;
	wire [4-1:0] node22086;
	wire [4-1:0] node22089;
	wire [4-1:0] node22090;
	wire [4-1:0] node22091;
	wire [4-1:0] node22093;
	wire [4-1:0] node22097;
	wire [4-1:0] node22098;
	wire [4-1:0] node22101;
	wire [4-1:0] node22104;
	wire [4-1:0] node22105;
	wire [4-1:0] node22106;
	wire [4-1:0] node22107;
	wire [4-1:0] node22109;
	wire [4-1:0] node22112;
	wire [4-1:0] node22113;
	wire [4-1:0] node22114;
	wire [4-1:0] node22118;
	wire [4-1:0] node22119;
	wire [4-1:0] node22122;
	wire [4-1:0] node22125;
	wire [4-1:0] node22126;
	wire [4-1:0] node22129;
	wire [4-1:0] node22132;
	wire [4-1:0] node22133;
	wire [4-1:0] node22134;
	wire [4-1:0] node22137;
	wire [4-1:0] node22140;
	wire [4-1:0] node22141;
	wire [4-1:0] node22142;
	wire [4-1:0] node22147;
	wire [4-1:0] node22148;
	wire [4-1:0] node22149;
	wire [4-1:0] node22150;
	wire [4-1:0] node22151;
	wire [4-1:0] node22152;
	wire [4-1:0] node22154;
	wire [4-1:0] node22157;
	wire [4-1:0] node22158;
	wire [4-1:0] node22161;
	wire [4-1:0] node22164;
	wire [4-1:0] node22165;
	wire [4-1:0] node22166;
	wire [4-1:0] node22169;
	wire [4-1:0] node22170;
	wire [4-1:0] node22174;
	wire [4-1:0] node22175;
	wire [4-1:0] node22176;
	wire [4-1:0] node22179;
	wire [4-1:0] node22182;
	wire [4-1:0] node22185;
	wire [4-1:0] node22186;
	wire [4-1:0] node22187;
	wire [4-1:0] node22188;
	wire [4-1:0] node22190;
	wire [4-1:0] node22193;
	wire [4-1:0] node22195;
	wire [4-1:0] node22198;
	wire [4-1:0] node22199;
	wire [4-1:0] node22201;
	wire [4-1:0] node22204;
	wire [4-1:0] node22206;
	wire [4-1:0] node22209;
	wire [4-1:0] node22210;
	wire [4-1:0] node22212;
	wire [4-1:0] node22215;
	wire [4-1:0] node22216;
	wire [4-1:0] node22218;
	wire [4-1:0] node22221;
	wire [4-1:0] node22222;
	wire [4-1:0] node22225;
	wire [4-1:0] node22228;
	wire [4-1:0] node22229;
	wire [4-1:0] node22230;
	wire [4-1:0] node22231;
	wire [4-1:0] node22233;
	wire [4-1:0] node22236;
	wire [4-1:0] node22237;
	wire [4-1:0] node22241;
	wire [4-1:0] node22242;
	wire [4-1:0] node22243;
	wire [4-1:0] node22245;
	wire [4-1:0] node22248;
	wire [4-1:0] node22249;
	wire [4-1:0] node22253;
	wire [4-1:0] node22254;
	wire [4-1:0] node22255;
	wire [4-1:0] node22259;
	wire [4-1:0] node22260;
	wire [4-1:0] node22264;
	wire [4-1:0] node22265;
	wire [4-1:0] node22266;
	wire [4-1:0] node22267;
	wire [4-1:0] node22269;
	wire [4-1:0] node22272;
	wire [4-1:0] node22273;
	wire [4-1:0] node22277;
	wire [4-1:0] node22278;
	wire [4-1:0] node22279;
	wire [4-1:0] node22283;
	wire [4-1:0] node22284;
	wire [4-1:0] node22288;
	wire [4-1:0] node22289;
	wire [4-1:0] node22290;
	wire [4-1:0] node22292;
	wire [4-1:0] node22295;
	wire [4-1:0] node22297;
	wire [4-1:0] node22300;
	wire [4-1:0] node22301;
	wire [4-1:0] node22303;
	wire [4-1:0] node22306;
	wire [4-1:0] node22307;
	wire [4-1:0] node22311;
	wire [4-1:0] node22312;
	wire [4-1:0] node22313;
	wire [4-1:0] node22314;
	wire [4-1:0] node22315;
	wire [4-1:0] node22317;
	wire [4-1:0] node22320;
	wire [4-1:0] node22322;
	wire [4-1:0] node22325;
	wire [4-1:0] node22326;
	wire [4-1:0] node22327;
	wire [4-1:0] node22329;
	wire [4-1:0] node22332;
	wire [4-1:0] node22334;
	wire [4-1:0] node22337;
	wire [4-1:0] node22339;
	wire [4-1:0] node22340;
	wire [4-1:0] node22344;
	wire [4-1:0] node22345;
	wire [4-1:0] node22346;
	wire [4-1:0] node22347;
	wire [4-1:0] node22349;
	wire [4-1:0] node22352;
	wire [4-1:0] node22353;
	wire [4-1:0] node22357;
	wire [4-1:0] node22358;
	wire [4-1:0] node22359;
	wire [4-1:0] node22363;
	wire [4-1:0] node22364;
	wire [4-1:0] node22368;
	wire [4-1:0] node22369;
	wire [4-1:0] node22370;
	wire [4-1:0] node22372;
	wire [4-1:0] node22375;
	wire [4-1:0] node22377;
	wire [4-1:0] node22380;
	wire [4-1:0] node22381;
	wire [4-1:0] node22382;
	wire [4-1:0] node22386;
	wire [4-1:0] node22387;
	wire [4-1:0] node22391;
	wire [4-1:0] node22392;
	wire [4-1:0] node22393;
	wire [4-1:0] node22394;
	wire [4-1:0] node22395;
	wire [4-1:0] node22396;
	wire [4-1:0] node22399;
	wire [4-1:0] node22402;
	wire [4-1:0] node22403;
	wire [4-1:0] node22406;
	wire [4-1:0] node22409;
	wire [4-1:0] node22410;
	wire [4-1:0] node22413;
	wire [4-1:0] node22414;
	wire [4-1:0] node22418;
	wire [4-1:0] node22419;
	wire [4-1:0] node22420;
	wire [4-1:0] node22421;
	wire [4-1:0] node22424;
	wire [4-1:0] node22427;
	wire [4-1:0] node22428;
	wire [4-1:0] node22432;
	wire [4-1:0] node22433;
	wire [4-1:0] node22434;
	wire [4-1:0] node22437;
	wire [4-1:0] node22440;
	wire [4-1:0] node22441;
	wire [4-1:0] node22445;
	wire [4-1:0] node22446;
	wire [4-1:0] node22447;
	wire [4-1:0] node22448;
	wire [4-1:0] node22451;
	wire [4-1:0] node22453;
	wire [4-1:0] node22456;
	wire [4-1:0] node22457;
	wire [4-1:0] node22458;
	wire [4-1:0] node22461;
	wire [4-1:0] node22464;
	wire [4-1:0] node22465;
	wire [4-1:0] node22468;
	wire [4-1:0] node22471;
	wire [4-1:0] node22472;
	wire [4-1:0] node22473;
	wire [4-1:0] node22477;
	wire [4-1:0] node22478;
	wire [4-1:0] node22479;
	wire [4-1:0] node22484;
	wire [4-1:0] node22485;
	wire [4-1:0] node22486;
	wire [4-1:0] node22487;
	wire [4-1:0] node22488;
	wire [4-1:0] node22489;
	wire [4-1:0] node22490;
	wire [4-1:0] node22491;
	wire [4-1:0] node22493;
	wire [4-1:0] node22496;
	wire [4-1:0] node22497;
	wire [4-1:0] node22500;
	wire [4-1:0] node22501;
	wire [4-1:0] node22505;
	wire [4-1:0] node22506;
	wire [4-1:0] node22507;
	wire [4-1:0] node22509;
	wire [4-1:0] node22512;
	wire [4-1:0] node22515;
	wire [4-1:0] node22516;
	wire [4-1:0] node22517;
	wire [4-1:0] node22520;
	wire [4-1:0] node22523;
	wire [4-1:0] node22526;
	wire [4-1:0] node22527;
	wire [4-1:0] node22528;
	wire [4-1:0] node22529;
	wire [4-1:0] node22531;
	wire [4-1:0] node22534;
	wire [4-1:0] node22536;
	wire [4-1:0] node22539;
	wire [4-1:0] node22540;
	wire [4-1:0] node22543;
	wire [4-1:0] node22544;
	wire [4-1:0] node22547;
	wire [4-1:0] node22550;
	wire [4-1:0] node22551;
	wire [4-1:0] node22552;
	wire [4-1:0] node22555;
	wire [4-1:0] node22558;
	wire [4-1:0] node22559;
	wire [4-1:0] node22561;
	wire [4-1:0] node22564;
	wire [4-1:0] node22565;
	wire [4-1:0] node22566;
	wire [4-1:0] node22569;
	wire [4-1:0] node22572;
	wire [4-1:0] node22573;
	wire [4-1:0] node22576;
	wire [4-1:0] node22579;
	wire [4-1:0] node22580;
	wire [4-1:0] node22581;
	wire [4-1:0] node22582;
	wire [4-1:0] node22583;
	wire [4-1:0] node22586;
	wire [4-1:0] node22587;
	wire [4-1:0] node22590;
	wire [4-1:0] node22593;
	wire [4-1:0] node22594;
	wire [4-1:0] node22595;
	wire [4-1:0] node22598;
	wire [4-1:0] node22601;
	wire [4-1:0] node22602;
	wire [4-1:0] node22605;
	wire [4-1:0] node22608;
	wire [4-1:0] node22609;
	wire [4-1:0] node22610;
	wire [4-1:0] node22612;
	wire [4-1:0] node22615;
	wire [4-1:0] node22617;
	wire [4-1:0] node22620;
	wire [4-1:0] node22621;
	wire [4-1:0] node22622;
	wire [4-1:0] node22625;
	wire [4-1:0] node22628;
	wire [4-1:0] node22629;
	wire [4-1:0] node22632;
	wire [4-1:0] node22635;
	wire [4-1:0] node22636;
	wire [4-1:0] node22637;
	wire [4-1:0] node22638;
	wire [4-1:0] node22640;
	wire [4-1:0] node22643;
	wire [4-1:0] node22645;
	wire [4-1:0] node22648;
	wire [4-1:0] node22650;
	wire [4-1:0] node22653;
	wire [4-1:0] node22654;
	wire [4-1:0] node22655;
	wire [4-1:0] node22657;
	wire [4-1:0] node22660;
	wire [4-1:0] node22662;
	wire [4-1:0] node22665;
	wire [4-1:0] node22666;
	wire [4-1:0] node22668;
	wire [4-1:0] node22671;
	wire [4-1:0] node22672;
	wire [4-1:0] node22673;
	wire [4-1:0] node22676;
	wire [4-1:0] node22679;
	wire [4-1:0] node22680;
	wire [4-1:0] node22683;
	wire [4-1:0] node22686;
	wire [4-1:0] node22687;
	wire [4-1:0] node22688;
	wire [4-1:0] node22689;
	wire [4-1:0] node22690;
	wire [4-1:0] node22692;
	wire [4-1:0] node22694;
	wire [4-1:0] node22697;
	wire [4-1:0] node22699;
	wire [4-1:0] node22702;
	wire [4-1:0] node22703;
	wire [4-1:0] node22704;
	wire [4-1:0] node22705;
	wire [4-1:0] node22708;
	wire [4-1:0] node22711;
	wire [4-1:0] node22712;
	wire [4-1:0] node22715;
	wire [4-1:0] node22718;
	wire [4-1:0] node22719;
	wire [4-1:0] node22720;
	wire [4-1:0] node22724;
	wire [4-1:0] node22727;
	wire [4-1:0] node22728;
	wire [4-1:0] node22729;
	wire [4-1:0] node22730;
	wire [4-1:0] node22734;
	wire [4-1:0] node22735;
	wire [4-1:0] node22736;
	wire [4-1:0] node22739;
	wire [4-1:0] node22742;
	wire [4-1:0] node22744;
	wire [4-1:0] node22747;
	wire [4-1:0] node22748;
	wire [4-1:0] node22749;
	wire [4-1:0] node22750;
	wire [4-1:0] node22754;
	wire [4-1:0] node22757;
	wire [4-1:0] node22758;
	wire [4-1:0] node22759;
	wire [4-1:0] node22762;
	wire [4-1:0] node22765;
	wire [4-1:0] node22766;
	wire [4-1:0] node22769;
	wire [4-1:0] node22772;
	wire [4-1:0] node22773;
	wire [4-1:0] node22774;
	wire [4-1:0] node22775;
	wire [4-1:0] node22777;
	wire [4-1:0] node22780;
	wire [4-1:0] node22781;
	wire [4-1:0] node22784;
	wire [4-1:0] node22785;
	wire [4-1:0] node22789;
	wire [4-1:0] node22790;
	wire [4-1:0] node22791;
	wire [4-1:0] node22793;
	wire [4-1:0] node22796;
	wire [4-1:0] node22799;
	wire [4-1:0] node22800;
	wire [4-1:0] node22802;
	wire [4-1:0] node22805;
	wire [4-1:0] node22808;
	wire [4-1:0] node22809;
	wire [4-1:0] node22810;
	wire [4-1:0] node22811;
	wire [4-1:0] node22813;
	wire [4-1:0] node22816;
	wire [4-1:0] node22818;
	wire [4-1:0] node22821;
	wire [4-1:0] node22822;
	wire [4-1:0] node22824;
	wire [4-1:0] node22827;
	wire [4-1:0] node22828;
	wire [4-1:0] node22831;
	wire [4-1:0] node22834;
	wire [4-1:0] node22835;
	wire [4-1:0] node22836;
	wire [4-1:0] node22838;
	wire [4-1:0] node22841;
	wire [4-1:0] node22843;
	wire [4-1:0] node22846;
	wire [4-1:0] node22847;
	wire [4-1:0] node22849;
	wire [4-1:0] node22852;
	wire [4-1:0] node22854;
	wire [4-1:0] node22857;
	wire [4-1:0] node22858;
	wire [4-1:0] node22859;
	wire [4-1:0] node22860;
	wire [4-1:0] node22861;
	wire [4-1:0] node22862;
	wire [4-1:0] node22863;
	wire [4-1:0] node22866;
	wire [4-1:0] node22869;
	wire [4-1:0] node22870;
	wire [4-1:0] node22871;
	wire [4-1:0] node22874;
	wire [4-1:0] node22877;
	wire [4-1:0] node22878;
	wire [4-1:0] node22881;
	wire [4-1:0] node22884;
	wire [4-1:0] node22885;
	wire [4-1:0] node22888;
	wire [4-1:0] node22891;
	wire [4-1:0] node22892;
	wire [4-1:0] node22893;
	wire [4-1:0] node22894;
	wire [4-1:0] node22895;
	wire [4-1:0] node22898;
	wire [4-1:0] node22901;
	wire [4-1:0] node22902;
	wire [4-1:0] node22903;
	wire [4-1:0] node22906;
	wire [4-1:0] node22909;
	wire [4-1:0] node22910;
	wire [4-1:0] node22913;
	wire [4-1:0] node22916;
	wire [4-1:0] node22917;
	wire [4-1:0] node22918;
	wire [4-1:0] node22919;
	wire [4-1:0] node22922;
	wire [4-1:0] node22926;
	wire [4-1:0] node22927;
	wire [4-1:0] node22928;
	wire [4-1:0] node22931;
	wire [4-1:0] node22934;
	wire [4-1:0] node22935;
	wire [4-1:0] node22939;
	wire [4-1:0] node22940;
	wire [4-1:0] node22941;
	wire [4-1:0] node22942;
	wire [4-1:0] node22945;
	wire [4-1:0] node22948;
	wire [4-1:0] node22949;
	wire [4-1:0] node22952;
	wire [4-1:0] node22955;
	wire [4-1:0] node22956;
	wire [4-1:0] node22957;
	wire [4-1:0] node22958;
	wire [4-1:0] node22961;
	wire [4-1:0] node22964;
	wire [4-1:0] node22965;
	wire [4-1:0] node22968;
	wire [4-1:0] node22971;
	wire [4-1:0] node22973;
	wire [4-1:0] node22976;
	wire [4-1:0] node22977;
	wire [4-1:0] node22978;
	wire [4-1:0] node22979;
	wire [4-1:0] node22980;
	wire [4-1:0] node22983;
	wire [4-1:0] node22986;
	wire [4-1:0] node22987;
	wire [4-1:0] node22990;
	wire [4-1:0] node22993;
	wire [4-1:0] node22994;
	wire [4-1:0] node22995;
	wire [4-1:0] node22996;
	wire [4-1:0] node22997;
	wire [4-1:0] node23001;
	wire [4-1:0] node23004;
	wire [4-1:0] node23005;
	wire [4-1:0] node23008;
	wire [4-1:0] node23011;
	wire [4-1:0] node23012;
	wire [4-1:0] node23015;
	wire [4-1:0] node23018;
	wire [4-1:0] node23019;
	wire [4-1:0] node23020;
	wire [4-1:0] node23021;
	wire [4-1:0] node23022;
	wire [4-1:0] node23025;
	wire [4-1:0] node23028;
	wire [4-1:0] node23030;
	wire [4-1:0] node23033;
	wire [4-1:0] node23034;
	wire [4-1:0] node23035;
	wire [4-1:0] node23039;
	wire [4-1:0] node23040;
	wire [4-1:0] node23041;
	wire [4-1:0] node23044;
	wire [4-1:0] node23048;
	wire [4-1:0] node23049;
	wire [4-1:0] node23050;
	wire [4-1:0] node23051;
	wire [4-1:0] node23052;
	wire [4-1:0] node23055;
	wire [4-1:0] node23058;
	wire [4-1:0] node23059;
	wire [4-1:0] node23062;
	wire [4-1:0] node23065;
	wire [4-1:0] node23067;
	wire [4-1:0] node23070;
	wire [4-1:0] node23071;
	wire [4-1:0] node23072;
	wire [4-1:0] node23073;
	wire [4-1:0] node23076;
	wire [4-1:0] node23079;
	wire [4-1:0] node23081;
	wire [4-1:0] node23084;
	wire [4-1:0] node23085;
	wire [4-1:0] node23086;
	wire [4-1:0] node23090;
	wire [4-1:0] node23091;
	wire [4-1:0] node23094;
	wire [4-1:0] node23097;
	wire [4-1:0] node23098;
	wire [4-1:0] node23099;
	wire [4-1:0] node23100;
	wire [4-1:0] node23101;
	wire [4-1:0] node23102;
	wire [4-1:0] node23103;
	wire [4-1:0] node23104;
	wire [4-1:0] node23107;
	wire [4-1:0] node23110;
	wire [4-1:0] node23111;
	wire [4-1:0] node23114;
	wire [4-1:0] node23117;
	wire [4-1:0] node23118;
	wire [4-1:0] node23119;
	wire [4-1:0] node23123;
	wire [4-1:0] node23124;
	wire [4-1:0] node23127;
	wire [4-1:0] node23130;
	wire [4-1:0] node23131;
	wire [4-1:0] node23132;
	wire [4-1:0] node23133;
	wire [4-1:0] node23136;
	wire [4-1:0] node23139;
	wire [4-1:0] node23140;
	wire [4-1:0] node23143;
	wire [4-1:0] node23146;
	wire [4-1:0] node23148;
	wire [4-1:0] node23149;
	wire [4-1:0] node23152;
	wire [4-1:0] node23155;
	wire [4-1:0] node23156;
	wire [4-1:0] node23157;
	wire [4-1:0] node23158;
	wire [4-1:0] node23159;
	wire [4-1:0] node23162;
	wire [4-1:0] node23165;
	wire [4-1:0] node23166;
	wire [4-1:0] node23169;
	wire [4-1:0] node23172;
	wire [4-1:0] node23173;
	wire [4-1:0] node23176;
	wire [4-1:0] node23179;
	wire [4-1:0] node23180;
	wire [4-1:0] node23181;
	wire [4-1:0] node23182;
	wire [4-1:0] node23185;
	wire [4-1:0] node23188;
	wire [4-1:0] node23189;
	wire [4-1:0] node23193;
	wire [4-1:0] node23194;
	wire [4-1:0] node23197;
	wire [4-1:0] node23200;
	wire [4-1:0] node23201;
	wire [4-1:0] node23202;
	wire [4-1:0] node23203;
	wire [4-1:0] node23204;
	wire [4-1:0] node23205;
	wire [4-1:0] node23208;
	wire [4-1:0] node23211;
	wire [4-1:0] node23212;
	wire [4-1:0] node23216;
	wire [4-1:0] node23217;
	wire [4-1:0] node23218;
	wire [4-1:0] node23221;
	wire [4-1:0] node23224;
	wire [4-1:0] node23225;
	wire [4-1:0] node23228;
	wire [4-1:0] node23231;
	wire [4-1:0] node23232;
	wire [4-1:0] node23233;
	wire [4-1:0] node23236;
	wire [4-1:0] node23239;
	wire [4-1:0] node23240;
	wire [4-1:0] node23241;
	wire [4-1:0] node23244;
	wire [4-1:0] node23247;
	wire [4-1:0] node23248;
	wire [4-1:0] node23251;
	wire [4-1:0] node23254;
	wire [4-1:0] node23255;
	wire [4-1:0] node23256;
	wire [4-1:0] node23257;
	wire [4-1:0] node23258;
	wire [4-1:0] node23261;
	wire [4-1:0] node23264;
	wire [4-1:0] node23265;
	wire [4-1:0] node23268;
	wire [4-1:0] node23271;
	wire [4-1:0] node23273;
	wire [4-1:0] node23274;
	wire [4-1:0] node23277;
	wire [4-1:0] node23280;
	wire [4-1:0] node23281;
	wire [4-1:0] node23282;
	wire [4-1:0] node23284;
	wire [4-1:0] node23287;
	wire [4-1:0] node23288;
	wire [4-1:0] node23292;
	wire [4-1:0] node23293;
	wire [4-1:0] node23296;
	wire [4-1:0] node23299;
	wire [4-1:0] node23300;
	wire [4-1:0] node23301;
	wire [4-1:0] node23302;
	wire [4-1:0] node23303;
	wire [4-1:0] node23304;
	wire [4-1:0] node23307;
	wire [4-1:0] node23308;
	wire [4-1:0] node23311;
	wire [4-1:0] node23314;
	wire [4-1:0] node23315;
	wire [4-1:0] node23317;
	wire [4-1:0] node23320;
	wire [4-1:0] node23321;
	wire [4-1:0] node23324;
	wire [4-1:0] node23327;
	wire [4-1:0] node23328;
	wire [4-1:0] node23329;
	wire [4-1:0] node23330;
	wire [4-1:0] node23333;
	wire [4-1:0] node23336;
	wire [4-1:0] node23338;
	wire [4-1:0] node23341;
	wire [4-1:0] node23343;
	wire [4-1:0] node23344;
	wire [4-1:0] node23348;
	wire [4-1:0] node23349;
	wire [4-1:0] node23350;
	wire [4-1:0] node23352;
	wire [4-1:0] node23353;
	wire [4-1:0] node23357;
	wire [4-1:0] node23358;
	wire [4-1:0] node23359;
	wire [4-1:0] node23362;
	wire [4-1:0] node23365;
	wire [4-1:0] node23368;
	wire [4-1:0] node23369;
	wire [4-1:0] node23370;
	wire [4-1:0] node23372;
	wire [4-1:0] node23375;
	wire [4-1:0] node23376;
	wire [4-1:0] node23379;
	wire [4-1:0] node23382;
	wire [4-1:0] node23383;
	wire [4-1:0] node23385;
	wire [4-1:0] node23388;
	wire [4-1:0] node23391;
	wire [4-1:0] node23392;
	wire [4-1:0] node23393;
	wire [4-1:0] node23394;
	wire [4-1:0] node23395;
	wire [4-1:0] node23397;
	wire [4-1:0] node23400;
	wire [4-1:0] node23401;
	wire [4-1:0] node23405;
	wire [4-1:0] node23406;
	wire [4-1:0] node23407;
	wire [4-1:0] node23411;
	wire [4-1:0] node23412;
	wire [4-1:0] node23415;
	wire [4-1:0] node23418;
	wire [4-1:0] node23419;
	wire [4-1:0] node23420;
	wire [4-1:0] node23421;
	wire [4-1:0] node23425;
	wire [4-1:0] node23427;
	wire [4-1:0] node23430;
	wire [4-1:0] node23432;
	wire [4-1:0] node23433;
	wire [4-1:0] node23436;
	wire [4-1:0] node23439;
	wire [4-1:0] node23440;
	wire [4-1:0] node23441;
	wire [4-1:0] node23442;
	wire [4-1:0] node23443;
	wire [4-1:0] node23447;
	wire [4-1:0] node23449;
	wire [4-1:0] node23452;
	wire [4-1:0] node23453;
	wire [4-1:0] node23456;
	wire [4-1:0] node23457;
	wire [4-1:0] node23460;
	wire [4-1:0] node23463;
	wire [4-1:0] node23464;
	wire [4-1:0] node23465;
	wire [4-1:0] node23466;
	wire [4-1:0] node23469;
	wire [4-1:0] node23472;
	wire [4-1:0] node23473;
	wire [4-1:0] node23476;
	wire [4-1:0] node23479;
	wire [4-1:0] node23480;
	wire [4-1:0] node23481;
	wire [4-1:0] node23486;
	wire [4-1:0] node23487;
	wire [4-1:0] node23488;
	wire [4-1:0] node23489;
	wire [4-1:0] node23490;
	wire [4-1:0] node23491;
	wire [4-1:0] node23492;
	wire [4-1:0] node23493;
	wire [4-1:0] node23495;
	wire [4-1:0] node23498;
	wire [4-1:0] node23500;
	wire [4-1:0] node23503;
	wire [4-1:0] node23504;
	wire [4-1:0] node23506;
	wire [4-1:0] node23509;
	wire [4-1:0] node23510;
	wire [4-1:0] node23514;
	wire [4-1:0] node23515;
	wire [4-1:0] node23516;
	wire [4-1:0] node23518;
	wire [4-1:0] node23521;
	wire [4-1:0] node23522;
	wire [4-1:0] node23526;
	wire [4-1:0] node23527;
	wire [4-1:0] node23528;
	wire [4-1:0] node23533;
	wire [4-1:0] node23534;
	wire [4-1:0] node23535;
	wire [4-1:0] node23536;
	wire [4-1:0] node23538;
	wire [4-1:0] node23541;
	wire [4-1:0] node23543;
	wire [4-1:0] node23546;
	wire [4-1:0] node23547;
	wire [4-1:0] node23549;
	wire [4-1:0] node23552;
	wire [4-1:0] node23554;
	wire [4-1:0] node23557;
	wire [4-1:0] node23558;
	wire [4-1:0] node23560;
	wire [4-1:0] node23563;
	wire [4-1:0] node23564;
	wire [4-1:0] node23568;
	wire [4-1:0] node23569;
	wire [4-1:0] node23570;
	wire [4-1:0] node23571;
	wire [4-1:0] node23573;
	wire [4-1:0] node23576;
	wire [4-1:0] node23577;
	wire [4-1:0] node23578;
	wire [4-1:0] node23582;
	wire [4-1:0] node23583;
	wire [4-1:0] node23586;
	wire [4-1:0] node23589;
	wire [4-1:0] node23590;
	wire [4-1:0] node23591;
	wire [4-1:0] node23594;
	wire [4-1:0] node23596;
	wire [4-1:0] node23599;
	wire [4-1:0] node23600;
	wire [4-1:0] node23601;
	wire [4-1:0] node23605;
	wire [4-1:0] node23606;
	wire [4-1:0] node23609;
	wire [4-1:0] node23612;
	wire [4-1:0] node23613;
	wire [4-1:0] node23614;
	wire [4-1:0] node23615;
	wire [4-1:0] node23616;
	wire [4-1:0] node23620;
	wire [4-1:0] node23623;
	wire [4-1:0] node23624;
	wire [4-1:0] node23625;
	wire [4-1:0] node23628;
	wire [4-1:0] node23631;
	wire [4-1:0] node23634;
	wire [4-1:0] node23635;
	wire [4-1:0] node23636;
	wire [4-1:0] node23637;
	wire [4-1:0] node23640;
	wire [4-1:0] node23643;
	wire [4-1:0] node23644;
	wire [4-1:0] node23648;
	wire [4-1:0] node23651;
	wire [4-1:0] node23652;
	wire [4-1:0] node23653;
	wire [4-1:0] node23654;
	wire [4-1:0] node23655;
	wire [4-1:0] node23656;
	wire [4-1:0] node23658;
	wire [4-1:0] node23661;
	wire [4-1:0] node23663;
	wire [4-1:0] node23666;
	wire [4-1:0] node23667;
	wire [4-1:0] node23669;
	wire [4-1:0] node23672;
	wire [4-1:0] node23673;
	wire [4-1:0] node23677;
	wire [4-1:0] node23678;
	wire [4-1:0] node23679;
	wire [4-1:0] node23681;
	wire [4-1:0] node23684;
	wire [4-1:0] node23685;
	wire [4-1:0] node23689;
	wire [4-1:0] node23690;
	wire [4-1:0] node23691;
	wire [4-1:0] node23695;
	wire [4-1:0] node23696;
	wire [4-1:0] node23700;
	wire [4-1:0] node23701;
	wire [4-1:0] node23702;
	wire [4-1:0] node23703;
	wire [4-1:0] node23705;
	wire [4-1:0] node23708;
	wire [4-1:0] node23710;
	wire [4-1:0] node23713;
	wire [4-1:0] node23714;
	wire [4-1:0] node23715;
	wire [4-1:0] node23719;
	wire [4-1:0] node23720;
	wire [4-1:0] node23724;
	wire [4-1:0] node23725;
	wire [4-1:0] node23727;
	wire [4-1:0] node23730;
	wire [4-1:0] node23731;
	wire [4-1:0] node23735;
	wire [4-1:0] node23736;
	wire [4-1:0] node23737;
	wire [4-1:0] node23738;
	wire [4-1:0] node23739;
	wire [4-1:0] node23742;
	wire [4-1:0] node23745;
	wire [4-1:0] node23747;
	wire [4-1:0] node23748;
	wire [4-1:0] node23752;
	wire [4-1:0] node23753;
	wire [4-1:0] node23754;
	wire [4-1:0] node23756;
	wire [4-1:0] node23759;
	wire [4-1:0] node23762;
	wire [4-1:0] node23763;
	wire [4-1:0] node23764;
	wire [4-1:0] node23767;
	wire [4-1:0] node23770;
	wire [4-1:0] node23773;
	wire [4-1:0] node23774;
	wire [4-1:0] node23775;
	wire [4-1:0] node23776;
	wire [4-1:0] node23779;
	wire [4-1:0] node23780;
	wire [4-1:0] node23783;
	wire [4-1:0] node23786;
	wire [4-1:0] node23787;
	wire [4-1:0] node23789;
	wire [4-1:0] node23792;
	wire [4-1:0] node23793;
	wire [4-1:0] node23797;
	wire [4-1:0] node23798;
	wire [4-1:0] node23799;
	wire [4-1:0] node23800;
	wire [4-1:0] node23804;
	wire [4-1:0] node23805;
	wire [4-1:0] node23808;
	wire [4-1:0] node23811;
	wire [4-1:0] node23812;
	wire [4-1:0] node23815;
	wire [4-1:0] node23818;
	wire [4-1:0] node23819;
	wire [4-1:0] node23820;
	wire [4-1:0] node23821;
	wire [4-1:0] node23822;
	wire [4-1:0] node23823;
	wire [4-1:0] node23824;
	wire [4-1:0] node23825;
	wire [4-1:0] node23828;
	wire [4-1:0] node23831;
	wire [4-1:0] node23832;
	wire [4-1:0] node23835;
	wire [4-1:0] node23838;
	wire [4-1:0] node23839;
	wire [4-1:0] node23840;
	wire [4-1:0] node23843;
	wire [4-1:0] node23846;
	wire [4-1:0] node23847;
	wire [4-1:0] node23851;
	wire [4-1:0] node23852;
	wire [4-1:0] node23853;
	wire [4-1:0] node23854;
	wire [4-1:0] node23857;
	wire [4-1:0] node23860;
	wire [4-1:0] node23861;
	wire [4-1:0] node23864;
	wire [4-1:0] node23867;
	wire [4-1:0] node23868;
	wire [4-1:0] node23869;
	wire [4-1:0] node23872;
	wire [4-1:0] node23875;
	wire [4-1:0] node23878;
	wire [4-1:0] node23879;
	wire [4-1:0] node23880;
	wire [4-1:0] node23881;
	wire [4-1:0] node23882;
	wire [4-1:0] node23885;
	wire [4-1:0] node23888;
	wire [4-1:0] node23889;
	wire [4-1:0] node23892;
	wire [4-1:0] node23895;
	wire [4-1:0] node23896;
	wire [4-1:0] node23897;
	wire [4-1:0] node23901;
	wire [4-1:0] node23902;
	wire [4-1:0] node23906;
	wire [4-1:0] node23907;
	wire [4-1:0] node23908;
	wire [4-1:0] node23909;
	wire [4-1:0] node23912;
	wire [4-1:0] node23915;
	wire [4-1:0] node23916;
	wire [4-1:0] node23920;
	wire [4-1:0] node23921;
	wire [4-1:0] node23922;
	wire [4-1:0] node23925;
	wire [4-1:0] node23928;
	wire [4-1:0] node23929;
	wire [4-1:0] node23933;
	wire [4-1:0] node23934;
	wire [4-1:0] node23935;
	wire [4-1:0] node23936;
	wire [4-1:0] node23937;
	wire [4-1:0] node23938;
	wire [4-1:0] node23941;
	wire [4-1:0] node23944;
	wire [4-1:0] node23945;
	wire [4-1:0] node23949;
	wire [4-1:0] node23950;
	wire [4-1:0] node23953;
	wire [4-1:0] node23956;
	wire [4-1:0] node23957;
	wire [4-1:0] node23958;
	wire [4-1:0] node23959;
	wire [4-1:0] node23962;
	wire [4-1:0] node23965;
	wire [4-1:0] node23966;
	wire [4-1:0] node23969;
	wire [4-1:0] node23972;
	wire [4-1:0] node23973;
	wire [4-1:0] node23974;
	wire [4-1:0] node23978;
	wire [4-1:0] node23979;
	wire [4-1:0] node23983;
	wire [4-1:0] node23984;
	wire [4-1:0] node23985;
	wire [4-1:0] node23986;
	wire [4-1:0] node23987;
	wire [4-1:0] node23990;
	wire [4-1:0] node23993;
	wire [4-1:0] node23995;
	wire [4-1:0] node23998;
	wire [4-1:0] node23999;
	wire [4-1:0] node24000;
	wire [4-1:0] node24003;
	wire [4-1:0] node24006;
	wire [4-1:0] node24007;
	wire [4-1:0] node24011;
	wire [4-1:0] node24012;
	wire [4-1:0] node24013;
	wire [4-1:0] node24014;
	wire [4-1:0] node24017;
	wire [4-1:0] node24020;
	wire [4-1:0] node24021;
	wire [4-1:0] node24024;
	wire [4-1:0] node24027;
	wire [4-1:0] node24028;
	wire [4-1:0] node24029;
	wire [4-1:0] node24032;
	wire [4-1:0] node24035;
	wire [4-1:0] node24036;
	wire [4-1:0] node24040;
	wire [4-1:0] node24041;
	wire [4-1:0] node24042;
	wire [4-1:0] node24043;
	wire [4-1:0] node24044;
	wire [4-1:0] node24045;
	wire [4-1:0] node24048;
	wire [4-1:0] node24051;
	wire [4-1:0] node24052;
	wire [4-1:0] node24053;
	wire [4-1:0] node24056;
	wire [4-1:0] node24059;
	wire [4-1:0] node24060;
	wire [4-1:0] node24063;
	wire [4-1:0] node24066;
	wire [4-1:0] node24067;
	wire [4-1:0] node24068;
	wire [4-1:0] node24069;
	wire [4-1:0] node24070;
	wire [4-1:0] node24074;
	wire [4-1:0] node24076;
	wire [4-1:0] node24079;
	wire [4-1:0] node24080;
	wire [4-1:0] node24083;
	wire [4-1:0] node24086;
	wire [4-1:0] node24087;
	wire [4-1:0] node24088;
	wire [4-1:0] node24091;
	wire [4-1:0] node24094;
	wire [4-1:0] node24096;
	wire [4-1:0] node24099;
	wire [4-1:0] node24100;
	wire [4-1:0] node24101;
	wire [4-1:0] node24102;
	wire [4-1:0] node24103;
	wire [4-1:0] node24106;
	wire [4-1:0] node24109;
	wire [4-1:0] node24111;
	wire [4-1:0] node24114;
	wire [4-1:0] node24115;
	wire [4-1:0] node24116;
	wire [4-1:0] node24119;
	wire [4-1:0] node24122;
	wire [4-1:0] node24123;
	wire [4-1:0] node24124;
	wire [4-1:0] node24128;
	wire [4-1:0] node24131;
	wire [4-1:0] node24132;
	wire [4-1:0] node24133;
	wire [4-1:0] node24134;
	wire [4-1:0] node24135;
	wire [4-1:0] node24138;
	wire [4-1:0] node24141;
	wire [4-1:0] node24142;
	wire [4-1:0] node24145;
	wire [4-1:0] node24148;
	wire [4-1:0] node24149;
	wire [4-1:0] node24150;
	wire [4-1:0] node24153;
	wire [4-1:0] node24156;
	wire [4-1:0] node24157;
	wire [4-1:0] node24161;
	wire [4-1:0] node24162;
	wire [4-1:0] node24165;
	wire [4-1:0] node24168;
	wire [4-1:0] node24169;
	wire [4-1:0] node24170;
	wire [4-1:0] node24171;
	wire [4-1:0] node24172;
	wire [4-1:0] node24175;
	wire [4-1:0] node24178;
	wire [4-1:0] node24179;
	wire [4-1:0] node24180;
	wire [4-1:0] node24181;
	wire [4-1:0] node24185;
	wire [4-1:0] node24187;
	wire [4-1:0] node24191;
	wire [4-1:0] node24192;
	wire [4-1:0] node24193;
	wire [4-1:0] node24195;
	wire [4-1:0] node24198;
	wire [4-1:0] node24200;
	wire [4-1:0] node24203;
	wire [4-1:0] node24204;
	wire [4-1:0] node24205;
	wire [4-1:0] node24208;
	wire [4-1:0] node24211;
	wire [4-1:0] node24212;
	wire [4-1:0] node24215;
	wire [4-1:0] node24218;
	wire [4-1:0] node24219;
	wire [4-1:0] node24220;
	wire [4-1:0] node24221;
	wire [4-1:0] node24222;
	wire [4-1:0] node24225;
	wire [4-1:0] node24228;
	wire [4-1:0] node24229;
	wire [4-1:0] node24232;
	wire [4-1:0] node24235;
	wire [4-1:0] node24236;
	wire [4-1:0] node24239;
	wire [4-1:0] node24242;
	wire [4-1:0] node24243;
	wire [4-1:0] node24244;
	wire [4-1:0] node24245;
	wire [4-1:0] node24248;
	wire [4-1:0] node24251;
	wire [4-1:0] node24252;
	wire [4-1:0] node24255;
	wire [4-1:0] node24258;
	wire [4-1:0] node24259;
	wire [4-1:0] node24260;
	wire [4-1:0] node24263;
	wire [4-1:0] node24266;
	wire [4-1:0] node24267;
	wire [4-1:0] node24270;
	wire [4-1:0] node24273;
	wire [4-1:0] node24274;
	wire [4-1:0] node24275;
	wire [4-1:0] node24276;
	wire [4-1:0] node24277;
	wire [4-1:0] node24278;
	wire [4-1:0] node24279;
	wire [4-1:0] node24280;
	wire [4-1:0] node24281;
	wire [4-1:0] node24282;
	wire [4-1:0] node24285;
	wire [4-1:0] node24286;
	wire [4-1:0] node24289;
	wire [4-1:0] node24290;
	wire [4-1:0] node24293;
	wire [4-1:0] node24296;
	wire [4-1:0] node24297;
	wire [4-1:0] node24298;
	wire [4-1:0] node24301;
	wire [4-1:0] node24302;
	wire [4-1:0] node24305;
	wire [4-1:0] node24308;
	wire [4-1:0] node24309;
	wire [4-1:0] node24310;
	wire [4-1:0] node24313;
	wire [4-1:0] node24316;
	wire [4-1:0] node24317;
	wire [4-1:0] node24320;
	wire [4-1:0] node24323;
	wire [4-1:0] node24324;
	wire [4-1:0] node24325;
	wire [4-1:0] node24328;
	wire [4-1:0] node24329;
	wire [4-1:0] node24332;
	wire [4-1:0] node24333;
	wire [4-1:0] node24337;
	wire [4-1:0] node24338;
	wire [4-1:0] node24339;
	wire [4-1:0] node24342;
	wire [4-1:0] node24343;
	wire [4-1:0] node24346;
	wire [4-1:0] node24349;
	wire [4-1:0] node24350;
	wire [4-1:0] node24353;
	wire [4-1:0] node24354;
	wire [4-1:0] node24357;
	wire [4-1:0] node24360;
	wire [4-1:0] node24361;
	wire [4-1:0] node24362;
	wire [4-1:0] node24363;
	wire [4-1:0] node24366;
	wire [4-1:0] node24367;
	wire [4-1:0] node24370;
	wire [4-1:0] node24371;
	wire [4-1:0] node24372;
	wire [4-1:0] node24375;
	wire [4-1:0] node24378;
	wire [4-1:0] node24379;
	wire [4-1:0] node24383;
	wire [4-1:0] node24384;
	wire [4-1:0] node24385;
	wire [4-1:0] node24388;
	wire [4-1:0] node24389;
	wire [4-1:0] node24392;
	wire [4-1:0] node24395;
	wire [4-1:0] node24396;
	wire [4-1:0] node24399;
	wire [4-1:0] node24400;
	wire [4-1:0] node24404;
	wire [4-1:0] node24405;
	wire [4-1:0] node24406;
	wire [4-1:0] node24408;
	wire [4-1:0] node24411;
	wire [4-1:0] node24413;
	wire [4-1:0] node24416;
	wire [4-1:0] node24417;
	wire [4-1:0] node24418;
	wire [4-1:0] node24419;
	wire [4-1:0] node24423;
	wire [4-1:0] node24425;
	wire [4-1:0] node24428;
	wire [4-1:0] node24429;
	wire [4-1:0] node24430;
	wire [4-1:0] node24434;
	wire [4-1:0] node24435;
	wire [4-1:0] node24439;
	wire [4-1:0] node24440;
	wire [4-1:0] node24441;
	wire [4-1:0] node24442;
	wire [4-1:0] node24443;
	wire [4-1:0] node24444;
	wire [4-1:0] node24445;
	wire [4-1:0] node24446;
	wire [4-1:0] node24449;
	wire [4-1:0] node24452;
	wire [4-1:0] node24453;
	wire [4-1:0] node24456;
	wire [4-1:0] node24459;
	wire [4-1:0] node24460;
	wire [4-1:0] node24461;
	wire [4-1:0] node24464;
	wire [4-1:0] node24467;
	wire [4-1:0] node24469;
	wire [4-1:0] node24472;
	wire [4-1:0] node24473;
	wire [4-1:0] node24474;
	wire [4-1:0] node24477;
	wire [4-1:0] node24479;
	wire [4-1:0] node24482;
	wire [4-1:0] node24483;
	wire [4-1:0] node24484;
	wire [4-1:0] node24487;
	wire [4-1:0] node24490;
	wire [4-1:0] node24491;
	wire [4-1:0] node24494;
	wire [4-1:0] node24497;
	wire [4-1:0] node24498;
	wire [4-1:0] node24499;
	wire [4-1:0] node24500;
	wire [4-1:0] node24503;
	wire [4-1:0] node24505;
	wire [4-1:0] node24508;
	wire [4-1:0] node24510;
	wire [4-1:0] node24513;
	wire [4-1:0] node24514;
	wire [4-1:0] node24515;
	wire [4-1:0] node24516;
	wire [4-1:0] node24519;
	wire [4-1:0] node24522;
	wire [4-1:0] node24523;
	wire [4-1:0] node24526;
	wire [4-1:0] node24529;
	wire [4-1:0] node24530;
	wire [4-1:0] node24531;
	wire [4-1:0] node24534;
	wire [4-1:0] node24537;
	wire [4-1:0] node24538;
	wire [4-1:0] node24541;
	wire [4-1:0] node24544;
	wire [4-1:0] node24545;
	wire [4-1:0] node24546;
	wire [4-1:0] node24547;
	wire [4-1:0] node24548;
	wire [4-1:0] node24550;
	wire [4-1:0] node24554;
	wire [4-1:0] node24556;
	wire [4-1:0] node24557;
	wire [4-1:0] node24561;
	wire [4-1:0] node24562;
	wire [4-1:0] node24563;
	wire [4-1:0] node24566;
	wire [4-1:0] node24569;
	wire [4-1:0] node24572;
	wire [4-1:0] node24573;
	wire [4-1:0] node24574;
	wire [4-1:0] node24575;
	wire [4-1:0] node24577;
	wire [4-1:0] node24581;
	wire [4-1:0] node24582;
	wire [4-1:0] node24584;
	wire [4-1:0] node24587;
	wire [4-1:0] node24590;
	wire [4-1:0] node24591;
	wire [4-1:0] node24592;
	wire [4-1:0] node24594;
	wire [4-1:0] node24597;
	wire [4-1:0] node24600;
	wire [4-1:0] node24601;
	wire [4-1:0] node24604;
	wire [4-1:0] node24605;
	wire [4-1:0] node24609;
	wire [4-1:0] node24610;
	wire [4-1:0] node24611;
	wire [4-1:0] node24612;
	wire [4-1:0] node24613;
	wire [4-1:0] node24615;
	wire [4-1:0] node24618;
	wire [4-1:0] node24621;
	wire [4-1:0] node24622;
	wire [4-1:0] node24624;
	wire [4-1:0] node24627;
	wire [4-1:0] node24629;
	wire [4-1:0] node24632;
	wire [4-1:0] node24633;
	wire [4-1:0] node24634;
	wire [4-1:0] node24635;
	wire [4-1:0] node24638;
	wire [4-1:0] node24641;
	wire [4-1:0] node24642;
	wire [4-1:0] node24646;
	wire [4-1:0] node24647;
	wire [4-1:0] node24648;
	wire [4-1:0] node24649;
	wire [4-1:0] node24652;
	wire [4-1:0] node24655;
	wire [4-1:0] node24656;
	wire [4-1:0] node24659;
	wire [4-1:0] node24662;
	wire [4-1:0] node24663;
	wire [4-1:0] node24664;
	wire [4-1:0] node24667;
	wire [4-1:0] node24670;
	wire [4-1:0] node24671;
	wire [4-1:0] node24674;
	wire [4-1:0] node24677;
	wire [4-1:0] node24678;
	wire [4-1:0] node24679;
	wire [4-1:0] node24680;
	wire [4-1:0] node24681;
	wire [4-1:0] node24684;
	wire [4-1:0] node24687;
	wire [4-1:0] node24688;
	wire [4-1:0] node24689;
	wire [4-1:0] node24692;
	wire [4-1:0] node24695;
	wire [4-1:0] node24696;
	wire [4-1:0] node24699;
	wire [4-1:0] node24702;
	wire [4-1:0] node24703;
	wire [4-1:0] node24704;
	wire [4-1:0] node24705;
	wire [4-1:0] node24708;
	wire [4-1:0] node24711;
	wire [4-1:0] node24712;
	wire [4-1:0] node24715;
	wire [4-1:0] node24718;
	wire [4-1:0] node24719;
	wire [4-1:0] node24721;
	wire [4-1:0] node24724;
	wire [4-1:0] node24725;
	wire [4-1:0] node24728;
	wire [4-1:0] node24731;
	wire [4-1:0] node24732;
	wire [4-1:0] node24733;
	wire [4-1:0] node24734;
	wire [4-1:0] node24735;
	wire [4-1:0] node24738;
	wire [4-1:0] node24741;
	wire [4-1:0] node24743;
	wire [4-1:0] node24746;
	wire [4-1:0] node24747;
	wire [4-1:0] node24750;
	wire [4-1:0] node24753;
	wire [4-1:0] node24754;
	wire [4-1:0] node24755;
	wire [4-1:0] node24756;
	wire [4-1:0] node24759;
	wire [4-1:0] node24762;
	wire [4-1:0] node24763;
	wire [4-1:0] node24767;
	wire [4-1:0] node24768;
	wire [4-1:0] node24771;
	wire [4-1:0] node24774;
	wire [4-1:0] node24775;
	wire [4-1:0] node24776;
	wire [4-1:0] node24777;
	wire [4-1:0] node24778;
	wire [4-1:0] node24779;
	wire [4-1:0] node24782;
	wire [4-1:0] node24783;
	wire [4-1:0] node24787;
	wire [4-1:0] node24788;
	wire [4-1:0] node24789;
	wire [4-1:0] node24792;
	wire [4-1:0] node24795;
	wire [4-1:0] node24797;
	wire [4-1:0] node24800;
	wire [4-1:0] node24801;
	wire [4-1:0] node24802;
	wire [4-1:0] node24804;
	wire [4-1:0] node24807;
	wire [4-1:0] node24808;
	wire [4-1:0] node24812;
	wire [4-1:0] node24813;
	wire [4-1:0] node24815;
	wire [4-1:0] node24818;
	wire [4-1:0] node24820;
	wire [4-1:0] node24823;
	wire [4-1:0] node24824;
	wire [4-1:0] node24825;
	wire [4-1:0] node24826;
	wire [4-1:0] node24829;
	wire [4-1:0] node24830;
	wire [4-1:0] node24834;
	wire [4-1:0] node24835;
	wire [4-1:0] node24836;
	wire [4-1:0] node24840;
	wire [4-1:0] node24841;
	wire [4-1:0] node24844;
	wire [4-1:0] node24847;
	wire [4-1:0] node24848;
	wire [4-1:0] node24849;
	wire [4-1:0] node24851;
	wire [4-1:0] node24854;
	wire [4-1:0] node24855;
	wire [4-1:0] node24859;
	wire [4-1:0] node24860;
	wire [4-1:0] node24862;
	wire [4-1:0] node24865;
	wire [4-1:0] node24867;
	wire [4-1:0] node24870;
	wire [4-1:0] node24871;
	wire [4-1:0] node24872;
	wire [4-1:0] node24873;
	wire [4-1:0] node24874;
	wire [4-1:0] node24876;
	wire [4-1:0] node24879;
	wire [4-1:0] node24882;
	wire [4-1:0] node24883;
	wire [4-1:0] node24886;
	wire [4-1:0] node24887;
	wire [4-1:0] node24891;
	wire [4-1:0] node24892;
	wire [4-1:0] node24893;
	wire [4-1:0] node24894;
	wire [4-1:0] node24895;
	wire [4-1:0] node24898;
	wire [4-1:0] node24901;
	wire [4-1:0] node24902;
	wire [4-1:0] node24906;
	wire [4-1:0] node24907;
	wire [4-1:0] node24908;
	wire [4-1:0] node24911;
	wire [4-1:0] node24914;
	wire [4-1:0] node24915;
	wire [4-1:0] node24916;
	wire [4-1:0] node24919;
	wire [4-1:0] node24922;
	wire [4-1:0] node24923;
	wire [4-1:0] node24926;
	wire [4-1:0] node24929;
	wire [4-1:0] node24930;
	wire [4-1:0] node24931;
	wire [4-1:0] node24932;
	wire [4-1:0] node24935;
	wire [4-1:0] node24938;
	wire [4-1:0] node24939;
	wire [4-1:0] node24942;
	wire [4-1:0] node24945;
	wire [4-1:0] node24946;
	wire [4-1:0] node24949;
	wire [4-1:0] node24952;
	wire [4-1:0] node24953;
	wire [4-1:0] node24954;
	wire [4-1:0] node24955;
	wire [4-1:0] node24957;
	wire [4-1:0] node24960;
	wire [4-1:0] node24963;
	wire [4-1:0] node24964;
	wire [4-1:0] node24965;
	wire [4-1:0] node24969;
	wire [4-1:0] node24970;
	wire [4-1:0] node24973;
	wire [4-1:0] node24976;
	wire [4-1:0] node24977;
	wire [4-1:0] node24978;
	wire [4-1:0] node24980;
	wire [4-1:0] node24983;
	wire [4-1:0] node24985;
	wire [4-1:0] node24988;
	wire [4-1:0] node24989;
	wire [4-1:0] node24990;
	wire [4-1:0] node24994;
	wire [4-1:0] node24996;
	wire [4-1:0] node24999;
	wire [4-1:0] node25000;
	wire [4-1:0] node25001;
	wire [4-1:0] node25002;
	wire [4-1:0] node25003;
	wire [4-1:0] node25006;
	wire [4-1:0] node25007;
	wire [4-1:0] node25009;
	wire [4-1:0] node25012;
	wire [4-1:0] node25013;
	wire [4-1:0] node25017;
	wire [4-1:0] node25018;
	wire [4-1:0] node25019;
	wire [4-1:0] node25020;
	wire [4-1:0] node25021;
	wire [4-1:0] node25022;
	wire [4-1:0] node25023;
	wire [4-1:0] node25026;
	wire [4-1:0] node25029;
	wire [4-1:0] node25030;
	wire [4-1:0] node25034;
	wire [4-1:0] node25035;
	wire [4-1:0] node25038;
	wire [4-1:0] node25041;
	wire [4-1:0] node25042;
	wire [4-1:0] node25043;
	wire [4-1:0] node25044;
	wire [4-1:0] node25047;
	wire [4-1:0] node25050;
	wire [4-1:0] node25051;
	wire [4-1:0] node25054;
	wire [4-1:0] node25057;
	wire [4-1:0] node25058;
	wire [4-1:0] node25059;
	wire [4-1:0] node25062;
	wire [4-1:0] node25065;
	wire [4-1:0] node25066;
	wire [4-1:0] node25069;
	wire [4-1:0] node25072;
	wire [4-1:0] node25073;
	wire [4-1:0] node25074;
	wire [4-1:0] node25075;
	wire [4-1:0] node25078;
	wire [4-1:0] node25081;
	wire [4-1:0] node25082;
	wire [4-1:0] node25083;
	wire [4-1:0] node25086;
	wire [4-1:0] node25089;
	wire [4-1:0] node25090;
	wire [4-1:0] node25094;
	wire [4-1:0] node25095;
	wire [4-1:0] node25098;
	wire [4-1:0] node25101;
	wire [4-1:0] node25102;
	wire [4-1:0] node25104;
	wire [4-1:0] node25107;
	wire [4-1:0] node25108;
	wire [4-1:0] node25112;
	wire [4-1:0] node25113;
	wire [4-1:0] node25114;
	wire [4-1:0] node25117;
	wire [4-1:0] node25118;
	wire [4-1:0] node25120;
	wire [4-1:0] node25123;
	wire [4-1:0] node25124;
	wire [4-1:0] node25128;
	wire [4-1:0] node25129;
	wire [4-1:0] node25130;
	wire [4-1:0] node25131;
	wire [4-1:0] node25134;
	wire [4-1:0] node25137;
	wire [4-1:0] node25138;
	wire [4-1:0] node25141;
	wire [4-1:0] node25144;
	wire [4-1:0] node25145;
	wire [4-1:0] node25147;
	wire [4-1:0] node25150;
	wire [4-1:0] node25152;
	wire [4-1:0] node25155;
	wire [4-1:0] node25156;
	wire [4-1:0] node25157;
	wire [4-1:0] node25158;
	wire [4-1:0] node25161;
	wire [4-1:0] node25162;
	wire [4-1:0] node25164;
	wire [4-1:0] node25167;
	wire [4-1:0] node25168;
	wire [4-1:0] node25172;
	wire [4-1:0] node25173;
	wire [4-1:0] node25174;
	wire [4-1:0] node25175;
	wire [4-1:0] node25178;
	wire [4-1:0] node25181;
	wire [4-1:0] node25182;
	wire [4-1:0] node25185;
	wire [4-1:0] node25188;
	wire [4-1:0] node25189;
	wire [4-1:0] node25190;
	wire [4-1:0] node25194;
	wire [4-1:0] node25196;
	wire [4-1:0] node25199;
	wire [4-1:0] node25200;
	wire [4-1:0] node25201;
	wire [4-1:0] node25204;
	wire [4-1:0] node25205;
	wire [4-1:0] node25207;
	wire [4-1:0] node25210;
	wire [4-1:0] node25211;
	wire [4-1:0] node25215;
	wire [4-1:0] node25216;
	wire [4-1:0] node25217;
	wire [4-1:0] node25218;
	wire [4-1:0] node25221;
	wire [4-1:0] node25224;
	wire [4-1:0] node25225;
	wire [4-1:0] node25228;
	wire [4-1:0] node25231;
	wire [4-1:0] node25232;
	wire [4-1:0] node25234;
	wire [4-1:0] node25237;
	wire [4-1:0] node25239;
	wire [4-1:0] node25242;
	wire [4-1:0] node25243;
	wire [4-1:0] node25244;
	wire [4-1:0] node25245;
	wire [4-1:0] node25246;
	wire [4-1:0] node25247;
	wire [4-1:0] node25248;
	wire [4-1:0] node25251;
	wire [4-1:0] node25252;
	wire [4-1:0] node25253;
	wire [4-1:0] node25254;
	wire [4-1:0] node25257;
	wire [4-1:0] node25260;
	wire [4-1:0] node25261;
	wire [4-1:0] node25262;
	wire [4-1:0] node25265;
	wire [4-1:0] node25268;
	wire [4-1:0] node25269;
	wire [4-1:0] node25272;
	wire [4-1:0] node25275;
	wire [4-1:0] node25278;
	wire [4-1:0] node25279;
	wire [4-1:0] node25282;
	wire [4-1:0] node25283;
	wire [4-1:0] node25284;
	wire [4-1:0] node25287;
	wire [4-1:0] node25290;
	wire [4-1:0] node25293;
	wire [4-1:0] node25294;
	wire [4-1:0] node25295;
	wire [4-1:0] node25298;
	wire [4-1:0] node25299;
	wire [4-1:0] node25300;
	wire [4-1:0] node25303;
	wire [4-1:0] node25306;
	wire [4-1:0] node25309;
	wire [4-1:0] node25310;
	wire [4-1:0] node25313;
	wire [4-1:0] node25314;
	wire [4-1:0] node25315;
	wire [4-1:0] node25316;
	wire [4-1:0] node25319;
	wire [4-1:0] node25322;
	wire [4-1:0] node25323;
	wire [4-1:0] node25324;
	wire [4-1:0] node25327;
	wire [4-1:0] node25330;
	wire [4-1:0] node25331;
	wire [4-1:0] node25334;
	wire [4-1:0] node25337;
	wire [4-1:0] node25340;
	wire [4-1:0] node25341;
	wire [4-1:0] node25342;
	wire [4-1:0] node25343;
	wire [4-1:0] node25344;
	wire [4-1:0] node25345;
	wire [4-1:0] node25348;
	wire [4-1:0] node25351;
	wire [4-1:0] node25352;
	wire [4-1:0] node25353;
	wire [4-1:0] node25356;
	wire [4-1:0] node25359;
	wire [4-1:0] node25360;
	wire [4-1:0] node25363;
	wire [4-1:0] node25366;
	wire [4-1:0] node25367;
	wire [4-1:0] node25370;
	wire [4-1:0] node25373;
	wire [4-1:0] node25374;
	wire [4-1:0] node25375;
	wire [4-1:0] node25376;
	wire [4-1:0] node25377;
	wire [4-1:0] node25380;
	wire [4-1:0] node25383;
	wire [4-1:0] node25384;
	wire [4-1:0] node25385;
	wire [4-1:0] node25388;
	wire [4-1:0] node25391;
	wire [4-1:0] node25392;
	wire [4-1:0] node25395;
	wire [4-1:0] node25398;
	wire [4-1:0] node25399;
	wire [4-1:0] node25400;
	wire [4-1:0] node25403;
	wire [4-1:0] node25406;
	wire [4-1:0] node25407;
	wire [4-1:0] node25408;
	wire [4-1:0] node25411;
	wire [4-1:0] node25414;
	wire [4-1:0] node25415;
	wire [4-1:0] node25418;
	wire [4-1:0] node25421;
	wire [4-1:0] node25422;
	wire [4-1:0] node25425;
	wire [4-1:0] node25428;
	wire [4-1:0] node25429;
	wire [4-1:0] node25430;
	wire [4-1:0] node25431;
	wire [4-1:0] node25432;
	wire [4-1:0] node25433;
	wire [4-1:0] node25434;
	wire [4-1:0] node25437;
	wire [4-1:0] node25440;
	wire [4-1:0] node25441;
	wire [4-1:0] node25444;
	wire [4-1:0] node25447;
	wire [4-1:0] node25448;
	wire [4-1:0] node25449;
	wire [4-1:0] node25452;
	wire [4-1:0] node25455;
	wire [4-1:0] node25456;
	wire [4-1:0] node25459;
	wire [4-1:0] node25462;
	wire [4-1:0] node25463;
	wire [4-1:0] node25464;
	wire [4-1:0] node25467;
	wire [4-1:0] node25470;
	wire [4-1:0] node25471;
	wire [4-1:0] node25474;
	wire [4-1:0] node25477;
	wire [4-1:0] node25478;
	wire [4-1:0] node25479;
	wire [4-1:0] node25480;
	wire [4-1:0] node25481;
	wire [4-1:0] node25484;
	wire [4-1:0] node25487;
	wire [4-1:0] node25489;
	wire [4-1:0] node25492;
	wire [4-1:0] node25493;
	wire [4-1:0] node25496;
	wire [4-1:0] node25499;
	wire [4-1:0] node25500;
	wire [4-1:0] node25501;
	wire [4-1:0] node25502;
	wire [4-1:0] node25505;
	wire [4-1:0] node25508;
	wire [4-1:0] node25509;
	wire [4-1:0] node25512;
	wire [4-1:0] node25515;
	wire [4-1:0] node25516;
	wire [4-1:0] node25519;
	wire [4-1:0] node25522;
	wire [4-1:0] node25523;
	wire [4-1:0] node25524;
	wire [4-1:0] node25527;
	wire [4-1:0] node25530;
	wire [4-1:0] node25531;
	wire [4-1:0] node25532;
	wire [4-1:0] node25533;
	wire [4-1:0] node25536;
	wire [4-1:0] node25539;
	wire [4-1:0] node25540;
	wire [4-1:0] node25543;
	wire [4-1:0] node25546;
	wire [4-1:0] node25547;
	wire [4-1:0] node25550;
	wire [4-1:0] node25553;
	wire [4-1:0] node25554;
	wire [4-1:0] node25555;
	wire [4-1:0] node25556;
	wire [4-1:0] node25557;
	wire [4-1:0] node25558;
	wire [4-1:0] node25559;
	wire [4-1:0] node25560;
	wire [4-1:0] node25563;
	wire [4-1:0] node25566;
	wire [4-1:0] node25567;
	wire [4-1:0] node25568;
	wire [4-1:0] node25572;
	wire [4-1:0] node25573;
	wire [4-1:0] node25576;
	wire [4-1:0] node25579;
	wire [4-1:0] node25580;
	wire [4-1:0] node25581;
	wire [4-1:0] node25584;
	wire [4-1:0] node25587;
	wire [4-1:0] node25588;
	wire [4-1:0] node25591;
	wire [4-1:0] node25594;
	wire [4-1:0] node25595;
	wire [4-1:0] node25596;
	wire [4-1:0] node25599;
	wire [4-1:0] node25602;
	wire [4-1:0] node25603;
	wire [4-1:0] node25606;
	wire [4-1:0] node25609;
	wire [4-1:0] node25610;
	wire [4-1:0] node25611;
	wire [4-1:0] node25612;
	wire [4-1:0] node25616;
	wire [4-1:0] node25617;
	wire [4-1:0] node25621;
	wire [4-1:0] node25622;
	wire [4-1:0] node25623;
	wire [4-1:0] node25627;
	wire [4-1:0] node25628;
	wire [4-1:0] node25632;
	wire [4-1:0] node25633;
	wire [4-1:0] node25634;
	wire [4-1:0] node25635;
	wire [4-1:0] node25636;
	wire [4-1:0] node25639;
	wire [4-1:0] node25642;
	wire [4-1:0] node25643;
	wire [4-1:0] node25646;
	wire [4-1:0] node25649;
	wire [4-1:0] node25650;
	wire [4-1:0] node25651;
	wire [4-1:0] node25652;
	wire [4-1:0] node25653;
	wire [4-1:0] node25656;
	wire [4-1:0] node25660;
	wire [4-1:0] node25661;
	wire [4-1:0] node25664;
	wire [4-1:0] node25667;
	wire [4-1:0] node25668;
	wire [4-1:0] node25669;
	wire [4-1:0] node25673;
	wire [4-1:0] node25674;
	wire [4-1:0] node25675;
	wire [4-1:0] node25678;
	wire [4-1:0] node25681;
	wire [4-1:0] node25682;
	wire [4-1:0] node25685;
	wire [4-1:0] node25688;
	wire [4-1:0] node25689;
	wire [4-1:0] node25690;
	wire [4-1:0] node25693;
	wire [4-1:0] node25696;
	wire [4-1:0] node25697;
	wire [4-1:0] node25698;
	wire [4-1:0] node25699;
	wire [4-1:0] node25700;
	wire [4-1:0] node25703;
	wire [4-1:0] node25706;
	wire [4-1:0] node25707;
	wire [4-1:0] node25710;
	wire [4-1:0] node25713;
	wire [4-1:0] node25714;
	wire [4-1:0] node25717;
	wire [4-1:0] node25720;
	wire [4-1:0] node25721;
	wire [4-1:0] node25722;
	wire [4-1:0] node25725;
	wire [4-1:0] node25728;
	wire [4-1:0] node25729;
	wire [4-1:0] node25732;
	wire [4-1:0] node25735;
	wire [4-1:0] node25736;
	wire [4-1:0] node25737;
	wire [4-1:0] node25738;
	wire [4-1:0] node25739;
	wire [4-1:0] node25740;
	wire [4-1:0] node25741;
	wire [4-1:0] node25742;
	wire [4-1:0] node25745;
	wire [4-1:0] node25749;
	wire [4-1:0] node25750;
	wire [4-1:0] node25753;
	wire [4-1:0] node25756;
	wire [4-1:0] node25757;
	wire [4-1:0] node25760;
	wire [4-1:0] node25763;
	wire [4-1:0] node25764;
	wire [4-1:0] node25767;
	wire [4-1:0] node25770;
	wire [4-1:0] node25771;
	wire [4-1:0] node25772;
	wire [4-1:0] node25773;
	wire [4-1:0] node25777;
	wire [4-1:0] node25778;
	wire [4-1:0] node25782;
	wire [4-1:0] node25783;
	wire [4-1:0] node25785;
	wire [4-1:0] node25788;
	wire [4-1:0] node25789;
	wire [4-1:0] node25793;
	wire [4-1:0] node25794;
	wire [4-1:0] node25795;
	wire [4-1:0] node25796;
	wire [4-1:0] node25797;
	wire [4-1:0] node25798;
	wire [4-1:0] node25801;
	wire [4-1:0] node25804;
	wire [4-1:0] node25805;
	wire [4-1:0] node25806;
	wire [4-1:0] node25809;
	wire [4-1:0] node25812;
	wire [4-1:0] node25813;
	wire [4-1:0] node25816;
	wire [4-1:0] node25819;
	wire [4-1:0] node25820;
	wire [4-1:0] node25822;
	wire [4-1:0] node25823;
	wire [4-1:0] node25826;
	wire [4-1:0] node25829;
	wire [4-1:0] node25830;
	wire [4-1:0] node25833;
	wire [4-1:0] node25836;
	wire [4-1:0] node25837;
	wire [4-1:0] node25840;
	wire [4-1:0] node25843;
	wire [4-1:0] node25844;
	wire [4-1:0] node25845;
	wire [4-1:0] node25848;
	wire [4-1:0] node25851;
	wire [4-1:0] node25852;
	wire [4-1:0] node25853;
	wire [4-1:0] node25854;
	wire [4-1:0] node25856;
	wire [4-1:0] node25859;
	wire [4-1:0] node25860;
	wire [4-1:0] node25863;
	wire [4-1:0] node25866;
	wire [4-1:0] node25867;
	wire [4-1:0] node25868;
	wire [4-1:0] node25871;
	wire [4-1:0] node25874;
	wire [4-1:0] node25875;
	wire [4-1:0] node25878;
	wire [4-1:0] node25881;
	wire [4-1:0] node25882;
	wire [4-1:0] node25883;
	wire [4-1:0] node25886;
	wire [4-1:0] node25889;
	wire [4-1:0] node25890;
	wire [4-1:0] node25894;
	wire [4-1:0] node25895;
	wire [4-1:0] node25896;
	wire [4-1:0] node25897;
	wire [4-1:0] node25898;
	wire [4-1:0] node25899;
	wire [4-1:0] node25900;
	wire [4-1:0] node25901;
	wire [4-1:0] node25903;
	wire [4-1:0] node25906;
	wire [4-1:0] node25907;
	wire [4-1:0] node25910;
	wire [4-1:0] node25913;
	wire [4-1:0] node25914;
	wire [4-1:0] node25916;
	wire [4-1:0] node25919;
	wire [4-1:0] node25920;
	wire [4-1:0] node25923;
	wire [4-1:0] node25926;
	wire [4-1:0] node25927;
	wire [4-1:0] node25928;
	wire [4-1:0] node25930;
	wire [4-1:0] node25933;
	wire [4-1:0] node25936;
	wire [4-1:0] node25937;
	wire [4-1:0] node25940;
	wire [4-1:0] node25941;
	wire [4-1:0] node25942;
	wire [4-1:0] node25945;
	wire [4-1:0] node25948;
	wire [4-1:0] node25949;
	wire [4-1:0] node25952;
	wire [4-1:0] node25955;
	wire [4-1:0] node25956;
	wire [4-1:0] node25957;
	wire [4-1:0] node25958;
	wire [4-1:0] node25959;
	wire [4-1:0] node25963;
	wire [4-1:0] node25964;
	wire [4-1:0] node25965;
	wire [4-1:0] node25968;
	wire [4-1:0] node25971;
	wire [4-1:0] node25972;
	wire [4-1:0] node25975;
	wire [4-1:0] node25978;
	wire [4-1:0] node25979;
	wire [4-1:0] node25980;
	wire [4-1:0] node25983;
	wire [4-1:0] node25986;
	wire [4-1:0] node25987;
	wire [4-1:0] node25990;
	wire [4-1:0] node25993;
	wire [4-1:0] node25994;
	wire [4-1:0] node25995;
	wire [4-1:0] node25996;
	wire [4-1:0] node25999;
	wire [4-1:0] node26002;
	wire [4-1:0] node26005;
	wire [4-1:0] node26006;
	wire [4-1:0] node26007;
	wire [4-1:0] node26010;
	wire [4-1:0] node26013;
	wire [4-1:0] node26014;
	wire [4-1:0] node26017;
	wire [4-1:0] node26020;
	wire [4-1:0] node26021;
	wire [4-1:0] node26022;
	wire [4-1:0] node26023;
	wire [4-1:0] node26024;
	wire [4-1:0] node26026;
	wire [4-1:0] node26029;
	wire [4-1:0] node26031;
	wire [4-1:0] node26034;
	wire [4-1:0] node26035;
	wire [4-1:0] node26037;
	wire [4-1:0] node26040;
	wire [4-1:0] node26041;
	wire [4-1:0] node26045;
	wire [4-1:0] node26046;
	wire [4-1:0] node26047;
	wire [4-1:0] node26048;
	wire [4-1:0] node26051;
	wire [4-1:0] node26054;
	wire [4-1:0] node26055;
	wire [4-1:0] node26058;
	wire [4-1:0] node26061;
	wire [4-1:0] node26062;
	wire [4-1:0] node26063;
	wire [4-1:0] node26066;
	wire [4-1:0] node26069;
	wire [4-1:0] node26070;
	wire [4-1:0] node26073;
	wire [4-1:0] node26076;
	wire [4-1:0] node26077;
	wire [4-1:0] node26078;
	wire [4-1:0] node26079;
	wire [4-1:0] node26081;
	wire [4-1:0] node26084;
	wire [4-1:0] node26085;
	wire [4-1:0] node26089;
	wire [4-1:0] node26090;
	wire [4-1:0] node26091;
	wire [4-1:0] node26094;
	wire [4-1:0] node26097;
	wire [4-1:0] node26098;
	wire [4-1:0] node26101;
	wire [4-1:0] node26104;
	wire [4-1:0] node26105;
	wire [4-1:0] node26106;
	wire [4-1:0] node26107;
	wire [4-1:0] node26110;
	wire [4-1:0] node26113;
	wire [4-1:0] node26114;
	wire [4-1:0] node26115;
	wire [4-1:0] node26118;
	wire [4-1:0] node26121;
	wire [4-1:0] node26123;
	wire [4-1:0] node26126;
	wire [4-1:0] node26127;
	wire [4-1:0] node26128;
	wire [4-1:0] node26131;
	wire [4-1:0] node26134;
	wire [4-1:0] node26135;
	wire [4-1:0] node26138;
	wire [4-1:0] node26141;
	wire [4-1:0] node26142;
	wire [4-1:0] node26143;
	wire [4-1:0] node26144;
	wire [4-1:0] node26145;
	wire [4-1:0] node26146;
	wire [4-1:0] node26147;
	wire [4-1:0] node26149;
	wire [4-1:0] node26152;
	wire [4-1:0] node26153;
	wire [4-1:0] node26156;
	wire [4-1:0] node26159;
	wire [4-1:0] node26160;
	wire [4-1:0] node26163;
	wire [4-1:0] node26164;
	wire [4-1:0] node26167;
	wire [4-1:0] node26170;
	wire [4-1:0] node26171;
	wire [4-1:0] node26172;
	wire [4-1:0] node26173;
	wire [4-1:0] node26178;
	wire [4-1:0] node26180;
	wire [4-1:0] node26183;
	wire [4-1:0] node26184;
	wire [4-1:0] node26185;
	wire [4-1:0] node26186;
	wire [4-1:0] node26188;
	wire [4-1:0] node26191;
	wire [4-1:0] node26192;
	wire [4-1:0] node26195;
	wire [4-1:0] node26198;
	wire [4-1:0] node26199;
	wire [4-1:0] node26201;
	wire [4-1:0] node26204;
	wire [4-1:0] node26205;
	wire [4-1:0] node26209;
	wire [4-1:0] node26210;
	wire [4-1:0] node26211;
	wire [4-1:0] node26214;
	wire [4-1:0] node26215;
	wire [4-1:0] node26218;
	wire [4-1:0] node26221;
	wire [4-1:0] node26222;
	wire [4-1:0] node26224;
	wire [4-1:0] node26227;
	wire [4-1:0] node26228;
	wire [4-1:0] node26231;
	wire [4-1:0] node26234;
	wire [4-1:0] node26235;
	wire [4-1:0] node26236;
	wire [4-1:0] node26237;
	wire [4-1:0] node26238;
	wire [4-1:0] node26240;
	wire [4-1:0] node26243;
	wire [4-1:0] node26244;
	wire [4-1:0] node26247;
	wire [4-1:0] node26250;
	wire [4-1:0] node26251;
	wire [4-1:0] node26252;
	wire [4-1:0] node26256;
	wire [4-1:0] node26259;
	wire [4-1:0] node26260;
	wire [4-1:0] node26261;
	wire [4-1:0] node26264;
	wire [4-1:0] node26265;
	wire [4-1:0] node26269;
	wire [4-1:0] node26270;
	wire [4-1:0] node26271;
	wire [4-1:0] node26275;
	wire [4-1:0] node26276;
	wire [4-1:0] node26280;
	wire [4-1:0] node26281;
	wire [4-1:0] node26282;
	wire [4-1:0] node26283;
	wire [4-1:0] node26284;
	wire [4-1:0] node26287;
	wire [4-1:0] node26290;
	wire [4-1:0] node26291;
	wire [4-1:0] node26294;
	wire [4-1:0] node26297;
	wire [4-1:0] node26298;
	wire [4-1:0] node26301;
	wire [4-1:0] node26304;
	wire [4-1:0] node26305;
	wire [4-1:0] node26306;
	wire [4-1:0] node26307;
	wire [4-1:0] node26311;
	wire [4-1:0] node26314;
	wire [4-1:0] node26315;
	wire [4-1:0] node26316;
	wire [4-1:0] node26320;
	wire [4-1:0] node26321;
	wire [4-1:0] node26325;
	wire [4-1:0] node26326;
	wire [4-1:0] node26327;
	wire [4-1:0] node26328;
	wire [4-1:0] node26329;
	wire [4-1:0] node26330;
	wire [4-1:0] node26332;
	wire [4-1:0] node26335;
	wire [4-1:0] node26338;
	wire [4-1:0] node26339;
	wire [4-1:0] node26340;
	wire [4-1:0] node26343;
	wire [4-1:0] node26346;
	wire [4-1:0] node26348;
	wire [4-1:0] node26351;
	wire [4-1:0] node26352;
	wire [4-1:0] node26353;
	wire [4-1:0] node26355;
	wire [4-1:0] node26358;
	wire [4-1:0] node26359;
	wire [4-1:0] node26363;
	wire [4-1:0] node26366;
	wire [4-1:0] node26367;
	wire [4-1:0] node26368;
	wire [4-1:0] node26369;
	wire [4-1:0] node26371;
	wire [4-1:0] node26374;
	wire [4-1:0] node26375;
	wire [4-1:0] node26378;
	wire [4-1:0] node26381;
	wire [4-1:0] node26382;
	wire [4-1:0] node26384;
	wire [4-1:0] node26387;
	wire [4-1:0] node26389;
	wire [4-1:0] node26392;
	wire [4-1:0] node26393;
	wire [4-1:0] node26394;
	wire [4-1:0] node26395;
	wire [4-1:0] node26398;
	wire [4-1:0] node26402;
	wire [4-1:0] node26403;
	wire [4-1:0] node26407;
	wire [4-1:0] node26408;
	wire [4-1:0] node26409;
	wire [4-1:0] node26410;
	wire [4-1:0] node26411;
	wire [4-1:0] node26413;
	wire [4-1:0] node26416;
	wire [4-1:0] node26417;
	wire [4-1:0] node26420;
	wire [4-1:0] node26423;
	wire [4-1:0] node26425;
	wire [4-1:0] node26427;
	wire [4-1:0] node26430;
	wire [4-1:0] node26431;
	wire [4-1:0] node26432;
	wire [4-1:0] node26433;
	wire [4-1:0] node26437;
	wire [4-1:0] node26438;
	wire [4-1:0] node26441;
	wire [4-1:0] node26444;
	wire [4-1:0] node26445;
	wire [4-1:0] node26446;
	wire [4-1:0] node26450;
	wire [4-1:0] node26453;
	wire [4-1:0] node26454;
	wire [4-1:0] node26455;
	wire [4-1:0] node26456;
	wire [4-1:0] node26457;
	wire [4-1:0] node26460;
	wire [4-1:0] node26464;
	wire [4-1:0] node26465;
	wire [4-1:0] node26466;
	wire [4-1:0] node26469;
	wire [4-1:0] node26472;
	wire [4-1:0] node26474;
	wire [4-1:0] node26477;
	wire [4-1:0] node26478;
	wire [4-1:0] node26479;
	wire [4-1:0] node26480;
	wire [4-1:0] node26484;
	wire [4-1:0] node26485;
	wire [4-1:0] node26489;
	wire [4-1:0] node26492;
	wire [4-1:0] node26493;
	wire [4-1:0] node26494;
	wire [4-1:0] node26495;
	wire [4-1:0] node26496;
	wire [4-1:0] node26497;
	wire [4-1:0] node26498;
	wire [4-1:0] node26499;
	wire [4-1:0] node26502;
	wire [4-1:0] node26505;
	wire [4-1:0] node26506;
	wire [4-1:0] node26509;
	wire [4-1:0] node26512;
	wire [4-1:0] node26513;
	wire [4-1:0] node26514;
	wire [4-1:0] node26517;
	wire [4-1:0] node26520;
	wire [4-1:0] node26521;
	wire [4-1:0] node26525;
	wire [4-1:0] node26526;
	wire [4-1:0] node26527;
	wire [4-1:0] node26528;
	wire [4-1:0] node26531;
	wire [4-1:0] node26534;
	wire [4-1:0] node26535;
	wire [4-1:0] node26538;
	wire [4-1:0] node26541;
	wire [4-1:0] node26542;
	wire [4-1:0] node26543;
	wire [4-1:0] node26544;
	wire [4-1:0] node26547;
	wire [4-1:0] node26550;
	wire [4-1:0] node26551;
	wire [4-1:0] node26554;
	wire [4-1:0] node26557;
	wire [4-1:0] node26558;
	wire [4-1:0] node26559;
	wire [4-1:0] node26562;
	wire [4-1:0] node26565;
	wire [4-1:0] node26567;
	wire [4-1:0] node26570;
	wire [4-1:0] node26571;
	wire [4-1:0] node26572;
	wire [4-1:0] node26573;
	wire [4-1:0] node26574;
	wire [4-1:0] node26575;
	wire [4-1:0] node26579;
	wire [4-1:0] node26580;
	wire [4-1:0] node26583;
	wire [4-1:0] node26586;
	wire [4-1:0] node26587;
	wire [4-1:0] node26588;
	wire [4-1:0] node26591;
	wire [4-1:0] node26594;
	wire [4-1:0] node26595;
	wire [4-1:0] node26598;
	wire [4-1:0] node26601;
	wire [4-1:0] node26602;
	wire [4-1:0] node26603;
	wire [4-1:0] node26605;
	wire [4-1:0] node26608;
	wire [4-1:0] node26609;
	wire [4-1:0] node26612;
	wire [4-1:0] node26615;
	wire [4-1:0] node26616;
	wire [4-1:0] node26617;
	wire [4-1:0] node26620;
	wire [4-1:0] node26623;
	wire [4-1:0] node26624;
	wire [4-1:0] node26628;
	wire [4-1:0] node26629;
	wire [4-1:0] node26630;
	wire [4-1:0] node26633;
	wire [4-1:0] node26636;
	wire [4-1:0] node26637;
	wire [4-1:0] node26638;
	wire [4-1:0] node26639;
	wire [4-1:0] node26642;
	wire [4-1:0] node26645;
	wire [4-1:0] node26647;
	wire [4-1:0] node26650;
	wire [4-1:0] node26651;
	wire [4-1:0] node26655;
	wire [4-1:0] node26656;
	wire [4-1:0] node26657;
	wire [4-1:0] node26658;
	wire [4-1:0] node26659;
	wire [4-1:0] node26660;
	wire [4-1:0] node26663;
	wire [4-1:0] node26666;
	wire [4-1:0] node26668;
	wire [4-1:0] node26669;
	wire [4-1:0] node26672;
	wire [4-1:0] node26675;
	wire [4-1:0] node26676;
	wire [4-1:0] node26677;
	wire [4-1:0] node26678;
	wire [4-1:0] node26681;
	wire [4-1:0] node26685;
	wire [4-1:0] node26686;
	wire [4-1:0] node26687;
	wire [4-1:0] node26690;
	wire [4-1:0] node26693;
	wire [4-1:0] node26694;
	wire [4-1:0] node26697;
	wire [4-1:0] node26700;
	wire [4-1:0] node26701;
	wire [4-1:0] node26702;
	wire [4-1:0] node26703;
	wire [4-1:0] node26706;
	wire [4-1:0] node26709;
	wire [4-1:0] node26710;
	wire [4-1:0] node26711;
	wire [4-1:0] node26714;
	wire [4-1:0] node26717;
	wire [4-1:0] node26718;
	wire [4-1:0] node26721;
	wire [4-1:0] node26724;
	wire [4-1:0] node26725;
	wire [4-1:0] node26726;
	wire [4-1:0] node26727;
	wire [4-1:0] node26730;
	wire [4-1:0] node26733;
	wire [4-1:0] node26734;
	wire [4-1:0] node26737;
	wire [4-1:0] node26740;
	wire [4-1:0] node26742;
	wire [4-1:0] node26743;
	wire [4-1:0] node26746;
	wire [4-1:0] node26749;
	wire [4-1:0] node26750;
	wire [4-1:0] node26751;
	wire [4-1:0] node26752;
	wire [4-1:0] node26755;
	wire [4-1:0] node26758;
	wire [4-1:0] node26759;
	wire [4-1:0] node26762;
	wire [4-1:0] node26765;
	wire [4-1:0] node26766;
	wire [4-1:0] node26767;
	wire [4-1:0] node26768;
	wire [4-1:0] node26771;
	wire [4-1:0] node26774;
	wire [4-1:0] node26775;
	wire [4-1:0] node26778;
	wire [4-1:0] node26781;
	wire [4-1:0] node26782;
	wire [4-1:0] node26783;
	wire [4-1:0] node26786;
	wire [4-1:0] node26789;
	wire [4-1:0] node26790;
	wire [4-1:0] node26793;
	wire [4-1:0] node26796;
	wire [4-1:0] node26797;
	wire [4-1:0] node26798;
	wire [4-1:0] node26799;
	wire [4-1:0] node26800;
	wire [4-1:0] node26801;
	wire [4-1:0] node26802;
	wire [4-1:0] node26804;
	wire [4-1:0] node26807;
	wire [4-1:0] node26809;
	wire [4-1:0] node26812;
	wire [4-1:0] node26813;
	wire [4-1:0] node26815;
	wire [4-1:0] node26818;
	wire [4-1:0] node26819;
	wire [4-1:0] node26823;
	wire [4-1:0] node26824;
	wire [4-1:0] node26825;
	wire [4-1:0] node26828;
	wire [4-1:0] node26831;
	wire [4-1:0] node26832;
	wire [4-1:0] node26835;
	wire [4-1:0] node26838;
	wire [4-1:0] node26839;
	wire [4-1:0] node26840;
	wire [4-1:0] node26842;
	wire [4-1:0] node26845;
	wire [4-1:0] node26846;
	wire [4-1:0] node26850;
	wire [4-1:0] node26851;
	wire [4-1:0] node26853;
	wire [4-1:0] node26856;
	wire [4-1:0] node26857;
	wire [4-1:0] node26861;
	wire [4-1:0] node26862;
	wire [4-1:0] node26863;
	wire [4-1:0] node26864;
	wire [4-1:0] node26865;
	wire [4-1:0] node26869;
	wire [4-1:0] node26870;
	wire [4-1:0] node26873;
	wire [4-1:0] node26876;
	wire [4-1:0] node26877;
	wire [4-1:0] node26878;
	wire [4-1:0] node26879;
	wire [4-1:0] node26883;
	wire [4-1:0] node26884;
	wire [4-1:0] node26888;
	wire [4-1:0] node26889;
	wire [4-1:0] node26890;
	wire [4-1:0] node26894;
	wire [4-1:0] node26895;
	wire [4-1:0] node26899;
	wire [4-1:0] node26900;
	wire [4-1:0] node26901;
	wire [4-1:0] node26902;
	wire [4-1:0] node26906;
	wire [4-1:0] node26907;
	wire [4-1:0] node26911;
	wire [4-1:0] node26912;
	wire [4-1:0] node26913;
	wire [4-1:0] node26917;
	wire [4-1:0] node26918;
	wire [4-1:0] node26922;
	wire [4-1:0] node26923;
	wire [4-1:0] node26924;
	wire [4-1:0] node26925;
	wire [4-1:0] node26926;
	wire [4-1:0] node26927;
	wire [4-1:0] node26930;
	wire [4-1:0] node26933;
	wire [4-1:0] node26934;
	wire [4-1:0] node26937;
	wire [4-1:0] node26940;
	wire [4-1:0] node26941;
	wire [4-1:0] node26942;
	wire [4-1:0] node26943;
	wire [4-1:0] node26946;
	wire [4-1:0] node26950;
	wire [4-1:0] node26951;
	wire [4-1:0] node26954;
	wire [4-1:0] node26957;
	wire [4-1:0] node26958;
	wire [4-1:0] node26959;
	wire [4-1:0] node26960;
	wire [4-1:0] node26964;
	wire [4-1:0] node26965;
	wire [4-1:0] node26969;
	wire [4-1:0] node26970;
	wire [4-1:0] node26971;
	wire [4-1:0] node26975;
	wire [4-1:0] node26976;
	wire [4-1:0] node26980;
	wire [4-1:0] node26981;
	wire [4-1:0] node26982;
	wire [4-1:0] node26983;
	wire [4-1:0] node26984;
	wire [4-1:0] node26988;
	wire [4-1:0] node26989;
	wire [4-1:0] node26993;
	wire [4-1:0] node26994;
	wire [4-1:0] node26995;
	wire [4-1:0] node26999;
	wire [4-1:0] node27000;
	wire [4-1:0] node27004;
	wire [4-1:0] node27005;
	wire [4-1:0] node27006;
	wire [4-1:0] node27007;
	wire [4-1:0] node27010;
	wire [4-1:0] node27013;
	wire [4-1:0] node27014;
	wire [4-1:0] node27015;
	wire [4-1:0] node27018;
	wire [4-1:0] node27021;
	wire [4-1:0] node27022;
	wire [4-1:0] node27025;
	wire [4-1:0] node27028;
	wire [4-1:0] node27029;
	wire [4-1:0] node27032;
	wire [4-1:0] node27035;
	wire [4-1:0] node27036;
	wire [4-1:0] node27037;
	wire [4-1:0] node27038;
	wire [4-1:0] node27039;
	wire [4-1:0] node27040;
	wire [4-1:0] node27041;
	wire [4-1:0] node27044;
	wire [4-1:0] node27045;
	wire [4-1:0] node27047;
	wire [4-1:0] node27050;
	wire [4-1:0] node27051;
	wire [4-1:0] node27055;
	wire [4-1:0] node27056;
	wire [4-1:0] node27057;
	wire [4-1:0] node27058;
	wire [4-1:0] node27061;
	wire [4-1:0] node27064;
	wire [4-1:0] node27065;
	wire [4-1:0] node27068;
	wire [4-1:0] node27071;
	wire [4-1:0] node27072;
	wire [4-1:0] node27073;
	wire [4-1:0] node27077;
	wire [4-1:0] node27079;
	wire [4-1:0] node27082;
	wire [4-1:0] node27083;
	wire [4-1:0] node27084;
	wire [4-1:0] node27087;
	wire [4-1:0] node27088;
	wire [4-1:0] node27090;
	wire [4-1:0] node27093;
	wire [4-1:0] node27094;
	wire [4-1:0] node27098;
	wire [4-1:0] node27099;
	wire [4-1:0] node27100;
	wire [4-1:0] node27101;
	wire [4-1:0] node27104;
	wire [4-1:0] node27107;
	wire [4-1:0] node27108;
	wire [4-1:0] node27111;
	wire [4-1:0] node27114;
	wire [4-1:0] node27115;
	wire [4-1:0] node27117;
	wire [4-1:0] node27120;
	wire [4-1:0] node27122;
	wire [4-1:0] node27125;
	wire [4-1:0] node27126;
	wire [4-1:0] node27127;
	wire [4-1:0] node27128;
	wire [4-1:0] node27131;
	wire [4-1:0] node27132;
	wire [4-1:0] node27134;
	wire [4-1:0] node27137;
	wire [4-1:0] node27138;
	wire [4-1:0] node27142;
	wire [4-1:0] node27143;
	wire [4-1:0] node27144;
	wire [4-1:0] node27145;
	wire [4-1:0] node27146;
	wire [4-1:0] node27149;
	wire [4-1:0] node27152;
	wire [4-1:0] node27153;
	wire [4-1:0] node27154;
	wire [4-1:0] node27157;
	wire [4-1:0] node27160;
	wire [4-1:0] node27161;
	wire [4-1:0] node27162;
	wire [4-1:0] node27165;
	wire [4-1:0] node27168;
	wire [4-1:0] node27170;
	wire [4-1:0] node27173;
	wire [4-1:0] node27174;
	wire [4-1:0] node27177;
	wire [4-1:0] node27180;
	wire [4-1:0] node27181;
	wire [4-1:0] node27183;
	wire [4-1:0] node27186;
	wire [4-1:0] node27188;
	wire [4-1:0] node27191;
	wire [4-1:0] node27192;
	wire [4-1:0] node27193;
	wire [4-1:0] node27196;
	wire [4-1:0] node27197;
	wire [4-1:0] node27199;
	wire [4-1:0] node27202;
	wire [4-1:0] node27203;
	wire [4-1:0] node27207;
	wire [4-1:0] node27208;
	wire [4-1:0] node27209;
	wire [4-1:0] node27210;
	wire [4-1:0] node27213;
	wire [4-1:0] node27216;
	wire [4-1:0] node27217;
	wire [4-1:0] node27218;
	wire [4-1:0] node27220;
	wire [4-1:0] node27223;
	wire [4-1:0] node27224;
	wire [4-1:0] node27227;
	wire [4-1:0] node27230;
	wire [4-1:0] node27231;
	wire [4-1:0] node27232;
	wire [4-1:0] node27235;
	wire [4-1:0] node27238;
	wire [4-1:0] node27239;
	wire [4-1:0] node27242;
	wire [4-1:0] node27245;
	wire [4-1:0] node27246;
	wire [4-1:0] node27247;
	wire [4-1:0] node27251;
	wire [4-1:0] node27252;
	wire [4-1:0] node27256;
	wire [4-1:0] node27257;
	wire [4-1:0] node27258;
	wire [4-1:0] node27259;
	wire [4-1:0] node27260;
	wire [4-1:0] node27262;
	wire [4-1:0] node27265;
	wire [4-1:0] node27267;
	wire [4-1:0] node27270;
	wire [4-1:0] node27271;
	wire [4-1:0] node27273;
	wire [4-1:0] node27276;
	wire [4-1:0] node27278;
	wire [4-1:0] node27281;
	wire [4-1:0] node27282;
	wire [4-1:0] node27283;
	wire [4-1:0] node27284;
	wire [4-1:0] node27285;
	wire [4-1:0] node27286;
	wire [4-1:0] node27289;
	wire [4-1:0] node27292;
	wire [4-1:0] node27293;
	wire [4-1:0] node27294;
	wire [4-1:0] node27297;
	wire [4-1:0] node27300;
	wire [4-1:0] node27301;
	wire [4-1:0] node27302;
	wire [4-1:0] node27305;
	wire [4-1:0] node27308;
	wire [4-1:0] node27309;
	wire [4-1:0] node27312;
	wire [4-1:0] node27315;
	wire [4-1:0] node27316;
	wire [4-1:0] node27319;
	wire [4-1:0] node27322;
	wire [4-1:0] node27323;
	wire [4-1:0] node27324;
	wire [4-1:0] node27327;
	wire [4-1:0] node27330;
	wire [4-1:0] node27331;
	wire [4-1:0] node27334;
	wire [4-1:0] node27337;
	wire [4-1:0] node27338;
	wire [4-1:0] node27339;
	wire [4-1:0] node27340;
	wire [4-1:0] node27341;
	wire [4-1:0] node27342;
	wire [4-1:0] node27343;
	wire [4-1:0] node27346;
	wire [4-1:0] node27349;
	wire [4-1:0] node27350;
	wire [4-1:0] node27354;
	wire [4-1:0] node27356;
	wire [4-1:0] node27359;
	wire [4-1:0] node27360;
	wire [4-1:0] node27363;
	wire [4-1:0] node27366;
	wire [4-1:0] node27367;
	wire [4-1:0] node27368;
	wire [4-1:0] node27371;
	wire [4-1:0] node27374;
	wire [4-1:0] node27375;
	wire [4-1:0] node27378;
	wire [4-1:0] node27381;
	wire [4-1:0] node27382;
	wire [4-1:0] node27383;
	wire [4-1:0] node27384;
	wire [4-1:0] node27387;
	wire [4-1:0] node27390;
	wire [4-1:0] node27391;
	wire [4-1:0] node27394;
	wire [4-1:0] node27397;
	wire [4-1:0] node27398;
	wire [4-1:0] node27401;
	wire [4-1:0] node27404;
	wire [4-1:0] node27405;
	wire [4-1:0] node27406;
	wire [4-1:0] node27407;
	wire [4-1:0] node27408;
	wire [4-1:0] node27409;
	wire [4-1:0] node27412;
	wire [4-1:0] node27415;
	wire [4-1:0] node27416;
	wire [4-1:0] node27417;
	wire [4-1:0] node27420;
	wire [4-1:0] node27423;
	wire [4-1:0] node27424;
	wire [4-1:0] node27427;
	wire [4-1:0] node27430;
	wire [4-1:0] node27431;
	wire [4-1:0] node27432;
	wire [4-1:0] node27435;
	wire [4-1:0] node27438;
	wire [4-1:0] node27439;
	wire [4-1:0] node27440;
	wire [4-1:0] node27441;
	wire [4-1:0] node27442;
	wire [4-1:0] node27446;
	wire [4-1:0] node27447;
	wire [4-1:0] node27450;
	wire [4-1:0] node27453;
	wire [4-1:0] node27454;
	wire [4-1:0] node27457;
	wire [4-1:0] node27460;
	wire [4-1:0] node27461;
	wire [4-1:0] node27464;
	wire [4-1:0] node27467;
	wire [4-1:0] node27468;
	wire [4-1:0] node27469;
	wire [4-1:0] node27470;
	wire [4-1:0] node27474;
	wire [4-1:0] node27476;
	wire [4-1:0] node27479;
	wire [4-1:0] node27480;
	wire [4-1:0] node27482;
	wire [4-1:0] node27485;
	wire [4-1:0] node27486;
	wire [4-1:0] node27490;
	wire [4-1:0] node27491;
	wire [4-1:0] node27492;
	wire [4-1:0] node27493;
	wire [4-1:0] node27494;
	wire [4-1:0] node27495;
	wire [4-1:0] node27498;
	wire [4-1:0] node27501;
	wire [4-1:0] node27502;
	wire [4-1:0] node27503;
	wire [4-1:0] node27504;
	wire [4-1:0] node27508;
	wire [4-1:0] node27511;
	wire [4-1:0] node27512;
	wire [4-1:0] node27515;
	wire [4-1:0] node27518;
	wire [4-1:0] node27519;
	wire [4-1:0] node27520;
	wire [4-1:0] node27523;
	wire [4-1:0] node27526;
	wire [4-1:0] node27527;
	wire [4-1:0] node27528;
	wire [4-1:0] node27531;
	wire [4-1:0] node27534;
	wire [4-1:0] node27535;
	wire [4-1:0] node27538;
	wire [4-1:0] node27541;
	wire [4-1:0] node27542;
	wire [4-1:0] node27543;
	wire [4-1:0] node27544;
	wire [4-1:0] node27547;
	wire [4-1:0] node27550;
	wire [4-1:0] node27551;
	wire [4-1:0] node27554;
	wire [4-1:0] node27557;
	wire [4-1:0] node27558;
	wire [4-1:0] node27561;
	wire [4-1:0] node27564;
	wire [4-1:0] node27565;
	wire [4-1:0] node27566;
	wire [4-1:0] node27567;
	wire [4-1:0] node27570;
	wire [4-1:0] node27573;
	wire [4-1:0] node27574;
	wire [4-1:0] node27575;
	wire [4-1:0] node27578;
	wire [4-1:0] node27581;
	wire [4-1:0] node27582;
	wire [4-1:0] node27585;
	wire [4-1:0] node27588;
	wire [4-1:0] node27589;
	wire [4-1:0] node27590;
	wire [4-1:0] node27591;
	wire [4-1:0] node27592;
	wire [4-1:0] node27595;
	wire [4-1:0] node27598;
	wire [4-1:0] node27599;
	wire [4-1:0] node27602;
	wire [4-1:0] node27605;
	wire [4-1:0] node27606;
	wire [4-1:0] node27607;
	wire [4-1:0] node27610;
	wire [4-1:0] node27613;
	wire [4-1:0] node27614;
	wire [4-1:0] node27615;
	wire [4-1:0] node27618;
	wire [4-1:0] node27621;
	wire [4-1:0] node27622;
	wire [4-1:0] node27625;
	wire [4-1:0] node27628;
	wire [4-1:0] node27629;
	wire [4-1:0] node27630;
	wire [4-1:0] node27633;
	wire [4-1:0] node27636;
	wire [4-1:0] node27637;
	wire [4-1:0] node27640;
	wire [4-1:0] node27643;
	wire [4-1:0] node27644;
	wire [4-1:0] node27645;
	wire [4-1:0] node27646;
	wire [4-1:0] node27647;
	wire [4-1:0] node27648;
	wire [4-1:0] node27649;
	wire [4-1:0] node27650;
	wire [4-1:0] node27651;
	wire [4-1:0] node27652;
	wire [4-1:0] node27653;
	wire [4-1:0] node27656;
	wire [4-1:0] node27659;
	wire [4-1:0] node27660;
	wire [4-1:0] node27663;
	wire [4-1:0] node27666;
	wire [4-1:0] node27667;
	wire [4-1:0] node27670;
	wire [4-1:0] node27673;
	wire [4-1:0] node27674;
	wire [4-1:0] node27675;
	wire [4-1:0] node27676;
	wire [4-1:0] node27679;
	wire [4-1:0] node27682;
	wire [4-1:0] node27683;
	wire [4-1:0] node27686;
	wire [4-1:0] node27689;
	wire [4-1:0] node27690;
	wire [4-1:0] node27693;
	wire [4-1:0] node27696;
	wire [4-1:0] node27697;
	wire [4-1:0] node27698;
	wire [4-1:0] node27701;
	wire [4-1:0] node27704;
	wire [4-1:0] node27705;
	wire [4-1:0] node27708;
	wire [4-1:0] node27711;
	wire [4-1:0] node27712;
	wire [4-1:0] node27713;
	wire [4-1:0] node27714;
	wire [4-1:0] node27717;
	wire [4-1:0] node27720;
	wire [4-1:0] node27721;
	wire [4-1:0] node27724;
	wire [4-1:0] node27727;
	wire [4-1:0] node27728;
	wire [4-1:0] node27729;
	wire [4-1:0] node27732;
	wire [4-1:0] node27735;
	wire [4-1:0] node27736;
	wire [4-1:0] node27737;
	wire [4-1:0] node27740;
	wire [4-1:0] node27743;
	wire [4-1:0] node27745;
	wire [4-1:0] node27748;
	wire [4-1:0] node27749;
	wire [4-1:0] node27750;
	wire [4-1:0] node27751;
	wire [4-1:0] node27752;
	wire [4-1:0] node27753;
	wire [4-1:0] node27756;
	wire [4-1:0] node27759;
	wire [4-1:0] node27760;
	wire [4-1:0] node27763;
	wire [4-1:0] node27766;
	wire [4-1:0] node27767;
	wire [4-1:0] node27768;
	wire [4-1:0] node27771;
	wire [4-1:0] node27774;
	wire [4-1:0] node27775;
	wire [4-1:0] node27776;
	wire [4-1:0] node27779;
	wire [4-1:0] node27782;
	wire [4-1:0] node27783;
	wire [4-1:0] node27786;
	wire [4-1:0] node27789;
	wire [4-1:0] node27790;
	wire [4-1:0] node27791;
	wire [4-1:0] node27792;
	wire [4-1:0] node27795;
	wire [4-1:0] node27798;
	wire [4-1:0] node27799;
	wire [4-1:0] node27802;
	wire [4-1:0] node27805;
	wire [4-1:0] node27806;
	wire [4-1:0] node27809;
	wire [4-1:0] node27812;
	wire [4-1:0] node27813;
	wire [4-1:0] node27814;
	wire [4-1:0] node27815;
	wire [4-1:0] node27816;
	wire [4-1:0] node27819;
	wire [4-1:0] node27822;
	wire [4-1:0] node27823;
	wire [4-1:0] node27826;
	wire [4-1:0] node27829;
	wire [4-1:0] node27830;
	wire [4-1:0] node27831;
	wire [4-1:0] node27832;
	wire [4-1:0] node27835;
	wire [4-1:0] node27838;
	wire [4-1:0] node27839;
	wire [4-1:0] node27842;
	wire [4-1:0] node27845;
	wire [4-1:0] node27846;
	wire [4-1:0] node27849;
	wire [4-1:0] node27852;
	wire [4-1:0] node27853;
	wire [4-1:0] node27854;
	wire [4-1:0] node27855;
	wire [4-1:0] node27858;
	wire [4-1:0] node27861;
	wire [4-1:0] node27862;
	wire [4-1:0] node27865;
	wire [4-1:0] node27868;
	wire [4-1:0] node27869;
	wire [4-1:0] node27870;
	wire [4-1:0] node27874;
	wire [4-1:0] node27875;
	wire [4-1:0] node27878;
	wire [4-1:0] node27881;
	wire [4-1:0] node27882;
	wire [4-1:0] node27883;
	wire [4-1:0] node27884;
	wire [4-1:0] node27888;
	wire [4-1:0] node27890;
	wire [4-1:0] node27893;
	wire [4-1:0] node27894;
	wire [4-1:0] node27896;
	wire [4-1:0] node27899;
	wire [4-1:0] node27901;
	wire [4-1:0] node27904;
	wire [4-1:0] node27905;
	wire [4-1:0] node27906;
	wire [4-1:0] node27909;
	wire [4-1:0] node27912;
	wire [4-1:0] node27913;
	wire [4-1:0] node27914;
	wire [4-1:0] node27915;
	wire [4-1:0] node27916;
	wire [4-1:0] node27917;
	wire [4-1:0] node27920;
	wire [4-1:0] node27923;
	wire [4-1:0] node27924;
	wire [4-1:0] node27927;
	wire [4-1:0] node27930;
	wire [4-1:0] node27931;
	wire [4-1:0] node27932;
	wire [4-1:0] node27933;
	wire [4-1:0] node27936;
	wire [4-1:0] node27939;
	wire [4-1:0] node27940;
	wire [4-1:0] node27943;
	wire [4-1:0] node27946;
	wire [4-1:0] node27947;
	wire [4-1:0] node27950;
	wire [4-1:0] node27953;
	wire [4-1:0] node27954;
	wire [4-1:0] node27955;
	wire [4-1:0] node27956;
	wire [4-1:0] node27959;
	wire [4-1:0] node27962;
	wire [4-1:0] node27963;
	wire [4-1:0] node27964;
	wire [4-1:0] node27966;
	wire [4-1:0] node27970;
	wire [4-1:0] node27972;
	wire [4-1:0] node27973;
	wire [4-1:0] node27976;
	wire [4-1:0] node27979;
	wire [4-1:0] node27980;
	wire [4-1:0] node27981;
	wire [4-1:0] node27984;
	wire [4-1:0] node27987;
	wire [4-1:0] node27988;
	wire [4-1:0] node27991;
	wire [4-1:0] node27994;
	wire [4-1:0] node27995;
	wire [4-1:0] node27996;
	wire [4-1:0] node27997;
	wire [4-1:0] node27998;
	wire [4-1:0] node27999;
	wire [4-1:0] node28000;
	wire [4-1:0] node28003;
	wire [4-1:0] node28006;
	wire [4-1:0] node28007;
	wire [4-1:0] node28010;
	wire [4-1:0] node28013;
	wire [4-1:0] node28014;
	wire [4-1:0] node28015;
	wire [4-1:0] node28018;
	wire [4-1:0] node28021;
	wire [4-1:0] node28022;
	wire [4-1:0] node28025;
	wire [4-1:0] node28028;
	wire [4-1:0] node28029;
	wire [4-1:0] node28030;
	wire [4-1:0] node28034;
	wire [4-1:0] node28035;
	wire [4-1:0] node28038;
	wire [4-1:0] node28041;
	wire [4-1:0] node28042;
	wire [4-1:0] node28045;
	wire [4-1:0] node28048;
	wire [4-1:0] node28049;
	wire [4-1:0] node28052;
	wire [4-1:0] node28055;
	wire [4-1:0] node28056;
	wire [4-1:0] node28057;
	wire [4-1:0] node28058;
	wire [4-1:0] node28059;
	wire [4-1:0] node28060;
	wire [4-1:0] node28061;
	wire [4-1:0] node28065;
	wire [4-1:0] node28067;
	wire [4-1:0] node28070;
	wire [4-1:0] node28071;
	wire [4-1:0] node28072;
	wire [4-1:0] node28076;
	wire [4-1:0] node28078;
	wire [4-1:0] node28081;
	wire [4-1:0] node28082;
	wire [4-1:0] node28083;
	wire [4-1:0] node28084;
	wire [4-1:0] node28085;
	wire [4-1:0] node28089;
	wire [4-1:0] node28090;
	wire [4-1:0] node28094;
	wire [4-1:0] node28095;
	wire [4-1:0] node28097;
	wire [4-1:0] node28100;
	wire [4-1:0] node28102;
	wire [4-1:0] node28105;
	wire [4-1:0] node28106;
	wire [4-1:0] node28107;
	wire [4-1:0] node28108;
	wire [4-1:0] node28109;
	wire [4-1:0] node28112;
	wire [4-1:0] node28115;
	wire [4-1:0] node28116;
	wire [4-1:0] node28119;
	wire [4-1:0] node28122;
	wire [4-1:0] node28123;
	wire [4-1:0] node28124;
	wire [4-1:0] node28125;
	wire [4-1:0] node28128;
	wire [4-1:0] node28132;
	wire [4-1:0] node28133;
	wire [4-1:0] node28134;
	wire [4-1:0] node28138;
	wire [4-1:0] node28139;
	wire [4-1:0] node28142;
	wire [4-1:0] node28145;
	wire [4-1:0] node28146;
	wire [4-1:0] node28147;
	wire [4-1:0] node28148;
	wire [4-1:0] node28149;
	wire [4-1:0] node28152;
	wire [4-1:0] node28155;
	wire [4-1:0] node28156;
	wire [4-1:0] node28159;
	wire [4-1:0] node28162;
	wire [4-1:0] node28163;
	wire [4-1:0] node28164;
	wire [4-1:0] node28167;
	wire [4-1:0] node28170;
	wire [4-1:0] node28171;
	wire [4-1:0] node28174;
	wire [4-1:0] node28177;
	wire [4-1:0] node28178;
	wire [4-1:0] node28179;
	wire [4-1:0] node28182;
	wire [4-1:0] node28185;
	wire [4-1:0] node28186;
	wire [4-1:0] node28187;
	wire [4-1:0] node28190;
	wire [4-1:0] node28193;
	wire [4-1:0] node28194;
	wire [4-1:0] node28197;
	wire [4-1:0] node28200;
	wire [4-1:0] node28201;
	wire [4-1:0] node28202;
	wire [4-1:0] node28203;
	wire [4-1:0] node28204;
	wire [4-1:0] node28205;
	wire [4-1:0] node28209;
	wire [4-1:0] node28210;
	wire [4-1:0] node28214;
	wire [4-1:0] node28215;
	wire [4-1:0] node28216;
	wire [4-1:0] node28220;
	wire [4-1:0] node28221;
	wire [4-1:0] node28225;
	wire [4-1:0] node28226;
	wire [4-1:0] node28227;
	wire [4-1:0] node28228;
	wire [4-1:0] node28232;
	wire [4-1:0] node28233;
	wire [4-1:0] node28237;
	wire [4-1:0] node28238;
	wire [4-1:0] node28239;
	wire [4-1:0] node28243;
	wire [4-1:0] node28244;
	wire [4-1:0] node28248;
	wire [4-1:0] node28249;
	wire [4-1:0] node28250;
	wire [4-1:0] node28251;
	wire [4-1:0] node28252;
	wire [4-1:0] node28254;
	wire [4-1:0] node28255;
	wire [4-1:0] node28258;
	wire [4-1:0] node28261;
	wire [4-1:0] node28262;
	wire [4-1:0] node28263;
	wire [4-1:0] node28266;
	wire [4-1:0] node28269;
	wire [4-1:0] node28271;
	wire [4-1:0] node28274;
	wire [4-1:0] node28275;
	wire [4-1:0] node28276;
	wire [4-1:0] node28278;
	wire [4-1:0] node28282;
	wire [4-1:0] node28283;
	wire [4-1:0] node28284;
	wire [4-1:0] node28287;
	wire [4-1:0] node28290;
	wire [4-1:0] node28291;
	wire [4-1:0] node28294;
	wire [4-1:0] node28297;
	wire [4-1:0] node28298;
	wire [4-1:0] node28299;
	wire [4-1:0] node28302;
	wire [4-1:0] node28305;
	wire [4-1:0] node28306;
	wire [4-1:0] node28309;
	wire [4-1:0] node28312;
	wire [4-1:0] node28313;
	wire [4-1:0] node28315;
	wire [4-1:0] node28316;
	wire [4-1:0] node28320;
	wire [4-1:0] node28321;
	wire [4-1:0] node28322;
	wire [4-1:0] node28326;
	wire [4-1:0] node28327;
	wire [4-1:0] node28331;
	wire [4-1:0] node28332;
	wire [4-1:0] node28333;
	wire [4-1:0] node28337;
	wire [4-1:0] node28338;
	wire [4-1:0] node28342;
	wire [4-1:0] node28343;
	wire [4-1:0] node28344;
	wire [4-1:0] node28345;
	wire [4-1:0] node28346;
	wire [4-1:0] node28347;
	wire [4-1:0] node28348;
	wire [4-1:0] node28349;
	wire [4-1:0] node28350;
	wire [4-1:0] node28351;
	wire [4-1:0] node28352;
	wire [4-1:0] node28353;
	wire [4-1:0] node28354;
	wire [4-1:0] node28355;
	wire [4-1:0] node28356;
	wire [4-1:0] node28360;
	wire [4-1:0] node28361;
	wire [4-1:0] node28365;
	wire [4-1:0] node28367;
	wire [4-1:0] node28369;
	wire [4-1:0] node28372;
	wire [4-1:0] node28373;
	wire [4-1:0] node28374;
	wire [4-1:0] node28375;
	wire [4-1:0] node28379;
	wire [4-1:0] node28381;
	wire [4-1:0] node28384;
	wire [4-1:0] node28385;
	wire [4-1:0] node28386;
	wire [4-1:0] node28390;
	wire [4-1:0] node28391;
	wire [4-1:0] node28395;
	wire [4-1:0] node28396;
	wire [4-1:0] node28397;
	wire [4-1:0] node28398;
	wire [4-1:0] node28399;
	wire [4-1:0] node28402;
	wire [4-1:0] node28405;
	wire [4-1:0] node28407;
	wire [4-1:0] node28410;
	wire [4-1:0] node28411;
	wire [4-1:0] node28412;
	wire [4-1:0] node28415;
	wire [4-1:0] node28418;
	wire [4-1:0] node28419;
	wire [4-1:0] node28422;
	wire [4-1:0] node28425;
	wire [4-1:0] node28426;
	wire [4-1:0] node28427;
	wire [4-1:0] node28428;
	wire [4-1:0] node28431;
	wire [4-1:0] node28435;
	wire [4-1:0] node28436;
	wire [4-1:0] node28439;
	wire [4-1:0] node28442;
	wire [4-1:0] node28443;
	wire [4-1:0] node28444;
	wire [4-1:0] node28445;
	wire [4-1:0] node28446;
	wire [4-1:0] node28449;
	wire [4-1:0] node28452;
	wire [4-1:0] node28453;
	wire [4-1:0] node28454;
	wire [4-1:0] node28457;
	wire [4-1:0] node28460;
	wire [4-1:0] node28461;
	wire [4-1:0] node28464;
	wire [4-1:0] node28467;
	wire [4-1:0] node28468;
	wire [4-1:0] node28469;
	wire [4-1:0] node28470;
	wire [4-1:0] node28474;
	wire [4-1:0] node28477;
	wire [4-1:0] node28478;
	wire [4-1:0] node28479;
	wire [4-1:0] node28483;
	wire [4-1:0] node28484;
	wire [4-1:0] node28488;
	wire [4-1:0] node28489;
	wire [4-1:0] node28490;
	wire [4-1:0] node28491;
	wire [4-1:0] node28493;
	wire [4-1:0] node28496;
	wire [4-1:0] node28497;
	wire [4-1:0] node28500;
	wire [4-1:0] node28503;
	wire [4-1:0] node28505;
	wire [4-1:0] node28506;
	wire [4-1:0] node28509;
	wire [4-1:0] node28512;
	wire [4-1:0] node28513;
	wire [4-1:0] node28514;
	wire [4-1:0] node28515;
	wire [4-1:0] node28518;
	wire [4-1:0] node28521;
	wire [4-1:0] node28522;
	wire [4-1:0] node28525;
	wire [4-1:0] node28528;
	wire [4-1:0] node28529;
	wire [4-1:0] node28532;
	wire [4-1:0] node28535;
	wire [4-1:0] node28536;
	wire [4-1:0] node28537;
	wire [4-1:0] node28538;
	wire [4-1:0] node28539;
	wire [4-1:0] node28540;
	wire [4-1:0] node28541;
	wire [4-1:0] node28545;
	wire [4-1:0] node28546;
	wire [4-1:0] node28549;
	wire [4-1:0] node28552;
	wire [4-1:0] node28553;
	wire [4-1:0] node28556;
	wire [4-1:0] node28557;
	wire [4-1:0] node28561;
	wire [4-1:0] node28562;
	wire [4-1:0] node28563;
	wire [4-1:0] node28566;
	wire [4-1:0] node28568;
	wire [4-1:0] node28571;
	wire [4-1:0] node28572;
	wire [4-1:0] node28575;
	wire [4-1:0] node28577;
	wire [4-1:0] node28580;
	wire [4-1:0] node28581;
	wire [4-1:0] node28582;
	wire [4-1:0] node28583;
	wire [4-1:0] node28587;
	wire [4-1:0] node28588;
	wire [4-1:0] node28591;
	wire [4-1:0] node28592;
	wire [4-1:0] node28595;
	wire [4-1:0] node28598;
	wire [4-1:0] node28599;
	wire [4-1:0] node28600;
	wire [4-1:0] node28601;
	wire [4-1:0] node28604;
	wire [4-1:0] node28607;
	wire [4-1:0] node28608;
	wire [4-1:0] node28612;
	wire [4-1:0] node28613;
	wire [4-1:0] node28614;
	wire [4-1:0] node28617;
	wire [4-1:0] node28620;
	wire [4-1:0] node28621;
	wire [4-1:0] node28625;
	wire [4-1:0] node28626;
	wire [4-1:0] node28627;
	wire [4-1:0] node28628;
	wire [4-1:0] node28629;
	wire [4-1:0] node28630;
	wire [4-1:0] node28633;
	wire [4-1:0] node28636;
	wire [4-1:0] node28638;
	wire [4-1:0] node28641;
	wire [4-1:0] node28642;
	wire [4-1:0] node28645;
	wire [4-1:0] node28648;
	wire [4-1:0] node28649;
	wire [4-1:0] node28650;
	wire [4-1:0] node28654;
	wire [4-1:0] node28655;
	wire [4-1:0] node28656;
	wire [4-1:0] node28659;
	wire [4-1:0] node28662;
	wire [4-1:0] node28663;
	wire [4-1:0] node28666;
	wire [4-1:0] node28669;
	wire [4-1:0] node28670;
	wire [4-1:0] node28671;
	wire [4-1:0] node28672;
	wire [4-1:0] node28674;
	wire [4-1:0] node28678;
	wire [4-1:0] node28679;
	wire [4-1:0] node28680;
	wire [4-1:0] node28684;
	wire [4-1:0] node28685;
	wire [4-1:0] node28689;
	wire [4-1:0] node28690;
	wire [4-1:0] node28691;
	wire [4-1:0] node28692;
	wire [4-1:0] node28696;
	wire [4-1:0] node28697;
	wire [4-1:0] node28701;
	wire [4-1:0] node28702;
	wire [4-1:0] node28703;
	wire [4-1:0] node28706;
	wire [4-1:0] node28709;
	wire [4-1:0] node28710;
	wire [4-1:0] node28713;
	wire [4-1:0] node28716;
	wire [4-1:0] node28717;
	wire [4-1:0] node28718;
	wire [4-1:0] node28719;
	wire [4-1:0] node28720;
	wire [4-1:0] node28721;
	wire [4-1:0] node28722;
	wire [4-1:0] node28723;
	wire [4-1:0] node28726;
	wire [4-1:0] node28729;
	wire [4-1:0] node28731;
	wire [4-1:0] node28734;
	wire [4-1:0] node28735;
	wire [4-1:0] node28736;
	wire [4-1:0] node28739;
	wire [4-1:0] node28742;
	wire [4-1:0] node28743;
	wire [4-1:0] node28746;
	wire [4-1:0] node28749;
	wire [4-1:0] node28750;
	wire [4-1:0] node28751;
	wire [4-1:0] node28754;
	wire [4-1:0] node28757;
	wire [4-1:0] node28758;
	wire [4-1:0] node28759;
	wire [4-1:0] node28762;
	wire [4-1:0] node28765;
	wire [4-1:0] node28766;
	wire [4-1:0] node28769;
	wire [4-1:0] node28772;
	wire [4-1:0] node28773;
	wire [4-1:0] node28774;
	wire [4-1:0] node28776;
	wire [4-1:0] node28779;
	wire [4-1:0] node28780;
	wire [4-1:0] node28784;
	wire [4-1:0] node28785;
	wire [4-1:0] node28787;
	wire [4-1:0] node28790;
	wire [4-1:0] node28792;
	wire [4-1:0] node28795;
	wire [4-1:0] node28796;
	wire [4-1:0] node28797;
	wire [4-1:0] node28798;
	wire [4-1:0] node28799;
	wire [4-1:0] node28800;
	wire [4-1:0] node28804;
	wire [4-1:0] node28807;
	wire [4-1:0] node28808;
	wire [4-1:0] node28809;
	wire [4-1:0] node28813;
	wire [4-1:0] node28816;
	wire [4-1:0] node28817;
	wire [4-1:0] node28818;
	wire [4-1:0] node28820;
	wire [4-1:0] node28824;
	wire [4-1:0] node28825;
	wire [4-1:0] node28829;
	wire [4-1:0] node28830;
	wire [4-1:0] node28831;
	wire [4-1:0] node28832;
	wire [4-1:0] node28834;
	wire [4-1:0] node28837;
	wire [4-1:0] node28839;
	wire [4-1:0] node28842;
	wire [4-1:0] node28843;
	wire [4-1:0] node28846;
	wire [4-1:0] node28849;
	wire [4-1:0] node28850;
	wire [4-1:0] node28851;
	wire [4-1:0] node28852;
	wire [4-1:0] node28855;
	wire [4-1:0] node28858;
	wire [4-1:0] node28860;
	wire [4-1:0] node28863;
	wire [4-1:0] node28864;
	wire [4-1:0] node28865;
	wire [4-1:0] node28868;
	wire [4-1:0] node28871;
	wire [4-1:0] node28872;
	wire [4-1:0] node28875;
	wire [4-1:0] node28878;
	wire [4-1:0] node28879;
	wire [4-1:0] node28880;
	wire [4-1:0] node28881;
	wire [4-1:0] node28882;
	wire [4-1:0] node28883;
	wire [4-1:0] node28884;
	wire [4-1:0] node28887;
	wire [4-1:0] node28890;
	wire [4-1:0] node28891;
	wire [4-1:0] node28895;
	wire [4-1:0] node28896;
	wire [4-1:0] node28897;
	wire [4-1:0] node28900;
	wire [4-1:0] node28903;
	wire [4-1:0] node28904;
	wire [4-1:0] node28907;
	wire [4-1:0] node28910;
	wire [4-1:0] node28911;
	wire [4-1:0] node28912;
	wire [4-1:0] node28913;
	wire [4-1:0] node28916;
	wire [4-1:0] node28919;
	wire [4-1:0] node28922;
	wire [4-1:0] node28923;
	wire [4-1:0] node28924;
	wire [4-1:0] node28928;
	wire [4-1:0] node28929;
	wire [4-1:0] node28933;
	wire [4-1:0] node28934;
	wire [4-1:0] node28935;
	wire [4-1:0] node28936;
	wire [4-1:0] node28939;
	wire [4-1:0] node28941;
	wire [4-1:0] node28944;
	wire [4-1:0] node28945;
	wire [4-1:0] node28948;
	wire [4-1:0] node28950;
	wire [4-1:0] node28953;
	wire [4-1:0] node28954;
	wire [4-1:0] node28955;
	wire [4-1:0] node28958;
	wire [4-1:0] node28961;
	wire [4-1:0] node28963;
	wire [4-1:0] node28965;
	wire [4-1:0] node28968;
	wire [4-1:0] node28969;
	wire [4-1:0] node28970;
	wire [4-1:0] node28971;
	wire [4-1:0] node28972;
	wire [4-1:0] node28975;
	wire [4-1:0] node28978;
	wire [4-1:0] node28979;
	wire [4-1:0] node28980;
	wire [4-1:0] node28983;
	wire [4-1:0] node28986;
	wire [4-1:0] node28988;
	wire [4-1:0] node28991;
	wire [4-1:0] node28992;
	wire [4-1:0] node28993;
	wire [4-1:0] node28994;
	wire [4-1:0] node28998;
	wire [4-1:0] node28999;
	wire [4-1:0] node29003;
	wire [4-1:0] node29004;
	wire [4-1:0] node29005;
	wire [4-1:0] node29009;
	wire [4-1:0] node29010;
	wire [4-1:0] node29014;
	wire [4-1:0] node29015;
	wire [4-1:0] node29016;
	wire [4-1:0] node29017;
	wire [4-1:0] node29020;
	wire [4-1:0] node29023;
	wire [4-1:0] node29024;
	wire [4-1:0] node29025;
	wire [4-1:0] node29028;
	wire [4-1:0] node29031;
	wire [4-1:0] node29033;
	wire [4-1:0] node29036;
	wire [4-1:0] node29037;
	wire [4-1:0] node29038;
	wire [4-1:0] node29039;
	wire [4-1:0] node29043;
	wire [4-1:0] node29044;
	wire [4-1:0] node29048;
	wire [4-1:0] node29049;
	wire [4-1:0] node29051;
	wire [4-1:0] node29054;
	wire [4-1:0] node29055;
	wire [4-1:0] node29059;
	wire [4-1:0] node29060;
	wire [4-1:0] node29061;
	wire [4-1:0] node29062;
	wire [4-1:0] node29063;
	wire [4-1:0] node29064;
	wire [4-1:0] node29065;
	wire [4-1:0] node29066;
	wire [4-1:0] node29068;
	wire [4-1:0] node29072;
	wire [4-1:0] node29073;
	wire [4-1:0] node29074;
	wire [4-1:0] node29078;
	wire [4-1:0] node29079;
	wire [4-1:0] node29083;
	wire [4-1:0] node29084;
	wire [4-1:0] node29085;
	wire [4-1:0] node29086;
	wire [4-1:0] node29089;
	wire [4-1:0] node29093;
	wire [4-1:0] node29094;
	wire [4-1:0] node29095;
	wire [4-1:0] node29099;
	wire [4-1:0] node29100;
	wire [4-1:0] node29104;
	wire [4-1:0] node29105;
	wire [4-1:0] node29106;
	wire [4-1:0] node29107;
	wire [4-1:0] node29109;
	wire [4-1:0] node29112;
	wire [4-1:0] node29113;
	wire [4-1:0] node29116;
	wire [4-1:0] node29119;
	wire [4-1:0] node29121;
	wire [4-1:0] node29124;
	wire [4-1:0] node29125;
	wire [4-1:0] node29126;
	wire [4-1:0] node29127;
	wire [4-1:0] node29131;
	wire [4-1:0] node29133;
	wire [4-1:0] node29136;
	wire [4-1:0] node29138;
	wire [4-1:0] node29139;
	wire [4-1:0] node29143;
	wire [4-1:0] node29144;
	wire [4-1:0] node29145;
	wire [4-1:0] node29146;
	wire [4-1:0] node29147;
	wire [4-1:0] node29148;
	wire [4-1:0] node29151;
	wire [4-1:0] node29154;
	wire [4-1:0] node29155;
	wire [4-1:0] node29159;
	wire [4-1:0] node29160;
	wire [4-1:0] node29161;
	wire [4-1:0] node29164;
	wire [4-1:0] node29167;
	wire [4-1:0] node29168;
	wire [4-1:0] node29171;
	wire [4-1:0] node29174;
	wire [4-1:0] node29175;
	wire [4-1:0] node29176;
	wire [4-1:0] node29177;
	wire [4-1:0] node29181;
	wire [4-1:0] node29182;
	wire [4-1:0] node29185;
	wire [4-1:0] node29188;
	wire [4-1:0] node29189;
	wire [4-1:0] node29190;
	wire [4-1:0] node29193;
	wire [4-1:0] node29196;
	wire [4-1:0] node29197;
	wire [4-1:0] node29201;
	wire [4-1:0] node29202;
	wire [4-1:0] node29203;
	wire [4-1:0] node29204;
	wire [4-1:0] node29207;
	wire [4-1:0] node29210;
	wire [4-1:0] node29211;
	wire [4-1:0] node29214;
	wire [4-1:0] node29216;
	wire [4-1:0] node29219;
	wire [4-1:0] node29220;
	wire [4-1:0] node29221;
	wire [4-1:0] node29224;
	wire [4-1:0] node29227;
	wire [4-1:0] node29228;
	wire [4-1:0] node29231;
	wire [4-1:0] node29233;
	wire [4-1:0] node29236;
	wire [4-1:0] node29237;
	wire [4-1:0] node29238;
	wire [4-1:0] node29239;
	wire [4-1:0] node29240;
	wire [4-1:0] node29241;
	wire [4-1:0] node29244;
	wire [4-1:0] node29247;
	wire [4-1:0] node29248;
	wire [4-1:0] node29249;
	wire [4-1:0] node29252;
	wire [4-1:0] node29255;
	wire [4-1:0] node29256;
	wire [4-1:0] node29259;
	wire [4-1:0] node29262;
	wire [4-1:0] node29263;
	wire [4-1:0] node29264;
	wire [4-1:0] node29267;
	wire [4-1:0] node29270;
	wire [4-1:0] node29271;
	wire [4-1:0] node29273;
	wire [4-1:0] node29276;
	wire [4-1:0] node29277;
	wire [4-1:0] node29280;
	wire [4-1:0] node29283;
	wire [4-1:0] node29284;
	wire [4-1:0] node29285;
	wire [4-1:0] node29286;
	wire [4-1:0] node29289;
	wire [4-1:0] node29290;
	wire [4-1:0] node29294;
	wire [4-1:0] node29295;
	wire [4-1:0] node29298;
	wire [4-1:0] node29300;
	wire [4-1:0] node29303;
	wire [4-1:0] node29304;
	wire [4-1:0] node29305;
	wire [4-1:0] node29306;
	wire [4-1:0] node29309;
	wire [4-1:0] node29312;
	wire [4-1:0] node29314;
	wire [4-1:0] node29317;
	wire [4-1:0] node29318;
	wire [4-1:0] node29319;
	wire [4-1:0] node29323;
	wire [4-1:0] node29325;
	wire [4-1:0] node29328;
	wire [4-1:0] node29329;
	wire [4-1:0] node29330;
	wire [4-1:0] node29331;
	wire [4-1:0] node29332;
	wire [4-1:0] node29333;
	wire [4-1:0] node29337;
	wire [4-1:0] node29338;
	wire [4-1:0] node29342;
	wire [4-1:0] node29343;
	wire [4-1:0] node29345;
	wire [4-1:0] node29348;
	wire [4-1:0] node29350;
	wire [4-1:0] node29353;
	wire [4-1:0] node29354;
	wire [4-1:0] node29356;
	wire [4-1:0] node29358;
	wire [4-1:0] node29361;
	wire [4-1:0] node29362;
	wire [4-1:0] node29363;
	wire [4-1:0] node29367;
	wire [4-1:0] node29368;
	wire [4-1:0] node29372;
	wire [4-1:0] node29373;
	wire [4-1:0] node29374;
	wire [4-1:0] node29375;
	wire [4-1:0] node29377;
	wire [4-1:0] node29380;
	wire [4-1:0] node29382;
	wire [4-1:0] node29385;
	wire [4-1:0] node29386;
	wire [4-1:0] node29387;
	wire [4-1:0] node29390;
	wire [4-1:0] node29394;
	wire [4-1:0] node29395;
	wire [4-1:0] node29396;
	wire [4-1:0] node29397;
	wire [4-1:0] node29401;
	wire [4-1:0] node29404;
	wire [4-1:0] node29405;
	wire [4-1:0] node29406;
	wire [4-1:0] node29410;
	wire [4-1:0] node29413;
	wire [4-1:0] node29414;
	wire [4-1:0] node29415;
	wire [4-1:0] node29416;
	wire [4-1:0] node29417;
	wire [4-1:0] node29418;
	wire [4-1:0] node29419;
	wire [4-1:0] node29420;
	wire [4-1:0] node29423;
	wire [4-1:0] node29427;
	wire [4-1:0] node29428;
	wire [4-1:0] node29429;
	wire [4-1:0] node29432;
	wire [4-1:0] node29435;
	wire [4-1:0] node29436;
	wire [4-1:0] node29439;
	wire [4-1:0] node29442;
	wire [4-1:0] node29443;
	wire [4-1:0] node29444;
	wire [4-1:0] node29445;
	wire [4-1:0] node29449;
	wire [4-1:0] node29450;
	wire [4-1:0] node29453;
	wire [4-1:0] node29456;
	wire [4-1:0] node29457;
	wire [4-1:0] node29458;
	wire [4-1:0] node29461;
	wire [4-1:0] node29464;
	wire [4-1:0] node29465;
	wire [4-1:0] node29468;
	wire [4-1:0] node29471;
	wire [4-1:0] node29472;
	wire [4-1:0] node29473;
	wire [4-1:0] node29474;
	wire [4-1:0] node29476;
	wire [4-1:0] node29479;
	wire [4-1:0] node29482;
	wire [4-1:0] node29483;
	wire [4-1:0] node29484;
	wire [4-1:0] node29488;
	wire [4-1:0] node29489;
	wire [4-1:0] node29493;
	wire [4-1:0] node29494;
	wire [4-1:0] node29496;
	wire [4-1:0] node29497;
	wire [4-1:0] node29501;
	wire [4-1:0] node29502;
	wire [4-1:0] node29503;
	wire [4-1:0] node29508;
	wire [4-1:0] node29509;
	wire [4-1:0] node29510;
	wire [4-1:0] node29511;
	wire [4-1:0] node29512;
	wire [4-1:0] node29513;
	wire [4-1:0] node29516;
	wire [4-1:0] node29519;
	wire [4-1:0] node29520;
	wire [4-1:0] node29523;
	wire [4-1:0] node29526;
	wire [4-1:0] node29527;
	wire [4-1:0] node29528;
	wire [4-1:0] node29531;
	wire [4-1:0] node29534;
	wire [4-1:0] node29535;
	wire [4-1:0] node29538;
	wire [4-1:0] node29541;
	wire [4-1:0] node29542;
	wire [4-1:0] node29543;
	wire [4-1:0] node29544;
	wire [4-1:0] node29547;
	wire [4-1:0] node29550;
	wire [4-1:0] node29551;
	wire [4-1:0] node29554;
	wire [4-1:0] node29557;
	wire [4-1:0] node29558;
	wire [4-1:0] node29559;
	wire [4-1:0] node29562;
	wire [4-1:0] node29565;
	wire [4-1:0] node29566;
	wire [4-1:0] node29570;
	wire [4-1:0] node29571;
	wire [4-1:0] node29572;
	wire [4-1:0] node29574;
	wire [4-1:0] node29575;
	wire [4-1:0] node29578;
	wire [4-1:0] node29581;
	wire [4-1:0] node29582;
	wire [4-1:0] node29583;
	wire [4-1:0] node29586;
	wire [4-1:0] node29589;
	wire [4-1:0] node29591;
	wire [4-1:0] node29594;
	wire [4-1:0] node29595;
	wire [4-1:0] node29596;
	wire [4-1:0] node29597;
	wire [4-1:0] node29600;
	wire [4-1:0] node29603;
	wire [4-1:0] node29604;
	wire [4-1:0] node29608;
	wire [4-1:0] node29609;
	wire [4-1:0] node29610;
	wire [4-1:0] node29613;
	wire [4-1:0] node29616;
	wire [4-1:0] node29617;
	wire [4-1:0] node29621;
	wire [4-1:0] node29622;
	wire [4-1:0] node29623;
	wire [4-1:0] node29624;
	wire [4-1:0] node29625;
	wire [4-1:0] node29626;
	wire [4-1:0] node29628;
	wire [4-1:0] node29631;
	wire [4-1:0] node29633;
	wire [4-1:0] node29636;
	wire [4-1:0] node29637;
	wire [4-1:0] node29640;
	wire [4-1:0] node29643;
	wire [4-1:0] node29644;
	wire [4-1:0] node29645;
	wire [4-1:0] node29647;
	wire [4-1:0] node29651;
	wire [4-1:0] node29652;
	wire [4-1:0] node29655;
	wire [4-1:0] node29657;
	wire [4-1:0] node29660;
	wire [4-1:0] node29661;
	wire [4-1:0] node29662;
	wire [4-1:0] node29663;
	wire [4-1:0] node29666;
	wire [4-1:0] node29669;
	wire [4-1:0] node29670;
	wire [4-1:0] node29672;
	wire [4-1:0] node29675;
	wire [4-1:0] node29676;
	wire [4-1:0] node29679;
	wire [4-1:0] node29682;
	wire [4-1:0] node29683;
	wire [4-1:0] node29684;
	wire [4-1:0] node29685;
	wire [4-1:0] node29689;
	wire [4-1:0] node29692;
	wire [4-1:0] node29693;
	wire [4-1:0] node29697;
	wire [4-1:0] node29698;
	wire [4-1:0] node29699;
	wire [4-1:0] node29700;
	wire [4-1:0] node29701;
	wire [4-1:0] node29704;
	wire [4-1:0] node29707;
	wire [4-1:0] node29708;
	wire [4-1:0] node29709;
	wire [4-1:0] node29712;
	wire [4-1:0] node29715;
	wire [4-1:0] node29716;
	wire [4-1:0] node29720;
	wire [4-1:0] node29721;
	wire [4-1:0] node29722;
	wire [4-1:0] node29723;
	wire [4-1:0] node29726;
	wire [4-1:0] node29729;
	wire [4-1:0] node29730;
	wire [4-1:0] node29734;
	wire [4-1:0] node29735;
	wire [4-1:0] node29738;
	wire [4-1:0] node29741;
	wire [4-1:0] node29742;
	wire [4-1:0] node29743;
	wire [4-1:0] node29745;
	wire [4-1:0] node29748;
	wire [4-1:0] node29749;
	wire [4-1:0] node29750;
	wire [4-1:0] node29754;
	wire [4-1:0] node29755;
	wire [4-1:0] node29759;
	wire [4-1:0] node29760;
	wire [4-1:0] node29761;
	wire [4-1:0] node29762;
	wire [4-1:0] node29766;
	wire [4-1:0] node29768;
	wire [4-1:0] node29771;
	wire [4-1:0] node29772;
	wire [4-1:0] node29776;
	wire [4-1:0] node29777;
	wire [4-1:0] node29778;
	wire [4-1:0] node29779;
	wire [4-1:0] node29780;
	wire [4-1:0] node29781;
	wire [4-1:0] node29782;
	wire [4-1:0] node29784;
	wire [4-1:0] node29785;
	wire [4-1:0] node29789;
	wire [4-1:0] node29791;
	wire [4-1:0] node29792;
	wire [4-1:0] node29795;
	wire [4-1:0] node29798;
	wire [4-1:0] node29799;
	wire [4-1:0] node29800;
	wire [4-1:0] node29801;
	wire [4-1:0] node29805;
	wire [4-1:0] node29807;
	wire [4-1:0] node29810;
	wire [4-1:0] node29811;
	wire [4-1:0] node29813;
	wire [4-1:0] node29816;
	wire [4-1:0] node29818;
	wire [4-1:0] node29821;
	wire [4-1:0] node29822;
	wire [4-1:0] node29823;
	wire [4-1:0] node29824;
	wire [4-1:0] node29825;
	wire [4-1:0] node29829;
	wire [4-1:0] node29830;
	wire [4-1:0] node29833;
	wire [4-1:0] node29836;
	wire [4-1:0] node29838;
	wire [4-1:0] node29839;
	wire [4-1:0] node29843;
	wire [4-1:0] node29844;
	wire [4-1:0] node29845;
	wire [4-1:0] node29846;
	wire [4-1:0] node29850;
	wire [4-1:0] node29851;
	wire [4-1:0] node29855;
	wire [4-1:0] node29856;
	wire [4-1:0] node29858;
	wire [4-1:0] node29861;
	wire [4-1:0] node29863;
	wire [4-1:0] node29866;
	wire [4-1:0] node29867;
	wire [4-1:0] node29868;
	wire [4-1:0] node29869;
	wire [4-1:0] node29870;
	wire [4-1:0] node29872;
	wire [4-1:0] node29876;
	wire [4-1:0] node29877;
	wire [4-1:0] node29878;
	wire [4-1:0] node29879;
	wire [4-1:0] node29882;
	wire [4-1:0] node29885;
	wire [4-1:0] node29886;
	wire [4-1:0] node29889;
	wire [4-1:0] node29892;
	wire [4-1:0] node29893;
	wire [4-1:0] node29897;
	wire [4-1:0] node29898;
	wire [4-1:0] node29899;
	wire [4-1:0] node29901;
	wire [4-1:0] node29904;
	wire [4-1:0] node29905;
	wire [4-1:0] node29909;
	wire [4-1:0] node29910;
	wire [4-1:0] node29912;
	wire [4-1:0] node29915;
	wire [4-1:0] node29917;
	wire [4-1:0] node29920;
	wire [4-1:0] node29921;
	wire [4-1:0] node29922;
	wire [4-1:0] node29924;
	wire [4-1:0] node29925;
	wire [4-1:0] node29929;
	wire [4-1:0] node29930;
	wire [4-1:0] node29931;
	wire [4-1:0] node29934;
	wire [4-1:0] node29937;
	wire [4-1:0] node29938;
	wire [4-1:0] node29942;
	wire [4-1:0] node29943;
	wire [4-1:0] node29944;
	wire [4-1:0] node29945;
	wire [4-1:0] node29949;
	wire [4-1:0] node29950;
	wire [4-1:0] node29954;
	wire [4-1:0] node29955;
	wire [4-1:0] node29957;
	wire [4-1:0] node29960;
	wire [4-1:0] node29961;
	wire [4-1:0] node29965;
	wire [4-1:0] node29966;
	wire [4-1:0] node29967;
	wire [4-1:0] node29968;
	wire [4-1:0] node29969;
	wire [4-1:0] node29971;
	wire [4-1:0] node29974;
	wire [4-1:0] node29975;
	wire [4-1:0] node29977;
	wire [4-1:0] node29980;
	wire [4-1:0] node29983;
	wire [4-1:0] node29984;
	wire [4-1:0] node29985;
	wire [4-1:0] node29986;
	wire [4-1:0] node29990;
	wire [4-1:0] node29992;
	wire [4-1:0] node29995;
	wire [4-1:0] node29996;
	wire [4-1:0] node29997;
	wire [4-1:0] node30001;
	wire [4-1:0] node30003;
	wire [4-1:0] node30006;
	wire [4-1:0] node30007;
	wire [4-1:0] node30008;
	wire [4-1:0] node30010;
	wire [4-1:0] node30012;
	wire [4-1:0] node30015;
	wire [4-1:0] node30016;
	wire [4-1:0] node30019;
	wire [4-1:0] node30020;
	wire [4-1:0] node30024;
	wire [4-1:0] node30025;
	wire [4-1:0] node30026;
	wire [4-1:0] node30028;
	wire [4-1:0] node30031;
	wire [4-1:0] node30032;
	wire [4-1:0] node30036;
	wire [4-1:0] node30037;
	wire [4-1:0] node30038;
	wire [4-1:0] node30042;
	wire [4-1:0] node30044;
	wire [4-1:0] node30047;
	wire [4-1:0] node30048;
	wire [4-1:0] node30049;
	wire [4-1:0] node30050;
	wire [4-1:0] node30052;
	wire [4-1:0] node30054;
	wire [4-1:0] node30057;
	wire [4-1:0] node30058;
	wire [4-1:0] node30059;
	wire [4-1:0] node30060;
	wire [4-1:0] node30063;
	wire [4-1:0] node30066;
	wire [4-1:0] node30068;
	wire [4-1:0] node30071;
	wire [4-1:0] node30072;
	wire [4-1:0] node30076;
	wire [4-1:0] node30077;
	wire [4-1:0] node30078;
	wire [4-1:0] node30079;
	wire [4-1:0] node30084;
	wire [4-1:0] node30085;
	wire [4-1:0] node30086;
	wire [4-1:0] node30090;
	wire [4-1:0] node30092;
	wire [4-1:0] node30095;
	wire [4-1:0] node30096;
	wire [4-1:0] node30097;
	wire [4-1:0] node30098;
	wire [4-1:0] node30099;
	wire [4-1:0] node30103;
	wire [4-1:0] node30104;
	wire [4-1:0] node30107;
	wire [4-1:0] node30110;
	wire [4-1:0] node30111;
	wire [4-1:0] node30113;
	wire [4-1:0] node30117;
	wire [4-1:0] node30118;
	wire [4-1:0] node30119;
	wire [4-1:0] node30120;
	wire [4-1:0] node30124;
	wire [4-1:0] node30125;
	wire [4-1:0] node30129;
	wire [4-1:0] node30130;
	wire [4-1:0] node30132;
	wire [4-1:0] node30135;
	wire [4-1:0] node30136;
	wire [4-1:0] node30140;
	wire [4-1:0] node30141;
	wire [4-1:0] node30142;
	wire [4-1:0] node30143;
	wire [4-1:0] node30144;
	wire [4-1:0] node30145;
	wire [4-1:0] node30146;
	wire [4-1:0] node30148;
	wire [4-1:0] node30152;
	wire [4-1:0] node30153;
	wire [4-1:0] node30155;
	wire [4-1:0] node30158;
	wire [4-1:0] node30161;
	wire [4-1:0] node30162;
	wire [4-1:0] node30163;
	wire [4-1:0] node30165;
	wire [4-1:0] node30168;
	wire [4-1:0] node30170;
	wire [4-1:0] node30173;
	wire [4-1:0] node30175;
	wire [4-1:0] node30177;
	wire [4-1:0] node30180;
	wire [4-1:0] node30181;
	wire [4-1:0] node30182;
	wire [4-1:0] node30183;
	wire [4-1:0] node30184;
	wire [4-1:0] node30188;
	wire [4-1:0] node30189;
	wire [4-1:0] node30192;
	wire [4-1:0] node30195;
	wire [4-1:0] node30197;
	wire [4-1:0] node30198;
	wire [4-1:0] node30202;
	wire [4-1:0] node30203;
	wire [4-1:0] node30204;
	wire [4-1:0] node30207;
	wire [4-1:0] node30208;
	wire [4-1:0] node30212;
	wire [4-1:0] node30213;
	wire [4-1:0] node30214;
	wire [4-1:0] node30218;
	wire [4-1:0] node30220;
	wire [4-1:0] node30223;
	wire [4-1:0] node30224;
	wire [4-1:0] node30225;
	wire [4-1:0] node30226;
	wire [4-1:0] node30228;
	wire [4-1:0] node30229;
	wire [4-1:0] node30233;
	wire [4-1:0] node30234;
	wire [4-1:0] node30237;
	wire [4-1:0] node30239;
	wire [4-1:0] node30242;
	wire [4-1:0] node30243;
	wire [4-1:0] node30244;
	wire [4-1:0] node30246;
	wire [4-1:0] node30249;
	wire [4-1:0] node30250;
	wire [4-1:0] node30254;
	wire [4-1:0] node30255;
	wire [4-1:0] node30257;
	wire [4-1:0] node30260;
	wire [4-1:0] node30262;
	wire [4-1:0] node30265;
	wire [4-1:0] node30266;
	wire [4-1:0] node30267;
	wire [4-1:0] node30269;
	wire [4-1:0] node30271;
	wire [4-1:0] node30274;
	wire [4-1:0] node30275;
	wire [4-1:0] node30278;
	wire [4-1:0] node30280;
	wire [4-1:0] node30283;
	wire [4-1:0] node30284;
	wire [4-1:0] node30285;
	wire [4-1:0] node30286;
	wire [4-1:0] node30290;
	wire [4-1:0] node30291;
	wire [4-1:0] node30295;
	wire [4-1:0] node30296;
	wire [4-1:0] node30297;
	wire [4-1:0] node30301;
	wire [4-1:0] node30302;
	wire [4-1:0] node30306;
	wire [4-1:0] node30307;
	wire [4-1:0] node30308;
	wire [4-1:0] node30309;
	wire [4-1:0] node30310;
	wire [4-1:0] node30312;
	wire [4-1:0] node30314;
	wire [4-1:0] node30317;
	wire [4-1:0] node30318;
	wire [4-1:0] node30320;
	wire [4-1:0] node30323;
	wire [4-1:0] node30326;
	wire [4-1:0] node30327;
	wire [4-1:0] node30328;
	wire [4-1:0] node30330;
	wire [4-1:0] node30333;
	wire [4-1:0] node30335;
	wire [4-1:0] node30338;
	wire [4-1:0] node30339;
	wire [4-1:0] node30340;
	wire [4-1:0] node30344;
	wire [4-1:0] node30346;
	wire [4-1:0] node30349;
	wire [4-1:0] node30350;
	wire [4-1:0] node30351;
	wire [4-1:0] node30352;
	wire [4-1:0] node30353;
	wire [4-1:0] node30357;
	wire [4-1:0] node30358;
	wire [4-1:0] node30361;
	wire [4-1:0] node30364;
	wire [4-1:0] node30366;
	wire [4-1:0] node30367;
	wire [4-1:0] node30371;
	wire [4-1:0] node30372;
	wire [4-1:0] node30373;
	wire [4-1:0] node30375;
	wire [4-1:0] node30378;
	wire [4-1:0] node30381;
	wire [4-1:0] node30382;
	wire [4-1:0] node30383;
	wire [4-1:0] node30387;
	wire [4-1:0] node30389;
	wire [4-1:0] node30392;
	wire [4-1:0] node30393;
	wire [4-1:0] node30394;
	wire [4-1:0] node30395;
	wire [4-1:0] node30396;
	wire [4-1:0] node30399;
	wire [4-1:0] node30401;
	wire [4-1:0] node30404;
	wire [4-1:0] node30406;
	wire [4-1:0] node30408;
	wire [4-1:0] node30411;
	wire [4-1:0] node30412;
	wire [4-1:0] node30413;
	wire [4-1:0] node30414;
	wire [4-1:0] node30418;
	wire [4-1:0] node30419;
	wire [4-1:0] node30423;
	wire [4-1:0] node30424;
	wire [4-1:0] node30426;
	wire [4-1:0] node30429;
	wire [4-1:0] node30431;
	wire [4-1:0] node30434;
	wire [4-1:0] node30435;
	wire [4-1:0] node30436;
	wire [4-1:0] node30437;
	wire [4-1:0] node30439;
	wire [4-1:0] node30443;
	wire [4-1:0] node30444;
	wire [4-1:0] node30445;
	wire [4-1:0] node30448;
	wire [4-1:0] node30451;
	wire [4-1:0] node30452;
	wire [4-1:0] node30456;
	wire [4-1:0] node30457;
	wire [4-1:0] node30458;
	wire [4-1:0] node30460;
	wire [4-1:0] node30463;
	wire [4-1:0] node30464;
	wire [4-1:0] node30468;
	wire [4-1:0] node30469;
	wire [4-1:0] node30471;
	wire [4-1:0] node30474;
	wire [4-1:0] node30475;
	wire [4-1:0] node30479;
	wire [4-1:0] node30480;
	wire [4-1:0] node30481;
	wire [4-1:0] node30482;
	wire [4-1:0] node30483;
	wire [4-1:0] node30484;
	wire [4-1:0] node30485;
	wire [4-1:0] node30486;
	wire [4-1:0] node30487;
	wire [4-1:0] node30488;
	wire [4-1:0] node30489;
	wire [4-1:0] node30492;
	wire [4-1:0] node30496;
	wire [4-1:0] node30497;
	wire [4-1:0] node30498;
	wire [4-1:0] node30501;
	wire [4-1:0] node30504;
	wire [4-1:0] node30505;
	wire [4-1:0] node30508;
	wire [4-1:0] node30511;
	wire [4-1:0] node30512;
	wire [4-1:0] node30513;
	wire [4-1:0] node30515;
	wire [4-1:0] node30518;
	wire [4-1:0] node30521;
	wire [4-1:0] node30522;
	wire [4-1:0] node30523;
	wire [4-1:0] node30526;
	wire [4-1:0] node30529;
	wire [4-1:0] node30531;
	wire [4-1:0] node30534;
	wire [4-1:0] node30535;
	wire [4-1:0] node30536;
	wire [4-1:0] node30537;
	wire [4-1:0] node30539;
	wire [4-1:0] node30542;
	wire [4-1:0] node30543;
	wire [4-1:0] node30547;
	wire [4-1:0] node30548;
	wire [4-1:0] node30551;
	wire [4-1:0] node30552;
	wire [4-1:0] node30556;
	wire [4-1:0] node30557;
	wire [4-1:0] node30558;
	wire [4-1:0] node30559;
	wire [4-1:0] node30562;
	wire [4-1:0] node30565;
	wire [4-1:0] node30566;
	wire [4-1:0] node30569;
	wire [4-1:0] node30572;
	wire [4-1:0] node30574;
	wire [4-1:0] node30575;
	wire [4-1:0] node30578;
	wire [4-1:0] node30581;
	wire [4-1:0] node30582;
	wire [4-1:0] node30583;
	wire [4-1:0] node30584;
	wire [4-1:0] node30586;
	wire [4-1:0] node30587;
	wire [4-1:0] node30591;
	wire [4-1:0] node30592;
	wire [4-1:0] node30593;
	wire [4-1:0] node30597;
	wire [4-1:0] node30598;
	wire [4-1:0] node30602;
	wire [4-1:0] node30603;
	wire [4-1:0] node30604;
	wire [4-1:0] node30605;
	wire [4-1:0] node30609;
	wire [4-1:0] node30611;
	wire [4-1:0] node30614;
	wire [4-1:0] node30616;
	wire [4-1:0] node30617;
	wire [4-1:0] node30621;
	wire [4-1:0] node30622;
	wire [4-1:0] node30623;
	wire [4-1:0] node30624;
	wire [4-1:0] node30626;
	wire [4-1:0] node30629;
	wire [4-1:0] node30631;
	wire [4-1:0] node30634;
	wire [4-1:0] node30635;
	wire [4-1:0] node30638;
	wire [4-1:0] node30641;
	wire [4-1:0] node30642;
	wire [4-1:0] node30643;
	wire [4-1:0] node30644;
	wire [4-1:0] node30649;
	wire [4-1:0] node30650;
	wire [4-1:0] node30651;
	wire [4-1:0] node30655;
	wire [4-1:0] node30656;
	wire [4-1:0] node30660;
	wire [4-1:0] node30661;
	wire [4-1:0] node30662;
	wire [4-1:0] node30663;
	wire [4-1:0] node30664;
	wire [4-1:0] node30665;
	wire [4-1:0] node30667;
	wire [4-1:0] node30670;
	wire [4-1:0] node30671;
	wire [4-1:0] node30675;
	wire [4-1:0] node30676;
	wire [4-1:0] node30679;
	wire [4-1:0] node30680;
	wire [4-1:0] node30684;
	wire [4-1:0] node30685;
	wire [4-1:0] node30688;
	wire [4-1:0] node30689;
	wire [4-1:0] node30692;
	wire [4-1:0] node30693;
	wire [4-1:0] node30697;
	wire [4-1:0] node30698;
	wire [4-1:0] node30699;
	wire [4-1:0] node30700;
	wire [4-1:0] node30701;
	wire [4-1:0] node30705;
	wire [4-1:0] node30708;
	wire [4-1:0] node30709;
	wire [4-1:0] node30711;
	wire [4-1:0] node30714;
	wire [4-1:0] node30715;
	wire [4-1:0] node30718;
	wire [4-1:0] node30721;
	wire [4-1:0] node30722;
	wire [4-1:0] node30723;
	wire [4-1:0] node30724;
	wire [4-1:0] node30727;
	wire [4-1:0] node30730;
	wire [4-1:0] node30731;
	wire [4-1:0] node30734;
	wire [4-1:0] node30737;
	wire [4-1:0] node30738;
	wire [4-1:0] node30739;
	wire [4-1:0] node30742;
	wire [4-1:0] node30745;
	wire [4-1:0] node30747;
	wire [4-1:0] node30750;
	wire [4-1:0] node30751;
	wire [4-1:0] node30752;
	wire [4-1:0] node30753;
	wire [4-1:0] node30754;
	wire [4-1:0] node30755;
	wire [4-1:0] node30759;
	wire [4-1:0] node30760;
	wire [4-1:0] node30763;
	wire [4-1:0] node30766;
	wire [4-1:0] node30767;
	wire [4-1:0] node30769;
	wire [4-1:0] node30772;
	wire [4-1:0] node30773;
	wire [4-1:0] node30776;
	wire [4-1:0] node30779;
	wire [4-1:0] node30780;
	wire [4-1:0] node30781;
	wire [4-1:0] node30782;
	wire [4-1:0] node30786;
	wire [4-1:0] node30787;
	wire [4-1:0] node30790;
	wire [4-1:0] node30793;
	wire [4-1:0] node30794;
	wire [4-1:0] node30796;
	wire [4-1:0] node30799;
	wire [4-1:0] node30802;
	wire [4-1:0] node30803;
	wire [4-1:0] node30804;
	wire [4-1:0] node30805;
	wire [4-1:0] node30806;
	wire [4-1:0] node30809;
	wire [4-1:0] node30812;
	wire [4-1:0] node30814;
	wire [4-1:0] node30817;
	wire [4-1:0] node30818;
	wire [4-1:0] node30819;
	wire [4-1:0] node30822;
	wire [4-1:0] node30825;
	wire [4-1:0] node30826;
	wire [4-1:0] node30829;
	wire [4-1:0] node30832;
	wire [4-1:0] node30833;
	wire [4-1:0] node30834;
	wire [4-1:0] node30836;
	wire [4-1:0] node30839;
	wire [4-1:0] node30842;
	wire [4-1:0] node30843;
	wire [4-1:0] node30846;
	wire [4-1:0] node30849;
	wire [4-1:0] node30850;
	wire [4-1:0] node30851;
	wire [4-1:0] node30852;
	wire [4-1:0] node30853;
	wire [4-1:0] node30854;
	wire [4-1:0] node30855;
	wire [4-1:0] node30857;
	wire [4-1:0] node30860;
	wire [4-1:0] node30861;
	wire [4-1:0] node30865;
	wire [4-1:0] node30866;
	wire [4-1:0] node30868;
	wire [4-1:0] node30871;
	wire [4-1:0] node30872;
	wire [4-1:0] node30876;
	wire [4-1:0] node30877;
	wire [4-1:0] node30878;
	wire [4-1:0] node30879;
	wire [4-1:0] node30883;
	wire [4-1:0] node30884;
	wire [4-1:0] node30888;
	wire [4-1:0] node30889;
	wire [4-1:0] node30891;
	wire [4-1:0] node30894;
	wire [4-1:0] node30896;
	wire [4-1:0] node30899;
	wire [4-1:0] node30900;
	wire [4-1:0] node30901;
	wire [4-1:0] node30902;
	wire [4-1:0] node30905;
	wire [4-1:0] node30908;
	wire [4-1:0] node30909;
	wire [4-1:0] node30910;
	wire [4-1:0] node30913;
	wire [4-1:0] node30916;
	wire [4-1:0] node30917;
	wire [4-1:0] node30921;
	wire [4-1:0] node30922;
	wire [4-1:0] node30923;
	wire [4-1:0] node30924;
	wire [4-1:0] node30928;
	wire [4-1:0] node30929;
	wire [4-1:0] node30933;
	wire [4-1:0] node30934;
	wire [4-1:0] node30935;
	wire [4-1:0] node30938;
	wire [4-1:0] node30942;
	wire [4-1:0] node30943;
	wire [4-1:0] node30944;
	wire [4-1:0] node30945;
	wire [4-1:0] node30946;
	wire [4-1:0] node30950;
	wire [4-1:0] node30951;
	wire [4-1:0] node30952;
	wire [4-1:0] node30955;
	wire [4-1:0] node30958;
	wire [4-1:0] node30959;
	wire [4-1:0] node30962;
	wire [4-1:0] node30965;
	wire [4-1:0] node30966;
	wire [4-1:0] node30967;
	wire [4-1:0] node30970;
	wire [4-1:0] node30973;
	wire [4-1:0] node30974;
	wire [4-1:0] node30977;
	wire [4-1:0] node30980;
	wire [4-1:0] node30981;
	wire [4-1:0] node30982;
	wire [4-1:0] node30983;
	wire [4-1:0] node30984;
	wire [4-1:0] node30987;
	wire [4-1:0] node30990;
	wire [4-1:0] node30991;
	wire [4-1:0] node30994;
	wire [4-1:0] node30997;
	wire [4-1:0] node30998;
	wire [4-1:0] node30999;
	wire [4-1:0] node31002;
	wire [4-1:0] node31005;
	wire [4-1:0] node31006;
	wire [4-1:0] node31009;
	wire [4-1:0] node31012;
	wire [4-1:0] node31013;
	wire [4-1:0] node31014;
	wire [4-1:0] node31016;
	wire [4-1:0] node31019;
	wire [4-1:0] node31020;
	wire [4-1:0] node31024;
	wire [4-1:0] node31025;
	wire [4-1:0] node31026;
	wire [4-1:0] node31030;
	wire [4-1:0] node31032;
	wire [4-1:0] node31035;
	wire [4-1:0] node31036;
	wire [4-1:0] node31037;
	wire [4-1:0] node31038;
	wire [4-1:0] node31039;
	wire [4-1:0] node31040;
	wire [4-1:0] node31042;
	wire [4-1:0] node31045;
	wire [4-1:0] node31046;
	wire [4-1:0] node31050;
	wire [4-1:0] node31051;
	wire [4-1:0] node31054;
	wire [4-1:0] node31056;
	wire [4-1:0] node31059;
	wire [4-1:0] node31060;
	wire [4-1:0] node31062;
	wire [4-1:0] node31063;
	wire [4-1:0] node31067;
	wire [4-1:0] node31068;
	wire [4-1:0] node31070;
	wire [4-1:0] node31073;
	wire [4-1:0] node31075;
	wire [4-1:0] node31078;
	wire [4-1:0] node31079;
	wire [4-1:0] node31080;
	wire [4-1:0] node31081;
	wire [4-1:0] node31084;
	wire [4-1:0] node31087;
	wire [4-1:0] node31088;
	wire [4-1:0] node31089;
	wire [4-1:0] node31092;
	wire [4-1:0] node31095;
	wire [4-1:0] node31096;
	wire [4-1:0] node31099;
	wire [4-1:0] node31102;
	wire [4-1:0] node31103;
	wire [4-1:0] node31104;
	wire [4-1:0] node31105;
	wire [4-1:0] node31108;
	wire [4-1:0] node31111;
	wire [4-1:0] node31112;
	wire [4-1:0] node31115;
	wire [4-1:0] node31118;
	wire [4-1:0] node31119;
	wire [4-1:0] node31120;
	wire [4-1:0] node31123;
	wire [4-1:0] node31126;
	wire [4-1:0] node31127;
	wire [4-1:0] node31130;
	wire [4-1:0] node31133;
	wire [4-1:0] node31134;
	wire [4-1:0] node31135;
	wire [4-1:0] node31136;
	wire [4-1:0] node31137;
	wire [4-1:0] node31138;
	wire [4-1:0] node31141;
	wire [4-1:0] node31144;
	wire [4-1:0] node31145;
	wire [4-1:0] node31149;
	wire [4-1:0] node31150;
	wire [4-1:0] node31151;
	wire [4-1:0] node31155;
	wire [4-1:0] node31156;
	wire [4-1:0] node31159;
	wire [4-1:0] node31162;
	wire [4-1:0] node31163;
	wire [4-1:0] node31164;
	wire [4-1:0] node31165;
	wire [4-1:0] node31169;
	wire [4-1:0] node31170;
	wire [4-1:0] node31174;
	wire [4-1:0] node31176;
	wire [4-1:0] node31177;
	wire [4-1:0] node31180;
	wire [4-1:0] node31183;
	wire [4-1:0] node31184;
	wire [4-1:0] node31185;
	wire [4-1:0] node31186;
	wire [4-1:0] node31187;
	wire [4-1:0] node31190;
	wire [4-1:0] node31193;
	wire [4-1:0] node31194;
	wire [4-1:0] node31197;
	wire [4-1:0] node31200;
	wire [4-1:0] node31201;
	wire [4-1:0] node31202;
	wire [4-1:0] node31205;
	wire [4-1:0] node31208;
	wire [4-1:0] node31210;
	wire [4-1:0] node31213;
	wire [4-1:0] node31214;
	wire [4-1:0] node31215;
	wire [4-1:0] node31218;
	wire [4-1:0] node31221;
	wire [4-1:0] node31222;
	wire [4-1:0] node31225;
	wire [4-1:0] node31228;
	wire [4-1:0] node31229;
	wire [4-1:0] node31230;
	wire [4-1:0] node31231;
	wire [4-1:0] node31232;
	wire [4-1:0] node31233;
	wire [4-1:0] node31234;
	wire [4-1:0] node31235;
	wire [4-1:0] node31238;
	wire [4-1:0] node31241;
	wire [4-1:0] node31242;
	wire [4-1:0] node31245;
	wire [4-1:0] node31248;
	wire [4-1:0] node31249;
	wire [4-1:0] node31250;
	wire [4-1:0] node31251;
	wire [4-1:0] node31254;
	wire [4-1:0] node31257;
	wire [4-1:0] node31258;
	wire [4-1:0] node31261;
	wire [4-1:0] node31264;
	wire [4-1:0] node31265;
	wire [4-1:0] node31266;
	wire [4-1:0] node31269;
	wire [4-1:0] node31272;
	wire [4-1:0] node31273;
	wire [4-1:0] node31276;
	wire [4-1:0] node31279;
	wire [4-1:0] node31280;
	wire [4-1:0] node31281;
	wire [4-1:0] node31282;
	wire [4-1:0] node31285;
	wire [4-1:0] node31288;
	wire [4-1:0] node31290;
	wire [4-1:0] node31293;
	wire [4-1:0] node31294;
	wire [4-1:0] node31295;
	wire [4-1:0] node31298;
	wire [4-1:0] node31301;
	wire [4-1:0] node31302;
	wire [4-1:0] node31305;
	wire [4-1:0] node31308;
	wire [4-1:0] node31309;
	wire [4-1:0] node31310;
	wire [4-1:0] node31311;
	wire [4-1:0] node31312;
	wire [4-1:0] node31315;
	wire [4-1:0] node31318;
	wire [4-1:0] node31319;
	wire [4-1:0] node31320;
	wire [4-1:0] node31324;
	wire [4-1:0] node31325;
	wire [4-1:0] node31328;
	wire [4-1:0] node31331;
	wire [4-1:0] node31332;
	wire [4-1:0] node31333;
	wire [4-1:0] node31334;
	wire [4-1:0] node31337;
	wire [4-1:0] node31340;
	wire [4-1:0] node31341;
	wire [4-1:0] node31344;
	wire [4-1:0] node31347;
	wire [4-1:0] node31348;
	wire [4-1:0] node31351;
	wire [4-1:0] node31354;
	wire [4-1:0] node31355;
	wire [4-1:0] node31356;
	wire [4-1:0] node31357;
	wire [4-1:0] node31358;
	wire [4-1:0] node31361;
	wire [4-1:0] node31364;
	wire [4-1:0] node31365;
	wire [4-1:0] node31369;
	wire [4-1:0] node31370;
	wire [4-1:0] node31373;
	wire [4-1:0] node31376;
	wire [4-1:0] node31377;
	wire [4-1:0] node31378;
	wire [4-1:0] node31380;
	wire [4-1:0] node31383;
	wire [4-1:0] node31384;
	wire [4-1:0] node31387;
	wire [4-1:0] node31390;
	wire [4-1:0] node31391;
	wire [4-1:0] node31394;
	wire [4-1:0] node31397;
	wire [4-1:0] node31398;
	wire [4-1:0] node31399;
	wire [4-1:0] node31400;
	wire [4-1:0] node31401;
	wire [4-1:0] node31403;
	wire [4-1:0] node31405;
	wire [4-1:0] node31408;
	wire [4-1:0] node31409;
	wire [4-1:0] node31412;
	wire [4-1:0] node31415;
	wire [4-1:0] node31416;
	wire [4-1:0] node31417;
	wire [4-1:0] node31418;
	wire [4-1:0] node31421;
	wire [4-1:0] node31424;
	wire [4-1:0] node31425;
	wire [4-1:0] node31428;
	wire [4-1:0] node31431;
	wire [4-1:0] node31432;
	wire [4-1:0] node31433;
	wire [4-1:0] node31436;
	wire [4-1:0] node31439;
	wire [4-1:0] node31440;
	wire [4-1:0] node31443;
	wire [4-1:0] node31446;
	wire [4-1:0] node31447;
	wire [4-1:0] node31448;
	wire [4-1:0] node31449;
	wire [4-1:0] node31452;
	wire [4-1:0] node31455;
	wire [4-1:0] node31456;
	wire [4-1:0] node31459;
	wire [4-1:0] node31462;
	wire [4-1:0] node31463;
	wire [4-1:0] node31466;
	wire [4-1:0] node31469;
	wire [4-1:0] node31470;
	wire [4-1:0] node31471;
	wire [4-1:0] node31472;
	wire [4-1:0] node31474;
	wire [4-1:0] node31475;
	wire [4-1:0] node31479;
	wire [4-1:0] node31480;
	wire [4-1:0] node31481;
	wire [4-1:0] node31484;
	wire [4-1:0] node31488;
	wire [4-1:0] node31489;
	wire [4-1:0] node31492;
	wire [4-1:0] node31495;
	wire [4-1:0] node31496;
	wire [4-1:0] node31497;
	wire [4-1:0] node31498;
	wire [4-1:0] node31499;
	wire [4-1:0] node31502;
	wire [4-1:0] node31505;
	wire [4-1:0] node31506;
	wire [4-1:0] node31509;
	wire [4-1:0] node31512;
	wire [4-1:0] node31514;
	wire [4-1:0] node31517;
	wire [4-1:0] node31518;
	wire [4-1:0] node31521;
	wire [4-1:0] node31524;
	wire [4-1:0] node31525;
	wire [4-1:0] node31526;
	wire [4-1:0] node31527;
	wire [4-1:0] node31528;
	wire [4-1:0] node31529;
	wire [4-1:0] node31530;
	wire [4-1:0] node31533;
	wire [4-1:0] node31536;
	wire [4-1:0] node31537;
	wire [4-1:0] node31540;
	wire [4-1:0] node31543;
	wire [4-1:0] node31544;
	wire [4-1:0] node31545;
	wire [4-1:0] node31548;
	wire [4-1:0] node31551;
	wire [4-1:0] node31552;
	wire [4-1:0] node31555;
	wire [4-1:0] node31558;
	wire [4-1:0] node31559;
	wire [4-1:0] node31560;
	wire [4-1:0] node31561;
	wire [4-1:0] node31562;
	wire [4-1:0] node31565;
	wire [4-1:0] node31568;
	wire [4-1:0] node31569;
	wire [4-1:0] node31572;
	wire [4-1:0] node31575;
	wire [4-1:0] node31576;
	wire [4-1:0] node31579;
	wire [4-1:0] node31582;
	wire [4-1:0] node31583;
	wire [4-1:0] node31584;
	wire [4-1:0] node31587;
	wire [4-1:0] node31590;
	wire [4-1:0] node31591;
	wire [4-1:0] node31594;
	wire [4-1:0] node31597;
	wire [4-1:0] node31598;
	wire [4-1:0] node31599;
	wire [4-1:0] node31600;
	wire [4-1:0] node31601;
	wire [4-1:0] node31605;
	wire [4-1:0] node31606;
	wire [4-1:0] node31609;
	wire [4-1:0] node31612;
	wire [4-1:0] node31613;
	wire [4-1:0] node31614;
	wire [4-1:0] node31617;
	wire [4-1:0] node31620;
	wire [4-1:0] node31621;
	wire [4-1:0] node31624;
	wire [4-1:0] node31627;
	wire [4-1:0] node31628;
	wire [4-1:0] node31629;
	wire [4-1:0] node31631;
	wire [4-1:0] node31634;
	wire [4-1:0] node31635;
	wire [4-1:0] node31636;
	wire [4-1:0] node31639;
	wire [4-1:0] node31642;
	wire [4-1:0] node31643;
	wire [4-1:0] node31646;
	wire [4-1:0] node31649;
	wire [4-1:0] node31650;
	wire [4-1:0] node31651;
	wire [4-1:0] node31654;
	wire [4-1:0] node31657;
	wire [4-1:0] node31658;
	wire [4-1:0] node31661;
	wire [4-1:0] node31664;
	wire [4-1:0] node31665;
	wire [4-1:0] node31666;
	wire [4-1:0] node31667;
	wire [4-1:0] node31668;
	wire [4-1:0] node31671;
	wire [4-1:0] node31673;
	wire [4-1:0] node31676;
	wire [4-1:0] node31677;
	wire [4-1:0] node31680;
	wire [4-1:0] node31682;
	wire [4-1:0] node31685;
	wire [4-1:0] node31686;
	wire [4-1:0] node31687;
	wire [4-1:0] node31690;
	wire [4-1:0] node31692;
	wire [4-1:0] node31695;
	wire [4-1:0] node31696;
	wire [4-1:0] node31699;
	wire [4-1:0] node31701;
	wire [4-1:0] node31704;
	wire [4-1:0] node31705;
	wire [4-1:0] node31706;
	wire [4-1:0] node31707;
	wire [4-1:0] node31711;
	wire [4-1:0] node31712;
	wire [4-1:0] node31713;
	wire [4-1:0] node31714;
	wire [4-1:0] node31717;
	wire [4-1:0] node31720;
	wire [4-1:0] node31721;
	wire [4-1:0] node31724;
	wire [4-1:0] node31727;
	wire [4-1:0] node31728;
	wire [4-1:0] node31731;
	wire [4-1:0] node31734;
	wire [4-1:0] node31735;
	wire [4-1:0] node31736;
	wire [4-1:0] node31737;
	wire [4-1:0] node31738;
	wire [4-1:0] node31741;
	wire [4-1:0] node31744;
	wire [4-1:0] node31745;
	wire [4-1:0] node31749;
	wire [4-1:0] node31750;
	wire [4-1:0] node31753;
	wire [4-1:0] node31756;
	wire [4-1:0] node31757;
	wire [4-1:0] node31758;
	wire [4-1:0] node31761;
	wire [4-1:0] node31764;
	wire [4-1:0] node31765;
	wire [4-1:0] node31768;
	wire [4-1:0] node31771;
	wire [4-1:0] node31772;
	wire [4-1:0] node31773;
	wire [4-1:0] node31774;
	wire [4-1:0] node31775;
	wire [4-1:0] node31776;
	wire [4-1:0] node31777;
	wire [4-1:0] node31778;
	wire [4-1:0] node31779;
	wire [4-1:0] node31780;
	wire [4-1:0] node31783;
	wire [4-1:0] node31786;
	wire [4-1:0] node31788;
	wire [4-1:0] node31791;
	wire [4-1:0] node31792;
	wire [4-1:0] node31793;
	wire [4-1:0] node31796;
	wire [4-1:0] node31799;
	wire [4-1:0] node31800;
	wire [4-1:0] node31804;
	wire [4-1:0] node31805;
	wire [4-1:0] node31806;
	wire [4-1:0] node31809;
	wire [4-1:0] node31812;
	wire [4-1:0] node31815;
	wire [4-1:0] node31816;
	wire [4-1:0] node31817;
	wire [4-1:0] node31818;
	wire [4-1:0] node31819;
	wire [4-1:0] node31824;
	wire [4-1:0] node31825;
	wire [4-1:0] node31827;
	wire [4-1:0] node31830;
	wire [4-1:0] node31831;
	wire [4-1:0] node31835;
	wire [4-1:0] node31836;
	wire [4-1:0] node31837;
	wire [4-1:0] node31838;
	wire [4-1:0] node31841;
	wire [4-1:0] node31845;
	wire [4-1:0] node31846;
	wire [4-1:0] node31848;
	wire [4-1:0] node31851;
	wire [4-1:0] node31852;
	wire [4-1:0] node31856;
	wire [4-1:0] node31857;
	wire [4-1:0] node31858;
	wire [4-1:0] node31859;
	wire [4-1:0] node31860;
	wire [4-1:0] node31863;
	wire [4-1:0] node31866;
	wire [4-1:0] node31867;
	wire [4-1:0] node31868;
	wire [4-1:0] node31872;
	wire [4-1:0] node31873;
	wire [4-1:0] node31876;
	wire [4-1:0] node31879;
	wire [4-1:0] node31880;
	wire [4-1:0] node31881;
	wire [4-1:0] node31884;
	wire [4-1:0] node31887;
	wire [4-1:0] node31888;
	wire [4-1:0] node31891;
	wire [4-1:0] node31894;
	wire [4-1:0] node31895;
	wire [4-1:0] node31896;
	wire [4-1:0] node31898;
	wire [4-1:0] node31901;
	wire [4-1:0] node31902;
	wire [4-1:0] node31905;
	wire [4-1:0] node31908;
	wire [4-1:0] node31909;
	wire [4-1:0] node31910;
	wire [4-1:0] node31913;
	wire [4-1:0] node31916;
	wire [4-1:0] node31917;
	wire [4-1:0] node31918;
	wire [4-1:0] node31922;
	wire [4-1:0] node31925;
	wire [4-1:0] node31926;
	wire [4-1:0] node31927;
	wire [4-1:0] node31928;
	wire [4-1:0] node31929;
	wire [4-1:0] node31930;
	wire [4-1:0] node31933;
	wire [4-1:0] node31934;
	wire [4-1:0] node31938;
	wire [4-1:0] node31941;
	wire [4-1:0] node31942;
	wire [4-1:0] node31943;
	wire [4-1:0] node31944;
	wire [4-1:0] node31948;
	wire [4-1:0] node31949;
	wire [4-1:0] node31953;
	wire [4-1:0] node31954;
	wire [4-1:0] node31957;
	wire [4-1:0] node31960;
	wire [4-1:0] node31961;
	wire [4-1:0] node31962;
	wire [4-1:0] node31963;
	wire [4-1:0] node31965;
	wire [4-1:0] node31968;
	wire [4-1:0] node31970;
	wire [4-1:0] node31974;
	wire [4-1:0] node31975;
	wire [4-1:0] node31976;
	wire [4-1:0] node31977;
	wire [4-1:0] node31981;
	wire [4-1:0] node31983;
	wire [4-1:0] node31987;
	wire [4-1:0] node31988;
	wire [4-1:0] node31989;
	wire [4-1:0] node31990;
	wire [4-1:0] node31992;
	wire [4-1:0] node31995;
	wire [4-1:0] node31997;
	wire [4-1:0] node32000;
	wire [4-1:0] node32001;
	wire [4-1:0] node32004;
	wire [4-1:0] node32005;
	wire [4-1:0] node32009;
	wire [4-1:0] node32010;
	wire [4-1:0] node32011;
	wire [4-1:0] node32012;
	wire [4-1:0] node32015;
	wire [4-1:0] node32018;
	wire [4-1:0] node32019;
	wire [4-1:0] node32020;
	wire [4-1:0] node32023;
	wire [4-1:0] node32026;
	wire [4-1:0] node32027;
	wire [4-1:0] node32030;
	wire [4-1:0] node32033;
	wire [4-1:0] node32034;
	wire [4-1:0] node32036;
	wire [4-1:0] node32039;
	wire [4-1:0] node32040;
	wire [4-1:0] node32043;
	wire [4-1:0] node32046;
	wire [4-1:0] node32047;
	wire [4-1:0] node32048;
	wire [4-1:0] node32049;
	wire [4-1:0] node32050;
	wire [4-1:0] node32051;
	wire [4-1:0] node32052;
	wire [4-1:0] node32055;
	wire [4-1:0] node32056;
	wire [4-1:0] node32060;
	wire [4-1:0] node32061;
	wire [4-1:0] node32062;
	wire [4-1:0] node32066;
	wire [4-1:0] node32067;
	wire [4-1:0] node32071;
	wire [4-1:0] node32072;
	wire [4-1:0] node32073;
	wire [4-1:0] node32074;
	wire [4-1:0] node32077;
	wire [4-1:0] node32080;
	wire [4-1:0] node32081;
	wire [4-1:0] node32085;
	wire [4-1:0] node32088;
	wire [4-1:0] node32089;
	wire [4-1:0] node32090;
	wire [4-1:0] node32092;
	wire [4-1:0] node32095;
	wire [4-1:0] node32096;
	wire [4-1:0] node32099;
	wire [4-1:0] node32102;
	wire [4-1:0] node32103;
	wire [4-1:0] node32105;
	wire [4-1:0] node32108;
	wire [4-1:0] node32111;
	wire [4-1:0] node32112;
	wire [4-1:0] node32113;
	wire [4-1:0] node32114;
	wire [4-1:0] node32115;
	wire [4-1:0] node32116;
	wire [4-1:0] node32119;
	wire [4-1:0] node32123;
	wire [4-1:0] node32124;
	wire [4-1:0] node32128;
	wire [4-1:0] node32129;
	wire [4-1:0] node32130;
	wire [4-1:0] node32131;
	wire [4-1:0] node32134;
	wire [4-1:0] node32137;
	wire [4-1:0] node32140;
	wire [4-1:0] node32141;
	wire [4-1:0] node32145;
	wire [4-1:0] node32146;
	wire [4-1:0] node32147;
	wire [4-1:0] node32148;
	wire [4-1:0] node32149;
	wire [4-1:0] node32152;
	wire [4-1:0] node32155;
	wire [4-1:0] node32156;
	wire [4-1:0] node32160;
	wire [4-1:0] node32162;
	wire [4-1:0] node32165;
	wire [4-1:0] node32166;
	wire [4-1:0] node32167;
	wire [4-1:0] node32168;
	wire [4-1:0] node32173;
	wire [4-1:0] node32174;
	wire [4-1:0] node32175;
	wire [4-1:0] node32180;
	wire [4-1:0] node32181;
	wire [4-1:0] node32182;
	wire [4-1:0] node32183;
	wire [4-1:0] node32184;
	wire [4-1:0] node32185;
	wire [4-1:0] node32186;
	wire [4-1:0] node32190;
	wire [4-1:0] node32193;
	wire [4-1:0] node32194;
	wire [4-1:0] node32195;
	wire [4-1:0] node32198;
	wire [4-1:0] node32201;
	wire [4-1:0] node32202;
	wire [4-1:0] node32205;
	wire [4-1:0] node32208;
	wire [4-1:0] node32209;
	wire [4-1:0] node32210;
	wire [4-1:0] node32213;
	wire [4-1:0] node32216;
	wire [4-1:0] node32219;
	wire [4-1:0] node32220;
	wire [4-1:0] node32221;
	wire [4-1:0] node32223;
	wire [4-1:0] node32226;
	wire [4-1:0] node32229;
	wire [4-1:0] node32230;
	wire [4-1:0] node32232;
	wire [4-1:0] node32235;
	wire [4-1:0] node32236;
	wire [4-1:0] node32239;
	wire [4-1:0] node32242;
	wire [4-1:0] node32243;
	wire [4-1:0] node32244;
	wire [4-1:0] node32245;
	wire [4-1:0] node32246;
	wire [4-1:0] node32247;
	wire [4-1:0] node32251;
	wire [4-1:0] node32252;
	wire [4-1:0] node32256;
	wire [4-1:0] node32257;
	wire [4-1:0] node32261;
	wire [4-1:0] node32262;
	wire [4-1:0] node32263;
	wire [4-1:0] node32266;
	wire [4-1:0] node32269;
	wire [4-1:0] node32270;
	wire [4-1:0] node32273;
	wire [4-1:0] node32276;
	wire [4-1:0] node32277;
	wire [4-1:0] node32278;
	wire [4-1:0] node32279;
	wire [4-1:0] node32282;
	wire [4-1:0] node32283;
	wire [4-1:0] node32287;
	wire [4-1:0] node32288;
	wire [4-1:0] node32289;
	wire [4-1:0] node32292;
	wire [4-1:0] node32295;
	wire [4-1:0] node32296;
	wire [4-1:0] node32299;
	wire [4-1:0] node32302;
	wire [4-1:0] node32303;
	wire [4-1:0] node32305;
	wire [4-1:0] node32306;
	wire [4-1:0] node32310;
	wire [4-1:0] node32313;
	wire [4-1:0] node32314;
	wire [4-1:0] node32315;
	wire [4-1:0] node32316;
	wire [4-1:0] node32317;
	wire [4-1:0] node32318;
	wire [4-1:0] node32319;
	wire [4-1:0] node32320;
	wire [4-1:0] node32321;
	wire [4-1:0] node32325;
	wire [4-1:0] node32328;
	wire [4-1:0] node32330;
	wire [4-1:0] node32332;
	wire [4-1:0] node32335;
	wire [4-1:0] node32336;
	wire [4-1:0] node32337;
	wire [4-1:0] node32338;
	wire [4-1:0] node32342;
	wire [4-1:0] node32343;
	wire [4-1:0] node32347;
	wire [4-1:0] node32348;
	wire [4-1:0] node32350;
	wire [4-1:0] node32354;
	wire [4-1:0] node32355;
	wire [4-1:0] node32356;
	wire [4-1:0] node32357;
	wire [4-1:0] node32358;
	wire [4-1:0] node32363;
	wire [4-1:0] node32364;
	wire [4-1:0] node32365;
	wire [4-1:0] node32368;
	wire [4-1:0] node32372;
	wire [4-1:0] node32373;
	wire [4-1:0] node32374;
	wire [4-1:0] node32375;
	wire [4-1:0] node32378;
	wire [4-1:0] node32381;
	wire [4-1:0] node32382;
	wire [4-1:0] node32385;
	wire [4-1:0] node32388;
	wire [4-1:0] node32389;
	wire [4-1:0] node32392;
	wire [4-1:0] node32395;
	wire [4-1:0] node32396;
	wire [4-1:0] node32397;
	wire [4-1:0] node32398;
	wire [4-1:0] node32399;
	wire [4-1:0] node32401;
	wire [4-1:0] node32404;
	wire [4-1:0] node32405;
	wire [4-1:0] node32408;
	wire [4-1:0] node32411;
	wire [4-1:0] node32412;
	wire [4-1:0] node32415;
	wire [4-1:0] node32418;
	wire [4-1:0] node32419;
	wire [4-1:0] node32420;
	wire [4-1:0] node32421;
	wire [4-1:0] node32424;
	wire [4-1:0] node32429;
	wire [4-1:0] node32430;
	wire [4-1:0] node32431;
	wire [4-1:0] node32432;
	wire [4-1:0] node32436;
	wire [4-1:0] node32437;
	wire [4-1:0] node32441;
	wire [4-1:0] node32442;
	wire [4-1:0] node32443;
	wire [4-1:0] node32447;
	wire [4-1:0] node32448;
	wire [4-1:0] node32452;
	wire [4-1:0] node32453;
	wire [4-1:0] node32454;
	wire [4-1:0] node32455;
	wire [4-1:0] node32456;
	wire [4-1:0] node32457;
	wire [4-1:0] node32460;
	wire [4-1:0] node32463;
	wire [4-1:0] node32464;
	wire [4-1:0] node32465;
	wire [4-1:0] node32468;
	wire [4-1:0] node32471;
	wire [4-1:0] node32472;
	wire [4-1:0] node32475;
	wire [4-1:0] node32478;
	wire [4-1:0] node32479;
	wire [4-1:0] node32480;
	wire [4-1:0] node32482;
	wire [4-1:0] node32485;
	wire [4-1:0] node32486;
	wire [4-1:0] node32490;
	wire [4-1:0] node32492;
	wire [4-1:0] node32493;
	wire [4-1:0] node32496;
	wire [4-1:0] node32499;
	wire [4-1:0] node32500;
	wire [4-1:0] node32501;
	wire [4-1:0] node32503;
	wire [4-1:0] node32504;
	wire [4-1:0] node32508;
	wire [4-1:0] node32509;
	wire [4-1:0] node32510;
	wire [4-1:0] node32513;
	wire [4-1:0] node32517;
	wire [4-1:0] node32518;
	wire [4-1:0] node32519;
	wire [4-1:0] node32523;
	wire [4-1:0] node32524;
	wire [4-1:0] node32528;
	wire [4-1:0] node32529;
	wire [4-1:0] node32530;
	wire [4-1:0] node32531;
	wire [4-1:0] node32533;
	wire [4-1:0] node32536;
	wire [4-1:0] node32537;
	wire [4-1:0] node32538;
	wire [4-1:0] node32541;
	wire [4-1:0] node32544;
	wire [4-1:0] node32545;
	wire [4-1:0] node32548;
	wire [4-1:0] node32551;
	wire [4-1:0] node32552;
	wire [4-1:0] node32553;
	wire [4-1:0] node32555;
	wire [4-1:0] node32558;
	wire [4-1:0] node32559;
	wire [4-1:0] node32563;
	wire [4-1:0] node32564;
	wire [4-1:0] node32567;
	wire [4-1:0] node32570;
	wire [4-1:0] node32571;
	wire [4-1:0] node32572;
	wire [4-1:0] node32573;
	wire [4-1:0] node32574;
	wire [4-1:0] node32578;
	wire [4-1:0] node32579;
	wire [4-1:0] node32583;
	wire [4-1:0] node32584;
	wire [4-1:0] node32585;
	wire [4-1:0] node32588;
	wire [4-1:0] node32591;
	wire [4-1:0] node32594;
	wire [4-1:0] node32595;
	wire [4-1:0] node32596;
	wire [4-1:0] node32600;
	wire [4-1:0] node32603;
	wire [4-1:0] node32604;
	wire [4-1:0] node32605;
	wire [4-1:0] node32606;
	wire [4-1:0] node32607;
	wire [4-1:0] node32608;
	wire [4-1:0] node32609;
	wire [4-1:0] node32610;
	wire [4-1:0] node32613;
	wire [4-1:0] node32616;
	wire [4-1:0] node32617;
	wire [4-1:0] node32620;
	wire [4-1:0] node32623;
	wire [4-1:0] node32624;
	wire [4-1:0] node32627;
	wire [4-1:0] node32630;
	wire [4-1:0] node32631;
	wire [4-1:0] node32632;
	wire [4-1:0] node32634;
	wire [4-1:0] node32637;
	wire [4-1:0] node32640;
	wire [4-1:0] node32641;
	wire [4-1:0] node32643;
	wire [4-1:0] node32646;
	wire [4-1:0] node32647;
	wire [4-1:0] node32651;
	wire [4-1:0] node32652;
	wire [4-1:0] node32653;
	wire [4-1:0] node32654;
	wire [4-1:0] node32657;
	wire [4-1:0] node32661;
	wire [4-1:0] node32662;
	wire [4-1:0] node32663;
	wire [4-1:0] node32667;
	wire [4-1:0] node32668;
	wire [4-1:0] node32672;
	wire [4-1:0] node32673;
	wire [4-1:0] node32674;
	wire [4-1:0] node32675;
	wire [4-1:0] node32676;
	wire [4-1:0] node32678;
	wire [4-1:0] node32681;
	wire [4-1:0] node32682;
	wire [4-1:0] node32685;
	wire [4-1:0] node32688;
	wire [4-1:0] node32689;
	wire [4-1:0] node32693;
	wire [4-1:0] node32694;
	wire [4-1:0] node32695;
	wire [4-1:0] node32697;
	wire [4-1:0] node32700;
	wire [4-1:0] node32701;
	wire [4-1:0] node32706;
	wire [4-1:0] node32707;
	wire [4-1:0] node32708;
	wire [4-1:0] node32709;
	wire [4-1:0] node32712;
	wire [4-1:0] node32715;
	wire [4-1:0] node32716;
	wire [4-1:0] node32719;
	wire [4-1:0] node32722;
	wire [4-1:0] node32725;
	wire [4-1:0] node32726;
	wire [4-1:0] node32727;
	wire [4-1:0] node32728;
	wire [4-1:0] node32729;
	wire [4-1:0] node32730;
	wire [4-1:0] node32732;
	wire [4-1:0] node32735;
	wire [4-1:0] node32736;
	wire [4-1:0] node32739;
	wire [4-1:0] node32742;
	wire [4-1:0] node32743;
	wire [4-1:0] node32746;
	wire [4-1:0] node32749;
	wire [4-1:0] node32750;
	wire [4-1:0] node32751;
	wire [4-1:0] node32752;
	wire [4-1:0] node32756;
	wire [4-1:0] node32759;
	wire [4-1:0] node32760;
	wire [4-1:0] node32763;
	wire [4-1:0] node32765;
	wire [4-1:0] node32768;
	wire [4-1:0] node32769;
	wire [4-1:0] node32770;
	wire [4-1:0] node32771;
	wire [4-1:0] node32774;
	wire [4-1:0] node32778;
	wire [4-1:0] node32779;
	wire [4-1:0] node32780;
	wire [4-1:0] node32784;
	wire [4-1:0] node32785;
	wire [4-1:0] node32789;
	wire [4-1:0] node32790;
	wire [4-1:0] node32791;
	wire [4-1:0] node32792;
	wire [4-1:0] node32793;
	wire [4-1:0] node32795;
	wire [4-1:0] node32798;
	wire [4-1:0] node32799;
	wire [4-1:0] node32803;
	wire [4-1:0] node32804;
	wire [4-1:0] node32807;
	wire [4-1:0] node32810;
	wire [4-1:0] node32811;
	wire [4-1:0] node32812;
	wire [4-1:0] node32813;
	wire [4-1:0] node32817;
	wire [4-1:0] node32819;
	wire [4-1:0] node32823;
	wire [4-1:0] node32824;
	wire [4-1:0] node32825;
	wire [4-1:0] node32826;
	wire [4-1:0] node32829;
	wire [4-1:0] node32833;
	wire [4-1:0] node32834;
	wire [4-1:0] node32835;
	wire [4-1:0] node32838;
	wire [4-1:0] node32842;
	wire [4-1:0] node32843;
	wire [4-1:0] node32844;
	wire [4-1:0] node32845;
	wire [4-1:0] node32846;
	wire [4-1:0] node32847;
	wire [4-1:0] node32848;
	wire [4-1:0] node32849;
	wire [4-1:0] node32850;
	wire [4-1:0] node32851;
	wire [4-1:0] node32852;
	wire [4-1:0] node32854;
	wire [4-1:0] node32857;
	wire [4-1:0] node32859;
	wire [4-1:0] node32862;
	wire [4-1:0] node32863;
	wire [4-1:0] node32866;
	wire [4-1:0] node32867;
	wire [4-1:0] node32871;
	wire [4-1:0] node32872;
	wire [4-1:0] node32873;
	wire [4-1:0] node32874;
	wire [4-1:0] node32879;
	wire [4-1:0] node32880;
	wire [4-1:0] node32882;
	wire [4-1:0] node32885;
	wire [4-1:0] node32887;
	wire [4-1:0] node32890;
	wire [4-1:0] node32891;
	wire [4-1:0] node32892;
	wire [4-1:0] node32893;
	wire [4-1:0] node32896;
	wire [4-1:0] node32899;
	wire [4-1:0] node32900;
	wire [4-1:0] node32903;
	wire [4-1:0] node32906;
	wire [4-1:0] node32907;
	wire [4-1:0] node32909;
	wire [4-1:0] node32911;
	wire [4-1:0] node32914;
	wire [4-1:0] node32915;
	wire [4-1:0] node32916;
	wire [4-1:0] node32920;
	wire [4-1:0] node32921;
	wire [4-1:0] node32925;
	wire [4-1:0] node32926;
	wire [4-1:0] node32927;
	wire [4-1:0] node32928;
	wire [4-1:0] node32929;
	wire [4-1:0] node32932;
	wire [4-1:0] node32935;
	wire [4-1:0] node32936;
	wire [4-1:0] node32938;
	wire [4-1:0] node32941;
	wire [4-1:0] node32942;
	wire [4-1:0] node32946;
	wire [4-1:0] node32947;
	wire [4-1:0] node32948;
	wire [4-1:0] node32949;
	wire [4-1:0] node32953;
	wire [4-1:0] node32955;
	wire [4-1:0] node32958;
	wire [4-1:0] node32959;
	wire [4-1:0] node32961;
	wire [4-1:0] node32964;
	wire [4-1:0] node32965;
	wire [4-1:0] node32969;
	wire [4-1:0] node32970;
	wire [4-1:0] node32971;
	wire [4-1:0] node32972;
	wire [4-1:0] node32974;
	wire [4-1:0] node32977;
	wire [4-1:0] node32980;
	wire [4-1:0] node32981;
	wire [4-1:0] node32983;
	wire [4-1:0] node32986;
	wire [4-1:0] node32989;
	wire [4-1:0] node32990;
	wire [4-1:0] node32991;
	wire [4-1:0] node32994;
	wire [4-1:0] node32996;
	wire [4-1:0] node32999;
	wire [4-1:0] node33000;
	wire [4-1:0] node33001;
	wire [4-1:0] node33005;
	wire [4-1:0] node33006;
	wire [4-1:0] node33010;
	wire [4-1:0] node33011;
	wire [4-1:0] node33012;
	wire [4-1:0] node33013;
	wire [4-1:0] node33014;
	wire [4-1:0] node33015;
	wire [4-1:0] node33017;
	wire [4-1:0] node33021;
	wire [4-1:0] node33022;
	wire [4-1:0] node33025;
	wire [4-1:0] node33028;
	wire [4-1:0] node33029;
	wire [4-1:0] node33030;
	wire [4-1:0] node33031;
	wire [4-1:0] node33036;
	wire [4-1:0] node33037;
	wire [4-1:0] node33038;
	wire [4-1:0] node33043;
	wire [4-1:0] node33044;
	wire [4-1:0] node33045;
	wire [4-1:0] node33046;
	wire [4-1:0] node33049;
	wire [4-1:0] node33050;
	wire [4-1:0] node33054;
	wire [4-1:0] node33055;
	wire [4-1:0] node33058;
	wire [4-1:0] node33059;
	wire [4-1:0] node33063;
	wire [4-1:0] node33064;
	wire [4-1:0] node33066;
	wire [4-1:0] node33069;
	wire [4-1:0] node33070;
	wire [4-1:0] node33073;
	wire [4-1:0] node33074;
	wire [4-1:0] node33078;
	wire [4-1:0] node33079;
	wire [4-1:0] node33080;
	wire [4-1:0] node33081;
	wire [4-1:0] node33083;
	wire [4-1:0] node33086;
	wire [4-1:0] node33087;
	wire [4-1:0] node33088;
	wire [4-1:0] node33092;
	wire [4-1:0] node33093;
	wire [4-1:0] node33096;
	wire [4-1:0] node33099;
	wire [4-1:0] node33100;
	wire [4-1:0] node33101;
	wire [4-1:0] node33102;
	wire [4-1:0] node33105;
	wire [4-1:0] node33108;
	wire [4-1:0] node33109;
	wire [4-1:0] node33112;
	wire [4-1:0] node33115;
	wire [4-1:0] node33116;
	wire [4-1:0] node33119;
	wire [4-1:0] node33120;
	wire [4-1:0] node33123;
	wire [4-1:0] node33126;
	wire [4-1:0] node33127;
	wire [4-1:0] node33128;
	wire [4-1:0] node33129;
	wire [4-1:0] node33130;
	wire [4-1:0] node33134;
	wire [4-1:0] node33136;
	wire [4-1:0] node33139;
	wire [4-1:0] node33140;
	wire [4-1:0] node33142;
	wire [4-1:0] node33145;
	wire [4-1:0] node33146;
	wire [4-1:0] node33150;
	wire [4-1:0] node33151;
	wire [4-1:0] node33152;
	wire [4-1:0] node33153;
	wire [4-1:0] node33157;
	wire [4-1:0] node33160;
	wire [4-1:0] node33161;
	wire [4-1:0] node33162;
	wire [4-1:0] node33165;
	wire [4-1:0] node33168;
	wire [4-1:0] node33169;
	wire [4-1:0] node33173;
	wire [4-1:0] node33174;
	wire [4-1:0] node33175;
	wire [4-1:0] node33176;
	wire [4-1:0] node33177;
	wire [4-1:0] node33178;
	wire [4-1:0] node33179;
	wire [4-1:0] node33180;
	wire [4-1:0] node33184;
	wire [4-1:0] node33187;
	wire [4-1:0] node33188;
	wire [4-1:0] node33189;
	wire [4-1:0] node33193;
	wire [4-1:0] node33194;
	wire [4-1:0] node33198;
	wire [4-1:0] node33199;
	wire [4-1:0] node33200;
	wire [4-1:0] node33201;
	wire [4-1:0] node33205;
	wire [4-1:0] node33206;
	wire [4-1:0] node33210;
	wire [4-1:0] node33211;
	wire [4-1:0] node33212;
	wire [4-1:0] node33216;
	wire [4-1:0] node33219;
	wire [4-1:0] node33220;
	wire [4-1:0] node33221;
	wire [4-1:0] node33222;
	wire [4-1:0] node33225;
	wire [4-1:0] node33226;
	wire [4-1:0] node33230;
	wire [4-1:0] node33231;
	wire [4-1:0] node33233;
	wire [4-1:0] node33236;
	wire [4-1:0] node33238;
	wire [4-1:0] node33241;
	wire [4-1:0] node33242;
	wire [4-1:0] node33244;
	wire [4-1:0] node33245;
	wire [4-1:0] node33248;
	wire [4-1:0] node33251;
	wire [4-1:0] node33253;
	wire [4-1:0] node33255;
	wire [4-1:0] node33258;
	wire [4-1:0] node33259;
	wire [4-1:0] node33260;
	wire [4-1:0] node33261;
	wire [4-1:0] node33262;
	wire [4-1:0] node33265;
	wire [4-1:0] node33267;
	wire [4-1:0] node33270;
	wire [4-1:0] node33271;
	wire [4-1:0] node33272;
	wire [4-1:0] node33276;
	wire [4-1:0] node33279;
	wire [4-1:0] node33280;
	wire [4-1:0] node33282;
	wire [4-1:0] node33283;
	wire [4-1:0] node33288;
	wire [4-1:0] node33289;
	wire [4-1:0] node33290;
	wire [4-1:0] node33291;
	wire [4-1:0] node33292;
	wire [4-1:0] node33296;
	wire [4-1:0] node33298;
	wire [4-1:0] node33301;
	wire [4-1:0] node33302;
	wire [4-1:0] node33303;
	wire [4-1:0] node33307;
	wire [4-1:0] node33310;
	wire [4-1:0] node33311;
	wire [4-1:0] node33312;
	wire [4-1:0] node33313;
	wire [4-1:0] node33317;
	wire [4-1:0] node33319;
	wire [4-1:0] node33322;
	wire [4-1:0] node33323;
	wire [4-1:0] node33324;
	wire [4-1:0] node33327;
	wire [4-1:0] node33331;
	wire [4-1:0] node33332;
	wire [4-1:0] node33333;
	wire [4-1:0] node33334;
	wire [4-1:0] node33335;
	wire [4-1:0] node33337;
	wire [4-1:0] node33339;
	wire [4-1:0] node33342;
	wire [4-1:0] node33343;
	wire [4-1:0] node33344;
	wire [4-1:0] node33348;
	wire [4-1:0] node33349;
	wire [4-1:0] node33353;
	wire [4-1:0] node33354;
	wire [4-1:0] node33355;
	wire [4-1:0] node33356;
	wire [4-1:0] node33360;
	wire [4-1:0] node33362;
	wire [4-1:0] node33365;
	wire [4-1:0] node33367;
	wire [4-1:0] node33368;
	wire [4-1:0] node33372;
	wire [4-1:0] node33373;
	wire [4-1:0] node33374;
	wire [4-1:0] node33375;
	wire [4-1:0] node33376;
	wire [4-1:0] node33380;
	wire [4-1:0] node33381;
	wire [4-1:0] node33384;
	wire [4-1:0] node33387;
	wire [4-1:0] node33388;
	wire [4-1:0] node33389;
	wire [4-1:0] node33392;
	wire [4-1:0] node33395;
	wire [4-1:0] node33396;
	wire [4-1:0] node33399;
	wire [4-1:0] node33402;
	wire [4-1:0] node33403;
	wire [4-1:0] node33404;
	wire [4-1:0] node33407;
	wire [4-1:0] node33409;
	wire [4-1:0] node33412;
	wire [4-1:0] node33413;
	wire [4-1:0] node33414;
	wire [4-1:0] node33418;
	wire [4-1:0] node33421;
	wire [4-1:0] node33422;
	wire [4-1:0] node33423;
	wire [4-1:0] node33424;
	wire [4-1:0] node33426;
	wire [4-1:0] node33428;
	wire [4-1:0] node33431;
	wire [4-1:0] node33432;
	wire [4-1:0] node33434;
	wire [4-1:0] node33437;
	wire [4-1:0] node33438;
	wire [4-1:0] node33442;
	wire [4-1:0] node33443;
	wire [4-1:0] node33444;
	wire [4-1:0] node33447;
	wire [4-1:0] node33448;
	wire [4-1:0] node33452;
	wire [4-1:0] node33453;
	wire [4-1:0] node33455;
	wire [4-1:0] node33458;
	wire [4-1:0] node33460;
	wire [4-1:0] node33463;
	wire [4-1:0] node33464;
	wire [4-1:0] node33465;
	wire [4-1:0] node33467;
	wire [4-1:0] node33470;
	wire [4-1:0] node33471;
	wire [4-1:0] node33474;
	wire [4-1:0] node33477;
	wire [4-1:0] node33478;
	wire [4-1:0] node33479;
	wire [4-1:0] node33483;
	wire [4-1:0] node33485;
	wire [4-1:0] node33486;
	wire [4-1:0] node33490;
	wire [4-1:0] node33491;
	wire [4-1:0] node33492;
	wire [4-1:0] node33493;
	wire [4-1:0] node33494;
	wire [4-1:0] node33495;
	wire [4-1:0] node33496;
	wire [4-1:0] node33497;
	wire [4-1:0] node33499;
	wire [4-1:0] node33502;
	wire [4-1:0] node33505;
	wire [4-1:0] node33506;
	wire [4-1:0] node33508;
	wire [4-1:0] node33511;
	wire [4-1:0] node33514;
	wire [4-1:0] node33515;
	wire [4-1:0] node33516;
	wire [4-1:0] node33518;
	wire [4-1:0] node33521;
	wire [4-1:0] node33523;
	wire [4-1:0] node33526;
	wire [4-1:0] node33527;
	wire [4-1:0] node33530;
	wire [4-1:0] node33532;
	wire [4-1:0] node33535;
	wire [4-1:0] node33536;
	wire [4-1:0] node33537;
	wire [4-1:0] node33538;
	wire [4-1:0] node33539;
	wire [4-1:0] node33543;
	wire [4-1:0] node33546;
	wire [4-1:0] node33547;
	wire [4-1:0] node33548;
	wire [4-1:0] node33551;
	wire [4-1:0] node33554;
	wire [4-1:0] node33555;
	wire [4-1:0] node33559;
	wire [4-1:0] node33560;
	wire [4-1:0] node33561;
	wire [4-1:0] node33562;
	wire [4-1:0] node33566;
	wire [4-1:0] node33569;
	wire [4-1:0] node33570;
	wire [4-1:0] node33572;
	wire [4-1:0] node33575;
	wire [4-1:0] node33578;
	wire [4-1:0] node33579;
	wire [4-1:0] node33580;
	wire [4-1:0] node33581;
	wire [4-1:0] node33582;
	wire [4-1:0] node33583;
	wire [4-1:0] node33587;
	wire [4-1:0] node33588;
	wire [4-1:0] node33592;
	wire [4-1:0] node33593;
	wire [4-1:0] node33596;
	wire [4-1:0] node33597;
	wire [4-1:0] node33601;
	wire [4-1:0] node33602;
	wire [4-1:0] node33603;
	wire [4-1:0] node33604;
	wire [4-1:0] node33608;
	wire [4-1:0] node33609;
	wire [4-1:0] node33612;
	wire [4-1:0] node33615;
	wire [4-1:0] node33616;
	wire [4-1:0] node33617;
	wire [4-1:0] node33621;
	wire [4-1:0] node33622;
	wire [4-1:0] node33625;
	wire [4-1:0] node33628;
	wire [4-1:0] node33629;
	wire [4-1:0] node33630;
	wire [4-1:0] node33631;
	wire [4-1:0] node33634;
	wire [4-1:0] node33637;
	wire [4-1:0] node33638;
	wire [4-1:0] node33639;
	wire [4-1:0] node33642;
	wire [4-1:0] node33645;
	wire [4-1:0] node33646;
	wire [4-1:0] node33650;
	wire [4-1:0] node33651;
	wire [4-1:0] node33652;
	wire [4-1:0] node33653;
	wire [4-1:0] node33656;
	wire [4-1:0] node33659;
	wire [4-1:0] node33661;
	wire [4-1:0] node33664;
	wire [4-1:0] node33665;
	wire [4-1:0] node33667;
	wire [4-1:0] node33670;
	wire [4-1:0] node33671;
	wire [4-1:0] node33675;
	wire [4-1:0] node33676;
	wire [4-1:0] node33677;
	wire [4-1:0] node33678;
	wire [4-1:0] node33679;
	wire [4-1:0] node33680;
	wire [4-1:0] node33681;
	wire [4-1:0] node33684;
	wire [4-1:0] node33687;
	wire [4-1:0] node33688;
	wire [4-1:0] node33692;
	wire [4-1:0] node33693;
	wire [4-1:0] node33694;
	wire [4-1:0] node33698;
	wire [4-1:0] node33699;
	wire [4-1:0] node33703;
	wire [4-1:0] node33704;
	wire [4-1:0] node33705;
	wire [4-1:0] node33707;
	wire [4-1:0] node33710;
	wire [4-1:0] node33711;
	wire [4-1:0] node33714;
	wire [4-1:0] node33717;
	wire [4-1:0] node33718;
	wire [4-1:0] node33721;
	wire [4-1:0] node33722;
	wire [4-1:0] node33725;
	wire [4-1:0] node33728;
	wire [4-1:0] node33729;
	wire [4-1:0] node33730;
	wire [4-1:0] node33731;
	wire [4-1:0] node33732;
	wire [4-1:0] node33735;
	wire [4-1:0] node33738;
	wire [4-1:0] node33739;
	wire [4-1:0] node33742;
	wire [4-1:0] node33745;
	wire [4-1:0] node33746;
	wire [4-1:0] node33747;
	wire [4-1:0] node33751;
	wire [4-1:0] node33752;
	wire [4-1:0] node33755;
	wire [4-1:0] node33758;
	wire [4-1:0] node33759;
	wire [4-1:0] node33760;
	wire [4-1:0] node33761;
	wire [4-1:0] node33764;
	wire [4-1:0] node33767;
	wire [4-1:0] node33770;
	wire [4-1:0] node33771;
	wire [4-1:0] node33772;
	wire [4-1:0] node33775;
	wire [4-1:0] node33778;
	wire [4-1:0] node33779;
	wire [4-1:0] node33782;
	wire [4-1:0] node33785;
	wire [4-1:0] node33786;
	wire [4-1:0] node33787;
	wire [4-1:0] node33788;
	wire [4-1:0] node33789;
	wire [4-1:0] node33790;
	wire [4-1:0] node33794;
	wire [4-1:0] node33795;
	wire [4-1:0] node33798;
	wire [4-1:0] node33801;
	wire [4-1:0] node33802;
	wire [4-1:0] node33805;
	wire [4-1:0] node33806;
	wire [4-1:0] node33810;
	wire [4-1:0] node33811;
	wire [4-1:0] node33812;
	wire [4-1:0] node33815;
	wire [4-1:0] node33816;
	wire [4-1:0] node33820;
	wire [4-1:0] node33821;
	wire [4-1:0] node33822;
	wire [4-1:0] node33826;
	wire [4-1:0] node33829;
	wire [4-1:0] node33830;
	wire [4-1:0] node33831;
	wire [4-1:0] node33832;
	wire [4-1:0] node33833;
	wire [4-1:0] node33837;
	wire [4-1:0] node33839;
	wire [4-1:0] node33842;
	wire [4-1:0] node33843;
	wire [4-1:0] node33844;
	wire [4-1:0] node33848;
	wire [4-1:0] node33849;
	wire [4-1:0] node33852;
	wire [4-1:0] node33855;
	wire [4-1:0] node33856;
	wire [4-1:0] node33857;
	wire [4-1:0] node33859;
	wire [4-1:0] node33862;
	wire [4-1:0] node33864;
	wire [4-1:0] node33867;
	wire [4-1:0] node33869;
	wire [4-1:0] node33871;
	wire [4-1:0] node33874;
	wire [4-1:0] node33875;
	wire [4-1:0] node33876;
	wire [4-1:0] node33877;
	wire [4-1:0] node33878;
	wire [4-1:0] node33879;
	wire [4-1:0] node33880;
	wire [4-1:0] node33881;
	wire [4-1:0] node33884;
	wire [4-1:0] node33887;
	wire [4-1:0] node33888;
	wire [4-1:0] node33891;
	wire [4-1:0] node33894;
	wire [4-1:0] node33895;
	wire [4-1:0] node33897;
	wire [4-1:0] node33900;
	wire [4-1:0] node33901;
	wire [4-1:0] node33905;
	wire [4-1:0] node33906;
	wire [4-1:0] node33907;
	wire [4-1:0] node33908;
	wire [4-1:0] node33911;
	wire [4-1:0] node33914;
	wire [4-1:0] node33915;
	wire [4-1:0] node33918;
	wire [4-1:0] node33921;
	wire [4-1:0] node33922;
	wire [4-1:0] node33923;
	wire [4-1:0] node33926;
	wire [4-1:0] node33929;
	wire [4-1:0] node33930;
	wire [4-1:0] node33933;
	wire [4-1:0] node33936;
	wire [4-1:0] node33937;
	wire [4-1:0] node33938;
	wire [4-1:0] node33939;
	wire [4-1:0] node33940;
	wire [4-1:0] node33945;
	wire [4-1:0] node33946;
	wire [4-1:0] node33947;
	wire [4-1:0] node33950;
	wire [4-1:0] node33953;
	wire [4-1:0] node33955;
	wire [4-1:0] node33958;
	wire [4-1:0] node33959;
	wire [4-1:0] node33960;
	wire [4-1:0] node33961;
	wire [4-1:0] node33965;
	wire [4-1:0] node33967;
	wire [4-1:0] node33970;
	wire [4-1:0] node33971;
	wire [4-1:0] node33972;
	wire [4-1:0] node33976;
	wire [4-1:0] node33977;
	wire [4-1:0] node33980;
	wire [4-1:0] node33983;
	wire [4-1:0] node33984;
	wire [4-1:0] node33985;
	wire [4-1:0] node33986;
	wire [4-1:0] node33987;
	wire [4-1:0] node33988;
	wire [4-1:0] node33991;
	wire [4-1:0] node33994;
	wire [4-1:0] node33995;
	wire [4-1:0] node33998;
	wire [4-1:0] node34001;
	wire [4-1:0] node34002;
	wire [4-1:0] node34004;
	wire [4-1:0] node34007;
	wire [4-1:0] node34008;
	wire [4-1:0] node34011;
	wire [4-1:0] node34014;
	wire [4-1:0] node34015;
	wire [4-1:0] node34016;
	wire [4-1:0] node34019;
	wire [4-1:0] node34020;
	wire [4-1:0] node34024;
	wire [4-1:0] node34025;
	wire [4-1:0] node34026;
	wire [4-1:0] node34029;
	wire [4-1:0] node34032;
	wire [4-1:0] node34034;
	wire [4-1:0] node34037;
	wire [4-1:0] node34038;
	wire [4-1:0] node34039;
	wire [4-1:0] node34040;
	wire [4-1:0] node34041;
	wire [4-1:0] node34045;
	wire [4-1:0] node34046;
	wire [4-1:0] node34050;
	wire [4-1:0] node34051;
	wire [4-1:0] node34054;
	wire [4-1:0] node34056;
	wire [4-1:0] node34059;
	wire [4-1:0] node34060;
	wire [4-1:0] node34061;
	wire [4-1:0] node34062;
	wire [4-1:0] node34066;
	wire [4-1:0] node34068;
	wire [4-1:0] node34071;
	wire [4-1:0] node34072;
	wire [4-1:0] node34073;
	wire [4-1:0] node34076;
	wire [4-1:0] node34079;
	wire [4-1:0] node34080;
	wire [4-1:0] node34084;
	wire [4-1:0] node34085;
	wire [4-1:0] node34086;
	wire [4-1:0] node34087;
	wire [4-1:0] node34088;
	wire [4-1:0] node34089;
	wire [4-1:0] node34092;
	wire [4-1:0] node34094;
	wire [4-1:0] node34097;
	wire [4-1:0] node34098;
	wire [4-1:0] node34099;
	wire [4-1:0] node34103;
	wire [4-1:0] node34106;
	wire [4-1:0] node34107;
	wire [4-1:0] node34108;
	wire [4-1:0] node34110;
	wire [4-1:0] node34113;
	wire [4-1:0] node34114;
	wire [4-1:0] node34117;
	wire [4-1:0] node34120;
	wire [4-1:0] node34121;
	wire [4-1:0] node34122;
	wire [4-1:0] node34125;
	wire [4-1:0] node34128;
	wire [4-1:0] node34130;
	wire [4-1:0] node34133;
	wire [4-1:0] node34134;
	wire [4-1:0] node34135;
	wire [4-1:0] node34136;
	wire [4-1:0] node34137;
	wire [4-1:0] node34141;
	wire [4-1:0] node34142;
	wire [4-1:0] node34145;
	wire [4-1:0] node34148;
	wire [4-1:0] node34149;
	wire [4-1:0] node34152;
	wire [4-1:0] node34153;
	wire [4-1:0] node34156;
	wire [4-1:0] node34159;
	wire [4-1:0] node34160;
	wire [4-1:0] node34161;
	wire [4-1:0] node34162;
	wire [4-1:0] node34166;
	wire [4-1:0] node34169;
	wire [4-1:0] node34170;
	wire [4-1:0] node34171;
	wire [4-1:0] node34174;
	wire [4-1:0] node34177;
	wire [4-1:0] node34178;
	wire [4-1:0] node34181;
	wire [4-1:0] node34184;
	wire [4-1:0] node34185;
	wire [4-1:0] node34186;
	wire [4-1:0] node34187;
	wire [4-1:0] node34188;
	wire [4-1:0] node34189;
	wire [4-1:0] node34193;
	wire [4-1:0] node34196;
	wire [4-1:0] node34197;
	wire [4-1:0] node34200;
	wire [4-1:0] node34201;
	wire [4-1:0] node34205;
	wire [4-1:0] node34206;
	wire [4-1:0] node34207;
	wire [4-1:0] node34210;
	wire [4-1:0] node34211;
	wire [4-1:0] node34215;
	wire [4-1:0] node34216;
	wire [4-1:0] node34217;
	wire [4-1:0] node34221;
	wire [4-1:0] node34222;
	wire [4-1:0] node34226;
	wire [4-1:0] node34227;
	wire [4-1:0] node34228;
	wire [4-1:0] node34229;
	wire [4-1:0] node34231;
	wire [4-1:0] node34234;
	wire [4-1:0] node34237;
	wire [4-1:0] node34238;
	wire [4-1:0] node34241;
	wire [4-1:0] node34243;
	wire [4-1:0] node34246;
	wire [4-1:0] node34247;
	wire [4-1:0] node34248;
	wire [4-1:0] node34250;
	wire [4-1:0] node34253;
	wire [4-1:0] node34255;
	wire [4-1:0] node34258;
	wire [4-1:0] node34259;
	wire [4-1:0] node34260;
	wire [4-1:0] node34264;
	wire [4-1:0] node34266;
	wire [4-1:0] node34269;
	wire [4-1:0] node34270;
	wire [4-1:0] node34271;
	wire [4-1:0] node34272;
	wire [4-1:0] node34273;
	wire [4-1:0] node34274;
	wire [4-1:0] node34275;
	wire [4-1:0] node34276;
	wire [4-1:0] node34277;
	wire [4-1:0] node34280;
	wire [4-1:0] node34283;
	wire [4-1:0] node34284;
	wire [4-1:0] node34287;
	wire [4-1:0] node34290;
	wire [4-1:0] node34291;
	wire [4-1:0] node34292;
	wire [4-1:0] node34295;
	wire [4-1:0] node34298;
	wire [4-1:0] node34301;
	wire [4-1:0] node34302;
	wire [4-1:0] node34303;
	wire [4-1:0] node34304;
	wire [4-1:0] node34307;
	wire [4-1:0] node34310;
	wire [4-1:0] node34313;
	wire [4-1:0] node34314;
	wire [4-1:0] node34315;
	wire [4-1:0] node34318;
	wire [4-1:0] node34321;
	wire [4-1:0] node34324;
	wire [4-1:0] node34325;
	wire [4-1:0] node34326;
	wire [4-1:0] node34327;
	wire [4-1:0] node34329;
	wire [4-1:0] node34330;
	wire [4-1:0] node34333;
	wire [4-1:0] node34336;
	wire [4-1:0] node34337;
	wire [4-1:0] node34338;
	wire [4-1:0] node34342;
	wire [4-1:0] node34343;
	wire [4-1:0] node34346;
	wire [4-1:0] node34349;
	wire [4-1:0] node34350;
	wire [4-1:0] node34351;
	wire [4-1:0] node34354;
	wire [4-1:0] node34357;
	wire [4-1:0] node34358;
	wire [4-1:0] node34361;
	wire [4-1:0] node34364;
	wire [4-1:0] node34365;
	wire [4-1:0] node34366;
	wire [4-1:0] node34367;
	wire [4-1:0] node34370;
	wire [4-1:0] node34373;
	wire [4-1:0] node34375;
	wire [4-1:0] node34376;
	wire [4-1:0] node34379;
	wire [4-1:0] node34382;
	wire [4-1:0] node34383;
	wire [4-1:0] node34384;
	wire [4-1:0] node34387;
	wire [4-1:0] node34390;
	wire [4-1:0] node34391;
	wire [4-1:0] node34392;
	wire [4-1:0] node34396;
	wire [4-1:0] node34397;
	wire [4-1:0] node34400;
	wire [4-1:0] node34403;
	wire [4-1:0] node34404;
	wire [4-1:0] node34405;
	wire [4-1:0] node34406;
	wire [4-1:0] node34407;
	wire [4-1:0] node34408;
	wire [4-1:0] node34411;
	wire [4-1:0] node34414;
	wire [4-1:0] node34415;
	wire [4-1:0] node34418;
	wire [4-1:0] node34421;
	wire [4-1:0] node34422;
	wire [4-1:0] node34423;
	wire [4-1:0] node34424;
	wire [4-1:0] node34427;
	wire [4-1:0] node34430;
	wire [4-1:0] node34431;
	wire [4-1:0] node34434;
	wire [4-1:0] node34437;
	wire [4-1:0] node34438;
	wire [4-1:0] node34439;
	wire [4-1:0] node34442;
	wire [4-1:0] node34445;
	wire [4-1:0] node34447;
	wire [4-1:0] node34450;
	wire [4-1:0] node34451;
	wire [4-1:0] node34452;
	wire [4-1:0] node34453;
	wire [4-1:0] node34456;
	wire [4-1:0] node34459;
	wire [4-1:0] node34460;
	wire [4-1:0] node34463;
	wire [4-1:0] node34466;
	wire [4-1:0] node34467;
	wire [4-1:0] node34468;
	wire [4-1:0] node34472;
	wire [4-1:0] node34475;
	wire [4-1:0] node34476;
	wire [4-1:0] node34477;
	wire [4-1:0] node34478;
	wire [4-1:0] node34480;
	wire [4-1:0] node34483;
	wire [4-1:0] node34485;
	wire [4-1:0] node34488;
	wire [4-1:0] node34489;
	wire [4-1:0] node34490;
	wire [4-1:0] node34493;
	wire [4-1:0] node34496;
	wire [4-1:0] node34499;
	wire [4-1:0] node34500;
	wire [4-1:0] node34501;
	wire [4-1:0] node34502;
	wire [4-1:0] node34505;
	wire [4-1:0] node34508;
	wire [4-1:0] node34511;
	wire [4-1:0] node34512;
	wire [4-1:0] node34513;
	wire [4-1:0] node34516;
	wire [4-1:0] node34519;
	wire [4-1:0] node34522;
	wire [4-1:0] node34523;
	wire [4-1:0] node34524;
	wire [4-1:0] node34525;
	wire [4-1:0] node34526;
	wire [4-1:0] node34527;
	wire [4-1:0] node34528;
	wire [4-1:0] node34533;
	wire [4-1:0] node34534;
	wire [4-1:0] node34536;
	wire [4-1:0] node34540;
	wire [4-1:0] node34541;
	wire [4-1:0] node34542;
	wire [4-1:0] node34544;
	wire [4-1:0] node34548;
	wire [4-1:0] node34549;
	wire [4-1:0] node34550;
	wire [4-1:0] node34555;
	wire [4-1:0] node34556;
	wire [4-1:0] node34557;
	wire [4-1:0] node34558;
	wire [4-1:0] node34560;
	wire [4-1:0] node34563;
	wire [4-1:0] node34565;
	wire [4-1:0] node34568;
	wire [4-1:0] node34569;
	wire [4-1:0] node34570;
	wire [4-1:0] node34574;
	wire [4-1:0] node34576;
	wire [4-1:0] node34579;
	wire [4-1:0] node34580;
	wire [4-1:0] node34581;
	wire [4-1:0] node34582;
	wire [4-1:0] node34585;
	wire [4-1:0] node34588;
	wire [4-1:0] node34589;
	wire [4-1:0] node34593;
	wire [4-1:0] node34594;
	wire [4-1:0] node34595;
	wire [4-1:0] node34598;
	wire [4-1:0] node34601;
	wire [4-1:0] node34602;
	wire [4-1:0] node34605;
	wire [4-1:0] node34608;
	wire [4-1:0] node34609;
	wire [4-1:0] node34610;
	wire [4-1:0] node34611;
	wire [4-1:0] node34612;
	wire [4-1:0] node34613;
	wire [4-1:0] node34616;
	wire [4-1:0] node34619;
	wire [4-1:0] node34620;
	wire [4-1:0] node34621;
	wire [4-1:0] node34624;
	wire [4-1:0] node34627;
	wire [4-1:0] node34628;
	wire [4-1:0] node34631;
	wire [4-1:0] node34634;
	wire [4-1:0] node34635;
	wire [4-1:0] node34636;
	wire [4-1:0] node34637;
	wire [4-1:0] node34640;
	wire [4-1:0] node34643;
	wire [4-1:0] node34644;
	wire [4-1:0] node34647;
	wire [4-1:0] node34650;
	wire [4-1:0] node34651;
	wire [4-1:0] node34652;
	wire [4-1:0] node34655;
	wire [4-1:0] node34658;
	wire [4-1:0] node34659;
	wire [4-1:0] node34662;
	wire [4-1:0] node34665;
	wire [4-1:0] node34666;
	wire [4-1:0] node34667;
	wire [4-1:0] node34668;
	wire [4-1:0] node34669;
	wire [4-1:0] node34673;
	wire [4-1:0] node34674;
	wire [4-1:0] node34678;
	wire [4-1:0] node34680;
	wire [4-1:0] node34681;
	wire [4-1:0] node34685;
	wire [4-1:0] node34686;
	wire [4-1:0] node34687;
	wire [4-1:0] node34689;
	wire [4-1:0] node34692;
	wire [4-1:0] node34693;
	wire [4-1:0] node34696;
	wire [4-1:0] node34699;
	wire [4-1:0] node34700;
	wire [4-1:0] node34701;
	wire [4-1:0] node34704;
	wire [4-1:0] node34707;
	wire [4-1:0] node34708;
	wire [4-1:0] node34711;
	wire [4-1:0] node34714;
	wire [4-1:0] node34715;
	wire [4-1:0] node34716;
	wire [4-1:0] node34717;
	wire [4-1:0] node34718;
	wire [4-1:0] node34721;
	wire [4-1:0] node34724;
	wire [4-1:0] node34725;
	wire [4-1:0] node34728;
	wire [4-1:0] node34731;
	wire [4-1:0] node34732;
	wire [4-1:0] node34734;
	wire [4-1:0] node34735;
	wire [4-1:0] node34738;
	wire [4-1:0] node34741;
	wire [4-1:0] node34742;
	wire [4-1:0] node34743;
	wire [4-1:0] node34746;
	wire [4-1:0] node34749;
	wire [4-1:0] node34751;
	wire [4-1:0] node34754;
	wire [4-1:0] node34755;
	wire [4-1:0] node34756;
	wire [4-1:0] node34757;
	wire [4-1:0] node34760;
	wire [4-1:0] node34763;
	wire [4-1:0] node34764;
	wire [4-1:0] node34767;
	wire [4-1:0] node34770;
	wire [4-1:0] node34771;
	wire [4-1:0] node34772;
	wire [4-1:0] node34773;
	wire [4-1:0] node34776;
	wire [4-1:0] node34779;
	wire [4-1:0] node34780;
	wire [4-1:0] node34783;
	wire [4-1:0] node34786;
	wire [4-1:0] node34787;
	wire [4-1:0] node34788;
	wire [4-1:0] node34791;
	wire [4-1:0] node34794;
	wire [4-1:0] node34795;
	wire [4-1:0] node34799;
	wire [4-1:0] node34800;
	wire [4-1:0] node34801;
	wire [4-1:0] node34802;
	wire [4-1:0] node34803;
	wire [4-1:0] node34804;
	wire [4-1:0] node34805;
	wire [4-1:0] node34806;
	wire [4-1:0] node34810;
	wire [4-1:0] node34813;
	wire [4-1:0] node34814;
	wire [4-1:0] node34815;
	wire [4-1:0] node34819;
	wire [4-1:0] node34822;
	wire [4-1:0] node34823;
	wire [4-1:0] node34824;
	wire [4-1:0] node34825;
	wire [4-1:0] node34828;
	wire [4-1:0] node34831;
	wire [4-1:0] node34833;
	wire [4-1:0] node34836;
	wire [4-1:0] node34837;
	wire [4-1:0] node34838;
	wire [4-1:0] node34843;
	wire [4-1:0] node34844;
	wire [4-1:0] node34845;
	wire [4-1:0] node34846;
	wire [4-1:0] node34849;
	wire [4-1:0] node34851;
	wire [4-1:0] node34854;
	wire [4-1:0] node34855;
	wire [4-1:0] node34856;
	wire [4-1:0] node34861;
	wire [4-1:0] node34862;
	wire [4-1:0] node34863;
	wire [4-1:0] node34864;
	wire [4-1:0] node34867;
	wire [4-1:0] node34870;
	wire [4-1:0] node34871;
	wire [4-1:0] node34872;
	wire [4-1:0] node34875;
	wire [4-1:0] node34879;
	wire [4-1:0] node34881;
	wire [4-1:0] node34882;
	wire [4-1:0] node34886;
	wire [4-1:0] node34887;
	wire [4-1:0] node34888;
	wire [4-1:0] node34889;
	wire [4-1:0] node34890;
	wire [4-1:0] node34891;
	wire [4-1:0] node34895;
	wire [4-1:0] node34898;
	wire [4-1:0] node34899;
	wire [4-1:0] node34900;
	wire [4-1:0] node34904;
	wire [4-1:0] node34907;
	wire [4-1:0] node34908;
	wire [4-1:0] node34909;
	wire [4-1:0] node34910;
	wire [4-1:0] node34911;
	wire [4-1:0] node34914;
	wire [4-1:0] node34917;
	wire [4-1:0] node34918;
	wire [4-1:0] node34922;
	wire [4-1:0] node34923;
	wire [4-1:0] node34926;
	wire [4-1:0] node34929;
	wire [4-1:0] node34930;
	wire [4-1:0] node34931;
	wire [4-1:0] node34936;
	wire [4-1:0] node34937;
	wire [4-1:0] node34938;
	wire [4-1:0] node34939;
	wire [4-1:0] node34942;
	wire [4-1:0] node34944;
	wire [4-1:0] node34947;
	wire [4-1:0] node34948;
	wire [4-1:0] node34950;
	wire [4-1:0] node34954;
	wire [4-1:0] node34955;
	wire [4-1:0] node34956;
	wire [4-1:0] node34957;
	wire [4-1:0] node34960;
	wire [4-1:0] node34963;
	wire [4-1:0] node34964;
	wire [4-1:0] node34967;
	wire [4-1:0] node34970;
	wire [4-1:0] node34971;
	wire [4-1:0] node34973;
	wire [4-1:0] node34977;
	wire [4-1:0] node34978;
	wire [4-1:0] node34979;
	wire [4-1:0] node34980;
	wire [4-1:0] node34981;
	wire [4-1:0] node34982;
	wire [4-1:0] node34983;
	wire [4-1:0] node34987;
	wire [4-1:0] node34990;
	wire [4-1:0] node34991;
	wire [4-1:0] node34992;
	wire [4-1:0] node34996;
	wire [4-1:0] node34999;
	wire [4-1:0] node35000;
	wire [4-1:0] node35001;
	wire [4-1:0] node35002;
	wire [4-1:0] node35006;
	wire [4-1:0] node35007;
	wire [4-1:0] node35010;
	wire [4-1:0] node35013;
	wire [4-1:0] node35014;
	wire [4-1:0] node35015;
	wire [4-1:0] node35020;
	wire [4-1:0] node35021;
	wire [4-1:0] node35022;
	wire [4-1:0] node35023;
	wire [4-1:0] node35026;
	wire [4-1:0] node35028;
	wire [4-1:0] node35031;
	wire [4-1:0] node35032;
	wire [4-1:0] node35034;
	wire [4-1:0] node35038;
	wire [4-1:0] node35039;
	wire [4-1:0] node35040;
	wire [4-1:0] node35041;
	wire [4-1:0] node35044;
	wire [4-1:0] node35047;
	wire [4-1:0] node35048;
	wire [4-1:0] node35051;
	wire [4-1:0] node35054;
	wire [4-1:0] node35055;
	wire [4-1:0] node35057;
	wire [4-1:0] node35061;
	wire [4-1:0] node35062;
	wire [4-1:0] node35063;
	wire [4-1:0] node35064;
	wire [4-1:0] node35065;
	wire [4-1:0] node35066;
	wire [4-1:0] node35070;
	wire [4-1:0] node35073;
	wire [4-1:0] node35074;
	wire [4-1:0] node35076;
	wire [4-1:0] node35079;
	wire [4-1:0] node35082;
	wire [4-1:0] node35083;
	wire [4-1:0] node35084;
	wire [4-1:0] node35085;
	wire [4-1:0] node35089;
	wire [4-1:0] node35090;
	wire [4-1:0] node35094;
	wire [4-1:0] node35095;
	wire [4-1:0] node35097;
	wire [4-1:0] node35101;
	wire [4-1:0] node35102;
	wire [4-1:0] node35103;
	wire [4-1:0] node35104;
	wire [4-1:0] node35107;
	wire [4-1:0] node35109;
	wire [4-1:0] node35112;
	wire [4-1:0] node35114;
	wire [4-1:0] node35115;
	wire [4-1:0] node35119;
	wire [4-1:0] node35120;
	wire [4-1:0] node35121;
	wire [4-1:0] node35122;
	wire [4-1:0] node35125;
	wire [4-1:0] node35128;
	wire [4-1:0] node35130;
	wire [4-1:0] node35133;
	wire [4-1:0] node35134;
	wire [4-1:0] node35136;
	wire [4-1:0] node35137;
	wire [4-1:0] node35142;
	wire [4-1:0] node35143;
	wire [4-1:0] node35144;
	wire [4-1:0] node35145;
	wire [4-1:0] node35146;
	wire [4-1:0] node35147;
	wire [4-1:0] node35148;
	wire [4-1:0] node35149;
	wire [4-1:0] node35150;
	wire [4-1:0] node35153;
	wire [4-1:0] node35154;
	wire [4-1:0] node35156;
	wire [4-1:0] node35159;
	wire [4-1:0] node35162;
	wire [4-1:0] node35163;
	wire [4-1:0] node35164;
	wire [4-1:0] node35165;
	wire [4-1:0] node35169;
	wire [4-1:0] node35171;
	wire [4-1:0] node35174;
	wire [4-1:0] node35175;
	wire [4-1:0] node35177;
	wire [4-1:0] node35181;
	wire [4-1:0] node35182;
	wire [4-1:0] node35183;
	wire [4-1:0] node35185;
	wire [4-1:0] node35186;
	wire [4-1:0] node35189;
	wire [4-1:0] node35192;
	wire [4-1:0] node35193;
	wire [4-1:0] node35194;
	wire [4-1:0] node35197;
	wire [4-1:0] node35201;
	wire [4-1:0] node35202;
	wire [4-1:0] node35203;
	wire [4-1:0] node35204;
	wire [4-1:0] node35208;
	wire [4-1:0] node35209;
	wire [4-1:0] node35213;
	wire [4-1:0] node35214;
	wire [4-1:0] node35218;
	wire [4-1:0] node35219;
	wire [4-1:0] node35220;
	wire [4-1:0] node35221;
	wire [4-1:0] node35222;
	wire [4-1:0] node35223;
	wire [4-1:0] node35228;
	wire [4-1:0] node35229;
	wire [4-1:0] node35232;
	wire [4-1:0] node35234;
	wire [4-1:0] node35237;
	wire [4-1:0] node35238;
	wire [4-1:0] node35239;
	wire [4-1:0] node35241;
	wire [4-1:0] node35244;
	wire [4-1:0] node35247;
	wire [4-1:0] node35248;
	wire [4-1:0] node35250;
	wire [4-1:0] node35253;
	wire [4-1:0] node35254;
	wire [4-1:0] node35258;
	wire [4-1:0] node35259;
	wire [4-1:0] node35260;
	wire [4-1:0] node35261;
	wire [4-1:0] node35264;
	wire [4-1:0] node35267;
	wire [4-1:0] node35268;
	wire [4-1:0] node35269;
	wire [4-1:0] node35272;
	wire [4-1:0] node35275;
	wire [4-1:0] node35276;
	wire [4-1:0] node35279;
	wire [4-1:0] node35282;
	wire [4-1:0] node35283;
	wire [4-1:0] node35285;
	wire [4-1:0] node35286;
	wire [4-1:0] node35289;
	wire [4-1:0] node35292;
	wire [4-1:0] node35293;
	wire [4-1:0] node35294;
	wire [4-1:0] node35297;
	wire [4-1:0] node35300;
	wire [4-1:0] node35301;
	wire [4-1:0] node35304;
	wire [4-1:0] node35307;
	wire [4-1:0] node35308;
	wire [4-1:0] node35309;
	wire [4-1:0] node35310;
	wire [4-1:0] node35311;
	wire [4-1:0] node35313;
	wire [4-1:0] node35316;
	wire [4-1:0] node35318;
	wire [4-1:0] node35321;
	wire [4-1:0] node35322;
	wire [4-1:0] node35323;
	wire [4-1:0] node35324;
	wire [4-1:0] node35328;
	wire [4-1:0] node35331;
	wire [4-1:0] node35332;
	wire [4-1:0] node35333;
	wire [4-1:0] node35337;
	wire [4-1:0] node35339;
	wire [4-1:0] node35342;
	wire [4-1:0] node35343;
	wire [4-1:0] node35344;
	wire [4-1:0] node35345;
	wire [4-1:0] node35346;
	wire [4-1:0] node35349;
	wire [4-1:0] node35352;
	wire [4-1:0] node35353;
	wire [4-1:0] node35356;
	wire [4-1:0] node35359;
	wire [4-1:0] node35360;
	wire [4-1:0] node35362;
	wire [4-1:0] node35365;
	wire [4-1:0] node35366;
	wire [4-1:0] node35369;
	wire [4-1:0] node35372;
	wire [4-1:0] node35373;
	wire [4-1:0] node35374;
	wire [4-1:0] node35375;
	wire [4-1:0] node35378;
	wire [4-1:0] node35381;
	wire [4-1:0] node35382;
	wire [4-1:0] node35385;
	wire [4-1:0] node35388;
	wire [4-1:0] node35389;
	wire [4-1:0] node35392;
	wire [4-1:0] node35395;
	wire [4-1:0] node35396;
	wire [4-1:0] node35397;
	wire [4-1:0] node35398;
	wire [4-1:0] node35399;
	wire [4-1:0] node35402;
	wire [4-1:0] node35405;
	wire [4-1:0] node35406;
	wire [4-1:0] node35407;
	wire [4-1:0] node35410;
	wire [4-1:0] node35413;
	wire [4-1:0] node35414;
	wire [4-1:0] node35417;
	wire [4-1:0] node35420;
	wire [4-1:0] node35421;
	wire [4-1:0] node35422;
	wire [4-1:0] node35423;
	wire [4-1:0] node35427;
	wire [4-1:0] node35428;
	wire [4-1:0] node35432;
	wire [4-1:0] node35433;
	wire [4-1:0] node35435;
	wire [4-1:0] node35438;
	wire [4-1:0] node35441;
	wire [4-1:0] node35442;
	wire [4-1:0] node35443;
	wire [4-1:0] node35444;
	wire [4-1:0] node35445;
	wire [4-1:0] node35449;
	wire [4-1:0] node35450;
	wire [4-1:0] node35454;
	wire [4-1:0] node35455;
	wire [4-1:0] node35458;
	wire [4-1:0] node35459;
	wire [4-1:0] node35463;
	wire [4-1:0] node35464;
	wire [4-1:0] node35466;
	wire [4-1:0] node35469;
	wire [4-1:0] node35470;
	wire [4-1:0] node35472;
	wire [4-1:0] node35475;
	wire [4-1:0] node35476;
	wire [4-1:0] node35480;
	wire [4-1:0] node35481;
	wire [4-1:0] node35482;
	wire [4-1:0] node35483;
	wire [4-1:0] node35484;
	wire [4-1:0] node35485;
	wire [4-1:0] node35486;
	wire [4-1:0] node35489;
	wire [4-1:0] node35490;
	wire [4-1:0] node35493;
	wire [4-1:0] node35496;
	wire [4-1:0] node35497;
	wire [4-1:0] node35498;
	wire [4-1:0] node35501;
	wire [4-1:0] node35504;
	wire [4-1:0] node35505;
	wire [4-1:0] node35508;
	wire [4-1:0] node35511;
	wire [4-1:0] node35512;
	wire [4-1:0] node35513;
	wire [4-1:0] node35514;
	wire [4-1:0] node35517;
	wire [4-1:0] node35520;
	wire [4-1:0] node35521;
	wire [4-1:0] node35524;
	wire [4-1:0] node35527;
	wire [4-1:0] node35528;
	wire [4-1:0] node35529;
	wire [4-1:0] node35532;
	wire [4-1:0] node35535;
	wire [4-1:0] node35537;
	wire [4-1:0] node35540;
	wire [4-1:0] node35541;
	wire [4-1:0] node35542;
	wire [4-1:0] node35543;
	wire [4-1:0] node35545;
	wire [4-1:0] node35548;
	wire [4-1:0] node35549;
	wire [4-1:0] node35552;
	wire [4-1:0] node35555;
	wire [4-1:0] node35556;
	wire [4-1:0] node35557;
	wire [4-1:0] node35560;
	wire [4-1:0] node35563;
	wire [4-1:0] node35564;
	wire [4-1:0] node35568;
	wire [4-1:0] node35569;
	wire [4-1:0] node35570;
	wire [4-1:0] node35571;
	wire [4-1:0] node35574;
	wire [4-1:0] node35577;
	wire [4-1:0] node35578;
	wire [4-1:0] node35581;
	wire [4-1:0] node35584;
	wire [4-1:0] node35585;
	wire [4-1:0] node35586;
	wire [4-1:0] node35589;
	wire [4-1:0] node35592;
	wire [4-1:0] node35593;
	wire [4-1:0] node35597;
	wire [4-1:0] node35598;
	wire [4-1:0] node35599;
	wire [4-1:0] node35600;
	wire [4-1:0] node35601;
	wire [4-1:0] node35603;
	wire [4-1:0] node35606;
	wire [4-1:0] node35607;
	wire [4-1:0] node35611;
	wire [4-1:0] node35612;
	wire [4-1:0] node35613;
	wire [4-1:0] node35616;
	wire [4-1:0] node35619;
	wire [4-1:0] node35620;
	wire [4-1:0] node35623;
	wire [4-1:0] node35626;
	wire [4-1:0] node35627;
	wire [4-1:0] node35629;
	wire [4-1:0] node35630;
	wire [4-1:0] node35633;
	wire [4-1:0] node35636;
	wire [4-1:0] node35637;
	wire [4-1:0] node35638;
	wire [4-1:0] node35641;
	wire [4-1:0] node35645;
	wire [4-1:0] node35646;
	wire [4-1:0] node35647;
	wire [4-1:0] node35648;
	wire [4-1:0] node35649;
	wire [4-1:0] node35652;
	wire [4-1:0] node35655;
	wire [4-1:0] node35656;
	wire [4-1:0] node35660;
	wire [4-1:0] node35661;
	wire [4-1:0] node35664;
	wire [4-1:0] node35665;
	wire [4-1:0] node35668;
	wire [4-1:0] node35671;
	wire [4-1:0] node35672;
	wire [4-1:0] node35673;
	wire [4-1:0] node35674;
	wire [4-1:0] node35677;
	wire [4-1:0] node35680;
	wire [4-1:0] node35681;
	wire [4-1:0] node35684;
	wire [4-1:0] node35687;
	wire [4-1:0] node35688;
	wire [4-1:0] node35689;
	wire [4-1:0] node35692;
	wire [4-1:0] node35695;
	wire [4-1:0] node35696;
	wire [4-1:0] node35699;
	wire [4-1:0] node35702;
	wire [4-1:0] node35703;
	wire [4-1:0] node35704;
	wire [4-1:0] node35705;
	wire [4-1:0] node35706;
	wire [4-1:0] node35707;
	wire [4-1:0] node35708;
	wire [4-1:0] node35711;
	wire [4-1:0] node35714;
	wire [4-1:0] node35715;
	wire [4-1:0] node35718;
	wire [4-1:0] node35721;
	wire [4-1:0] node35722;
	wire [4-1:0] node35723;
	wire [4-1:0] node35727;
	wire [4-1:0] node35728;
	wire [4-1:0] node35731;
	wire [4-1:0] node35734;
	wire [4-1:0] node35735;
	wire [4-1:0] node35736;
	wire [4-1:0] node35737;
	wire [4-1:0] node35740;
	wire [4-1:0] node35743;
	wire [4-1:0] node35744;
	wire [4-1:0] node35747;
	wire [4-1:0] node35750;
	wire [4-1:0] node35751;
	wire [4-1:0] node35752;
	wire [4-1:0] node35755;
	wire [4-1:0] node35758;
	wire [4-1:0] node35759;
	wire [4-1:0] node35762;
	wire [4-1:0] node35765;
	wire [4-1:0] node35766;
	wire [4-1:0] node35767;
	wire [4-1:0] node35768;
	wire [4-1:0] node35769;
	wire [4-1:0] node35772;
	wire [4-1:0] node35775;
	wire [4-1:0] node35776;
	wire [4-1:0] node35779;
	wire [4-1:0] node35782;
	wire [4-1:0] node35783;
	wire [4-1:0] node35784;
	wire [4-1:0] node35787;
	wire [4-1:0] node35790;
	wire [4-1:0] node35791;
	wire [4-1:0] node35794;
	wire [4-1:0] node35797;
	wire [4-1:0] node35798;
	wire [4-1:0] node35799;
	wire [4-1:0] node35802;
	wire [4-1:0] node35803;
	wire [4-1:0] node35806;
	wire [4-1:0] node35809;
	wire [4-1:0] node35810;
	wire [4-1:0] node35811;
	wire [4-1:0] node35814;
	wire [4-1:0] node35817;
	wire [4-1:0] node35819;
	wire [4-1:0] node35822;
	wire [4-1:0] node35823;
	wire [4-1:0] node35824;
	wire [4-1:0] node35825;
	wire [4-1:0] node35826;
	wire [4-1:0] node35827;
	wire [4-1:0] node35830;
	wire [4-1:0] node35833;
	wire [4-1:0] node35834;
	wire [4-1:0] node35837;
	wire [4-1:0] node35840;
	wire [4-1:0] node35841;
	wire [4-1:0] node35843;
	wire [4-1:0] node35846;
	wire [4-1:0] node35849;
	wire [4-1:0] node35850;
	wire [4-1:0] node35851;
	wire [4-1:0] node35852;
	wire [4-1:0] node35855;
	wire [4-1:0] node35858;
	wire [4-1:0] node35861;
	wire [4-1:0] node35862;
	wire [4-1:0] node35863;
	wire [4-1:0] node35866;
	wire [4-1:0] node35869;
	wire [4-1:0] node35872;
	wire [4-1:0] node35873;
	wire [4-1:0] node35874;
	wire [4-1:0] node35875;
	wire [4-1:0] node35877;
	wire [4-1:0] node35880;
	wire [4-1:0] node35881;
	wire [4-1:0] node35885;
	wire [4-1:0] node35886;
	wire [4-1:0] node35887;
	wire [4-1:0] node35890;
	wire [4-1:0] node35893;
	wire [4-1:0] node35894;
	wire [4-1:0] node35897;
	wire [4-1:0] node35900;
	wire [4-1:0] node35901;
	wire [4-1:0] node35902;
	wire [4-1:0] node35903;
	wire [4-1:0] node35906;
	wire [4-1:0] node35909;
	wire [4-1:0] node35911;
	wire [4-1:0] node35914;
	wire [4-1:0] node35915;
	wire [4-1:0] node35917;
	wire [4-1:0] node35920;
	wire [4-1:0] node35923;
	wire [4-1:0] node35924;
	wire [4-1:0] node35925;
	wire [4-1:0] node35926;
	wire [4-1:0] node35927;
	wire [4-1:0] node35928;
	wire [4-1:0] node35929;
	wire [4-1:0] node35930;
	wire [4-1:0] node35931;
	wire [4-1:0] node35934;
	wire [4-1:0] node35937;
	wire [4-1:0] node35938;
	wire [4-1:0] node35941;
	wire [4-1:0] node35944;
	wire [4-1:0] node35945;
	wire [4-1:0] node35948;
	wire [4-1:0] node35951;
	wire [4-1:0] node35952;
	wire [4-1:0] node35953;
	wire [4-1:0] node35955;
	wire [4-1:0] node35959;
	wire [4-1:0] node35960;
	wire [4-1:0] node35963;
	wire [4-1:0] node35966;
	wire [4-1:0] node35967;
	wire [4-1:0] node35968;
	wire [4-1:0] node35969;
	wire [4-1:0] node35972;
	wire [4-1:0] node35975;
	wire [4-1:0] node35976;
	wire [4-1:0] node35977;
	wire [4-1:0] node35980;
	wire [4-1:0] node35984;
	wire [4-1:0] node35985;
	wire [4-1:0] node35986;
	wire [4-1:0] node35987;
	wire [4-1:0] node35990;
	wire [4-1:0] node35993;
	wire [4-1:0] node35994;
	wire [4-1:0] node35997;
	wire [4-1:0] node36000;
	wire [4-1:0] node36001;
	wire [4-1:0] node36002;
	wire [4-1:0] node36005;
	wire [4-1:0] node36008;
	wire [4-1:0] node36009;
	wire [4-1:0] node36012;
	wire [4-1:0] node36015;
	wire [4-1:0] node36016;
	wire [4-1:0] node36017;
	wire [4-1:0] node36018;
	wire [4-1:0] node36019;
	wire [4-1:0] node36020;
	wire [4-1:0] node36024;
	wire [4-1:0] node36027;
	wire [4-1:0] node36028;
	wire [4-1:0] node36032;
	wire [4-1:0] node36033;
	wire [4-1:0] node36034;
	wire [4-1:0] node36035;
	wire [4-1:0] node36038;
	wire [4-1:0] node36041;
	wire [4-1:0] node36043;
	wire [4-1:0] node36046;
	wire [4-1:0] node36047;
	wire [4-1:0] node36048;
	wire [4-1:0] node36052;
	wire [4-1:0] node36055;
	wire [4-1:0] node36056;
	wire [4-1:0] node36057;
	wire [4-1:0] node36058;
	wire [4-1:0] node36061;
	wire [4-1:0] node36062;
	wire [4-1:0] node36066;
	wire [4-1:0] node36067;
	wire [4-1:0] node36069;
	wire [4-1:0] node36073;
	wire [4-1:0] node36074;
	wire [4-1:0] node36077;
	wire [4-1:0] node36078;
	wire [4-1:0] node36079;
	wire [4-1:0] node36083;
	wire [4-1:0] node36084;
	wire [4-1:0] node36088;
	wire [4-1:0] node36089;
	wire [4-1:0] node36090;
	wire [4-1:0] node36091;
	wire [4-1:0] node36092;
	wire [4-1:0] node36093;
	wire [4-1:0] node36094;
	wire [4-1:0] node36097;
	wire [4-1:0] node36100;
	wire [4-1:0] node36101;
	wire [4-1:0] node36104;
	wire [4-1:0] node36107;
	wire [4-1:0] node36108;
	wire [4-1:0] node36111;
	wire [4-1:0] node36112;
	wire [4-1:0] node36115;
	wire [4-1:0] node36118;
	wire [4-1:0] node36119;
	wire [4-1:0] node36120;
	wire [4-1:0] node36123;
	wire [4-1:0] node36124;
	wire [4-1:0] node36127;
	wire [4-1:0] node36130;
	wire [4-1:0] node36131;
	wire [4-1:0] node36134;
	wire [4-1:0] node36135;
	wire [4-1:0] node36138;
	wire [4-1:0] node36141;
	wire [4-1:0] node36142;
	wire [4-1:0] node36143;
	wire [4-1:0] node36144;
	wire [4-1:0] node36145;
	wire [4-1:0] node36148;
	wire [4-1:0] node36151;
	wire [4-1:0] node36152;
	wire [4-1:0] node36155;
	wire [4-1:0] node36158;
	wire [4-1:0] node36159;
	wire [4-1:0] node36160;
	wire [4-1:0] node36164;
	wire [4-1:0] node36165;
	wire [4-1:0] node36168;
	wire [4-1:0] node36171;
	wire [4-1:0] node36172;
	wire [4-1:0] node36173;
	wire [4-1:0] node36174;
	wire [4-1:0] node36178;
	wire [4-1:0] node36181;
	wire [4-1:0] node36182;
	wire [4-1:0] node36183;
	wire [4-1:0] node36187;
	wire [4-1:0] node36190;
	wire [4-1:0] node36191;
	wire [4-1:0] node36192;
	wire [4-1:0] node36193;
	wire [4-1:0] node36194;
	wire [4-1:0] node36195;
	wire [4-1:0] node36198;
	wire [4-1:0] node36201;
	wire [4-1:0] node36202;
	wire [4-1:0] node36205;
	wire [4-1:0] node36208;
	wire [4-1:0] node36209;
	wire [4-1:0] node36210;
	wire [4-1:0] node36213;
	wire [4-1:0] node36217;
	wire [4-1:0] node36218;
	wire [4-1:0] node36219;
	wire [4-1:0] node36220;
	wire [4-1:0] node36224;
	wire [4-1:0] node36227;
	wire [4-1:0] node36228;
	wire [4-1:0] node36231;
	wire [4-1:0] node36234;
	wire [4-1:0] node36235;
	wire [4-1:0] node36236;
	wire [4-1:0] node36237;
	wire [4-1:0] node36240;
	wire [4-1:0] node36243;
	wire [4-1:0] node36244;
	wire [4-1:0] node36245;
	wire [4-1:0] node36248;
	wire [4-1:0] node36251;
	wire [4-1:0] node36253;
	wire [4-1:0] node36256;
	wire [4-1:0] node36257;
	wire [4-1:0] node36258;
	wire [4-1:0] node36260;
	wire [4-1:0] node36263;
	wire [4-1:0] node36266;
	wire [4-1:0] node36267;
	wire [4-1:0] node36268;
	wire [4-1:0] node36273;
	wire [4-1:0] node36274;
	wire [4-1:0] node36275;
	wire [4-1:0] node36276;
	wire [4-1:0] node36277;
	wire [4-1:0] node36278;
	wire [4-1:0] node36279;
	wire [4-1:0] node36281;
	wire [4-1:0] node36284;
	wire [4-1:0] node36285;
	wire [4-1:0] node36288;
	wire [4-1:0] node36291;
	wire [4-1:0] node36292;
	wire [4-1:0] node36293;
	wire [4-1:0] node36297;
	wire [4-1:0] node36298;
	wire [4-1:0] node36302;
	wire [4-1:0] node36303;
	wire [4-1:0] node36304;
	wire [4-1:0] node36307;
	wire [4-1:0] node36308;
	wire [4-1:0] node36312;
	wire [4-1:0] node36313;
	wire [4-1:0] node36316;
	wire [4-1:0] node36318;
	wire [4-1:0] node36321;
	wire [4-1:0] node36322;
	wire [4-1:0] node36323;
	wire [4-1:0] node36324;
	wire [4-1:0] node36327;
	wire [4-1:0] node36330;
	wire [4-1:0] node36331;
	wire [4-1:0] node36332;
	wire [4-1:0] node36336;
	wire [4-1:0] node36338;
	wire [4-1:0] node36341;
	wire [4-1:0] node36342;
	wire [4-1:0] node36343;
	wire [4-1:0] node36346;
	wire [4-1:0] node36348;
	wire [4-1:0] node36351;
	wire [4-1:0] node36352;
	wire [4-1:0] node36353;
	wire [4-1:0] node36357;
	wire [4-1:0] node36359;
	wire [4-1:0] node36362;
	wire [4-1:0] node36363;
	wire [4-1:0] node36364;
	wire [4-1:0] node36365;
	wire [4-1:0] node36366;
	wire [4-1:0] node36369;
	wire [4-1:0] node36372;
	wire [4-1:0] node36373;
	wire [4-1:0] node36374;
	wire [4-1:0] node36377;
	wire [4-1:0] node36380;
	wire [4-1:0] node36383;
	wire [4-1:0] node36384;
	wire [4-1:0] node36385;
	wire [4-1:0] node36387;
	wire [4-1:0] node36390;
	wire [4-1:0] node36391;
	wire [4-1:0] node36395;
	wire [4-1:0] node36396;
	wire [4-1:0] node36399;
	wire [4-1:0] node36400;
	wire [4-1:0] node36404;
	wire [4-1:0] node36405;
	wire [4-1:0] node36406;
	wire [4-1:0] node36407;
	wire [4-1:0] node36408;
	wire [4-1:0] node36411;
	wire [4-1:0] node36414;
	wire [4-1:0] node36416;
	wire [4-1:0] node36419;
	wire [4-1:0] node36420;
	wire [4-1:0] node36423;
	wire [4-1:0] node36425;
	wire [4-1:0] node36428;
	wire [4-1:0] node36429;
	wire [4-1:0] node36430;
	wire [4-1:0] node36433;
	wire [4-1:0] node36436;
	wire [4-1:0] node36437;
	wire [4-1:0] node36439;
	wire [4-1:0] node36442;
	wire [4-1:0] node36444;
	wire [4-1:0] node36447;
	wire [4-1:0] node36448;
	wire [4-1:0] node36449;
	wire [4-1:0] node36450;
	wire [4-1:0] node36451;
	wire [4-1:0] node36452;
	wire [4-1:0] node36455;
	wire [4-1:0] node36458;
	wire [4-1:0] node36460;
	wire [4-1:0] node36461;
	wire [4-1:0] node36464;
	wire [4-1:0] node36467;
	wire [4-1:0] node36468;
	wire [4-1:0] node36469;
	wire [4-1:0] node36471;
	wire [4-1:0] node36475;
	wire [4-1:0] node36476;
	wire [4-1:0] node36477;
	wire [4-1:0] node36481;
	wire [4-1:0] node36482;
	wire [4-1:0] node36485;
	wire [4-1:0] node36488;
	wire [4-1:0] node36489;
	wire [4-1:0] node36490;
	wire [4-1:0] node36491;
	wire [4-1:0] node36494;
	wire [4-1:0] node36497;
	wire [4-1:0] node36499;
	wire [4-1:0] node36500;
	wire [4-1:0] node36503;
	wire [4-1:0] node36506;
	wire [4-1:0] node36507;
	wire [4-1:0] node36508;
	wire [4-1:0] node36509;
	wire [4-1:0] node36512;
	wire [4-1:0] node36515;
	wire [4-1:0] node36517;
	wire [4-1:0] node36520;
	wire [4-1:0] node36521;
	wire [4-1:0] node36522;
	wire [4-1:0] node36525;
	wire [4-1:0] node36528;
	wire [4-1:0] node36529;
	wire [4-1:0] node36532;
	wire [4-1:0] node36535;
	wire [4-1:0] node36536;
	wire [4-1:0] node36537;
	wire [4-1:0] node36538;
	wire [4-1:0] node36539;
	wire [4-1:0] node36540;
	wire [4-1:0] node36543;
	wire [4-1:0] node36546;
	wire [4-1:0] node36547;
	wire [4-1:0] node36551;
	wire [4-1:0] node36552;
	wire [4-1:0] node36553;
	wire [4-1:0] node36557;
	wire [4-1:0] node36560;
	wire [4-1:0] node36561;
	wire [4-1:0] node36562;
	wire [4-1:0] node36565;
	wire [4-1:0] node36568;
	wire [4-1:0] node36569;
	wire [4-1:0] node36571;
	wire [4-1:0] node36574;
	wire [4-1:0] node36577;
	wire [4-1:0] node36578;
	wire [4-1:0] node36579;
	wire [4-1:0] node36580;
	wire [4-1:0] node36581;
	wire [4-1:0] node36585;
	wire [4-1:0] node36586;
	wire [4-1:0] node36590;
	wire [4-1:0] node36591;
	wire [4-1:0] node36592;
	wire [4-1:0] node36595;
	wire [4-1:0] node36598;
	wire [4-1:0] node36599;
	wire [4-1:0] node36602;
	wire [4-1:0] node36605;
	wire [4-1:0] node36606;
	wire [4-1:0] node36607;
	wire [4-1:0] node36608;
	wire [4-1:0] node36611;
	wire [4-1:0] node36614;
	wire [4-1:0] node36615;
	wire [4-1:0] node36618;
	wire [4-1:0] node36621;
	wire [4-1:0] node36622;
	wire [4-1:0] node36623;
	wire [4-1:0] node36626;
	wire [4-1:0] node36629;
	wire [4-1:0] node36630;
	wire [4-1:0] node36633;
	wire [4-1:0] node36636;
	wire [4-1:0] node36637;
	wire [4-1:0] node36638;
	wire [4-1:0] node36639;
	wire [4-1:0] node36640;
	wire [4-1:0] node36641;
	wire [4-1:0] node36642;
	wire [4-1:0] node36643;
	wire [4-1:0] node36644;
	wire [4-1:0] node36645;
	wire [4-1:0] node36648;
	wire [4-1:0] node36651;
	wire [4-1:0] node36652;
	wire [4-1:0] node36655;
	wire [4-1:0] node36658;
	wire [4-1:0] node36659;
	wire [4-1:0] node36660;
	wire [4-1:0] node36664;
	wire [4-1:0] node36665;
	wire [4-1:0] node36668;
	wire [4-1:0] node36671;
	wire [4-1:0] node36672;
	wire [4-1:0] node36673;
	wire [4-1:0] node36676;
	wire [4-1:0] node36679;
	wire [4-1:0] node36680;
	wire [4-1:0] node36681;
	wire [4-1:0] node36685;
	wire [4-1:0] node36686;
	wire [4-1:0] node36689;
	wire [4-1:0] node36692;
	wire [4-1:0] node36693;
	wire [4-1:0] node36694;
	wire [4-1:0] node36695;
	wire [4-1:0] node36699;
	wire [4-1:0] node36701;
	wire [4-1:0] node36704;
	wire [4-1:0] node36705;
	wire [4-1:0] node36706;
	wire [4-1:0] node36710;
	wire [4-1:0] node36711;
	wire [4-1:0] node36715;
	wire [4-1:0] node36716;
	wire [4-1:0] node36717;
	wire [4-1:0] node36718;
	wire [4-1:0] node36721;
	wire [4-1:0] node36724;
	wire [4-1:0] node36725;
	wire [4-1:0] node36726;
	wire [4-1:0] node36727;
	wire [4-1:0] node36730;
	wire [4-1:0] node36733;
	wire [4-1:0] node36734;
	wire [4-1:0] node36737;
	wire [4-1:0] node36740;
	wire [4-1:0] node36741;
	wire [4-1:0] node36744;
	wire [4-1:0] node36747;
	wire [4-1:0] node36748;
	wire [4-1:0] node36749;
	wire [4-1:0] node36750;
	wire [4-1:0] node36753;
	wire [4-1:0] node36756;
	wire [4-1:0] node36757;
	wire [4-1:0] node36760;
	wire [4-1:0] node36763;
	wire [4-1:0] node36764;
	wire [4-1:0] node36765;
	wire [4-1:0] node36768;
	wire [4-1:0] node36771;
	wire [4-1:0] node36772;
	wire [4-1:0] node36775;
	wire [4-1:0] node36778;
	wire [4-1:0] node36779;
	wire [4-1:0] node36780;
	wire [4-1:0] node36781;
	wire [4-1:0] node36782;
	wire [4-1:0] node36783;
	wire [4-1:0] node36784;
	wire [4-1:0] node36788;
	wire [4-1:0] node36791;
	wire [4-1:0] node36792;
	wire [4-1:0] node36794;
	wire [4-1:0] node36797;
	wire [4-1:0] node36800;
	wire [4-1:0] node36801;
	wire [4-1:0] node36802;
	wire [4-1:0] node36803;
	wire [4-1:0] node36807;
	wire [4-1:0] node36809;
	wire [4-1:0] node36812;
	wire [4-1:0] node36814;
	wire [4-1:0] node36815;
	wire [4-1:0] node36818;
	wire [4-1:0] node36821;
	wire [4-1:0] node36822;
	wire [4-1:0] node36823;
	wire [4-1:0] node36824;
	wire [4-1:0] node36828;
	wire [4-1:0] node36829;
	wire [4-1:0] node36833;
	wire [4-1:0] node36834;
	wire [4-1:0] node36836;
	wire [4-1:0] node36839;
	wire [4-1:0] node36842;
	wire [4-1:0] node36843;
	wire [4-1:0] node36844;
	wire [4-1:0] node36845;
	wire [4-1:0] node36846;
	wire [4-1:0] node36849;
	wire [4-1:0] node36852;
	wire [4-1:0] node36853;
	wire [4-1:0] node36856;
	wire [4-1:0] node36859;
	wire [4-1:0] node36860;
	wire [4-1:0] node36863;
	wire [4-1:0] node36866;
	wire [4-1:0] node36867;
	wire [4-1:0] node36868;
	wire [4-1:0] node36871;
	wire [4-1:0] node36874;
	wire [4-1:0] node36875;
	wire [4-1:0] node36876;
	wire [4-1:0] node36879;
	wire [4-1:0] node36882;
	wire [4-1:0] node36883;
	wire [4-1:0] node36886;
	wire [4-1:0] node36889;
	wire [4-1:0] node36890;
	wire [4-1:0] node36891;
	wire [4-1:0] node36892;
	wire [4-1:0] node36893;
	wire [4-1:0] node36894;
	wire [4-1:0] node36896;
	wire [4-1:0] node36899;
	wire [4-1:0] node36901;
	wire [4-1:0] node36902;
	wire [4-1:0] node36906;
	wire [4-1:0] node36907;
	wire [4-1:0] node36908;
	wire [4-1:0] node36909;
	wire [4-1:0] node36912;
	wire [4-1:0] node36915;
	wire [4-1:0] node36916;
	wire [4-1:0] node36919;
	wire [4-1:0] node36922;
	wire [4-1:0] node36923;
	wire [4-1:0] node36926;
	wire [4-1:0] node36929;
	wire [4-1:0] node36930;
	wire [4-1:0] node36931;
	wire [4-1:0] node36934;
	wire [4-1:0] node36937;
	wire [4-1:0] node36938;
	wire [4-1:0] node36940;
	wire [4-1:0] node36941;
	wire [4-1:0] node36944;
	wire [4-1:0] node36947;
	wire [4-1:0] node36948;
	wire [4-1:0] node36949;
	wire [4-1:0] node36952;
	wire [4-1:0] node36955;
	wire [4-1:0] node36956;
	wire [4-1:0] node36959;
	wire [4-1:0] node36962;
	wire [4-1:0] node36963;
	wire [4-1:0] node36964;
	wire [4-1:0] node36965;
	wire [4-1:0] node36966;
	wire [4-1:0] node36970;
	wire [4-1:0] node36973;
	wire [4-1:0] node36974;
	wire [4-1:0] node36976;
	wire [4-1:0] node36979;
	wire [4-1:0] node36980;
	wire [4-1:0] node36983;
	wire [4-1:0] node36986;
	wire [4-1:0] node36987;
	wire [4-1:0] node36988;
	wire [4-1:0] node36989;
	wire [4-1:0] node36994;
	wire [4-1:0] node36995;
	wire [4-1:0] node36999;
	wire [4-1:0] node37000;
	wire [4-1:0] node37001;
	wire [4-1:0] node37002;
	wire [4-1:0] node37003;
	wire [4-1:0] node37004;
	wire [4-1:0] node37007;
	wire [4-1:0] node37010;
	wire [4-1:0] node37011;
	wire [4-1:0] node37012;
	wire [4-1:0] node37017;
	wire [4-1:0] node37018;
	wire [4-1:0] node37019;
	wire [4-1:0] node37022;
	wire [4-1:0] node37025;
	wire [4-1:0] node37026;
	wire [4-1:0] node37029;
	wire [4-1:0] node37032;
	wire [4-1:0] node37033;
	wire [4-1:0] node37035;
	wire [4-1:0] node37036;
	wire [4-1:0] node37039;
	wire [4-1:0] node37041;
	wire [4-1:0] node37044;
	wire [4-1:0] node37045;
	wire [4-1:0] node37046;
	wire [4-1:0] node37047;
	wire [4-1:0] node37050;
	wire [4-1:0] node37053;
	wire [4-1:0] node37054;
	wire [4-1:0] node37057;
	wire [4-1:0] node37060;
	wire [4-1:0] node37061;
	wire [4-1:0] node37064;
	wire [4-1:0] node37067;
	wire [4-1:0] node37068;
	wire [4-1:0] node37069;
	wire [4-1:0] node37070;
	wire [4-1:0] node37072;
	wire [4-1:0] node37075;
	wire [4-1:0] node37076;
	wire [4-1:0] node37079;
	wire [4-1:0] node37082;
	wire [4-1:0] node37083;
	wire [4-1:0] node37084;
	wire [4-1:0] node37088;
	wire [4-1:0] node37091;
	wire [4-1:0] node37092;
	wire [4-1:0] node37093;
	wire [4-1:0] node37094;
	wire [4-1:0] node37099;
	wire [4-1:0] node37100;
	wire [4-1:0] node37101;
	wire [4-1:0] node37106;
	wire [4-1:0] node37107;
	wire [4-1:0] node37108;
	wire [4-1:0] node37109;
	wire [4-1:0] node37110;
	wire [4-1:0] node37111;
	wire [4-1:0] node37112;
	wire [4-1:0] node37113;
	wire [4-1:0] node37115;
	wire [4-1:0] node37118;
	wire [4-1:0] node37119;
	wire [4-1:0] node37122;
	wire [4-1:0] node37125;
	wire [4-1:0] node37126;
	wire [4-1:0] node37127;
	wire [4-1:0] node37131;
	wire [4-1:0] node37132;
	wire [4-1:0] node37135;
	wire [4-1:0] node37138;
	wire [4-1:0] node37139;
	wire [4-1:0] node37140;
	wire [4-1:0] node37142;
	wire [4-1:0] node37145;
	wire [4-1:0] node37146;
	wire [4-1:0] node37150;
	wire [4-1:0] node37151;
	wire [4-1:0] node37152;
	wire [4-1:0] node37156;
	wire [4-1:0] node37157;
	wire [4-1:0] node37161;
	wire [4-1:0] node37162;
	wire [4-1:0] node37163;
	wire [4-1:0] node37164;
	wire [4-1:0] node37166;
	wire [4-1:0] node37169;
	wire [4-1:0] node37170;
	wire [4-1:0] node37174;
	wire [4-1:0] node37176;
	wire [4-1:0] node37179;
	wire [4-1:0] node37180;
	wire [4-1:0] node37181;
	wire [4-1:0] node37182;
	wire [4-1:0] node37185;
	wire [4-1:0] node37188;
	wire [4-1:0] node37189;
	wire [4-1:0] node37192;
	wire [4-1:0] node37195;
	wire [4-1:0] node37196;
	wire [4-1:0] node37197;
	wire [4-1:0] node37200;
	wire [4-1:0] node37203;
	wire [4-1:0] node37204;
	wire [4-1:0] node37207;
	wire [4-1:0] node37210;
	wire [4-1:0] node37211;
	wire [4-1:0] node37212;
	wire [4-1:0] node37215;
	wire [4-1:0] node37218;
	wire [4-1:0] node37219;
	wire [4-1:0] node37220;
	wire [4-1:0] node37221;
	wire [4-1:0] node37224;
	wire [4-1:0] node37227;
	wire [4-1:0] node37228;
	wire [4-1:0] node37229;
	wire [4-1:0] node37232;
	wire [4-1:0] node37235;
	wire [4-1:0] node37236;
	wire [4-1:0] node37239;
	wire [4-1:0] node37242;
	wire [4-1:0] node37243;
	wire [4-1:0] node37244;
	wire [4-1:0] node37247;
	wire [4-1:0] node37251;
	wire [4-1:0] node37252;
	wire [4-1:0] node37253;
	wire [4-1:0] node37254;
	wire [4-1:0] node37255;
	wire [4-1:0] node37256;
	wire [4-1:0] node37260;
	wire [4-1:0] node37261;
	wire [4-1:0] node37265;
	wire [4-1:0] node37266;
	wire [4-1:0] node37267;
	wire [4-1:0] node37271;
	wire [4-1:0] node37273;
	wire [4-1:0] node37276;
	wire [4-1:0] node37277;
	wire [4-1:0] node37278;
	wire [4-1:0] node37279;
	wire [4-1:0] node37280;
	wire [4-1:0] node37285;
	wire [4-1:0] node37286;
	wire [4-1:0] node37289;
	wire [4-1:0] node37291;
	wire [4-1:0] node37294;
	wire [4-1:0] node37295;
	wire [4-1:0] node37296;
	wire [4-1:0] node37299;
	wire [4-1:0] node37302;
	wire [4-1:0] node37303;
	wire [4-1:0] node37306;
	wire [4-1:0] node37309;
	wire [4-1:0] node37310;
	wire [4-1:0] node37311;
	wire [4-1:0] node37312;
	wire [4-1:0] node37316;
	wire [4-1:0] node37317;
	wire [4-1:0] node37321;
	wire [4-1:0] node37322;
	wire [4-1:0] node37323;
	wire [4-1:0] node37327;
	wire [4-1:0] node37328;
	wire [4-1:0] node37332;
	wire [4-1:0] node37333;
	wire [4-1:0] node37334;
	wire [4-1:0] node37335;
	wire [4-1:0] node37336;
	wire [4-1:0] node37337;
	wire [4-1:0] node37338;
	wire [4-1:0] node37339;
	wire [4-1:0] node37342;
	wire [4-1:0] node37345;
	wire [4-1:0] node37346;
	wire [4-1:0] node37349;
	wire [4-1:0] node37352;
	wire [4-1:0] node37353;
	wire [4-1:0] node37354;
	wire [4-1:0] node37357;
	wire [4-1:0] node37361;
	wire [4-1:0] node37362;
	wire [4-1:0] node37363;
	wire [4-1:0] node37364;
	wire [4-1:0] node37367;
	wire [4-1:0] node37371;
	wire [4-1:0] node37372;
	wire [4-1:0] node37373;
	wire [4-1:0] node37377;
	wire [4-1:0] node37378;
	wire [4-1:0] node37381;
	wire [4-1:0] node37384;
	wire [4-1:0] node37385;
	wire [4-1:0] node37386;
	wire [4-1:0] node37387;
	wire [4-1:0] node37388;
	wire [4-1:0] node37391;
	wire [4-1:0] node37394;
	wire [4-1:0] node37395;
	wire [4-1:0] node37398;
	wire [4-1:0] node37401;
	wire [4-1:0] node37402;
	wire [4-1:0] node37403;
	wire [4-1:0] node37407;
	wire [4-1:0] node37408;
	wire [4-1:0] node37411;
	wire [4-1:0] node37414;
	wire [4-1:0] node37415;
	wire [4-1:0] node37416;
	wire [4-1:0] node37419;
	wire [4-1:0] node37422;
	wire [4-1:0] node37423;
	wire [4-1:0] node37426;
	wire [4-1:0] node37428;
	wire [4-1:0] node37431;
	wire [4-1:0] node37432;
	wire [4-1:0] node37433;
	wire [4-1:0] node37434;
	wire [4-1:0] node37435;
	wire [4-1:0] node37439;
	wire [4-1:0] node37440;
	wire [4-1:0] node37444;
	wire [4-1:0] node37445;
	wire [4-1:0] node37446;
	wire [4-1:0] node37450;
	wire [4-1:0] node37451;
	wire [4-1:0] node37455;
	wire [4-1:0] node37456;
	wire [4-1:0] node37457;
	wire [4-1:0] node37458;
	wire [4-1:0] node37461;
	wire [4-1:0] node37464;
	wire [4-1:0] node37465;
	wire [4-1:0] node37466;
	wire [4-1:0] node37469;
	wire [4-1:0] node37472;
	wire [4-1:0] node37474;
	wire [4-1:0] node37477;
	wire [4-1:0] node37478;
	wire [4-1:0] node37479;
	wire [4-1:0] node37480;
	wire [4-1:0] node37483;
	wire [4-1:0] node37486;
	wire [4-1:0] node37487;
	wire [4-1:0] node37490;
	wire [4-1:0] node37493;
	wire [4-1:0] node37494;
	wire [4-1:0] node37498;
	wire [4-1:0] node37499;
	wire [4-1:0] node37500;
	wire [4-1:0] node37501;
	wire [4-1:0] node37502;
	wire [4-1:0] node37503;
	wire [4-1:0] node37507;
	wire [4-1:0] node37510;
	wire [4-1:0] node37511;
	wire [4-1:0] node37512;
	wire [4-1:0] node37516;
	wire [4-1:0] node37518;
	wire [4-1:0] node37521;
	wire [4-1:0] node37522;
	wire [4-1:0] node37523;
	wire [4-1:0] node37524;
	wire [4-1:0] node37527;
	wire [4-1:0] node37530;
	wire [4-1:0] node37531;
	wire [4-1:0] node37532;
	wire [4-1:0] node37536;
	wire [4-1:0] node37537;
	wire [4-1:0] node37540;
	wire [4-1:0] node37543;
	wire [4-1:0] node37544;
	wire [4-1:0] node37545;
	wire [4-1:0] node37547;
	wire [4-1:0] node37550;
	wire [4-1:0] node37551;
	wire [4-1:0] node37554;
	wire [4-1:0] node37557;
	wire [4-1:0] node37558;
	wire [4-1:0] node37561;
	wire [4-1:0] node37564;
	wire [4-1:0] node37565;
	wire [4-1:0] node37566;
	wire [4-1:0] node37567;
	wire [4-1:0] node37568;
	wire [4-1:0] node37571;
	wire [4-1:0] node37574;
	wire [4-1:0] node37575;
	wire [4-1:0] node37576;
	wire [4-1:0] node37579;
	wire [4-1:0] node37582;
	wire [4-1:0] node37583;
	wire [4-1:0] node37586;
	wire [4-1:0] node37589;
	wire [4-1:0] node37590;
	wire [4-1:0] node37593;
	wire [4-1:0] node37596;
	wire [4-1:0] node37597;
	wire [4-1:0] node37600;
	wire [4-1:0] node37603;
	wire [4-1:0] node37604;
	wire [4-1:0] node37605;
	wire [4-1:0] node37606;
	wire [4-1:0] node37607;
	wire [4-1:0] node37608;
	wire [4-1:0] node37609;
	wire [4-1:0] node37610;
	wire [4-1:0] node37611;
	wire [4-1:0] node37612;
	wire [4-1:0] node37613;
	wire [4-1:0] node37614;
	wire [4-1:0] node37615;
	wire [4-1:0] node37619;
	wire [4-1:0] node37621;
	wire [4-1:0] node37624;
	wire [4-1:0] node37625;
	wire [4-1:0] node37628;
	wire [4-1:0] node37629;
	wire [4-1:0] node37632;
	wire [4-1:0] node37635;
	wire [4-1:0] node37636;
	wire [4-1:0] node37637;
	wire [4-1:0] node37639;
	wire [4-1:0] node37642;
	wire [4-1:0] node37645;
	wire [4-1:0] node37646;
	wire [4-1:0] node37648;
	wire [4-1:0] node37651;
	wire [4-1:0] node37654;
	wire [4-1:0] node37655;
	wire [4-1:0] node37656;
	wire [4-1:0] node37657;
	wire [4-1:0] node37658;
	wire [4-1:0] node37662;
	wire [4-1:0] node37665;
	wire [4-1:0] node37666;
	wire [4-1:0] node37667;
	wire [4-1:0] node37670;
	wire [4-1:0] node37673;
	wire [4-1:0] node37674;
	wire [4-1:0] node37678;
	wire [4-1:0] node37679;
	wire [4-1:0] node37680;
	wire [4-1:0] node37681;
	wire [4-1:0] node37685;
	wire [4-1:0] node37686;
	wire [4-1:0] node37689;
	wire [4-1:0] node37692;
	wire [4-1:0] node37693;
	wire [4-1:0] node37696;
	wire [4-1:0] node37699;
	wire [4-1:0] node37700;
	wire [4-1:0] node37701;
	wire [4-1:0] node37702;
	wire [4-1:0] node37703;
	wire [4-1:0] node37705;
	wire [4-1:0] node37708;
	wire [4-1:0] node37709;
	wire [4-1:0] node37713;
	wire [4-1:0] node37714;
	wire [4-1:0] node37715;
	wire [4-1:0] node37719;
	wire [4-1:0] node37720;
	wire [4-1:0] node37724;
	wire [4-1:0] node37725;
	wire [4-1:0] node37726;
	wire [4-1:0] node37729;
	wire [4-1:0] node37731;
	wire [4-1:0] node37734;
	wire [4-1:0] node37736;
	wire [4-1:0] node37739;
	wire [4-1:0] node37740;
	wire [4-1:0] node37741;
	wire [4-1:0] node37742;
	wire [4-1:0] node37743;
	wire [4-1:0] node37748;
	wire [4-1:0] node37749;
	wire [4-1:0] node37750;
	wire [4-1:0] node37754;
	wire [4-1:0] node37755;
	wire [4-1:0] node37759;
	wire [4-1:0] node37760;
	wire [4-1:0] node37762;
	wire [4-1:0] node37764;
	wire [4-1:0] node37767;
	wire [4-1:0] node37768;
	wire [4-1:0] node37770;
	wire [4-1:0] node37773;
	wire [4-1:0] node37775;
	wire [4-1:0] node37778;
	wire [4-1:0] node37779;
	wire [4-1:0] node37780;
	wire [4-1:0] node37781;
	wire [4-1:0] node37782;
	wire [4-1:0] node37783;
	wire [4-1:0] node37787;
	wire [4-1:0] node37788;
	wire [4-1:0] node37792;
	wire [4-1:0] node37793;
	wire [4-1:0] node37794;
	wire [4-1:0] node37795;
	wire [4-1:0] node37799;
	wire [4-1:0] node37800;
	wire [4-1:0] node37804;
	wire [4-1:0] node37805;
	wire [4-1:0] node37806;
	wire [4-1:0] node37810;
	wire [4-1:0] node37811;
	wire [4-1:0] node37814;
	wire [4-1:0] node37817;
	wire [4-1:0] node37818;
	wire [4-1:0] node37819;
	wire [4-1:0] node37820;
	wire [4-1:0] node37821;
	wire [4-1:0] node37824;
	wire [4-1:0] node37827;
	wire [4-1:0] node37828;
	wire [4-1:0] node37831;
	wire [4-1:0] node37834;
	wire [4-1:0] node37835;
	wire [4-1:0] node37836;
	wire [4-1:0] node37839;
	wire [4-1:0] node37842;
	wire [4-1:0] node37845;
	wire [4-1:0] node37846;
	wire [4-1:0] node37847;
	wire [4-1:0] node37848;
	wire [4-1:0] node37852;
	wire [4-1:0] node37853;
	wire [4-1:0] node37857;
	wire [4-1:0] node37858;
	wire [4-1:0] node37859;
	wire [4-1:0] node37863;
	wire [4-1:0] node37864;
	wire [4-1:0] node37867;
	wire [4-1:0] node37870;
	wire [4-1:0] node37871;
	wire [4-1:0] node37872;
	wire [4-1:0] node37873;
	wire [4-1:0] node37874;
	wire [4-1:0] node37878;
	wire [4-1:0] node37879;
	wire [4-1:0] node37880;
	wire [4-1:0] node37883;
	wire [4-1:0] node37887;
	wire [4-1:0] node37888;
	wire [4-1:0] node37889;
	wire [4-1:0] node37892;
	wire [4-1:0] node37894;
	wire [4-1:0] node37897;
	wire [4-1:0] node37898;
	wire [4-1:0] node37901;
	wire [4-1:0] node37904;
	wire [4-1:0] node37905;
	wire [4-1:0] node37906;
	wire [4-1:0] node37907;
	wire [4-1:0] node37908;
	wire [4-1:0] node37911;
	wire [4-1:0] node37914;
	wire [4-1:0] node37915;
	wire [4-1:0] node37919;
	wire [4-1:0] node37920;
	wire [4-1:0] node37923;
	wire [4-1:0] node37925;
	wire [4-1:0] node37928;
	wire [4-1:0] node37929;
	wire [4-1:0] node37930;
	wire [4-1:0] node37933;
	wire [4-1:0] node37936;
	wire [4-1:0] node37938;
	wire [4-1:0] node37939;
	wire [4-1:0] node37943;
	wire [4-1:0] node37944;
	wire [4-1:0] node37945;
	wire [4-1:0] node37946;
	wire [4-1:0] node37947;
	wire [4-1:0] node37948;
	wire [4-1:0] node37949;
	wire [4-1:0] node37950;
	wire [4-1:0] node37954;
	wire [4-1:0] node37956;
	wire [4-1:0] node37959;
	wire [4-1:0] node37960;
	wire [4-1:0] node37962;
	wire [4-1:0] node37966;
	wire [4-1:0] node37967;
	wire [4-1:0] node37968;
	wire [4-1:0] node37970;
	wire [4-1:0] node37973;
	wire [4-1:0] node37974;
	wire [4-1:0] node37978;
	wire [4-1:0] node37980;
	wire [4-1:0] node37982;
	wire [4-1:0] node37985;
	wire [4-1:0] node37986;
	wire [4-1:0] node37987;
	wire [4-1:0] node37989;
	wire [4-1:0] node37990;
	wire [4-1:0] node37993;
	wire [4-1:0] node37996;
	wire [4-1:0] node37997;
	wire [4-1:0] node37998;
	wire [4-1:0] node38002;
	wire [4-1:0] node38003;
	wire [4-1:0] node38006;
	wire [4-1:0] node38009;
	wire [4-1:0] node38010;
	wire [4-1:0] node38011;
	wire [4-1:0] node38012;
	wire [4-1:0] node38016;
	wire [4-1:0] node38017;
	wire [4-1:0] node38021;
	wire [4-1:0] node38022;
	wire [4-1:0] node38023;
	wire [4-1:0] node38027;
	wire [4-1:0] node38028;
	wire [4-1:0] node38032;
	wire [4-1:0] node38033;
	wire [4-1:0] node38034;
	wire [4-1:0] node38035;
	wire [4-1:0] node38036;
	wire [4-1:0] node38039;
	wire [4-1:0] node38042;
	wire [4-1:0] node38043;
	wire [4-1:0] node38045;
	wire [4-1:0] node38048;
	wire [4-1:0] node38050;
	wire [4-1:0] node38053;
	wire [4-1:0] node38054;
	wire [4-1:0] node38055;
	wire [4-1:0] node38058;
	wire [4-1:0] node38061;
	wire [4-1:0] node38062;
	wire [4-1:0] node38063;
	wire [4-1:0] node38066;
	wire [4-1:0] node38069;
	wire [4-1:0] node38070;
	wire [4-1:0] node38073;
	wire [4-1:0] node38076;
	wire [4-1:0] node38077;
	wire [4-1:0] node38078;
	wire [4-1:0] node38079;
	wire [4-1:0] node38081;
	wire [4-1:0] node38084;
	wire [4-1:0] node38085;
	wire [4-1:0] node38088;
	wire [4-1:0] node38091;
	wire [4-1:0] node38092;
	wire [4-1:0] node38095;
	wire [4-1:0] node38098;
	wire [4-1:0] node38099;
	wire [4-1:0] node38100;
	wire [4-1:0] node38101;
	wire [4-1:0] node38104;
	wire [4-1:0] node38108;
	wire [4-1:0] node38109;
	wire [4-1:0] node38110;
	wire [4-1:0] node38114;
	wire [4-1:0] node38115;
	wire [4-1:0] node38119;
	wire [4-1:0] node38120;
	wire [4-1:0] node38121;
	wire [4-1:0] node38122;
	wire [4-1:0] node38123;
	wire [4-1:0] node38124;
	wire [4-1:0] node38127;
	wire [4-1:0] node38130;
	wire [4-1:0] node38131;
	wire [4-1:0] node38132;
	wire [4-1:0] node38135;
	wire [4-1:0] node38138;
	wire [4-1:0] node38139;
	wire [4-1:0] node38142;
	wire [4-1:0] node38145;
	wire [4-1:0] node38146;
	wire [4-1:0] node38147;
	wire [4-1:0] node38149;
	wire [4-1:0] node38152;
	wire [4-1:0] node38154;
	wire [4-1:0] node38157;
	wire [4-1:0] node38158;
	wire [4-1:0] node38161;
	wire [4-1:0] node38163;
	wire [4-1:0] node38166;
	wire [4-1:0] node38167;
	wire [4-1:0] node38168;
	wire [4-1:0] node38170;
	wire [4-1:0] node38173;
	wire [4-1:0] node38174;
	wire [4-1:0] node38175;
	wire [4-1:0] node38179;
	wire [4-1:0] node38182;
	wire [4-1:0] node38183;
	wire [4-1:0] node38184;
	wire [4-1:0] node38188;
	wire [4-1:0] node38189;
	wire [4-1:0] node38190;
	wire [4-1:0] node38194;
	wire [4-1:0] node38195;
	wire [4-1:0] node38199;
	wire [4-1:0] node38200;
	wire [4-1:0] node38201;
	wire [4-1:0] node38202;
	wire [4-1:0] node38203;
	wire [4-1:0] node38204;
	wire [4-1:0] node38207;
	wire [4-1:0] node38210;
	wire [4-1:0] node38211;
	wire [4-1:0] node38214;
	wire [4-1:0] node38217;
	wire [4-1:0] node38218;
	wire [4-1:0] node38219;
	wire [4-1:0] node38222;
	wire [4-1:0] node38225;
	wire [4-1:0] node38226;
	wire [4-1:0] node38230;
	wire [4-1:0] node38231;
	wire [4-1:0] node38233;
	wire [4-1:0] node38234;
	wire [4-1:0] node38237;
	wire [4-1:0] node38240;
	wire [4-1:0] node38241;
	wire [4-1:0] node38242;
	wire [4-1:0] node38246;
	wire [4-1:0] node38247;
	wire [4-1:0] node38251;
	wire [4-1:0] node38252;
	wire [4-1:0] node38253;
	wire [4-1:0] node38255;
	wire [4-1:0] node38258;
	wire [4-1:0] node38259;
	wire [4-1:0] node38263;
	wire [4-1:0] node38264;
	wire [4-1:0] node38265;
	wire [4-1:0] node38268;
	wire [4-1:0] node38271;
	wire [4-1:0] node38272;
	wire [4-1:0] node38273;
	wire [4-1:0] node38277;
	wire [4-1:0] node38278;
	wire [4-1:0] node38281;
	wire [4-1:0] node38284;
	wire [4-1:0] node38285;
	wire [4-1:0] node38286;
	wire [4-1:0] node38287;
	wire [4-1:0] node38288;
	wire [4-1:0] node38289;
	wire [4-1:0] node38290;
	wire [4-1:0] node38291;
	wire [4-1:0] node38292;
	wire [4-1:0] node38295;
	wire [4-1:0] node38299;
	wire [4-1:0] node38300;
	wire [4-1:0] node38301;
	wire [4-1:0] node38304;
	wire [4-1:0] node38307;
	wire [4-1:0] node38308;
	wire [4-1:0] node38311;
	wire [4-1:0] node38314;
	wire [4-1:0] node38315;
	wire [4-1:0] node38316;
	wire [4-1:0] node38319;
	wire [4-1:0] node38322;
	wire [4-1:0] node38323;
	wire [4-1:0] node38324;
	wire [4-1:0] node38327;
	wire [4-1:0] node38330;
	wire [4-1:0] node38331;
	wire [4-1:0] node38334;
	wire [4-1:0] node38337;
	wire [4-1:0] node38338;
	wire [4-1:0] node38339;
	wire [4-1:0] node38340;
	wire [4-1:0] node38341;
	wire [4-1:0] node38344;
	wire [4-1:0] node38347;
	wire [4-1:0] node38349;
	wire [4-1:0] node38352;
	wire [4-1:0] node38353;
	wire [4-1:0] node38356;
	wire [4-1:0] node38359;
	wire [4-1:0] node38360;
	wire [4-1:0] node38361;
	wire [4-1:0] node38362;
	wire [4-1:0] node38365;
	wire [4-1:0] node38369;
	wire [4-1:0] node38370;
	wire [4-1:0] node38371;
	wire [4-1:0] node38374;
	wire [4-1:0] node38377;
	wire [4-1:0] node38378;
	wire [4-1:0] node38381;
	wire [4-1:0] node38384;
	wire [4-1:0] node38385;
	wire [4-1:0] node38386;
	wire [4-1:0] node38387;
	wire [4-1:0] node38388;
	wire [4-1:0] node38389;
	wire [4-1:0] node38392;
	wire [4-1:0] node38395;
	wire [4-1:0] node38396;
	wire [4-1:0] node38399;
	wire [4-1:0] node38402;
	wire [4-1:0] node38403;
	wire [4-1:0] node38404;
	wire [4-1:0] node38407;
	wire [4-1:0] node38410;
	wire [4-1:0] node38411;
	wire [4-1:0] node38415;
	wire [4-1:0] node38416;
	wire [4-1:0] node38418;
	wire [4-1:0] node38419;
	wire [4-1:0] node38423;
	wire [4-1:0] node38424;
	wire [4-1:0] node38425;
	wire [4-1:0] node38429;
	wire [4-1:0] node38430;
	wire [4-1:0] node38433;
	wire [4-1:0] node38436;
	wire [4-1:0] node38437;
	wire [4-1:0] node38438;
	wire [4-1:0] node38439;
	wire [4-1:0] node38441;
	wire [4-1:0] node38444;
	wire [4-1:0] node38445;
	wire [4-1:0] node38448;
	wire [4-1:0] node38451;
	wire [4-1:0] node38452;
	wire [4-1:0] node38453;
	wire [4-1:0] node38456;
	wire [4-1:0] node38459;
	wire [4-1:0] node38460;
	wire [4-1:0] node38464;
	wire [4-1:0] node38465;
	wire [4-1:0] node38466;
	wire [4-1:0] node38467;
	wire [4-1:0] node38470;
	wire [4-1:0] node38473;
	wire [4-1:0] node38474;
	wire [4-1:0] node38477;
	wire [4-1:0] node38480;
	wire [4-1:0] node38481;
	wire [4-1:0] node38484;
	wire [4-1:0] node38487;
	wire [4-1:0] node38488;
	wire [4-1:0] node38489;
	wire [4-1:0] node38490;
	wire [4-1:0] node38491;
	wire [4-1:0] node38492;
	wire [4-1:0] node38495;
	wire [4-1:0] node38498;
	wire [4-1:0] node38499;
	wire [4-1:0] node38500;
	wire [4-1:0] node38504;
	wire [4-1:0] node38507;
	wire [4-1:0] node38508;
	wire [4-1:0] node38509;
	wire [4-1:0] node38512;
	wire [4-1:0] node38513;
	wire [4-1:0] node38517;
	wire [4-1:0] node38518;
	wire [4-1:0] node38521;
	wire [4-1:0] node38522;
	wire [4-1:0] node38526;
	wire [4-1:0] node38527;
	wire [4-1:0] node38528;
	wire [4-1:0] node38529;
	wire [4-1:0] node38531;
	wire [4-1:0] node38534;
	wire [4-1:0] node38535;
	wire [4-1:0] node38538;
	wire [4-1:0] node38541;
	wire [4-1:0] node38542;
	wire [4-1:0] node38543;
	wire [4-1:0] node38546;
	wire [4-1:0] node38549;
	wire [4-1:0] node38550;
	wire [4-1:0] node38554;
	wire [4-1:0] node38555;
	wire [4-1:0] node38556;
	wire [4-1:0] node38557;
	wire [4-1:0] node38560;
	wire [4-1:0] node38563;
	wire [4-1:0] node38564;
	wire [4-1:0] node38567;
	wire [4-1:0] node38570;
	wire [4-1:0] node38571;
	wire [4-1:0] node38572;
	wire [4-1:0] node38575;
	wire [4-1:0] node38578;
	wire [4-1:0] node38579;
	wire [4-1:0] node38582;
	wire [4-1:0] node38585;
	wire [4-1:0] node38586;
	wire [4-1:0] node38587;
	wire [4-1:0] node38588;
	wire [4-1:0] node38589;
	wire [4-1:0] node38590;
	wire [4-1:0] node38593;
	wire [4-1:0] node38596;
	wire [4-1:0] node38597;
	wire [4-1:0] node38600;
	wire [4-1:0] node38603;
	wire [4-1:0] node38604;
	wire [4-1:0] node38605;
	wire [4-1:0] node38608;
	wire [4-1:0] node38611;
	wire [4-1:0] node38612;
	wire [4-1:0] node38615;
	wire [4-1:0] node38618;
	wire [4-1:0] node38619;
	wire [4-1:0] node38620;
	wire [4-1:0] node38622;
	wire [4-1:0] node38625;
	wire [4-1:0] node38626;
	wire [4-1:0] node38630;
	wire [4-1:0] node38631;
	wire [4-1:0] node38632;
	wire [4-1:0] node38635;
	wire [4-1:0] node38638;
	wire [4-1:0] node38639;
	wire [4-1:0] node38642;
	wire [4-1:0] node38645;
	wire [4-1:0] node38646;
	wire [4-1:0] node38647;
	wire [4-1:0] node38649;
	wire [4-1:0] node38651;
	wire [4-1:0] node38654;
	wire [4-1:0] node38655;
	wire [4-1:0] node38656;
	wire [4-1:0] node38659;
	wire [4-1:0] node38663;
	wire [4-1:0] node38664;
	wire [4-1:0] node38666;
	wire [4-1:0] node38667;
	wire [4-1:0] node38670;
	wire [4-1:0] node38673;
	wire [4-1:0] node38674;
	wire [4-1:0] node38675;
	wire [4-1:0] node38678;
	wire [4-1:0] node38681;
	wire [4-1:0] node38682;
	wire [4-1:0] node38686;
	wire [4-1:0] node38687;
	wire [4-1:0] node38688;
	wire [4-1:0] node38689;
	wire [4-1:0] node38690;
	wire [4-1:0] node38691;
	wire [4-1:0] node38692;
	wire [4-1:0] node38693;
	wire [4-1:0] node38696;
	wire [4-1:0] node38699;
	wire [4-1:0] node38700;
	wire [4-1:0] node38704;
	wire [4-1:0] node38705;
	wire [4-1:0] node38706;
	wire [4-1:0] node38709;
	wire [4-1:0] node38712;
	wire [4-1:0] node38713;
	wire [4-1:0] node38717;
	wire [4-1:0] node38718;
	wire [4-1:0] node38719;
	wire [4-1:0] node38720;
	wire [4-1:0] node38723;
	wire [4-1:0] node38726;
	wire [4-1:0] node38727;
	wire [4-1:0] node38731;
	wire [4-1:0] node38732;
	wire [4-1:0] node38733;
	wire [4-1:0] node38736;
	wire [4-1:0] node38739;
	wire [4-1:0] node38740;
	wire [4-1:0] node38743;
	wire [4-1:0] node38746;
	wire [4-1:0] node38747;
	wire [4-1:0] node38748;
	wire [4-1:0] node38749;
	wire [4-1:0] node38752;
	wire [4-1:0] node38755;
	wire [4-1:0] node38756;
	wire [4-1:0] node38759;
	wire [4-1:0] node38762;
	wire [4-1:0] node38763;
	wire [4-1:0] node38764;
	wire [4-1:0] node38766;
	wire [4-1:0] node38769;
	wire [4-1:0] node38770;
	wire [4-1:0] node38773;
	wire [4-1:0] node38776;
	wire [4-1:0] node38777;
	wire [4-1:0] node38778;
	wire [4-1:0] node38781;
	wire [4-1:0] node38784;
	wire [4-1:0] node38785;
	wire [4-1:0] node38788;
	wire [4-1:0] node38791;
	wire [4-1:0] node38792;
	wire [4-1:0] node38793;
	wire [4-1:0] node38794;
	wire [4-1:0] node38795;
	wire [4-1:0] node38798;
	wire [4-1:0] node38801;
	wire [4-1:0] node38802;
	wire [4-1:0] node38803;
	wire [4-1:0] node38806;
	wire [4-1:0] node38809;
	wire [4-1:0] node38810;
	wire [4-1:0] node38813;
	wire [4-1:0] node38816;
	wire [4-1:0] node38817;
	wire [4-1:0] node38818;
	wire [4-1:0] node38819;
	wire [4-1:0] node38823;
	wire [4-1:0] node38826;
	wire [4-1:0] node38827;
	wire [4-1:0] node38830;
	wire [4-1:0] node38832;
	wire [4-1:0] node38835;
	wire [4-1:0] node38836;
	wire [4-1:0] node38837;
	wire [4-1:0] node38838;
	wire [4-1:0] node38841;
	wire [4-1:0] node38844;
	wire [4-1:0] node38845;
	wire [4-1:0] node38848;
	wire [4-1:0] node38850;
	wire [4-1:0] node38853;
	wire [4-1:0] node38854;
	wire [4-1:0] node38855;
	wire [4-1:0] node38856;
	wire [4-1:0] node38860;
	wire [4-1:0] node38863;
	wire [4-1:0] node38864;
	wire [4-1:0] node38867;
	wire [4-1:0] node38869;
	wire [4-1:0] node38872;
	wire [4-1:0] node38873;
	wire [4-1:0] node38874;
	wire [4-1:0] node38875;
	wire [4-1:0] node38876;
	wire [4-1:0] node38877;
	wire [4-1:0] node38878;
	wire [4-1:0] node38881;
	wire [4-1:0] node38884;
	wire [4-1:0] node38886;
	wire [4-1:0] node38889;
	wire [4-1:0] node38890;
	wire [4-1:0] node38893;
	wire [4-1:0] node38894;
	wire [4-1:0] node38897;
	wire [4-1:0] node38900;
	wire [4-1:0] node38901;
	wire [4-1:0] node38902;
	wire [4-1:0] node38903;
	wire [4-1:0] node38906;
	wire [4-1:0] node38909;
	wire [4-1:0] node38910;
	wire [4-1:0] node38913;
	wire [4-1:0] node38916;
	wire [4-1:0] node38917;
	wire [4-1:0] node38918;
	wire [4-1:0] node38922;
	wire [4-1:0] node38923;
	wire [4-1:0] node38927;
	wire [4-1:0] node38928;
	wire [4-1:0] node38929;
	wire [4-1:0] node38930;
	wire [4-1:0] node38933;
	wire [4-1:0] node38936;
	wire [4-1:0] node38937;
	wire [4-1:0] node38939;
	wire [4-1:0] node38942;
	wire [4-1:0] node38944;
	wire [4-1:0] node38947;
	wire [4-1:0] node38948;
	wire [4-1:0] node38949;
	wire [4-1:0] node38950;
	wire [4-1:0] node38953;
	wire [4-1:0] node38956;
	wire [4-1:0] node38958;
	wire [4-1:0] node38961;
	wire [4-1:0] node38962;
	wire [4-1:0] node38963;
	wire [4-1:0] node38967;
	wire [4-1:0] node38969;
	wire [4-1:0] node38972;
	wire [4-1:0] node38973;
	wire [4-1:0] node38974;
	wire [4-1:0] node38975;
	wire [4-1:0] node38976;
	wire [4-1:0] node38977;
	wire [4-1:0] node38980;
	wire [4-1:0] node38983;
	wire [4-1:0] node38984;
	wire [4-1:0] node38987;
	wire [4-1:0] node38990;
	wire [4-1:0] node38991;
	wire [4-1:0] node38992;
	wire [4-1:0] node38995;
	wire [4-1:0] node38998;
	wire [4-1:0] node38999;
	wire [4-1:0] node39002;
	wire [4-1:0] node39005;
	wire [4-1:0] node39006;
	wire [4-1:0] node39007;
	wire [4-1:0] node39008;
	wire [4-1:0] node39011;
	wire [4-1:0] node39015;
	wire [4-1:0] node39016;
	wire [4-1:0] node39018;
	wire [4-1:0] node39021;
	wire [4-1:0] node39022;
	wire [4-1:0] node39025;
	wire [4-1:0] node39028;
	wire [4-1:0] node39029;
	wire [4-1:0] node39030;
	wire [4-1:0] node39031;
	wire [4-1:0] node39032;
	wire [4-1:0] node39035;
	wire [4-1:0] node39038;
	wire [4-1:0] node39039;
	wire [4-1:0] node39042;
	wire [4-1:0] node39045;
	wire [4-1:0] node39046;
	wire [4-1:0] node39047;
	wire [4-1:0] node39050;
	wire [4-1:0] node39053;
	wire [4-1:0] node39054;
	wire [4-1:0] node39057;
	wire [4-1:0] node39060;
	wire [4-1:0] node39061;
	wire [4-1:0] node39062;
	wire [4-1:0] node39063;
	wire [4-1:0] node39067;
	wire [4-1:0] node39068;
	wire [4-1:0] node39071;
	wire [4-1:0] node39074;
	wire [4-1:0] node39075;
	wire [4-1:0] node39078;
	wire [4-1:0] node39079;
	wire [4-1:0] node39082;
	wire [4-1:0] node39085;
	wire [4-1:0] node39086;
	wire [4-1:0] node39087;
	wire [4-1:0] node39088;
	wire [4-1:0] node39089;
	wire [4-1:0] node39090;
	wire [4-1:0] node39091;
	wire [4-1:0] node39092;
	wire [4-1:0] node39093;
	wire [4-1:0] node39096;
	wire [4-1:0] node39097;
	wire [4-1:0] node39101;
	wire [4-1:0] node39103;
	wire [4-1:0] node39105;
	wire [4-1:0] node39108;
	wire [4-1:0] node39109;
	wire [4-1:0] node39110;
	wire [4-1:0] node39111;
	wire [4-1:0] node39115;
	wire [4-1:0] node39116;
	wire [4-1:0] node39120;
	wire [4-1:0] node39121;
	wire [4-1:0] node39123;
	wire [4-1:0] node39126;
	wire [4-1:0] node39128;
	wire [4-1:0] node39131;
	wire [4-1:0] node39132;
	wire [4-1:0] node39133;
	wire [4-1:0] node39135;
	wire [4-1:0] node39136;
	wire [4-1:0] node39140;
	wire [4-1:0] node39141;
	wire [4-1:0] node39144;
	wire [4-1:0] node39145;
	wire [4-1:0] node39149;
	wire [4-1:0] node39150;
	wire [4-1:0] node39151;
	wire [4-1:0] node39152;
	wire [4-1:0] node39157;
	wire [4-1:0] node39158;
	wire [4-1:0] node39159;
	wire [4-1:0] node39163;
	wire [4-1:0] node39166;
	wire [4-1:0] node39167;
	wire [4-1:0] node39168;
	wire [4-1:0] node39169;
	wire [4-1:0] node39170;
	wire [4-1:0] node39173;
	wire [4-1:0] node39174;
	wire [4-1:0] node39178;
	wire [4-1:0] node39179;
	wire [4-1:0] node39180;
	wire [4-1:0] node39184;
	wire [4-1:0] node39185;
	wire [4-1:0] node39189;
	wire [4-1:0] node39190;
	wire [4-1:0] node39191;
	wire [4-1:0] node39192;
	wire [4-1:0] node39196;
	wire [4-1:0] node39199;
	wire [4-1:0] node39200;
	wire [4-1:0] node39203;
	wire [4-1:0] node39205;
	wire [4-1:0] node39208;
	wire [4-1:0] node39209;
	wire [4-1:0] node39210;
	wire [4-1:0] node39211;
	wire [4-1:0] node39213;
	wire [4-1:0] node39216;
	wire [4-1:0] node39219;
	wire [4-1:0] node39220;
	wire [4-1:0] node39223;
	wire [4-1:0] node39224;
	wire [4-1:0] node39228;
	wire [4-1:0] node39229;
	wire [4-1:0] node39230;
	wire [4-1:0] node39231;
	wire [4-1:0] node39235;
	wire [4-1:0] node39238;
	wire [4-1:0] node39239;
	wire [4-1:0] node39240;
	wire [4-1:0] node39244;
	wire [4-1:0] node39246;
	wire [4-1:0] node39249;
	wire [4-1:0] node39250;
	wire [4-1:0] node39251;
	wire [4-1:0] node39252;
	wire [4-1:0] node39253;
	wire [4-1:0] node39254;
	wire [4-1:0] node39256;
	wire [4-1:0] node39259;
	wire [4-1:0] node39262;
	wire [4-1:0] node39263;
	wire [4-1:0] node39264;
	wire [4-1:0] node39268;
	wire [4-1:0] node39271;
	wire [4-1:0] node39272;
	wire [4-1:0] node39273;
	wire [4-1:0] node39274;
	wire [4-1:0] node39277;
	wire [4-1:0] node39280;
	wire [4-1:0] node39281;
	wire [4-1:0] node39285;
	wire [4-1:0] node39286;
	wire [4-1:0] node39287;
	wire [4-1:0] node39291;
	wire [4-1:0] node39292;
	wire [4-1:0] node39296;
	wire [4-1:0] node39297;
	wire [4-1:0] node39298;
	wire [4-1:0] node39299;
	wire [4-1:0] node39300;
	wire [4-1:0] node39304;
	wire [4-1:0] node39305;
	wire [4-1:0] node39308;
	wire [4-1:0] node39311;
	wire [4-1:0] node39312;
	wire [4-1:0] node39313;
	wire [4-1:0] node39317;
	wire [4-1:0] node39318;
	wire [4-1:0] node39322;
	wire [4-1:0] node39323;
	wire [4-1:0] node39324;
	wire [4-1:0] node39327;
	wire [4-1:0] node39328;
	wire [4-1:0] node39331;
	wire [4-1:0] node39334;
	wire [4-1:0] node39335;
	wire [4-1:0] node39336;
	wire [4-1:0] node39340;
	wire [4-1:0] node39341;
	wire [4-1:0] node39345;
	wire [4-1:0] node39346;
	wire [4-1:0] node39347;
	wire [4-1:0] node39348;
	wire [4-1:0] node39349;
	wire [4-1:0] node39350;
	wire [4-1:0] node39353;
	wire [4-1:0] node39356;
	wire [4-1:0] node39357;
	wire [4-1:0] node39361;
	wire [4-1:0] node39362;
	wire [4-1:0] node39363;
	wire [4-1:0] node39366;
	wire [4-1:0] node39369;
	wire [4-1:0] node39370;
	wire [4-1:0] node39373;
	wire [4-1:0] node39376;
	wire [4-1:0] node39377;
	wire [4-1:0] node39378;
	wire [4-1:0] node39379;
	wire [4-1:0] node39383;
	wire [4-1:0] node39385;
	wire [4-1:0] node39388;
	wire [4-1:0] node39389;
	wire [4-1:0] node39390;
	wire [4-1:0] node39394;
	wire [4-1:0] node39397;
	wire [4-1:0] node39398;
	wire [4-1:0] node39399;
	wire [4-1:0] node39400;
	wire [4-1:0] node39403;
	wire [4-1:0] node39404;
	wire [4-1:0] node39407;
	wire [4-1:0] node39410;
	wire [4-1:0] node39411;
	wire [4-1:0] node39412;
	wire [4-1:0] node39415;
	wire [4-1:0] node39418;
	wire [4-1:0] node39419;
	wire [4-1:0] node39422;
	wire [4-1:0] node39425;
	wire [4-1:0] node39426;
	wire [4-1:0] node39427;
	wire [4-1:0] node39428;
	wire [4-1:0] node39432;
	wire [4-1:0] node39435;
	wire [4-1:0] node39436;
	wire [4-1:0] node39437;
	wire [4-1:0] node39441;
	wire [4-1:0] node39444;
	wire [4-1:0] node39445;
	wire [4-1:0] node39446;
	wire [4-1:0] node39447;
	wire [4-1:0] node39448;
	wire [4-1:0] node39449;
	wire [4-1:0] node39450;
	wire [4-1:0] node39452;
	wire [4-1:0] node39455;
	wire [4-1:0] node39456;
	wire [4-1:0] node39459;
	wire [4-1:0] node39462;
	wire [4-1:0] node39463;
	wire [4-1:0] node39466;
	wire [4-1:0] node39469;
	wire [4-1:0] node39470;
	wire [4-1:0] node39471;
	wire [4-1:0] node39473;
	wire [4-1:0] node39476;
	wire [4-1:0] node39477;
	wire [4-1:0] node39481;
	wire [4-1:0] node39483;
	wire [4-1:0] node39484;
	wire [4-1:0] node39488;
	wire [4-1:0] node39489;
	wire [4-1:0] node39490;
	wire [4-1:0] node39491;
	wire [4-1:0] node39494;
	wire [4-1:0] node39497;
	wire [4-1:0] node39498;
	wire [4-1:0] node39499;
	wire [4-1:0] node39503;
	wire [4-1:0] node39504;
	wire [4-1:0] node39507;
	wire [4-1:0] node39510;
	wire [4-1:0] node39511;
	wire [4-1:0] node39512;
	wire [4-1:0] node39514;
	wire [4-1:0] node39518;
	wire [4-1:0] node39519;
	wire [4-1:0] node39523;
	wire [4-1:0] node39524;
	wire [4-1:0] node39525;
	wire [4-1:0] node39526;
	wire [4-1:0] node39527;
	wire [4-1:0] node39530;
	wire [4-1:0] node39532;
	wire [4-1:0] node39535;
	wire [4-1:0] node39536;
	wire [4-1:0] node39537;
	wire [4-1:0] node39541;
	wire [4-1:0] node39543;
	wire [4-1:0] node39546;
	wire [4-1:0] node39547;
	wire [4-1:0] node39549;
	wire [4-1:0] node39551;
	wire [4-1:0] node39554;
	wire [4-1:0] node39555;
	wire [4-1:0] node39557;
	wire [4-1:0] node39560;
	wire [4-1:0] node39561;
	wire [4-1:0] node39565;
	wire [4-1:0] node39566;
	wire [4-1:0] node39567;
	wire [4-1:0] node39568;
	wire [4-1:0] node39569;
	wire [4-1:0] node39574;
	wire [4-1:0] node39575;
	wire [4-1:0] node39576;
	wire [4-1:0] node39580;
	wire [4-1:0] node39582;
	wire [4-1:0] node39585;
	wire [4-1:0] node39586;
	wire [4-1:0] node39588;
	wire [4-1:0] node39590;
	wire [4-1:0] node39593;
	wire [4-1:0] node39594;
	wire [4-1:0] node39598;
	wire [4-1:0] node39599;
	wire [4-1:0] node39600;
	wire [4-1:0] node39601;
	wire [4-1:0] node39602;
	wire [4-1:0] node39603;
	wire [4-1:0] node39605;
	wire [4-1:0] node39608;
	wire [4-1:0] node39609;
	wire [4-1:0] node39613;
	wire [4-1:0] node39614;
	wire [4-1:0] node39615;
	wire [4-1:0] node39618;
	wire [4-1:0] node39621;
	wire [4-1:0] node39623;
	wire [4-1:0] node39626;
	wire [4-1:0] node39627;
	wire [4-1:0] node39628;
	wire [4-1:0] node39629;
	wire [4-1:0] node39632;
	wire [4-1:0] node39635;
	wire [4-1:0] node39636;
	wire [4-1:0] node39639;
	wire [4-1:0] node39642;
	wire [4-1:0] node39643;
	wire [4-1:0] node39645;
	wire [4-1:0] node39648;
	wire [4-1:0] node39649;
	wire [4-1:0] node39653;
	wire [4-1:0] node39654;
	wire [4-1:0] node39655;
	wire [4-1:0] node39656;
	wire [4-1:0] node39659;
	wire [4-1:0] node39662;
	wire [4-1:0] node39663;
	wire [4-1:0] node39666;
	wire [4-1:0] node39669;
	wire [4-1:0] node39670;
	wire [4-1:0] node39671;
	wire [4-1:0] node39674;
	wire [4-1:0] node39677;
	wire [4-1:0] node39678;
	wire [4-1:0] node39679;
	wire [4-1:0] node39684;
	wire [4-1:0] node39685;
	wire [4-1:0] node39686;
	wire [4-1:0] node39687;
	wire [4-1:0] node39688;
	wire [4-1:0] node39689;
	wire [4-1:0] node39693;
	wire [4-1:0] node39696;
	wire [4-1:0] node39697;
	wire [4-1:0] node39700;
	wire [4-1:0] node39702;
	wire [4-1:0] node39705;
	wire [4-1:0] node39706;
	wire [4-1:0] node39707;
	wire [4-1:0] node39708;
	wire [4-1:0] node39711;
	wire [4-1:0] node39714;
	wire [4-1:0] node39715;
	wire [4-1:0] node39719;
	wire [4-1:0] node39720;
	wire [4-1:0] node39721;
	wire [4-1:0] node39724;
	wire [4-1:0] node39727;
	wire [4-1:0] node39728;
	wire [4-1:0] node39731;
	wire [4-1:0] node39734;
	wire [4-1:0] node39735;
	wire [4-1:0] node39736;
	wire [4-1:0] node39737;
	wire [4-1:0] node39738;
	wire [4-1:0] node39742;
	wire [4-1:0] node39743;
	wire [4-1:0] node39746;
	wire [4-1:0] node39749;
	wire [4-1:0] node39750;
	wire [4-1:0] node39752;
	wire [4-1:0] node39755;
	wire [4-1:0] node39756;
	wire [4-1:0] node39759;
	wire [4-1:0] node39762;
	wire [4-1:0] node39763;
	wire [4-1:0] node39764;
	wire [4-1:0] node39767;
	wire [4-1:0] node39770;
	wire [4-1:0] node39771;
	wire [4-1:0] node39772;
	wire [4-1:0] node39775;
	wire [4-1:0] node39778;
	wire [4-1:0] node39780;
	wire [4-1:0] node39783;
	wire [4-1:0] node39784;
	wire [4-1:0] node39785;
	wire [4-1:0] node39786;
	wire [4-1:0] node39787;
	wire [4-1:0] node39788;
	wire [4-1:0] node39789;
	wire [4-1:0] node39790;
	wire [4-1:0] node39792;
	wire [4-1:0] node39795;
	wire [4-1:0] node39796;
	wire [4-1:0] node39799;
	wire [4-1:0] node39802;
	wire [4-1:0] node39803;
	wire [4-1:0] node39804;
	wire [4-1:0] node39809;
	wire [4-1:0] node39810;
	wire [4-1:0] node39811;
	wire [4-1:0] node39812;
	wire [4-1:0] node39815;
	wire [4-1:0] node39818;
	wire [4-1:0] node39819;
	wire [4-1:0] node39822;
	wire [4-1:0] node39825;
	wire [4-1:0] node39826;
	wire [4-1:0] node39827;
	wire [4-1:0] node39830;
	wire [4-1:0] node39833;
	wire [4-1:0] node39834;
	wire [4-1:0] node39837;
	wire [4-1:0] node39840;
	wire [4-1:0] node39841;
	wire [4-1:0] node39842;
	wire [4-1:0] node39843;
	wire [4-1:0] node39846;
	wire [4-1:0] node39849;
	wire [4-1:0] node39850;
	wire [4-1:0] node39851;
	wire [4-1:0] node39854;
	wire [4-1:0] node39857;
	wire [4-1:0] node39858;
	wire [4-1:0] node39861;
	wire [4-1:0] node39864;
	wire [4-1:0] node39865;
	wire [4-1:0] node39866;
	wire [4-1:0] node39869;
	wire [4-1:0] node39872;
	wire [4-1:0] node39875;
	wire [4-1:0] node39876;
	wire [4-1:0] node39877;
	wire [4-1:0] node39878;
	wire [4-1:0] node39879;
	wire [4-1:0] node39880;
	wire [4-1:0] node39883;
	wire [4-1:0] node39886;
	wire [4-1:0] node39888;
	wire [4-1:0] node39891;
	wire [4-1:0] node39892;
	wire [4-1:0] node39893;
	wire [4-1:0] node39896;
	wire [4-1:0] node39899;
	wire [4-1:0] node39900;
	wire [4-1:0] node39903;
	wire [4-1:0] node39906;
	wire [4-1:0] node39907;
	wire [4-1:0] node39908;
	wire [4-1:0] node39909;
	wire [4-1:0] node39913;
	wire [4-1:0] node39914;
	wire [4-1:0] node39917;
	wire [4-1:0] node39920;
	wire [4-1:0] node39921;
	wire [4-1:0] node39922;
	wire [4-1:0] node39926;
	wire [4-1:0] node39927;
	wire [4-1:0] node39930;
	wire [4-1:0] node39933;
	wire [4-1:0] node39934;
	wire [4-1:0] node39935;
	wire [4-1:0] node39936;
	wire [4-1:0] node39939;
	wire [4-1:0] node39942;
	wire [4-1:0] node39945;
	wire [4-1:0] node39946;
	wire [4-1:0] node39947;
	wire [4-1:0] node39950;
	wire [4-1:0] node39953;
	wire [4-1:0] node39956;
	wire [4-1:0] node39957;
	wire [4-1:0] node39958;
	wire [4-1:0] node39959;
	wire [4-1:0] node39960;
	wire [4-1:0] node39961;
	wire [4-1:0] node39962;
	wire [4-1:0] node39965;
	wire [4-1:0] node39969;
	wire [4-1:0] node39971;
	wire [4-1:0] node39972;
	wire [4-1:0] node39975;
	wire [4-1:0] node39978;
	wire [4-1:0] node39979;
	wire [4-1:0] node39980;
	wire [4-1:0] node39981;
	wire [4-1:0] node39984;
	wire [4-1:0] node39987;
	wire [4-1:0] node39988;
	wire [4-1:0] node39991;
	wire [4-1:0] node39994;
	wire [4-1:0] node39996;
	wire [4-1:0] node39997;
	wire [4-1:0] node40000;
	wire [4-1:0] node40003;
	wire [4-1:0] node40004;
	wire [4-1:0] node40005;
	wire [4-1:0] node40006;
	wire [4-1:0] node40009;
	wire [4-1:0] node40012;
	wire [4-1:0] node40015;
	wire [4-1:0] node40016;
	wire [4-1:0] node40017;
	wire [4-1:0] node40020;
	wire [4-1:0] node40023;
	wire [4-1:0] node40026;
	wire [4-1:0] node40027;
	wire [4-1:0] node40028;
	wire [4-1:0] node40029;
	wire [4-1:0] node40030;
	wire [4-1:0] node40031;
	wire [4-1:0] node40034;
	wire [4-1:0] node40037;
	wire [4-1:0] node40038;
	wire [4-1:0] node40041;
	wire [4-1:0] node40044;
	wire [4-1:0] node40045;
	wire [4-1:0] node40046;
	wire [4-1:0] node40049;
	wire [4-1:0] node40052;
	wire [4-1:0] node40053;
	wire [4-1:0] node40056;
	wire [4-1:0] node40059;
	wire [4-1:0] node40060;
	wire [4-1:0] node40062;
	wire [4-1:0] node40063;
	wire [4-1:0] node40066;
	wire [4-1:0] node40069;
	wire [4-1:0] node40070;
	wire [4-1:0] node40073;
	wire [4-1:0] node40074;
	wire [4-1:0] node40077;
	wire [4-1:0] node40080;
	wire [4-1:0] node40081;
	wire [4-1:0] node40082;
	wire [4-1:0] node40083;
	wire [4-1:0] node40086;
	wire [4-1:0] node40089;
	wire [4-1:0] node40092;
	wire [4-1:0] node40093;
	wire [4-1:0] node40094;
	wire [4-1:0] node40097;
	wire [4-1:0] node40100;
	wire [4-1:0] node40103;
	wire [4-1:0] node40104;
	wire [4-1:0] node40105;
	wire [4-1:0] node40106;
	wire [4-1:0] node40107;
	wire [4-1:0] node40108;
	wire [4-1:0] node40109;
	wire [4-1:0] node40112;
	wire [4-1:0] node40115;
	wire [4-1:0] node40116;
	wire [4-1:0] node40117;
	wire [4-1:0] node40120;
	wire [4-1:0] node40123;
	wire [4-1:0] node40125;
	wire [4-1:0] node40128;
	wire [4-1:0] node40129;
	wire [4-1:0] node40130;
	wire [4-1:0] node40131;
	wire [4-1:0] node40135;
	wire [4-1:0] node40136;
	wire [4-1:0] node40139;
	wire [4-1:0] node40142;
	wire [4-1:0] node40143;
	wire [4-1:0] node40146;
	wire [4-1:0] node40149;
	wire [4-1:0] node40150;
	wire [4-1:0] node40151;
	wire [4-1:0] node40152;
	wire [4-1:0] node40155;
	wire [4-1:0] node40158;
	wire [4-1:0] node40159;
	wire [4-1:0] node40162;
	wire [4-1:0] node40165;
	wire [4-1:0] node40166;
	wire [4-1:0] node40167;
	wire [4-1:0] node40168;
	wire [4-1:0] node40171;
	wire [4-1:0] node40174;
	wire [4-1:0] node40175;
	wire [4-1:0] node40178;
	wire [4-1:0] node40181;
	wire [4-1:0] node40182;
	wire [4-1:0] node40183;
	wire [4-1:0] node40186;
	wire [4-1:0] node40189;
	wire [4-1:0] node40190;
	wire [4-1:0] node40193;
	wire [4-1:0] node40196;
	wire [4-1:0] node40197;
	wire [4-1:0] node40198;
	wire [4-1:0] node40199;
	wire [4-1:0] node40200;
	wire [4-1:0] node40202;
	wire [4-1:0] node40205;
	wire [4-1:0] node40206;
	wire [4-1:0] node40210;
	wire [4-1:0] node40211;
	wire [4-1:0] node40212;
	wire [4-1:0] node40216;
	wire [4-1:0] node40217;
	wire [4-1:0] node40221;
	wire [4-1:0] node40222;
	wire [4-1:0] node40223;
	wire [4-1:0] node40224;
	wire [4-1:0] node40228;
	wire [4-1:0] node40229;
	wire [4-1:0] node40233;
	wire [4-1:0] node40235;
	wire [4-1:0] node40236;
	wire [4-1:0] node40239;
	wire [4-1:0] node40242;
	wire [4-1:0] node40243;
	wire [4-1:0] node40244;
	wire [4-1:0] node40245;
	wire [4-1:0] node40246;
	wire [4-1:0] node40249;
	wire [4-1:0] node40252;
	wire [4-1:0] node40253;
	wire [4-1:0] node40256;
	wire [4-1:0] node40259;
	wire [4-1:0] node40260;
	wire [4-1:0] node40261;
	wire [4-1:0] node40265;
	wire [4-1:0] node40266;
	wire [4-1:0] node40269;
	wire [4-1:0] node40272;
	wire [4-1:0] node40273;
	wire [4-1:0] node40274;
	wire [4-1:0] node40277;
	wire [4-1:0] node40280;
	wire [4-1:0] node40281;
	wire [4-1:0] node40284;
	wire [4-1:0] node40287;
	wire [4-1:0] node40288;
	wire [4-1:0] node40289;
	wire [4-1:0] node40290;
	wire [4-1:0] node40291;
	wire [4-1:0] node40292;
	wire [4-1:0] node40294;
	wire [4-1:0] node40298;
	wire [4-1:0] node40299;
	wire [4-1:0] node40302;
	wire [4-1:0] node40304;
	wire [4-1:0] node40307;
	wire [4-1:0] node40308;
	wire [4-1:0] node40309;
	wire [4-1:0] node40313;
	wire [4-1:0] node40314;
	wire [4-1:0] node40315;
	wire [4-1:0] node40319;
	wire [4-1:0] node40322;
	wire [4-1:0] node40323;
	wire [4-1:0] node40324;
	wire [4-1:0] node40325;
	wire [4-1:0] node40326;
	wire [4-1:0] node40329;
	wire [4-1:0] node40332;
	wire [4-1:0] node40333;
	wire [4-1:0] node40336;
	wire [4-1:0] node40339;
	wire [4-1:0] node40340;
	wire [4-1:0] node40342;
	wire [4-1:0] node40346;
	wire [4-1:0] node40347;
	wire [4-1:0] node40350;
	wire [4-1:0] node40353;
	wire [4-1:0] node40354;
	wire [4-1:0] node40355;
	wire [4-1:0] node40356;
	wire [4-1:0] node40357;
	wire [4-1:0] node40358;
	wire [4-1:0] node40362;
	wire [4-1:0] node40365;
	wire [4-1:0] node40367;
	wire [4-1:0] node40370;
	wire [4-1:0] node40371;
	wire [4-1:0] node40372;
	wire [4-1:0] node40376;
	wire [4-1:0] node40377;
	wire [4-1:0] node40380;
	wire [4-1:0] node40383;
	wire [4-1:0] node40384;
	wire [4-1:0] node40385;
	wire [4-1:0] node40386;
	wire [4-1:0] node40387;
	wire [4-1:0] node40392;
	wire [4-1:0] node40393;
	wire [4-1:0] node40394;
	wire [4-1:0] node40399;
	wire [4-1:0] node40400;
	wire [4-1:0] node40401;
	wire [4-1:0] node40402;
	wire [4-1:0] node40407;
	wire [4-1:0] node40408;
	wire [4-1:0] node40409;
	wire [4-1:0] node40414;
	wire [4-1:0] node40415;
	wire [4-1:0] node40416;
	wire [4-1:0] node40417;
	wire [4-1:0] node40418;
	wire [4-1:0] node40419;
	wire [4-1:0] node40420;
	wire [4-1:0] node40421;
	wire [4-1:0] node40422;
	wire [4-1:0] node40425;
	wire [4-1:0] node40428;
	wire [4-1:0] node40429;
	wire [4-1:0] node40431;
	wire [4-1:0] node40434;
	wire [4-1:0] node40435;
	wire [4-1:0] node40438;
	wire [4-1:0] node40441;
	wire [4-1:0] node40442;
	wire [4-1:0] node40443;
	wire [4-1:0] node40444;
	wire [4-1:0] node40447;
	wire [4-1:0] node40450;
	wire [4-1:0] node40451;
	wire [4-1:0] node40452;
	wire [4-1:0] node40456;
	wire [4-1:0] node40457;
	wire [4-1:0] node40460;
	wire [4-1:0] node40463;
	wire [4-1:0] node40464;
	wire [4-1:0] node40467;
	wire [4-1:0] node40470;
	wire [4-1:0] node40471;
	wire [4-1:0] node40472;
	wire [4-1:0] node40475;
	wire [4-1:0] node40477;
	wire [4-1:0] node40480;
	wire [4-1:0] node40481;
	wire [4-1:0] node40482;
	wire [4-1:0] node40485;
	wire [4-1:0] node40488;
	wire [4-1:0] node40489;
	wire [4-1:0] node40492;
	wire [4-1:0] node40495;
	wire [4-1:0] node40496;
	wire [4-1:0] node40497;
	wire [4-1:0] node40498;
	wire [4-1:0] node40499;
	wire [4-1:0] node40502;
	wire [4-1:0] node40505;
	wire [4-1:0] node40506;
	wire [4-1:0] node40508;
	wire [4-1:0] node40509;
	wire [4-1:0] node40512;
	wire [4-1:0] node40515;
	wire [4-1:0] node40516;
	wire [4-1:0] node40517;
	wire [4-1:0] node40520;
	wire [4-1:0] node40523;
	wire [4-1:0] node40525;
	wire [4-1:0] node40528;
	wire [4-1:0] node40529;
	wire [4-1:0] node40532;
	wire [4-1:0] node40534;
	wire [4-1:0] node40537;
	wire [4-1:0] node40538;
	wire [4-1:0] node40539;
	wire [4-1:0] node40542;
	wire [4-1:0] node40544;
	wire [4-1:0] node40547;
	wire [4-1:0] node40548;
	wire [4-1:0] node40549;
	wire [4-1:0] node40552;
	wire [4-1:0] node40555;
	wire [4-1:0] node40556;
	wire [4-1:0] node40559;
	wire [4-1:0] node40562;
	wire [4-1:0] node40563;
	wire [4-1:0] node40564;
	wire [4-1:0] node40565;
	wire [4-1:0] node40568;
	wire [4-1:0] node40571;
	wire [4-1:0] node40572;
	wire [4-1:0] node40573;
	wire [4-1:0] node40574;
	wire [4-1:0] node40575;
	wire [4-1:0] node40576;
	wire [4-1:0] node40579;
	wire [4-1:0] node40582;
	wire [4-1:0] node40583;
	wire [4-1:0] node40587;
	wire [4-1:0] node40588;
	wire [4-1:0] node40591;
	wire [4-1:0] node40594;
	wire [4-1:0] node40595;
	wire [4-1:0] node40597;
	wire [4-1:0] node40598;
	wire [4-1:0] node40601;
	wire [4-1:0] node40604;
	wire [4-1:0] node40605;
	wire [4-1:0] node40608;
	wire [4-1:0] node40611;
	wire [4-1:0] node40612;
	wire [4-1:0] node40613;
	wire [4-1:0] node40614;
	wire [4-1:0] node40615;
	wire [4-1:0] node40618;
	wire [4-1:0] node40621;
	wire [4-1:0] node40622;
	wire [4-1:0] node40625;
	wire [4-1:0] node40628;
	wire [4-1:0] node40629;
	wire [4-1:0] node40632;
	wire [4-1:0] node40635;
	wire [4-1:0] node40636;
	wire [4-1:0] node40637;
	wire [4-1:0] node40640;
	wire [4-1:0] node40643;
	wire [4-1:0] node40645;
	wire [4-1:0] node40648;
	wire [4-1:0] node40649;
	wire [4-1:0] node40650;
	wire [4-1:0] node40651;
	wire [4-1:0] node40652;
	wire [4-1:0] node40654;
	wire [4-1:0] node40657;
	wire [4-1:0] node40658;
	wire [4-1:0] node40661;
	wire [4-1:0] node40664;
	wire [4-1:0] node40665;
	wire [4-1:0] node40666;
	wire [4-1:0] node40667;
	wire [4-1:0] node40670;
	wire [4-1:0] node40673;
	wire [4-1:0] node40674;
	wire [4-1:0] node40677;
	wire [4-1:0] node40680;
	wire [4-1:0] node40681;
	wire [4-1:0] node40682;
	wire [4-1:0] node40685;
	wire [4-1:0] node40688;
	wire [4-1:0] node40689;
	wire [4-1:0] node40692;
	wire [4-1:0] node40695;
	wire [4-1:0] node40696;
	wire [4-1:0] node40697;
	wire [4-1:0] node40698;
	wire [4-1:0] node40701;
	wire [4-1:0] node40704;
	wire [4-1:0] node40705;
	wire [4-1:0] node40706;
	wire [4-1:0] node40711;
	wire [4-1:0] node40712;
	wire [4-1:0] node40715;
	wire [4-1:0] node40718;
	wire [4-1:0] node40719;
	wire [4-1:0] node40720;
	wire [4-1:0] node40721;
	wire [4-1:0] node40722;
	wire [4-1:0] node40723;
	wire [4-1:0] node40728;
	wire [4-1:0] node40729;
	wire [4-1:0] node40732;
	wire [4-1:0] node40735;
	wire [4-1:0] node40736;
	wire [4-1:0] node40737;
	wire [4-1:0] node40739;
	wire [4-1:0] node40742;
	wire [4-1:0] node40743;
	wire [4-1:0] node40746;
	wire [4-1:0] node40749;
	wire [4-1:0] node40750;
	wire [4-1:0] node40752;
	wire [4-1:0] node40755;
	wire [4-1:0] node40756;
	wire [4-1:0] node40760;
	wire [4-1:0] node40761;
	wire [4-1:0] node40762;
	wire [4-1:0] node40763;
	wire [4-1:0] node40766;
	wire [4-1:0] node40769;
	wire [4-1:0] node40770;
	wire [4-1:0] node40773;
	wire [4-1:0] node40776;
	wire [4-1:0] node40777;
	wire [4-1:0] node40778;
	wire [4-1:0] node40781;
	wire [4-1:0] node40784;
	wire [4-1:0] node40785;
	wire [4-1:0] node40788;
	wire [4-1:0] node40791;
	wire [4-1:0] node40792;
	wire [4-1:0] node40793;
	wire [4-1:0] node40794;
	wire [4-1:0] node40795;
	wire [4-1:0] node40796;
	wire [4-1:0] node40797;
	wire [4-1:0] node40799;
	wire [4-1:0] node40802;
	wire [4-1:0] node40803;
	wire [4-1:0] node40804;
	wire [4-1:0] node40808;
	wire [4-1:0] node40809;
	wire [4-1:0] node40812;
	wire [4-1:0] node40815;
	wire [4-1:0] node40816;
	wire [4-1:0] node40817;
	wire [4-1:0] node40820;
	wire [4-1:0] node40823;
	wire [4-1:0] node40824;
	wire [4-1:0] node40827;
	wire [4-1:0] node40830;
	wire [4-1:0] node40831;
	wire [4-1:0] node40832;
	wire [4-1:0] node40833;
	wire [4-1:0] node40836;
	wire [4-1:0] node40839;
	wire [4-1:0] node40840;
	wire [4-1:0] node40841;
	wire [4-1:0] node40844;
	wire [4-1:0] node40847;
	wire [4-1:0] node40848;
	wire [4-1:0] node40851;
	wire [4-1:0] node40854;
	wire [4-1:0] node40855;
	wire [4-1:0] node40856;
	wire [4-1:0] node40859;
	wire [4-1:0] node40862;
	wire [4-1:0] node40863;
	wire [4-1:0] node40864;
	wire [4-1:0] node40867;
	wire [4-1:0] node40870;
	wire [4-1:0] node40871;
	wire [4-1:0] node40874;
	wire [4-1:0] node40877;
	wire [4-1:0] node40878;
	wire [4-1:0] node40879;
	wire [4-1:0] node40880;
	wire [4-1:0] node40881;
	wire [4-1:0] node40884;
	wire [4-1:0] node40887;
	wire [4-1:0] node40888;
	wire [4-1:0] node40891;
	wire [4-1:0] node40894;
	wire [4-1:0] node40895;
	wire [4-1:0] node40896;
	wire [4-1:0] node40899;
	wire [4-1:0] node40902;
	wire [4-1:0] node40903;
	wire [4-1:0] node40906;
	wire [4-1:0] node40909;
	wire [4-1:0] node40910;
	wire [4-1:0] node40911;
	wire [4-1:0] node40912;
	wire [4-1:0] node40913;
	wire [4-1:0] node40916;
	wire [4-1:0] node40919;
	wire [4-1:0] node40920;
	wire [4-1:0] node40923;
	wire [4-1:0] node40926;
	wire [4-1:0] node40927;
	wire [4-1:0] node40928;
	wire [4-1:0] node40931;
	wire [4-1:0] node40934;
	wire [4-1:0] node40935;
	wire [4-1:0] node40938;
	wire [4-1:0] node40941;
	wire [4-1:0] node40942;
	wire [4-1:0] node40943;
	wire [4-1:0] node40944;
	wire [4-1:0] node40947;
	wire [4-1:0] node40950;
	wire [4-1:0] node40951;
	wire [4-1:0] node40954;
	wire [4-1:0] node40957;
	wire [4-1:0] node40958;
	wire [4-1:0] node40959;
	wire [4-1:0] node40962;
	wire [4-1:0] node40965;
	wire [4-1:0] node40967;
	wire [4-1:0] node40970;
	wire [4-1:0] node40971;
	wire [4-1:0] node40972;
	wire [4-1:0] node40973;
	wire [4-1:0] node40974;
	wire [4-1:0] node40977;
	wire [4-1:0] node40980;
	wire [4-1:0] node40981;
	wire [4-1:0] node40983;
	wire [4-1:0] node40984;
	wire [4-1:0] node40987;
	wire [4-1:0] node40990;
	wire [4-1:0] node40991;
	wire [4-1:0] node40992;
	wire [4-1:0] node40996;
	wire [4-1:0] node40997;
	wire [4-1:0] node41001;
	wire [4-1:0] node41002;
	wire [4-1:0] node41003;
	wire [4-1:0] node41004;
	wire [4-1:0] node41005;
	wire [4-1:0] node41008;
	wire [4-1:0] node41011;
	wire [4-1:0] node41012;
	wire [4-1:0] node41016;
	wire [4-1:0] node41018;
	wire [4-1:0] node41021;
	wire [4-1:0] node41022;
	wire [4-1:0] node41025;
	wire [4-1:0] node41028;
	wire [4-1:0] node41029;
	wire [4-1:0] node41030;
	wire [4-1:0] node41031;
	wire [4-1:0] node41034;
	wire [4-1:0] node41037;
	wire [4-1:0] node41038;
	wire [4-1:0] node41039;
	wire [4-1:0] node41042;
	wire [4-1:0] node41045;
	wire [4-1:0] node41046;
	wire [4-1:0] node41050;
	wire [4-1:0] node41051;
	wire [4-1:0] node41052;
	wire [4-1:0] node41055;
	wire [4-1:0] node41058;
	wire [4-1:0] node41059;
	wire [4-1:0] node41061;
	wire [4-1:0] node41062;
	wire [4-1:0] node41066;
	wire [4-1:0] node41068;
	wire [4-1:0] node41069;
	wire [4-1:0] node41072;
	wire [4-1:0] node41075;
	wire [4-1:0] node41076;
	wire [4-1:0] node41077;
	wire [4-1:0] node41078;
	wire [4-1:0] node41079;
	wire [4-1:0] node41080;
	wire [4-1:0] node41083;
	wire [4-1:0] node41087;
	wire [4-1:0] node41088;
	wire [4-1:0] node41089;
	wire [4-1:0] node41092;
	wire [4-1:0] node41096;
	wire [4-1:0] node41097;
	wire [4-1:0] node41098;
	wire [4-1:0] node41099;
	wire [4-1:0] node41102;
	wire [4-1:0] node41106;
	wire [4-1:0] node41107;
	wire [4-1:0] node41108;
	wire [4-1:0] node41111;
	wire [4-1:0] node41115;
	wire [4-1:0] node41116;
	wire [4-1:0] node41117;
	wire [4-1:0] node41118;
	wire [4-1:0] node41119;
	wire [4-1:0] node41120;
	wire [4-1:0] node41123;
	wire [4-1:0] node41127;
	wire [4-1:0] node41128;
	wire [4-1:0] node41129;
	wire [4-1:0] node41132;
	wire [4-1:0] node41136;
	wire [4-1:0] node41137;
	wire [4-1:0] node41138;
	wire [4-1:0] node41139;
	wire [4-1:0] node41142;
	wire [4-1:0] node41146;
	wire [4-1:0] node41147;
	wire [4-1:0] node41148;
	wire [4-1:0] node41151;
	wire [4-1:0] node41155;
	wire [4-1:0] node41156;
	wire [4-1:0] node41157;
	wire [4-1:0] node41158;
	wire [4-1:0] node41159;
	wire [4-1:0] node41160;
	wire [4-1:0] node41163;
	wire [4-1:0] node41166;
	wire [4-1:0] node41167;
	wire [4-1:0] node41170;
	wire [4-1:0] node41174;
	wire [4-1:0] node41175;
	wire [4-1:0] node41176;
	wire [4-1:0] node41177;
	wire [4-1:0] node41180;
	wire [4-1:0] node41183;
	wire [4-1:0] node41184;
	wire [4-1:0] node41187;
	wire [4-1:0] node41191;
	wire [4-1:0] node41192;
	wire [4-1:0] node41193;
	wire [4-1:0] node41194;
	wire [4-1:0] node41197;
	wire [4-1:0] node41201;
	wire [4-1:0] node41202;
	wire [4-1:0] node41203;
	wire [4-1:0] node41205;
	wire [4-1:0] node41208;
	wire [4-1:0] node41209;
	wire [4-1:0] node41212;
	wire [4-1:0] node41216;
	wire [4-1:0] node41217;
	wire [4-1:0] node41218;
	wire [4-1:0] node41219;
	wire [4-1:0] node41220;
	wire [4-1:0] node41221;
	wire [4-1:0] node41222;
	wire [4-1:0] node41223;
	wire [4-1:0] node41225;
	wire [4-1:0] node41228;
	wire [4-1:0] node41230;
	wire [4-1:0] node41233;
	wire [4-1:0] node41234;
	wire [4-1:0] node41235;
	wire [4-1:0] node41236;
	wire [4-1:0] node41239;
	wire [4-1:0] node41242;
	wire [4-1:0] node41243;
	wire [4-1:0] node41246;
	wire [4-1:0] node41249;
	wire [4-1:0] node41250;
	wire [4-1:0] node41253;
	wire [4-1:0] node41255;
	wire [4-1:0] node41258;
	wire [4-1:0] node41259;
	wire [4-1:0] node41260;
	wire [4-1:0] node41261;
	wire [4-1:0] node41263;
	wire [4-1:0] node41266;
	wire [4-1:0] node41267;
	wire [4-1:0] node41270;
	wire [4-1:0] node41273;
	wire [4-1:0] node41274;
	wire [4-1:0] node41275;
	wire [4-1:0] node41278;
	wire [4-1:0] node41281;
	wire [4-1:0] node41282;
	wire [4-1:0] node41285;
	wire [4-1:0] node41288;
	wire [4-1:0] node41289;
	wire [4-1:0] node41290;
	wire [4-1:0] node41292;
	wire [4-1:0] node41295;
	wire [4-1:0] node41296;
	wire [4-1:0] node41299;
	wire [4-1:0] node41302;
	wire [4-1:0] node41304;
	wire [4-1:0] node41307;
	wire [4-1:0] node41308;
	wire [4-1:0] node41309;
	wire [4-1:0] node41310;
	wire [4-1:0] node41311;
	wire [4-1:0] node41312;
	wire [4-1:0] node41315;
	wire [4-1:0] node41318;
	wire [4-1:0] node41319;
	wire [4-1:0] node41322;
	wire [4-1:0] node41325;
	wire [4-1:0] node41326;
	wire [4-1:0] node41329;
	wire [4-1:0] node41332;
	wire [4-1:0] node41333;
	wire [4-1:0] node41334;
	wire [4-1:0] node41335;
	wire [4-1:0] node41338;
	wire [4-1:0] node41342;
	wire [4-1:0] node41343;
	wire [4-1:0] node41344;
	wire [4-1:0] node41347;
	wire [4-1:0] node41350;
	wire [4-1:0] node41351;
	wire [4-1:0] node41354;
	wire [4-1:0] node41357;
	wire [4-1:0] node41358;
	wire [4-1:0] node41359;
	wire [4-1:0] node41361;
	wire [4-1:0] node41364;
	wire [4-1:0] node41365;
	wire [4-1:0] node41368;
	wire [4-1:0] node41371;
	wire [4-1:0] node41372;
	wire [4-1:0] node41373;
	wire [4-1:0] node41376;
	wire [4-1:0] node41379;
	wire [4-1:0] node41380;
	wire [4-1:0] node41383;
	wire [4-1:0] node41386;
	wire [4-1:0] node41387;
	wire [4-1:0] node41388;
	wire [4-1:0] node41391;
	wire [4-1:0] node41394;
	wire [4-1:0] node41395;
	wire [4-1:0] node41396;
	wire [4-1:0] node41397;
	wire [4-1:0] node41400;
	wire [4-1:0] node41403;
	wire [4-1:0] node41404;
	wire [4-1:0] node41405;
	wire [4-1:0] node41409;
	wire [4-1:0] node41410;
	wire [4-1:0] node41411;
	wire [4-1:0] node41414;
	wire [4-1:0] node41417;
	wire [4-1:0] node41418;
	wire [4-1:0] node41422;
	wire [4-1:0] node41423;
	wire [4-1:0] node41426;
	wire [4-1:0] node41429;
	wire [4-1:0] node41430;
	wire [4-1:0] node41431;
	wire [4-1:0] node41432;
	wire [4-1:0] node41433;
	wire [4-1:0] node41436;
	wire [4-1:0] node41440;
	wire [4-1:0] node41441;
	wire [4-1:0] node41442;
	wire [4-1:0] node41443;
	wire [4-1:0] node41444;
	wire [4-1:0] node41445;
	wire [4-1:0] node41448;
	wire [4-1:0] node41451;
	wire [4-1:0] node41452;
	wire [4-1:0] node41455;
	wire [4-1:0] node41458;
	wire [4-1:0] node41459;
	wire [4-1:0] node41462;
	wire [4-1:0] node41465;
	wire [4-1:0] node41466;
	wire [4-1:0] node41469;
	wire [4-1:0] node41473;
	wire [4-1:0] node41474;
	wire [4-1:0] node41475;
	wire [4-1:0] node41476;
	wire [4-1:0] node41477;
	wire [4-1:0] node41478;
	wire [4-1:0] node41481;
	wire [4-1:0] node41484;
	wire [4-1:0] node41485;
	wire [4-1:0] node41488;
	wire [4-1:0] node41491;
	wire [4-1:0] node41492;
	wire [4-1:0] node41493;
	wire [4-1:0] node41496;
	wire [4-1:0] node41499;
	wire [4-1:0] node41500;
	wire [4-1:0] node41503;
	wire [4-1:0] node41507;
	wire [4-1:0] node41508;
	wire [4-1:0] node41509;
	wire [4-1:0] node41512;
	wire [4-1:0] node41516;
	wire [4-1:0] node41517;
	wire [4-1:0] node41518;
	wire [4-1:0] node41519;
	wire [4-1:0] node41520;
	wire [4-1:0] node41521;
	wire [4-1:0] node41522;
	wire [4-1:0] node41523;
	wire [4-1:0] node41526;
	wire [4-1:0] node41529;
	wire [4-1:0] node41530;
	wire [4-1:0] node41533;
	wire [4-1:0] node41536;
	wire [4-1:0] node41537;
	wire [4-1:0] node41540;
	wire [4-1:0] node41543;
	wire [4-1:0] node41544;
	wire [4-1:0] node41545;
	wire [4-1:0] node41547;
	wire [4-1:0] node41550;
	wire [4-1:0] node41551;
	wire [4-1:0] node41555;
	wire [4-1:0] node41556;
	wire [4-1:0] node41557;
	wire [4-1:0] node41561;
	wire [4-1:0] node41562;
	wire [4-1:0] node41566;
	wire [4-1:0] node41567;
	wire [4-1:0] node41568;
	wire [4-1:0] node41569;
	wire [4-1:0] node41573;
	wire [4-1:0] node41574;
	wire [4-1:0] node41578;
	wire [4-1:0] node41579;
	wire [4-1:0] node41581;
	wire [4-1:0] node41584;
	wire [4-1:0] node41586;
	wire [4-1:0] node41589;
	wire [4-1:0] node41590;
	wire [4-1:0] node41591;
	wire [4-1:0] node41592;
	wire [4-1:0] node41593;
	wire [4-1:0] node41594;
	wire [4-1:0] node41595;
	wire [4-1:0] node41598;
	wire [4-1:0] node41601;
	wire [4-1:0] node41602;
	wire [4-1:0] node41605;
	wire [4-1:0] node41608;
	wire [4-1:0] node41609;
	wire [4-1:0] node41612;
	wire [4-1:0] node41615;
	wire [4-1:0] node41616;
	wire [4-1:0] node41617;
	wire [4-1:0] node41621;
	wire [4-1:0] node41622;
	wire [4-1:0] node41625;
	wire [4-1:0] node41628;
	wire [4-1:0] node41629;
	wire [4-1:0] node41632;
	wire [4-1:0] node41635;
	wire [4-1:0] node41636;
	wire [4-1:0] node41637;
	wire [4-1:0] node41638;
	wire [4-1:0] node41639;
	wire [4-1:0] node41642;
	wire [4-1:0] node41645;
	wire [4-1:0] node41646;
	wire [4-1:0] node41649;
	wire [4-1:0] node41652;
	wire [4-1:0] node41653;
	wire [4-1:0] node41654;
	wire [4-1:0] node41657;
	wire [4-1:0] node41660;
	wire [4-1:0] node41661;
	wire [4-1:0] node41664;
	wire [4-1:0] node41667;
	wire [4-1:0] node41668;
	wire [4-1:0] node41669;
	wire [4-1:0] node41670;
	wire [4-1:0] node41671;
	wire [4-1:0] node41674;
	wire [4-1:0] node41677;
	wire [4-1:0] node41678;
	wire [4-1:0] node41681;
	wire [4-1:0] node41684;
	wire [4-1:0] node41685;
	wire [4-1:0] node41689;
	wire [4-1:0] node41690;
	wire [4-1:0] node41691;
	wire [4-1:0] node41694;
	wire [4-1:0] node41697;
	wire [4-1:0] node41698;
	wire [4-1:0] node41699;
	wire [4-1:0] node41703;
	wire [4-1:0] node41704;
	wire [4-1:0] node41707;
	wire [4-1:0] node41710;
	wire [4-1:0] node41711;
	wire [4-1:0] node41712;
	wire [4-1:0] node41713;
	wire [4-1:0] node41714;
	wire [4-1:0] node41715;
	wire [4-1:0] node41718;
	wire [4-1:0] node41721;
	wire [4-1:0] node41722;
	wire [4-1:0] node41724;
	wire [4-1:0] node41725;
	wire [4-1:0] node41728;
	wire [4-1:0] node41731;
	wire [4-1:0] node41732;
	wire [4-1:0] node41733;
	wire [4-1:0] node41736;
	wire [4-1:0] node41739;
	wire [4-1:0] node41740;
	wire [4-1:0] node41743;
	wire [4-1:0] node41746;
	wire [4-1:0] node41747;
	wire [4-1:0] node41748;
	wire [4-1:0] node41751;
	wire [4-1:0] node41754;
	wire [4-1:0] node41755;
	wire [4-1:0] node41758;
	wire [4-1:0] node41761;
	wire [4-1:0] node41762;
	wire [4-1:0] node41765;
	wire [4-1:0] node41768;
	wire [4-1:0] node41769;
	wire [4-1:0] node41770;
	wire [4-1:0] node41771;
	wire [4-1:0] node41772;
	wire [4-1:0] node41775;
	wire [4-1:0] node41778;
	wire [4-1:0] node41779;
	wire [4-1:0] node41780;
	wire [4-1:0] node41783;
	wire [4-1:0] node41786;
	wire [4-1:0] node41787;
	wire [4-1:0] node41790;
	wire [4-1:0] node41793;
	wire [4-1:0] node41794;
	wire [4-1:0] node41795;
	wire [4-1:0] node41796;
	wire [4-1:0] node41799;
	wire [4-1:0] node41802;
	wire [4-1:0] node41803;
	wire [4-1:0] node41807;
	wire [4-1:0] node41808;
	wire [4-1:0] node41811;
	wire [4-1:0] node41814;
	wire [4-1:0] node41815;
	wire [4-1:0] node41818;
	wire [4-1:0] node41821;
	wire [4-1:0] node41822;
	wire [4-1:0] node41823;
	wire [4-1:0] node41824;
	wire [4-1:0] node41825;
	wire [4-1:0] node41826;
	wire [4-1:0] node41827;
	wire [4-1:0] node41828;
	wire [4-1:0] node41829;
	wire [4-1:0] node41830;
	wire [4-1:0] node41831;
	wire [4-1:0] node41832;
	wire [4-1:0] node41836;
	wire [4-1:0] node41837;
	wire [4-1:0] node41840;
	wire [4-1:0] node41843;
	wire [4-1:0] node41844;
	wire [4-1:0] node41847;
	wire [4-1:0] node41850;
	wire [4-1:0] node41851;
	wire [4-1:0] node41852;
	wire [4-1:0] node41853;
	wire [4-1:0] node41856;
	wire [4-1:0] node41859;
	wire [4-1:0] node41860;
	wire [4-1:0] node41863;
	wire [4-1:0] node41866;
	wire [4-1:0] node41867;
	wire [4-1:0] node41868;
	wire [4-1:0] node41871;
	wire [4-1:0] node41874;
	wire [4-1:0] node41875;
	wire [4-1:0] node41878;
	wire [4-1:0] node41881;
	wire [4-1:0] node41882;
	wire [4-1:0] node41883;
	wire [4-1:0] node41885;
	wire [4-1:0] node41886;
	wire [4-1:0] node41889;
	wire [4-1:0] node41892;
	wire [4-1:0] node41893;
	wire [4-1:0] node41894;
	wire [4-1:0] node41897;
	wire [4-1:0] node41900;
	wire [4-1:0] node41901;
	wire [4-1:0] node41904;
	wire [4-1:0] node41907;
	wire [4-1:0] node41908;
	wire [4-1:0] node41909;
	wire [4-1:0] node41911;
	wire [4-1:0] node41914;
	wire [4-1:0] node41916;
	wire [4-1:0] node41919;
	wire [4-1:0] node41920;
	wire [4-1:0] node41923;
	wire [4-1:0] node41925;
	wire [4-1:0] node41928;
	wire [4-1:0] node41929;
	wire [4-1:0] node41930;
	wire [4-1:0] node41931;
	wire [4-1:0] node41932;
	wire [4-1:0] node41935;
	wire [4-1:0] node41937;
	wire [4-1:0] node41940;
	wire [4-1:0] node41941;
	wire [4-1:0] node41943;
	wire [4-1:0] node41947;
	wire [4-1:0] node41948;
	wire [4-1:0] node41949;
	wire [4-1:0] node41950;
	wire [4-1:0] node41953;
	wire [4-1:0] node41956;
	wire [4-1:0] node41957;
	wire [4-1:0] node41961;
	wire [4-1:0] node41962;
	wire [4-1:0] node41965;
	wire [4-1:0] node41968;
	wire [4-1:0] node41969;
	wire [4-1:0] node41970;
	wire [4-1:0] node41971;
	wire [4-1:0] node41972;
	wire [4-1:0] node41976;
	wire [4-1:0] node41977;
	wire [4-1:0] node41981;
	wire [4-1:0] node41982;
	wire [4-1:0] node41983;
	wire [4-1:0] node41987;
	wire [4-1:0] node41988;
	wire [4-1:0] node41992;
	wire [4-1:0] node41993;
	wire [4-1:0] node41994;
	wire [4-1:0] node41996;
	wire [4-1:0] node41999;
	wire [4-1:0] node42000;
	wire [4-1:0] node42004;
	wire [4-1:0] node42005;
	wire [4-1:0] node42009;
	wire [4-1:0] node42010;
	wire [4-1:0] node42011;
	wire [4-1:0] node42012;
	wire [4-1:0] node42013;
	wire [4-1:0] node42014;
	wire [4-1:0] node42016;
	wire [4-1:0] node42019;
	wire [4-1:0] node42022;
	wire [4-1:0] node42023;
	wire [4-1:0] node42027;
	wire [4-1:0] node42028;
	wire [4-1:0] node42029;
	wire [4-1:0] node42030;
	wire [4-1:0] node42034;
	wire [4-1:0] node42035;
	wire [4-1:0] node42039;
	wire [4-1:0] node42040;
	wire [4-1:0] node42043;
	wire [4-1:0] node42044;
	wire [4-1:0] node42048;
	wire [4-1:0] node42049;
	wire [4-1:0] node42050;
	wire [4-1:0] node42051;
	wire [4-1:0] node42054;
	wire [4-1:0] node42057;
	wire [4-1:0] node42058;
	wire [4-1:0] node42062;
	wire [4-1:0] node42063;
	wire [4-1:0] node42064;
	wire [4-1:0] node42065;
	wire [4-1:0] node42069;
	wire [4-1:0] node42070;
	wire [4-1:0] node42074;
	wire [4-1:0] node42075;
	wire [4-1:0] node42076;
	wire [4-1:0] node42080;
	wire [4-1:0] node42081;
	wire [4-1:0] node42085;
	wire [4-1:0] node42086;
	wire [4-1:0] node42087;
	wire [4-1:0] node42088;
	wire [4-1:0] node42089;
	wire [4-1:0] node42090;
	wire [4-1:0] node42094;
	wire [4-1:0] node42097;
	wire [4-1:0] node42098;
	wire [4-1:0] node42099;
	wire [4-1:0] node42103;
	wire [4-1:0] node42106;
	wire [4-1:0] node42107;
	wire [4-1:0] node42108;
	wire [4-1:0] node42109;
	wire [4-1:0] node42113;
	wire [4-1:0] node42116;
	wire [4-1:0] node42117;
	wire [4-1:0] node42118;
	wire [4-1:0] node42122;
	wire [4-1:0] node42125;
	wire [4-1:0] node42126;
	wire [4-1:0] node42127;
	wire [4-1:0] node42128;
	wire [4-1:0] node42131;
	wire [4-1:0] node42134;
	wire [4-1:0] node42135;
	wire [4-1:0] node42136;
	wire [4-1:0] node42139;
	wire [4-1:0] node42142;
	wire [4-1:0] node42143;
	wire [4-1:0] node42146;
	wire [4-1:0] node42149;
	wire [4-1:0] node42150;
	wire [4-1:0] node42151;
	wire [4-1:0] node42152;
	wire [4-1:0] node42155;
	wire [4-1:0] node42158;
	wire [4-1:0] node42159;
	wire [4-1:0] node42163;
	wire [4-1:0] node42164;
	wire [4-1:0] node42165;
	wire [4-1:0] node42168;
	wire [4-1:0] node42171;
	wire [4-1:0] node42172;
	wire [4-1:0] node42176;
	wire [4-1:0] node42177;
	wire [4-1:0] node42178;
	wire [4-1:0] node42179;
	wire [4-1:0] node42180;
	wire [4-1:0] node42181;
	wire [4-1:0] node42182;
	wire [4-1:0] node42183;
	wire [4-1:0] node42187;
	wire [4-1:0] node42188;
	wire [4-1:0] node42192;
	wire [4-1:0] node42193;
	wire [4-1:0] node42196;
	wire [4-1:0] node42197;
	wire [4-1:0] node42201;
	wire [4-1:0] node42202;
	wire [4-1:0] node42203;
	wire [4-1:0] node42207;
	wire [4-1:0] node42208;
	wire [4-1:0] node42211;
	wire [4-1:0] node42214;
	wire [4-1:0] node42215;
	wire [4-1:0] node42216;
	wire [4-1:0] node42217;
	wire [4-1:0] node42219;
	wire [4-1:0] node42222;
	wire [4-1:0] node42224;
	wire [4-1:0] node42227;
	wire [4-1:0] node42228;
	wire [4-1:0] node42231;
	wire [4-1:0] node42234;
	wire [4-1:0] node42235;
	wire [4-1:0] node42236;
	wire [4-1:0] node42237;
	wire [4-1:0] node42240;
	wire [4-1:0] node42243;
	wire [4-1:0] node42244;
	wire [4-1:0] node42247;
	wire [4-1:0] node42250;
	wire [4-1:0] node42251;
	wire [4-1:0] node42254;
	wire [4-1:0] node42257;
	wire [4-1:0] node42258;
	wire [4-1:0] node42259;
	wire [4-1:0] node42260;
	wire [4-1:0] node42261;
	wire [4-1:0] node42262;
	wire [4-1:0] node42266;
	wire [4-1:0] node42267;
	wire [4-1:0] node42271;
	wire [4-1:0] node42273;
	wire [4-1:0] node42276;
	wire [4-1:0] node42277;
	wire [4-1:0] node42278;
	wire [4-1:0] node42280;
	wire [4-1:0] node42283;
	wire [4-1:0] node42285;
	wire [4-1:0] node42288;
	wire [4-1:0] node42289;
	wire [4-1:0] node42291;
	wire [4-1:0] node42295;
	wire [4-1:0] node42296;
	wire [4-1:0] node42297;
	wire [4-1:0] node42298;
	wire [4-1:0] node42302;
	wire [4-1:0] node42303;
	wire [4-1:0] node42307;
	wire [4-1:0] node42308;
	wire [4-1:0] node42309;
	wire [4-1:0] node42313;
	wire [4-1:0] node42314;
	wire [4-1:0] node42318;
	wire [4-1:0] node42319;
	wire [4-1:0] node42320;
	wire [4-1:0] node42321;
	wire [4-1:0] node42322;
	wire [4-1:0] node42323;
	wire [4-1:0] node42324;
	wire [4-1:0] node42328;
	wire [4-1:0] node42329;
	wire [4-1:0] node42332;
	wire [4-1:0] node42335;
	wire [4-1:0] node42336;
	wire [4-1:0] node42339;
	wire [4-1:0] node42342;
	wire [4-1:0] node42343;
	wire [4-1:0] node42344;
	wire [4-1:0] node42347;
	wire [4-1:0] node42348;
	wire [4-1:0] node42352;
	wire [4-1:0] node42353;
	wire [4-1:0] node42356;
	wire [4-1:0] node42357;
	wire [4-1:0] node42361;
	wire [4-1:0] node42362;
	wire [4-1:0] node42363;
	wire [4-1:0] node42364;
	wire [4-1:0] node42366;
	wire [4-1:0] node42369;
	wire [4-1:0] node42370;
	wire [4-1:0] node42374;
	wire [4-1:0] node42375;
	wire [4-1:0] node42376;
	wire [4-1:0] node42380;
	wire [4-1:0] node42382;
	wire [4-1:0] node42385;
	wire [4-1:0] node42386;
	wire [4-1:0] node42387;
	wire [4-1:0] node42389;
	wire [4-1:0] node42392;
	wire [4-1:0] node42393;
	wire [4-1:0] node42397;
	wire [4-1:0] node42398;
	wire [4-1:0] node42400;
	wire [4-1:0] node42403;
	wire [4-1:0] node42404;
	wire [4-1:0] node42408;
	wire [4-1:0] node42409;
	wire [4-1:0] node42410;
	wire [4-1:0] node42411;
	wire [4-1:0] node42412;
	wire [4-1:0] node42416;
	wire [4-1:0] node42417;
	wire [4-1:0] node42418;
	wire [4-1:0] node42421;
	wire [4-1:0] node42424;
	wire [4-1:0] node42425;
	wire [4-1:0] node42428;
	wire [4-1:0] node42431;
	wire [4-1:0] node42432;
	wire [4-1:0] node42433;
	wire [4-1:0] node42434;
	wire [4-1:0] node42437;
	wire [4-1:0] node42440;
	wire [4-1:0] node42442;
	wire [4-1:0] node42445;
	wire [4-1:0] node42446;
	wire [4-1:0] node42448;
	wire [4-1:0] node42451;
	wire [4-1:0] node42452;
	wire [4-1:0] node42455;
	wire [4-1:0] node42458;
	wire [4-1:0] node42459;
	wire [4-1:0] node42460;
	wire [4-1:0] node42461;
	wire [4-1:0] node42465;
	wire [4-1:0] node42466;
	wire [4-1:0] node42470;
	wire [4-1:0] node42471;
	wire [4-1:0] node42472;
	wire [4-1:0] node42476;
	wire [4-1:0] node42477;
	wire [4-1:0] node42481;
	wire [4-1:0] node42482;
	wire [4-1:0] node42483;
	wire [4-1:0] node42484;
	wire [4-1:0] node42485;
	wire [4-1:0] node42486;
	wire [4-1:0] node42487;
	wire [4-1:0] node42488;
	wire [4-1:0] node42490;
	wire [4-1:0] node42493;
	wire [4-1:0] node42496;
	wire [4-1:0] node42497;
	wire [4-1:0] node42499;
	wire [4-1:0] node42502;
	wire [4-1:0] node42505;
	wire [4-1:0] node42506;
	wire [4-1:0] node42507;
	wire [4-1:0] node42508;
	wire [4-1:0] node42512;
	wire [4-1:0] node42513;
	wire [4-1:0] node42516;
	wire [4-1:0] node42519;
	wire [4-1:0] node42520;
	wire [4-1:0] node42521;
	wire [4-1:0] node42525;
	wire [4-1:0] node42526;
	wire [4-1:0] node42529;
	wire [4-1:0] node42532;
	wire [4-1:0] node42533;
	wire [4-1:0] node42534;
	wire [4-1:0] node42535;
	wire [4-1:0] node42536;
	wire [4-1:0] node42539;
	wire [4-1:0] node42542;
	wire [4-1:0] node42543;
	wire [4-1:0] node42546;
	wire [4-1:0] node42549;
	wire [4-1:0] node42550;
	wire [4-1:0] node42553;
	wire [4-1:0] node42554;
	wire [4-1:0] node42558;
	wire [4-1:0] node42559;
	wire [4-1:0] node42560;
	wire [4-1:0] node42562;
	wire [4-1:0] node42565;
	wire [4-1:0] node42566;
	wire [4-1:0] node42569;
	wire [4-1:0] node42572;
	wire [4-1:0] node42573;
	wire [4-1:0] node42575;
	wire [4-1:0] node42578;
	wire [4-1:0] node42579;
	wire [4-1:0] node42582;
	wire [4-1:0] node42585;
	wire [4-1:0] node42586;
	wire [4-1:0] node42587;
	wire [4-1:0] node42588;
	wire [4-1:0] node42589;
	wire [4-1:0] node42592;
	wire [4-1:0] node42594;
	wire [4-1:0] node42597;
	wire [4-1:0] node42598;
	wire [4-1:0] node42599;
	wire [4-1:0] node42603;
	wire [4-1:0] node42604;
	wire [4-1:0] node42607;
	wire [4-1:0] node42610;
	wire [4-1:0] node42611;
	wire [4-1:0] node42612;
	wire [4-1:0] node42615;
	wire [4-1:0] node42617;
	wire [4-1:0] node42620;
	wire [4-1:0] node42621;
	wire [4-1:0] node42622;
	wire [4-1:0] node42625;
	wire [4-1:0] node42629;
	wire [4-1:0] node42630;
	wire [4-1:0] node42631;
	wire [4-1:0] node42633;
	wire [4-1:0] node42634;
	wire [4-1:0] node42638;
	wire [4-1:0] node42639;
	wire [4-1:0] node42642;
	wire [4-1:0] node42645;
	wire [4-1:0] node42646;
	wire [4-1:0] node42647;
	wire [4-1:0] node42648;
	wire [4-1:0] node42651;
	wire [4-1:0] node42654;
	wire [4-1:0] node42656;
	wire [4-1:0] node42659;
	wire [4-1:0] node42660;
	wire [4-1:0] node42663;
	wire [4-1:0] node42666;
	wire [4-1:0] node42667;
	wire [4-1:0] node42668;
	wire [4-1:0] node42669;
	wire [4-1:0] node42670;
	wire [4-1:0] node42671;
	wire [4-1:0] node42672;
	wire [4-1:0] node42675;
	wire [4-1:0] node42678;
	wire [4-1:0] node42679;
	wire [4-1:0] node42682;
	wire [4-1:0] node42685;
	wire [4-1:0] node42686;
	wire [4-1:0] node42689;
	wire [4-1:0] node42691;
	wire [4-1:0] node42694;
	wire [4-1:0] node42695;
	wire [4-1:0] node42696;
	wire [4-1:0] node42697;
	wire [4-1:0] node42700;
	wire [4-1:0] node42703;
	wire [4-1:0] node42704;
	wire [4-1:0] node42708;
	wire [4-1:0] node42710;
	wire [4-1:0] node42711;
	wire [4-1:0] node42714;
	wire [4-1:0] node42717;
	wire [4-1:0] node42718;
	wire [4-1:0] node42719;
	wire [4-1:0] node42720;
	wire [4-1:0] node42722;
	wire [4-1:0] node42725;
	wire [4-1:0] node42727;
	wire [4-1:0] node42730;
	wire [4-1:0] node42731;
	wire [4-1:0] node42734;
	wire [4-1:0] node42736;
	wire [4-1:0] node42739;
	wire [4-1:0] node42740;
	wire [4-1:0] node42742;
	wire [4-1:0] node42743;
	wire [4-1:0] node42746;
	wire [4-1:0] node42749;
	wire [4-1:0] node42750;
	wire [4-1:0] node42751;
	wire [4-1:0] node42754;
	wire [4-1:0] node42757;
	wire [4-1:0] node42758;
	wire [4-1:0] node42762;
	wire [4-1:0] node42763;
	wire [4-1:0] node42764;
	wire [4-1:0] node42765;
	wire [4-1:0] node42766;
	wire [4-1:0] node42768;
	wire [4-1:0] node42771;
	wire [4-1:0] node42772;
	wire [4-1:0] node42775;
	wire [4-1:0] node42778;
	wire [4-1:0] node42779;
	wire [4-1:0] node42780;
	wire [4-1:0] node42783;
	wire [4-1:0] node42786;
	wire [4-1:0] node42787;
	wire [4-1:0] node42791;
	wire [4-1:0] node42792;
	wire [4-1:0] node42793;
	wire [4-1:0] node42794;
	wire [4-1:0] node42797;
	wire [4-1:0] node42800;
	wire [4-1:0] node42801;
	wire [4-1:0] node42804;
	wire [4-1:0] node42807;
	wire [4-1:0] node42808;
	wire [4-1:0] node42809;
	wire [4-1:0] node42812;
	wire [4-1:0] node42815;
	wire [4-1:0] node42816;
	wire [4-1:0] node42820;
	wire [4-1:0] node42821;
	wire [4-1:0] node42822;
	wire [4-1:0] node42823;
	wire [4-1:0] node42824;
	wire [4-1:0] node42827;
	wire [4-1:0] node42830;
	wire [4-1:0] node42832;
	wire [4-1:0] node42835;
	wire [4-1:0] node42836;
	wire [4-1:0] node42837;
	wire [4-1:0] node42840;
	wire [4-1:0] node42843;
	wire [4-1:0] node42845;
	wire [4-1:0] node42848;
	wire [4-1:0] node42849;
	wire [4-1:0] node42850;
	wire [4-1:0] node42851;
	wire [4-1:0] node42855;
	wire [4-1:0] node42856;
	wire [4-1:0] node42859;
	wire [4-1:0] node42862;
	wire [4-1:0] node42863;
	wire [4-1:0] node42864;
	wire [4-1:0] node42867;
	wire [4-1:0] node42870;
	wire [4-1:0] node42871;
	wire [4-1:0] node42875;
	wire [4-1:0] node42876;
	wire [4-1:0] node42877;
	wire [4-1:0] node42878;
	wire [4-1:0] node42879;
	wire [4-1:0] node42880;
	wire [4-1:0] node42881;
	wire [4-1:0] node42882;
	wire [4-1:0] node42885;
	wire [4-1:0] node42888;
	wire [4-1:0] node42889;
	wire [4-1:0] node42892;
	wire [4-1:0] node42895;
	wire [4-1:0] node42896;
	wire [4-1:0] node42900;
	wire [4-1:0] node42901;
	wire [4-1:0] node42902;
	wire [4-1:0] node42905;
	wire [4-1:0] node42908;
	wire [4-1:0] node42909;
	wire [4-1:0] node42912;
	wire [4-1:0] node42913;
	wire [4-1:0] node42916;
	wire [4-1:0] node42919;
	wire [4-1:0] node42920;
	wire [4-1:0] node42921;
	wire [4-1:0] node42922;
	wire [4-1:0] node42925;
	wire [4-1:0] node42927;
	wire [4-1:0] node42930;
	wire [4-1:0] node42931;
	wire [4-1:0] node42932;
	wire [4-1:0] node42935;
	wire [4-1:0] node42938;
	wire [4-1:0] node42939;
	wire [4-1:0] node42943;
	wire [4-1:0] node42944;
	wire [4-1:0] node42945;
	wire [4-1:0] node42948;
	wire [4-1:0] node42951;
	wire [4-1:0] node42952;
	wire [4-1:0] node42955;
	wire [4-1:0] node42958;
	wire [4-1:0] node42959;
	wire [4-1:0] node42960;
	wire [4-1:0] node42961;
	wire [4-1:0] node42962;
	wire [4-1:0] node42963;
	wire [4-1:0] node42967;
	wire [4-1:0] node42968;
	wire [4-1:0] node42972;
	wire [4-1:0] node42973;
	wire [4-1:0] node42974;
	wire [4-1:0] node42978;
	wire [4-1:0] node42979;
	wire [4-1:0] node42982;
	wire [4-1:0] node42985;
	wire [4-1:0] node42986;
	wire [4-1:0] node42987;
	wire [4-1:0] node42990;
	wire [4-1:0] node42993;
	wire [4-1:0] node42994;
	wire [4-1:0] node42997;
	wire [4-1:0] node43000;
	wire [4-1:0] node43001;
	wire [4-1:0] node43002;
	wire [4-1:0] node43003;
	wire [4-1:0] node43006;
	wire [4-1:0] node43008;
	wire [4-1:0] node43011;
	wire [4-1:0] node43012;
	wire [4-1:0] node43014;
	wire [4-1:0] node43017;
	wire [4-1:0] node43020;
	wire [4-1:0] node43021;
	wire [4-1:0] node43022;
	wire [4-1:0] node43026;
	wire [4-1:0] node43029;
	wire [4-1:0] node43030;
	wire [4-1:0] node43031;
	wire [4-1:0] node43032;
	wire [4-1:0] node43033;
	wire [4-1:0] node43034;
	wire [4-1:0] node43035;
	wire [4-1:0] node43038;
	wire [4-1:0] node43041;
	wire [4-1:0] node43042;
	wire [4-1:0] node43046;
	wire [4-1:0] node43047;
	wire [4-1:0] node43050;
	wire [4-1:0] node43053;
	wire [4-1:0] node43054;
	wire [4-1:0] node43055;
	wire [4-1:0] node43056;
	wire [4-1:0] node43059;
	wire [4-1:0] node43062;
	wire [4-1:0] node43063;
	wire [4-1:0] node43066;
	wire [4-1:0] node43069;
	wire [4-1:0] node43070;
	wire [4-1:0] node43073;
	wire [4-1:0] node43076;
	wire [4-1:0] node43077;
	wire [4-1:0] node43078;
	wire [4-1:0] node43079;
	wire [4-1:0] node43081;
	wire [4-1:0] node43085;
	wire [4-1:0] node43086;
	wire [4-1:0] node43090;
	wire [4-1:0] node43091;
	wire [4-1:0] node43092;
	wire [4-1:0] node43094;
	wire [4-1:0] node43097;
	wire [4-1:0] node43098;
	wire [4-1:0] node43102;
	wire [4-1:0] node43105;
	wire [4-1:0] node43106;
	wire [4-1:0] node43107;
	wire [4-1:0] node43108;
	wire [4-1:0] node43109;
	wire [4-1:0] node43110;
	wire [4-1:0] node43113;
	wire [4-1:0] node43116;
	wire [4-1:0] node43117;
	wire [4-1:0] node43121;
	wire [4-1:0] node43122;
	wire [4-1:0] node43123;
	wire [4-1:0] node43126;
	wire [4-1:0] node43129;
	wire [4-1:0] node43130;
	wire [4-1:0] node43133;
	wire [4-1:0] node43136;
	wire [4-1:0] node43137;
	wire [4-1:0] node43138;
	wire [4-1:0] node43139;
	wire [4-1:0] node43142;
	wire [4-1:0] node43145;
	wire [4-1:0] node43146;
	wire [4-1:0] node43149;
	wire [4-1:0] node43152;
	wire [4-1:0] node43153;
	wire [4-1:0] node43154;
	wire [4-1:0] node43158;
	wire [4-1:0] node43159;
	wire [4-1:0] node43163;
	wire [4-1:0] node43164;
	wire [4-1:0] node43165;
	wire [4-1:0] node43166;
	wire [4-1:0] node43168;
	wire [4-1:0] node43172;
	wire [4-1:0] node43173;
	wire [4-1:0] node43174;
	wire [4-1:0] node43177;
	wire [4-1:0] node43180;
	wire [4-1:0] node43181;
	wire [4-1:0] node43184;
	wire [4-1:0] node43187;
	wire [4-1:0] node43188;
	wire [4-1:0] node43190;
	wire [4-1:0] node43193;
	wire [4-1:0] node43194;
	wire [4-1:0] node43195;
	wire [4-1:0] node43198;
	wire [4-1:0] node43201;
	wire [4-1:0] node43202;
	wire [4-1:0] node43205;
	wire [4-1:0] node43208;
	wire [4-1:0] node43209;
	wire [4-1:0] node43210;
	wire [4-1:0] node43211;
	wire [4-1:0] node43212;
	wire [4-1:0] node43213;
	wire [4-1:0] node43214;
	wire [4-1:0] node43215;
	wire [4-1:0] node43216;
	wire [4-1:0] node43217;
	wire [4-1:0] node43221;
	wire [4-1:0] node43222;
	wire [4-1:0] node43225;
	wire [4-1:0] node43228;
	wire [4-1:0] node43229;
	wire [4-1:0] node43230;
	wire [4-1:0] node43233;
	wire [4-1:0] node43236;
	wire [4-1:0] node43237;
	wire [4-1:0] node43240;
	wire [4-1:0] node43243;
	wire [4-1:0] node43244;
	wire [4-1:0] node43245;
	wire [4-1:0] node43246;
	wire [4-1:0] node43249;
	wire [4-1:0] node43252;
	wire [4-1:0] node43253;
	wire [4-1:0] node43256;
	wire [4-1:0] node43259;
	wire [4-1:0] node43260;
	wire [4-1:0] node43261;
	wire [4-1:0] node43264;
	wire [4-1:0] node43267;
	wire [4-1:0] node43268;
	wire [4-1:0] node43271;
	wire [4-1:0] node43274;
	wire [4-1:0] node43275;
	wire [4-1:0] node43276;
	wire [4-1:0] node43277;
	wire [4-1:0] node43279;
	wire [4-1:0] node43282;
	wire [4-1:0] node43283;
	wire [4-1:0] node43286;
	wire [4-1:0] node43289;
	wire [4-1:0] node43290;
	wire [4-1:0] node43291;
	wire [4-1:0] node43296;
	wire [4-1:0] node43297;
	wire [4-1:0] node43298;
	wire [4-1:0] node43299;
	wire [4-1:0] node43302;
	wire [4-1:0] node43305;
	wire [4-1:0] node43306;
	wire [4-1:0] node43309;
	wire [4-1:0] node43312;
	wire [4-1:0] node43313;
	wire [4-1:0] node43314;
	wire [4-1:0] node43317;
	wire [4-1:0] node43320;
	wire [4-1:0] node43323;
	wire [4-1:0] node43324;
	wire [4-1:0] node43325;
	wire [4-1:0] node43326;
	wire [4-1:0] node43327;
	wire [4-1:0] node43328;
	wire [4-1:0] node43332;
	wire [4-1:0] node43333;
	wire [4-1:0] node43337;
	wire [4-1:0] node43338;
	wire [4-1:0] node43339;
	wire [4-1:0] node43344;
	wire [4-1:0] node43345;
	wire [4-1:0] node43346;
	wire [4-1:0] node43347;
	wire [4-1:0] node43351;
	wire [4-1:0] node43354;
	wire [4-1:0] node43355;
	wire [4-1:0] node43357;
	wire [4-1:0] node43360;
	wire [4-1:0] node43362;
	wire [4-1:0] node43365;
	wire [4-1:0] node43366;
	wire [4-1:0] node43367;
	wire [4-1:0] node43368;
	wire [4-1:0] node43369;
	wire [4-1:0] node43372;
	wire [4-1:0] node43375;
	wire [4-1:0] node43376;
	wire [4-1:0] node43379;
	wire [4-1:0] node43382;
	wire [4-1:0] node43383;
	wire [4-1:0] node43385;
	wire [4-1:0] node43388;
	wire [4-1:0] node43389;
	wire [4-1:0] node43393;
	wire [4-1:0] node43394;
	wire [4-1:0] node43395;
	wire [4-1:0] node43398;
	wire [4-1:0] node43400;
	wire [4-1:0] node43403;
	wire [4-1:0] node43404;
	wire [4-1:0] node43407;
	wire [4-1:0] node43409;
	wire [4-1:0] node43412;
	wire [4-1:0] node43413;
	wire [4-1:0] node43414;
	wire [4-1:0] node43415;
	wire [4-1:0] node43416;
	wire [4-1:0] node43417;
	wire [4-1:0] node43418;
	wire [4-1:0] node43421;
	wire [4-1:0] node43424;
	wire [4-1:0] node43425;
	wire [4-1:0] node43428;
	wire [4-1:0] node43431;
	wire [4-1:0] node43433;
	wire [4-1:0] node43435;
	wire [4-1:0] node43438;
	wire [4-1:0] node43439;
	wire [4-1:0] node43440;
	wire [4-1:0] node43442;
	wire [4-1:0] node43445;
	wire [4-1:0] node43446;
	wire [4-1:0] node43449;
	wire [4-1:0] node43452;
	wire [4-1:0] node43453;
	wire [4-1:0] node43456;
	wire [4-1:0] node43457;
	wire [4-1:0] node43461;
	wire [4-1:0] node43462;
	wire [4-1:0] node43463;
	wire [4-1:0] node43464;
	wire [4-1:0] node43465;
	wire [4-1:0] node43469;
	wire [4-1:0] node43470;
	wire [4-1:0] node43474;
	wire [4-1:0] node43475;
	wire [4-1:0] node43476;
	wire [4-1:0] node43479;
	wire [4-1:0] node43482;
	wire [4-1:0] node43483;
	wire [4-1:0] node43486;
	wire [4-1:0] node43489;
	wire [4-1:0] node43490;
	wire [4-1:0] node43491;
	wire [4-1:0] node43493;
	wire [4-1:0] node43496;
	wire [4-1:0] node43497;
	wire [4-1:0] node43500;
	wire [4-1:0] node43503;
	wire [4-1:0] node43504;
	wire [4-1:0] node43508;
	wire [4-1:0] node43509;
	wire [4-1:0] node43510;
	wire [4-1:0] node43511;
	wire [4-1:0] node43512;
	wire [4-1:0] node43514;
	wire [4-1:0] node43517;
	wire [4-1:0] node43519;
	wire [4-1:0] node43522;
	wire [4-1:0] node43523;
	wire [4-1:0] node43524;
	wire [4-1:0] node43528;
	wire [4-1:0] node43529;
	wire [4-1:0] node43532;
	wire [4-1:0] node43535;
	wire [4-1:0] node43536;
	wire [4-1:0] node43537;
	wire [4-1:0] node43539;
	wire [4-1:0] node43542;
	wire [4-1:0] node43545;
	wire [4-1:0] node43546;
	wire [4-1:0] node43548;
	wire [4-1:0] node43552;
	wire [4-1:0] node43553;
	wire [4-1:0] node43554;
	wire [4-1:0] node43556;
	wire [4-1:0] node43557;
	wire [4-1:0] node43560;
	wire [4-1:0] node43563;
	wire [4-1:0] node43564;
	wire [4-1:0] node43565;
	wire [4-1:0] node43568;
	wire [4-1:0] node43571;
	wire [4-1:0] node43574;
	wire [4-1:0] node43575;
	wire [4-1:0] node43576;
	wire [4-1:0] node43577;
	wire [4-1:0] node43580;
	wire [4-1:0] node43583;
	wire [4-1:0] node43584;
	wire [4-1:0] node43587;
	wire [4-1:0] node43590;
	wire [4-1:0] node43591;
	wire [4-1:0] node43593;
	wire [4-1:0] node43597;
	wire [4-1:0] node43598;
	wire [4-1:0] node43599;
	wire [4-1:0] node43600;
	wire [4-1:0] node43601;
	wire [4-1:0] node43602;
	wire [4-1:0] node43603;
	wire [4-1:0] node43604;
	wire [4-1:0] node43607;
	wire [4-1:0] node43611;
	wire [4-1:0] node43612;
	wire [4-1:0] node43613;
	wire [4-1:0] node43616;
	wire [4-1:0] node43619;
	wire [4-1:0] node43621;
	wire [4-1:0] node43624;
	wire [4-1:0] node43625;
	wire [4-1:0] node43626;
	wire [4-1:0] node43629;
	wire [4-1:0] node43632;
	wire [4-1:0] node43633;
	wire [4-1:0] node43636;
	wire [4-1:0] node43639;
	wire [4-1:0] node43640;
	wire [4-1:0] node43641;
	wire [4-1:0] node43642;
	wire [4-1:0] node43643;
	wire [4-1:0] node43646;
	wire [4-1:0] node43649;
	wire [4-1:0] node43650;
	wire [4-1:0] node43653;
	wire [4-1:0] node43656;
	wire [4-1:0] node43657;
	wire [4-1:0] node43661;
	wire [4-1:0] node43662;
	wire [4-1:0] node43663;
	wire [4-1:0] node43664;
	wire [4-1:0] node43668;
	wire [4-1:0] node43669;
	wire [4-1:0] node43672;
	wire [4-1:0] node43675;
	wire [4-1:0] node43678;
	wire [4-1:0] node43679;
	wire [4-1:0] node43680;
	wire [4-1:0] node43681;
	wire [4-1:0] node43682;
	wire [4-1:0] node43683;
	wire [4-1:0] node43686;
	wire [4-1:0] node43689;
	wire [4-1:0] node43690;
	wire [4-1:0] node43693;
	wire [4-1:0] node43696;
	wire [4-1:0] node43697;
	wire [4-1:0] node43700;
	wire [4-1:0] node43702;
	wire [4-1:0] node43705;
	wire [4-1:0] node43706;
	wire [4-1:0] node43707;
	wire [4-1:0] node43711;
	wire [4-1:0] node43712;
	wire [4-1:0] node43713;
	wire [4-1:0] node43716;
	wire [4-1:0] node43719;
	wire [4-1:0] node43720;
	wire [4-1:0] node43723;
	wire [4-1:0] node43726;
	wire [4-1:0] node43727;
	wire [4-1:0] node43728;
	wire [4-1:0] node43730;
	wire [4-1:0] node43733;
	wire [4-1:0] node43734;
	wire [4-1:0] node43738;
	wire [4-1:0] node43739;
	wire [4-1:0] node43740;
	wire [4-1:0] node43744;
	wire [4-1:0] node43745;
	wire [4-1:0] node43749;
	wire [4-1:0] node43750;
	wire [4-1:0] node43751;
	wire [4-1:0] node43752;
	wire [4-1:0] node43753;
	wire [4-1:0] node43754;
	wire [4-1:0] node43755;
	wire [4-1:0] node43758;
	wire [4-1:0] node43762;
	wire [4-1:0] node43763;
	wire [4-1:0] node43764;
	wire [4-1:0] node43768;
	wire [4-1:0] node43771;
	wire [4-1:0] node43772;
	wire [4-1:0] node43773;
	wire [4-1:0] node43776;
	wire [4-1:0] node43779;
	wire [4-1:0] node43780;
	wire [4-1:0] node43783;
	wire [4-1:0] node43786;
	wire [4-1:0] node43787;
	wire [4-1:0] node43788;
	wire [4-1:0] node43789;
	wire [4-1:0] node43792;
	wire [4-1:0] node43794;
	wire [4-1:0] node43797;
	wire [4-1:0] node43798;
	wire [4-1:0] node43802;
	wire [4-1:0] node43803;
	wire [4-1:0] node43804;
	wire [4-1:0] node43805;
	wire [4-1:0] node43809;
	wire [4-1:0] node43810;
	wire [4-1:0] node43814;
	wire [4-1:0] node43817;
	wire [4-1:0] node43818;
	wire [4-1:0] node43819;
	wire [4-1:0] node43820;
	wire [4-1:0] node43822;
	wire [4-1:0] node43823;
	wire [4-1:0] node43827;
	wire [4-1:0] node43829;
	wire [4-1:0] node43832;
	wire [4-1:0] node43833;
	wire [4-1:0] node43834;
	wire [4-1:0] node43837;
	wire [4-1:0] node43839;
	wire [4-1:0] node43842;
	wire [4-1:0] node43845;
	wire [4-1:0] node43846;
	wire [4-1:0] node43847;
	wire [4-1:0] node43848;
	wire [4-1:0] node43849;
	wire [4-1:0] node43854;
	wire [4-1:0] node43855;
	wire [4-1:0] node43859;
	wire [4-1:0] node43860;
	wire [4-1:0] node43861;
	wire [4-1:0] node43863;
	wire [4-1:0] node43866;
	wire [4-1:0] node43869;
	wire [4-1:0] node43870;
	wire [4-1:0] node43874;
	wire [4-1:0] node43875;
	wire [4-1:0] node43876;
	wire [4-1:0] node43877;
	wire [4-1:0] node43878;
	wire [4-1:0] node43879;
	wire [4-1:0] node43880;
	wire [4-1:0] node43881;
	wire [4-1:0] node43883;
	wire [4-1:0] node43887;
	wire [4-1:0] node43888;
	wire [4-1:0] node43891;
	wire [4-1:0] node43892;
	wire [4-1:0] node43896;
	wire [4-1:0] node43897;
	wire [4-1:0] node43898;
	wire [4-1:0] node43899;
	wire [4-1:0] node43903;
	wire [4-1:0] node43904;
	wire [4-1:0] node43908;
	wire [4-1:0] node43909;
	wire [4-1:0] node43912;
	wire [4-1:0] node43913;
	wire [4-1:0] node43917;
	wire [4-1:0] node43918;
	wire [4-1:0] node43919;
	wire [4-1:0] node43920;
	wire [4-1:0] node43921;
	wire [4-1:0] node43925;
	wire [4-1:0] node43926;
	wire [4-1:0] node43929;
	wire [4-1:0] node43932;
	wire [4-1:0] node43933;
	wire [4-1:0] node43935;
	wire [4-1:0] node43938;
	wire [4-1:0] node43939;
	wire [4-1:0] node43942;
	wire [4-1:0] node43945;
	wire [4-1:0] node43946;
	wire [4-1:0] node43947;
	wire [4-1:0] node43950;
	wire [4-1:0] node43953;
	wire [4-1:0] node43956;
	wire [4-1:0] node43957;
	wire [4-1:0] node43958;
	wire [4-1:0] node43959;
	wire [4-1:0] node43960;
	wire [4-1:0] node43961;
	wire [4-1:0] node43965;
	wire [4-1:0] node43967;
	wire [4-1:0] node43970;
	wire [4-1:0] node43971;
	wire [4-1:0] node43972;
	wire [4-1:0] node43975;
	wire [4-1:0] node43978;
	wire [4-1:0] node43980;
	wire [4-1:0] node43983;
	wire [4-1:0] node43984;
	wire [4-1:0] node43985;
	wire [4-1:0] node43988;
	wire [4-1:0] node43991;
	wire [4-1:0] node43994;
	wire [4-1:0] node43995;
	wire [4-1:0] node43996;
	wire [4-1:0] node43997;
	wire [4-1:0] node43998;
	wire [4-1:0] node44001;
	wire [4-1:0] node44004;
	wire [4-1:0] node44007;
	wire [4-1:0] node44008;
	wire [4-1:0] node44009;
	wire [4-1:0] node44013;
	wire [4-1:0] node44014;
	wire [4-1:0] node44018;
	wire [4-1:0] node44019;
	wire [4-1:0] node44020;
	wire [4-1:0] node44023;
	wire [4-1:0] node44024;
	wire [4-1:0] node44028;
	wire [4-1:0] node44029;
	wire [4-1:0] node44032;
	wire [4-1:0] node44033;
	wire [4-1:0] node44037;
	wire [4-1:0] node44038;
	wire [4-1:0] node44039;
	wire [4-1:0] node44040;
	wire [4-1:0] node44041;
	wire [4-1:0] node44042;
	wire [4-1:0] node44043;
	wire [4-1:0] node44046;
	wire [4-1:0] node44049;
	wire [4-1:0] node44052;
	wire [4-1:0] node44053;
	wire [4-1:0] node44054;
	wire [4-1:0] node44059;
	wire [4-1:0] node44060;
	wire [4-1:0] node44061;
	wire [4-1:0] node44062;
	wire [4-1:0] node44067;
	wire [4-1:0] node44068;
	wire [4-1:0] node44070;
	wire [4-1:0] node44073;
	wire [4-1:0] node44074;
	wire [4-1:0] node44077;
	wire [4-1:0] node44080;
	wire [4-1:0] node44081;
	wire [4-1:0] node44082;
	wire [4-1:0] node44083;
	wire [4-1:0] node44084;
	wire [4-1:0] node44088;
	wire [4-1:0] node44090;
	wire [4-1:0] node44093;
	wire [4-1:0] node44094;
	wire [4-1:0] node44095;
	wire [4-1:0] node44098;
	wire [4-1:0] node44101;
	wire [4-1:0] node44103;
	wire [4-1:0] node44106;
	wire [4-1:0] node44107;
	wire [4-1:0] node44108;
	wire [4-1:0] node44111;
	wire [4-1:0] node44114;
	wire [4-1:0] node44117;
	wire [4-1:0] node44118;
	wire [4-1:0] node44119;
	wire [4-1:0] node44120;
	wire [4-1:0] node44121;
	wire [4-1:0] node44124;
	wire [4-1:0] node44125;
	wire [4-1:0] node44128;
	wire [4-1:0] node44131;
	wire [4-1:0] node44132;
	wire [4-1:0] node44133;
	wire [4-1:0] node44137;
	wire [4-1:0] node44139;
	wire [4-1:0] node44142;
	wire [4-1:0] node44143;
	wire [4-1:0] node44144;
	wire [4-1:0] node44147;
	wire [4-1:0] node44150;
	wire [4-1:0] node44153;
	wire [4-1:0] node44154;
	wire [4-1:0] node44155;
	wire [4-1:0] node44156;
	wire [4-1:0] node44157;
	wire [4-1:0] node44160;
	wire [4-1:0] node44163;
	wire [4-1:0] node44166;
	wire [4-1:0] node44167;
	wire [4-1:0] node44168;
	wire [4-1:0] node44172;
	wire [4-1:0] node44173;
	wire [4-1:0] node44177;
	wire [4-1:0] node44178;
	wire [4-1:0] node44179;
	wire [4-1:0] node44180;
	wire [4-1:0] node44183;
	wire [4-1:0] node44186;
	wire [4-1:0] node44187;
	wire [4-1:0] node44191;
	wire [4-1:0] node44192;
	wire [4-1:0] node44193;
	wire [4-1:0] node44196;
	wire [4-1:0] node44199;
	wire [4-1:0] node44200;
	wire [4-1:0] node44203;
	wire [4-1:0] node44206;
	wire [4-1:0] node44207;
	wire [4-1:0] node44208;
	wire [4-1:0] node44209;
	wire [4-1:0] node44210;
	wire [4-1:0] node44211;
	wire [4-1:0] node44212;
	wire [4-1:0] node44213;
	wire [4-1:0] node44216;
	wire [4-1:0] node44219;
	wire [4-1:0] node44222;
	wire [4-1:0] node44223;
	wire [4-1:0] node44224;
	wire [4-1:0] node44228;
	wire [4-1:0] node44231;
	wire [4-1:0] node44232;
	wire [4-1:0] node44233;
	wire [4-1:0] node44234;
	wire [4-1:0] node44238;
	wire [4-1:0] node44239;
	wire [4-1:0] node44243;
	wire [4-1:0] node44244;
	wire [4-1:0] node44245;
	wire [4-1:0] node44249;
	wire [4-1:0] node44252;
	wire [4-1:0] node44253;
	wire [4-1:0] node44254;
	wire [4-1:0] node44255;
	wire [4-1:0] node44256;
	wire [4-1:0] node44260;
	wire [4-1:0] node44261;
	wire [4-1:0] node44264;
	wire [4-1:0] node44267;
	wire [4-1:0] node44268;
	wire [4-1:0] node44269;
	wire [4-1:0] node44272;
	wire [4-1:0] node44275;
	wire [4-1:0] node44276;
	wire [4-1:0] node44279;
	wire [4-1:0] node44282;
	wire [4-1:0] node44283;
	wire [4-1:0] node44284;
	wire [4-1:0] node44287;
	wire [4-1:0] node44290;
	wire [4-1:0] node44293;
	wire [4-1:0] node44294;
	wire [4-1:0] node44295;
	wire [4-1:0] node44296;
	wire [4-1:0] node44297;
	wire [4-1:0] node44298;
	wire [4-1:0] node44302;
	wire [4-1:0] node44304;
	wire [4-1:0] node44307;
	wire [4-1:0] node44308;
	wire [4-1:0] node44309;
	wire [4-1:0] node44312;
	wire [4-1:0] node44315;
	wire [4-1:0] node44316;
	wire [4-1:0] node44319;
	wire [4-1:0] node44322;
	wire [4-1:0] node44323;
	wire [4-1:0] node44324;
	wire [4-1:0] node44327;
	wire [4-1:0] node44330;
	wire [4-1:0] node44333;
	wire [4-1:0] node44334;
	wire [4-1:0] node44335;
	wire [4-1:0] node44336;
	wire [4-1:0] node44339;
	wire [4-1:0] node44340;
	wire [4-1:0] node44345;
	wire [4-1:0] node44346;
	wire [4-1:0] node44349;
	wire [4-1:0] node44350;
	wire [4-1:0] node44354;
	wire [4-1:0] node44355;
	wire [4-1:0] node44356;
	wire [4-1:0] node44357;
	wire [4-1:0] node44358;
	wire [4-1:0] node44359;
	wire [4-1:0] node44360;
	wire [4-1:0] node44363;
	wire [4-1:0] node44366;
	wire [4-1:0] node44369;
	wire [4-1:0] node44370;
	wire [4-1:0] node44373;
	wire [4-1:0] node44374;
	wire [4-1:0] node44378;
	wire [4-1:0] node44379;
	wire [4-1:0] node44381;
	wire [4-1:0] node44382;
	wire [4-1:0] node44385;
	wire [4-1:0] node44388;
	wire [4-1:0] node44389;
	wire [4-1:0] node44390;
	wire [4-1:0] node44393;
	wire [4-1:0] node44397;
	wire [4-1:0] node44398;
	wire [4-1:0] node44399;
	wire [4-1:0] node44400;
	wire [4-1:0] node44401;
	wire [4-1:0] node44404;
	wire [4-1:0] node44407;
	wire [4-1:0] node44408;
	wire [4-1:0] node44411;
	wire [4-1:0] node44414;
	wire [4-1:0] node44415;
	wire [4-1:0] node44416;
	wire [4-1:0] node44419;
	wire [4-1:0] node44422;
	wire [4-1:0] node44424;
	wire [4-1:0] node44427;
	wire [4-1:0] node44428;
	wire [4-1:0] node44429;
	wire [4-1:0] node44432;
	wire [4-1:0] node44435;
	wire [4-1:0] node44438;
	wire [4-1:0] node44439;
	wire [4-1:0] node44440;
	wire [4-1:0] node44441;
	wire [4-1:0] node44442;
	wire [4-1:0] node44443;
	wire [4-1:0] node44446;
	wire [4-1:0] node44449;
	wire [4-1:0] node44451;
	wire [4-1:0] node44454;
	wire [4-1:0] node44455;
	wire [4-1:0] node44458;
	wire [4-1:0] node44459;
	wire [4-1:0] node44462;
	wire [4-1:0] node44465;
	wire [4-1:0] node44466;
	wire [4-1:0] node44467;
	wire [4-1:0] node44470;
	wire [4-1:0] node44473;
	wire [4-1:0] node44476;
	wire [4-1:0] node44477;
	wire [4-1:0] node44478;
	wire [4-1:0] node44479;
	wire [4-1:0] node44480;
	wire [4-1:0] node44484;
	wire [4-1:0] node44487;
	wire [4-1:0] node44489;
	wire [4-1:0] node44490;
	wire [4-1:0] node44494;
	wire [4-1:0] node44495;
	wire [4-1:0] node44496;
	wire [4-1:0] node44497;
	wire [4-1:0] node44500;
	wire [4-1:0] node44503;
	wire [4-1:0] node44504;
	wire [4-1:0] node44507;
	wire [4-1:0] node44510;
	wire [4-1:0] node44511;
	wire [4-1:0] node44512;
	wire [4-1:0] node44515;
	wire [4-1:0] node44518;
	wire [4-1:0] node44520;
	wire [4-1:0] node44523;
	wire [4-1:0] node44524;
	wire [4-1:0] node44525;
	wire [4-1:0] node44526;
	wire [4-1:0] node44527;
	wire [4-1:0] node44528;
	wire [4-1:0] node44529;
	wire [4-1:0] node44530;
	wire [4-1:0] node44531;
	wire [4-1:0] node44532;
	wire [4-1:0] node44533;
	wire [4-1:0] node44536;
	wire [4-1:0] node44539;
	wire [4-1:0] node44540;
	wire [4-1:0] node44543;
	wire [4-1:0] node44546;
	wire [4-1:0] node44547;
	wire [4-1:0] node44548;
	wire [4-1:0] node44551;
	wire [4-1:0] node44554;
	wire [4-1:0] node44555;
	wire [4-1:0] node44559;
	wire [4-1:0] node44560;
	wire [4-1:0] node44561;
	wire [4-1:0] node44562;
	wire [4-1:0] node44565;
	wire [4-1:0] node44568;
	wire [4-1:0] node44569;
	wire [4-1:0] node44572;
	wire [4-1:0] node44575;
	wire [4-1:0] node44576;
	wire [4-1:0] node44577;
	wire [4-1:0] node44580;
	wire [4-1:0] node44584;
	wire [4-1:0] node44585;
	wire [4-1:0] node44588;
	wire [4-1:0] node44591;
	wire [4-1:0] node44592;
	wire [4-1:0] node44593;
	wire [4-1:0] node44594;
	wire [4-1:0] node44595;
	wire [4-1:0] node44597;
	wire [4-1:0] node44600;
	wire [4-1:0] node44601;
	wire [4-1:0] node44605;
	wire [4-1:0] node44606;
	wire [4-1:0] node44608;
	wire [4-1:0] node44612;
	wire [4-1:0] node44613;
	wire [4-1:0] node44614;
	wire [4-1:0] node44616;
	wire [4-1:0] node44619;
	wire [4-1:0] node44621;
	wire [4-1:0] node44624;
	wire [4-1:0] node44625;
	wire [4-1:0] node44627;
	wire [4-1:0] node44630;
	wire [4-1:0] node44632;
	wire [4-1:0] node44635;
	wire [4-1:0] node44636;
	wire [4-1:0] node44637;
	wire [4-1:0] node44640;
	wire [4-1:0] node44643;
	wire [4-1:0] node44644;
	wire [4-1:0] node44645;
	wire [4-1:0] node44648;
	wire [4-1:0] node44651;
	wire [4-1:0] node44653;
	wire [4-1:0] node44654;
	wire [4-1:0] node44657;
	wire [4-1:0] node44660;
	wire [4-1:0] node44661;
	wire [4-1:0] node44662;
	wire [4-1:0] node44663;
	wire [4-1:0] node44664;
	wire [4-1:0] node44666;
	wire [4-1:0] node44669;
	wire [4-1:0] node44670;
	wire [4-1:0] node44671;
	wire [4-1:0] node44674;
	wire [4-1:0] node44677;
	wire [4-1:0] node44679;
	wire [4-1:0] node44682;
	wire [4-1:0] node44683;
	wire [4-1:0] node44686;
	wire [4-1:0] node44689;
	wire [4-1:0] node44690;
	wire [4-1:0] node44691;
	wire [4-1:0] node44693;
	wire [4-1:0] node44696;
	wire [4-1:0] node44698;
	wire [4-1:0] node44699;
	wire [4-1:0] node44702;
	wire [4-1:0] node44705;
	wire [4-1:0] node44706;
	wire [4-1:0] node44707;
	wire [4-1:0] node44708;
	wire [4-1:0] node44711;
	wire [4-1:0] node44714;
	wire [4-1:0] node44715;
	wire [4-1:0] node44718;
	wire [4-1:0] node44721;
	wire [4-1:0] node44722;
	wire [4-1:0] node44723;
	wire [4-1:0] node44727;
	wire [4-1:0] node44728;
	wire [4-1:0] node44731;
	wire [4-1:0] node44734;
	wire [4-1:0] node44735;
	wire [4-1:0] node44736;
	wire [4-1:0] node44738;
	wire [4-1:0] node44741;
	wire [4-1:0] node44743;
	wire [4-1:0] node44746;
	wire [4-1:0] node44747;
	wire [4-1:0] node44749;
	wire [4-1:0] node44752;
	wire [4-1:0] node44754;
	wire [4-1:0] node44757;
	wire [4-1:0] node44758;
	wire [4-1:0] node44759;
	wire [4-1:0] node44760;
	wire [4-1:0] node44761;
	wire [4-1:0] node44762;
	wire [4-1:0] node44766;
	wire [4-1:0] node44767;
	wire [4-1:0] node44771;
	wire [4-1:0] node44772;
	wire [4-1:0] node44773;
	wire [4-1:0] node44777;
	wire [4-1:0] node44778;
	wire [4-1:0] node44782;
	wire [4-1:0] node44783;
	wire [4-1:0] node44784;
	wire [4-1:0] node44785;
	wire [4-1:0] node44786;
	wire [4-1:0] node44787;
	wire [4-1:0] node44790;
	wire [4-1:0] node44793;
	wire [4-1:0] node44795;
	wire [4-1:0] node44798;
	wire [4-1:0] node44799;
	wire [4-1:0] node44800;
	wire [4-1:0] node44803;
	wire [4-1:0] node44806;
	wire [4-1:0] node44808;
	wire [4-1:0] node44811;
	wire [4-1:0] node44812;
	wire [4-1:0] node44813;
	wire [4-1:0] node44814;
	wire [4-1:0] node44817;
	wire [4-1:0] node44821;
	wire [4-1:0] node44822;
	wire [4-1:0] node44823;
	wire [4-1:0] node44826;
	wire [4-1:0] node44829;
	wire [4-1:0] node44830;
	wire [4-1:0] node44834;
	wire [4-1:0] node44835;
	wire [4-1:0] node44836;
	wire [4-1:0] node44839;
	wire [4-1:0] node44842;
	wire [4-1:0] node44843;
	wire [4-1:0] node44844;
	wire [4-1:0] node44845;
	wire [4-1:0] node44848;
	wire [4-1:0] node44851;
	wire [4-1:0] node44853;
	wire [4-1:0] node44856;
	wire [4-1:0] node44857;
	wire [4-1:0] node44860;
	wire [4-1:0] node44863;
	wire [4-1:0] node44864;
	wire [4-1:0] node44865;
	wire [4-1:0] node44866;
	wire [4-1:0] node44867;
	wire [4-1:0] node44868;
	wire [4-1:0] node44869;
	wire [4-1:0] node44872;
	wire [4-1:0] node44875;
	wire [4-1:0] node44876;
	wire [4-1:0] node44879;
	wire [4-1:0] node44882;
	wire [4-1:0] node44883;
	wire [4-1:0] node44884;
	wire [4-1:0] node44887;
	wire [4-1:0] node44890;
	wire [4-1:0] node44891;
	wire [4-1:0] node44894;
	wire [4-1:0] node44897;
	wire [4-1:0] node44898;
	wire [4-1:0] node44899;
	wire [4-1:0] node44902;
	wire [4-1:0] node44905;
	wire [4-1:0] node44906;
	wire [4-1:0] node44909;
	wire [4-1:0] node44912;
	wire [4-1:0] node44913;
	wire [4-1:0] node44914;
	wire [4-1:0] node44915;
	wire [4-1:0] node44918;
	wire [4-1:0] node44921;
	wire [4-1:0] node44922;
	wire [4-1:0] node44925;
	wire [4-1:0] node44928;
	wire [4-1:0] node44929;
	wire [4-1:0] node44930;
	wire [4-1:0] node44933;
	wire [4-1:0] node44936;
	wire [4-1:0] node44937;
	wire [4-1:0] node44939;
	wire [4-1:0] node44943;
	wire [4-1:0] node44944;
	wire [4-1:0] node44945;
	wire [4-1:0] node44946;
	wire [4-1:0] node44947;
	wire [4-1:0] node44948;
	wire [4-1:0] node44952;
	wire [4-1:0] node44954;
	wire [4-1:0] node44957;
	wire [4-1:0] node44958;
	wire [4-1:0] node44961;
	wire [4-1:0] node44964;
	wire [4-1:0] node44965;
	wire [4-1:0] node44968;
	wire [4-1:0] node44971;
	wire [4-1:0] node44972;
	wire [4-1:0] node44973;
	wire [4-1:0] node44974;
	wire [4-1:0] node44975;
	wire [4-1:0] node44979;
	wire [4-1:0] node44980;
	wire [4-1:0] node44983;
	wire [4-1:0] node44986;
	wire [4-1:0] node44988;
	wire [4-1:0] node44989;
	wire [4-1:0] node44992;
	wire [4-1:0] node44995;
	wire [4-1:0] node44996;
	wire [4-1:0] node44997;
	wire [4-1:0] node44998;
	wire [4-1:0] node45001;
	wire [4-1:0] node45004;
	wire [4-1:0] node45005;
	wire [4-1:0] node45008;
	wire [4-1:0] node45011;
	wire [4-1:0] node45012;
	wire [4-1:0] node45013;
	wire [4-1:0] node45016;
	wire [4-1:0] node45020;
	wire [4-1:0] node45021;
	wire [4-1:0] node45022;
	wire [4-1:0] node45023;
	wire [4-1:0] node45024;
	wire [4-1:0] node45028;
	wire [4-1:0] node45031;
	wire [4-1:0] node45032;
	wire [4-1:0] node45034;
	wire [4-1:0] node45037;
	wire [4-1:0] node45038;
	wire [4-1:0] node45041;
	wire [4-1:0] node45044;
	wire [4-1:0] node45045;
	wire [4-1:0] node45046;
	wire [4-1:0] node45047;
	wire [4-1:0] node45052;
	wire [4-1:0] node45053;
	wire [4-1:0] node45054;
	wire [4-1:0] node45059;
	wire [4-1:0] node45060;
	wire [4-1:0] node45061;
	wire [4-1:0] node45062;
	wire [4-1:0] node45063;
	wire [4-1:0] node45064;
	wire [4-1:0] node45065;
	wire [4-1:0] node45066;
	wire [4-1:0] node45070;
	wire [4-1:0] node45071;
	wire [4-1:0] node45075;
	wire [4-1:0] node45076;
	wire [4-1:0] node45077;
	wire [4-1:0] node45081;
	wire [4-1:0] node45082;
	wire [4-1:0] node45086;
	wire [4-1:0] node45087;
	wire [4-1:0] node45088;
	wire [4-1:0] node45089;
	wire [4-1:0] node45093;
	wire [4-1:0] node45094;
	wire [4-1:0] node45098;
	wire [4-1:0] node45099;
	wire [4-1:0] node45100;
	wire [4-1:0] node45104;
	wire [4-1:0] node45105;
	wire [4-1:0] node45109;
	wire [4-1:0] node45110;
	wire [4-1:0] node45111;
	wire [4-1:0] node45112;
	wire [4-1:0] node45113;
	wire [4-1:0] node45114;
	wire [4-1:0] node45117;
	wire [4-1:0] node45120;
	wire [4-1:0] node45121;
	wire [4-1:0] node45122;
	wire [4-1:0] node45125;
	wire [4-1:0] node45128;
	wire [4-1:0] node45129;
	wire [4-1:0] node45132;
	wire [4-1:0] node45135;
	wire [4-1:0] node45136;
	wire [4-1:0] node45137;
	wire [4-1:0] node45138;
	wire [4-1:0] node45141;
	wire [4-1:0] node45144;
	wire [4-1:0] node45145;
	wire [4-1:0] node45148;
	wire [4-1:0] node45151;
	wire [4-1:0] node45152;
	wire [4-1:0] node45155;
	wire [4-1:0] node45158;
	wire [4-1:0] node45159;
	wire [4-1:0] node45160;
	wire [4-1:0] node45161;
	wire [4-1:0] node45164;
	wire [4-1:0] node45167;
	wire [4-1:0] node45168;
	wire [4-1:0] node45171;
	wire [4-1:0] node45174;
	wire [4-1:0] node45175;
	wire [4-1:0] node45176;
	wire [4-1:0] node45179;
	wire [4-1:0] node45182;
	wire [4-1:0] node45184;
	wire [4-1:0] node45185;
	wire [4-1:0] node45188;
	wire [4-1:0] node45191;
	wire [4-1:0] node45192;
	wire [4-1:0] node45193;
	wire [4-1:0] node45194;
	wire [4-1:0] node45195;
	wire [4-1:0] node45198;
	wire [4-1:0] node45201;
	wire [4-1:0] node45202;
	wire [4-1:0] node45205;
	wire [4-1:0] node45208;
	wire [4-1:0] node45209;
	wire [4-1:0] node45210;
	wire [4-1:0] node45211;
	wire [4-1:0] node45214;
	wire [4-1:0] node45217;
	wire [4-1:0] node45218;
	wire [4-1:0] node45221;
	wire [4-1:0] node45224;
	wire [4-1:0] node45225;
	wire [4-1:0] node45228;
	wire [4-1:0] node45231;
	wire [4-1:0] node45232;
	wire [4-1:0] node45233;
	wire [4-1:0] node45236;
	wire [4-1:0] node45239;
	wire [4-1:0] node45240;
	wire [4-1:0] node45243;
	wire [4-1:0] node45246;
	wire [4-1:0] node45247;
	wire [4-1:0] node45248;
	wire [4-1:0] node45249;
	wire [4-1:0] node45250;
	wire [4-1:0] node45252;
	wire [4-1:0] node45255;
	wire [4-1:0] node45257;
	wire [4-1:0] node45260;
	wire [4-1:0] node45261;
	wire [4-1:0] node45263;
	wire [4-1:0] node45266;
	wire [4-1:0] node45268;
	wire [4-1:0] node45271;
	wire [4-1:0] node45272;
	wire [4-1:0] node45273;
	wire [4-1:0] node45274;
	wire [4-1:0] node45275;
	wire [4-1:0] node45277;
	wire [4-1:0] node45281;
	wire [4-1:0] node45282;
	wire [4-1:0] node45283;
	wire [4-1:0] node45287;
	wire [4-1:0] node45288;
	wire [4-1:0] node45291;
	wire [4-1:0] node45294;
	wire [4-1:0] node45295;
	wire [4-1:0] node45296;
	wire [4-1:0] node45299;
	wire [4-1:0] node45302;
	wire [4-1:0] node45303;
	wire [4-1:0] node45306;
	wire [4-1:0] node45309;
	wire [4-1:0] node45310;
	wire [4-1:0] node45311;
	wire [4-1:0] node45314;
	wire [4-1:0] node45317;
	wire [4-1:0] node45318;
	wire [4-1:0] node45321;
	wire [4-1:0] node45324;
	wire [4-1:0] node45325;
	wire [4-1:0] node45326;
	wire [4-1:0] node45327;
	wire [4-1:0] node45331;
	wire [4-1:0] node45332;
	wire [4-1:0] node45336;
	wire [4-1:0] node45337;
	wire [4-1:0] node45338;
	wire [4-1:0] node45342;
	wire [4-1:0] node45343;
	wire [4-1:0] node45347;
	wire [4-1:0] node45348;
	wire [4-1:0] node45349;
	wire [4-1:0] node45350;
	wire [4-1:0] node45351;
	wire [4-1:0] node45355;
	wire [4-1:0] node45356;
	wire [4-1:0] node45361;
	wire [4-1:0] node45362;
	wire [4-1:0] node45363;
	wire [4-1:0] node45364;
	wire [4-1:0] node45368;
	wire [4-1:0] node45369;
	wire [4-1:0] node45374;
	wire [4-1:0] node45375;
	wire [4-1:0] node45376;
	wire [4-1:0] node45377;
	wire [4-1:0] node45378;
	wire [4-1:0] node45379;
	wire [4-1:0] node45380;
	wire [4-1:0] node45381;
	wire [4-1:0] node45382;
	wire [4-1:0] node45383;
	wire [4-1:0] node45384;
	wire [4-1:0] node45385;
	wire [4-1:0] node45386;
	wire [4-1:0] node45387;
	wire [4-1:0] node45390;
	wire [4-1:0] node45393;
	wire [4-1:0] node45395;
	wire [4-1:0] node45398;
	wire [4-1:0] node45399;
	wire [4-1:0] node45403;
	wire [4-1:0] node45404;
	wire [4-1:0] node45405;
	wire [4-1:0] node45408;
	wire [4-1:0] node45411;
	wire [4-1:0] node45412;
	wire [4-1:0] node45415;
	wire [4-1:0] node45418;
	wire [4-1:0] node45419;
	wire [4-1:0] node45422;
	wire [4-1:0] node45425;
	wire [4-1:0] node45426;
	wire [4-1:0] node45427;
	wire [4-1:0] node45430;
	wire [4-1:0] node45433;
	wire [4-1:0] node45434;
	wire [4-1:0] node45437;
	wire [4-1:0] node45440;
	wire [4-1:0] node45441;
	wire [4-1:0] node45442;
	wire [4-1:0] node45443;
	wire [4-1:0] node45444;
	wire [4-1:0] node45445;
	wire [4-1:0] node45447;
	wire [4-1:0] node45450;
	wire [4-1:0] node45451;
	wire [4-1:0] node45454;
	wire [4-1:0] node45457;
	wire [4-1:0] node45458;
	wire [4-1:0] node45461;
	wire [4-1:0] node45464;
	wire [4-1:0] node45465;
	wire [4-1:0] node45468;
	wire [4-1:0] node45471;
	wire [4-1:0] node45472;
	wire [4-1:0] node45475;
	wire [4-1:0] node45478;
	wire [4-1:0] node45479;
	wire [4-1:0] node45480;
	wire [4-1:0] node45481;
	wire [4-1:0] node45482;
	wire [4-1:0] node45485;
	wire [4-1:0] node45488;
	wire [4-1:0] node45489;
	wire [4-1:0] node45492;
	wire [4-1:0] node45495;
	wire [4-1:0] node45496;
	wire [4-1:0] node45497;
	wire [4-1:0] node45500;
	wire [4-1:0] node45503;
	wire [4-1:0] node45504;
	wire [4-1:0] node45505;
	wire [4-1:0] node45508;
	wire [4-1:0] node45511;
	wire [4-1:0] node45512;
	wire [4-1:0] node45515;
	wire [4-1:0] node45518;
	wire [4-1:0] node45519;
	wire [4-1:0] node45520;
	wire [4-1:0] node45521;
	wire [4-1:0] node45524;
	wire [4-1:0] node45527;
	wire [4-1:0] node45528;
	wire [4-1:0] node45531;
	wire [4-1:0] node45534;
	wire [4-1:0] node45535;
	wire [4-1:0] node45536;
	wire [4-1:0] node45537;
	wire [4-1:0] node45540;
	wire [4-1:0] node45543;
	wire [4-1:0] node45544;
	wire [4-1:0] node45547;
	wire [4-1:0] node45550;
	wire [4-1:0] node45551;
	wire [4-1:0] node45552;
	wire [4-1:0] node45555;
	wire [4-1:0] node45558;
	wire [4-1:0] node45559;
	wire [4-1:0] node45562;
	wire [4-1:0] node45565;
	wire [4-1:0] node45566;
	wire [4-1:0] node45567;
	wire [4-1:0] node45568;
	wire [4-1:0] node45569;
	wire [4-1:0] node45570;
	wire [4-1:0] node45571;
	wire [4-1:0] node45572;
	wire [4-1:0] node45575;
	wire [4-1:0] node45578;
	wire [4-1:0] node45579;
	wire [4-1:0] node45583;
	wire [4-1:0] node45584;
	wire [4-1:0] node45587;
	wire [4-1:0] node45590;
	wire [4-1:0] node45591;
	wire [4-1:0] node45594;
	wire [4-1:0] node45595;
	wire [4-1:0] node45599;
	wire [4-1:0] node45600;
	wire [4-1:0] node45601;
	wire [4-1:0] node45604;
	wire [4-1:0] node45605;
	wire [4-1:0] node45609;
	wire [4-1:0] node45610;
	wire [4-1:0] node45612;
	wire [4-1:0] node45615;
	wire [4-1:0] node45618;
	wire [4-1:0] node45619;
	wire [4-1:0] node45620;
	wire [4-1:0] node45621;
	wire [4-1:0] node45624;
	wire [4-1:0] node45625;
	wire [4-1:0] node45629;
	wire [4-1:0] node45630;
	wire [4-1:0] node45633;
	wire [4-1:0] node45634;
	wire [4-1:0] node45638;
	wire [4-1:0] node45639;
	wire [4-1:0] node45640;
	wire [4-1:0] node45643;
	wire [4-1:0] node45644;
	wire [4-1:0] node45648;
	wire [4-1:0] node45649;
	wire [4-1:0] node45651;
	wire [4-1:0] node45654;
	wire [4-1:0] node45657;
	wire [4-1:0] node45658;
	wire [4-1:0] node45659;
	wire [4-1:0] node45660;
	wire [4-1:0] node45661;
	wire [4-1:0] node45662;
	wire [4-1:0] node45665;
	wire [4-1:0] node45668;
	wire [4-1:0] node45669;
	wire [4-1:0] node45672;
	wire [4-1:0] node45675;
	wire [4-1:0] node45676;
	wire [4-1:0] node45677;
	wire [4-1:0] node45680;
	wire [4-1:0] node45683;
	wire [4-1:0] node45684;
	wire [4-1:0] node45685;
	wire [4-1:0] node45688;
	wire [4-1:0] node45692;
	wire [4-1:0] node45693;
	wire [4-1:0] node45694;
	wire [4-1:0] node45696;
	wire [4-1:0] node45699;
	wire [4-1:0] node45702;
	wire [4-1:0] node45703;
	wire [4-1:0] node45706;
	wire [4-1:0] node45707;
	wire [4-1:0] node45711;
	wire [4-1:0] node45712;
	wire [4-1:0] node45713;
	wire [4-1:0] node45714;
	wire [4-1:0] node45715;
	wire [4-1:0] node45716;
	wire [4-1:0] node45719;
	wire [4-1:0] node45722;
	wire [4-1:0] node45723;
	wire [4-1:0] node45726;
	wire [4-1:0] node45729;
	wire [4-1:0] node45730;
	wire [4-1:0] node45733;
	wire [4-1:0] node45736;
	wire [4-1:0] node45737;
	wire [4-1:0] node45738;
	wire [4-1:0] node45739;
	wire [4-1:0] node45742;
	wire [4-1:0] node45745;
	wire [4-1:0] node45746;
	wire [4-1:0] node45749;
	wire [4-1:0] node45752;
	wire [4-1:0] node45754;
	wire [4-1:0] node45757;
	wire [4-1:0] node45758;
	wire [4-1:0] node45760;
	wire [4-1:0] node45761;
	wire [4-1:0] node45762;
	wire [4-1:0] node45767;
	wire [4-1:0] node45768;
	wire [4-1:0] node45771;
	wire [4-1:0] node45774;
	wire [4-1:0] node45775;
	wire [4-1:0] node45776;
	wire [4-1:0] node45777;
	wire [4-1:0] node45778;
	wire [4-1:0] node45779;
	wire [4-1:0] node45780;
	wire [4-1:0] node45782;
	wire [4-1:0] node45785;
	wire [4-1:0] node45786;
	wire [4-1:0] node45789;
	wire [4-1:0] node45792;
	wire [4-1:0] node45793;
	wire [4-1:0] node45794;
	wire [4-1:0] node45797;
	wire [4-1:0] node45800;
	wire [4-1:0] node45801;
	wire [4-1:0] node45804;
	wire [4-1:0] node45807;
	wire [4-1:0] node45808;
	wire [4-1:0] node45809;
	wire [4-1:0] node45811;
	wire [4-1:0] node45814;
	wire [4-1:0] node45815;
	wire [4-1:0] node45818;
	wire [4-1:0] node45821;
	wire [4-1:0] node45822;
	wire [4-1:0] node45824;
	wire [4-1:0] node45827;
	wire [4-1:0] node45828;
	wire [4-1:0] node45831;
	wire [4-1:0] node45834;
	wire [4-1:0] node45835;
	wire [4-1:0] node45836;
	wire [4-1:0] node45837;
	wire [4-1:0] node45839;
	wire [4-1:0] node45842;
	wire [4-1:0] node45844;
	wire [4-1:0] node45847;
	wire [4-1:0] node45848;
	wire [4-1:0] node45850;
	wire [4-1:0] node45853;
	wire [4-1:0] node45854;
	wire [4-1:0] node45857;
	wire [4-1:0] node45860;
	wire [4-1:0] node45861;
	wire [4-1:0] node45862;
	wire [4-1:0] node45865;
	wire [4-1:0] node45866;
	wire [4-1:0] node45869;
	wire [4-1:0] node45872;
	wire [4-1:0] node45873;
	wire [4-1:0] node45874;
	wire [4-1:0] node45877;
	wire [4-1:0] node45880;
	wire [4-1:0] node45881;
	wire [4-1:0] node45884;
	wire [4-1:0] node45887;
	wire [4-1:0] node45888;
	wire [4-1:0] node45889;
	wire [4-1:0] node45890;
	wire [4-1:0] node45891;
	wire [4-1:0] node45892;
	wire [4-1:0] node45894;
	wire [4-1:0] node45897;
	wire [4-1:0] node45898;
	wire [4-1:0] node45901;
	wire [4-1:0] node45904;
	wire [4-1:0] node45905;
	wire [4-1:0] node45906;
	wire [4-1:0] node45909;
	wire [4-1:0] node45912;
	wire [4-1:0] node45913;
	wire [4-1:0] node45916;
	wire [4-1:0] node45919;
	wire [4-1:0] node45920;
	wire [4-1:0] node45921;
	wire [4-1:0] node45922;
	wire [4-1:0] node45926;
	wire [4-1:0] node45927;
	wire [4-1:0] node45930;
	wire [4-1:0] node45933;
	wire [4-1:0] node45934;
	wire [4-1:0] node45935;
	wire [4-1:0] node45938;
	wire [4-1:0] node45941;
	wire [4-1:0] node45942;
	wire [4-1:0] node45946;
	wire [4-1:0] node45947;
	wire [4-1:0] node45948;
	wire [4-1:0] node45949;
	wire [4-1:0] node45952;
	wire [4-1:0] node45955;
	wire [4-1:0] node45956;
	wire [4-1:0] node45957;
	wire [4-1:0] node45960;
	wire [4-1:0] node45964;
	wire [4-1:0] node45965;
	wire [4-1:0] node45967;
	wire [4-1:0] node45968;
	wire [4-1:0] node45971;
	wire [4-1:0] node45974;
	wire [4-1:0] node45975;
	wire [4-1:0] node45976;
	wire [4-1:0] node45979;
	wire [4-1:0] node45982;
	wire [4-1:0] node45983;
	wire [4-1:0] node45986;
	wire [4-1:0] node45989;
	wire [4-1:0] node45990;
	wire [4-1:0] node45991;
	wire [4-1:0] node45992;
	wire [4-1:0] node45993;
	wire [4-1:0] node45996;
	wire [4-1:0] node45999;
	wire [4-1:0] node46000;
	wire [4-1:0] node46003;
	wire [4-1:0] node46006;
	wire [4-1:0] node46007;
	wire [4-1:0] node46008;
	wire [4-1:0] node46011;
	wire [4-1:0] node46014;
	wire [4-1:0] node46015;
	wire [4-1:0] node46018;
	wire [4-1:0] node46021;
	wire [4-1:0] node46022;
	wire [4-1:0] node46023;
	wire [4-1:0] node46024;
	wire [4-1:0] node46027;
	wire [4-1:0] node46030;
	wire [4-1:0] node46031;
	wire [4-1:0] node46034;
	wire [4-1:0] node46037;
	wire [4-1:0] node46038;
	wire [4-1:0] node46039;
	wire [4-1:0] node46042;
	wire [4-1:0] node46045;
	wire [4-1:0] node46046;
	wire [4-1:0] node46049;
	wire [4-1:0] node46052;
	wire [4-1:0] node46053;
	wire [4-1:0] node46054;
	wire [4-1:0] node46055;
	wire [4-1:0] node46056;
	wire [4-1:0] node46057;
	wire [4-1:0] node46058;
	wire [4-1:0] node46061;
	wire [4-1:0] node46064;
	wire [4-1:0] node46065;
	wire [4-1:0] node46068;
	wire [4-1:0] node46071;
	wire [4-1:0] node46072;
	wire [4-1:0] node46073;
	wire [4-1:0] node46076;
	wire [4-1:0] node46079;
	wire [4-1:0] node46080;
	wire [4-1:0] node46084;
	wire [4-1:0] node46085;
	wire [4-1:0] node46086;
	wire [4-1:0] node46087;
	wire [4-1:0] node46090;
	wire [4-1:0] node46093;
	wire [4-1:0] node46094;
	wire [4-1:0] node46097;
	wire [4-1:0] node46100;
	wire [4-1:0] node46101;
	wire [4-1:0] node46102;
	wire [4-1:0] node46103;
	wire [4-1:0] node46106;
	wire [4-1:0] node46109;
	wire [4-1:0] node46110;
	wire [4-1:0] node46113;
	wire [4-1:0] node46116;
	wire [4-1:0] node46117;
	wire [4-1:0] node46120;
	wire [4-1:0] node46123;
	wire [4-1:0] node46124;
	wire [4-1:0] node46125;
	wire [4-1:0] node46126;
	wire [4-1:0] node46127;
	wire [4-1:0] node46130;
	wire [4-1:0] node46133;
	wire [4-1:0] node46134;
	wire [4-1:0] node46137;
	wire [4-1:0] node46140;
	wire [4-1:0] node46141;
	wire [4-1:0] node46142;
	wire [4-1:0] node46143;
	wire [4-1:0] node46146;
	wire [4-1:0] node46149;
	wire [4-1:0] node46150;
	wire [4-1:0] node46153;
	wire [4-1:0] node46156;
	wire [4-1:0] node46157;
	wire [4-1:0] node46160;
	wire [4-1:0] node46163;
	wire [4-1:0] node46164;
	wire [4-1:0] node46165;
	wire [4-1:0] node46166;
	wire [4-1:0] node46167;
	wire [4-1:0] node46170;
	wire [4-1:0] node46173;
	wire [4-1:0] node46174;
	wire [4-1:0] node46177;
	wire [4-1:0] node46180;
	wire [4-1:0] node46181;
	wire [4-1:0] node46182;
	wire [4-1:0] node46185;
	wire [4-1:0] node46188;
	wire [4-1:0] node46189;
	wire [4-1:0] node46192;
	wire [4-1:0] node46195;
	wire [4-1:0] node46196;
	wire [4-1:0] node46198;
	wire [4-1:0] node46201;
	wire [4-1:0] node46202;
	wire [4-1:0] node46203;
	wire [4-1:0] node46207;
	wire [4-1:0] node46209;
	wire [4-1:0] node46212;
	wire [4-1:0] node46213;
	wire [4-1:0] node46214;
	wire [4-1:0] node46215;
	wire [4-1:0] node46216;
	wire [4-1:0] node46219;
	wire [4-1:0] node46222;
	wire [4-1:0] node46223;
	wire [4-1:0] node46224;
	wire [4-1:0] node46227;
	wire [4-1:0] node46230;
	wire [4-1:0] node46231;
	wire [4-1:0] node46232;
	wire [4-1:0] node46235;
	wire [4-1:0] node46238;
	wire [4-1:0] node46239;
	wire [4-1:0] node46242;
	wire [4-1:0] node46245;
	wire [4-1:0] node46246;
	wire [4-1:0] node46247;
	wire [4-1:0] node46250;
	wire [4-1:0] node46253;
	wire [4-1:0] node46254;
	wire [4-1:0] node46255;
	wire [4-1:0] node46258;
	wire [4-1:0] node46261;
	wire [4-1:0] node46262;
	wire [4-1:0] node46265;
	wire [4-1:0] node46268;
	wire [4-1:0] node46269;
	wire [4-1:0] node46270;
	wire [4-1:0] node46271;
	wire [4-1:0] node46272;
	wire [4-1:0] node46275;
	wire [4-1:0] node46278;
	wire [4-1:0] node46279;
	wire [4-1:0] node46282;
	wire [4-1:0] node46285;
	wire [4-1:0] node46286;
	wire [4-1:0] node46287;
	wire [4-1:0] node46291;
	wire [4-1:0] node46292;
	wire [4-1:0] node46295;
	wire [4-1:0] node46298;
	wire [4-1:0] node46299;
	wire [4-1:0] node46300;
	wire [4-1:0] node46301;
	wire [4-1:0] node46304;
	wire [4-1:0] node46307;
	wire [4-1:0] node46308;
	wire [4-1:0] node46309;
	wire [4-1:0] node46312;
	wire [4-1:0] node46315;
	wire [4-1:0] node46316;
	wire [4-1:0] node46319;
	wire [4-1:0] node46322;
	wire [4-1:0] node46323;
	wire [4-1:0] node46324;
	wire [4-1:0] node46327;
	wire [4-1:0] node46330;
	wire [4-1:0] node46332;
	wire [4-1:0] node46334;
	wire [4-1:0] node46337;
	wire [4-1:0] node46338;
	wire [4-1:0] node46339;
	wire [4-1:0] node46340;
	wire [4-1:0] node46341;
	wire [4-1:0] node46342;
	wire [4-1:0] node46343;
	wire [4-1:0] node46344;
	wire [4-1:0] node46346;
	wire [4-1:0] node46347;
	wire [4-1:0] node46350;
	wire [4-1:0] node46353;
	wire [4-1:0] node46355;
	wire [4-1:0] node46356;
	wire [4-1:0] node46359;
	wire [4-1:0] node46362;
	wire [4-1:0] node46363;
	wire [4-1:0] node46365;
	wire [4-1:0] node46367;
	wire [4-1:0] node46370;
	wire [4-1:0] node46372;
	wire [4-1:0] node46373;
	wire [4-1:0] node46376;
	wire [4-1:0] node46379;
	wire [4-1:0] node46380;
	wire [4-1:0] node46381;
	wire [4-1:0] node46382;
	wire [4-1:0] node46385;
	wire [4-1:0] node46388;
	wire [4-1:0] node46390;
	wire [4-1:0] node46392;
	wire [4-1:0] node46395;
	wire [4-1:0] node46396;
	wire [4-1:0] node46397;
	wire [4-1:0] node46398;
	wire [4-1:0] node46402;
	wire [4-1:0] node46404;
	wire [4-1:0] node46407;
	wire [4-1:0] node46408;
	wire [4-1:0] node46412;
	wire [4-1:0] node46413;
	wire [4-1:0] node46414;
	wire [4-1:0] node46415;
	wire [4-1:0] node46416;
	wire [4-1:0] node46418;
	wire [4-1:0] node46421;
	wire [4-1:0] node46423;
	wire [4-1:0] node46426;
	wire [4-1:0] node46427;
	wire [4-1:0] node46429;
	wire [4-1:0] node46432;
	wire [4-1:0] node46434;
	wire [4-1:0] node46437;
	wire [4-1:0] node46438;
	wire [4-1:0] node46439;
	wire [4-1:0] node46441;
	wire [4-1:0] node46444;
	wire [4-1:0] node46446;
	wire [4-1:0] node46449;
	wire [4-1:0] node46450;
	wire [4-1:0] node46452;
	wire [4-1:0] node46456;
	wire [4-1:0] node46457;
	wire [4-1:0] node46458;
	wire [4-1:0] node46459;
	wire [4-1:0] node46460;
	wire [4-1:0] node46464;
	wire [4-1:0] node46465;
	wire [4-1:0] node46468;
	wire [4-1:0] node46471;
	wire [4-1:0] node46472;
	wire [4-1:0] node46473;
	wire [4-1:0] node46476;
	wire [4-1:0] node46479;
	wire [4-1:0] node46480;
	wire [4-1:0] node46483;
	wire [4-1:0] node46486;
	wire [4-1:0] node46487;
	wire [4-1:0] node46490;
	wire [4-1:0] node46493;
	wire [4-1:0] node46494;
	wire [4-1:0] node46495;
	wire [4-1:0] node46496;
	wire [4-1:0] node46497;
	wire [4-1:0] node46499;
	wire [4-1:0] node46502;
	wire [4-1:0] node46503;
	wire [4-1:0] node46506;
	wire [4-1:0] node46509;
	wire [4-1:0] node46510;
	wire [4-1:0] node46513;
	wire [4-1:0] node46516;
	wire [4-1:0] node46517;
	wire [4-1:0] node46518;
	wire [4-1:0] node46519;
	wire [4-1:0] node46520;
	wire [4-1:0] node46523;
	wire [4-1:0] node46526;
	wire [4-1:0] node46527;
	wire [4-1:0] node46530;
	wire [4-1:0] node46533;
	wire [4-1:0] node46534;
	wire [4-1:0] node46536;
	wire [4-1:0] node46539;
	wire [4-1:0] node46540;
	wire [4-1:0] node46543;
	wire [4-1:0] node46546;
	wire [4-1:0] node46547;
	wire [4-1:0] node46548;
	wire [4-1:0] node46549;
	wire [4-1:0] node46552;
	wire [4-1:0] node46555;
	wire [4-1:0] node46556;
	wire [4-1:0] node46559;
	wire [4-1:0] node46562;
	wire [4-1:0] node46563;
	wire [4-1:0] node46564;
	wire [4-1:0] node46567;
	wire [4-1:0] node46570;
	wire [4-1:0] node46571;
	wire [4-1:0] node46574;
	wire [4-1:0] node46577;
	wire [4-1:0] node46578;
	wire [4-1:0] node46579;
	wire [4-1:0] node46580;
	wire [4-1:0] node46581;
	wire [4-1:0] node46582;
	wire [4-1:0] node46585;
	wire [4-1:0] node46588;
	wire [4-1:0] node46589;
	wire [4-1:0] node46592;
	wire [4-1:0] node46595;
	wire [4-1:0] node46596;
	wire [4-1:0] node46597;
	wire [4-1:0] node46600;
	wire [4-1:0] node46603;
	wire [4-1:0] node46605;
	wire [4-1:0] node46608;
	wire [4-1:0] node46609;
	wire [4-1:0] node46612;
	wire [4-1:0] node46615;
	wire [4-1:0] node46616;
	wire [4-1:0] node46617;
	wire [4-1:0] node46618;
	wire [4-1:0] node46619;
	wire [4-1:0] node46622;
	wire [4-1:0] node46625;
	wire [4-1:0] node46626;
	wire [4-1:0] node46629;
	wire [4-1:0] node46632;
	wire [4-1:0] node46633;
	wire [4-1:0] node46636;
	wire [4-1:0] node46639;
	wire [4-1:0] node46640;
	wire [4-1:0] node46642;
	wire [4-1:0] node46645;
	wire [4-1:0] node46646;
	wire [4-1:0] node46647;
	wire [4-1:0] node46650;
	wire [4-1:0] node46653;
	wire [4-1:0] node46654;
	wire [4-1:0] node46658;
	wire [4-1:0] node46659;
	wire [4-1:0] node46660;
	wire [4-1:0] node46661;
	wire [4-1:0] node46662;
	wire [4-1:0] node46663;
	wire [4-1:0] node46665;
	wire [4-1:0] node46668;
	wire [4-1:0] node46670;
	wire [4-1:0] node46673;
	wire [4-1:0] node46674;
	wire [4-1:0] node46676;
	wire [4-1:0] node46679;
	wire [4-1:0] node46681;
	wire [4-1:0] node46684;
	wire [4-1:0] node46685;
	wire [4-1:0] node46686;
	wire [4-1:0] node46687;
	wire [4-1:0] node46689;
	wire [4-1:0] node46693;
	wire [4-1:0] node46695;
	wire [4-1:0] node46697;
	wire [4-1:0] node46700;
	wire [4-1:0] node46701;
	wire [4-1:0] node46702;
	wire [4-1:0] node46705;
	wire [4-1:0] node46708;
	wire [4-1:0] node46709;
	wire [4-1:0] node46710;
	wire [4-1:0] node46713;
	wire [4-1:0] node46716;
	wire [4-1:0] node46717;
	wire [4-1:0] node46720;
	wire [4-1:0] node46723;
	wire [4-1:0] node46724;
	wire [4-1:0] node46725;
	wire [4-1:0] node46727;
	wire [4-1:0] node46728;
	wire [4-1:0] node46731;
	wire [4-1:0] node46734;
	wire [4-1:0] node46736;
	wire [4-1:0] node46737;
	wire [4-1:0] node46738;
	wire [4-1:0] node46741;
	wire [4-1:0] node46745;
	wire [4-1:0] node46746;
	wire [4-1:0] node46748;
	wire [4-1:0] node46749;
	wire [4-1:0] node46752;
	wire [4-1:0] node46755;
	wire [4-1:0] node46757;
	wire [4-1:0] node46758;
	wire [4-1:0] node46759;
	wire [4-1:0] node46762;
	wire [4-1:0] node46765;
	wire [4-1:0] node46766;
	wire [4-1:0] node46769;
	wire [4-1:0] node46772;
	wire [4-1:0] node46773;
	wire [4-1:0] node46774;
	wire [4-1:0] node46775;
	wire [4-1:0] node46776;
	wire [4-1:0] node46779;
	wire [4-1:0] node46782;
	wire [4-1:0] node46783;
	wire [4-1:0] node46784;
	wire [4-1:0] node46787;
	wire [4-1:0] node46790;
	wire [4-1:0] node46791;
	wire [4-1:0] node46792;
	wire [4-1:0] node46795;
	wire [4-1:0] node46798;
	wire [4-1:0] node46799;
	wire [4-1:0] node46802;
	wire [4-1:0] node46805;
	wire [4-1:0] node46806;
	wire [4-1:0] node46807;
	wire [4-1:0] node46808;
	wire [4-1:0] node46809;
	wire [4-1:0] node46813;
	wire [4-1:0] node46815;
	wire [4-1:0] node46818;
	wire [4-1:0] node46819;
	wire [4-1:0] node46820;
	wire [4-1:0] node46824;
	wire [4-1:0] node46825;
	wire [4-1:0] node46829;
	wire [4-1:0] node46830;
	wire [4-1:0] node46832;
	wire [4-1:0] node46833;
	wire [4-1:0] node46837;
	wire [4-1:0] node46838;
	wire [4-1:0] node46840;
	wire [4-1:0] node46844;
	wire [4-1:0] node46845;
	wire [4-1:0] node46846;
	wire [4-1:0] node46847;
	wire [4-1:0] node46848;
	wire [4-1:0] node46849;
	wire [4-1:0] node46852;
	wire [4-1:0] node46855;
	wire [4-1:0] node46856;
	wire [4-1:0] node46859;
	wire [4-1:0] node46862;
	wire [4-1:0] node46863;
	wire [4-1:0] node46866;
	wire [4-1:0] node46869;
	wire [4-1:0] node46870;
	wire [4-1:0] node46872;
	wire [4-1:0] node46874;
	wire [4-1:0] node46877;
	wire [4-1:0] node46878;
	wire [4-1:0] node46880;
	wire [4-1:0] node46883;
	wire [4-1:0] node46884;
	wire [4-1:0] node46888;
	wire [4-1:0] node46889;
	wire [4-1:0] node46890;
	wire [4-1:0] node46891;
	wire [4-1:0] node46893;
	wire [4-1:0] node46897;
	wire [4-1:0] node46898;
	wire [4-1:0] node46899;
	wire [4-1:0] node46902;
	wire [4-1:0] node46906;
	wire [4-1:0] node46907;
	wire [4-1:0] node46908;
	wire [4-1:0] node46909;
	wire [4-1:0] node46912;
	wire [4-1:0] node46916;
	wire [4-1:0] node46917;
	wire [4-1:0] node46918;
	wire [4-1:0] node46921;
	wire [4-1:0] node46925;
	wire [4-1:0] node46926;
	wire [4-1:0] node46927;
	wire [4-1:0] node46928;
	wire [4-1:0] node46929;
	wire [4-1:0] node46930;
	wire [4-1:0] node46931;
	wire [4-1:0] node46933;
	wire [4-1:0] node46936;
	wire [4-1:0] node46938;
	wire [4-1:0] node46941;
	wire [4-1:0] node46942;
	wire [4-1:0] node46944;
	wire [4-1:0] node46947;
	wire [4-1:0] node46949;
	wire [4-1:0] node46952;
	wire [4-1:0] node46953;
	wire [4-1:0] node46954;
	wire [4-1:0] node46957;
	wire [4-1:0] node46960;
	wire [4-1:0] node46961;
	wire [4-1:0] node46962;
	wire [4-1:0] node46965;
	wire [4-1:0] node46968;
	wire [4-1:0] node46969;
	wire [4-1:0] node46972;
	wire [4-1:0] node46975;
	wire [4-1:0] node46976;
	wire [4-1:0] node46977;
	wire [4-1:0] node46978;
	wire [4-1:0] node46980;
	wire [4-1:0] node46983;
	wire [4-1:0] node46984;
	wire [4-1:0] node46986;
	wire [4-1:0] node46989;
	wire [4-1:0] node46991;
	wire [4-1:0] node46994;
	wire [4-1:0] node46995;
	wire [4-1:0] node46996;
	wire [4-1:0] node46999;
	wire [4-1:0] node47002;
	wire [4-1:0] node47003;
	wire [4-1:0] node47004;
	wire [4-1:0] node47007;
	wire [4-1:0] node47010;
	wire [4-1:0] node47011;
	wire [4-1:0] node47015;
	wire [4-1:0] node47016;
	wire [4-1:0] node47017;
	wire [4-1:0] node47018;
	wire [4-1:0] node47022;
	wire [4-1:0] node47023;
	wire [4-1:0] node47027;
	wire [4-1:0] node47028;
	wire [4-1:0] node47029;
	wire [4-1:0] node47033;
	wire [4-1:0] node47034;
	wire [4-1:0] node47038;
	wire [4-1:0] node47039;
	wire [4-1:0] node47040;
	wire [4-1:0] node47041;
	wire [4-1:0] node47042;
	wire [4-1:0] node47043;
	wire [4-1:0] node47046;
	wire [4-1:0] node47049;
	wire [4-1:0] node47050;
	wire [4-1:0] node47054;
	wire [4-1:0] node47055;
	wire [4-1:0] node47056;
	wire [4-1:0] node47059;
	wire [4-1:0] node47062;
	wire [4-1:0] node47063;
	wire [4-1:0] node47066;
	wire [4-1:0] node47069;
	wire [4-1:0] node47070;
	wire [4-1:0] node47071;
	wire [4-1:0] node47072;
	wire [4-1:0] node47075;
	wire [4-1:0] node47078;
	wire [4-1:0] node47079;
	wire [4-1:0] node47082;
	wire [4-1:0] node47085;
	wire [4-1:0] node47086;
	wire [4-1:0] node47087;
	wire [4-1:0] node47091;
	wire [4-1:0] node47092;
	wire [4-1:0] node47093;
	wire [4-1:0] node47096;
	wire [4-1:0] node47100;
	wire [4-1:0] node47101;
	wire [4-1:0] node47102;
	wire [4-1:0] node47103;
	wire [4-1:0] node47104;
	wire [4-1:0] node47107;
	wire [4-1:0] node47110;
	wire [4-1:0] node47111;
	wire [4-1:0] node47112;
	wire [4-1:0] node47115;
	wire [4-1:0] node47119;
	wire [4-1:0] node47120;
	wire [4-1:0] node47121;
	wire [4-1:0] node47122;
	wire [4-1:0] node47126;
	wire [4-1:0] node47127;
	wire [4-1:0] node47130;
	wire [4-1:0] node47133;
	wire [4-1:0] node47134;
	wire [4-1:0] node47135;
	wire [4-1:0] node47138;
	wire [4-1:0] node47141;
	wire [4-1:0] node47142;
	wire [4-1:0] node47145;
	wire [4-1:0] node47148;
	wire [4-1:0] node47149;
	wire [4-1:0] node47150;
	wire [4-1:0] node47151;
	wire [4-1:0] node47152;
	wire [4-1:0] node47156;
	wire [4-1:0] node47157;
	wire [4-1:0] node47160;
	wire [4-1:0] node47163;
	wire [4-1:0] node47164;
	wire [4-1:0] node47165;
	wire [4-1:0] node47169;
	wire [4-1:0] node47170;
	wire [4-1:0] node47173;
	wire [4-1:0] node47176;
	wire [4-1:0] node47177;
	wire [4-1:0] node47178;
	wire [4-1:0] node47180;
	wire [4-1:0] node47183;
	wire [4-1:0] node47186;
	wire [4-1:0] node47187;
	wire [4-1:0] node47189;
	wire [4-1:0] node47192;
	wire [4-1:0] node47195;
	wire [4-1:0] node47196;
	wire [4-1:0] node47197;
	wire [4-1:0] node47198;
	wire [4-1:0] node47199;
	wire [4-1:0] node47200;
	wire [4-1:0] node47201;
	wire [4-1:0] node47202;
	wire [4-1:0] node47205;
	wire [4-1:0] node47208;
	wire [4-1:0] node47209;
	wire [4-1:0] node47212;
	wire [4-1:0] node47215;
	wire [4-1:0] node47217;
	wire [4-1:0] node47219;
	wire [4-1:0] node47222;
	wire [4-1:0] node47223;
	wire [4-1:0] node47224;
	wire [4-1:0] node47226;
	wire [4-1:0] node47229;
	wire [4-1:0] node47231;
	wire [4-1:0] node47234;
	wire [4-1:0] node47235;
	wire [4-1:0] node47236;
	wire [4-1:0] node47239;
	wire [4-1:0] node47242;
	wire [4-1:0] node47243;
	wire [4-1:0] node47246;
	wire [4-1:0] node47249;
	wire [4-1:0] node47250;
	wire [4-1:0] node47251;
	wire [4-1:0] node47253;
	wire [4-1:0] node47254;
	wire [4-1:0] node47258;
	wire [4-1:0] node47259;
	wire [4-1:0] node47260;
	wire [4-1:0] node47263;
	wire [4-1:0] node47266;
	wire [4-1:0] node47267;
	wire [4-1:0] node47270;
	wire [4-1:0] node47273;
	wire [4-1:0] node47274;
	wire [4-1:0] node47275;
	wire [4-1:0] node47276;
	wire [4-1:0] node47280;
	wire [4-1:0] node47281;
	wire [4-1:0] node47284;
	wire [4-1:0] node47287;
	wire [4-1:0] node47288;
	wire [4-1:0] node47289;
	wire [4-1:0] node47292;
	wire [4-1:0] node47295;
	wire [4-1:0] node47296;
	wire [4-1:0] node47299;
	wire [4-1:0] node47302;
	wire [4-1:0] node47303;
	wire [4-1:0] node47304;
	wire [4-1:0] node47305;
	wire [4-1:0] node47306;
	wire [4-1:0] node47307;
	wire [4-1:0] node47310;
	wire [4-1:0] node47313;
	wire [4-1:0] node47314;
	wire [4-1:0] node47317;
	wire [4-1:0] node47320;
	wire [4-1:0] node47321;
	wire [4-1:0] node47322;
	wire [4-1:0] node47326;
	wire [4-1:0] node47328;
	wire [4-1:0] node47331;
	wire [4-1:0] node47332;
	wire [4-1:0] node47333;
	wire [4-1:0] node47334;
	wire [4-1:0] node47337;
	wire [4-1:0] node47340;
	wire [4-1:0] node47341;
	wire [4-1:0] node47344;
	wire [4-1:0] node47347;
	wire [4-1:0] node47348;
	wire [4-1:0] node47349;
	wire [4-1:0] node47352;
	wire [4-1:0] node47355;
	wire [4-1:0] node47356;
	wire [4-1:0] node47359;
	wire [4-1:0] node47362;
	wire [4-1:0] node47363;
	wire [4-1:0] node47364;
	wire [4-1:0] node47365;
	wire [4-1:0] node47368;
	wire [4-1:0] node47371;
	wire [4-1:0] node47372;
	wire [4-1:0] node47375;
	wire [4-1:0] node47378;
	wire [4-1:0] node47379;
	wire [4-1:0] node47381;
	wire [4-1:0] node47382;
	wire [4-1:0] node47385;
	wire [4-1:0] node47388;
	wire [4-1:0] node47389;
	wire [4-1:0] node47390;
	wire [4-1:0] node47393;
	wire [4-1:0] node47397;
	wire [4-1:0] node47398;
	wire [4-1:0] node47399;
	wire [4-1:0] node47400;
	wire [4-1:0] node47401;
	wire [4-1:0] node47402;
	wire [4-1:0] node47405;
	wire [4-1:0] node47408;
	wire [4-1:0] node47409;
	wire [4-1:0] node47413;
	wire [4-1:0] node47414;
	wire [4-1:0] node47415;
	wire [4-1:0] node47418;
	wire [4-1:0] node47421;
	wire [4-1:0] node47422;
	wire [4-1:0] node47425;
	wire [4-1:0] node47428;
	wire [4-1:0] node47429;
	wire [4-1:0] node47430;
	wire [4-1:0] node47431;
	wire [4-1:0] node47435;
	wire [4-1:0] node47436;
	wire [4-1:0] node47439;
	wire [4-1:0] node47442;
	wire [4-1:0] node47443;
	wire [4-1:0] node47444;
	wire [4-1:0] node47447;
	wire [4-1:0] node47450;
	wire [4-1:0] node47452;
	wire [4-1:0] node47455;
	wire [4-1:0] node47456;
	wire [4-1:0] node47457;
	wire [4-1:0] node47458;
	wire [4-1:0] node47459;
	wire [4-1:0] node47462;
	wire [4-1:0] node47465;
	wire [4-1:0] node47466;
	wire [4-1:0] node47469;
	wire [4-1:0] node47472;
	wire [4-1:0] node47473;
	wire [4-1:0] node47474;
	wire [4-1:0] node47477;
	wire [4-1:0] node47480;
	wire [4-1:0] node47481;
	wire [4-1:0] node47484;
	wire [4-1:0] node47487;
	wire [4-1:0] node47488;
	wire [4-1:0] node47489;
	wire [4-1:0] node47490;
	wire [4-1:0] node47493;
	wire [4-1:0] node47496;
	wire [4-1:0] node47497;
	wire [4-1:0] node47500;
	wire [4-1:0] node47503;
	wire [4-1:0] node47504;
	wire [4-1:0] node47505;
	wire [4-1:0] node47508;
	wire [4-1:0] node47511;
	wire [4-1:0] node47512;
	wire [4-1:0] node47515;
	wire [4-1:0] node47518;
	wire [4-1:0] node47519;
	wire [4-1:0] node47520;
	wire [4-1:0] node47521;
	wire [4-1:0] node47522;
	wire [4-1:0] node47523;
	wire [4-1:0] node47524;
	wire [4-1:0] node47525;
	wire [4-1:0] node47526;
	wire [4-1:0] node47527;
	wire [4-1:0] node47531;
	wire [4-1:0] node47532;
	wire [4-1:0] node47536;
	wire [4-1:0] node47537;
	wire [4-1:0] node47539;
	wire [4-1:0] node47542;
	wire [4-1:0] node47544;
	wire [4-1:0] node47547;
	wire [4-1:0] node47548;
	wire [4-1:0] node47549;
	wire [4-1:0] node47550;
	wire [4-1:0] node47551;
	wire [4-1:0] node47554;
	wire [4-1:0] node47557;
	wire [4-1:0] node47558;
	wire [4-1:0] node47561;
	wire [4-1:0] node47564;
	wire [4-1:0] node47565;
	wire [4-1:0] node47567;
	wire [4-1:0] node47570;
	wire [4-1:0] node47571;
	wire [4-1:0] node47574;
	wire [4-1:0] node47577;
	wire [4-1:0] node47578;
	wire [4-1:0] node47579;
	wire [4-1:0] node47580;
	wire [4-1:0] node47584;
	wire [4-1:0] node47585;
	wire [4-1:0] node47589;
	wire [4-1:0] node47590;
	wire [4-1:0] node47593;
	wire [4-1:0] node47596;
	wire [4-1:0] node47597;
	wire [4-1:0] node47598;
	wire [4-1:0] node47601;
	wire [4-1:0] node47604;
	wire [4-1:0] node47605;
	wire [4-1:0] node47606;
	wire [4-1:0] node47609;
	wire [4-1:0] node47612;
	wire [4-1:0] node47613;
	wire [4-1:0] node47614;
	wire [4-1:0] node47617;
	wire [4-1:0] node47620;
	wire [4-1:0] node47621;
	wire [4-1:0] node47622;
	wire [4-1:0] node47626;
	wire [4-1:0] node47627;
	wire [4-1:0] node47630;
	wire [4-1:0] node47633;
	wire [4-1:0] node47634;
	wire [4-1:0] node47635;
	wire [4-1:0] node47636;
	wire [4-1:0] node47638;
	wire [4-1:0] node47641;
	wire [4-1:0] node47642;
	wire [4-1:0] node47646;
	wire [4-1:0] node47647;
	wire [4-1:0] node47649;
	wire [4-1:0] node47652;
	wire [4-1:0] node47654;
	wire [4-1:0] node47657;
	wire [4-1:0] node47658;
	wire [4-1:0] node47659;
	wire [4-1:0] node47660;
	wire [4-1:0] node47664;
	wire [4-1:0] node47666;
	wire [4-1:0] node47669;
	wire [4-1:0] node47670;
	wire [4-1:0] node47672;
	wire [4-1:0] node47675;
	wire [4-1:0] node47676;
	wire [4-1:0] node47680;
	wire [4-1:0] node47681;
	wire [4-1:0] node47682;
	wire [4-1:0] node47683;
	wire [4-1:0] node47684;
	wire [4-1:0] node47685;
	wire [4-1:0] node47686;
	wire [4-1:0] node47690;
	wire [4-1:0] node47691;
	wire [4-1:0] node47695;
	wire [4-1:0] node47696;
	wire [4-1:0] node47698;
	wire [4-1:0] node47701;
	wire [4-1:0] node47703;
	wire [4-1:0] node47706;
	wire [4-1:0] node47707;
	wire [4-1:0] node47708;
	wire [4-1:0] node47709;
	wire [4-1:0] node47712;
	wire [4-1:0] node47715;
	wire [4-1:0] node47716;
	wire [4-1:0] node47719;
	wire [4-1:0] node47722;
	wire [4-1:0] node47723;
	wire [4-1:0] node47724;
	wire [4-1:0] node47727;
	wire [4-1:0] node47730;
	wire [4-1:0] node47732;
	wire [4-1:0] node47735;
	wire [4-1:0] node47736;
	wire [4-1:0] node47737;
	wire [4-1:0] node47739;
	wire [4-1:0] node47742;
	wire [4-1:0] node47743;
	wire [4-1:0] node47747;
	wire [4-1:0] node47748;
	wire [4-1:0] node47749;
	wire [4-1:0] node47753;
	wire [4-1:0] node47755;
	wire [4-1:0] node47758;
	wire [4-1:0] node47759;
	wire [4-1:0] node47760;
	wire [4-1:0] node47761;
	wire [4-1:0] node47762;
	wire [4-1:0] node47763;
	wire [4-1:0] node47764;
	wire [4-1:0] node47767;
	wire [4-1:0] node47770;
	wire [4-1:0] node47771;
	wire [4-1:0] node47774;
	wire [4-1:0] node47777;
	wire [4-1:0] node47778;
	wire [4-1:0] node47779;
	wire [4-1:0] node47783;
	wire [4-1:0] node47784;
	wire [4-1:0] node47787;
	wire [4-1:0] node47790;
	wire [4-1:0] node47791;
	wire [4-1:0] node47792;
	wire [4-1:0] node47795;
	wire [4-1:0] node47798;
	wire [4-1:0] node47800;
	wire [4-1:0] node47803;
	wire [4-1:0] node47804;
	wire [4-1:0] node47805;
	wire [4-1:0] node47806;
	wire [4-1:0] node47807;
	wire [4-1:0] node47810;
	wire [4-1:0] node47813;
	wire [4-1:0] node47814;
	wire [4-1:0] node47817;
	wire [4-1:0] node47820;
	wire [4-1:0] node47821;
	wire [4-1:0] node47823;
	wire [4-1:0] node47826;
	wire [4-1:0] node47829;
	wire [4-1:0] node47830;
	wire [4-1:0] node47831;
	wire [4-1:0] node47832;
	wire [4-1:0] node47835;
	wire [4-1:0] node47838;
	wire [4-1:0] node47839;
	wire [4-1:0] node47842;
	wire [4-1:0] node47845;
	wire [4-1:0] node47846;
	wire [4-1:0] node47847;
	wire [4-1:0] node47850;
	wire [4-1:0] node47853;
	wire [4-1:0] node47854;
	wire [4-1:0] node47857;
	wire [4-1:0] node47860;
	wire [4-1:0] node47861;
	wire [4-1:0] node47862;
	wire [4-1:0] node47863;
	wire [4-1:0] node47864;
	wire [4-1:0] node47865;
	wire [4-1:0] node47868;
	wire [4-1:0] node47871;
	wire [4-1:0] node47872;
	wire [4-1:0] node47875;
	wire [4-1:0] node47878;
	wire [4-1:0] node47880;
	wire [4-1:0] node47881;
	wire [4-1:0] node47884;
	wire [4-1:0] node47887;
	wire [4-1:0] node47888;
	wire [4-1:0] node47890;
	wire [4-1:0] node47891;
	wire [4-1:0] node47894;
	wire [4-1:0] node47897;
	wire [4-1:0] node47898;
	wire [4-1:0] node47899;
	wire [4-1:0] node47902;
	wire [4-1:0] node47905;
	wire [4-1:0] node47906;
	wire [4-1:0] node47910;
	wire [4-1:0] node47911;
	wire [4-1:0] node47912;
	wire [4-1:0] node47913;
	wire [4-1:0] node47916;
	wire [4-1:0] node47919;
	wire [4-1:0] node47920;
	wire [4-1:0] node47923;
	wire [4-1:0] node47926;
	wire [4-1:0] node47927;
	wire [4-1:0] node47928;
	wire [4-1:0] node47929;
	wire [4-1:0] node47932;
	wire [4-1:0] node47935;
	wire [4-1:0] node47936;
	wire [4-1:0] node47939;
	wire [4-1:0] node47942;
	wire [4-1:0] node47943;
	wire [4-1:0] node47944;
	wire [4-1:0] node47947;
	wire [4-1:0] node47950;
	wire [4-1:0] node47951;
	wire [4-1:0] node47954;
	wire [4-1:0] node47957;
	wire [4-1:0] node47958;
	wire [4-1:0] node47959;
	wire [4-1:0] node47960;
	wire [4-1:0] node47961;
	wire [4-1:0] node47962;
	wire [4-1:0] node47963;
	wire [4-1:0] node47966;
	wire [4-1:0] node47969;
	wire [4-1:0] node47970;
	wire [4-1:0] node47971;
	wire [4-1:0] node47974;
	wire [4-1:0] node47977;
	wire [4-1:0] node47978;
	wire [4-1:0] node47981;
	wire [4-1:0] node47984;
	wire [4-1:0] node47985;
	wire [4-1:0] node47986;
	wire [4-1:0] node47987;
	wire [4-1:0] node47990;
	wire [4-1:0] node47993;
	wire [4-1:0] node47994;
	wire [4-1:0] node47997;
	wire [4-1:0] node48000;
	wire [4-1:0] node48001;
	wire [4-1:0] node48002;
	wire [4-1:0] node48003;
	wire [4-1:0] node48006;
	wire [4-1:0] node48009;
	wire [4-1:0] node48011;
	wire [4-1:0] node48014;
	wire [4-1:0] node48015;
	wire [4-1:0] node48018;
	wire [4-1:0] node48021;
	wire [4-1:0] node48022;
	wire [4-1:0] node48023;
	wire [4-1:0] node48024;
	wire [4-1:0] node48025;
	wire [4-1:0] node48028;
	wire [4-1:0] node48031;
	wire [4-1:0] node48032;
	wire [4-1:0] node48035;
	wire [4-1:0] node48038;
	wire [4-1:0] node48039;
	wire [4-1:0] node48040;
	wire [4-1:0] node48041;
	wire [4-1:0] node48045;
	wire [4-1:0] node48047;
	wire [4-1:0] node48050;
	wire [4-1:0] node48051;
	wire [4-1:0] node48054;
	wire [4-1:0] node48057;
	wire [4-1:0] node48058;
	wire [4-1:0] node48061;
	wire [4-1:0] node48064;
	wire [4-1:0] node48065;
	wire [4-1:0] node48066;
	wire [4-1:0] node48067;
	wire [4-1:0] node48070;
	wire [4-1:0] node48073;
	wire [4-1:0] node48074;
	wire [4-1:0] node48077;
	wire [4-1:0] node48080;
	wire [4-1:0] node48081;
	wire [4-1:0] node48082;
	wire [4-1:0] node48083;
	wire [4-1:0] node48086;
	wire [4-1:0] node48089;
	wire [4-1:0] node48090;
	wire [4-1:0] node48093;
	wire [4-1:0] node48096;
	wire [4-1:0] node48097;
	wire [4-1:0] node48098;
	wire [4-1:0] node48100;
	wire [4-1:0] node48101;
	wire [4-1:0] node48104;
	wire [4-1:0] node48107;
	wire [4-1:0] node48108;
	wire [4-1:0] node48109;
	wire [4-1:0] node48112;
	wire [4-1:0] node48115;
	wire [4-1:0] node48116;
	wire [4-1:0] node48119;
	wire [4-1:0] node48122;
	wire [4-1:0] node48123;
	wire [4-1:0] node48124;
	wire [4-1:0] node48127;
	wire [4-1:0] node48130;
	wire [4-1:0] node48131;
	wire [4-1:0] node48133;
	wire [4-1:0] node48136;
	wire [4-1:0] node48137;
	wire [4-1:0] node48140;
	wire [4-1:0] node48143;
	wire [4-1:0] node48144;
	wire [4-1:0] node48145;
	wire [4-1:0] node48146;
	wire [4-1:0] node48147;
	wire [4-1:0] node48148;
	wire [4-1:0] node48151;
	wire [4-1:0] node48154;
	wire [4-1:0] node48157;
	wire [4-1:0] node48158;
	wire [4-1:0] node48159;
	wire [4-1:0] node48160;
	wire [4-1:0] node48163;
	wire [4-1:0] node48166;
	wire [4-1:0] node48167;
	wire [4-1:0] node48170;
	wire [4-1:0] node48173;
	wire [4-1:0] node48174;
	wire [4-1:0] node48177;
	wire [4-1:0] node48180;
	wire [4-1:0] node48181;
	wire [4-1:0] node48182;
	wire [4-1:0] node48183;
	wire [4-1:0] node48186;
	wire [4-1:0] node48189;
	wire [4-1:0] node48192;
	wire [4-1:0] node48193;
	wire [4-1:0] node48194;
	wire [4-1:0] node48195;
	wire [4-1:0] node48198;
	wire [4-1:0] node48201;
	wire [4-1:0] node48202;
	wire [4-1:0] node48205;
	wire [4-1:0] node48208;
	wire [4-1:0] node48209;
	wire [4-1:0] node48212;
	wire [4-1:0] node48215;
	wire [4-1:0] node48216;
	wire [4-1:0] node48217;
	wire [4-1:0] node48218;
	wire [4-1:0] node48219;
	wire [4-1:0] node48222;
	wire [4-1:0] node48225;
	wire [4-1:0] node48226;
	wire [4-1:0] node48229;
	wire [4-1:0] node48232;
	wire [4-1:0] node48233;
	wire [4-1:0] node48236;
	wire [4-1:0] node48239;
	wire [4-1:0] node48240;
	wire [4-1:0] node48241;
	wire [4-1:0] node48242;
	wire [4-1:0] node48243;
	wire [4-1:0] node48244;
	wire [4-1:0] node48248;
	wire [4-1:0] node48249;
	wire [4-1:0] node48252;
	wire [4-1:0] node48255;
	wire [4-1:0] node48256;
	wire [4-1:0] node48259;
	wire [4-1:0] node48262;
	wire [4-1:0] node48263;
	wire [4-1:0] node48264;
	wire [4-1:0] node48265;
	wire [4-1:0] node48268;
	wire [4-1:0] node48271;
	wire [4-1:0] node48272;
	wire [4-1:0] node48276;
	wire [4-1:0] node48277;
	wire [4-1:0] node48278;
	wire [4-1:0] node48281;
	wire [4-1:0] node48284;
	wire [4-1:0] node48285;
	wire [4-1:0] node48288;
	wire [4-1:0] node48291;
	wire [4-1:0] node48292;
	wire [4-1:0] node48295;
	wire [4-1:0] node48298;
	wire [4-1:0] node48299;
	wire [4-1:0] node48300;
	wire [4-1:0] node48301;
	wire [4-1:0] node48302;
	wire [4-1:0] node48303;
	wire [4-1:0] node48304;
	wire [4-1:0] node48305;
	wire [4-1:0] node48306;
	wire [4-1:0] node48307;
	wire [4-1:0] node48310;
	wire [4-1:0] node48313;
	wire [4-1:0] node48314;
	wire [4-1:0] node48317;
	wire [4-1:0] node48320;
	wire [4-1:0] node48322;
	wire [4-1:0] node48323;
	wire [4-1:0] node48327;
	wire [4-1:0] node48328;
	wire [4-1:0] node48329;
	wire [4-1:0] node48330;
	wire [4-1:0] node48333;
	wire [4-1:0] node48336;
	wire [4-1:0] node48338;
	wire [4-1:0] node48341;
	wire [4-1:0] node48342;
	wire [4-1:0] node48343;
	wire [4-1:0] node48346;
	wire [4-1:0] node48349;
	wire [4-1:0] node48350;
	wire [4-1:0] node48353;
	wire [4-1:0] node48356;
	wire [4-1:0] node48357;
	wire [4-1:0] node48358;
	wire [4-1:0] node48359;
	wire [4-1:0] node48360;
	wire [4-1:0] node48363;
	wire [4-1:0] node48366;
	wire [4-1:0] node48367;
	wire [4-1:0] node48370;
	wire [4-1:0] node48373;
	wire [4-1:0] node48374;
	wire [4-1:0] node48377;
	wire [4-1:0] node48380;
	wire [4-1:0] node48381;
	wire [4-1:0] node48382;
	wire [4-1:0] node48383;
	wire [4-1:0] node48386;
	wire [4-1:0] node48389;
	wire [4-1:0] node48390;
	wire [4-1:0] node48393;
	wire [4-1:0] node48396;
	wire [4-1:0] node48397;
	wire [4-1:0] node48399;
	wire [4-1:0] node48402;
	wire [4-1:0] node48404;
	wire [4-1:0] node48407;
	wire [4-1:0] node48408;
	wire [4-1:0] node48409;
	wire [4-1:0] node48412;
	wire [4-1:0] node48415;
	wire [4-1:0] node48416;
	wire [4-1:0] node48417;
	wire [4-1:0] node48418;
	wire [4-1:0] node48421;
	wire [4-1:0] node48424;
	wire [4-1:0] node48425;
	wire [4-1:0] node48426;
	wire [4-1:0] node48429;
	wire [4-1:0] node48432;
	wire [4-1:0] node48433;
	wire [4-1:0] node48436;
	wire [4-1:0] node48439;
	wire [4-1:0] node48440;
	wire [4-1:0] node48443;
	wire [4-1:0] node48446;
	wire [4-1:0] node48447;
	wire [4-1:0] node48448;
	wire [4-1:0] node48449;
	wire [4-1:0] node48450;
	wire [4-1:0] node48454;
	wire [4-1:0] node48455;
	wire [4-1:0] node48459;
	wire [4-1:0] node48460;
	wire [4-1:0] node48461;
	wire [4-1:0] node48465;
	wire [4-1:0] node48466;
	wire [4-1:0] node48470;
	wire [4-1:0] node48471;
	wire [4-1:0] node48472;
	wire [4-1:0] node48473;
	wire [4-1:0] node48477;
	wire [4-1:0] node48478;
	wire [4-1:0] node48482;
	wire [4-1:0] node48483;
	wire [4-1:0] node48484;
	wire [4-1:0] node48488;
	wire [4-1:0] node48489;
	wire [4-1:0] node48493;
	wire [4-1:0] node48494;
	wire [4-1:0] node48495;
	wire [4-1:0] node48496;
	wire [4-1:0] node48497;
	wire [4-1:0] node48498;
	wire [4-1:0] node48499;
	wire [4-1:0] node48502;
	wire [4-1:0] node48505;
	wire [4-1:0] node48506;
	wire [4-1:0] node48509;
	wire [4-1:0] node48512;
	wire [4-1:0] node48513;
	wire [4-1:0] node48516;
	wire [4-1:0] node48519;
	wire [4-1:0] node48520;
	wire [4-1:0] node48523;
	wire [4-1:0] node48526;
	wire [4-1:0] node48527;
	wire [4-1:0] node48530;
	wire [4-1:0] node48533;
	wire [4-1:0] node48534;
	wire [4-1:0] node48535;
	wire [4-1:0] node48536;
	wire [4-1:0] node48537;
	wire [4-1:0] node48540;
	wire [4-1:0] node48543;
	wire [4-1:0] node48544;
	wire [4-1:0] node48547;
	wire [4-1:0] node48550;
	wire [4-1:0] node48551;
	wire [4-1:0] node48552;
	wire [4-1:0] node48555;
	wire [4-1:0] node48558;
	wire [4-1:0] node48559;
	wire [4-1:0] node48562;
	wire [4-1:0] node48565;
	wire [4-1:0] node48566;
	wire [4-1:0] node48567;
	wire [4-1:0] node48570;
	wire [4-1:0] node48573;
	wire [4-1:0] node48574;
	wire [4-1:0] node48575;
	wire [4-1:0] node48576;
	wire [4-1:0] node48579;
	wire [4-1:0] node48582;
	wire [4-1:0] node48583;
	wire [4-1:0] node48587;
	wire [4-1:0] node48588;
	wire [4-1:0] node48591;
	wire [4-1:0] node48594;
	wire [4-1:0] node48595;
	wire [4-1:0] node48596;
	wire [4-1:0] node48597;
	wire [4-1:0] node48598;
	wire [4-1:0] node48599;
	wire [4-1:0] node48600;
	wire [4-1:0] node48601;
	wire [4-1:0] node48603;
	wire [4-1:0] node48606;
	wire [4-1:0] node48609;
	wire [4-1:0] node48610;
	wire [4-1:0] node48611;
	wire [4-1:0] node48615;
	wire [4-1:0] node48616;
	wire [4-1:0] node48620;
	wire [4-1:0] node48621;
	wire [4-1:0] node48622;
	wire [4-1:0] node48625;
	wire [4-1:0] node48626;
	wire [4-1:0] node48630;
	wire [4-1:0] node48631;
	wire [4-1:0] node48632;
	wire [4-1:0] node48636;
	wire [4-1:0] node48639;
	wire [4-1:0] node48640;
	wire [4-1:0] node48641;
	wire [4-1:0] node48644;
	wire [4-1:0] node48647;
	wire [4-1:0] node48648;
	wire [4-1:0] node48649;
	wire [4-1:0] node48652;
	wire [4-1:0] node48655;
	wire [4-1:0] node48656;
	wire [4-1:0] node48657;
	wire [4-1:0] node48661;
	wire [4-1:0] node48663;
	wire [4-1:0] node48666;
	wire [4-1:0] node48667;
	wire [4-1:0] node48668;
	wire [4-1:0] node48669;
	wire [4-1:0] node48670;
	wire [4-1:0] node48673;
	wire [4-1:0] node48676;
	wire [4-1:0] node48677;
	wire [4-1:0] node48680;
	wire [4-1:0] node48683;
	wire [4-1:0] node48684;
	wire [4-1:0] node48685;
	wire [4-1:0] node48688;
	wire [4-1:0] node48691;
	wire [4-1:0] node48693;
	wire [4-1:0] node48696;
	wire [4-1:0] node48697;
	wire [4-1:0] node48698;
	wire [4-1:0] node48699;
	wire [4-1:0] node48702;
	wire [4-1:0] node48705;
	wire [4-1:0] node48706;
	wire [4-1:0] node48707;
	wire [4-1:0] node48711;
	wire [4-1:0] node48712;
	wire [4-1:0] node48715;
	wire [4-1:0] node48718;
	wire [4-1:0] node48719;
	wire [4-1:0] node48720;
	wire [4-1:0] node48721;
	wire [4-1:0] node48724;
	wire [4-1:0] node48728;
	wire [4-1:0] node48730;
	wire [4-1:0] node48731;
	wire [4-1:0] node48734;
	wire [4-1:0] node48737;
	wire [4-1:0] node48738;
	wire [4-1:0] node48739;
	wire [4-1:0] node48740;
	wire [4-1:0] node48741;
	wire [4-1:0] node48745;
	wire [4-1:0] node48748;
	wire [4-1:0] node48749;
	wire [4-1:0] node48751;
	wire [4-1:0] node48754;
	wire [4-1:0] node48755;
	wire [4-1:0] node48756;
	wire [4-1:0] node48758;
	wire [4-1:0] node48761;
	wire [4-1:0] node48762;
	wire [4-1:0] node48765;
	wire [4-1:0] node48768;
	wire [4-1:0] node48769;
	wire [4-1:0] node48772;
	wire [4-1:0] node48775;
	wire [4-1:0] node48776;
	wire [4-1:0] node48777;
	wire [4-1:0] node48778;
	wire [4-1:0] node48783;
	wire [4-1:0] node48784;
	wire [4-1:0] node48785;
	wire [4-1:0] node48790;
	wire [4-1:0] node48791;
	wire [4-1:0] node48792;
	wire [4-1:0] node48793;
	wire [4-1:0] node48794;
	wire [4-1:0] node48796;
	wire [4-1:0] node48799;
	wire [4-1:0] node48800;
	wire [4-1:0] node48803;
	wire [4-1:0] node48806;
	wire [4-1:0] node48807;
	wire [4-1:0] node48808;
	wire [4-1:0] node48812;
	wire [4-1:0] node48815;
	wire [4-1:0] node48816;
	wire [4-1:0] node48817;
	wire [4-1:0] node48818;
	wire [4-1:0] node48823;
	wire [4-1:0] node48824;
	wire [4-1:0] node48825;
	wire [4-1:0] node48830;
	wire [4-1:0] node48831;
	wire [4-1:0] node48832;
	wire [4-1:0] node48833;
	wire [4-1:0] node48834;
	wire [4-1:0] node48836;
	wire [4-1:0] node48839;
	wire [4-1:0] node48840;
	wire [4-1:0] node48844;
	wire [4-1:0] node48845;
	wire [4-1:0] node48847;
	wire [4-1:0] node48850;
	wire [4-1:0] node48851;
	wire [4-1:0] node48855;
	wire [4-1:0] node48856;
	wire [4-1:0] node48857;
	wire [4-1:0] node48858;
	wire [4-1:0] node48862;
	wire [4-1:0] node48864;
	wire [4-1:0] node48867;
	wire [4-1:0] node48868;
	wire [4-1:0] node48870;
	wire [4-1:0] node48873;
	wire [4-1:0] node48875;
	wire [4-1:0] node48878;
	wire [4-1:0] node48879;
	wire [4-1:0] node48880;
	wire [4-1:0] node48881;
	wire [4-1:0] node48882;
	wire [4-1:0] node48885;
	wire [4-1:0] node48888;
	wire [4-1:0] node48889;
	wire [4-1:0] node48892;
	wire [4-1:0] node48895;
	wire [4-1:0] node48896;
	wire [4-1:0] node48899;
	wire [4-1:0] node48902;
	wire [4-1:0] node48903;
	wire [4-1:0] node48906;
	wire [4-1:0] node48909;
	wire [4-1:0] node48910;
	wire [4-1:0] node48911;
	wire [4-1:0] node48912;
	wire [4-1:0] node48913;
	wire [4-1:0] node48914;
	wire [4-1:0] node48915;
	wire [4-1:0] node48916;
	wire [4-1:0] node48917;
	wire [4-1:0] node48918;
	wire [4-1:0] node48919;
	wire [4-1:0] node48923;
	wire [4-1:0] node48924;
	wire [4-1:0] node48927;
	wire [4-1:0] node48929;
	wire [4-1:0] node48932;
	wire [4-1:0] node48933;
	wire [4-1:0] node48935;
	wire [4-1:0] node48938;
	wire [4-1:0] node48939;
	wire [4-1:0] node48940;
	wire [4-1:0] node48944;
	wire [4-1:0] node48945;
	wire [4-1:0] node48948;
	wire [4-1:0] node48951;
	wire [4-1:0] node48952;
	wire [4-1:0] node48953;
	wire [4-1:0] node48956;
	wire [4-1:0] node48957;
	wire [4-1:0] node48959;
	wire [4-1:0] node48963;
	wire [4-1:0] node48964;
	wire [4-1:0] node48966;
	wire [4-1:0] node48967;
	wire [4-1:0] node48971;
	wire [4-1:0] node48972;
	wire [4-1:0] node48976;
	wire [4-1:0] node48977;
	wire [4-1:0] node48978;
	wire [4-1:0] node48979;
	wire [4-1:0] node48980;
	wire [4-1:0] node48983;
	wire [4-1:0] node48984;
	wire [4-1:0] node48987;
	wire [4-1:0] node48990;
	wire [4-1:0] node48991;
	wire [4-1:0] node48992;
	wire [4-1:0] node48995;
	wire [4-1:0] node48998;
	wire [4-1:0] node48999;
	wire [4-1:0] node49003;
	wire [4-1:0] node49004;
	wire [4-1:0] node49005;
	wire [4-1:0] node49007;
	wire [4-1:0] node49010;
	wire [4-1:0] node49012;
	wire [4-1:0] node49015;
	wire [4-1:0] node49016;
	wire [4-1:0] node49018;
	wire [4-1:0] node49021;
	wire [4-1:0] node49022;
	wire [4-1:0] node49026;
	wire [4-1:0] node49027;
	wire [4-1:0] node49028;
	wire [4-1:0] node49029;
	wire [4-1:0] node49032;
	wire [4-1:0] node49035;
	wire [4-1:0] node49036;
	wire [4-1:0] node49037;
	wire [4-1:0] node49041;
	wire [4-1:0] node49042;
	wire [4-1:0] node49045;
	wire [4-1:0] node49048;
	wire [4-1:0] node49049;
	wire [4-1:0] node49050;
	wire [4-1:0] node49052;
	wire [4-1:0] node49056;
	wire [4-1:0] node49057;
	wire [4-1:0] node49061;
	wire [4-1:0] node49062;
	wire [4-1:0] node49063;
	wire [4-1:0] node49064;
	wire [4-1:0] node49065;
	wire [4-1:0] node49067;
	wire [4-1:0] node49070;
	wire [4-1:0] node49071;
	wire [4-1:0] node49072;
	wire [4-1:0] node49076;
	wire [4-1:0] node49079;
	wire [4-1:0] node49080;
	wire [4-1:0] node49081;
	wire [4-1:0] node49085;
	wire [4-1:0] node49087;
	wire [4-1:0] node49089;
	wire [4-1:0] node49092;
	wire [4-1:0] node49093;
	wire [4-1:0] node49094;
	wire [4-1:0] node49095;
	wire [4-1:0] node49096;
	wire [4-1:0] node49100;
	wire [4-1:0] node49101;
	wire [4-1:0] node49105;
	wire [4-1:0] node49106;
	wire [4-1:0] node49107;
	wire [4-1:0] node49111;
	wire [4-1:0] node49114;
	wire [4-1:0] node49115;
	wire [4-1:0] node49116;
	wire [4-1:0] node49118;
	wire [4-1:0] node49121;
	wire [4-1:0] node49123;
	wire [4-1:0] node49126;
	wire [4-1:0] node49127;
	wire [4-1:0] node49128;
	wire [4-1:0] node49132;
	wire [4-1:0] node49133;
	wire [4-1:0] node49137;
	wire [4-1:0] node49138;
	wire [4-1:0] node49139;
	wire [4-1:0] node49140;
	wire [4-1:0] node49142;
	wire [4-1:0] node49145;
	wire [4-1:0] node49147;
	wire [4-1:0] node49150;
	wire [4-1:0] node49151;
	wire [4-1:0] node49152;
	wire [4-1:0] node49153;
	wire [4-1:0] node49156;
	wire [4-1:0] node49159;
	wire [4-1:0] node49161;
	wire [4-1:0] node49164;
	wire [4-1:0] node49165;
	wire [4-1:0] node49169;
	wire [4-1:0] node49170;
	wire [4-1:0] node49171;
	wire [4-1:0] node49172;
	wire [4-1:0] node49173;
	wire [4-1:0] node49176;
	wire [4-1:0] node49179;
	wire [4-1:0] node49180;
	wire [4-1:0] node49183;
	wire [4-1:0] node49186;
	wire [4-1:0] node49187;
	wire [4-1:0] node49190;
	wire [4-1:0] node49191;
	wire [4-1:0] node49195;
	wire [4-1:0] node49196;
	wire [4-1:0] node49197;
	wire [4-1:0] node49198;
	wire [4-1:0] node49202;
	wire [4-1:0] node49203;
	wire [4-1:0] node49206;
	wire [4-1:0] node49209;
	wire [4-1:0] node49212;
	wire [4-1:0] node49213;
	wire [4-1:0] node49214;
	wire [4-1:0] node49215;
	wire [4-1:0] node49216;
	wire [4-1:0] node49217;
	wire [4-1:0] node49220;
	wire [4-1:0] node49221;
	wire [4-1:0] node49223;
	wire [4-1:0] node49226;
	wire [4-1:0] node49229;
	wire [4-1:0] node49230;
	wire [4-1:0] node49231;
	wire [4-1:0] node49234;
	wire [4-1:0] node49236;
	wire [4-1:0] node49239;
	wire [4-1:0] node49240;
	wire [4-1:0] node49243;
	wire [4-1:0] node49246;
	wire [4-1:0] node49247;
	wire [4-1:0] node49248;
	wire [4-1:0] node49249;
	wire [4-1:0] node49250;
	wire [4-1:0] node49253;
	wire [4-1:0] node49256;
	wire [4-1:0] node49257;
	wire [4-1:0] node49261;
	wire [4-1:0] node49262;
	wire [4-1:0] node49263;
	wire [4-1:0] node49266;
	wire [4-1:0] node49269;
	wire [4-1:0] node49270;
	wire [4-1:0] node49274;
	wire [4-1:0] node49275;
	wire [4-1:0] node49276;
	wire [4-1:0] node49279;
	wire [4-1:0] node49280;
	wire [4-1:0] node49283;
	wire [4-1:0] node49286;
	wire [4-1:0] node49287;
	wire [4-1:0] node49289;
	wire [4-1:0] node49292;
	wire [4-1:0] node49295;
	wire [4-1:0] node49296;
	wire [4-1:0] node49297;
	wire [4-1:0] node49298;
	wire [4-1:0] node49301;
	wire [4-1:0] node49302;
	wire [4-1:0] node49304;
	wire [4-1:0] node49307;
	wire [4-1:0] node49310;
	wire [4-1:0] node49311;
	wire [4-1:0] node49312;
	wire [4-1:0] node49315;
	wire [4-1:0] node49317;
	wire [4-1:0] node49320;
	wire [4-1:0] node49321;
	wire [4-1:0] node49322;
	wire [4-1:0] node49326;
	wire [4-1:0] node49328;
	wire [4-1:0] node49331;
	wire [4-1:0] node49332;
	wire [4-1:0] node49333;
	wire [4-1:0] node49334;
	wire [4-1:0] node49336;
	wire [4-1:0] node49339;
	wire [4-1:0] node49342;
	wire [4-1:0] node49343;
	wire [4-1:0] node49345;
	wire [4-1:0] node49348;
	wire [4-1:0] node49349;
	wire [4-1:0] node49353;
	wire [4-1:0] node49354;
	wire [4-1:0] node49355;
	wire [4-1:0] node49358;
	wire [4-1:0] node49359;
	wire [4-1:0] node49362;
	wire [4-1:0] node49365;
	wire [4-1:0] node49366;
	wire [4-1:0] node49367;
	wire [4-1:0] node49370;
	wire [4-1:0] node49373;
	wire [4-1:0] node49376;
	wire [4-1:0] node49377;
	wire [4-1:0] node49378;
	wire [4-1:0] node49379;
	wire [4-1:0] node49380;
	wire [4-1:0] node49381;
	wire [4-1:0] node49383;
	wire [4-1:0] node49386;
	wire [4-1:0] node49387;
	wire [4-1:0] node49390;
	wire [4-1:0] node49393;
	wire [4-1:0] node49394;
	wire [4-1:0] node49395;
	wire [4-1:0] node49398;
	wire [4-1:0] node49401;
	wire [4-1:0] node49404;
	wire [4-1:0] node49405;
	wire [4-1:0] node49406;
	wire [4-1:0] node49407;
	wire [4-1:0] node49410;
	wire [4-1:0] node49414;
	wire [4-1:0] node49415;
	wire [4-1:0] node49417;
	wire [4-1:0] node49420;
	wire [4-1:0] node49421;
	wire [4-1:0] node49425;
	wire [4-1:0] node49426;
	wire [4-1:0] node49427;
	wire [4-1:0] node49428;
	wire [4-1:0] node49432;
	wire [4-1:0] node49434;
	wire [4-1:0] node49435;
	wire [4-1:0] node49439;
	wire [4-1:0] node49440;
	wire [4-1:0] node49441;
	wire [4-1:0] node49442;
	wire [4-1:0] node49446;
	wire [4-1:0] node49448;
	wire [4-1:0] node49451;
	wire [4-1:0] node49452;
	wire [4-1:0] node49456;
	wire [4-1:0] node49457;
	wire [4-1:0] node49458;
	wire [4-1:0] node49459;
	wire [4-1:0] node49460;
	wire [4-1:0] node49463;
	wire [4-1:0] node49464;
	wire [4-1:0] node49467;
	wire [4-1:0] node49470;
	wire [4-1:0] node49471;
	wire [4-1:0] node49472;
	wire [4-1:0] node49475;
	wire [4-1:0] node49478;
	wire [4-1:0] node49480;
	wire [4-1:0] node49483;
	wire [4-1:0] node49484;
	wire [4-1:0] node49487;
	wire [4-1:0] node49488;
	wire [4-1:0] node49489;
	wire [4-1:0] node49492;
	wire [4-1:0] node49496;
	wire [4-1:0] node49497;
	wire [4-1:0] node49498;
	wire [4-1:0] node49499;
	wire [4-1:0] node49501;
	wire [4-1:0] node49504;
	wire [4-1:0] node49507;
	wire [4-1:0] node49509;
	wire [4-1:0] node49510;
	wire [4-1:0] node49513;
	wire [4-1:0] node49516;
	wire [4-1:0] node49517;
	wire [4-1:0] node49518;
	wire [4-1:0] node49519;
	wire [4-1:0] node49523;
	wire [4-1:0] node49525;
	wire [4-1:0] node49528;
	wire [4-1:0] node49529;
	wire [4-1:0] node49530;
	wire [4-1:0] node49534;
	wire [4-1:0] node49535;
	wire [4-1:0] node49539;
	wire [4-1:0] node49540;
	wire [4-1:0] node49541;
	wire [4-1:0] node49542;
	wire [4-1:0] node49543;
	wire [4-1:0] node49544;
	wire [4-1:0] node49545;
	wire [4-1:0] node49546;
	wire [4-1:0] node49549;
	wire [4-1:0] node49552;
	wire [4-1:0] node49554;
	wire [4-1:0] node49557;
	wire [4-1:0] node49558;
	wire [4-1:0] node49559;
	wire [4-1:0] node49562;
	wire [4-1:0] node49565;
	wire [4-1:0] node49566;
	wire [4-1:0] node49570;
	wire [4-1:0] node49571;
	wire [4-1:0] node49572;
	wire [4-1:0] node49573;
	wire [4-1:0] node49576;
	wire [4-1:0] node49579;
	wire [4-1:0] node49580;
	wire [4-1:0] node49583;
	wire [4-1:0] node49586;
	wire [4-1:0] node49587;
	wire [4-1:0] node49588;
	wire [4-1:0] node49592;
	wire [4-1:0] node49593;
	wire [4-1:0] node49596;
	wire [4-1:0] node49599;
	wire [4-1:0] node49600;
	wire [4-1:0] node49601;
	wire [4-1:0] node49602;
	wire [4-1:0] node49605;
	wire [4-1:0] node49608;
	wire [4-1:0] node49609;
	wire [4-1:0] node49610;
	wire [4-1:0] node49614;
	wire [4-1:0] node49615;
	wire [4-1:0] node49618;
	wire [4-1:0] node49621;
	wire [4-1:0] node49622;
	wire [4-1:0] node49624;
	wire [4-1:0] node49625;
	wire [4-1:0] node49629;
	wire [4-1:0] node49630;
	wire [4-1:0] node49634;
	wire [4-1:0] node49635;
	wire [4-1:0] node49636;
	wire [4-1:0] node49637;
	wire [4-1:0] node49639;
	wire [4-1:0] node49642;
	wire [4-1:0] node49644;
	wire [4-1:0] node49645;
	wire [4-1:0] node49649;
	wire [4-1:0] node49650;
	wire [4-1:0] node49651;
	wire [4-1:0] node49652;
	wire [4-1:0] node49655;
	wire [4-1:0] node49658;
	wire [4-1:0] node49660;
	wire [4-1:0] node49663;
	wire [4-1:0] node49664;
	wire [4-1:0] node49667;
	wire [4-1:0] node49670;
	wire [4-1:0] node49671;
	wire [4-1:0] node49672;
	wire [4-1:0] node49673;
	wire [4-1:0] node49675;
	wire [4-1:0] node49678;
	wire [4-1:0] node49680;
	wire [4-1:0] node49683;
	wire [4-1:0] node49684;
	wire [4-1:0] node49685;
	wire [4-1:0] node49688;
	wire [4-1:0] node49691;
	wire [4-1:0] node49692;
	wire [4-1:0] node49696;
	wire [4-1:0] node49697;
	wire [4-1:0] node49698;
	wire [4-1:0] node49701;
	wire [4-1:0] node49702;
	wire [4-1:0] node49705;
	wire [4-1:0] node49708;
	wire [4-1:0] node49709;
	wire [4-1:0] node49710;
	wire [4-1:0] node49713;
	wire [4-1:0] node49716;
	wire [4-1:0] node49717;
	wire [4-1:0] node49720;
	wire [4-1:0] node49723;
	wire [4-1:0] node49724;
	wire [4-1:0] node49725;
	wire [4-1:0] node49726;
	wire [4-1:0] node49727;
	wire [4-1:0] node49729;
	wire [4-1:0] node49732;
	wire [4-1:0] node49733;
	wire [4-1:0] node49734;
	wire [4-1:0] node49738;
	wire [4-1:0] node49739;
	wire [4-1:0] node49742;
	wire [4-1:0] node49745;
	wire [4-1:0] node49746;
	wire [4-1:0] node49747;
	wire [4-1:0] node49749;
	wire [4-1:0] node49753;
	wire [4-1:0] node49754;
	wire [4-1:0] node49757;
	wire [4-1:0] node49760;
	wire [4-1:0] node49761;
	wire [4-1:0] node49762;
	wire [4-1:0] node49763;
	wire [4-1:0] node49765;
	wire [4-1:0] node49768;
	wire [4-1:0] node49769;
	wire [4-1:0] node49772;
	wire [4-1:0] node49775;
	wire [4-1:0] node49776;
	wire [4-1:0] node49778;
	wire [4-1:0] node49781;
	wire [4-1:0] node49782;
	wire [4-1:0] node49785;
	wire [4-1:0] node49788;
	wire [4-1:0] node49789;
	wire [4-1:0] node49790;
	wire [4-1:0] node49791;
	wire [4-1:0] node49794;
	wire [4-1:0] node49797;
	wire [4-1:0] node49798;
	wire [4-1:0] node49799;
	wire [4-1:0] node49802;
	wire [4-1:0] node49805;
	wire [4-1:0] node49806;
	wire [4-1:0] node49809;
	wire [4-1:0] node49812;
	wire [4-1:0] node49813;
	wire [4-1:0] node49814;
	wire [4-1:0] node49817;
	wire [4-1:0] node49820;
	wire [4-1:0] node49823;
	wire [4-1:0] node49824;
	wire [4-1:0] node49825;
	wire [4-1:0] node49826;
	wire [4-1:0] node49827;
	wire [4-1:0] node49828;
	wire [4-1:0] node49831;
	wire [4-1:0] node49834;
	wire [4-1:0] node49835;
	wire [4-1:0] node49838;
	wire [4-1:0] node49841;
	wire [4-1:0] node49842;
	wire [4-1:0] node49843;
	wire [4-1:0] node49846;
	wire [4-1:0] node49849;
	wire [4-1:0] node49852;
	wire [4-1:0] node49853;
	wire [4-1:0] node49854;
	wire [4-1:0] node49856;
	wire [4-1:0] node49859;
	wire [4-1:0] node49861;
	wire [4-1:0] node49864;
	wire [4-1:0] node49865;
	wire [4-1:0] node49866;
	wire [4-1:0] node49869;
	wire [4-1:0] node49872;
	wire [4-1:0] node49875;
	wire [4-1:0] node49876;
	wire [4-1:0] node49877;
	wire [4-1:0] node49879;
	wire [4-1:0] node49882;
	wire [4-1:0] node49884;
	wire [4-1:0] node49885;
	wire [4-1:0] node49889;
	wire [4-1:0] node49890;
	wire [4-1:0] node49891;
	wire [4-1:0] node49892;
	wire [4-1:0] node49895;
	wire [4-1:0] node49898;
	wire [4-1:0] node49900;
	wire [4-1:0] node49903;
	wire [4-1:0] node49904;
	wire [4-1:0] node49908;
	wire [4-1:0] node49909;
	wire [4-1:0] node49910;
	wire [4-1:0] node49911;
	wire [4-1:0] node49912;
	wire [4-1:0] node49913;
	wire [4-1:0] node49915;
	wire [4-1:0] node49918;
	wire [4-1:0] node49920;
	wire [4-1:0] node49923;
	wire [4-1:0] node49924;
	wire [4-1:0] node49926;
	wire [4-1:0] node49929;
	wire [4-1:0] node49931;
	wire [4-1:0] node49934;
	wire [4-1:0] node49935;
	wire [4-1:0] node49936;
	wire [4-1:0] node49938;
	wire [4-1:0] node49941;
	wire [4-1:0] node49943;
	wire [4-1:0] node49946;
	wire [4-1:0] node49947;
	wire [4-1:0] node49949;
	wire [4-1:0] node49952;
	wire [4-1:0] node49954;
	wire [4-1:0] node49957;
	wire [4-1:0] node49958;
	wire [4-1:0] node49961;
	wire [4-1:0] node49964;
	wire [4-1:0] node49965;
	wire [4-1:0] node49966;
	wire [4-1:0] node49967;
	wire [4-1:0] node49968;
	wire [4-1:0] node49971;
	wire [4-1:0] node49974;
	wire [4-1:0] node49975;
	wire [4-1:0] node49976;
	wire [4-1:0] node49977;
	wire [4-1:0] node49980;
	wire [4-1:0] node49983;
	wire [4-1:0] node49984;
	wire [4-1:0] node49987;
	wire [4-1:0] node49990;
	wire [4-1:0] node49991;
	wire [4-1:0] node49992;
	wire [4-1:0] node49993;
	wire [4-1:0] node49996;
	wire [4-1:0] node49999;
	wire [4-1:0] node50000;
	wire [4-1:0] node50003;
	wire [4-1:0] node50006;
	wire [4-1:0] node50007;
	wire [4-1:0] node50008;
	wire [4-1:0] node50011;
	wire [4-1:0] node50014;
	wire [4-1:0] node50015;
	wire [4-1:0] node50016;
	wire [4-1:0] node50019;
	wire [4-1:0] node50022;
	wire [4-1:0] node50023;
	wire [4-1:0] node50026;
	wire [4-1:0] node50029;
	wire [4-1:0] node50030;
	wire [4-1:0] node50031;
	wire [4-1:0] node50032;
	wire [4-1:0] node50033;
	wire [4-1:0] node50037;
	wire [4-1:0] node50038;
	wire [4-1:0] node50042;
	wire [4-1:0] node50043;
	wire [4-1:0] node50044;
	wire [4-1:0] node50048;
	wire [4-1:0] node50050;
	wire [4-1:0] node50053;
	wire [4-1:0] node50054;
	wire [4-1:0] node50055;
	wire [4-1:0] node50057;
	wire [4-1:0] node50060;
	wire [4-1:0] node50062;
	wire [4-1:0] node50065;
	wire [4-1:0] node50066;
	wire [4-1:0] node50067;
	wire [4-1:0] node50071;
	wire [4-1:0] node50072;
	wire [4-1:0] node50076;
	wire [4-1:0] node50077;
	wire [4-1:0] node50080;
	wire [4-1:0] node50083;
	wire [4-1:0] node50084;
	wire [4-1:0] node50085;
	wire [4-1:0] node50086;
	wire [4-1:0] node50087;
	wire [4-1:0] node50088;
	wire [4-1:0] node50089;
	wire [4-1:0] node50090;
	wire [4-1:0] node50091;
	wire [4-1:0] node50092;
	wire [4-1:0] node50093;
	wire [4-1:0] node50096;
	wire [4-1:0] node50100;
	wire [4-1:0] node50101;
	wire [4-1:0] node50102;
	wire [4-1:0] node50105;
	wire [4-1:0] node50108;
	wire [4-1:0] node50109;
	wire [4-1:0] node50113;
	wire [4-1:0] node50114;
	wire [4-1:0] node50115;
	wire [4-1:0] node50116;
	wire [4-1:0] node50119;
	wire [4-1:0] node50122;
	wire [4-1:0] node50124;
	wire [4-1:0] node50127;
	wire [4-1:0] node50128;
	wire [4-1:0] node50131;
	wire [4-1:0] node50134;
	wire [4-1:0] node50135;
	wire [4-1:0] node50136;
	wire [4-1:0] node50137;
	wire [4-1:0] node50138;
	wire [4-1:0] node50141;
	wire [4-1:0] node50144;
	wire [4-1:0] node50145;
	wire [4-1:0] node50149;
	wire [4-1:0] node50150;
	wire [4-1:0] node50151;
	wire [4-1:0] node50154;
	wire [4-1:0] node50157;
	wire [4-1:0] node50158;
	wire [4-1:0] node50161;
	wire [4-1:0] node50164;
	wire [4-1:0] node50165;
	wire [4-1:0] node50166;
	wire [4-1:0] node50170;
	wire [4-1:0] node50171;
	wire [4-1:0] node50172;
	wire [4-1:0] node50176;
	wire [4-1:0] node50177;
	wire [4-1:0] node50181;
	wire [4-1:0] node50182;
	wire [4-1:0] node50183;
	wire [4-1:0] node50185;
	wire [4-1:0] node50188;
	wire [4-1:0] node50190;
	wire [4-1:0] node50193;
	wire [4-1:0] node50194;
	wire [4-1:0] node50196;
	wire [4-1:0] node50199;
	wire [4-1:0] node50201;
	wire [4-1:0] node50204;
	wire [4-1:0] node50205;
	wire [4-1:0] node50206;
	wire [4-1:0] node50207;
	wire [4-1:0] node50208;
	wire [4-1:0] node50210;
	wire [4-1:0] node50213;
	wire [4-1:0] node50215;
	wire [4-1:0] node50218;
	wire [4-1:0] node50219;
	wire [4-1:0] node50221;
	wire [4-1:0] node50224;
	wire [4-1:0] node50227;
	wire [4-1:0] node50228;
	wire [4-1:0] node50229;
	wire [4-1:0] node50231;
	wire [4-1:0] node50234;
	wire [4-1:0] node50237;
	wire [4-1:0] node50238;
	wire [4-1:0] node50240;
	wire [4-1:0] node50243;
	wire [4-1:0] node50245;
	wire [4-1:0] node50248;
	wire [4-1:0] node50249;
	wire [4-1:0] node50250;
	wire [4-1:0] node50251;
	wire [4-1:0] node50254;
	wire [4-1:0] node50257;
	wire [4-1:0] node50258;
	wire [4-1:0] node50261;
	wire [4-1:0] node50264;
	wire [4-1:0] node50265;
	wire [4-1:0] node50266;
	wire [4-1:0] node50267;
	wire [4-1:0] node50268;
	wire [4-1:0] node50271;
	wire [4-1:0] node50274;
	wire [4-1:0] node50275;
	wire [4-1:0] node50279;
	wire [4-1:0] node50280;
	wire [4-1:0] node50281;
	wire [4-1:0] node50284;
	wire [4-1:0] node50287;
	wire [4-1:0] node50289;
	wire [4-1:0] node50292;
	wire [4-1:0] node50293;
	wire [4-1:0] node50294;
	wire [4-1:0] node50297;
	wire [4-1:0] node50300;
	wire [4-1:0] node50301;
	wire [4-1:0] node50304;
	wire [4-1:0] node50307;
	wire [4-1:0] node50308;
	wire [4-1:0] node50309;
	wire [4-1:0] node50310;
	wire [4-1:0] node50311;
	wire [4-1:0] node50312;
	wire [4-1:0] node50316;
	wire [4-1:0] node50317;
	wire [4-1:0] node50321;
	wire [4-1:0] node50322;
	wire [4-1:0] node50323;
	wire [4-1:0] node50327;
	wire [4-1:0] node50328;
	wire [4-1:0] node50332;
	wire [4-1:0] node50333;
	wire [4-1:0] node50334;
	wire [4-1:0] node50335;
	wire [4-1:0] node50339;
	wire [4-1:0] node50340;
	wire [4-1:0] node50344;
	wire [4-1:0] node50345;
	wire [4-1:0] node50346;
	wire [4-1:0] node50350;
	wire [4-1:0] node50351;
	wire [4-1:0] node50355;
	wire [4-1:0] node50356;
	wire [4-1:0] node50357;
	wire [4-1:0] node50358;
	wire [4-1:0] node50359;
	wire [4-1:0] node50361;
	wire [4-1:0] node50362;
	wire [4-1:0] node50365;
	wire [4-1:0] node50368;
	wire [4-1:0] node50369;
	wire [4-1:0] node50370;
	wire [4-1:0] node50373;
	wire [4-1:0] node50376;
	wire [4-1:0] node50377;
	wire [4-1:0] node50380;
	wire [4-1:0] node50383;
	wire [4-1:0] node50384;
	wire [4-1:0] node50385;
	wire [4-1:0] node50386;
	wire [4-1:0] node50389;
	wire [4-1:0] node50392;
	wire [4-1:0] node50393;
	wire [4-1:0] node50397;
	wire [4-1:0] node50398;
	wire [4-1:0] node50399;
	wire [4-1:0] node50402;
	wire [4-1:0] node50405;
	wire [4-1:0] node50406;
	wire [4-1:0] node50409;
	wire [4-1:0] node50412;
	wire [4-1:0] node50413;
	wire [4-1:0] node50414;
	wire [4-1:0] node50417;
	wire [4-1:0] node50420;
	wire [4-1:0] node50421;
	wire [4-1:0] node50423;
	wire [4-1:0] node50424;
	wire [4-1:0] node50428;
	wire [4-1:0] node50429;
	wire [4-1:0] node50432;
	wire [4-1:0] node50435;
	wire [4-1:0] node50436;
	wire [4-1:0] node50437;
	wire [4-1:0] node50438;
	wire [4-1:0] node50439;
	wire [4-1:0] node50440;
	wire [4-1:0] node50443;
	wire [4-1:0] node50447;
	wire [4-1:0] node50448;
	wire [4-1:0] node50449;
	wire [4-1:0] node50452;
	wire [4-1:0] node50455;
	wire [4-1:0] node50456;
	wire [4-1:0] node50459;
	wire [4-1:0] node50462;
	wire [4-1:0] node50463;
	wire [4-1:0] node50466;
	wire [4-1:0] node50469;
	wire [4-1:0] node50470;
	wire [4-1:0] node50471;
	wire [4-1:0] node50472;
	wire [4-1:0] node50476;
	wire [4-1:0] node50477;
	wire [4-1:0] node50481;
	wire [4-1:0] node50482;
	wire [4-1:0] node50483;
	wire [4-1:0] node50487;
	wire [4-1:0] node50488;
	wire [4-1:0] node50492;
	wire [4-1:0] node50493;
	wire [4-1:0] node50494;
	wire [4-1:0] node50495;
	wire [4-1:0] node50496;
	wire [4-1:0] node50497;
	wire [4-1:0] node50498;
	wire [4-1:0] node50499;
	wire [4-1:0] node50500;
	wire [4-1:0] node50503;
	wire [4-1:0] node50507;
	wire [4-1:0] node50508;
	wire [4-1:0] node50509;
	wire [4-1:0] node50513;
	wire [4-1:0] node50515;
	wire [4-1:0] node50518;
	wire [4-1:0] node50519;
	wire [4-1:0] node50520;
	wire [4-1:0] node50522;
	wire [4-1:0] node50525;
	wire [4-1:0] node50528;
	wire [4-1:0] node50529;
	wire [4-1:0] node50530;
	wire [4-1:0] node50534;
	wire [4-1:0] node50537;
	wire [4-1:0] node50538;
	wire [4-1:0] node50539;
	wire [4-1:0] node50540;
	wire [4-1:0] node50541;
	wire [4-1:0] node50545;
	wire [4-1:0] node50546;
	wire [4-1:0] node50549;
	wire [4-1:0] node50552;
	wire [4-1:0] node50554;
	wire [4-1:0] node50555;
	wire [4-1:0] node50558;
	wire [4-1:0] node50561;
	wire [4-1:0] node50562;
	wire [4-1:0] node50563;
	wire [4-1:0] node50564;
	wire [4-1:0] node50568;
	wire [4-1:0] node50569;
	wire [4-1:0] node50572;
	wire [4-1:0] node50575;
	wire [4-1:0] node50576;
	wire [4-1:0] node50577;
	wire [4-1:0] node50580;
	wire [4-1:0] node50583;
	wire [4-1:0] node50585;
	wire [4-1:0] node50588;
	wire [4-1:0] node50589;
	wire [4-1:0] node50590;
	wire [4-1:0] node50591;
	wire [4-1:0] node50594;
	wire [4-1:0] node50597;
	wire [4-1:0] node50598;
	wire [4-1:0] node50601;
	wire [4-1:0] node50604;
	wire [4-1:0] node50605;
	wire [4-1:0] node50608;
	wire [4-1:0] node50611;
	wire [4-1:0] node50612;
	wire [4-1:0] node50613;
	wire [4-1:0] node50614;
	wire [4-1:0] node50615;
	wire [4-1:0] node50618;
	wire [4-1:0] node50622;
	wire [4-1:0] node50623;
	wire [4-1:0] node50624;
	wire [4-1:0] node50625;
	wire [4-1:0] node50628;
	wire [4-1:0] node50631;
	wire [4-1:0] node50632;
	wire [4-1:0] node50635;
	wire [4-1:0] node50639;
	wire [4-1:0] node50640;
	wire [4-1:0] node50641;
	wire [4-1:0] node50645;
	wire [4-1:0] node50646;
	wire [4-1:0] node50650;
	wire [4-1:0] node50651;
	wire [4-1:0] node50652;
	wire [4-1:0] node50653;
	wire [4-1:0] node50656;
	wire [4-1:0] node50659;
	wire [4-1:0] node50660;
	wire [4-1:0] node50661;
	wire [4-1:0] node50664;
	wire [4-1:0] node50667;
	wire [4-1:0] node50668;
	wire [4-1:0] node50670;
	wire [4-1:0] node50671;
	wire [4-1:0] node50672;
	wire [4-1:0] node50675;
	wire [4-1:0] node50678;
	wire [4-1:0] node50679;
	wire [4-1:0] node50682;
	wire [4-1:0] node50685;
	wire [4-1:0] node50686;
	wire [4-1:0] node50689;
	wire [4-1:0] node50692;
	wire [4-1:0] node50693;
	wire [4-1:0] node50694;
	wire [4-1:0] node50695;
	wire [4-1:0] node50696;
	wire [4-1:0] node50700;
	wire [4-1:0] node50701;
	wire [4-1:0] node50705;
	wire [4-1:0] node50706;
	wire [4-1:0] node50707;
	wire [4-1:0] node50711;
	wire [4-1:0] node50712;
	wire [4-1:0] node50716;
	wire [4-1:0] node50717;
	wire [4-1:0] node50718;
	wire [4-1:0] node50719;
	wire [4-1:0] node50720;
	wire [4-1:0] node50723;
	wire [4-1:0] node50726;
	wire [4-1:0] node50727;
	wire [4-1:0] node50730;
	wire [4-1:0] node50733;
	wire [4-1:0] node50734;
	wire [4-1:0] node50735;
	wire [4-1:0] node50736;
	wire [4-1:0] node50740;
	wire [4-1:0] node50741;
	wire [4-1:0] node50744;
	wire [4-1:0] node50747;
	wire [4-1:0] node50748;
	wire [4-1:0] node50749;
	wire [4-1:0] node50752;
	wire [4-1:0] node50755;
	wire [4-1:0] node50756;
	wire [4-1:0] node50759;
	wire [4-1:0] node50762;
	wire [4-1:0] node50763;
	wire [4-1:0] node50766;
	wire [4-1:0] node50769;
	wire [4-1:0] node50770;
	wire [4-1:0] node50771;
	wire [4-1:0] node50772;
	wire [4-1:0] node50773;
	wire [4-1:0] node50774;
	wire [4-1:0] node50775;
	wire [4-1:0] node50776;
	wire [4-1:0] node50777;
	wire [4-1:0] node50778;
	wire [4-1:0] node50781;
	wire [4-1:0] node50784;
	wire [4-1:0] node50785;
	wire [4-1:0] node50788;
	wire [4-1:0] node50791;
	wire [4-1:0] node50792;
	wire [4-1:0] node50795;
	wire [4-1:0] node50798;
	wire [4-1:0] node50799;
	wire [4-1:0] node50800;
	wire [4-1:0] node50803;
	wire [4-1:0] node50806;
	wire [4-1:0] node50807;
	wire [4-1:0] node50810;
	wire [4-1:0] node50813;
	wire [4-1:0] node50814;
	wire [4-1:0] node50817;
	wire [4-1:0] node50820;
	wire [4-1:0] node50821;
	wire [4-1:0] node50822;
	wire [4-1:0] node50823;
	wire [4-1:0] node50824;
	wire [4-1:0] node50828;
	wire [4-1:0] node50829;
	wire [4-1:0] node50833;
	wire [4-1:0] node50834;
	wire [4-1:0] node50835;
	wire [4-1:0] node50839;
	wire [4-1:0] node50840;
	wire [4-1:0] node50844;
	wire [4-1:0] node50845;
	wire [4-1:0] node50846;
	wire [4-1:0] node50848;
	wire [4-1:0] node50849;
	wire [4-1:0] node50853;
	wire [4-1:0] node50855;
	wire [4-1:0] node50856;
	wire [4-1:0] node50860;
	wire [4-1:0] node50861;
	wire [4-1:0] node50862;
	wire [4-1:0] node50864;
	wire [4-1:0] node50867;
	wire [4-1:0] node50870;
	wire [4-1:0] node50871;
	wire [4-1:0] node50875;
	wire [4-1:0] node50876;
	wire [4-1:0] node50877;
	wire [4-1:0] node50878;
	wire [4-1:0] node50879;
	wire [4-1:0] node50880;
	wire [4-1:0] node50884;
	wire [4-1:0] node50885;
	wire [4-1:0] node50889;
	wire [4-1:0] node50890;
	wire [4-1:0] node50891;
	wire [4-1:0] node50895;
	wire [4-1:0] node50896;
	wire [4-1:0] node50900;
	wire [4-1:0] node50901;
	wire [4-1:0] node50902;
	wire [4-1:0] node50903;
	wire [4-1:0] node50906;
	wire [4-1:0] node50909;
	wire [4-1:0] node50910;
	wire [4-1:0] node50913;
	wire [4-1:0] node50916;
	wire [4-1:0] node50917;
	wire [4-1:0] node50918;
	wire [4-1:0] node50921;
	wire [4-1:0] node50924;
	wire [4-1:0] node50925;
	wire [4-1:0] node50928;
	wire [4-1:0] node50931;
	wire [4-1:0] node50932;
	wire [4-1:0] node50933;
	wire [4-1:0] node50934;
	wire [4-1:0] node50938;
	wire [4-1:0] node50939;
	wire [4-1:0] node50943;
	wire [4-1:0] node50944;
	wire [4-1:0] node50945;
	wire [4-1:0] node50949;
	wire [4-1:0] node50950;
	wire [4-1:0] node50954;
	wire [4-1:0] node50955;
	wire [4-1:0] node50956;
	wire [4-1:0] node50957;
	wire [4-1:0] node50958;
	wire [4-1:0] node50960;
	wire [4-1:0] node50963;
	wire [4-1:0] node50965;
	wire [4-1:0] node50968;
	wire [4-1:0] node50969;
	wire [4-1:0] node50971;
	wire [4-1:0] node50974;
	wire [4-1:0] node50976;
	wire [4-1:0] node50979;
	wire [4-1:0] node50980;
	wire [4-1:0] node50981;
	wire [4-1:0] node50982;
	wire [4-1:0] node50983;
	wire [4-1:0] node50987;
	wire [4-1:0] node50988;
	wire [4-1:0] node50992;
	wire [4-1:0] node50993;
	wire [4-1:0] node50994;
	wire [4-1:0] node50999;
	wire [4-1:0] node51000;
	wire [4-1:0] node51001;
	wire [4-1:0] node51002;
	wire [4-1:0] node51005;
	wire [4-1:0] node51008;
	wire [4-1:0] node51009;
	wire [4-1:0] node51010;
	wire [4-1:0] node51014;
	wire [4-1:0] node51016;
	wire [4-1:0] node51019;
	wire [4-1:0] node51020;
	wire [4-1:0] node51023;
	wire [4-1:0] node51026;
	wire [4-1:0] node51027;
	wire [4-1:0] node51028;
	wire [4-1:0] node51029;
	wire [4-1:0] node51033;
	wire [4-1:0] node51034;
	wire [4-1:0] node51038;
	wire [4-1:0] node51039;
	wire [4-1:0] node51040;
	wire [4-1:0] node51044;
	wire [4-1:0] node51045;
	wire [4-1:0] node51049;
	wire [4-1:0] node51050;
	wire [4-1:0] node51051;
	wire [4-1:0] node51052;
	wire [4-1:0] node51053;
	wire [4-1:0] node51057;
	wire [4-1:0] node51058;
	wire [4-1:0] node51063;
	wire [4-1:0] node51064;
	wire [4-1:0] node51065;
	wire [4-1:0] node51066;
	wire [4-1:0] node51070;
	wire [4-1:0] node51071;
	wire [4-1:0] node51076;
	wire [4-1:0] node51077;
	wire [4-1:0] node51078;
	wire [4-1:0] node51079;
	wire [4-1:0] node51080;
	wire [4-1:0] node51081;
	wire [4-1:0] node51082;
	wire [4-1:0] node51083;
	wire [4-1:0] node51084;
	wire [4-1:0] node51085;
	wire [4-1:0] node51086;
	wire [4-1:0] node51087;
	wire [4-1:0] node51089;
	wire [4-1:0] node51093;
	wire [4-1:0] node51094;
	wire [4-1:0] node51096;
	wire [4-1:0] node51099;
	wire [4-1:0] node51101;
	wire [4-1:0] node51104;
	wire [4-1:0] node51105;
	wire [4-1:0] node51106;
	wire [4-1:0] node51109;
	wire [4-1:0] node51112;
	wire [4-1:0] node51113;
	wire [4-1:0] node51114;
	wire [4-1:0] node51117;
	wire [4-1:0] node51121;
	wire [4-1:0] node51122;
	wire [4-1:0] node51123;
	wire [4-1:0] node51125;
	wire [4-1:0] node51128;
	wire [4-1:0] node51130;
	wire [4-1:0] node51133;
	wire [4-1:0] node51134;
	wire [4-1:0] node51136;
	wire [4-1:0] node51139;
	wire [4-1:0] node51142;
	wire [4-1:0] node51143;
	wire [4-1:0] node51144;
	wire [4-1:0] node51147;
	wire [4-1:0] node51150;
	wire [4-1:0] node51151;
	wire [4-1:0] node51152;
	wire [4-1:0] node51155;
	wire [4-1:0] node51158;
	wire [4-1:0] node51159;
	wire [4-1:0] node51162;
	wire [4-1:0] node51165;
	wire [4-1:0] node51166;
	wire [4-1:0] node51167;
	wire [4-1:0] node51168;
	wire [4-1:0] node51170;
	wire [4-1:0] node51173;
	wire [4-1:0] node51175;
	wire [4-1:0] node51178;
	wire [4-1:0] node51179;
	wire [4-1:0] node51181;
	wire [4-1:0] node51184;
	wire [4-1:0] node51186;
	wire [4-1:0] node51189;
	wire [4-1:0] node51190;
	wire [4-1:0] node51191;
	wire [4-1:0] node51192;
	wire [4-1:0] node51195;
	wire [4-1:0] node51198;
	wire [4-1:0] node51199;
	wire [4-1:0] node51200;
	wire [4-1:0] node51203;
	wire [4-1:0] node51206;
	wire [4-1:0] node51207;
	wire [4-1:0] node51208;
	wire [4-1:0] node51212;
	wire [4-1:0] node51213;
	wire [4-1:0] node51216;
	wire [4-1:0] node51219;
	wire [4-1:0] node51220;
	wire [4-1:0] node51221;
	wire [4-1:0] node51224;
	wire [4-1:0] node51227;
	wire [4-1:0] node51228;
	wire [4-1:0] node51229;
	wire [4-1:0] node51232;
	wire [4-1:0] node51235;
	wire [4-1:0] node51236;
	wire [4-1:0] node51239;
	wire [4-1:0] node51242;
	wire [4-1:0] node51243;
	wire [4-1:0] node51244;
	wire [4-1:0] node51245;
	wire [4-1:0] node51248;
	wire [4-1:0] node51251;
	wire [4-1:0] node51252;
	wire [4-1:0] node51253;
	wire [4-1:0] node51254;
	wire [4-1:0] node51255;
	wire [4-1:0] node51256;
	wire [4-1:0] node51259;
	wire [4-1:0] node51262;
	wire [4-1:0] node51263;
	wire [4-1:0] node51266;
	wire [4-1:0] node51269;
	wire [4-1:0] node51270;
	wire [4-1:0] node51273;
	wire [4-1:0] node51276;
	wire [4-1:0] node51277;
	wire [4-1:0] node51278;
	wire [4-1:0] node51279;
	wire [4-1:0] node51282;
	wire [4-1:0] node51285;
	wire [4-1:0] node51286;
	wire [4-1:0] node51289;
	wire [4-1:0] node51292;
	wire [4-1:0] node51293;
	wire [4-1:0] node51294;
	wire [4-1:0] node51297;
	wire [4-1:0] node51300;
	wire [4-1:0] node51302;
	wire [4-1:0] node51305;
	wire [4-1:0] node51306;
	wire [4-1:0] node51307;
	wire [4-1:0] node51308;
	wire [4-1:0] node51309;
	wire [4-1:0] node51313;
	wire [4-1:0] node51314;
	wire [4-1:0] node51317;
	wire [4-1:0] node51320;
	wire [4-1:0] node51321;
	wire [4-1:0] node51325;
	wire [4-1:0] node51326;
	wire [4-1:0] node51329;
	wire [4-1:0] node51332;
	wire [4-1:0] node51333;
	wire [4-1:0] node51334;
	wire [4-1:0] node51335;
	wire [4-1:0] node51336;
	wire [4-1:0] node51337;
	wire [4-1:0] node51340;
	wire [4-1:0] node51343;
	wire [4-1:0] node51344;
	wire [4-1:0] node51347;
	wire [4-1:0] node51350;
	wire [4-1:0] node51351;
	wire [4-1:0] node51352;
	wire [4-1:0] node51355;
	wire [4-1:0] node51358;
	wire [4-1:0] node51359;
	wire [4-1:0] node51362;
	wire [4-1:0] node51365;
	wire [4-1:0] node51366;
	wire [4-1:0] node51367;
	wire [4-1:0] node51370;
	wire [4-1:0] node51373;
	wire [4-1:0] node51374;
	wire [4-1:0] node51377;
	wire [4-1:0] node51380;
	wire [4-1:0] node51381;
	wire [4-1:0] node51382;
	wire [4-1:0] node51385;
	wire [4-1:0] node51388;
	wire [4-1:0] node51389;
	wire [4-1:0] node51390;
	wire [4-1:0] node51393;
	wire [4-1:0] node51396;
	wire [4-1:0] node51397;
	wire [4-1:0] node51398;
	wire [4-1:0] node51401;
	wire [4-1:0] node51404;
	wire [4-1:0] node51405;
	wire [4-1:0] node51408;
	wire [4-1:0] node51411;
	wire [4-1:0] node51412;
	wire [4-1:0] node51413;
	wire [4-1:0] node51414;
	wire [4-1:0] node51415;
	wire [4-1:0] node51418;
	wire [4-1:0] node51421;
	wire [4-1:0] node51422;
	wire [4-1:0] node51423;
	wire [4-1:0] node51424;
	wire [4-1:0] node51425;
	wire [4-1:0] node51428;
	wire [4-1:0] node51431;
	wire [4-1:0] node51432;
	wire [4-1:0] node51433;
	wire [4-1:0] node51436;
	wire [4-1:0] node51439;
	wire [4-1:0] node51440;
	wire [4-1:0] node51443;
	wire [4-1:0] node51446;
	wire [4-1:0] node51447;
	wire [4-1:0] node51448;
	wire [4-1:0] node51451;
	wire [4-1:0] node51454;
	wire [4-1:0] node51455;
	wire [4-1:0] node51458;
	wire [4-1:0] node51461;
	wire [4-1:0] node51462;
	wire [4-1:0] node51463;
	wire [4-1:0] node51464;
	wire [4-1:0] node51465;
	wire [4-1:0] node51469;
	wire [4-1:0] node51470;
	wire [4-1:0] node51473;
	wire [4-1:0] node51476;
	wire [4-1:0] node51477;
	wire [4-1:0] node51478;
	wire [4-1:0] node51481;
	wire [4-1:0] node51484;
	wire [4-1:0] node51486;
	wire [4-1:0] node51489;
	wire [4-1:0] node51490;
	wire [4-1:0] node51491;
	wire [4-1:0] node51494;
	wire [4-1:0] node51497;
	wire [4-1:0] node51498;
	wire [4-1:0] node51499;
	wire [4-1:0] node51502;
	wire [4-1:0] node51506;
	wire [4-1:0] node51507;
	wire [4-1:0] node51508;
	wire [4-1:0] node51509;
	wire [4-1:0] node51510;
	wire [4-1:0] node51511;
	wire [4-1:0] node51515;
	wire [4-1:0] node51516;
	wire [4-1:0] node51517;
	wire [4-1:0] node51520;
	wire [4-1:0] node51524;
	wire [4-1:0] node51525;
	wire [4-1:0] node51526;
	wire [4-1:0] node51527;
	wire [4-1:0] node51530;
	wire [4-1:0] node51534;
	wire [4-1:0] node51535;
	wire [4-1:0] node51536;
	wire [4-1:0] node51539;
	wire [4-1:0] node51543;
	wire [4-1:0] node51544;
	wire [4-1:0] node51545;
	wire [4-1:0] node51546;
	wire [4-1:0] node51547;
	wire [4-1:0] node51550;
	wire [4-1:0] node51554;
	wire [4-1:0] node51555;
	wire [4-1:0] node51557;
	wire [4-1:0] node51561;
	wire [4-1:0] node51562;
	wire [4-1:0] node51563;
	wire [4-1:0] node51564;
	wire [4-1:0] node51569;
	wire [4-1:0] node51570;
	wire [4-1:0] node51571;
	wire [4-1:0] node51574;
	wire [4-1:0] node51578;
	wire [4-1:0] node51579;
	wire [4-1:0] node51580;
	wire [4-1:0] node51581;
	wire [4-1:0] node51583;
	wire [4-1:0] node51584;
	wire [4-1:0] node51587;
	wire [4-1:0] node51590;
	wire [4-1:0] node51591;
	wire [4-1:0] node51592;
	wire [4-1:0] node51595;
	wire [4-1:0] node51598;
	wire [4-1:0] node51599;
	wire [4-1:0] node51602;
	wire [4-1:0] node51605;
	wire [4-1:0] node51606;
	wire [4-1:0] node51607;
	wire [4-1:0] node51608;
	wire [4-1:0] node51611;
	wire [4-1:0] node51614;
	wire [4-1:0] node51616;
	wire [4-1:0] node51619;
	wire [4-1:0] node51620;
	wire [4-1:0] node51621;
	wire [4-1:0] node51625;
	wire [4-1:0] node51626;
	wire [4-1:0] node51629;
	wire [4-1:0] node51632;
	wire [4-1:0] node51633;
	wire [4-1:0] node51634;
	wire [4-1:0] node51637;
	wire [4-1:0] node51640;
	wire [4-1:0] node51641;
	wire [4-1:0] node51644;
	wire [4-1:0] node51647;
	wire [4-1:0] node51648;
	wire [4-1:0] node51649;
	wire [4-1:0] node51650;
	wire [4-1:0] node51651;
	wire [4-1:0] node51652;
	wire [4-1:0] node51653;
	wire [4-1:0] node51656;
	wire [4-1:0] node51659;
	wire [4-1:0] node51660;
	wire [4-1:0] node51663;
	wire [4-1:0] node51667;
	wire [4-1:0] node51668;
	wire [4-1:0] node51669;
	wire [4-1:0] node51670;
	wire [4-1:0] node51673;
	wire [4-1:0] node51676;
	wire [4-1:0] node51677;
	wire [4-1:0] node51680;
	wire [4-1:0] node51684;
	wire [4-1:0] node51685;
	wire [4-1:0] node51686;
	wire [4-1:0] node51687;
	wire [4-1:0] node51690;
	wire [4-1:0] node51694;
	wire [4-1:0] node51695;
	wire [4-1:0] node51696;
	wire [4-1:0] node51698;
	wire [4-1:0] node51701;
	wire [4-1:0] node51702;
	wire [4-1:0] node51705;
	wire [4-1:0] node51709;
	wire [4-1:0] node51710;
	wire [4-1:0] node51711;
	wire [4-1:0] node51712;
	wire [4-1:0] node51713;
	wire [4-1:0] node51714;
	wire [4-1:0] node51715;
	wire [4-1:0] node51718;
	wire [4-1:0] node51721;
	wire [4-1:0] node51722;
	wire [4-1:0] node51725;
	wire [4-1:0] node51728;
	wire [4-1:0] node51729;
	wire [4-1:0] node51732;
	wire [4-1:0] node51735;
	wire [4-1:0] node51736;
	wire [4-1:0] node51737;
	wire [4-1:0] node51738;
	wire [4-1:0] node51741;
	wire [4-1:0] node51744;
	wire [4-1:0] node51745;
	wire [4-1:0] node51748;
	wire [4-1:0] node51751;
	wire [4-1:0] node51752;
	wire [4-1:0] node51753;
	wire [4-1:0] node51756;
	wire [4-1:0] node51759;
	wire [4-1:0] node51760;
	wire [4-1:0] node51763;
	wire [4-1:0] node51766;
	wire [4-1:0] node51767;
	wire [4-1:0] node51768;
	wire [4-1:0] node51771;
	wire [4-1:0] node51774;
	wire [4-1:0] node51775;
	wire [4-1:0] node51778;
	wire [4-1:0] node51781;
	wire [4-1:0] node51782;
	wire [4-1:0] node51783;
	wire [4-1:0] node51784;
	wire [4-1:0] node51785;
	wire [4-1:0] node51788;
	wire [4-1:0] node51792;
	wire [4-1:0] node51793;
	wire [4-1:0] node51794;
	wire [4-1:0] node51797;
	wire [4-1:0] node51801;
	wire [4-1:0] node51802;
	wire [4-1:0] node51803;
	wire [4-1:0] node51804;
	wire [4-1:0] node51805;
	wire [4-1:0] node51808;
	wire [4-1:0] node51811;
	wire [4-1:0] node51813;
	wire [4-1:0] node51817;
	wire [4-1:0] node51818;
	wire [4-1:0] node51819;
	wire [4-1:0] node51821;
	wire [4-1:0] node51824;
	wire [4-1:0] node51825;
	wire [4-1:0] node51828;
	wire [4-1:0] node51832;
	wire [4-1:0] node51833;
	wire [4-1:0] node51834;
	wire [4-1:0] node51835;
	wire [4-1:0] node51836;
	wire [4-1:0] node51837;
	wire [4-1:0] node51838;
	wire [4-1:0] node51840;
	wire [4-1:0] node51842;
	wire [4-1:0] node51844;
	wire [4-1:0] node51847;
	wire [4-1:0] node51848;
	wire [4-1:0] node51849;
	wire [4-1:0] node51851;
	wire [4-1:0] node51855;
	wire [4-1:0] node51857;
	wire [4-1:0] node51859;
	wire [4-1:0] node51862;
	wire [4-1:0] node51863;
	wire [4-1:0] node51864;
	wire [4-1:0] node51865;
	wire [4-1:0] node51866;
	wire [4-1:0] node51869;
	wire [4-1:0] node51872;
	wire [4-1:0] node51873;
	wire [4-1:0] node51876;
	wire [4-1:0] node51879;
	wire [4-1:0] node51880;
	wire [4-1:0] node51881;
	wire [4-1:0] node51884;
	wire [4-1:0] node51888;
	wire [4-1:0] node51889;
	wire [4-1:0] node51890;
	wire [4-1:0] node51893;
	wire [4-1:0] node51896;
	wire [4-1:0] node51897;
	wire [4-1:0] node51898;
	wire [4-1:0] node51901;
	wire [4-1:0] node51904;
	wire [4-1:0] node51905;
	wire [4-1:0] node51909;
	wire [4-1:0] node51910;
	wire [4-1:0] node51911;
	wire [4-1:0] node51912;
	wire [4-1:0] node51913;
	wire [4-1:0] node51916;
	wire [4-1:0] node51919;
	wire [4-1:0] node51920;
	wire [4-1:0] node51921;
	wire [4-1:0] node51924;
	wire [4-1:0] node51928;
	wire [4-1:0] node51929;
	wire [4-1:0] node51930;
	wire [4-1:0] node51933;
	wire [4-1:0] node51936;
	wire [4-1:0] node51937;
	wire [4-1:0] node51938;
	wire [4-1:0] node51941;
	wire [4-1:0] node51944;
	wire [4-1:0] node51945;
	wire [4-1:0] node51948;
	wire [4-1:0] node51951;
	wire [4-1:0] node51952;
	wire [4-1:0] node51953;
	wire [4-1:0] node51954;
	wire [4-1:0] node51956;
	wire [4-1:0] node51959;
	wire [4-1:0] node51961;
	wire [4-1:0] node51964;
	wire [4-1:0] node51965;
	wire [4-1:0] node51967;
	wire [4-1:0] node51970;
	wire [4-1:0] node51971;
	wire [4-1:0] node51975;
	wire [4-1:0] node51976;
	wire [4-1:0] node51977;
	wire [4-1:0] node51978;
	wire [4-1:0] node51981;
	wire [4-1:0] node51984;
	wire [4-1:0] node51985;
	wire [4-1:0] node51988;
	wire [4-1:0] node51991;
	wire [4-1:0] node51992;
	wire [4-1:0] node51993;
	wire [4-1:0] node51996;
	wire [4-1:0] node51999;
	wire [4-1:0] node52000;
	wire [4-1:0] node52003;
	wire [4-1:0] node52006;
	wire [4-1:0] node52007;
	wire [4-1:0] node52008;
	wire [4-1:0] node52009;
	wire [4-1:0] node52011;
	wire [4-1:0] node52012;
	wire [4-1:0] node52013;
	wire [4-1:0] node52016;
	wire [4-1:0] node52019;
	wire [4-1:0] node52020;
	wire [4-1:0] node52023;
	wire [4-1:0] node52026;
	wire [4-1:0] node52028;
	wire [4-1:0] node52029;
	wire [4-1:0] node52030;
	wire [4-1:0] node52033;
	wire [4-1:0] node52036;
	wire [4-1:0] node52038;
	wire [4-1:0] node52041;
	wire [4-1:0] node52042;
	wire [4-1:0] node52044;
	wire [4-1:0] node52045;
	wire [4-1:0] node52046;
	wire [4-1:0] node52049;
	wire [4-1:0] node52052;
	wire [4-1:0] node52054;
	wire [4-1:0] node52057;
	wire [4-1:0] node52059;
	wire [4-1:0] node52060;
	wire [4-1:0] node52063;
	wire [4-1:0] node52066;
	wire [4-1:0] node52067;
	wire [4-1:0] node52068;
	wire [4-1:0] node52069;
	wire [4-1:0] node52072;
	wire [4-1:0] node52075;
	wire [4-1:0] node52076;
	wire [4-1:0] node52079;
	wire [4-1:0] node52082;
	wire [4-1:0] node52083;
	wire [4-1:0] node52084;
	wire [4-1:0] node52085;
	wire [4-1:0] node52088;
	wire [4-1:0] node52091;
	wire [4-1:0] node52092;
	wire [4-1:0] node52095;
	wire [4-1:0] node52098;
	wire [4-1:0] node52099;
	wire [4-1:0] node52100;
	wire [4-1:0] node52102;
	wire [4-1:0] node52105;
	wire [4-1:0] node52106;
	wire [4-1:0] node52109;
	wire [4-1:0] node52112;
	wire [4-1:0] node52113;
	wire [4-1:0] node52117;
	wire [4-1:0] node52118;
	wire [4-1:0] node52119;
	wire [4-1:0] node52120;
	wire [4-1:0] node52121;
	wire [4-1:0] node52123;
	wire [4-1:0] node52125;
	wire [4-1:0] node52128;
	wire [4-1:0] node52129;
	wire [4-1:0] node52130;
	wire [4-1:0] node52133;
	wire [4-1:0] node52136;
	wire [4-1:0] node52137;
	wire [4-1:0] node52141;
	wire [4-1:0] node52142;
	wire [4-1:0] node52143;
	wire [4-1:0] node52145;
	wire [4-1:0] node52148;
	wire [4-1:0] node52149;
	wire [4-1:0] node52152;
	wire [4-1:0] node52155;
	wire [4-1:0] node52156;
	wire [4-1:0] node52157;
	wire [4-1:0] node52158;
	wire [4-1:0] node52164;
	wire [4-1:0] node52165;
	wire [4-1:0] node52166;
	wire [4-1:0] node52168;
	wire [4-1:0] node52170;
	wire [4-1:0] node52173;
	wire [4-1:0] node52174;
	wire [4-1:0] node52175;
	wire [4-1:0] node52177;
	wire [4-1:0] node52180;
	wire [4-1:0] node52181;
	wire [4-1:0] node52185;
	wire [4-1:0] node52186;
	wire [4-1:0] node52190;
	wire [4-1:0] node52191;
	wire [4-1:0] node52192;
	wire [4-1:0] node52194;
	wire [4-1:0] node52197;
	wire [4-1:0] node52198;
	wire [4-1:0] node52201;
	wire [4-1:0] node52204;
	wire [4-1:0] node52206;
	wire [4-1:0] node52207;
	wire [4-1:0] node52211;
	wire [4-1:0] node52212;
	wire [4-1:0] node52213;
	wire [4-1:0] node52214;
	wire [4-1:0] node52215;
	wire [4-1:0] node52217;
	wire [4-1:0] node52220;
	wire [4-1:0] node52222;
	wire [4-1:0] node52225;
	wire [4-1:0] node52226;
	wire [4-1:0] node52228;
	wire [4-1:0] node52231;
	wire [4-1:0] node52233;
	wire [4-1:0] node52236;
	wire [4-1:0] node52237;
	wire [4-1:0] node52238;
	wire [4-1:0] node52239;
	wire [4-1:0] node52240;
	wire [4-1:0] node52244;
	wire [4-1:0] node52246;
	wire [4-1:0] node52249;
	wire [4-1:0] node52250;
	wire [4-1:0] node52253;
	wire [4-1:0] node52256;
	wire [4-1:0] node52257;
	wire [4-1:0] node52258;
	wire [4-1:0] node52261;
	wire [4-1:0] node52264;
	wire [4-1:0] node52265;
	wire [4-1:0] node52269;
	wire [4-1:0] node52270;
	wire [4-1:0] node52271;
	wire [4-1:0] node52272;
	wire [4-1:0] node52273;
	wire [4-1:0] node52278;
	wire [4-1:0] node52279;
	wire [4-1:0] node52281;
	wire [4-1:0] node52285;
	wire [4-1:0] node52286;
	wire [4-1:0] node52287;
	wire [4-1:0] node52289;
	wire [4-1:0] node52293;
	wire [4-1:0] node52294;
	wire [4-1:0] node52295;
	wire [4-1:0] node52300;
	wire [4-1:0] node52301;
	wire [4-1:0] node52302;
	wire [4-1:0] node52303;
	wire [4-1:0] node52304;
	wire [4-1:0] node52305;
	wire [4-1:0] node52308;
	wire [4-1:0] node52311;
	wire [4-1:0] node52312;
	wire [4-1:0] node52313;
	wire [4-1:0] node52314;
	wire [4-1:0] node52315;
	wire [4-1:0] node52318;
	wire [4-1:0] node52321;
	wire [4-1:0] node52322;
	wire [4-1:0] node52325;
	wire [4-1:0] node52328;
	wire [4-1:0] node52329;
	wire [4-1:0] node52330;
	wire [4-1:0] node52333;
	wire [4-1:0] node52336;
	wire [4-1:0] node52337;
	wire [4-1:0] node52340;
	wire [4-1:0] node52343;
	wire [4-1:0] node52344;
	wire [4-1:0] node52347;
	wire [4-1:0] node52350;
	wire [4-1:0] node52351;
	wire [4-1:0] node52352;
	wire [4-1:0] node52353;
	wire [4-1:0] node52354;
	wire [4-1:0] node52357;
	wire [4-1:0] node52361;
	wire [4-1:0] node52362;
	wire [4-1:0] node52363;
	wire [4-1:0] node52366;
	wire [4-1:0] node52369;
	wire [4-1:0] node52370;
	wire [4-1:0] node52373;
	wire [4-1:0] node52376;
	wire [4-1:0] node52377;
	wire [4-1:0] node52378;
	wire [4-1:0] node52379;
	wire [4-1:0] node52383;
	wire [4-1:0] node52384;
	wire [4-1:0] node52388;
	wire [4-1:0] node52389;
	wire [4-1:0] node52391;
	wire [4-1:0] node52394;
	wire [4-1:0] node52396;
	wire [4-1:0] node52399;
	wire [4-1:0] node52400;
	wire [4-1:0] node52401;
	wire [4-1:0] node52402;
	wire [4-1:0] node52403;
	wire [4-1:0] node52404;
	wire [4-1:0] node52407;
	wire [4-1:0] node52410;
	wire [4-1:0] node52411;
	wire [4-1:0] node52412;
	wire [4-1:0] node52415;
	wire [4-1:0] node52418;
	wire [4-1:0] node52420;
	wire [4-1:0] node52423;
	wire [4-1:0] node52424;
	wire [4-1:0] node52427;
	wire [4-1:0] node52430;
	wire [4-1:0] node52431;
	wire [4-1:0] node52432;
	wire [4-1:0] node52433;
	wire [4-1:0] node52434;
	wire [4-1:0] node52437;
	wire [4-1:0] node52440;
	wire [4-1:0] node52441;
	wire [4-1:0] node52444;
	wire [4-1:0] node52447;
	wire [4-1:0] node52448;
	wire [4-1:0] node52449;
	wire [4-1:0] node52453;
	wire [4-1:0] node52455;
	wire [4-1:0] node52458;
	wire [4-1:0] node52459;
	wire [4-1:0] node52460;
	wire [4-1:0] node52463;
	wire [4-1:0] node52466;
	wire [4-1:0] node52467;
	wire [4-1:0] node52470;
	wire [4-1:0] node52473;
	wire [4-1:0] node52474;
	wire [4-1:0] node52475;
	wire [4-1:0] node52476;
	wire [4-1:0] node52477;
	wire [4-1:0] node52480;
	wire [4-1:0] node52483;
	wire [4-1:0] node52484;
	wire [4-1:0] node52487;
	wire [4-1:0] node52490;
	wire [4-1:0] node52491;
	wire [4-1:0] node52492;
	wire [4-1:0] node52495;
	wire [4-1:0] node52498;
	wire [4-1:0] node52499;
	wire [4-1:0] node52502;
	wire [4-1:0] node52505;
	wire [4-1:0] node52506;
	wire [4-1:0] node52507;
	wire [4-1:0] node52509;
	wire [4-1:0] node52510;
	wire [4-1:0] node52514;
	wire [4-1:0] node52515;
	wire [4-1:0] node52519;
	wire [4-1:0] node52520;
	wire [4-1:0] node52521;
	wire [4-1:0] node52525;
	wire [4-1:0] node52526;
	wire [4-1:0] node52530;
	wire [4-1:0] node52531;
	wire [4-1:0] node52532;
	wire [4-1:0] node52533;
	wire [4-1:0] node52534;
	wire [4-1:0] node52535;
	wire [4-1:0] node52536;
	wire [4-1:0] node52537;
	wire [4-1:0] node52540;
	wire [4-1:0] node52543;
	wire [4-1:0] node52544;
	wire [4-1:0] node52548;
	wire [4-1:0] node52549;
	wire [4-1:0] node52553;
	wire [4-1:0] node52554;
	wire [4-1:0] node52556;
	wire [4-1:0] node52560;
	wire [4-1:0] node52561;
	wire [4-1:0] node52562;
	wire [4-1:0] node52563;
	wire [4-1:0] node52567;
	wire [4-1:0] node52568;
	wire [4-1:0] node52569;
	wire [4-1:0] node52572;
	wire [4-1:0] node52575;
	wire [4-1:0] node52576;
	wire [4-1:0] node52579;
	wire [4-1:0] node52583;
	wire [4-1:0] node52584;
	wire [4-1:0] node52585;
	wire [4-1:0] node52586;
	wire [4-1:0] node52587;
	wire [4-1:0] node52590;
	wire [4-1:0] node52593;
	wire [4-1:0] node52595;
	wire [4-1:0] node52598;
	wire [4-1:0] node52600;
	wire [4-1:0] node52601;
	wire [4-1:0] node52605;
	wire [4-1:0] node52606;
	wire [4-1:0] node52607;
	wire [4-1:0] node52608;
	wire [4-1:0] node52612;
	wire [4-1:0] node52613;
	wire [4-1:0] node52616;
	wire [4-1:0] node52619;
	wire [4-1:0] node52620;
	wire [4-1:0] node52622;
	wire [4-1:0] node52626;
	wire [4-1:0] node52627;
	wire [4-1:0] node52628;
	wire [4-1:0] node52629;
	wire [4-1:0] node52630;
	wire [4-1:0] node52632;
	wire [4-1:0] node52635;
	wire [4-1:0] node52636;
	wire [4-1:0] node52639;
	wire [4-1:0] node52640;
	wire [4-1:0] node52644;
	wire [4-1:0] node52645;
	wire [4-1:0] node52646;
	wire [4-1:0] node52648;
	wire [4-1:0] node52651;
	wire [4-1:0] node52653;
	wire [4-1:0] node52656;
	wire [4-1:0] node52657;
	wire [4-1:0] node52659;
	wire [4-1:0] node52662;
	wire [4-1:0] node52663;
	wire [4-1:0] node52667;
	wire [4-1:0] node52668;
	wire [4-1:0] node52669;
	wire [4-1:0] node52670;
	wire [4-1:0] node52671;
	wire [4-1:0] node52675;
	wire [4-1:0] node52676;
	wire [4-1:0] node52680;
	wire [4-1:0] node52681;
	wire [4-1:0] node52682;
	wire [4-1:0] node52687;
	wire [4-1:0] node52688;
	wire [4-1:0] node52689;
	wire [4-1:0] node52690;
	wire [4-1:0] node52694;
	wire [4-1:0] node52695;
	wire [4-1:0] node52698;
	wire [4-1:0] node52701;
	wire [4-1:0] node52702;
	wire [4-1:0] node52703;
	wire [4-1:0] node52706;
	wire [4-1:0] node52709;
	wire [4-1:0] node52710;
	wire [4-1:0] node52713;
	wire [4-1:0] node52716;
	wire [4-1:0] node52717;
	wire [4-1:0] node52718;
	wire [4-1:0] node52719;
	wire [4-1:0] node52720;
	wire [4-1:0] node52723;
	wire [4-1:0] node52726;
	wire [4-1:0] node52727;
	wire [4-1:0] node52730;
	wire [4-1:0] node52733;
	wire [4-1:0] node52734;
	wire [4-1:0] node52735;
	wire [4-1:0] node52736;
	wire [4-1:0] node52739;
	wire [4-1:0] node52742;
	wire [4-1:0] node52743;
	wire [4-1:0] node52746;
	wire [4-1:0] node52749;
	wire [4-1:0] node52751;
	wire [4-1:0] node52752;
	wire [4-1:0] node52756;
	wire [4-1:0] node52757;
	wire [4-1:0] node52758;
	wire [4-1:0] node52759;
	wire [4-1:0] node52763;
	wire [4-1:0] node52764;
	wire [4-1:0] node52768;
	wire [4-1:0] node52769;
	wire [4-1:0] node52770;
	wire [4-1:0] node52771;
	wire [4-1:0] node52776;
	wire [4-1:0] node52777;
	wire [4-1:0] node52781;
	wire [4-1:0] node52782;
	wire [4-1:0] node52783;
	wire [4-1:0] node52784;
	wire [4-1:0] node52785;
	wire [4-1:0] node52786;
	wire [4-1:0] node52787;
	wire [4-1:0] node52790;
	wire [4-1:0] node52793;
	wire [4-1:0] node52794;
	wire [4-1:0] node52797;
	wire [4-1:0] node52800;
	wire [4-1:0] node52801;
	wire [4-1:0] node52802;
	wire [4-1:0] node52803;
	wire [4-1:0] node52806;
	wire [4-1:0] node52809;
	wire [4-1:0] node52810;
	wire [4-1:0] node52811;
	wire [4-1:0] node52812;
	wire [4-1:0] node52815;
	wire [4-1:0] node52818;
	wire [4-1:0] node52819;
	wire [4-1:0] node52823;
	wire [4-1:0] node52824;
	wire [4-1:0] node52825;
	wire [4-1:0] node52828;
	wire [4-1:0] node52831;
	wire [4-1:0] node52832;
	wire [4-1:0] node52833;
	wire [4-1:0] node52836;
	wire [4-1:0] node52839;
	wire [4-1:0] node52840;
	wire [4-1:0] node52843;
	wire [4-1:0] node52846;
	wire [4-1:0] node52847;
	wire [4-1:0] node52848;
	wire [4-1:0] node52849;
	wire [4-1:0] node52850;
	wire [4-1:0] node52851;
	wire [4-1:0] node52854;
	wire [4-1:0] node52857;
	wire [4-1:0] node52858;
	wire [4-1:0] node52861;
	wire [4-1:0] node52864;
	wire [4-1:0] node52865;
	wire [4-1:0] node52868;
	wire [4-1:0] node52871;
	wire [4-1:0] node52872;
	wire [4-1:0] node52875;
	wire [4-1:0] node52878;
	wire [4-1:0] node52879;
	wire [4-1:0] node52880;
	wire [4-1:0] node52883;
	wire [4-1:0] node52886;
	wire [4-1:0] node52887;
	wire [4-1:0] node52890;
	wire [4-1:0] node52893;
	wire [4-1:0] node52894;
	wire [4-1:0] node52897;
	wire [4-1:0] node52900;
	wire [4-1:0] node52901;
	wire [4-1:0] node52902;
	wire [4-1:0] node52903;
	wire [4-1:0] node52904;
	wire [4-1:0] node52905;
	wire [4-1:0] node52906;
	wire [4-1:0] node52909;
	wire [4-1:0] node52912;
	wire [4-1:0] node52913;
	wire [4-1:0] node52916;
	wire [4-1:0] node52919;
	wire [4-1:0] node52920;
	wire [4-1:0] node52921;
	wire [4-1:0] node52924;
	wire [4-1:0] node52927;
	wire [4-1:0] node52928;
	wire [4-1:0] node52929;
	wire [4-1:0] node52932;
	wire [4-1:0] node52935;
	wire [4-1:0] node52936;
	wire [4-1:0] node52939;
	wire [4-1:0] node52943;
	wire [4-1:0] node52944;
	wire [4-1:0] node52945;
	wire [4-1:0] node52946;
	wire [4-1:0] node52949;
	wire [4-1:0] node52952;
	wire [4-1:0] node52953;
	wire [4-1:0] node52954;
	wire [4-1:0] node52957;
	wire [4-1:0] node52960;
	wire [4-1:0] node52961;
	wire [4-1:0] node52964;
	wire [4-1:0] node52968;
	wire [4-1:0] node52969;
	wire [4-1:0] node52970;
	wire [4-1:0] node52974;
	wire [4-1:0] node52975;
	wire [4-1:0] node52979;
	wire [4-1:0] node52980;
	wire [4-1:0] node52981;
	wire [4-1:0] node52982;
	wire [4-1:0] node52983;
	wire [4-1:0] node52984;
	wire [4-1:0] node52988;
	wire [4-1:0] node52990;
	wire [4-1:0] node52993;
	wire [4-1:0] node52994;
	wire [4-1:0] node52996;
	wire [4-1:0] node52999;
	wire [4-1:0] node53001;
	wire [4-1:0] node53004;
	wire [4-1:0] node53005;
	wire [4-1:0] node53006;
	wire [4-1:0] node53007;
	wire [4-1:0] node53008;
	wire [4-1:0] node53009;
	wire [4-1:0] node53012;
	wire [4-1:0] node53015;
	wire [4-1:0] node53016;
	wire [4-1:0] node53019;
	wire [4-1:0] node53022;
	wire [4-1:0] node53023;
	wire [4-1:0] node53024;
	wire [4-1:0] node53025;
	wire [4-1:0] node53026;
	wire [4-1:0] node53029;
	wire [4-1:0] node53033;
	wire [4-1:0] node53034;
	wire [4-1:0] node53035;
	wire [4-1:0] node53038;
	wire [4-1:0] node53041;
	wire [4-1:0] node53043;
	wire [4-1:0] node53046;
	wire [4-1:0] node53047;
	wire [4-1:0] node53048;
	wire [4-1:0] node53052;
	wire [4-1:0] node53053;
	wire [4-1:0] node53056;
	wire [4-1:0] node53059;
	wire [4-1:0] node53060;
	wire [4-1:0] node53061;
	wire [4-1:0] node53062;
	wire [4-1:0] node53063;
	wire [4-1:0] node53066;
	wire [4-1:0] node53069;
	wire [4-1:0] node53070;
	wire [4-1:0] node53071;
	wire [4-1:0] node53074;
	wire [4-1:0] node53077;
	wire [4-1:0] node53078;
	wire [4-1:0] node53081;
	wire [4-1:0] node53084;
	wire [4-1:0] node53085;
	wire [4-1:0] node53086;
	wire [4-1:0] node53088;
	wire [4-1:0] node53091;
	wire [4-1:0] node53092;
	wire [4-1:0] node53096;
	wire [4-1:0] node53097;
	wire [4-1:0] node53100;
	wire [4-1:0] node53103;
	wire [4-1:0] node53104;
	wire [4-1:0] node53105;
	wire [4-1:0] node53108;
	wire [4-1:0] node53111;
	wire [4-1:0] node53112;
	wire [4-1:0] node53115;
	wire [4-1:0] node53118;
	wire [4-1:0] node53119;
	wire [4-1:0] node53120;
	wire [4-1:0] node53123;
	wire [4-1:0] node53126;
	wire [4-1:0] node53127;
	wire [4-1:0] node53130;
	wire [4-1:0] node53133;
	wire [4-1:0] node53134;
	wire [4-1:0] node53135;
	wire [4-1:0] node53139;
	wire [4-1:0] node53140;
	wire [4-1:0] node53144;
	wire [4-1:0] node53145;
	wire [4-1:0] node53146;
	wire [4-1:0] node53147;
	wire [4-1:0] node53148;
	wire [4-1:0] node53149;
	wire [4-1:0] node53150;
	wire [4-1:0] node53151;
	wire [4-1:0] node53152;
	wire [4-1:0] node53153;
	wire [4-1:0] node53156;
	wire [4-1:0] node53159;
	wire [4-1:0] node53160;
	wire [4-1:0] node53161;
	wire [4-1:0] node53164;
	wire [4-1:0] node53167;
	wire [4-1:0] node53168;
	wire [4-1:0] node53169;
	wire [4-1:0] node53173;
	wire [4-1:0] node53175;
	wire [4-1:0] node53178;
	wire [4-1:0] node53179;
	wire [4-1:0] node53180;
	wire [4-1:0] node53183;
	wire [4-1:0] node53186;
	wire [4-1:0] node53187;
	wire [4-1:0] node53188;
	wire [4-1:0] node53191;
	wire [4-1:0] node53194;
	wire [4-1:0] node53195;
	wire [4-1:0] node53198;
	wire [4-1:0] node53201;
	wire [4-1:0] node53202;
	wire [4-1:0] node53203;
	wire [4-1:0] node53204;
	wire [4-1:0] node53205;
	wire [4-1:0] node53208;
	wire [4-1:0] node53211;
	wire [4-1:0] node53212;
	wire [4-1:0] node53213;
	wire [4-1:0] node53216;
	wire [4-1:0] node53219;
	wire [4-1:0] node53220;
	wire [4-1:0] node53223;
	wire [4-1:0] node53226;
	wire [4-1:0] node53227;
	wire [4-1:0] node53230;
	wire [4-1:0] node53233;
	wire [4-1:0] node53234;
	wire [4-1:0] node53235;
	wire [4-1:0] node53236;
	wire [4-1:0] node53239;
	wire [4-1:0] node53242;
	wire [4-1:0] node53244;
	wire [4-1:0] node53245;
	wire [4-1:0] node53248;
	wire [4-1:0] node53251;
	wire [4-1:0] node53252;
	wire [4-1:0] node53255;
	wire [4-1:0] node53258;
	wire [4-1:0] node53259;
	wire [4-1:0] node53260;
	wire [4-1:0] node53261;
	wire [4-1:0] node53262;
	wire [4-1:0] node53265;
	wire [4-1:0] node53268;
	wire [4-1:0] node53269;
	wire [4-1:0] node53270;
	wire [4-1:0] node53273;
	wire [4-1:0] node53276;
	wire [4-1:0] node53277;
	wire [4-1:0] node53280;
	wire [4-1:0] node53283;
	wire [4-1:0] node53284;
	wire [4-1:0] node53285;
	wire [4-1:0] node53288;
	wire [4-1:0] node53291;
	wire [4-1:0] node53292;
	wire [4-1:0] node53295;
	wire [4-1:0] node53298;
	wire [4-1:0] node53299;
	wire [4-1:0] node53300;
	wire [4-1:0] node53301;
	wire [4-1:0] node53304;
	wire [4-1:0] node53307;
	wire [4-1:0] node53308;
	wire [4-1:0] node53309;
	wire [4-1:0] node53312;
	wire [4-1:0] node53315;
	wire [4-1:0] node53316;
	wire [4-1:0] node53319;
	wire [4-1:0] node53322;
	wire [4-1:0] node53323;
	wire [4-1:0] node53324;
	wire [4-1:0] node53327;
	wire [4-1:0] node53330;
	wire [4-1:0] node53331;
	wire [4-1:0] node53334;
	wire [4-1:0] node53337;
	wire [4-1:0] node53338;
	wire [4-1:0] node53339;
	wire [4-1:0] node53340;
	wire [4-1:0] node53344;
	wire [4-1:0] node53345;
	wire [4-1:0] node53349;
	wire [4-1:0] node53350;
	wire [4-1:0] node53351;
	wire [4-1:0] node53355;
	wire [4-1:0] node53357;
	wire [4-1:0] node53360;
	wire [4-1:0] node53361;
	wire [4-1:0] node53362;
	wire [4-1:0] node53363;
	wire [4-1:0] node53364;
	wire [4-1:0] node53367;
	wire [4-1:0] node53370;
	wire [4-1:0] node53371;
	wire [4-1:0] node53372;
	wire [4-1:0] node53373;
	wire [4-1:0] node53374;
	wire [4-1:0] node53375;
	wire [4-1:0] node53379;
	wire [4-1:0] node53380;
	wire [4-1:0] node53384;
	wire [4-1:0] node53385;
	wire [4-1:0] node53388;
	wire [4-1:0] node53391;
	wire [4-1:0] node53392;
	wire [4-1:0] node53395;
	wire [4-1:0] node53398;
	wire [4-1:0] node53399;
	wire [4-1:0] node53402;
	wire [4-1:0] node53405;
	wire [4-1:0] node53406;
	wire [4-1:0] node53407;
	wire [4-1:0] node53410;
	wire [4-1:0] node53413;
	wire [4-1:0] node53414;
	wire [4-1:0] node53415;
	wire [4-1:0] node53416;
	wire [4-1:0] node53419;
	wire [4-1:0] node53422;
	wire [4-1:0] node53423;
	wire [4-1:0] node53424;
	wire [4-1:0] node53427;
	wire [4-1:0] node53430;
	wire [4-1:0] node53431;
	wire [4-1:0] node53434;
	wire [4-1:0] node53437;
	wire [4-1:0] node53438;
	wire [4-1:0] node53439;
	wire [4-1:0] node53442;
	wire [4-1:0] node53445;
	wire [4-1:0] node53446;
	wire [4-1:0] node53447;
	wire [4-1:0] node53450;
	wire [4-1:0] node53453;
	wire [4-1:0] node53454;
	wire [4-1:0] node53457;
	wire [4-1:0] node53460;
	wire [4-1:0] node53461;
	wire [4-1:0] node53464;
	wire [4-1:0] node53467;
	wire [4-1:0] node53468;
	wire [4-1:0] node53469;
	wire [4-1:0] node53470;
	wire [4-1:0] node53471;
	wire [4-1:0] node53472;
	wire [4-1:0] node53473;
	wire [4-1:0] node53474;
	wire [4-1:0] node53477;
	wire [4-1:0] node53480;
	wire [4-1:0] node53481;
	wire [4-1:0] node53482;
	wire [4-1:0] node53483;
	wire [4-1:0] node53486;
	wire [4-1:0] node53490;
	wire [4-1:0] node53491;
	wire [4-1:0] node53492;
	wire [4-1:0] node53496;
	wire [4-1:0] node53498;
	wire [4-1:0] node53501;
	wire [4-1:0] node53502;
	wire [4-1:0] node53505;
	wire [4-1:0] node53508;
	wire [4-1:0] node53509;
	wire [4-1:0] node53510;
	wire [4-1:0] node53511;
	wire [4-1:0] node53512;
	wire [4-1:0] node53513;
	wire [4-1:0] node53517;
	wire [4-1:0] node53518;
	wire [4-1:0] node53521;
	wire [4-1:0] node53524;
	wire [4-1:0] node53525;
	wire [4-1:0] node53528;
	wire [4-1:0] node53531;
	wire [4-1:0] node53532;
	wire [4-1:0] node53533;
	wire [4-1:0] node53536;
	wire [4-1:0] node53539;
	wire [4-1:0] node53540;
	wire [4-1:0] node53541;
	wire [4-1:0] node53544;
	wire [4-1:0] node53547;
	wire [4-1:0] node53548;
	wire [4-1:0] node53551;
	wire [4-1:0] node53554;
	wire [4-1:0] node53555;
	wire [4-1:0] node53556;
	wire [4-1:0] node53557;
	wire [4-1:0] node53560;
	wire [4-1:0] node53563;
	wire [4-1:0] node53564;
	wire [4-1:0] node53567;
	wire [4-1:0] node53570;
	wire [4-1:0] node53571;
	wire [4-1:0] node53574;
	wire [4-1:0] node53577;
	wire [4-1:0] node53578;
	wire [4-1:0] node53579;
	wire [4-1:0] node53580;
	wire [4-1:0] node53581;
	wire [4-1:0] node53584;
	wire [4-1:0] node53587;
	wire [4-1:0] node53588;
	wire [4-1:0] node53589;
	wire [4-1:0] node53592;
	wire [4-1:0] node53595;
	wire [4-1:0] node53596;
	wire [4-1:0] node53599;
	wire [4-1:0] node53602;
	wire [4-1:0] node53603;
	wire [4-1:0] node53604;
	wire [4-1:0] node53605;
	wire [4-1:0] node53608;
	wire [4-1:0] node53611;
	wire [4-1:0] node53612;
	wire [4-1:0] node53615;
	wire [4-1:0] node53618;
	wire [4-1:0] node53619;
	wire [4-1:0] node53620;
	wire [4-1:0] node53623;
	wire [4-1:0] node53626;
	wire [4-1:0] node53627;
	wire [4-1:0] node53630;
	wire [4-1:0] node53633;
	wire [4-1:0] node53634;
	wire [4-1:0] node53635;
	wire [4-1:0] node53638;
	wire [4-1:0] node53641;
	wire [4-1:0] node53642;
	wire [4-1:0] node53643;
	wire [4-1:0] node53644;
	wire [4-1:0] node53646;
	wire [4-1:0] node53649;
	wire [4-1:0] node53650;
	wire [4-1:0] node53654;
	wire [4-1:0] node53655;
	wire [4-1:0] node53656;
	wire [4-1:0] node53659;
	wire [4-1:0] node53662;
	wire [4-1:0] node53663;
	wire [4-1:0] node53667;
	wire [4-1:0] node53668;
	wire [4-1:0] node53669;
	wire [4-1:0] node53670;
	wire [4-1:0] node53673;
	wire [4-1:0] node53676;
	wire [4-1:0] node53677;
	wire [4-1:0] node53680;
	wire [4-1:0] node53683;
	wire [4-1:0] node53684;
	wire [4-1:0] node53685;
	wire [4-1:0] node53688;
	wire [4-1:0] node53691;
	wire [4-1:0] node53692;
	wire [4-1:0] node53695;
	wire [4-1:0] node53698;
	wire [4-1:0] node53699;
	wire [4-1:0] node53702;
	wire [4-1:0] node53705;
	wire [4-1:0] node53706;
	wire [4-1:0] node53707;
	wire [4-1:0] node53711;
	wire [4-1:0] node53712;
	wire [4-1:0] node53716;
	wire [4-1:0] node53717;
	wire [4-1:0] node53718;
	wire [4-1:0] node53719;
	wire [4-1:0] node53720;
	wire [4-1:0] node53721;
	wire [4-1:0] node53722;
	wire [4-1:0] node53723;
	wire [4-1:0] node53724;
	wire [4-1:0] node53725;
	wire [4-1:0] node53728;
	wire [4-1:0] node53731;
	wire [4-1:0] node53732;
	wire [4-1:0] node53733;
	wire [4-1:0] node53736;
	wire [4-1:0] node53739;
	wire [4-1:0] node53740;
	wire [4-1:0] node53743;
	wire [4-1:0] node53746;
	wire [4-1:0] node53747;
	wire [4-1:0] node53748;
	wire [4-1:0] node53751;
	wire [4-1:0] node53754;
	wire [4-1:0] node53755;
	wire [4-1:0] node53758;
	wire [4-1:0] node53761;
	wire [4-1:0] node53762;
	wire [4-1:0] node53763;
	wire [4-1:0] node53766;
	wire [4-1:0] node53769;
	wire [4-1:0] node53770;
	wire [4-1:0] node53773;
	wire [4-1:0] node53777;
	wire [4-1:0] node53778;
	wire [4-1:0] node53779;
	wire [4-1:0] node53780;
	wire [4-1:0] node53783;
	wire [4-1:0] node53786;
	wire [4-1:0] node53787;
	wire [4-1:0] node53790;
	wire [4-1:0] node53794;
	wire [4-1:0] node53795;
	wire [4-1:0] node53796;
	wire [4-1:0] node53800;
	wire [4-1:0] node53801;
	wire [4-1:0] node53805;
	wire [4-1:0] node53806;
	wire [4-1:0] node53807;
	wire [4-1:0] node53808;
	wire [4-1:0] node53809;
	wire [4-1:0] node53813;
	wire [4-1:0] node53814;
	wire [4-1:0] node53819;
	wire [4-1:0] node53820;
	wire [4-1:0] node53821;
	wire [4-1:0] node53822;
	wire [4-1:0] node53826;
	wire [4-1:0] node53827;
	wire [4-1:0] node53832;
	wire [4-1:0] node53833;
	wire [4-1:0] node53834;
	wire [4-1:0] node53835;
	wire [4-1:0] node53839;
	wire [4-1:0] node53840;
	wire [4-1:0] node53844;
	wire [4-1:0] node53845;

	assign outp = (inp[14]) ? node28342 : node1;
		assign node1 = (inp[8]) ? node18103 : node2;
			assign node2 = (inp[3]) ? node8530 : node3;
				assign node3 = (inp[6]) ? node5683 : node4;
					assign node4 = (inp[11]) ? node2588 : node5;
						assign node5 = (inp[9]) ? node1279 : node6;
							assign node6 = (inp[10]) ? node652 : node7;
								assign node7 = (inp[13]) ? node327 : node8;
									assign node8 = (inp[2]) ? node182 : node9;
										assign node9 = (inp[5]) ? node95 : node10;
											assign node10 = (inp[0]) ? node48 : node11;
												assign node11 = (inp[7]) ? node25 : node12;
													assign node12 = (inp[12]) ? node20 : node13;
														assign node13 = (inp[15]) ? node15 : 4'b0000;
															assign node15 = (inp[4]) ? node17 : 4'b0000;
																assign node17 = (inp[1]) ? 4'b0110 : 4'b0010;
														assign node20 = (inp[4]) ? 4'b0000 : node21;
															assign node21 = (inp[1]) ? 4'b0011 : 4'b0010;
													assign node25 = (inp[12]) ? node35 : node26;
														assign node26 = (inp[4]) ? node30 : node27;
															assign node27 = (inp[15]) ? 4'b0110 : 4'b0010;
															assign node30 = (inp[15]) ? node32 : 4'b0010;
																assign node32 = (inp[1]) ? 4'b0001 : 4'b0000;
														assign node35 = (inp[15]) ? node41 : node36;
															assign node36 = (inp[1]) ? 4'b0000 : node37;
																assign node37 = (inp[4]) ? 4'b0100 : 4'b0000;
															assign node41 = (inp[4]) ? node45 : node42;
																assign node42 = (inp[1]) ? 4'b0000 : 4'b0100;
																assign node45 = (inp[1]) ? 4'b0110 : 4'b0111;
												assign node48 = (inp[15]) ? node68 : node49;
													assign node49 = (inp[12]) ? node53 : node50;
														assign node50 = (inp[7]) ? 4'b0010 : 4'b0000;
														assign node53 = (inp[7]) ? node61 : node54;
															assign node54 = (inp[1]) ? node58 : node55;
																assign node55 = (inp[4]) ? 4'b0110 : 4'b0010;
																assign node58 = (inp[4]) ? 4'b0111 : 4'b0011;
															assign node61 = (inp[1]) ? node65 : node62;
																assign node62 = (inp[4]) ? 4'b0101 : 4'b0001;
																assign node65 = (inp[4]) ? 4'b0000 : 4'b0100;
													assign node68 = (inp[7]) ? node84 : node69;
														assign node69 = (inp[1]) ? node77 : node70;
															assign node70 = (inp[12]) ? node74 : node71;
																assign node71 = (inp[4]) ? 4'b0010 : 4'b0000;
																assign node74 = (inp[4]) ? 4'b0001 : 4'b0010;
															assign node77 = (inp[12]) ? node81 : node78;
																assign node78 = (inp[4]) ? 4'b0111 : 4'b0001;
																assign node81 = (inp[4]) ? 4'b0000 : 4'b0010;
														assign node84 = (inp[12]) ? node90 : node85;
															assign node85 = (inp[4]) ? 4'b0001 : node86;
																assign node86 = (inp[1]) ? 4'b0111 : 4'b0110;
															assign node90 = (inp[4]) ? 4'b0111 : node91;
																assign node91 = (inp[1]) ? 4'b0001 : 4'b0101;
											assign node95 = (inp[1]) ? node139 : node96;
												assign node96 = (inp[0]) ? node114 : node97;
													assign node97 = (inp[7]) ? node101 : node98;
														assign node98 = (inp[4]) ? 4'b0110 : 4'b0010;
														assign node101 = (inp[12]) ? node107 : node102;
															assign node102 = (inp[4]) ? node104 : 4'b0111;
																assign node104 = (inp[15]) ? 4'b0000 : 4'b0011;
															assign node107 = (inp[4]) ? node111 : node108;
																assign node108 = (inp[15]) ? 4'b0000 : 4'b0101;
																assign node111 = (inp[15]) ? 4'b0110 : 4'b0000;
													assign node114 = (inp[4]) ? node124 : node115;
														assign node115 = (inp[7]) ? node119 : node116;
															assign node116 = (inp[12]) ? 4'b0010 : 4'b0000;
															assign node119 = (inp[12]) ? node121 : 4'b0111;
																assign node121 = (inp[15]) ? 4'b0000 : 4'b0100;
														assign node124 = (inp[12]) ? node132 : node125;
															assign node125 = (inp[7]) ? node129 : node126;
																assign node126 = (inp[15]) ? 4'b0111 : 4'b0001;
																assign node129 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node132 = (inp[15]) ? node136 : node133;
																assign node133 = (inp[7]) ? 4'b0001 : 4'b0111;
																assign node136 = (inp[7]) ? 4'b0111 : 4'b0001;
												assign node139 = (inp[7]) ? node159 : node140;
													assign node140 = (inp[12]) ? node152 : node141;
														assign node141 = (inp[15]) ? node147 : node142;
															assign node142 = (inp[4]) ? node144 : 4'b0100;
																assign node144 = (inp[0]) ? 4'b0101 : 4'b0100;
															assign node147 = (inp[4]) ? 4'b0111 : node148;
																assign node148 = (inp[0]) ? 4'b0101 : 4'b0100;
														assign node152 = (inp[4]) ? node154 : 4'b0111;
															assign node154 = (inp[15]) ? node156 : 4'b0010;
																assign node156 = (inp[0]) ? 4'b0101 : 4'b0100;
													assign node159 = (inp[15]) ? node171 : node160;
														assign node160 = (inp[12]) ? node166 : node161;
															assign node161 = (inp[4]) ? node163 : 4'b0111;
																assign node163 = (inp[0]) ? 4'b0110 : 4'b0111;
															assign node166 = (inp[4]) ? 4'b0000 : node167;
																assign node167 = (inp[0]) ? 4'b0101 : 4'b0100;
														assign node171 = (inp[4]) ? node177 : node172;
															assign node172 = (inp[12]) ? node174 : 4'b0010;
																assign node174 = (inp[0]) ? 4'b0000 : 4'b0001;
															assign node177 = (inp[12]) ? node179 : 4'b0101;
																assign node179 = (inp[0]) ? 4'b0011 : 4'b0010;
										assign node182 = (inp[1]) ? node248 : node183;
											assign node183 = (inp[7]) ? node207 : node184;
												assign node184 = (inp[4]) ? node188 : node185;
													assign node185 = (inp[12]) ? 4'b0110 : 4'b0100;
													assign node188 = (inp[5]) ? node198 : node189;
														assign node189 = (inp[12]) ? node193 : node190;
															assign node190 = (inp[15]) ? 4'b0111 : 4'b0101;
															assign node193 = (inp[15]) ? node195 : 4'b0011;
																assign node195 = (inp[0]) ? 4'b0100 : 4'b0101;
														assign node198 = (inp[15]) ? node204 : node199;
															assign node199 = (inp[12]) ? 4'b0010 : node200;
																assign node200 = (inp[0]) ? 4'b0100 : 4'b0101;
															assign node204 = (inp[12]) ? 4'b0100 : 4'b0010;
												assign node207 = (inp[12]) ? node231 : node208;
													assign node208 = (inp[4]) ? node220 : node209;
														assign node209 = (inp[15]) ? node213 : node210;
															assign node210 = (inp[0]) ? 4'b0110 : 4'b0111;
															assign node213 = (inp[0]) ? node217 : node214;
																assign node214 = (inp[5]) ? 4'b0011 : 4'b0010;
																assign node217 = (inp[5]) ? 4'b0010 : 4'b0011;
														assign node220 = (inp[15]) ? node226 : node221;
															assign node221 = (inp[0]) ? 4'b0111 : node222;
																assign node222 = (inp[5]) ? 4'b0110 : 4'b0111;
															assign node226 = (inp[5]) ? 4'b0101 : node227;
																assign node227 = (inp[0]) ? 4'b0100 : 4'b0101;
													assign node231 = (inp[4]) ? node241 : node232;
														assign node232 = (inp[5]) ? node238 : node233;
															assign node233 = (inp[15]) ? 4'b0001 : node234;
																assign node234 = (inp[0]) ? 4'b0101 : 4'b0100;
															assign node238 = (inp[15]) ? 4'b0100 : 4'b0000;
														assign node241 = (inp[15]) ? node245 : node242;
															assign node242 = (inp[5]) ? 4'b0100 : 4'b0000;
															assign node245 = (inp[0]) ? 4'b0011 : 4'b0010;
											assign node248 = (inp[5]) ? node286 : node249;
												assign node249 = (inp[15]) ? node267 : node250;
													assign node250 = (inp[12]) ? node258 : node251;
														assign node251 = (inp[4]) ? node255 : node252;
															assign node252 = (inp[7]) ? 4'b0110 : 4'b0100;
															assign node255 = (inp[7]) ? 4'b0111 : 4'b0101;
														assign node258 = (inp[7]) ? node264 : node259;
															assign node259 = (inp[4]) ? node261 : 4'b0111;
																assign node261 = (inp[0]) ? 4'b0011 : 4'b0010;
															assign node264 = (inp[4]) ? 4'b0101 : 4'b0000;
													assign node267 = (inp[4]) ? node279 : node268;
														assign node268 = (inp[12]) ? node274 : node269;
															assign node269 = (inp[7]) ? 4'b0011 : node270;
																assign node270 = (inp[0]) ? 4'b0101 : 4'b0100;
															assign node274 = (inp[7]) ? node276 : 4'b0110;
																assign node276 = (inp[0]) ? 4'b0101 : 4'b0100;
														assign node279 = (inp[7]) ? node283 : node280;
															assign node280 = (inp[12]) ? 4'b0101 : 4'b0010;
															assign node283 = (inp[12]) ? 4'b0010 : 4'b0100;
												assign node286 = (inp[12]) ? node306 : node287;
													assign node287 = (inp[0]) ? node295 : node288;
														assign node288 = (inp[7]) ? node292 : node289;
															assign node289 = (inp[15]) ? 4'b0010 : 4'b0000;
															assign node292 = (inp[15]) ? 4'b0000 : 4'b0011;
														assign node295 = (inp[7]) ? node299 : node296;
															assign node296 = (inp[4]) ? 4'b0011 : 4'b0001;
															assign node299 = (inp[4]) ? node303 : node300;
																assign node300 = (inp[15]) ? 4'b0110 : 4'b0010;
																assign node303 = (inp[15]) ? 4'b0000 : 4'b0011;
													assign node306 = (inp[7]) ? node316 : node307;
														assign node307 = (inp[15]) ? node313 : node308;
															assign node308 = (inp[4]) ? 4'b0111 : node309;
																assign node309 = (inp[0]) ? 4'b0010 : 4'b0011;
															assign node313 = (inp[4]) ? 4'b0000 : 4'b0010;
														assign node316 = (inp[4]) ? node322 : node317;
															assign node317 = (inp[15]) ? node319 : 4'b0001;
																assign node319 = (inp[0]) ? 4'b0100 : 4'b0101;
															assign node322 = (inp[15]) ? node324 : 4'b0100;
																assign node324 = (inp[0]) ? 4'b0110 : 4'b0111;
									assign node327 = (inp[2]) ? node483 : node328;
										assign node328 = (inp[5]) ? node390 : node329;
											assign node329 = (inp[12]) ? node353 : node330;
												assign node330 = (inp[15]) ? node334 : node331;
													assign node331 = (inp[7]) ? 4'b0110 : 4'b0100;
													assign node334 = (inp[1]) ? node346 : node335;
														assign node335 = (inp[7]) ? node339 : node336;
															assign node336 = (inp[4]) ? 4'b0111 : 4'b0101;
															assign node339 = (inp[4]) ? node343 : node340;
																assign node340 = (inp[0]) ? 4'b0010 : 4'b0011;
																assign node343 = (inp[0]) ? 4'b0100 : 4'b0101;
														assign node346 = (inp[7]) ? node350 : node347;
															assign node347 = (inp[4]) ? 4'b0010 : 4'b0100;
															assign node350 = (inp[4]) ? 4'b0100 : 4'b0010;
												assign node353 = (inp[7]) ? node373 : node354;
													assign node354 = (inp[15]) ? node366 : node355;
														assign node355 = (inp[4]) ? node359 : node356;
															assign node356 = (inp[1]) ? 4'b0111 : 4'b0110;
															assign node359 = (inp[1]) ? node363 : node360;
																assign node360 = (inp[0]) ? 4'b0011 : 4'b0010;
																assign node363 = (inp[0]) ? 4'b0010 : 4'b0011;
														assign node366 = (inp[4]) ? node368 : 4'b0111;
															assign node368 = (inp[0]) ? node370 : 4'b0101;
																assign node370 = (inp[1]) ? 4'b0101 : 4'b0100;
													assign node373 = (inp[15]) ? node381 : node374;
														assign node374 = (inp[1]) ? node378 : node375;
															assign node375 = (inp[4]) ? 4'b0001 : 4'b0101;
															assign node378 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node381 = (inp[4]) ? node385 : node382;
															assign node382 = (inp[1]) ? 4'b0101 : 4'b0000;
															assign node385 = (inp[1]) ? 4'b0010 : node386;
																assign node386 = (inp[0]) ? 4'b0011 : 4'b0010;
											assign node390 = (inp[1]) ? node440 : node391;
												assign node391 = (inp[0]) ? node411 : node392;
													assign node392 = (inp[7]) ? node400 : node393;
														assign node393 = (inp[12]) ? node397 : node394;
															assign node394 = (inp[15]) ? 4'b0101 : 4'b0100;
															assign node397 = (inp[15]) ? 4'b0100 : 4'b0011;
														assign node400 = (inp[12]) ? node404 : node401;
															assign node401 = (inp[15]) ? 4'b0010 : 4'b0111;
															assign node404 = (inp[15]) ? node408 : node405;
																assign node405 = (inp[4]) ? 4'b0100 : 4'b0000;
																assign node408 = (inp[4]) ? 4'b0010 : 4'b0101;
													assign node411 = (inp[4]) ? node427 : node412;
														assign node412 = (inp[15]) ? node420 : node413;
															assign node413 = (inp[12]) ? node417 : node414;
																assign node414 = (inp[7]) ? 4'b0111 : 4'b0100;
																assign node417 = (inp[7]) ? 4'b0000 : 4'b0110;
															assign node420 = (inp[7]) ? node424 : node421;
																assign node421 = (inp[12]) ? 4'b0111 : 4'b0101;
																assign node424 = (inp[12]) ? 4'b0101 : 4'b0011;
														assign node427 = (inp[7]) ? node433 : node428;
															assign node428 = (inp[15]) ? node430 : 4'b0011;
																assign node430 = (inp[12]) ? 4'b0100 : 4'b0010;
															assign node433 = (inp[12]) ? node437 : node434;
																assign node434 = (inp[15]) ? 4'b0101 : 4'b0110;
																assign node437 = (inp[15]) ? 4'b0010 : 4'b0101;
												assign node440 = (inp[7]) ? node462 : node441;
													assign node441 = (inp[12]) ? node453 : node442;
														assign node442 = (inp[4]) ? node448 : node443;
															assign node443 = (inp[0]) ? node445 : 4'b0000;
																assign node445 = (inp[15]) ? 4'b0000 : 4'b0001;
															assign node448 = (inp[15]) ? node450 : 4'b0001;
																assign node450 = (inp[0]) ? 4'b0011 : 4'b0010;
														assign node453 = (inp[4]) ? node459 : node454;
															assign node454 = (inp[0]) ? node456 : 4'b0011;
																assign node456 = (inp[15]) ? 4'b0011 : 4'b0010;
															assign node459 = (inp[15]) ? 4'b0000 : 4'b0110;
													assign node462 = (inp[12]) ? node470 : node463;
														assign node463 = (inp[4]) ? 4'b0000 : node464;
															assign node464 = (inp[15]) ? 4'b0111 : node465;
																assign node465 = (inp[0]) ? 4'b0010 : 4'b0011;
														assign node470 = (inp[15]) ? node476 : node471;
															assign node471 = (inp[4]) ? node473 : 4'b0001;
																assign node473 = (inp[0]) ? 4'b0100 : 4'b0101;
															assign node476 = (inp[4]) ? node480 : node477;
																assign node477 = (inp[0]) ? 4'b0101 : 4'b0100;
																assign node480 = (inp[0]) ? 4'b0110 : 4'b0111;
										assign node483 = (inp[5]) ? node565 : node484;
											assign node484 = (inp[12]) ? node524 : node485;
												assign node485 = (inp[7]) ? node499 : node486;
													assign node486 = (inp[4]) ? node492 : node487;
														assign node487 = (inp[15]) ? 4'b0000 : node488;
															assign node488 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node492 = (inp[15]) ? node496 : node493;
															assign node493 = (inp[0]) ? 4'b0000 : 4'b0001;
															assign node496 = (inp[1]) ? 4'b0111 : 4'b0010;
													assign node499 = (inp[15]) ? node515 : node500;
														assign node500 = (inp[1]) ? node508 : node501;
															assign node501 = (inp[4]) ? node505 : node502;
																assign node502 = (inp[0]) ? 4'b0011 : 4'b0010;
																assign node505 = (inp[0]) ? 4'b0010 : 4'b0011;
															assign node508 = (inp[4]) ? node512 : node509;
																assign node509 = (inp[0]) ? 4'b0011 : 4'b0010;
																assign node512 = (inp[0]) ? 4'b0010 : 4'b0011;
														assign node515 = (inp[4]) ? node519 : node516;
															assign node516 = (inp[1]) ? 4'b0110 : 4'b0111;
															assign node519 = (inp[1]) ? node521 : 4'b0001;
																assign node521 = (inp[0]) ? 4'b0000 : 4'b0001;
												assign node524 = (inp[7]) ? node546 : node525;
													assign node525 = (inp[15]) ? node541 : node526;
														assign node526 = (inp[4]) ? node534 : node527;
															assign node527 = (inp[1]) ? node531 : node528;
																assign node528 = (inp[0]) ? 4'b0011 : 4'b0010;
																assign node531 = (inp[0]) ? 4'b0010 : 4'b0011;
															assign node534 = (inp[0]) ? node538 : node535;
																assign node535 = (inp[1]) ? 4'b0110 : 4'b0111;
																assign node538 = (inp[1]) ? 4'b0111 : 4'b0110;
														assign node541 = (inp[4]) ? node543 : 4'b0011;
															assign node543 = (inp[1]) ? 4'b0000 : 4'b0001;
													assign node546 = (inp[4]) ? node556 : node547;
														assign node547 = (inp[0]) ? node553 : node548;
															assign node548 = (inp[15]) ? node550 : 4'b0100;
																assign node550 = (inp[1]) ? 4'b0000 : 4'b0100;
															assign node553 = (inp[1]) ? 4'b0000 : 4'b0001;
														assign node556 = (inp[15]) ? node562 : node557;
															assign node557 = (inp[1]) ? node559 : 4'b0100;
																assign node559 = (inp[0]) ? 4'b0000 : 4'b0001;
															assign node562 = (inp[0]) ? 4'b0110 : 4'b0111;
											assign node565 = (inp[1]) ? node609 : node566;
												assign node566 = (inp[15]) ? node584 : node567;
													assign node567 = (inp[12]) ? node575 : node568;
														assign node568 = (inp[7]) ? 4'b0011 : node569;
															assign node569 = (inp[4]) ? 4'b0000 : node570;
																assign node570 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node575 = (inp[7]) ? node581 : node576;
															assign node576 = (inp[4]) ? 4'b0110 : node577;
																assign node577 = (inp[0]) ? 4'b0011 : 4'b0010;
															assign node581 = (inp[4]) ? 4'b0000 : 4'b0100;
													assign node584 = (inp[4]) ? node596 : node585;
														assign node585 = (inp[12]) ? node591 : node586;
															assign node586 = (inp[7]) ? node588 : 4'b0000;
																assign node588 = (inp[0]) ? 4'b0111 : 4'b0110;
															assign node591 = (inp[7]) ? node593 : 4'b0010;
																assign node593 = (inp[0]) ? 4'b0000 : 4'b0001;
														assign node596 = (inp[0]) ? node604 : node597;
															assign node597 = (inp[12]) ? node601 : node598;
																assign node598 = (inp[7]) ? 4'b0000 : 4'b0111;
																assign node601 = (inp[7]) ? 4'b0111 : 4'b0001;
															assign node604 = (inp[7]) ? node606 : 4'b0111;
																assign node606 = (inp[12]) ? 4'b0111 : 4'b0001;
												assign node609 = (inp[7]) ? node633 : node610;
													assign node610 = (inp[12]) ? node622 : node611;
														assign node611 = (inp[4]) ? node617 : node612;
															assign node612 = (inp[15]) ? 4'b0100 : node613;
																assign node613 = (inp[0]) ? 4'b0101 : 4'b0100;
															assign node617 = (inp[15]) ? node619 : 4'b0100;
																assign node619 = (inp[0]) ? 4'b0110 : 4'b0111;
														assign node622 = (inp[15]) ? node630 : node623;
															assign node623 = (inp[0]) ? node627 : node624;
																assign node624 = (inp[4]) ? 4'b0011 : 4'b0111;
																assign node627 = (inp[4]) ? 4'b0010 : 4'b0110;
															assign node630 = (inp[4]) ? 4'b0101 : 4'b0111;
													assign node633 = (inp[12]) ? node645 : node634;
														assign node634 = (inp[4]) ? node642 : node635;
															assign node635 = (inp[0]) ? node639 : node636;
																assign node636 = (inp[15]) ? 4'b0011 : 4'b0111;
																assign node639 = (inp[15]) ? 4'b0010 : 4'b0110;
															assign node642 = (inp[15]) ? 4'b0101 : 4'b0111;
														assign node645 = (inp[4]) ? node649 : node646;
															assign node646 = (inp[15]) ? 4'b0001 : 4'b0101;
															assign node649 = (inp[15]) ? 4'b0011 : 4'b0001;
								assign node652 = (inp[13]) ? node960 : node653;
									assign node653 = (inp[2]) ? node815 : node654;
										assign node654 = (inp[5]) ? node728 : node655;
											assign node655 = (inp[12]) ? node683 : node656;
												assign node656 = (inp[7]) ? node670 : node657;
													assign node657 = (inp[15]) ? node659 : 4'b0001;
														assign node659 = (inp[4]) ? node665 : node660;
															assign node660 = (inp[1]) ? node662 : 4'b0001;
																assign node662 = (inp[0]) ? 4'b0000 : 4'b0001;
															assign node665 = (inp[1]) ? node667 : 4'b0011;
																assign node667 = (inp[0]) ? 4'b0110 : 4'b0111;
													assign node670 = (inp[15]) ? node672 : 4'b0011;
														assign node672 = (inp[4]) ? node678 : node673;
															assign node673 = (inp[1]) ? node675 : 4'b0111;
																assign node675 = (inp[0]) ? 4'b0110 : 4'b0111;
															assign node678 = (inp[0]) ? 4'b0000 : node679;
																assign node679 = (inp[1]) ? 4'b0000 : 4'b0001;
												assign node683 = (inp[7]) ? node701 : node684;
													assign node684 = (inp[15]) ? node692 : node685;
														assign node685 = (inp[1]) ? node689 : node686;
															assign node686 = (inp[4]) ? 4'b0111 : 4'b0011;
															assign node689 = (inp[4]) ? 4'b0110 : 4'b0010;
														assign node692 = (inp[4]) ? node696 : node693;
															assign node693 = (inp[0]) ? 4'b0011 : 4'b0010;
															assign node696 = (inp[1]) ? 4'b0001 : node697;
																assign node697 = (inp[0]) ? 4'b0000 : 4'b0001;
													assign node701 = (inp[15]) ? node715 : node702;
														assign node702 = (inp[0]) ? node710 : node703;
															assign node703 = (inp[4]) ? node707 : node704;
																assign node704 = (inp[1]) ? 4'b0100 : 4'b0001;
																assign node707 = (inp[1]) ? 4'b0001 : 4'b0101;
															assign node710 = (inp[1]) ? 4'b0001 : node711;
																assign node711 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node715 = (inp[4]) ? node723 : node716;
															assign node716 = (inp[0]) ? node720 : node717;
																assign node717 = (inp[1]) ? 4'b0001 : 4'b0101;
																assign node720 = (inp[1]) ? 4'b0000 : 4'b0100;
															assign node723 = (inp[0]) ? 4'b0110 : node724;
																assign node724 = (inp[1]) ? 4'b0111 : 4'b0110;
											assign node728 = (inp[1]) ? node772 : node729;
												assign node729 = (inp[12]) ? node749 : node730;
													assign node730 = (inp[15]) ? node740 : node731;
														assign node731 = (inp[7]) ? node735 : node732;
															assign node732 = (inp[4]) ? 4'b0000 : 4'b0001;
															assign node735 = (inp[0]) ? node737 : 4'b0010;
																assign node737 = (inp[4]) ? 4'b0011 : 4'b0010;
														assign node740 = (inp[4]) ? node744 : node741;
															assign node741 = (inp[7]) ? 4'b0110 : 4'b0001;
															assign node744 = (inp[7]) ? 4'b0001 : node745;
																assign node745 = (inp[0]) ? 4'b0110 : 4'b0111;
													assign node749 = (inp[4]) ? node757 : node750;
														assign node750 = (inp[7]) ? node752 : 4'b0011;
															assign node752 = (inp[15]) ? 4'b0001 : node753;
																assign node753 = (inp[0]) ? 4'b0101 : 4'b0100;
														assign node757 = (inp[0]) ? node765 : node758;
															assign node758 = (inp[15]) ? node762 : node759;
																assign node759 = (inp[7]) ? 4'b0001 : 4'b0111;
																assign node762 = (inp[7]) ? 4'b0111 : 4'b0000;
															assign node765 = (inp[7]) ? node769 : node766;
																assign node766 = (inp[15]) ? 4'b0000 : 4'b0110;
																assign node769 = (inp[15]) ? 4'b0110 : 4'b0000;
												assign node772 = (inp[12]) ? node796 : node773;
													assign node773 = (inp[7]) ? node785 : node774;
														assign node774 = (inp[4]) ? node780 : node775;
															assign node775 = (inp[15]) ? node777 : 4'b0101;
																assign node777 = (inp[0]) ? 4'b0100 : 4'b0101;
															assign node780 = (inp[15]) ? 4'b0110 : node781;
																assign node781 = (inp[0]) ? 4'b0100 : 4'b0101;
														assign node785 = (inp[15]) ? node791 : node786;
															assign node786 = (inp[4]) ? node788 : 4'b0110;
																assign node788 = (inp[0]) ? 4'b0111 : 4'b0110;
															assign node791 = (inp[4]) ? node793 : 4'b0011;
																assign node793 = (inp[0]) ? 4'b0100 : 4'b0101;
													assign node796 = (inp[4]) ? node804 : node797;
														assign node797 = (inp[7]) ? node799 : 4'b0110;
															assign node799 = (inp[15]) ? 4'b0000 : node800;
																assign node800 = (inp[0]) ? 4'b0100 : 4'b0101;
														assign node804 = (inp[15]) ? node810 : node805;
															assign node805 = (inp[7]) ? node807 : 4'b0011;
																assign node807 = (inp[0]) ? 4'b0001 : 4'b0000;
															assign node810 = (inp[7]) ? 4'b0011 : node811;
																assign node811 = (inp[0]) ? 4'b0100 : 4'b0101;
										assign node815 = (inp[5]) ? node883 : node816;
											assign node816 = (inp[12]) ? node846 : node817;
												assign node817 = (inp[7]) ? node831 : node818;
													assign node818 = (inp[4]) ? node826 : node819;
														assign node819 = (inp[0]) ? node821 : 4'b0101;
															assign node821 = (inp[15]) ? node823 : 4'b0101;
																assign node823 = (inp[1]) ? 4'b0100 : 4'b0101;
														assign node826 = (inp[15]) ? node828 : 4'b0100;
															assign node828 = (inp[1]) ? 4'b0011 : 4'b0110;
													assign node831 = (inp[4]) ? node839 : node832;
														assign node832 = (inp[15]) ? node834 : 4'b0111;
															assign node834 = (inp[0]) ? 4'b0010 : node835;
																assign node835 = (inp[1]) ? 4'b0010 : 4'b0011;
														assign node839 = (inp[15]) ? node841 : 4'b0110;
															assign node841 = (inp[0]) ? 4'b0101 : node842;
																assign node842 = (inp[1]) ? 4'b0101 : 4'b0100;
												assign node846 = (inp[7]) ? node866 : node847;
													assign node847 = (inp[4]) ? node855 : node848;
														assign node848 = (inp[1]) ? node850 : 4'b0111;
															assign node850 = (inp[15]) ? node852 : 4'b0110;
																assign node852 = (inp[0]) ? 4'b0111 : 4'b0110;
														assign node855 = (inp[15]) ? node863 : node856;
															assign node856 = (inp[0]) ? node860 : node857;
																assign node857 = (inp[1]) ? 4'b0011 : 4'b0010;
																assign node860 = (inp[1]) ? 4'b0010 : 4'b0011;
															assign node863 = (inp[0]) ? 4'b0101 : 4'b0100;
													assign node866 = (inp[15]) ? node874 : node867;
														assign node867 = (inp[1]) ? node871 : node868;
															assign node868 = (inp[4]) ? 4'b0001 : 4'b0101;
															assign node871 = (inp[4]) ? 4'b0100 : 4'b0001;
														assign node874 = (inp[4]) ? node878 : node875;
															assign node875 = (inp[0]) ? 4'b0100 : 4'b0000;
															assign node878 = (inp[1]) ? 4'b0011 : node879;
																assign node879 = (inp[0]) ? 4'b0010 : 4'b0011;
											assign node883 = (inp[1]) ? node923 : node884;
												assign node884 = (inp[12]) ? node906 : node885;
													assign node885 = (inp[7]) ? node895 : node886;
														assign node886 = (inp[15]) ? node892 : node887;
															assign node887 = (inp[0]) ? 4'b0101 : node888;
																assign node888 = (inp[4]) ? 4'b0100 : 4'b0101;
															assign node892 = (inp[4]) ? 4'b0011 : 4'b0101;
														assign node895 = (inp[4]) ? node901 : node896;
															assign node896 = (inp[0]) ? 4'b0011 : node897;
																assign node897 = (inp[15]) ? 4'b0010 : 4'b0110;
															assign node901 = (inp[15]) ? 4'b0100 : node902;
																assign node902 = (inp[0]) ? 4'b0110 : 4'b0111;
													assign node906 = (inp[7]) ? node914 : node907;
														assign node907 = (inp[15]) ? node911 : node908;
															assign node908 = (inp[4]) ? 4'b0011 : 4'b0111;
															assign node911 = (inp[4]) ? 4'b0101 : 4'b0111;
														assign node914 = (inp[4]) ? node918 : node915;
															assign node915 = (inp[15]) ? 4'b0101 : 4'b0001;
															assign node918 = (inp[15]) ? 4'b0011 : node919;
																assign node919 = (inp[0]) ? 4'b0101 : 4'b0100;
												assign node923 = (inp[15]) ? node945 : node924;
													assign node924 = (inp[12]) ? node936 : node925;
														assign node925 = (inp[7]) ? node931 : node926;
															assign node926 = (inp[0]) ? node928 : 4'b0001;
																assign node928 = (inp[4]) ? 4'b0001 : 4'b0000;
															assign node931 = (inp[4]) ? 4'b0010 : node932;
																assign node932 = (inp[0]) ? 4'b0011 : 4'b0010;
														assign node936 = (inp[7]) ? node942 : node937;
															assign node937 = (inp[4]) ? 4'b0110 : node938;
																assign node938 = (inp[0]) ? 4'b0011 : 4'b0010;
															assign node942 = (inp[4]) ? 4'b0100 : 4'b0000;
													assign node945 = (inp[7]) ? node951 : node946;
														assign node946 = (inp[12]) ? node948 : 4'b0000;
															assign node948 = (inp[4]) ? 4'b0001 : 4'b0011;
														assign node951 = (inp[12]) ? node955 : node952;
															assign node952 = (inp[4]) ? 4'b0001 : 4'b0111;
															assign node955 = (inp[0]) ? node957 : 4'b0100;
																assign node957 = (inp[4]) ? 4'b0111 : 4'b0101;
									assign node960 = (inp[2]) ? node1104 : node961;
										assign node961 = (inp[5]) ? node1025 : node962;
											assign node962 = (inp[7]) ? node992 : node963;
												assign node963 = (inp[12]) ? node971 : node964;
													assign node964 = (inp[15]) ? node966 : 4'b0101;
														assign node966 = (inp[4]) ? node968 : 4'b0100;
															assign node968 = (inp[1]) ? 4'b0011 : 4'b0110;
													assign node971 = (inp[4]) ? node981 : node972;
														assign node972 = (inp[0]) ? 4'b0110 : node973;
															assign node973 = (inp[1]) ? node977 : node974;
																assign node974 = (inp[15]) ? 4'b0110 : 4'b0111;
																assign node977 = (inp[15]) ? 4'b0111 : 4'b0110;
														assign node981 = (inp[15]) ? node987 : node982;
															assign node982 = (inp[1]) ? 4'b0010 : node983;
																assign node983 = (inp[0]) ? 4'b0010 : 4'b0011;
															assign node987 = (inp[1]) ? 4'b0100 : node988;
																assign node988 = (inp[0]) ? 4'b0101 : 4'b0100;
												assign node992 = (inp[12]) ? node1004 : node993;
													assign node993 = (inp[15]) ? node995 : 4'b0111;
														assign node995 = (inp[4]) ? node1001 : node996;
															assign node996 = (inp[0]) ? 4'b0011 : node997;
																assign node997 = (inp[1]) ? 4'b0011 : 4'b0010;
															assign node1001 = (inp[0]) ? 4'b0101 : 4'b0100;
													assign node1004 = (inp[4]) ? node1016 : node1005;
														assign node1005 = (inp[15]) ? node1011 : node1006;
															assign node1006 = (inp[1]) ? 4'b0001 : node1007;
																assign node1007 = (inp[0]) ? 4'b0100 : 4'b0101;
															assign node1011 = (inp[1]) ? node1013 : 4'b0001;
																assign node1013 = (inp[0]) ? 4'b0101 : 4'b0100;
														assign node1016 = (inp[15]) ? node1020 : node1017;
															assign node1017 = (inp[1]) ? 4'b0101 : 4'b0000;
															assign node1020 = (inp[0]) ? node1022 : 4'b0011;
																assign node1022 = (inp[1]) ? 4'b0011 : 4'b0010;
											assign node1025 = (inp[1]) ? node1061 : node1026;
												assign node1026 = (inp[12]) ? node1046 : node1027;
													assign node1027 = (inp[7]) ? node1037 : node1028;
														assign node1028 = (inp[15]) ? node1034 : node1029;
															assign node1029 = (inp[4]) ? node1031 : 4'b0101;
																assign node1031 = (inp[0]) ? 4'b0100 : 4'b0101;
															assign node1034 = (inp[4]) ? 4'b0011 : 4'b0100;
														assign node1037 = (inp[4]) ? node1043 : node1038;
															assign node1038 = (inp[15]) ? node1040 : 4'b0110;
																assign node1040 = (inp[0]) ? 4'b0010 : 4'b0011;
															assign node1043 = (inp[15]) ? 4'b0100 : 4'b0110;
													assign node1046 = (inp[7]) ? node1054 : node1047;
														assign node1047 = (inp[15]) ? node1051 : node1048;
															assign node1048 = (inp[4]) ? 4'b0010 : 4'b0111;
															assign node1051 = (inp[4]) ? 4'b0101 : 4'b0110;
														assign node1054 = (inp[4]) ? node1058 : node1055;
															assign node1055 = (inp[15]) ? 4'b0100 : 4'b0001;
															assign node1058 = (inp[15]) ? 4'b0011 : 4'b0101;
												assign node1061 = (inp[12]) ? node1083 : node1062;
													assign node1062 = (inp[7]) ? node1074 : node1063;
														assign node1063 = (inp[15]) ? node1069 : node1064;
															assign node1064 = (inp[4]) ? 4'b0000 : node1065;
																assign node1065 = (inp[0]) ? 4'b0000 : 4'b0001;
															assign node1069 = (inp[4]) ? node1071 : 4'b0001;
																assign node1071 = (inp[0]) ? 4'b0010 : 4'b0011;
														assign node1074 = (inp[4]) ? node1080 : node1075;
															assign node1075 = (inp[15]) ? 4'b0110 : node1076;
																assign node1076 = (inp[0]) ? 4'b0011 : 4'b0010;
															assign node1080 = (inp[15]) ? 4'b0001 : 4'b0011;
													assign node1083 = (inp[7]) ? node1093 : node1084;
														assign node1084 = (inp[4]) ? node1090 : node1085;
															assign node1085 = (inp[0]) ? node1087 : 4'b0010;
																assign node1087 = (inp[15]) ? 4'b0010 : 4'b0011;
															assign node1090 = (inp[15]) ? 4'b0001 : 4'b0111;
														assign node1093 = (inp[4]) ? node1099 : node1094;
															assign node1094 = (inp[15]) ? node1096 : 4'b0000;
																assign node1096 = (inp[0]) ? 4'b0100 : 4'b0101;
															assign node1099 = (inp[0]) ? 4'b0101 : node1100;
																assign node1100 = (inp[15]) ? 4'b0110 : 4'b0100;
										assign node1104 = (inp[5]) ? node1190 : node1105;
											assign node1105 = (inp[7]) ? node1151 : node1106;
												assign node1106 = (inp[12]) ? node1126 : node1107;
													assign node1107 = (inp[4]) ? node1117 : node1108;
														assign node1108 = (inp[0]) ? node1114 : node1109;
															assign node1109 = (inp[15]) ? node1111 : 4'b0001;
																assign node1111 = (inp[1]) ? 4'b0001 : 4'b0000;
															assign node1114 = (inp[15]) ? 4'b0001 : 4'b0000;
														assign node1117 = (inp[15]) ? node1121 : node1118;
															assign node1118 = (inp[0]) ? 4'b0001 : 4'b0000;
															assign node1121 = (inp[0]) ? node1123 : 4'b0011;
																assign node1123 = (inp[1]) ? 4'b0110 : 4'b0010;
													assign node1126 = (inp[4]) ? node1140 : node1127;
														assign node1127 = (inp[1]) ? node1135 : node1128;
															assign node1128 = (inp[0]) ? node1132 : node1129;
																assign node1129 = (inp[15]) ? 4'b0010 : 4'b0011;
																assign node1132 = (inp[15]) ? 4'b0011 : 4'b0010;
															assign node1135 = (inp[15]) ? 4'b0010 : node1136;
																assign node1136 = (inp[0]) ? 4'b0011 : 4'b0010;
														assign node1140 = (inp[15]) ? node1146 : node1141;
															assign node1141 = (inp[1]) ? 4'b0110 : node1142;
																assign node1142 = (inp[0]) ? 4'b0111 : 4'b0110;
															assign node1146 = (inp[1]) ? node1148 : 4'b0000;
																assign node1148 = (inp[0]) ? 4'b0000 : 4'b0001;
												assign node1151 = (inp[12]) ? node1171 : node1152;
													assign node1152 = (inp[4]) ? node1162 : node1153;
														assign node1153 = (inp[15]) ? node1157 : node1154;
															assign node1154 = (inp[0]) ? 4'b0010 : 4'b0011;
															assign node1157 = (inp[0]) ? 4'b0111 : node1158;
																assign node1158 = (inp[1]) ? 4'b0111 : 4'b0110;
														assign node1162 = (inp[15]) ? node1166 : node1163;
															assign node1163 = (inp[0]) ? 4'b0011 : 4'b0010;
															assign node1166 = (inp[1]) ? node1168 : 4'b0000;
																assign node1168 = (inp[0]) ? 4'b0001 : 4'b0000;
													assign node1171 = (inp[4]) ? node1179 : node1172;
														assign node1172 = (inp[15]) ? node1176 : node1173;
															assign node1173 = (inp[1]) ? 4'b0101 : 4'b0000;
															assign node1176 = (inp[1]) ? 4'b0001 : 4'b0101;
														assign node1179 = (inp[15]) ? node1185 : node1180;
															assign node1180 = (inp[1]) ? node1182 : 4'b0101;
																assign node1182 = (inp[0]) ? 4'b0001 : 4'b0000;
															assign node1185 = (inp[1]) ? 4'b0110 : node1186;
																assign node1186 = (inp[0]) ? 4'b0111 : 4'b0110;
											assign node1190 = (inp[1]) ? node1238 : node1191;
												assign node1191 = (inp[15]) ? node1213 : node1192;
													assign node1192 = (inp[12]) ? node1204 : node1193;
														assign node1193 = (inp[7]) ? node1199 : node1194;
															assign node1194 = (inp[4]) ? 4'b0001 : node1195;
																assign node1195 = (inp[0]) ? 4'b0000 : 4'b0001;
															assign node1199 = (inp[4]) ? 4'b0010 : node1200;
																assign node1200 = (inp[0]) ? 4'b0011 : 4'b0010;
														assign node1204 = (inp[7]) ? node1210 : node1205;
															assign node1205 = (inp[4]) ? 4'b0111 : node1206;
																assign node1206 = (inp[0]) ? 4'b0010 : 4'b0011;
															assign node1210 = (inp[4]) ? 4'b0001 : 4'b0101;
													assign node1213 = (inp[7]) ? node1227 : node1214;
														assign node1214 = (inp[0]) ? node1220 : node1215;
															assign node1215 = (inp[12]) ? node1217 : 4'b0000;
																assign node1217 = (inp[4]) ? 4'b0000 : 4'b0010;
															assign node1220 = (inp[4]) ? node1224 : node1221;
																assign node1221 = (inp[12]) ? 4'b0011 : 4'b0001;
																assign node1224 = (inp[12]) ? 4'b0001 : 4'b0110;
														assign node1227 = (inp[4]) ? node1235 : node1228;
															assign node1228 = (inp[12]) ? node1232 : node1229;
																assign node1229 = (inp[0]) ? 4'b0110 : 4'b0111;
																assign node1232 = (inp[0]) ? 4'b0001 : 4'b0000;
															assign node1235 = (inp[12]) ? 4'b0110 : 4'b0000;
												assign node1238 = (inp[12]) ? node1260 : node1239;
													assign node1239 = (inp[7]) ? node1251 : node1240;
														assign node1240 = (inp[4]) ? node1246 : node1241;
															assign node1241 = (inp[0]) ? node1243 : 4'b0101;
																assign node1243 = (inp[15]) ? 4'b0101 : 4'b0100;
															assign node1246 = (inp[15]) ? node1248 : 4'b0101;
																assign node1248 = (inp[0]) ? 4'b0111 : 4'b0110;
														assign node1251 = (inp[4]) ? node1257 : node1252;
															assign node1252 = (inp[15]) ? node1254 : 4'b0111;
																assign node1254 = (inp[0]) ? 4'b0011 : 4'b0010;
															assign node1257 = (inp[15]) ? 4'b0100 : 4'b0110;
													assign node1260 = (inp[7]) ? node1272 : node1261;
														assign node1261 = (inp[15]) ? node1269 : node1262;
															assign node1262 = (inp[0]) ? node1266 : node1263;
																assign node1263 = (inp[4]) ? 4'b0010 : 4'b0110;
																assign node1266 = (inp[4]) ? 4'b0011 : 4'b0111;
															assign node1269 = (inp[4]) ? 4'b0100 : 4'b0110;
														assign node1272 = (inp[15]) ? node1276 : node1273;
															assign node1273 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node1276 = (inp[4]) ? 4'b0010 : 4'b0000;
							assign node1279 = (inp[10]) ? node1891 : node1280;
								assign node1280 = (inp[13]) ? node1588 : node1281;
									assign node1281 = (inp[2]) ? node1435 : node1282;
										assign node1282 = (inp[5]) ? node1352 : node1283;
											assign node1283 = (inp[15]) ? node1309 : node1284;
												assign node1284 = (inp[12]) ? node1288 : node1285;
													assign node1285 = (inp[7]) ? 4'b0011 : 4'b0001;
													assign node1288 = (inp[7]) ? node1296 : node1289;
														assign node1289 = (inp[1]) ? node1293 : node1290;
															assign node1290 = (inp[4]) ? 4'b0111 : 4'b0011;
															assign node1293 = (inp[4]) ? 4'b0110 : 4'b0010;
														assign node1296 = (inp[0]) ? node1302 : node1297;
															assign node1297 = (inp[1]) ? 4'b0001 : node1298;
																assign node1298 = (inp[4]) ? 4'b0101 : 4'b0001;
															assign node1302 = (inp[1]) ? node1306 : node1303;
																assign node1303 = (inp[4]) ? 4'b0100 : 4'b0000;
																assign node1306 = (inp[4]) ? 4'b0001 : 4'b0101;
												assign node1309 = (inp[7]) ? node1331 : node1310;
													assign node1310 = (inp[1]) ? node1320 : node1311;
														assign node1311 = (inp[0]) ? 4'b0011 : node1312;
															assign node1312 = (inp[4]) ? node1316 : node1313;
																assign node1313 = (inp[12]) ? 4'b0011 : 4'b0001;
																assign node1316 = (inp[12]) ? 4'b0001 : 4'b0011;
														assign node1320 = (inp[12]) ? node1326 : node1321;
															assign node1321 = (inp[4]) ? node1323 : 4'b0001;
																assign node1323 = (inp[0]) ? 4'b0110 : 4'b0111;
															assign node1326 = (inp[4]) ? 4'b0001 : node1327;
																assign node1327 = (inp[0]) ? 4'b0011 : 4'b0010;
													assign node1331 = (inp[12]) ? node1343 : node1332;
														assign node1332 = (inp[4]) ? node1338 : node1333;
															assign node1333 = (inp[1]) ? node1335 : 4'b0111;
																assign node1335 = (inp[0]) ? 4'b0110 : 4'b0111;
															assign node1338 = (inp[1]) ? 4'b0000 : node1339;
																assign node1339 = (inp[0]) ? 4'b0000 : 4'b0001;
														assign node1343 = (inp[4]) ? node1347 : node1344;
															assign node1344 = (inp[0]) ? 4'b0100 : 4'b0101;
															assign node1347 = (inp[0]) ? 4'b0110 : node1348;
																assign node1348 = (inp[1]) ? 4'b0111 : 4'b0110;
											assign node1352 = (inp[1]) ? node1392 : node1353;
												assign node1353 = (inp[7]) ? node1371 : node1354;
													assign node1354 = (inp[4]) ? node1358 : node1355;
														assign node1355 = (inp[12]) ? 4'b0011 : 4'b0001;
														assign node1358 = (inp[0]) ? node1366 : node1359;
															assign node1359 = (inp[12]) ? node1363 : node1360;
																assign node1360 = (inp[15]) ? 4'b0111 : 4'b0001;
																assign node1363 = (inp[15]) ? 4'b0000 : 4'b0111;
															assign node1366 = (inp[15]) ? node1368 : 4'b0000;
																assign node1368 = (inp[12]) ? 4'b0000 : 4'b0110;
													assign node1371 = (inp[12]) ? node1381 : node1372;
														assign node1372 = (inp[4]) ? node1376 : node1373;
															assign node1373 = (inp[15]) ? 4'b0110 : 4'b0010;
															assign node1376 = (inp[15]) ? 4'b0001 : node1377;
																assign node1377 = (inp[0]) ? 4'b0011 : 4'b0010;
														assign node1381 = (inp[4]) ? node1387 : node1382;
															assign node1382 = (inp[15]) ? 4'b0001 : node1383;
																assign node1383 = (inp[0]) ? 4'b0101 : 4'b0100;
															assign node1387 = (inp[15]) ? 4'b0110 : node1388;
																assign node1388 = (inp[0]) ? 4'b0000 : 4'b0001;
												assign node1392 = (inp[7]) ? node1412 : node1393;
													assign node1393 = (inp[15]) ? node1401 : node1394;
														assign node1394 = (inp[12]) ? 4'b0011 : node1395;
															assign node1395 = (inp[4]) ? node1397 : 4'b0101;
																assign node1397 = (inp[0]) ? 4'b0100 : 4'b0101;
														assign node1401 = (inp[4]) ? node1407 : node1402;
															assign node1402 = (inp[12]) ? node1404 : 4'b0101;
																assign node1404 = (inp[0]) ? 4'b0111 : 4'b0110;
															assign node1407 = (inp[12]) ? node1409 : 4'b0110;
																assign node1409 = (inp[0]) ? 4'b0100 : 4'b0101;
													assign node1412 = (inp[12]) ? node1424 : node1413;
														assign node1413 = (inp[15]) ? node1419 : node1414;
															assign node1414 = (inp[0]) ? node1416 : 4'b0110;
																assign node1416 = (inp[4]) ? 4'b0111 : 4'b0110;
															assign node1419 = (inp[4]) ? node1421 : 4'b0011;
																assign node1421 = (inp[0]) ? 4'b0100 : 4'b0101;
														assign node1424 = (inp[4]) ? node1428 : node1425;
															assign node1425 = (inp[0]) ? 4'b0001 : 4'b0101;
															assign node1428 = (inp[15]) ? node1432 : node1429;
																assign node1429 = (inp[0]) ? 4'b0001 : 4'b0000;
																assign node1432 = (inp[0]) ? 4'b0010 : 4'b0011;
										assign node1435 = (inp[1]) ? node1509 : node1436;
											assign node1436 = (inp[12]) ? node1472 : node1437;
												assign node1437 = (inp[7]) ? node1449 : node1438;
													assign node1438 = (inp[4]) ? node1440 : 4'b0101;
														assign node1440 = (inp[15]) ? node1446 : node1441;
															assign node1441 = (inp[5]) ? node1443 : 4'b0100;
																assign node1443 = (inp[0]) ? 4'b0101 : 4'b0100;
															assign node1446 = (inp[5]) ? 4'b0011 : 4'b0110;
													assign node1449 = (inp[15]) ? node1463 : node1450;
														assign node1450 = (inp[0]) ? node1458 : node1451;
															assign node1451 = (inp[4]) ? node1455 : node1452;
																assign node1452 = (inp[5]) ? 4'b0110 : 4'b0111;
																assign node1455 = (inp[5]) ? 4'b0111 : 4'b0110;
															assign node1458 = (inp[4]) ? 4'b0110 : node1459;
																assign node1459 = (inp[5]) ? 4'b0110 : 4'b0111;
														assign node1463 = (inp[4]) ? node1469 : node1464;
															assign node1464 = (inp[0]) ? node1466 : 4'b0011;
																assign node1466 = (inp[5]) ? 4'b0011 : 4'b0010;
															assign node1469 = (inp[0]) ? 4'b0101 : 4'b0100;
												assign node1472 = (inp[7]) ? node1488 : node1473;
													assign node1473 = (inp[15]) ? node1481 : node1474;
														assign node1474 = (inp[4]) ? node1476 : 4'b0111;
															assign node1476 = (inp[5]) ? 4'b0011 : node1477;
																assign node1477 = (inp[0]) ? 4'b0011 : 4'b0010;
														assign node1481 = (inp[4]) ? node1483 : 4'b0111;
															assign node1483 = (inp[0]) ? 4'b0101 : node1484;
																assign node1484 = (inp[5]) ? 4'b0101 : 4'b0100;
													assign node1488 = (inp[4]) ? node1498 : node1489;
														assign node1489 = (inp[5]) ? node1495 : node1490;
															assign node1490 = (inp[15]) ? 4'b0000 : node1491;
																assign node1491 = (inp[0]) ? 4'b0100 : 4'b0101;
															assign node1495 = (inp[15]) ? 4'b0101 : 4'b0001;
														assign node1498 = (inp[15]) ? node1504 : node1499;
															assign node1499 = (inp[0]) ? node1501 : 4'b0100;
																assign node1501 = (inp[5]) ? 4'b0101 : 4'b0001;
															assign node1504 = (inp[0]) ? node1506 : 4'b0011;
																assign node1506 = (inp[5]) ? 4'b0011 : 4'b0010;
											assign node1509 = (inp[5]) ? node1545 : node1510;
												assign node1510 = (inp[15]) ? node1528 : node1511;
													assign node1511 = (inp[4]) ? node1519 : node1512;
														assign node1512 = (inp[7]) ? node1516 : node1513;
															assign node1513 = (inp[12]) ? 4'b0110 : 4'b0101;
															assign node1516 = (inp[12]) ? 4'b0001 : 4'b0111;
														assign node1519 = (inp[12]) ? node1523 : node1520;
															assign node1520 = (inp[7]) ? 4'b0110 : 4'b0100;
															assign node1523 = (inp[7]) ? 4'b0100 : node1524;
																assign node1524 = (inp[0]) ? 4'b0010 : 4'b0011;
													assign node1528 = (inp[4]) ? node1538 : node1529;
														assign node1529 = (inp[7]) ? node1535 : node1530;
															assign node1530 = (inp[12]) ? 4'b0110 : node1531;
																assign node1531 = (inp[0]) ? 4'b0100 : 4'b0101;
															assign node1535 = (inp[12]) ? 4'b0101 : 4'b0010;
														assign node1538 = (inp[12]) ? node1542 : node1539;
															assign node1539 = (inp[7]) ? 4'b0101 : 4'b0011;
															assign node1542 = (inp[7]) ? 4'b0011 : 4'b0100;
												assign node1545 = (inp[7]) ? node1565 : node1546;
													assign node1546 = (inp[12]) ? node1556 : node1547;
														assign node1547 = (inp[4]) ? node1553 : node1548;
															assign node1548 = (inp[0]) ? 4'b0000 : node1549;
																assign node1549 = (inp[15]) ? 4'b0000 : 4'b0001;
															assign node1553 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node1556 = (inp[15]) ? node1562 : node1557;
															assign node1557 = (inp[4]) ? 4'b0110 : node1558;
																assign node1558 = (inp[0]) ? 4'b0011 : 4'b0010;
															assign node1562 = (inp[4]) ? 4'b0001 : 4'b0011;
													assign node1565 = (inp[12]) ? node1575 : node1566;
														assign node1566 = (inp[15]) ? node1572 : node1567;
															assign node1567 = (inp[0]) ? node1569 : 4'b0010;
																assign node1569 = (inp[4]) ? 4'b0010 : 4'b0011;
															assign node1572 = (inp[4]) ? 4'b0001 : 4'b0111;
														assign node1575 = (inp[4]) ? node1581 : node1576;
															assign node1576 = (inp[15]) ? node1578 : 4'b0000;
																assign node1578 = (inp[0]) ? 4'b0101 : 4'b0100;
															assign node1581 = (inp[15]) ? node1585 : node1582;
																assign node1582 = (inp[0]) ? 4'b0100 : 4'b0101;
																assign node1585 = (inp[0]) ? 4'b0111 : 4'b0110;
									assign node1588 = (inp[2]) ? node1724 : node1589;
										assign node1589 = (inp[15]) ? node1645 : node1590;
											assign node1590 = (inp[5]) ? node1610 : node1591;
												assign node1591 = (inp[12]) ? node1595 : node1592;
													assign node1592 = (inp[7]) ? 4'b0111 : 4'b0101;
													assign node1595 = (inp[7]) ? node1601 : node1596;
														assign node1596 = (inp[4]) ? 4'b0011 : node1597;
															assign node1597 = (inp[1]) ? 4'b0110 : 4'b0111;
														assign node1601 = (inp[1]) ? node1607 : node1602;
															assign node1602 = (inp[4]) ? 4'b0000 : node1603;
																assign node1603 = (inp[0]) ? 4'b0100 : 4'b0101;
															assign node1607 = (inp[4]) ? 4'b0101 : 4'b0001;
												assign node1610 = (inp[1]) ? node1626 : node1611;
													assign node1611 = (inp[12]) ? node1619 : node1612;
														assign node1612 = (inp[7]) ? 4'b0110 : node1613;
															assign node1613 = (inp[4]) ? node1615 : 4'b0101;
																assign node1615 = (inp[0]) ? 4'b0100 : 4'b0101;
														assign node1619 = (inp[7]) ? node1623 : node1620;
															assign node1620 = (inp[4]) ? 4'b0010 : 4'b0111;
															assign node1623 = (inp[4]) ? 4'b0101 : 4'b0001;
													assign node1626 = (inp[12]) ? node1634 : node1627;
														assign node1627 = (inp[7]) ? 4'b0011 : node1628;
															assign node1628 = (inp[0]) ? 4'b0000 : node1629;
																assign node1629 = (inp[4]) ? 4'b0000 : 4'b0001;
														assign node1634 = (inp[4]) ? node1640 : node1635;
															assign node1635 = (inp[0]) ? 4'b0011 : node1636;
																assign node1636 = (inp[7]) ? 4'b0000 : 4'b0010;
															assign node1640 = (inp[7]) ? node1642 : 4'b0111;
																assign node1642 = (inp[0]) ? 4'b0101 : 4'b0100;
											assign node1645 = (inp[4]) ? node1683 : node1646;
												assign node1646 = (inp[7]) ? node1660 : node1647;
													assign node1647 = (inp[12]) ? node1653 : node1648;
														assign node1648 = (inp[1]) ? node1650 : 4'b0100;
															assign node1650 = (inp[5]) ? 4'b0001 : 4'b0100;
														assign node1653 = (inp[1]) ? node1655 : 4'b0110;
															assign node1655 = (inp[5]) ? 4'b0010 : node1656;
																assign node1656 = (inp[0]) ? 4'b0110 : 4'b0111;
													assign node1660 = (inp[12]) ? node1672 : node1661;
														assign node1661 = (inp[5]) ? node1667 : node1662;
															assign node1662 = (inp[0]) ? 4'b0011 : node1663;
																assign node1663 = (inp[1]) ? 4'b0011 : 4'b0010;
															assign node1667 = (inp[1]) ? 4'b0110 : node1668;
																assign node1668 = (inp[0]) ? 4'b0010 : 4'b0011;
														assign node1672 = (inp[5]) ? node1678 : node1673;
															assign node1673 = (inp[1]) ? node1675 : 4'b0001;
																assign node1675 = (inp[0]) ? 4'b0101 : 4'b0100;
															assign node1678 = (inp[0]) ? 4'b0100 : node1679;
																assign node1679 = (inp[1]) ? 4'b0101 : 4'b0100;
												assign node1683 = (inp[1]) ? node1701 : node1684;
													assign node1684 = (inp[12]) ? node1690 : node1685;
														assign node1685 = (inp[7]) ? 4'b0100 : node1686;
															assign node1686 = (inp[5]) ? 4'b0011 : 4'b0110;
														assign node1690 = (inp[7]) ? node1696 : node1691;
															assign node1691 = (inp[5]) ? 4'b0101 : node1692;
																assign node1692 = (inp[0]) ? 4'b0101 : 4'b0100;
															assign node1696 = (inp[0]) ? node1698 : 4'b0011;
																assign node1698 = (inp[5]) ? 4'b0011 : 4'b0010;
													assign node1701 = (inp[0]) ? node1715 : node1702;
														assign node1702 = (inp[12]) ? node1708 : node1703;
															assign node1703 = (inp[7]) ? node1705 : 4'b0011;
																assign node1705 = (inp[5]) ? 4'b0001 : 4'b0101;
															assign node1708 = (inp[7]) ? node1712 : node1709;
																assign node1709 = (inp[5]) ? 4'b0001 : 4'b0100;
																assign node1712 = (inp[5]) ? 4'b0110 : 4'b0011;
														assign node1715 = (inp[5]) ? node1717 : 4'b0011;
															assign node1717 = (inp[12]) ? node1721 : node1718;
																assign node1718 = (inp[7]) ? 4'b0001 : 4'b0010;
																assign node1721 = (inp[7]) ? 4'b0111 : 4'b0001;
										assign node1724 = (inp[5]) ? node1806 : node1725;
											assign node1725 = (inp[7]) ? node1767 : node1726;
												assign node1726 = (inp[12]) ? node1746 : node1727;
													assign node1727 = (inp[4]) ? node1737 : node1728;
														assign node1728 = (inp[15]) ? node1732 : node1729;
															assign node1729 = (inp[0]) ? 4'b0000 : 4'b0001;
															assign node1732 = (inp[0]) ? 4'b0001 : node1733;
																assign node1733 = (inp[1]) ? 4'b0001 : 4'b0000;
														assign node1737 = (inp[15]) ? node1741 : node1738;
															assign node1738 = (inp[0]) ? 4'b0001 : 4'b0000;
															assign node1741 = (inp[1]) ? 4'b0110 : node1742;
																assign node1742 = (inp[0]) ? 4'b0010 : 4'b0011;
													assign node1746 = (inp[15]) ? node1760 : node1747;
														assign node1747 = (inp[4]) ? node1755 : node1748;
															assign node1748 = (inp[1]) ? node1752 : node1749;
																assign node1749 = (inp[0]) ? 4'b0010 : 4'b0011;
																assign node1752 = (inp[0]) ? 4'b0011 : 4'b0010;
															assign node1755 = (inp[1]) ? 4'b0111 : node1756;
																assign node1756 = (inp[0]) ? 4'b0111 : 4'b0110;
														assign node1760 = (inp[4]) ? node1762 : 4'b0010;
															assign node1762 = (inp[0]) ? 4'b0000 : node1763;
																assign node1763 = (inp[1]) ? 4'b0001 : 4'b0000;
												assign node1767 = (inp[12]) ? node1787 : node1768;
													assign node1768 = (inp[4]) ? node1778 : node1769;
														assign node1769 = (inp[15]) ? node1773 : node1770;
															assign node1770 = (inp[0]) ? 4'b0010 : 4'b0011;
															assign node1773 = (inp[0]) ? 4'b0111 : node1774;
																assign node1774 = (inp[1]) ? 4'b0111 : 4'b0110;
														assign node1778 = (inp[15]) ? node1782 : node1779;
															assign node1779 = (inp[0]) ? 4'b0011 : 4'b0010;
															assign node1782 = (inp[0]) ? node1784 : 4'b0000;
																assign node1784 = (inp[1]) ? 4'b0001 : 4'b0000;
													assign node1787 = (inp[4]) ? node1795 : node1788;
														assign node1788 = (inp[15]) ? node1792 : node1789;
															assign node1789 = (inp[1]) ? 4'b0101 : 4'b0000;
															assign node1792 = (inp[1]) ? 4'b0001 : 4'b0101;
														assign node1795 = (inp[15]) ? node1801 : node1796;
															assign node1796 = (inp[1]) ? node1798 : 4'b0101;
																assign node1798 = (inp[0]) ? 4'b0001 : 4'b0000;
															assign node1801 = (inp[1]) ? 4'b0110 : node1802;
																assign node1802 = (inp[0]) ? 4'b0111 : 4'b0110;
											assign node1806 = (inp[1]) ? node1852 : node1807;
												assign node1807 = (inp[12]) ? node1827 : node1808;
													assign node1808 = (inp[15]) ? node1814 : node1809;
														assign node1809 = (inp[7]) ? 4'b0010 : node1810;
															assign node1810 = (inp[4]) ? 4'b0001 : 4'b0000;
														assign node1814 = (inp[7]) ? node1820 : node1815;
															assign node1815 = (inp[4]) ? 4'b0110 : node1816;
																assign node1816 = (inp[0]) ? 4'b0001 : 4'b0000;
															assign node1820 = (inp[4]) ? node1824 : node1821;
																assign node1821 = (inp[0]) ? 4'b0110 : 4'b0111;
																assign node1824 = (inp[0]) ? 4'b0000 : 4'b0001;
													assign node1827 = (inp[15]) ? node1837 : node1828;
														assign node1828 = (inp[7]) ? node1834 : node1829;
															assign node1829 = (inp[4]) ? 4'b0111 : node1830;
																assign node1830 = (inp[0]) ? 4'b0010 : 4'b0011;
															assign node1834 = (inp[4]) ? 4'b0001 : 4'b0101;
														assign node1837 = (inp[0]) ? node1845 : node1838;
															assign node1838 = (inp[4]) ? node1842 : node1839;
																assign node1839 = (inp[7]) ? 4'b0000 : 4'b0010;
																assign node1842 = (inp[7]) ? 4'b0110 : 4'b0000;
															assign node1845 = (inp[4]) ? node1849 : node1846;
																assign node1846 = (inp[7]) ? 4'b0001 : 4'b0011;
																assign node1849 = (inp[7]) ? 4'b0110 : 4'b0001;
												assign node1852 = (inp[7]) ? node1872 : node1853;
													assign node1853 = (inp[12]) ? node1861 : node1854;
														assign node1854 = (inp[4]) ? node1856 : 4'b0101;
															assign node1856 = (inp[15]) ? node1858 : 4'b0101;
																assign node1858 = (inp[0]) ? 4'b0111 : 4'b0110;
														assign node1861 = (inp[15]) ? node1869 : node1862;
															assign node1862 = (inp[0]) ? node1866 : node1863;
																assign node1863 = (inp[4]) ? 4'b0010 : 4'b0110;
																assign node1866 = (inp[4]) ? 4'b0011 : 4'b0111;
															assign node1869 = (inp[4]) ? 4'b0100 : 4'b0110;
													assign node1872 = (inp[12]) ? node1884 : node1873;
														assign node1873 = (inp[4]) ? node1881 : node1874;
															assign node1874 = (inp[15]) ? node1878 : node1875;
																assign node1875 = (inp[0]) ? 4'b0111 : 4'b0110;
																assign node1878 = (inp[0]) ? 4'b0011 : 4'b0010;
															assign node1881 = (inp[15]) ? 4'b0100 : 4'b0110;
														assign node1884 = (inp[4]) ? node1888 : node1885;
															assign node1885 = (inp[15]) ? 4'b0000 : 4'b0100;
															assign node1888 = (inp[15]) ? 4'b0010 : 4'b0000;
								assign node1891 = (inp[4]) ? node2211 : node1892;
									assign node1892 = (inp[5]) ? node2032 : node1893;
										assign node1893 = (inp[12]) ? node1947 : node1894;
											assign node1894 = (inp[7]) ? node1914 : node1895;
												assign node1895 = (inp[13]) ? node1899 : node1896;
													assign node1896 = (inp[2]) ? 4'b0100 : 4'b0000;
													assign node1899 = (inp[2]) ? node1905 : node1900;
														assign node1900 = (inp[15]) ? node1902 : 4'b0100;
															assign node1902 = (inp[1]) ? 4'b0100 : 4'b0101;
														assign node1905 = (inp[15]) ? node1909 : node1906;
															assign node1906 = (inp[0]) ? 4'b0001 : 4'b0000;
															assign node1909 = (inp[0]) ? 4'b0000 : node1910;
																assign node1910 = (inp[1]) ? 4'b0000 : 4'b0001;
												assign node1914 = (inp[15]) ? node1924 : node1915;
													assign node1915 = (inp[13]) ? node1919 : node1916;
														assign node1916 = (inp[2]) ? 4'b0110 : 4'b0010;
														assign node1919 = (inp[2]) ? node1921 : 4'b0110;
															assign node1921 = (inp[0]) ? 4'b0011 : 4'b0010;
													assign node1924 = (inp[2]) ? node1936 : node1925;
														assign node1925 = (inp[13]) ? node1931 : node1926;
															assign node1926 = (inp[0]) ? node1928 : 4'b0110;
																assign node1928 = (inp[1]) ? 4'b0111 : 4'b0110;
															assign node1931 = (inp[0]) ? 4'b0010 : node1932;
																assign node1932 = (inp[1]) ? 4'b0010 : 4'b0011;
														assign node1936 = (inp[13]) ? node1942 : node1937;
															assign node1937 = (inp[1]) ? 4'b0011 : node1938;
																assign node1938 = (inp[0]) ? 4'b0011 : 4'b0010;
															assign node1942 = (inp[1]) ? 4'b0110 : node1943;
																assign node1943 = (inp[0]) ? 4'b0110 : 4'b0111;
											assign node1947 = (inp[7]) ? node1985 : node1948;
												assign node1948 = (inp[1]) ? node1964 : node1949;
													assign node1949 = (inp[13]) ? node1953 : node1950;
														assign node1950 = (inp[2]) ? 4'b0110 : 4'b0010;
														assign node1953 = (inp[2]) ? node1957 : node1954;
															assign node1954 = (inp[15]) ? 4'b0111 : 4'b0110;
															assign node1957 = (inp[15]) ? node1961 : node1958;
																assign node1958 = (inp[0]) ? 4'b0011 : 4'b0010;
																assign node1961 = (inp[0]) ? 4'b0010 : 4'b0011;
													assign node1964 = (inp[15]) ? node1972 : node1965;
														assign node1965 = (inp[2]) ? node1969 : node1966;
															assign node1966 = (inp[13]) ? 4'b0111 : 4'b0011;
															assign node1969 = (inp[13]) ? 4'b0011 : 4'b0111;
														assign node1972 = (inp[2]) ? node1980 : node1973;
															assign node1973 = (inp[13]) ? node1977 : node1974;
																assign node1974 = (inp[0]) ? 4'b0010 : 4'b0011;
																assign node1977 = (inp[0]) ? 4'b0111 : 4'b0110;
															assign node1980 = (inp[13]) ? 4'b0011 : node1981;
																assign node1981 = (inp[0]) ? 4'b0110 : 4'b0111;
												assign node1985 = (inp[13]) ? node2013 : node1986;
													assign node1986 = (inp[0]) ? node2002 : node1987;
														assign node1987 = (inp[1]) ? node1995 : node1988;
															assign node1988 = (inp[2]) ? node1992 : node1989;
																assign node1989 = (inp[15]) ? 4'b0100 : 4'b0000;
																assign node1992 = (inp[15]) ? 4'b0001 : 4'b0100;
															assign node1995 = (inp[2]) ? node1999 : node1996;
																assign node1996 = (inp[15]) ? 4'b0000 : 4'b0101;
																assign node1999 = (inp[15]) ? 4'b0100 : 4'b0000;
														assign node2002 = (inp[15]) ? node2008 : node2003;
															assign node2003 = (inp[1]) ? 4'b0100 : node2004;
																assign node2004 = (inp[2]) ? 4'b0101 : 4'b0001;
															assign node2008 = (inp[2]) ? 4'b0001 : node2009;
																assign node2009 = (inp[1]) ? 4'b0001 : 4'b0101;
													assign node2013 = (inp[15]) ? node2023 : node2014;
														assign node2014 = (inp[1]) ? node2020 : node2015;
															assign node2015 = (inp[2]) ? 4'b0001 : node2016;
																assign node2016 = (inp[0]) ? 4'b0101 : 4'b0100;
															assign node2020 = (inp[2]) ? 4'b0100 : 4'b0000;
														assign node2023 = (inp[2]) ? node2029 : node2024;
															assign node2024 = (inp[1]) ? node2026 : 4'b0000;
																assign node2026 = (inp[0]) ? 4'b0100 : 4'b0101;
															assign node2029 = (inp[1]) ? 4'b0000 : 4'b0100;
										assign node2032 = (inp[1]) ? node2110 : node2033;
											assign node2033 = (inp[7]) ? node2063 : node2034;
												assign node2034 = (inp[12]) ? node2048 : node2035;
													assign node2035 = (inp[13]) ? node2039 : node2036;
														assign node2036 = (inp[2]) ? 4'b0100 : 4'b0000;
														assign node2039 = (inp[2]) ? node2043 : node2040;
															assign node2040 = (inp[15]) ? 4'b0101 : 4'b0100;
															assign node2043 = (inp[15]) ? node2045 : 4'b0000;
																assign node2045 = (inp[0]) ? 4'b0000 : 4'b0001;
													assign node2048 = (inp[13]) ? node2052 : node2049;
														assign node2049 = (inp[2]) ? 4'b0110 : 4'b0010;
														assign node2052 = (inp[2]) ? node2056 : node2053;
															assign node2053 = (inp[15]) ? 4'b0111 : 4'b0110;
															assign node2056 = (inp[15]) ? node2060 : node2057;
																assign node2057 = (inp[0]) ? 4'b0011 : 4'b0010;
																assign node2060 = (inp[0]) ? 4'b0010 : 4'b0011;
												assign node2063 = (inp[12]) ? node2085 : node2064;
													assign node2064 = (inp[13]) ? node2074 : node2065;
														assign node2065 = (inp[15]) ? node2069 : node2066;
															assign node2066 = (inp[2]) ? 4'b0111 : 4'b0011;
															assign node2069 = (inp[2]) ? node2071 : 4'b0111;
																assign node2071 = (inp[0]) ? 4'b0010 : 4'b0011;
														assign node2074 = (inp[0]) ? node2078 : node2075;
															assign node2075 = (inp[15]) ? 4'b0010 : 4'b0011;
															assign node2078 = (inp[2]) ? node2082 : node2079;
																assign node2079 = (inp[15]) ? 4'b0011 : 4'b0111;
																assign node2082 = (inp[15]) ? 4'b0111 : 4'b0010;
													assign node2085 = (inp[13]) ? node2101 : node2086;
														assign node2086 = (inp[0]) ? node2094 : node2087;
															assign node2087 = (inp[2]) ? node2091 : node2088;
																assign node2088 = (inp[15]) ? 4'b0000 : 4'b0101;
																assign node2091 = (inp[15]) ? 4'b0100 : 4'b0000;
															assign node2094 = (inp[2]) ? node2098 : node2095;
																assign node2095 = (inp[15]) ? 4'b0000 : 4'b0100;
																assign node2098 = (inp[15]) ? 4'b0100 : 4'b0000;
														assign node2101 = (inp[15]) ? node2105 : node2102;
															assign node2102 = (inp[2]) ? 4'b0100 : 4'b0000;
															assign node2105 = (inp[2]) ? node2107 : 4'b0101;
																assign node2107 = (inp[0]) ? 4'b0000 : 4'b0001;
											assign node2110 = (inp[12]) ? node2168 : node2111;
												assign node2111 = (inp[7]) ? node2139 : node2112;
													assign node2112 = (inp[0]) ? node2128 : node2113;
														assign node2113 = (inp[15]) ? node2121 : node2114;
															assign node2114 = (inp[13]) ? node2118 : node2115;
																assign node2115 = (inp[2]) ? 4'b0000 : 4'b0100;
																assign node2118 = (inp[2]) ? 4'b0100 : 4'b0000;
															assign node2121 = (inp[13]) ? node2125 : node2122;
																assign node2122 = (inp[2]) ? 4'b0001 : 4'b0100;
																assign node2125 = (inp[2]) ? 4'b0100 : 4'b0000;
														assign node2128 = (inp[13]) ? node2132 : node2129;
															assign node2129 = (inp[2]) ? 4'b0001 : 4'b0101;
															assign node2132 = (inp[15]) ? node2136 : node2133;
																assign node2133 = (inp[2]) ? 4'b0101 : 4'b0001;
																assign node2136 = (inp[2]) ? 4'b0100 : 4'b0000;
													assign node2139 = (inp[0]) ? node2155 : node2140;
														assign node2140 = (inp[13]) ? node2148 : node2141;
															assign node2141 = (inp[15]) ? node2145 : node2142;
																assign node2142 = (inp[2]) ? 4'b0011 : 4'b0111;
																assign node2145 = (inp[2]) ? 4'b0110 : 4'b0010;
															assign node2148 = (inp[2]) ? node2152 : node2149;
																assign node2149 = (inp[15]) ? 4'b0111 : 4'b0011;
																assign node2152 = (inp[15]) ? 4'b0011 : 4'b0111;
														assign node2155 = (inp[2]) ? node2161 : node2156;
															assign node2156 = (inp[15]) ? node2158 : 4'b0010;
																assign node2158 = (inp[13]) ? 4'b0111 : 4'b0010;
															assign node2161 = (inp[15]) ? node2165 : node2162;
																assign node2162 = (inp[13]) ? 4'b0110 : 4'b0010;
																assign node2165 = (inp[13]) ? 4'b0010 : 4'b0110;
												assign node2168 = (inp[7]) ? node2192 : node2169;
													assign node2169 = (inp[0]) ? node2179 : node2170;
														assign node2170 = (inp[2]) ? node2174 : node2171;
															assign node2171 = (inp[13]) ? 4'b0011 : 4'b0111;
															assign node2174 = (inp[13]) ? 4'b0111 : node2175;
																assign node2175 = (inp[15]) ? 4'b0010 : 4'b0011;
														assign node2179 = (inp[13]) ? node2185 : node2180;
															assign node2180 = (inp[2]) ? 4'b0010 : node2181;
																assign node2181 = (inp[15]) ? 4'b0110 : 4'b0111;
															assign node2185 = (inp[15]) ? node2189 : node2186;
																assign node2186 = (inp[2]) ? 4'b0110 : 4'b0010;
																assign node2189 = (inp[2]) ? 4'b0111 : 4'b0011;
													assign node2192 = (inp[15]) ? node2202 : node2193;
														assign node2193 = (inp[13]) ? node2199 : node2194;
															assign node2194 = (inp[2]) ? 4'b0001 : node2195;
																assign node2195 = (inp[0]) ? 4'b0101 : 4'b0100;
															assign node2199 = (inp[2]) ? 4'b0101 : 4'b0001;
														assign node2202 = (inp[0]) ? node2206 : node2203;
															assign node2203 = (inp[13]) ? 4'b0100 : 4'b0001;
															assign node2206 = (inp[13]) ? 4'b0001 : node2207;
																assign node2207 = (inp[2]) ? 4'b0100 : 4'b0000;
									assign node2211 = (inp[2]) ? node2411 : node2212;
										assign node2212 = (inp[0]) ? node2308 : node2213;
											assign node2213 = (inp[13]) ? node2265 : node2214;
												assign node2214 = (inp[12]) ? node2238 : node2215;
													assign node2215 = (inp[5]) ? node2229 : node2216;
														assign node2216 = (inp[1]) ? node2224 : node2217;
															assign node2217 = (inp[15]) ? node2221 : node2218;
																assign node2218 = (inp[7]) ? 4'b0010 : 4'b0000;
																assign node2221 = (inp[7]) ? 4'b0000 : 4'b0010;
															assign node2224 = (inp[15]) ? 4'b0110 : node2225;
																assign node2225 = (inp[7]) ? 4'b0010 : 4'b0000;
														assign node2229 = (inp[1]) ? 4'b0111 : node2230;
															assign node2230 = (inp[7]) ? node2234 : node2231;
																assign node2231 = (inp[15]) ? 4'b0110 : 4'b0000;
																assign node2234 = (inp[15]) ? 4'b0000 : 4'b0011;
													assign node2238 = (inp[1]) ? node2250 : node2239;
														assign node2239 = (inp[15]) ? node2245 : node2240;
															assign node2240 = (inp[7]) ? node2242 : 4'b0110;
																assign node2242 = (inp[5]) ? 4'b0000 : 4'b0100;
															assign node2245 = (inp[7]) ? 4'b0110 : node2246;
																assign node2246 = (inp[5]) ? 4'b0001 : 4'b0000;
														assign node2250 = (inp[15]) ? node2258 : node2251;
															assign node2251 = (inp[7]) ? node2255 : node2252;
																assign node2252 = (inp[5]) ? 4'b0010 : 4'b0111;
																assign node2255 = (inp[5]) ? 4'b0001 : 4'b0000;
															assign node2258 = (inp[7]) ? node2262 : node2259;
																assign node2259 = (inp[5]) ? 4'b0100 : 4'b0000;
																assign node2262 = (inp[5]) ? 4'b0010 : 4'b0110;
												assign node2265 = (inp[15]) ? node2285 : node2266;
													assign node2266 = (inp[5]) ? node2274 : node2267;
														assign node2267 = (inp[12]) ? node2271 : node2268;
															assign node2268 = (inp[7]) ? 4'b0110 : 4'b0100;
															assign node2271 = (inp[1]) ? 4'b0100 : 4'b0001;
														assign node2274 = (inp[7]) ? node2280 : node2275;
															assign node2275 = (inp[12]) ? node2277 : 4'b0001;
																assign node2277 = (inp[1]) ? 4'b0110 : 4'b0011;
															assign node2280 = (inp[12]) ? node2282 : 4'b0111;
																assign node2282 = (inp[1]) ? 4'b0101 : 4'b0100;
													assign node2285 = (inp[1]) ? node2297 : node2286;
														assign node2286 = (inp[12]) ? node2292 : node2287;
															assign node2287 = (inp[7]) ? 4'b0101 : node2288;
																assign node2288 = (inp[5]) ? 4'b0010 : 4'b0111;
															assign node2292 = (inp[7]) ? 4'b0010 : node2293;
																assign node2293 = (inp[5]) ? 4'b0100 : 4'b0101;
														assign node2297 = (inp[12]) ? node2301 : node2298;
															assign node2298 = (inp[7]) ? 4'b0000 : 4'b0010;
															assign node2301 = (inp[7]) ? node2305 : node2302;
																assign node2302 = (inp[5]) ? 4'b0000 : 4'b0101;
																assign node2305 = (inp[5]) ? 4'b0111 : 4'b0010;
											assign node2308 = (inp[13]) ? node2360 : node2309;
												assign node2309 = (inp[15]) ? node2335 : node2310;
													assign node2310 = (inp[7]) ? node2324 : node2311;
														assign node2311 = (inp[12]) ? node2317 : node2312;
															assign node2312 = (inp[5]) ? node2314 : 4'b0000;
																assign node2314 = (inp[1]) ? 4'b0101 : 4'b0001;
															assign node2317 = (inp[1]) ? node2321 : node2318;
																assign node2318 = (inp[5]) ? 4'b0111 : 4'b0110;
																assign node2321 = (inp[5]) ? 4'b0010 : 4'b0111;
														assign node2324 = (inp[12]) ? node2330 : node2325;
															assign node2325 = (inp[1]) ? node2327 : 4'b0010;
																assign node2327 = (inp[5]) ? 4'b0110 : 4'b0010;
															assign node2330 = (inp[1]) ? 4'b0000 : node2331;
																assign node2331 = (inp[5]) ? 4'b0001 : 4'b0101;
													assign node2335 = (inp[5]) ? node2347 : node2336;
														assign node2336 = (inp[7]) ? node2344 : node2337;
															assign node2337 = (inp[12]) ? node2341 : node2338;
																assign node2338 = (inp[1]) ? 4'b0111 : 4'b0010;
																assign node2341 = (inp[1]) ? 4'b0000 : 4'b0001;
															assign node2344 = (inp[12]) ? 4'b0111 : 4'b0001;
														assign node2347 = (inp[7]) ? node2353 : node2348;
															assign node2348 = (inp[12]) ? node2350 : 4'b0111;
																assign node2350 = (inp[1]) ? 4'b0101 : 4'b0001;
															assign node2353 = (inp[12]) ? node2357 : node2354;
																assign node2354 = (inp[1]) ? 4'b0101 : 4'b0000;
																assign node2357 = (inp[1]) ? 4'b0011 : 4'b0111;
												assign node2360 = (inp[1]) ? node2386 : node2361;
													assign node2361 = (inp[12]) ? node2375 : node2362;
														assign node2362 = (inp[7]) ? node2370 : node2363;
															assign node2363 = (inp[15]) ? node2367 : node2364;
																assign node2364 = (inp[5]) ? 4'b0101 : 4'b0100;
																assign node2367 = (inp[5]) ? 4'b0010 : 4'b0111;
															assign node2370 = (inp[15]) ? node2372 : 4'b0110;
																assign node2372 = (inp[5]) ? 4'b0101 : 4'b0100;
														assign node2375 = (inp[15]) ? node2381 : node2376;
															assign node2376 = (inp[7]) ? node2378 : 4'b0011;
																assign node2378 = (inp[5]) ? 4'b0101 : 4'b0001;
															assign node2381 = (inp[7]) ? node2383 : 4'b0100;
																assign node2383 = (inp[5]) ? 4'b0010 : 4'b0011;
													assign node2386 = (inp[15]) ? node2396 : node2387;
														assign node2387 = (inp[5]) ? node2393 : node2388;
															assign node2388 = (inp[12]) ? 4'b0100 : node2389;
																assign node2389 = (inp[7]) ? 4'b0110 : 4'b0100;
															assign node2393 = (inp[12]) ? 4'b0110 : 4'b0010;
														assign node2396 = (inp[7]) ? node2404 : node2397;
															assign node2397 = (inp[12]) ? node2401 : node2398;
																assign node2398 = (inp[5]) ? 4'b0011 : 4'b0010;
																assign node2401 = (inp[5]) ? 4'b0000 : 4'b0101;
															assign node2404 = (inp[12]) ? node2408 : node2405;
																assign node2405 = (inp[5]) ? 4'b0000 : 4'b0100;
																assign node2408 = (inp[5]) ? 4'b0110 : 4'b0010;
										assign node2411 = (inp[13]) ? node2493 : node2412;
											assign node2412 = (inp[15]) ? node2452 : node2413;
												assign node2413 = (inp[7]) ? node2433 : node2414;
													assign node2414 = (inp[12]) ? node2422 : node2415;
														assign node2415 = (inp[5]) ? node2417 : 4'b0101;
															assign node2417 = (inp[1]) ? 4'b0000 : node2418;
																assign node2418 = (inp[0]) ? 4'b0100 : 4'b0101;
														assign node2422 = (inp[5]) ? node2430 : node2423;
															assign node2423 = (inp[0]) ? node2427 : node2424;
																assign node2424 = (inp[1]) ? 4'b0010 : 4'b0011;
																assign node2427 = (inp[1]) ? 4'b0011 : 4'b0010;
															assign node2430 = (inp[0]) ? 4'b0010 : 4'b0111;
													assign node2433 = (inp[12]) ? node2441 : node2434;
														assign node2434 = (inp[5]) ? node2436 : 4'b0111;
															assign node2436 = (inp[1]) ? 4'b0011 : node2437;
																assign node2437 = (inp[0]) ? 4'b0111 : 4'b0110;
														assign node2441 = (inp[1]) ? node2447 : node2442;
															assign node2442 = (inp[5]) ? node2444 : 4'b0000;
																assign node2444 = (inp[0]) ? 4'b0100 : 4'b0101;
															assign node2447 = (inp[0]) ? 4'b0101 : node2448;
																assign node2448 = (inp[5]) ? 4'b0100 : 4'b0101;
												assign node2452 = (inp[1]) ? node2474 : node2453;
													assign node2453 = (inp[12]) ? node2463 : node2454;
														assign node2454 = (inp[7]) ? node2458 : node2455;
															assign node2455 = (inp[5]) ? 4'b0010 : 4'b0111;
															assign node2458 = (inp[5]) ? 4'b0101 : node2459;
																assign node2459 = (inp[0]) ? 4'b0100 : 4'b0101;
														assign node2463 = (inp[7]) ? node2469 : node2464;
															assign node2464 = (inp[0]) ? 4'b0100 : node2465;
																assign node2465 = (inp[5]) ? 4'b0100 : 4'b0101;
															assign node2469 = (inp[5]) ? 4'b0010 : node2470;
																assign node2470 = (inp[0]) ? 4'b0011 : 4'b0010;
													assign node2474 = (inp[12]) ? node2484 : node2475;
														assign node2475 = (inp[7]) ? node2481 : node2476;
															assign node2476 = (inp[5]) ? node2478 : 4'b0010;
																assign node2478 = (inp[0]) ? 4'b0011 : 4'b0010;
															assign node2481 = (inp[5]) ? 4'b0000 : 4'b0100;
														assign node2484 = (inp[7]) ? node2488 : node2485;
															assign node2485 = (inp[5]) ? 4'b0000 : 4'b0101;
															assign node2488 = (inp[5]) ? node2490 : 4'b0010;
																assign node2490 = (inp[0]) ? 4'b0110 : 4'b0111;
											assign node2493 = (inp[15]) ? node2543 : node2494;
												assign node2494 = (inp[0]) ? node2518 : node2495;
													assign node2495 = (inp[7]) ? node2507 : node2496;
														assign node2496 = (inp[12]) ? node2502 : node2497;
															assign node2497 = (inp[5]) ? node2499 : 4'b0001;
																assign node2499 = (inp[1]) ? 4'b0100 : 4'b0000;
															assign node2502 = (inp[5]) ? 4'b0011 : node2503;
																assign node2503 = (inp[1]) ? 4'b0110 : 4'b0111;
														assign node2507 = (inp[12]) ? node2513 : node2508;
															assign node2508 = (inp[5]) ? node2510 : 4'b0011;
																assign node2510 = (inp[1]) ? 4'b0111 : 4'b0011;
															assign node2513 = (inp[1]) ? 4'b0001 : node2514;
																assign node2514 = (inp[5]) ? 4'b0000 : 4'b0100;
													assign node2518 = (inp[7]) ? node2530 : node2519;
														assign node2519 = (inp[12]) ? node2525 : node2520;
															assign node2520 = (inp[5]) ? node2522 : 4'b0000;
																assign node2522 = (inp[1]) ? 4'b0100 : 4'b0000;
															assign node2525 = (inp[1]) ? node2527 : 4'b0110;
																assign node2527 = (inp[5]) ? 4'b0010 : 4'b0111;
														assign node2530 = (inp[12]) ? node2536 : node2531;
															assign node2531 = (inp[5]) ? node2533 : 4'b0010;
																assign node2533 = (inp[1]) ? 4'b0111 : 4'b0011;
															assign node2536 = (inp[5]) ? node2540 : node2537;
																assign node2537 = (inp[1]) ? 4'b0000 : 4'b0100;
																assign node2540 = (inp[1]) ? 4'b0001 : 4'b0000;
												assign node2543 = (inp[1]) ? node2567 : node2544;
													assign node2544 = (inp[0]) ? node2556 : node2545;
														assign node2545 = (inp[12]) ? node2553 : node2546;
															assign node2546 = (inp[7]) ? node2550 : node2547;
																assign node2547 = (inp[5]) ? 4'b0111 : 4'b0010;
																assign node2550 = (inp[5]) ? 4'b0000 : 4'b0001;
															assign node2553 = (inp[7]) ? 4'b0111 : 4'b0001;
														assign node2556 = (inp[12]) ? node2562 : node2557;
															assign node2557 = (inp[7]) ? 4'b0001 : node2558;
																assign node2558 = (inp[5]) ? 4'b0111 : 4'b0011;
															assign node2562 = (inp[7]) ? node2564 : 4'b0000;
																assign node2564 = (inp[5]) ? 4'b0111 : 4'b0110;
													assign node2567 = (inp[5]) ? node2579 : node2568;
														assign node2568 = (inp[12]) ? node2574 : node2569;
															assign node2569 = (inp[7]) ? node2571 : 4'b0111;
																assign node2571 = (inp[0]) ? 4'b0000 : 4'b0001;
															assign node2574 = (inp[7]) ? 4'b0111 : node2575;
																assign node2575 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node2579 = (inp[12]) ? node2585 : node2580;
															assign node2580 = (inp[7]) ? 4'b0101 : node2581;
																assign node2581 = (inp[0]) ? 4'b0110 : 4'b0111;
															assign node2585 = (inp[7]) ? 4'b0011 : 4'b0101;
						assign node2588 = (inp[10]) ? node4138 : node2589;
							assign node2589 = (inp[4]) ? node3361 : node2590;
								assign node2590 = (inp[0]) ? node2946 : node2591;
									assign node2591 = (inp[9]) ? node2779 : node2592;
										assign node2592 = (inp[13]) ? node2680 : node2593;
											assign node2593 = (inp[2]) ? node2639 : node2594;
												assign node2594 = (inp[7]) ? node2612 : node2595;
													assign node2595 = (inp[12]) ? node2603 : node2596;
														assign node2596 = (inp[1]) ? node2598 : 4'b0000;
															assign node2598 = (inp[5]) ? 4'b0100 : node2599;
																assign node2599 = (inp[15]) ? 4'b0001 : 4'b0000;
														assign node2603 = (inp[1]) ? node2605 : 4'b0010;
															assign node2605 = (inp[15]) ? node2609 : node2606;
																assign node2606 = (inp[5]) ? 4'b0111 : 4'b0011;
																assign node2609 = (inp[5]) ? 4'b0110 : 4'b0010;
													assign node2612 = (inp[12]) ? node2626 : node2613;
														assign node2613 = (inp[15]) ? node2619 : node2614;
															assign node2614 = (inp[5]) ? node2616 : 4'b0010;
																assign node2616 = (inp[1]) ? 4'b0111 : 4'b0011;
															assign node2619 = (inp[1]) ? node2623 : node2620;
																assign node2620 = (inp[5]) ? 4'b0111 : 4'b0110;
																assign node2623 = (inp[5]) ? 4'b0010 : 4'b0111;
														assign node2626 = (inp[5]) ? node2634 : node2627;
															assign node2627 = (inp[1]) ? node2631 : node2628;
																assign node2628 = (inp[15]) ? 4'b0101 : 4'b0001;
																assign node2631 = (inp[15]) ? 4'b0001 : 4'b0100;
															assign node2634 = (inp[15]) ? 4'b0000 : node2635;
																assign node2635 = (inp[1]) ? 4'b0101 : 4'b0100;
												assign node2639 = (inp[5]) ? node2661 : node2640;
													assign node2640 = (inp[7]) ? node2650 : node2641;
														assign node2641 = (inp[12]) ? node2645 : node2642;
															assign node2642 = (inp[15]) ? 4'b0101 : 4'b0100;
															assign node2645 = (inp[1]) ? node2647 : 4'b0110;
																assign node2647 = (inp[15]) ? 4'b0110 : 4'b0111;
														assign node2650 = (inp[12]) ? node2654 : node2651;
															assign node2651 = (inp[15]) ? 4'b0011 : 4'b0110;
															assign node2654 = (inp[1]) ? node2658 : node2655;
																assign node2655 = (inp[15]) ? 4'b0001 : 4'b0101;
																assign node2658 = (inp[15]) ? 4'b0101 : 4'b0000;
													assign node2661 = (inp[1]) ? node2671 : node2662;
														assign node2662 = (inp[7]) ? node2666 : node2663;
															assign node2663 = (inp[12]) ? 4'b0110 : 4'b0100;
															assign node2666 = (inp[12]) ? 4'b0100 : node2667;
																assign node2667 = (inp[15]) ? 4'b0010 : 4'b0111;
														assign node2671 = (inp[7]) ? node2675 : node2672;
															assign node2672 = (inp[12]) ? 4'b0010 : 4'b0001;
															assign node2675 = (inp[15]) ? node2677 : 4'b0010;
																assign node2677 = (inp[12]) ? 4'b0100 : 4'b0110;
											assign node2680 = (inp[2]) ? node2726 : node2681;
												assign node2681 = (inp[5]) ? node2701 : node2682;
													assign node2682 = (inp[7]) ? node2694 : node2683;
														assign node2683 = (inp[12]) ? node2689 : node2684;
															assign node2684 = (inp[15]) ? node2686 : 4'b0100;
																assign node2686 = (inp[1]) ? 4'b0100 : 4'b0101;
															assign node2689 = (inp[1]) ? 4'b0111 : node2690;
																assign node2690 = (inp[15]) ? 4'b0111 : 4'b0110;
														assign node2694 = (inp[15]) ? node2698 : node2695;
															assign node2695 = (inp[12]) ? 4'b0101 : 4'b0110;
															assign node2698 = (inp[12]) ? 4'b0000 : 4'b0010;
													assign node2701 = (inp[1]) ? node2713 : node2702;
														assign node2702 = (inp[15]) ? node2708 : node2703;
															assign node2703 = (inp[7]) ? 4'b0111 : node2704;
																assign node2704 = (inp[12]) ? 4'b0110 : 4'b0100;
															assign node2708 = (inp[7]) ? 4'b0101 : node2709;
																assign node2709 = (inp[12]) ? 4'b0111 : 4'b0101;
														assign node2713 = (inp[7]) ? node2721 : node2714;
															assign node2714 = (inp[12]) ? node2718 : node2715;
																assign node2715 = (inp[15]) ? 4'b0000 : 4'b0001;
																assign node2718 = (inp[15]) ? 4'b0011 : 4'b0010;
															assign node2721 = (inp[12]) ? node2723 : 4'b0111;
																assign node2723 = (inp[15]) ? 4'b0101 : 4'b0001;
												assign node2726 = (inp[15]) ? node2754 : node2727;
													assign node2727 = (inp[1]) ? node2739 : node2728;
														assign node2728 = (inp[7]) ? node2732 : node2729;
															assign node2729 = (inp[12]) ? 4'b0011 : 4'b0001;
															assign node2732 = (inp[12]) ? node2736 : node2733;
																assign node2733 = (inp[5]) ? 4'b0010 : 4'b0011;
																assign node2736 = (inp[5]) ? 4'b0100 : 4'b0001;
														assign node2739 = (inp[5]) ? node2747 : node2740;
															assign node2740 = (inp[12]) ? node2744 : node2741;
																assign node2741 = (inp[7]) ? 4'b0011 : 4'b0001;
																assign node2744 = (inp[7]) ? 4'b0100 : 4'b0010;
															assign node2747 = (inp[12]) ? node2751 : node2748;
																assign node2748 = (inp[7]) ? 4'b0110 : 4'b0101;
																assign node2751 = (inp[7]) ? 4'b0101 : 4'b0110;
													assign node2754 = (inp[12]) ? node2766 : node2755;
														assign node2755 = (inp[7]) ? node2761 : node2756;
															assign node2756 = (inp[5]) ? node2758 : 4'b0000;
																assign node2758 = (inp[1]) ? 4'b0100 : 4'b0000;
															assign node2761 = (inp[5]) ? node2763 : 4'b0110;
																assign node2763 = (inp[1]) ? 4'b0010 : 4'b0111;
														assign node2766 = (inp[7]) ? node2772 : node2767;
															assign node2767 = (inp[1]) ? node2769 : 4'b0010;
																assign node2769 = (inp[5]) ? 4'b0111 : 4'b0011;
															assign node2772 = (inp[5]) ? node2776 : node2773;
																assign node2773 = (inp[1]) ? 4'b0000 : 4'b0100;
																assign node2776 = (inp[1]) ? 4'b0001 : 4'b0000;
										assign node2779 = (inp[13]) ? node2851 : node2780;
											assign node2780 = (inp[2]) ? node2814 : node2781;
												assign node2781 = (inp[7]) ? node2795 : node2782;
													assign node2782 = (inp[12]) ? node2790 : node2783;
														assign node2783 = (inp[1]) ? node2785 : 4'b0001;
															assign node2785 = (inp[5]) ? 4'b0100 : node2786;
																assign node2786 = (inp[15]) ? 4'b0000 : 4'b0001;
														assign node2790 = (inp[1]) ? node2792 : 4'b0011;
															assign node2792 = (inp[15]) ? 4'b0111 : 4'b0010;
													assign node2795 = (inp[12]) ? node2807 : node2796;
														assign node2796 = (inp[5]) ? node2800 : node2797;
															assign node2797 = (inp[15]) ? 4'b0111 : 4'b0011;
															assign node2800 = (inp[1]) ? node2804 : node2801;
																assign node2801 = (inp[15]) ? 4'b0110 : 4'b0010;
																assign node2804 = (inp[15]) ? 4'b0011 : 4'b0110;
														assign node2807 = (inp[15]) ? 4'b0001 : node2808;
															assign node2808 = (inp[5]) ? node2810 : 4'b0101;
																assign node2810 = (inp[1]) ? 4'b0100 : 4'b0101;
												assign node2814 = (inp[7]) ? node2828 : node2815;
													assign node2815 = (inp[12]) ? node2821 : node2816;
														assign node2816 = (inp[15]) ? node2818 : 4'b0101;
															assign node2818 = (inp[1]) ? 4'b0100 : 4'b0101;
														assign node2821 = (inp[1]) ? node2823 : 4'b0111;
															assign node2823 = (inp[5]) ? 4'b0011 : node2824;
																assign node2824 = (inp[15]) ? 4'b0111 : 4'b0110;
													assign node2828 = (inp[12]) ? node2842 : node2829;
														assign node2829 = (inp[15]) ? node2837 : node2830;
															assign node2830 = (inp[1]) ? node2834 : node2831;
																assign node2831 = (inp[5]) ? 4'b0110 : 4'b0111;
																assign node2834 = (inp[5]) ? 4'b0011 : 4'b0111;
															assign node2837 = (inp[5]) ? node2839 : 4'b0010;
																assign node2839 = (inp[1]) ? 4'b0111 : 4'b0011;
														assign node2842 = (inp[15]) ? node2848 : node2843;
															assign node2843 = (inp[1]) ? node2845 : 4'b0100;
																assign node2845 = (inp[5]) ? 4'b0000 : 4'b0001;
															assign node2848 = (inp[5]) ? 4'b0101 : 4'b0100;
											assign node2851 = (inp[2]) ? node2901 : node2852;
												assign node2852 = (inp[5]) ? node2876 : node2853;
													assign node2853 = (inp[7]) ? node2865 : node2854;
														assign node2854 = (inp[12]) ? node2860 : node2855;
															assign node2855 = (inp[15]) ? node2857 : 4'b0101;
																assign node2857 = (inp[1]) ? 4'b0101 : 4'b0100;
															assign node2860 = (inp[15]) ? 4'b0110 : node2861;
																assign node2861 = (inp[1]) ? 4'b0110 : 4'b0111;
														assign node2865 = (inp[12]) ? node2869 : node2866;
															assign node2866 = (inp[15]) ? 4'b0011 : 4'b0111;
															assign node2869 = (inp[15]) ? node2873 : node2870;
																assign node2870 = (inp[1]) ? 4'b0001 : 4'b0100;
																assign node2873 = (inp[1]) ? 4'b0101 : 4'b0001;
													assign node2876 = (inp[15]) ? node2892 : node2877;
														assign node2877 = (inp[1]) ? node2885 : node2878;
															assign node2878 = (inp[12]) ? node2882 : node2879;
																assign node2879 = (inp[7]) ? 4'b0110 : 4'b0101;
																assign node2882 = (inp[7]) ? 4'b0001 : 4'b0111;
															assign node2885 = (inp[7]) ? node2889 : node2886;
																assign node2886 = (inp[12]) ? 4'b0011 : 4'b0000;
																assign node2889 = (inp[12]) ? 4'b0000 : 4'b0011;
														assign node2892 = (inp[7]) ? node2896 : node2893;
															assign node2893 = (inp[12]) ? 4'b0010 : 4'b0001;
															assign node2896 = (inp[12]) ? 4'b0100 : node2897;
																assign node2897 = (inp[1]) ? 4'b0110 : 4'b0010;
												assign node2901 = (inp[1]) ? node2923 : node2902;
													assign node2902 = (inp[15]) ? node2914 : node2903;
														assign node2903 = (inp[7]) ? node2907 : node2904;
															assign node2904 = (inp[12]) ? 4'b0010 : 4'b0000;
															assign node2907 = (inp[5]) ? node2911 : node2908;
																assign node2908 = (inp[12]) ? 4'b0000 : 4'b0010;
																assign node2911 = (inp[12]) ? 4'b0101 : 4'b0011;
														assign node2914 = (inp[7]) ? node2918 : node2915;
															assign node2915 = (inp[12]) ? 4'b0011 : 4'b0001;
															assign node2918 = (inp[5]) ? 4'b0001 : node2919;
																assign node2919 = (inp[12]) ? 4'b0101 : 4'b0111;
													assign node2923 = (inp[5]) ? node2933 : node2924;
														assign node2924 = (inp[7]) ? node2930 : node2925;
															assign node2925 = (inp[12]) ? node2927 : 4'b0000;
																assign node2927 = (inp[15]) ? 4'b0010 : 4'b0011;
															assign node2930 = (inp[12]) ? 4'b0101 : 4'b0111;
														assign node2933 = (inp[12]) ? node2941 : node2934;
															assign node2934 = (inp[7]) ? node2938 : node2935;
																assign node2935 = (inp[15]) ? 4'b0101 : 4'b0100;
																assign node2938 = (inp[15]) ? 4'b0011 : 4'b0111;
															assign node2941 = (inp[7]) ? 4'b0100 : node2942;
																assign node2942 = (inp[15]) ? 4'b0110 : 4'b0111;
									assign node2946 = (inp[9]) ? node3152 : node2947;
										assign node2947 = (inp[5]) ? node3043 : node2948;
											assign node2948 = (inp[12]) ? node2986 : node2949;
												assign node2949 = (inp[7]) ? node2965 : node2950;
													assign node2950 = (inp[15]) ? node2958 : node2951;
														assign node2951 = (inp[2]) ? node2955 : node2952;
															assign node2952 = (inp[13]) ? 4'b0101 : 4'b0001;
															assign node2955 = (inp[13]) ? 4'b0001 : 4'b0101;
														assign node2958 = (inp[2]) ? node2962 : node2959;
															assign node2959 = (inp[13]) ? 4'b0100 : 4'b0001;
															assign node2962 = (inp[13]) ? 4'b0001 : 4'b0101;
													assign node2965 = (inp[15]) ? node2973 : node2966;
														assign node2966 = (inp[2]) ? node2970 : node2967;
															assign node2967 = (inp[13]) ? 4'b0111 : 4'b0011;
															assign node2970 = (inp[13]) ? 4'b0011 : 4'b0111;
														assign node2973 = (inp[2]) ? node2979 : node2974;
															assign node2974 = (inp[13]) ? node2976 : 4'b0111;
																assign node2976 = (inp[1]) ? 4'b0011 : 4'b0010;
															assign node2979 = (inp[13]) ? node2983 : node2980;
																assign node2980 = (inp[1]) ? 4'b0010 : 4'b0011;
																assign node2983 = (inp[1]) ? 4'b0111 : 4'b0110;
												assign node2986 = (inp[7]) ? node3018 : node2987;
													assign node2987 = (inp[1]) ? node3003 : node2988;
														assign node2988 = (inp[15]) ? node2996 : node2989;
															assign node2989 = (inp[13]) ? node2993 : node2990;
																assign node2990 = (inp[2]) ? 4'b0111 : 4'b0011;
																assign node2993 = (inp[2]) ? 4'b0011 : 4'b0111;
															assign node2996 = (inp[13]) ? node3000 : node2997;
																assign node2997 = (inp[2]) ? 4'b0111 : 4'b0011;
																assign node3000 = (inp[2]) ? 4'b0010 : 4'b0110;
														assign node3003 = (inp[15]) ? node3011 : node3004;
															assign node3004 = (inp[13]) ? node3008 : node3005;
																assign node3005 = (inp[2]) ? 4'b0110 : 4'b0010;
																assign node3008 = (inp[2]) ? 4'b0010 : 4'b0110;
															assign node3011 = (inp[2]) ? node3015 : node3012;
																assign node3012 = (inp[13]) ? 4'b0111 : 4'b0010;
																assign node3015 = (inp[13]) ? 4'b0010 : 4'b0110;
													assign node3018 = (inp[15]) ? node3030 : node3019;
														assign node3019 = (inp[13]) ? node3023 : node3020;
															assign node3020 = (inp[1]) ? 4'b0100 : 4'b0101;
															assign node3023 = (inp[1]) ? node3027 : node3024;
																assign node3024 = (inp[2]) ? 4'b0000 : 4'b0101;
																assign node3027 = (inp[2]) ? 4'b0101 : 4'b0001;
														assign node3030 = (inp[1]) ? node3036 : node3031;
															assign node3031 = (inp[2]) ? 4'b0000 : node3032;
																assign node3032 = (inp[13]) ? 4'b0001 : 4'b0101;
															assign node3036 = (inp[2]) ? node3040 : node3037;
																assign node3037 = (inp[13]) ? 4'b0100 : 4'b0001;
																assign node3040 = (inp[13]) ? 4'b0001 : 4'b0101;
											assign node3043 = (inp[7]) ? node3097 : node3044;
												assign node3044 = (inp[12]) ? node3072 : node3045;
													assign node3045 = (inp[15]) ? node3057 : node3046;
														assign node3046 = (inp[1]) ? node3052 : node3047;
															assign node3047 = (inp[2]) ? node3049 : 4'b0101;
																assign node3049 = (inp[13]) ? 4'b0001 : 4'b0101;
															assign node3052 = (inp[13]) ? node3054 : 4'b0001;
																assign node3054 = (inp[2]) ? 4'b0101 : 4'b0001;
														assign node3057 = (inp[13]) ? node3065 : node3058;
															assign node3058 = (inp[2]) ? node3062 : node3059;
																assign node3059 = (inp[1]) ? 4'b0101 : 4'b0001;
																assign node3062 = (inp[1]) ? 4'b0000 : 4'b0101;
															assign node3065 = (inp[1]) ? node3069 : node3066;
																assign node3066 = (inp[2]) ? 4'b0000 : 4'b0100;
																assign node3069 = (inp[2]) ? 4'b0101 : 4'b0001;
													assign node3072 = (inp[1]) ? node3088 : node3073;
														assign node3073 = (inp[15]) ? node3081 : node3074;
															assign node3074 = (inp[13]) ? node3078 : node3075;
																assign node3075 = (inp[2]) ? 4'b0111 : 4'b0011;
																assign node3078 = (inp[2]) ? 4'b0011 : 4'b0111;
															assign node3081 = (inp[13]) ? node3085 : node3082;
																assign node3082 = (inp[2]) ? 4'b0111 : 4'b0011;
																assign node3085 = (inp[2]) ? 4'b0010 : 4'b0110;
														assign node3088 = (inp[2]) ? node3092 : node3089;
															assign node3089 = (inp[13]) ? 4'b0010 : 4'b0110;
															assign node3092 = (inp[13]) ? 4'b0110 : node3093;
																assign node3093 = (inp[15]) ? 4'b0011 : 4'b0010;
												assign node3097 = (inp[12]) ? node3121 : node3098;
													assign node3098 = (inp[15]) ? node3110 : node3099;
														assign node3099 = (inp[13]) ? node3105 : node3100;
															assign node3100 = (inp[2]) ? 4'b0010 : node3101;
																assign node3101 = (inp[1]) ? 4'b0110 : 4'b0010;
															assign node3105 = (inp[2]) ? 4'b0110 : node3106;
																assign node3106 = (inp[1]) ? 4'b0010 : 4'b0110;
														assign node3110 = (inp[1]) ? node3114 : node3111;
															assign node3111 = (inp[2]) ? 4'b0010 : 4'b0110;
															assign node3114 = (inp[13]) ? node3118 : node3115;
																assign node3115 = (inp[2]) ? 4'b0111 : 4'b0011;
																assign node3118 = (inp[2]) ? 4'b0010 : 4'b0110;
													assign node3121 = (inp[1]) ? node3137 : node3122;
														assign node3122 = (inp[15]) ? node3130 : node3123;
															assign node3123 = (inp[2]) ? node3127 : node3124;
																assign node3124 = (inp[13]) ? 4'b0001 : 4'b0100;
																assign node3127 = (inp[13]) ? 4'b0101 : 4'b0001;
															assign node3130 = (inp[13]) ? node3134 : node3131;
																assign node3131 = (inp[2]) ? 4'b0101 : 4'b0001;
																assign node3134 = (inp[2]) ? 4'b0000 : 4'b0100;
														assign node3137 = (inp[2]) ? node3145 : node3138;
															assign node3138 = (inp[13]) ? node3142 : node3139;
																assign node3139 = (inp[15]) ? 4'b0000 : 4'b0101;
																assign node3142 = (inp[15]) ? 4'b0101 : 4'b0000;
															assign node3145 = (inp[15]) ? node3149 : node3146;
																assign node3146 = (inp[13]) ? 4'b0100 : 4'b0000;
																assign node3149 = (inp[13]) ? 4'b0000 : 4'b0100;
										assign node3152 = (inp[5]) ? node3256 : node3153;
											assign node3153 = (inp[15]) ? node3207 : node3154;
												assign node3154 = (inp[12]) ? node3176 : node3155;
													assign node3155 = (inp[7]) ? node3171 : node3156;
														assign node3156 = (inp[1]) ? node3164 : node3157;
															assign node3157 = (inp[13]) ? node3161 : node3158;
																assign node3158 = (inp[2]) ? 4'b0100 : 4'b0000;
																assign node3161 = (inp[2]) ? 4'b0000 : 4'b0100;
															assign node3164 = (inp[2]) ? node3168 : node3165;
																assign node3165 = (inp[13]) ? 4'b0100 : 4'b0000;
																assign node3168 = (inp[13]) ? 4'b0000 : 4'b0100;
														assign node3171 = (inp[2]) ? 4'b0010 : node3172;
															assign node3172 = (inp[13]) ? 4'b0110 : 4'b0010;
													assign node3176 = (inp[7]) ? node3192 : node3177;
														assign node3177 = (inp[1]) ? node3185 : node3178;
															assign node3178 = (inp[2]) ? node3182 : node3179;
																assign node3179 = (inp[13]) ? 4'b0110 : 4'b0010;
																assign node3182 = (inp[13]) ? 4'b0010 : 4'b0110;
															assign node3185 = (inp[13]) ? node3189 : node3186;
																assign node3186 = (inp[2]) ? 4'b0111 : 4'b0011;
																assign node3189 = (inp[2]) ? 4'b0011 : 4'b0111;
														assign node3192 = (inp[13]) ? node3200 : node3193;
															assign node3193 = (inp[2]) ? node3197 : node3194;
																assign node3194 = (inp[1]) ? 4'b0101 : 4'b0000;
																assign node3197 = (inp[1]) ? 4'b0000 : 4'b0100;
															assign node3200 = (inp[1]) ? node3204 : node3201;
																assign node3201 = (inp[2]) ? 4'b0001 : 4'b0100;
																assign node3204 = (inp[2]) ? 4'b0100 : 4'b0000;
												assign node3207 = (inp[13]) ? node3231 : node3208;
													assign node3208 = (inp[2]) ? node3220 : node3209;
														assign node3209 = (inp[7]) ? node3215 : node3210;
															assign node3210 = (inp[12]) ? node3212 : 4'b0000;
																assign node3212 = (inp[1]) ? 4'b0011 : 4'b0010;
															assign node3215 = (inp[1]) ? 4'b0000 : node3216;
																assign node3216 = (inp[12]) ? 4'b0100 : 4'b0110;
														assign node3220 = (inp[7]) ? node3226 : node3221;
															assign node3221 = (inp[12]) ? node3223 : 4'b0100;
																assign node3223 = (inp[1]) ? 4'b0111 : 4'b0110;
															assign node3226 = (inp[12]) ? node3228 : 4'b0011;
																assign node3228 = (inp[1]) ? 4'b0100 : 4'b0001;
													assign node3231 = (inp[1]) ? node3241 : node3232;
														assign node3232 = (inp[12]) ? node3238 : node3233;
															assign node3233 = (inp[7]) ? node3235 : 4'b0101;
																assign node3235 = (inp[2]) ? 4'b0111 : 4'b0011;
															assign node3238 = (inp[7]) ? 4'b0100 : 4'b0111;
														assign node3241 = (inp[2]) ? node3249 : node3242;
															assign node3242 = (inp[7]) ? node3246 : node3243;
																assign node3243 = (inp[12]) ? 4'b0110 : 4'b0101;
																assign node3246 = (inp[12]) ? 4'b0101 : 4'b0010;
															assign node3249 = (inp[12]) ? node3253 : node3250;
																assign node3250 = (inp[7]) ? 4'b0110 : 4'b0000;
																assign node3253 = (inp[7]) ? 4'b0000 : 4'b0011;
											assign node3256 = (inp[7]) ? node3304 : node3257;
												assign node3257 = (inp[12]) ? node3283 : node3258;
													assign node3258 = (inp[15]) ? node3272 : node3259;
														assign node3259 = (inp[1]) ? node3265 : node3260;
															assign node3260 = (inp[13]) ? node3262 : 4'b0100;
																assign node3262 = (inp[2]) ? 4'b0000 : 4'b0100;
															assign node3265 = (inp[13]) ? node3269 : node3266;
																assign node3266 = (inp[2]) ? 4'b0000 : 4'b0100;
																assign node3269 = (inp[2]) ? 4'b0100 : 4'b0000;
														assign node3272 = (inp[2]) ? node3276 : node3273;
															assign node3273 = (inp[13]) ? 4'b0000 : 4'b0100;
															assign node3276 = (inp[13]) ? node3280 : node3277;
																assign node3277 = (inp[1]) ? 4'b0001 : 4'b0100;
																assign node3280 = (inp[1]) ? 4'b0100 : 4'b0001;
													assign node3283 = (inp[1]) ? node3295 : node3284;
														assign node3284 = (inp[13]) ? node3288 : node3285;
															assign node3285 = (inp[2]) ? 4'b0110 : 4'b0010;
															assign node3288 = (inp[2]) ? node3292 : node3289;
																assign node3289 = (inp[15]) ? 4'b0111 : 4'b0110;
																assign node3292 = (inp[15]) ? 4'b0011 : 4'b0010;
														assign node3295 = (inp[2]) ? node3299 : node3296;
															assign node3296 = (inp[13]) ? 4'b0011 : 4'b0111;
															assign node3299 = (inp[13]) ? 4'b0111 : node3300;
																assign node3300 = (inp[15]) ? 4'b0010 : 4'b0011;
												assign node3304 = (inp[12]) ? node3334 : node3305;
													assign node3305 = (inp[15]) ? node3321 : node3306;
														assign node3306 = (inp[1]) ? node3314 : node3307;
															assign node3307 = (inp[2]) ? node3311 : node3308;
																assign node3308 = (inp[13]) ? 4'b0111 : 4'b0011;
																assign node3311 = (inp[13]) ? 4'b0011 : 4'b0111;
															assign node3314 = (inp[13]) ? node3318 : node3315;
																assign node3315 = (inp[2]) ? 4'b0011 : 4'b0111;
																assign node3318 = (inp[2]) ? 4'b0111 : 4'b0011;
														assign node3321 = (inp[1]) ? node3329 : node3322;
															assign node3322 = (inp[13]) ? node3326 : node3323;
																assign node3323 = (inp[2]) ? 4'b0011 : 4'b0111;
																assign node3326 = (inp[2]) ? 4'b0110 : 4'b0010;
															assign node3329 = (inp[13]) ? 4'b0011 : node3330;
																assign node3330 = (inp[2]) ? 4'b0110 : 4'b0010;
													assign node3334 = (inp[1]) ? node3348 : node3335;
														assign node3335 = (inp[15]) ? node3341 : node3336;
															assign node3336 = (inp[2]) ? node3338 : 4'b0000;
																assign node3338 = (inp[13]) ? 4'b0100 : 4'b0000;
															assign node3341 = (inp[13]) ? node3345 : node3342;
																assign node3342 = (inp[2]) ? 4'b0100 : 4'b0000;
																assign node3345 = (inp[2]) ? 4'b0001 : 4'b0101;
														assign node3348 = (inp[2]) ? node3354 : node3349;
															assign node3349 = (inp[13]) ? 4'b0001 : node3350;
																assign node3350 = (inp[15]) ? 4'b0001 : 4'b0100;
															assign node3354 = (inp[15]) ? node3358 : node3355;
																assign node3355 = (inp[13]) ? 4'b0101 : 4'b0001;
																assign node3358 = (inp[13]) ? 4'b0001 : 4'b0101;
								assign node3361 = (inp[9]) ? node3765 : node3362;
									assign node3362 = (inp[2]) ? node3568 : node3363;
										assign node3363 = (inp[0]) ? node3459 : node3364;
											assign node3364 = (inp[13]) ? node3416 : node3365;
												assign node3365 = (inp[15]) ? node3391 : node3366;
													assign node3366 = (inp[12]) ? node3378 : node3367;
														assign node3367 = (inp[7]) ? node3373 : node3368;
															assign node3368 = (inp[5]) ? node3370 : 4'b0000;
																assign node3370 = (inp[1]) ? 4'b0101 : 4'b0001;
															assign node3373 = (inp[1]) ? node3375 : 4'b0010;
																assign node3375 = (inp[5]) ? 4'b0110 : 4'b0010;
														assign node3378 = (inp[7]) ? node3386 : node3379;
															assign node3379 = (inp[5]) ? node3383 : node3380;
																assign node3380 = (inp[1]) ? 4'b0111 : 4'b0110;
																assign node3383 = (inp[1]) ? 4'b0010 : 4'b0111;
															assign node3386 = (inp[1]) ? 4'b0000 : node3387;
																assign node3387 = (inp[5]) ? 4'b0001 : 4'b0101;
													assign node3391 = (inp[5]) ? node3403 : node3392;
														assign node3392 = (inp[7]) ? node3400 : node3393;
															assign node3393 = (inp[12]) ? node3397 : node3394;
																assign node3394 = (inp[1]) ? 4'b0111 : 4'b0010;
																assign node3397 = (inp[1]) ? 4'b0000 : 4'b0001;
															assign node3400 = (inp[12]) ? 4'b0111 : 4'b0001;
														assign node3403 = (inp[7]) ? node3409 : node3404;
															assign node3404 = (inp[12]) ? node3406 : 4'b0111;
																assign node3406 = (inp[1]) ? 4'b0101 : 4'b0001;
															assign node3409 = (inp[12]) ? node3413 : node3410;
																assign node3410 = (inp[1]) ? 4'b0101 : 4'b0000;
																assign node3413 = (inp[1]) ? 4'b0011 : 4'b0111;
												assign node3416 = (inp[1]) ? node3442 : node3417;
													assign node3417 = (inp[15]) ? node3427 : node3418;
														assign node3418 = (inp[12]) ? node3422 : node3419;
															assign node3419 = (inp[5]) ? 4'b0101 : 4'b0110;
															assign node3422 = (inp[7]) ? node3424 : 4'b0011;
																assign node3424 = (inp[5]) ? 4'b0101 : 4'b0001;
														assign node3427 = (inp[5]) ? node3435 : node3428;
															assign node3428 = (inp[7]) ? node3432 : node3429;
																assign node3429 = (inp[12]) ? 4'b0100 : 4'b0111;
																assign node3432 = (inp[12]) ? 4'b0011 : 4'b0100;
															assign node3435 = (inp[12]) ? node3439 : node3436;
																assign node3436 = (inp[7]) ? 4'b0101 : 4'b0010;
																assign node3439 = (inp[7]) ? 4'b0010 : 4'b0100;
													assign node3442 = (inp[7]) ? node3450 : node3443;
														assign node3443 = (inp[12]) ? node3445 : 4'b0001;
															assign node3445 = (inp[15]) ? 4'b0000 : node3446;
																assign node3446 = (inp[5]) ? 4'b0110 : 4'b0010;
														assign node3450 = (inp[15]) ? node3454 : node3451;
															assign node3451 = (inp[12]) ? 4'b0100 : 4'b0110;
															assign node3454 = (inp[12]) ? 4'b0010 : node3455;
																assign node3455 = (inp[5]) ? 4'b0000 : 4'b0100;
											assign node3459 = (inp[13]) ? node3515 : node3460;
												assign node3460 = (inp[15]) ? node3488 : node3461;
													assign node3461 = (inp[7]) ? node3475 : node3462;
														assign node3462 = (inp[12]) ? node3468 : node3463;
															assign node3463 = (inp[5]) ? node3465 : 4'b0001;
																assign node3465 = (inp[1]) ? 4'b0101 : 4'b0001;
															assign node3468 = (inp[5]) ? node3472 : node3469;
																assign node3469 = (inp[1]) ? 4'b0110 : 4'b0111;
																assign node3472 = (inp[1]) ? 4'b0011 : 4'b0111;
														assign node3475 = (inp[12]) ? node3481 : node3476;
															assign node3476 = (inp[5]) ? node3478 : 4'b0011;
																assign node3478 = (inp[1]) ? 4'b0110 : 4'b0010;
															assign node3481 = (inp[1]) ? node3485 : node3482;
																assign node3482 = (inp[5]) ? 4'b0001 : 4'b0101;
																assign node3485 = (inp[5]) ? 4'b0000 : 4'b0001;
													assign node3488 = (inp[1]) ? node3502 : node3489;
														assign node3489 = (inp[12]) ? node3495 : node3490;
															assign node3490 = (inp[7]) ? 4'b0001 : node3491;
																assign node3491 = (inp[5]) ? 4'b0111 : 4'b0011;
															assign node3495 = (inp[7]) ? node3499 : node3496;
																assign node3496 = (inp[5]) ? 4'b0000 : 4'b0001;
																assign node3499 = (inp[5]) ? 4'b0111 : 4'b0110;
														assign node3502 = (inp[12]) ? node3508 : node3503;
															assign node3503 = (inp[7]) ? 4'b0101 : node3504;
																assign node3504 = (inp[5]) ? 4'b0110 : 4'b0111;
															assign node3508 = (inp[7]) ? node3512 : node3509;
																assign node3509 = (inp[5]) ? 4'b0101 : 4'b0001;
																assign node3512 = (inp[5]) ? 4'b0011 : 4'b0111;
												assign node3515 = (inp[1]) ? node3537 : node3516;
													assign node3516 = (inp[12]) ? node3528 : node3517;
														assign node3517 = (inp[7]) ? node3523 : node3518;
															assign node3518 = (inp[15]) ? node3520 : 4'b0101;
																assign node3520 = (inp[5]) ? 4'b0011 : 4'b0110;
															assign node3523 = (inp[15]) ? 4'b0100 : node3524;
																assign node3524 = (inp[5]) ? 4'b0110 : 4'b0111;
														assign node3528 = (inp[7]) ? node3532 : node3529;
															assign node3529 = (inp[5]) ? 4'b0101 : 4'b0100;
															assign node3532 = (inp[15]) ? 4'b0011 : node3533;
																assign node3533 = (inp[5]) ? 4'b0101 : 4'b0000;
													assign node3537 = (inp[12]) ? node3553 : node3538;
														assign node3538 = (inp[5]) ? node3546 : node3539;
															assign node3539 = (inp[7]) ? node3543 : node3540;
																assign node3540 = (inp[15]) ? 4'b0011 : 4'b0101;
																assign node3543 = (inp[15]) ? 4'b0101 : 4'b0111;
															assign node3546 = (inp[7]) ? node3550 : node3547;
																assign node3547 = (inp[15]) ? 4'b0011 : 4'b0000;
																assign node3550 = (inp[15]) ? 4'b0001 : 4'b0011;
														assign node3553 = (inp[15]) ? node3561 : node3554;
															assign node3554 = (inp[7]) ? node3558 : node3555;
																assign node3555 = (inp[5]) ? 4'b0111 : 4'b0010;
																assign node3558 = (inp[5]) ? 4'b0100 : 4'b0101;
															assign node3561 = (inp[7]) ? node3565 : node3562;
																assign node3562 = (inp[5]) ? 4'b0001 : 4'b0100;
																assign node3565 = (inp[5]) ? 4'b0110 : 4'b0011;
										assign node3568 = (inp[13]) ? node3662 : node3569;
											assign node3569 = (inp[1]) ? node3613 : node3570;
												assign node3570 = (inp[12]) ? node3592 : node3571;
													assign node3571 = (inp[7]) ? node3583 : node3572;
														assign node3572 = (inp[15]) ? node3578 : node3573;
															assign node3573 = (inp[5]) ? 4'b0100 : node3574;
																assign node3574 = (inp[0]) ? 4'b0100 : 4'b0101;
															assign node3578 = (inp[5]) ? node3580 : 4'b0111;
																assign node3580 = (inp[0]) ? 4'b0011 : 4'b0010;
														assign node3583 = (inp[15]) ? node3587 : node3584;
															assign node3584 = (inp[5]) ? 4'b0111 : 4'b0110;
															assign node3587 = (inp[5]) ? node3589 : 4'b0100;
																assign node3589 = (inp[0]) ? 4'b0100 : 4'b0101;
													assign node3592 = (inp[0]) ? node3602 : node3593;
														assign node3593 = (inp[7]) ? node3597 : node3594;
															assign node3594 = (inp[15]) ? 4'b0100 : 4'b0010;
															assign node3597 = (inp[15]) ? 4'b0011 : node3598;
																assign node3598 = (inp[5]) ? 4'b0100 : 4'b0000;
														assign node3602 = (inp[7]) ? node3608 : node3603;
															assign node3603 = (inp[15]) ? node3605 : 4'b0011;
																assign node3605 = (inp[5]) ? 4'b0101 : 4'b0100;
															assign node3608 = (inp[15]) ? 4'b0011 : node3609;
																assign node3609 = (inp[5]) ? 4'b0100 : 4'b0001;
												assign node3613 = (inp[5]) ? node3639 : node3614;
													assign node3614 = (inp[12]) ? node3628 : node3615;
														assign node3615 = (inp[7]) ? node3621 : node3616;
															assign node3616 = (inp[15]) ? 4'b0010 : node3617;
																assign node3617 = (inp[0]) ? 4'b0100 : 4'b0101;
															assign node3621 = (inp[15]) ? node3625 : node3622;
																assign node3622 = (inp[0]) ? 4'b0110 : 4'b0111;
																assign node3625 = (inp[0]) ? 4'b0101 : 4'b0100;
														assign node3628 = (inp[7]) ? node3634 : node3629;
															assign node3629 = (inp[15]) ? node3631 : 4'b0011;
																assign node3631 = (inp[0]) ? 4'b0100 : 4'b0101;
															assign node3634 = (inp[15]) ? node3636 : 4'b0100;
																assign node3636 = (inp[0]) ? 4'b0011 : 4'b0010;
													assign node3639 = (inp[12]) ? node3651 : node3640;
														assign node3640 = (inp[15]) ? node3646 : node3641;
															assign node3641 = (inp[7]) ? node3643 : 4'b0000;
																assign node3643 = (inp[0]) ? 4'b0010 : 4'b0011;
															assign node3646 = (inp[7]) ? node3648 : 4'b0011;
																assign node3648 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node3651 = (inp[15]) ? node3657 : node3652;
															assign node3652 = (inp[7]) ? 4'b0101 : node3653;
																assign node3653 = (inp[0]) ? 4'b0110 : 4'b0111;
															assign node3657 = (inp[7]) ? 4'b0110 : node3658;
																assign node3658 = (inp[0]) ? 4'b0001 : 4'b0000;
											assign node3662 = (inp[0]) ? node3710 : node3663;
												assign node3663 = (inp[15]) ? node3685 : node3664;
													assign node3664 = (inp[7]) ? node3674 : node3665;
														assign node3665 = (inp[12]) ? node3669 : node3666;
															assign node3666 = (inp[1]) ? 4'b0100 : 4'b0000;
															assign node3669 = (inp[1]) ? node3671 : 4'b0110;
																assign node3671 = (inp[5]) ? 4'b0010 : 4'b0111;
														assign node3674 = (inp[12]) ? node3680 : node3675;
															assign node3675 = (inp[5]) ? node3677 : 4'b0010;
																assign node3677 = (inp[1]) ? 4'b0111 : 4'b0011;
															assign node3680 = (inp[1]) ? 4'b0001 : node3681;
																assign node3681 = (inp[5]) ? 4'b0000 : 4'b0100;
													assign node3685 = (inp[1]) ? node3695 : node3686;
														assign node3686 = (inp[12]) ? node3688 : 4'b0001;
															assign node3688 = (inp[7]) ? node3692 : node3689;
																assign node3689 = (inp[5]) ? 4'b0000 : 4'b0001;
																assign node3692 = (inp[5]) ? 4'b0111 : 4'b0110;
														assign node3695 = (inp[12]) ? node3703 : node3696;
															assign node3696 = (inp[7]) ? node3700 : node3697;
																assign node3697 = (inp[5]) ? 4'b0110 : 4'b0111;
																assign node3700 = (inp[5]) ? 4'b0101 : 4'b0000;
															assign node3703 = (inp[7]) ? node3707 : node3704;
																assign node3704 = (inp[5]) ? 4'b0101 : 4'b0001;
																assign node3707 = (inp[5]) ? 4'b0011 : 4'b0111;
												assign node3710 = (inp[1]) ? node3738 : node3711;
													assign node3711 = (inp[12]) ? node3727 : node3712;
														assign node3712 = (inp[5]) ? node3720 : node3713;
															assign node3713 = (inp[15]) ? node3717 : node3714;
																assign node3714 = (inp[7]) ? 4'b0010 : 4'b0000;
																assign node3717 = (inp[7]) ? 4'b0000 : 4'b0011;
															assign node3720 = (inp[15]) ? node3724 : node3721;
																assign node3721 = (inp[7]) ? 4'b0010 : 4'b0001;
																assign node3724 = (inp[7]) ? 4'b0001 : 4'b0110;
														assign node3727 = (inp[15]) ? node3735 : node3728;
															assign node3728 = (inp[7]) ? node3732 : node3729;
																assign node3729 = (inp[5]) ? 4'b0111 : 4'b0110;
																assign node3732 = (inp[5]) ? 4'b0001 : 4'b0101;
															assign node3735 = (inp[7]) ? 4'b0110 : 4'b0000;
													assign node3738 = (inp[7]) ? node3752 : node3739;
														assign node3739 = (inp[5]) ? node3745 : node3740;
															assign node3740 = (inp[12]) ? 4'b0001 : node3741;
																assign node3741 = (inp[15]) ? 4'b0110 : 4'b0000;
															assign node3745 = (inp[12]) ? node3749 : node3746;
																assign node3746 = (inp[15]) ? 4'b0110 : 4'b0101;
																assign node3749 = (inp[15]) ? 4'b0100 : 4'b0010;
														assign node3752 = (inp[5]) ? node3758 : node3753;
															assign node3753 = (inp[12]) ? 4'b0110 : node3754;
																assign node3754 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node3758 = (inp[12]) ? node3762 : node3759;
																assign node3759 = (inp[15]) ? 4'b0100 : 4'b0110;
																assign node3762 = (inp[15]) ? 4'b0010 : 4'b0000;
									assign node3765 = (inp[13]) ? node3935 : node3766;
										assign node3766 = (inp[2]) ? node3846 : node3767;
											assign node3767 = (inp[7]) ? node3813 : node3768;
												assign node3768 = (inp[5]) ? node3792 : node3769;
													assign node3769 = (inp[0]) ? node3781 : node3770;
														assign node3770 = (inp[15]) ? node3776 : node3771;
															assign node3771 = (inp[12]) ? node3773 : 4'b0001;
																assign node3773 = (inp[1]) ? 4'b0110 : 4'b0111;
															assign node3776 = (inp[12]) ? node3778 : 4'b0011;
																assign node3778 = (inp[1]) ? 4'b0001 : 4'b0000;
														assign node3781 = (inp[12]) ? node3787 : node3782;
															assign node3782 = (inp[15]) ? node3784 : 4'b0000;
																assign node3784 = (inp[1]) ? 4'b0110 : 4'b0010;
															assign node3787 = (inp[15]) ? 4'b0000 : node3788;
																assign node3788 = (inp[1]) ? 4'b0111 : 4'b0110;
													assign node3792 = (inp[12]) ? node3802 : node3793;
														assign node3793 = (inp[15]) ? node3797 : node3794;
															assign node3794 = (inp[1]) ? 4'b0100 : 4'b0000;
															assign node3797 = (inp[1]) ? node3799 : 4'b0110;
																assign node3799 = (inp[0]) ? 4'b0111 : 4'b0110;
														assign node3802 = (inp[15]) ? node3808 : node3803;
															assign node3803 = (inp[1]) ? node3805 : 4'b0110;
																assign node3805 = (inp[0]) ? 4'b0010 : 4'b0011;
															assign node3808 = (inp[1]) ? 4'b0100 : node3809;
																assign node3809 = (inp[0]) ? 4'b0001 : 4'b0000;
												assign node3813 = (inp[15]) ? node3831 : node3814;
													assign node3814 = (inp[12]) ? node3822 : node3815;
														assign node3815 = (inp[5]) ? node3819 : node3816;
															assign node3816 = (inp[0]) ? 4'b0010 : 4'b0011;
															assign node3819 = (inp[1]) ? 4'b0111 : 4'b0011;
														assign node3822 = (inp[1]) ? node3826 : node3823;
															assign node3823 = (inp[5]) ? 4'b0000 : 4'b0100;
															assign node3826 = (inp[5]) ? 4'b0001 : node3827;
																assign node3827 = (inp[0]) ? 4'b0000 : 4'b0001;
													assign node3831 = (inp[12]) ? node3843 : node3832;
														assign node3832 = (inp[1]) ? node3838 : node3833;
															assign node3833 = (inp[0]) ? 4'b0000 : node3834;
																assign node3834 = (inp[5]) ? 4'b0001 : 4'b0000;
															assign node3838 = (inp[5]) ? 4'b0100 : node3839;
																assign node3839 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node3843 = (inp[5]) ? 4'b0010 : 4'b0110;
											assign node3846 = (inp[1]) ? node3894 : node3847;
												assign node3847 = (inp[12]) ? node3873 : node3848;
													assign node3848 = (inp[0]) ? node3858 : node3849;
														assign node3849 = (inp[15]) ? node3853 : node3850;
															assign node3850 = (inp[7]) ? 4'b0110 : 4'b0101;
															assign node3853 = (inp[7]) ? node3855 : 4'b0110;
																assign node3855 = (inp[5]) ? 4'b0100 : 4'b0101;
														assign node3858 = (inp[5]) ? node3866 : node3859;
															assign node3859 = (inp[15]) ? node3863 : node3860;
																assign node3860 = (inp[7]) ? 4'b0111 : 4'b0101;
																assign node3863 = (inp[7]) ? 4'b0101 : 4'b0111;
															assign node3866 = (inp[7]) ? node3870 : node3867;
																assign node3867 = (inp[15]) ? 4'b0010 : 4'b0101;
																assign node3870 = (inp[15]) ? 4'b0101 : 4'b0110;
													assign node3873 = (inp[7]) ? node3885 : node3874;
														assign node3874 = (inp[15]) ? node3880 : node3875;
															assign node3875 = (inp[0]) ? node3877 : 4'b0011;
																assign node3877 = (inp[5]) ? 4'b0010 : 4'b0011;
															assign node3880 = (inp[5]) ? node3882 : 4'b0101;
																assign node3882 = (inp[0]) ? 4'b0100 : 4'b0101;
														assign node3885 = (inp[15]) ? node3889 : node3886;
															assign node3886 = (inp[0]) ? 4'b0000 : 4'b0001;
															assign node3889 = (inp[0]) ? 4'b0010 : node3890;
																assign node3890 = (inp[5]) ? 4'b0011 : 4'b0010;
												assign node3894 = (inp[7]) ? node3912 : node3895;
													assign node3895 = (inp[15]) ? node3907 : node3896;
														assign node3896 = (inp[12]) ? node3904 : node3897;
															assign node3897 = (inp[5]) ? node3901 : node3898;
																assign node3898 = (inp[0]) ? 4'b0101 : 4'b0100;
																assign node3901 = (inp[0]) ? 4'b0000 : 4'b0001;
															assign node3904 = (inp[5]) ? 4'b0110 : 4'b0010;
														assign node3907 = (inp[12]) ? node3909 : 4'b0010;
															assign node3909 = (inp[5]) ? 4'b0000 : 4'b0100;
													assign node3912 = (inp[12]) ? node3926 : node3913;
														assign node3913 = (inp[15]) ? node3919 : node3914;
															assign node3914 = (inp[0]) ? node3916 : 4'b0010;
																assign node3916 = (inp[5]) ? 4'b0011 : 4'b0111;
															assign node3919 = (inp[5]) ? node3923 : node3920;
																assign node3920 = (inp[0]) ? 4'b0100 : 4'b0101;
																assign node3923 = (inp[0]) ? 4'b0000 : 4'b0001;
														assign node3926 = (inp[15]) ? node3932 : node3927;
															assign node3927 = (inp[5]) ? 4'b0100 : node3928;
																assign node3928 = (inp[0]) ? 4'b0101 : 4'b0100;
															assign node3932 = (inp[5]) ? 4'b0111 : 4'b0010;
										assign node3935 = (inp[2]) ? node4041 : node3936;
											assign node3936 = (inp[0]) ? node3990 : node3937;
												assign node3937 = (inp[1]) ? node3963 : node3938;
													assign node3938 = (inp[12]) ? node3952 : node3939;
														assign node3939 = (inp[5]) ? node3945 : node3940;
															assign node3940 = (inp[15]) ? 4'b0101 : node3941;
																assign node3941 = (inp[7]) ? 4'b0111 : 4'b0101;
															assign node3945 = (inp[7]) ? node3949 : node3946;
																assign node3946 = (inp[15]) ? 4'b0011 : 4'b0100;
																assign node3949 = (inp[15]) ? 4'b0100 : 4'b0111;
														assign node3952 = (inp[15]) ? node3958 : node3953;
															assign node3953 = (inp[7]) ? node3955 : 4'b0010;
																assign node3955 = (inp[5]) ? 4'b0100 : 4'b0000;
															assign node3958 = (inp[7]) ? node3960 : 4'b0101;
																assign node3960 = (inp[5]) ? 4'b0011 : 4'b0010;
													assign node3963 = (inp[7]) ? node3979 : node3964;
														assign node3964 = (inp[5]) ? node3972 : node3965;
															assign node3965 = (inp[12]) ? node3969 : node3966;
																assign node3966 = (inp[15]) ? 4'b0011 : 4'b0101;
																assign node3969 = (inp[15]) ? 4'b0100 : 4'b0011;
															assign node3972 = (inp[12]) ? node3976 : node3973;
																assign node3973 = (inp[15]) ? 4'b0010 : 4'b0000;
																assign node3976 = (inp[15]) ? 4'b0001 : 4'b0111;
														assign node3979 = (inp[5]) ? node3983 : node3980;
															assign node3980 = (inp[15]) ? 4'b0101 : 4'b0111;
															assign node3983 = (inp[12]) ? node3987 : node3984;
																assign node3984 = (inp[15]) ? 4'b0001 : 4'b0011;
																assign node3987 = (inp[15]) ? 4'b0111 : 4'b0101;
												assign node3990 = (inp[12]) ? node4012 : node3991;
													assign node3991 = (inp[1]) ? node4001 : node3992;
														assign node3992 = (inp[7]) ? node3998 : node3993;
															assign node3993 = (inp[5]) ? node3995 : 4'b0111;
																assign node3995 = (inp[15]) ? 4'b0010 : 4'b0100;
															assign node3998 = (inp[15]) ? 4'b0101 : 4'b0111;
														assign node4001 = (inp[5]) ? node4009 : node4002;
															assign node4002 = (inp[15]) ? node4006 : node4003;
																assign node4003 = (inp[7]) ? 4'b0110 : 4'b0100;
																assign node4006 = (inp[7]) ? 4'b0100 : 4'b0010;
															assign node4009 = (inp[15]) ? 4'b0000 : 4'b0010;
													assign node4012 = (inp[1]) ? node4026 : node4013;
														assign node4013 = (inp[5]) ? node4019 : node4014;
															assign node4014 = (inp[15]) ? 4'b0010 : node4015;
																assign node4015 = (inp[7]) ? 4'b0001 : 4'b0010;
															assign node4019 = (inp[7]) ? node4023 : node4020;
																assign node4020 = (inp[15]) ? 4'b0100 : 4'b0011;
																assign node4023 = (inp[15]) ? 4'b0010 : 4'b0100;
														assign node4026 = (inp[15]) ? node4034 : node4027;
															assign node4027 = (inp[7]) ? node4031 : node4028;
																assign node4028 = (inp[5]) ? 4'b0110 : 4'b0011;
																assign node4031 = (inp[5]) ? 4'b0101 : 4'b0100;
															assign node4034 = (inp[7]) ? node4038 : node4035;
																assign node4035 = (inp[5]) ? 4'b0000 : 4'b0101;
																assign node4038 = (inp[5]) ? 4'b0111 : 4'b0010;
											assign node4041 = (inp[0]) ? node4095 : node4042;
												assign node4042 = (inp[15]) ? node4068 : node4043;
													assign node4043 = (inp[7]) ? node4055 : node4044;
														assign node4044 = (inp[12]) ? node4050 : node4045;
															assign node4045 = (inp[5]) ? node4047 : 4'b0001;
																assign node4047 = (inp[1]) ? 4'b0101 : 4'b0001;
															assign node4050 = (inp[5]) ? node4052 : 4'b0110;
																assign node4052 = (inp[1]) ? 4'b0011 : 4'b0111;
														assign node4055 = (inp[12]) ? node4061 : node4056;
															assign node4056 = (inp[1]) ? 4'b0110 : node4057;
																assign node4057 = (inp[5]) ? 4'b0010 : 4'b0011;
															assign node4061 = (inp[1]) ? node4065 : node4062;
																assign node4062 = (inp[5]) ? 4'b0001 : 4'b0101;
																assign node4065 = (inp[5]) ? 4'b0000 : 4'b0001;
													assign node4068 = (inp[5]) ? node4080 : node4069;
														assign node4069 = (inp[7]) ? node4075 : node4070;
															assign node4070 = (inp[12]) ? 4'b0000 : node4071;
																assign node4071 = (inp[1]) ? 4'b0110 : 4'b0010;
															assign node4075 = (inp[12]) ? node4077 : 4'b0001;
																assign node4077 = (inp[1]) ? 4'b0110 : 4'b0111;
														assign node4080 = (inp[7]) ? node4088 : node4081;
															assign node4081 = (inp[12]) ? node4085 : node4082;
																assign node4082 = (inp[1]) ? 4'b0111 : 4'b0110;
																assign node4085 = (inp[1]) ? 4'b0100 : 4'b0001;
															assign node4088 = (inp[12]) ? node4092 : node4089;
																assign node4089 = (inp[1]) ? 4'b0100 : 4'b0000;
																assign node4092 = (inp[1]) ? 4'b0010 : 4'b0110;
												assign node4095 = (inp[1]) ? node4119 : node4096;
													assign node4096 = (inp[12]) ? node4108 : node4097;
														assign node4097 = (inp[7]) ? node4103 : node4098;
															assign node4098 = (inp[15]) ? node4100 : 4'b0000;
																assign node4100 = (inp[5]) ? 4'b0111 : 4'b0010;
															assign node4103 = (inp[15]) ? node4105 : 4'b0011;
																assign node4105 = (inp[5]) ? 4'b0000 : 4'b0001;
														assign node4108 = (inp[15]) ? node4116 : node4109;
															assign node4109 = (inp[7]) ? node4113 : node4110;
																assign node4110 = (inp[5]) ? 4'b0110 : 4'b0111;
																assign node4113 = (inp[5]) ? 4'b0000 : 4'b0100;
															assign node4116 = (inp[7]) ? 4'b0111 : 4'b0001;
													assign node4119 = (inp[15]) ? node4131 : node4120;
														assign node4120 = (inp[7]) ? node4126 : node4121;
															assign node4121 = (inp[12]) ? node4123 : 4'b0001;
																assign node4123 = (inp[5]) ? 4'b0011 : 4'b0110;
															assign node4126 = (inp[12]) ? 4'b0001 : node4127;
																assign node4127 = (inp[5]) ? 4'b0111 : 4'b0011;
														assign node4131 = (inp[5]) ? 4'b0101 : node4132;
															assign node4132 = (inp[7]) ? node4134 : 4'b0111;
																assign node4134 = (inp[12]) ? 4'b0111 : 4'b0001;
							assign node4138 = (inp[5]) ? node4910 : node4139;
								assign node4139 = (inp[15]) ? node4553 : node4140;
									assign node4140 = (inp[1]) ? node4354 : node4141;
										assign node4141 = (inp[9]) ? node4245 : node4142;
											assign node4142 = (inp[0]) ? node4196 : node4143;
												assign node4143 = (inp[7]) ? node4171 : node4144;
													assign node4144 = (inp[12]) ? node4156 : node4145;
														assign node4145 = (inp[2]) ? node4149 : node4146;
															assign node4146 = (inp[13]) ? 4'b0101 : 4'b0001;
															assign node4149 = (inp[13]) ? node4153 : node4150;
																assign node4150 = (inp[4]) ? 4'b0100 : 4'b0101;
																assign node4153 = (inp[4]) ? 4'b0001 : 4'b0000;
														assign node4156 = (inp[13]) ? node4164 : node4157;
															assign node4157 = (inp[4]) ? node4161 : node4158;
																assign node4158 = (inp[2]) ? 4'b0111 : 4'b0011;
																assign node4161 = (inp[2]) ? 4'b0011 : 4'b0111;
															assign node4164 = (inp[4]) ? node4168 : node4165;
																assign node4165 = (inp[2]) ? 4'b0010 : 4'b0111;
																assign node4168 = (inp[2]) ? 4'b0111 : 4'b0010;
													assign node4171 = (inp[12]) ? node4181 : node4172;
														assign node4172 = (inp[2]) ? node4176 : node4173;
															assign node4173 = (inp[13]) ? 4'b0111 : 4'b0011;
															assign node4176 = (inp[13]) ? 4'b0010 : node4177;
																assign node4177 = (inp[4]) ? 4'b0110 : 4'b0111;
														assign node4181 = (inp[4]) ? node4189 : node4182;
															assign node4182 = (inp[13]) ? node4186 : node4183;
																assign node4183 = (inp[2]) ? 4'b0100 : 4'b0000;
																assign node4186 = (inp[2]) ? 4'b0000 : 4'b0100;
															assign node4189 = (inp[2]) ? node4193 : node4190;
																assign node4190 = (inp[13]) ? 4'b0000 : 4'b0100;
																assign node4193 = (inp[13]) ? 4'b0101 : 4'b0001;
												assign node4196 = (inp[2]) ? node4218 : node4197;
													assign node4197 = (inp[13]) ? node4209 : node4198;
														assign node4198 = (inp[12]) ? node4202 : node4199;
															assign node4199 = (inp[7]) ? 4'b0010 : 4'b0000;
															assign node4202 = (inp[4]) ? node4206 : node4203;
																assign node4203 = (inp[7]) ? 4'b0000 : 4'b0010;
																assign node4206 = (inp[7]) ? 4'b0100 : 4'b0110;
														assign node4209 = (inp[12]) ? node4213 : node4210;
															assign node4210 = (inp[7]) ? 4'b0110 : 4'b0100;
															assign node4213 = (inp[7]) ? 4'b0001 : node4214;
																assign node4214 = (inp[4]) ? 4'b0010 : 4'b0110;
													assign node4218 = (inp[4]) ? node4232 : node4219;
														assign node4219 = (inp[13]) ? node4225 : node4220;
															assign node4220 = (inp[7]) ? 4'b0110 : node4221;
																assign node4221 = (inp[12]) ? 4'b0110 : 4'b0100;
															assign node4225 = (inp[7]) ? node4229 : node4226;
																assign node4226 = (inp[12]) ? 4'b0010 : 4'b0000;
																assign node4229 = (inp[12]) ? 4'b0001 : 4'b0010;
														assign node4232 = (inp[12]) ? node4238 : node4233;
															assign node4233 = (inp[13]) ? node4235 : 4'b0111;
																assign node4235 = (inp[7]) ? 4'b0011 : 4'b0001;
															assign node4238 = (inp[7]) ? node4242 : node4239;
																assign node4239 = (inp[13]) ? 4'b0111 : 4'b0011;
																assign node4242 = (inp[13]) ? 4'b0100 : 4'b0000;
											assign node4245 = (inp[0]) ? node4299 : node4246;
												assign node4246 = (inp[7]) ? node4274 : node4247;
													assign node4247 = (inp[12]) ? node4259 : node4248;
														assign node4248 = (inp[2]) ? node4252 : node4249;
															assign node4249 = (inp[13]) ? 4'b0100 : 4'b0000;
															assign node4252 = (inp[13]) ? node4256 : node4253;
																assign node4253 = (inp[4]) ? 4'b0101 : 4'b0100;
																assign node4256 = (inp[4]) ? 4'b0000 : 4'b0001;
														assign node4259 = (inp[13]) ? node4267 : node4260;
															assign node4260 = (inp[4]) ? node4264 : node4261;
																assign node4261 = (inp[2]) ? 4'b0110 : 4'b0010;
																assign node4264 = (inp[2]) ? 4'b0010 : 4'b0110;
															assign node4267 = (inp[2]) ? node4271 : node4268;
																assign node4268 = (inp[4]) ? 4'b0011 : 4'b0110;
																assign node4271 = (inp[4]) ? 4'b0110 : 4'b0011;
													assign node4274 = (inp[12]) ? node4286 : node4275;
														assign node4275 = (inp[2]) ? node4279 : node4276;
															assign node4276 = (inp[13]) ? 4'b0110 : 4'b0010;
															assign node4279 = (inp[13]) ? node4283 : node4280;
																assign node4280 = (inp[4]) ? 4'b0111 : 4'b0110;
																assign node4283 = (inp[4]) ? 4'b0010 : 4'b0011;
														assign node4286 = (inp[4]) ? node4294 : node4287;
															assign node4287 = (inp[13]) ? node4291 : node4288;
																assign node4288 = (inp[2]) ? 4'b0101 : 4'b0001;
																assign node4291 = (inp[2]) ? 4'b0001 : 4'b0101;
															assign node4294 = (inp[2]) ? node4296 : 4'b0001;
																assign node4296 = (inp[13]) ? 4'b0100 : 4'b0000;
												assign node4299 = (inp[4]) ? node4331 : node4300;
													assign node4300 = (inp[12]) ? node4316 : node4301;
														assign node4301 = (inp[7]) ? node4309 : node4302;
															assign node4302 = (inp[13]) ? node4306 : node4303;
																assign node4303 = (inp[2]) ? 4'b0101 : 4'b0001;
																assign node4306 = (inp[2]) ? 4'b0001 : 4'b0101;
															assign node4309 = (inp[13]) ? node4313 : node4310;
																assign node4310 = (inp[2]) ? 4'b0111 : 4'b0011;
																assign node4313 = (inp[2]) ? 4'b0011 : 4'b0111;
														assign node4316 = (inp[7]) ? node4324 : node4317;
															assign node4317 = (inp[13]) ? node4321 : node4318;
																assign node4318 = (inp[2]) ? 4'b0111 : 4'b0011;
																assign node4321 = (inp[2]) ? 4'b0011 : 4'b0111;
															assign node4324 = (inp[13]) ? node4328 : node4325;
																assign node4325 = (inp[2]) ? 4'b0101 : 4'b0001;
																assign node4328 = (inp[2]) ? 4'b0000 : 4'b0101;
													assign node4331 = (inp[2]) ? node4343 : node4332;
														assign node4332 = (inp[7]) ? node4338 : node4333;
															assign node4333 = (inp[12]) ? node4335 : 4'b0001;
																assign node4335 = (inp[13]) ? 4'b0011 : 4'b0111;
															assign node4338 = (inp[12]) ? node4340 : 4'b0111;
																assign node4340 = (inp[13]) ? 4'b0000 : 4'b0101;
														assign node4343 = (inp[7]) ? node4347 : node4344;
															assign node4344 = (inp[13]) ? 4'b0110 : 4'b0010;
															assign node4347 = (inp[12]) ? node4351 : node4348;
																assign node4348 = (inp[13]) ? 4'b0010 : 4'b0110;
																assign node4351 = (inp[13]) ? 4'b0101 : 4'b0001;
										assign node4354 = (inp[9]) ? node4458 : node4355;
											assign node4355 = (inp[0]) ? node4405 : node4356;
												assign node4356 = (inp[7]) ? node4382 : node4357;
													assign node4357 = (inp[12]) ? node4369 : node4358;
														assign node4358 = (inp[2]) ? node4362 : node4359;
															assign node4359 = (inp[13]) ? 4'b0101 : 4'b0001;
															assign node4362 = (inp[13]) ? node4366 : node4363;
																assign node4363 = (inp[4]) ? 4'b0100 : 4'b0101;
																assign node4366 = (inp[4]) ? 4'b0001 : 4'b0000;
														assign node4369 = (inp[13]) ? node4377 : node4370;
															assign node4370 = (inp[4]) ? node4374 : node4371;
																assign node4371 = (inp[2]) ? 4'b0110 : 4'b0010;
																assign node4374 = (inp[2]) ? 4'b0010 : 4'b0110;
															assign node4377 = (inp[2]) ? node4379 : 4'b0110;
																assign node4379 = (inp[4]) ? 4'b0110 : 4'b0011;
													assign node4382 = (inp[12]) ? node4392 : node4383;
														assign node4383 = (inp[2]) ? node4387 : node4384;
															assign node4384 = (inp[13]) ? 4'b0111 : 4'b0011;
															assign node4387 = (inp[13]) ? node4389 : 4'b0111;
																assign node4389 = (inp[4]) ? 4'b0011 : 4'b0010;
														assign node4392 = (inp[4]) ? node4400 : node4393;
															assign node4393 = (inp[2]) ? node4397 : node4394;
																assign node4394 = (inp[13]) ? 4'b0001 : 4'b0101;
																assign node4397 = (inp[13]) ? 4'b0101 : 4'b0001;
															assign node4400 = (inp[2]) ? 4'b0100 : node4401;
																assign node4401 = (inp[13]) ? 4'b0101 : 4'b0001;
												assign node4405 = (inp[12]) ? node4431 : node4406;
													assign node4406 = (inp[7]) ? node4418 : node4407;
														assign node4407 = (inp[2]) ? node4411 : node4408;
															assign node4408 = (inp[13]) ? 4'b0100 : 4'b0000;
															assign node4411 = (inp[4]) ? node4415 : node4412;
																assign node4412 = (inp[13]) ? 4'b0000 : 4'b0100;
																assign node4415 = (inp[13]) ? 4'b0001 : 4'b0101;
														assign node4418 = (inp[4]) ? node4424 : node4419;
															assign node4419 = (inp[13]) ? node4421 : 4'b0110;
																assign node4421 = (inp[2]) ? 4'b0010 : 4'b0110;
															assign node4424 = (inp[2]) ? node4428 : node4425;
																assign node4425 = (inp[13]) ? 4'b0110 : 4'b0010;
																assign node4428 = (inp[13]) ? 4'b0011 : 4'b0111;
													assign node4431 = (inp[7]) ? node4447 : node4432;
														assign node4432 = (inp[4]) ? node4440 : node4433;
															assign node4433 = (inp[2]) ? node4437 : node4434;
																assign node4434 = (inp[13]) ? 4'b0111 : 4'b0011;
																assign node4437 = (inp[13]) ? 4'b0011 : 4'b0111;
															assign node4440 = (inp[2]) ? node4444 : node4441;
																assign node4441 = (inp[13]) ? 4'b0011 : 4'b0111;
																assign node4444 = (inp[13]) ? 4'b0110 : 4'b0010;
														assign node4447 = (inp[2]) ? node4453 : node4448;
															assign node4448 = (inp[13]) ? node4450 : 4'b0101;
																assign node4450 = (inp[4]) ? 4'b0100 : 4'b0000;
															assign node4453 = (inp[4]) ? node4455 : 4'b0000;
																assign node4455 = (inp[13]) ? 4'b0001 : 4'b0101;
											assign node4458 = (inp[0]) ? node4504 : node4459;
												assign node4459 = (inp[2]) ? node4477 : node4460;
													assign node4460 = (inp[13]) ? node4470 : node4461;
														assign node4461 = (inp[12]) ? node4465 : node4462;
															assign node4462 = (inp[7]) ? 4'b0010 : 4'b0000;
															assign node4465 = (inp[7]) ? node4467 : 4'b0011;
																assign node4467 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node4470 = (inp[12]) ? node4474 : node4471;
															assign node4471 = (inp[7]) ? 4'b0110 : 4'b0100;
															assign node4474 = (inp[7]) ? 4'b0000 : 4'b0010;
													assign node4477 = (inp[13]) ? node4491 : node4478;
														assign node4478 = (inp[4]) ? node4484 : node4479;
															assign node4479 = (inp[12]) ? 4'b0111 : node4480;
																assign node4480 = (inp[7]) ? 4'b0110 : 4'b0100;
															assign node4484 = (inp[12]) ? node4488 : node4485;
																assign node4485 = (inp[7]) ? 4'b0111 : 4'b0101;
																assign node4488 = (inp[7]) ? 4'b0101 : 4'b0011;
														assign node4491 = (inp[12]) ? node4499 : node4492;
															assign node4492 = (inp[4]) ? node4496 : node4493;
																assign node4493 = (inp[7]) ? 4'b0011 : 4'b0001;
																assign node4496 = (inp[7]) ? 4'b0010 : 4'b0000;
															assign node4499 = (inp[7]) ? node4501 : 4'b0111;
																assign node4501 = (inp[4]) ? 4'b0000 : 4'b0100;
												assign node4504 = (inp[12]) ? node4526 : node4505;
													assign node4505 = (inp[7]) ? node4517 : node4506;
														assign node4506 = (inp[2]) ? node4510 : node4507;
															assign node4507 = (inp[13]) ? 4'b0101 : 4'b0001;
															assign node4510 = (inp[4]) ? node4514 : node4511;
																assign node4511 = (inp[13]) ? 4'b0001 : 4'b0101;
																assign node4514 = (inp[13]) ? 4'b0000 : 4'b0100;
														assign node4517 = (inp[2]) ? node4521 : node4518;
															assign node4518 = (inp[13]) ? 4'b0111 : 4'b0011;
															assign node4521 = (inp[4]) ? node4523 : 4'b0011;
																assign node4523 = (inp[13]) ? 4'b0010 : 4'b0110;
													assign node4526 = (inp[7]) ? node4540 : node4527;
														assign node4527 = (inp[4]) ? node4533 : node4528;
															assign node4528 = (inp[2]) ? node4530 : 4'b0010;
																assign node4530 = (inp[13]) ? 4'b0010 : 4'b0110;
															assign node4533 = (inp[2]) ? node4537 : node4534;
																assign node4534 = (inp[13]) ? 4'b0010 : 4'b0110;
																assign node4537 = (inp[13]) ? 4'b0111 : 4'b0011;
														assign node4540 = (inp[13]) ? node4548 : node4541;
															assign node4541 = (inp[4]) ? node4545 : node4542;
																assign node4542 = (inp[2]) ? 4'b0001 : 4'b0100;
																assign node4545 = (inp[2]) ? 4'b0100 : 4'b0001;
															assign node4548 = (inp[4]) ? node4550 : 4'b0101;
																assign node4550 = (inp[2]) ? 4'b0000 : 4'b0101;
									assign node4553 = (inp[9]) ? node4723 : node4554;
										assign node4554 = (inp[13]) ? node4640 : node4555;
											assign node4555 = (inp[7]) ? node4601 : node4556;
												assign node4556 = (inp[2]) ? node4578 : node4557;
													assign node4557 = (inp[12]) ? node4567 : node4558;
														assign node4558 = (inp[4]) ? node4564 : node4559;
															assign node4559 = (inp[0]) ? 4'b0000 : node4560;
																assign node4560 = (inp[1]) ? 4'b0000 : 4'b0001;
															assign node4564 = (inp[1]) ? 4'b0110 : 4'b0010;
														assign node4567 = (inp[4]) ? node4573 : node4568;
															assign node4568 = (inp[0]) ? node4570 : 4'b0011;
																assign node4570 = (inp[1]) ? 4'b0011 : 4'b0010;
															assign node4573 = (inp[1]) ? node4575 : 4'b0000;
																assign node4575 = (inp[0]) ? 4'b0000 : 4'b0001;
													assign node4578 = (inp[12]) ? node4592 : node4579;
														assign node4579 = (inp[4]) ? node4585 : node4580;
															assign node4580 = (inp[1]) ? 4'b0100 : node4581;
																assign node4581 = (inp[0]) ? 4'b0100 : 4'b0101;
															assign node4585 = (inp[1]) ? node4589 : node4586;
																assign node4586 = (inp[0]) ? 4'b0111 : 4'b0110;
																assign node4589 = (inp[0]) ? 4'b0010 : 4'b0011;
														assign node4592 = (inp[4]) ? node4598 : node4593;
															assign node4593 = (inp[0]) ? node4595 : 4'b0111;
																assign node4595 = (inp[1]) ? 4'b0111 : 4'b0110;
															assign node4598 = (inp[0]) ? 4'b0101 : 4'b0100;
												assign node4601 = (inp[2]) ? node4619 : node4602;
													assign node4602 = (inp[4]) ? node4608 : node4603;
														assign node4603 = (inp[12]) ? node4605 : 4'b0110;
															assign node4605 = (inp[1]) ? 4'b0000 : 4'b0100;
														assign node4608 = (inp[12]) ? node4614 : node4609;
															assign node4609 = (inp[0]) ? node4611 : 4'b0000;
																assign node4611 = (inp[1]) ? 4'b0001 : 4'b0000;
															assign node4614 = (inp[1]) ? 4'b0110 : node4615;
																assign node4615 = (inp[0]) ? 4'b0111 : 4'b0110;
													assign node4619 = (inp[1]) ? node4629 : node4620;
														assign node4620 = (inp[12]) ? node4624 : node4621;
															assign node4621 = (inp[4]) ? 4'b0101 : 4'b0010;
															assign node4624 = (inp[4]) ? 4'b0010 : node4625;
																assign node4625 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node4629 = (inp[0]) ? node4635 : node4630;
															assign node4630 = (inp[4]) ? 4'b0011 : node4631;
																assign node4631 = (inp[12]) ? 4'b0100 : 4'b0010;
															assign node4635 = (inp[4]) ? node4637 : 4'b0100;
																assign node4637 = (inp[12]) ? 4'b0010 : 4'b0100;
											assign node4640 = (inp[7]) ? node4682 : node4641;
												assign node4641 = (inp[2]) ? node4667 : node4642;
													assign node4642 = (inp[1]) ? node4658 : node4643;
														assign node4643 = (inp[0]) ? node4651 : node4644;
															assign node4644 = (inp[12]) ? node4648 : node4645;
																assign node4645 = (inp[4]) ? 4'b0110 : 4'b0100;
																assign node4648 = (inp[4]) ? 4'b0101 : 4'b0110;
															assign node4651 = (inp[12]) ? node4655 : node4652;
																assign node4652 = (inp[4]) ? 4'b0111 : 4'b0101;
																assign node4655 = (inp[4]) ? 4'b0101 : 4'b0111;
														assign node4658 = (inp[12]) ? node4664 : node4659;
															assign node4659 = (inp[4]) ? node4661 : 4'b0101;
																assign node4661 = (inp[0]) ? 4'b0010 : 4'b0011;
															assign node4664 = (inp[4]) ? 4'b0100 : 4'b0110;
													assign node4667 = (inp[4]) ? node4675 : node4668;
														assign node4668 = (inp[12]) ? node4670 : 4'b0001;
															assign node4670 = (inp[0]) ? 4'b0011 : node4671;
																assign node4671 = (inp[1]) ? 4'b0010 : 4'b0011;
														assign node4675 = (inp[12]) ? 4'b0000 : node4676;
															assign node4676 = (inp[1]) ? node4678 : 4'b0010;
																assign node4678 = (inp[0]) ? 4'b0111 : 4'b0110;
												assign node4682 = (inp[12]) ? node4702 : node4683;
													assign node4683 = (inp[4]) ? node4695 : node4684;
														assign node4684 = (inp[2]) ? node4690 : node4685;
															assign node4685 = (inp[1]) ? node4687 : 4'b0011;
																assign node4687 = (inp[0]) ? 4'b0010 : 4'b0011;
															assign node4690 = (inp[1]) ? node4692 : 4'b0111;
																assign node4692 = (inp[0]) ? 4'b0110 : 4'b0111;
														assign node4695 = (inp[2]) ? node4697 : 4'b0101;
															assign node4697 = (inp[0]) ? 4'b0001 : node4698;
																assign node4698 = (inp[1]) ? 4'b0001 : 4'b0000;
													assign node4702 = (inp[4]) ? node4716 : node4703;
														assign node4703 = (inp[0]) ? node4709 : node4704;
															assign node4704 = (inp[1]) ? node4706 : 4'b0001;
																assign node4706 = (inp[2]) ? 4'b0001 : 4'b0101;
															assign node4709 = (inp[2]) ? node4713 : node4710;
																assign node4710 = (inp[1]) ? 4'b0101 : 4'b0000;
																assign node4713 = (inp[1]) ? 4'b0000 : 4'b0100;
														assign node4716 = (inp[2]) ? node4720 : node4717;
															assign node4717 = (inp[1]) ? 4'b0011 : 4'b0010;
															assign node4720 = (inp[0]) ? 4'b0111 : 4'b0110;
										assign node4723 = (inp[13]) ? node4815 : node4724;
											assign node4724 = (inp[2]) ? node4768 : node4725;
												assign node4725 = (inp[7]) ? node4751 : node4726;
													assign node4726 = (inp[0]) ? node4742 : node4727;
														assign node4727 = (inp[1]) ? node4735 : node4728;
															assign node4728 = (inp[12]) ? node4732 : node4729;
																assign node4729 = (inp[4]) ? 4'b0010 : 4'b0000;
																assign node4732 = (inp[4]) ? 4'b0001 : 4'b0010;
															assign node4735 = (inp[12]) ? node4739 : node4736;
																assign node4736 = (inp[4]) ? 4'b0111 : 4'b0001;
																assign node4739 = (inp[4]) ? 4'b0000 : 4'b0010;
														assign node4742 = (inp[12]) ? node4748 : node4743;
															assign node4743 = (inp[4]) ? node4745 : 4'b0001;
																assign node4745 = (inp[1]) ? 4'b0111 : 4'b0011;
															assign node4748 = (inp[4]) ? 4'b0001 : 4'b0010;
													assign node4751 = (inp[1]) ? node4763 : node4752;
														assign node4752 = (inp[4]) ? node4758 : node4753;
															assign node4753 = (inp[12]) ? 4'b0101 : node4754;
																assign node4754 = (inp[0]) ? 4'b0111 : 4'b0110;
															assign node4758 = (inp[12]) ? node4760 : 4'b0001;
																assign node4760 = (inp[0]) ? 4'b0110 : 4'b0111;
														assign node4763 = (inp[12]) ? node4765 : 4'b0111;
															assign node4765 = (inp[4]) ? 4'b0111 : 4'b0001;
												assign node4768 = (inp[7]) ? node4794 : node4769;
													assign node4769 = (inp[12]) ? node4783 : node4770;
														assign node4770 = (inp[4]) ? node4776 : node4771;
															assign node4771 = (inp[0]) ? 4'b0101 : node4772;
																assign node4772 = (inp[1]) ? 4'b0101 : 4'b0100;
															assign node4776 = (inp[1]) ? node4780 : node4777;
																assign node4777 = (inp[0]) ? 4'b0110 : 4'b0111;
																assign node4780 = (inp[0]) ? 4'b0011 : 4'b0010;
														assign node4783 = (inp[4]) ? node4789 : node4784;
															assign node4784 = (inp[0]) ? node4786 : 4'b0110;
																assign node4786 = (inp[1]) ? 4'b0110 : 4'b0111;
															assign node4789 = (inp[0]) ? 4'b0100 : node4790;
																assign node4790 = (inp[1]) ? 4'b0101 : 4'b0100;
													assign node4794 = (inp[4]) ? node4804 : node4795;
														assign node4795 = (inp[12]) ? node4801 : node4796;
															assign node4796 = (inp[0]) ? node4798 : 4'b0011;
																assign node4798 = (inp[1]) ? 4'b0010 : 4'b0011;
															assign node4801 = (inp[0]) ? 4'b0000 : 4'b0001;
														assign node4804 = (inp[12]) ? node4810 : node4805;
															assign node4805 = (inp[0]) ? node4807 : 4'b0100;
																assign node4807 = (inp[1]) ? 4'b0101 : 4'b0100;
															assign node4810 = (inp[0]) ? 4'b0011 : node4811;
																assign node4811 = (inp[1]) ? 4'b0010 : 4'b0011;
											assign node4815 = (inp[2]) ? node4859 : node4816;
												assign node4816 = (inp[7]) ? node4840 : node4817;
													assign node4817 = (inp[0]) ? node4827 : node4818;
														assign node4818 = (inp[12]) ? node4824 : node4819;
															assign node4819 = (inp[4]) ? 4'b0010 : node4820;
																assign node4820 = (inp[1]) ? 4'b0100 : 4'b0101;
															assign node4824 = (inp[4]) ? 4'b0101 : 4'b0111;
														assign node4827 = (inp[1]) ? node4835 : node4828;
															assign node4828 = (inp[12]) ? node4832 : node4829;
																assign node4829 = (inp[4]) ? 4'b0110 : 4'b0100;
																assign node4832 = (inp[4]) ? 4'b0100 : 4'b0110;
															assign node4835 = (inp[4]) ? node4837 : 4'b0100;
																assign node4837 = (inp[12]) ? 4'b0100 : 4'b0011;
													assign node4840 = (inp[0]) ? node4850 : node4841;
														assign node4841 = (inp[4]) ? node4847 : node4842;
															assign node4842 = (inp[12]) ? node4844 : 4'b0010;
																assign node4844 = (inp[1]) ? 4'b0100 : 4'b0000;
															assign node4847 = (inp[12]) ? 4'b0010 : 4'b0100;
														assign node4850 = (inp[4]) ? node4856 : node4851;
															assign node4851 = (inp[12]) ? 4'b0100 : node4852;
																assign node4852 = (inp[1]) ? 4'b0011 : 4'b0010;
															assign node4856 = (inp[12]) ? 4'b0011 : 4'b0100;
												assign node4859 = (inp[7]) ? node4883 : node4860;
													assign node4860 = (inp[4]) ? node4872 : node4861;
														assign node4861 = (inp[12]) ? node4867 : node4862;
															assign node4862 = (inp[1]) ? node4864 : 4'b0000;
																assign node4864 = (inp[0]) ? 4'b0001 : 4'b0000;
															assign node4867 = (inp[0]) ? 4'b0010 : node4868;
																assign node4868 = (inp[1]) ? 4'b0011 : 4'b0010;
														assign node4872 = (inp[12]) ? node4878 : node4873;
															assign node4873 = (inp[0]) ? 4'b0110 : node4874;
																assign node4874 = (inp[1]) ? 4'b0111 : 4'b0011;
															assign node4878 = (inp[1]) ? 4'b0001 : node4879;
																assign node4879 = (inp[0]) ? 4'b0000 : 4'b0001;
													assign node4883 = (inp[1]) ? node4895 : node4884;
														assign node4884 = (inp[12]) ? node4890 : node4885;
															assign node4885 = (inp[4]) ? node4887 : 4'b0110;
																assign node4887 = (inp[0]) ? 4'b0000 : 4'b0001;
															assign node4890 = (inp[4]) ? 4'b0110 : node4891;
																assign node4891 = (inp[0]) ? 4'b0101 : 4'b0100;
														assign node4895 = (inp[0]) ? node4903 : node4896;
															assign node4896 = (inp[4]) ? node4900 : node4897;
																assign node4897 = (inp[12]) ? 4'b0000 : 4'b0110;
																assign node4900 = (inp[12]) ? 4'b0111 : 4'b0000;
															assign node4903 = (inp[4]) ? node4907 : node4904;
																assign node4904 = (inp[12]) ? 4'b0001 : 4'b0111;
																assign node4907 = (inp[12]) ? 4'b0110 : 4'b0000;
								assign node4910 = (inp[4]) ? node5310 : node4911;
									assign node4911 = (inp[9]) ? node5111 : node4912;
										assign node4912 = (inp[2]) ? node5010 : node4913;
											assign node4913 = (inp[12]) ? node4965 : node4914;
												assign node4914 = (inp[7]) ? node4936 : node4915;
													assign node4915 = (inp[0]) ? node4927 : node4916;
														assign node4916 = (inp[1]) ? node4920 : node4917;
															assign node4917 = (inp[13]) ? 4'b0101 : 4'b0001;
															assign node4920 = (inp[13]) ? node4924 : node4921;
																assign node4921 = (inp[15]) ? 4'b0100 : 4'b0101;
																assign node4924 = (inp[15]) ? 4'b0001 : 4'b0000;
														assign node4927 = (inp[13]) ? node4931 : node4928;
															assign node4928 = (inp[1]) ? 4'b0100 : 4'b0000;
															assign node4931 = (inp[1]) ? 4'b0000 : node4932;
																assign node4932 = (inp[15]) ? 4'b0101 : 4'b0100;
													assign node4936 = (inp[0]) ? node4950 : node4937;
														assign node4937 = (inp[1]) ? node4943 : node4938;
															assign node4938 = (inp[15]) ? node4940 : 4'b0010;
																assign node4940 = (inp[13]) ? 4'b0010 : 4'b0110;
															assign node4943 = (inp[15]) ? node4947 : node4944;
																assign node4944 = (inp[13]) ? 4'b0011 : 4'b0110;
																assign node4947 = (inp[13]) ? 4'b0110 : 4'b0011;
														assign node4950 = (inp[15]) ? node4958 : node4951;
															assign node4951 = (inp[13]) ? node4955 : node4952;
																assign node4952 = (inp[1]) ? 4'b0111 : 4'b0011;
																assign node4955 = (inp[1]) ? 4'b0011 : 4'b0111;
															assign node4958 = (inp[1]) ? node4962 : node4959;
																assign node4959 = (inp[13]) ? 4'b0010 : 4'b0111;
																assign node4962 = (inp[13]) ? 4'b0111 : 4'b0010;
												assign node4965 = (inp[7]) ? node4989 : node4966;
													assign node4966 = (inp[1]) ? node4978 : node4967;
														assign node4967 = (inp[13]) ? node4971 : node4968;
															assign node4968 = (inp[0]) ? 4'b0010 : 4'b0011;
															assign node4971 = (inp[0]) ? node4975 : node4972;
																assign node4972 = (inp[15]) ? 4'b0110 : 4'b0111;
																assign node4975 = (inp[15]) ? 4'b0111 : 4'b0110;
														assign node4978 = (inp[13]) ? node4984 : node4979;
															assign node4979 = (inp[15]) ? 4'b0111 : node4980;
																assign node4980 = (inp[0]) ? 4'b0111 : 4'b0110;
															assign node4984 = (inp[0]) ? 4'b0011 : node4985;
																assign node4985 = (inp[15]) ? 4'b0010 : 4'b0011;
													assign node4989 = (inp[13]) ? node4999 : node4990;
														assign node4990 = (inp[15]) ? node4994 : node4991;
															assign node4991 = (inp[1]) ? 4'b0100 : 4'b0101;
															assign node4994 = (inp[1]) ? 4'b0001 : node4995;
																assign node4995 = (inp[0]) ? 4'b0000 : 4'b0001;
														assign node4999 = (inp[15]) ? node5005 : node5000;
															assign node5000 = (inp[1]) ? node5002 : 4'b0000;
																assign node5002 = (inp[0]) ? 4'b0001 : 4'b0000;
															assign node5005 = (inp[1]) ? 4'b0100 : node5006;
																assign node5006 = (inp[0]) ? 4'b0101 : 4'b0100;
											assign node5010 = (inp[0]) ? node5058 : node5011;
												assign node5011 = (inp[13]) ? node5031 : node5012;
													assign node5012 = (inp[1]) ? node5022 : node5013;
														assign node5013 = (inp[7]) ? node5017 : node5014;
															assign node5014 = (inp[12]) ? 4'b0111 : 4'b0101;
															assign node5017 = (inp[12]) ? node5019 : 4'b0110;
																assign node5019 = (inp[15]) ? 4'b0101 : 4'b0001;
														assign node5022 = (inp[7]) ? node5026 : node5023;
															assign node5023 = (inp[12]) ? 4'b0011 : 4'b0000;
															assign node5026 = (inp[15]) ? node5028 : 4'b0000;
																assign node5028 = (inp[12]) ? 4'b0101 : 4'b0111;
													assign node5031 = (inp[1]) ? node5047 : node5032;
														assign node5032 = (inp[7]) ? node5040 : node5033;
															assign node5033 = (inp[12]) ? node5037 : node5034;
																assign node5034 = (inp[15]) ? 4'b0001 : 4'b0000;
																assign node5037 = (inp[15]) ? 4'b0011 : 4'b0010;
															assign node5040 = (inp[12]) ? node5044 : node5041;
																assign node5041 = (inp[15]) ? 4'b0110 : 4'b0011;
																assign node5044 = (inp[15]) ? 4'b0001 : 4'b0101;
														assign node5047 = (inp[12]) ? node5053 : node5048;
															assign node5048 = (inp[7]) ? node5050 : 4'b0101;
																assign node5050 = (inp[15]) ? 4'b0011 : 4'b0111;
															assign node5053 = (inp[7]) ? 4'b0100 : node5054;
																assign node5054 = (inp[15]) ? 4'b0110 : 4'b0111;
												assign node5058 = (inp[7]) ? node5082 : node5059;
													assign node5059 = (inp[12]) ? node5073 : node5060;
														assign node5060 = (inp[15]) ? node5066 : node5061;
															assign node5061 = (inp[1]) ? node5063 : 4'b0100;
																assign node5063 = (inp[13]) ? 4'b0100 : 4'b0000;
															assign node5066 = (inp[13]) ? node5070 : node5067;
																assign node5067 = (inp[1]) ? 4'b0001 : 4'b0100;
																assign node5070 = (inp[1]) ? 4'b0100 : 4'b0001;
														assign node5073 = (inp[13]) ? node5077 : node5074;
															assign node5074 = (inp[1]) ? 4'b0010 : 4'b0110;
															assign node5077 = (inp[1]) ? 4'b0111 : node5078;
																assign node5078 = (inp[15]) ? 4'b0011 : 4'b0010;
													assign node5082 = (inp[12]) ? node5098 : node5083;
														assign node5083 = (inp[15]) ? node5091 : node5084;
															assign node5084 = (inp[1]) ? node5088 : node5085;
																assign node5085 = (inp[13]) ? 4'b0011 : 4'b0111;
																assign node5088 = (inp[13]) ? 4'b0111 : 4'b0011;
															assign node5091 = (inp[13]) ? node5095 : node5092;
																assign node5092 = (inp[1]) ? 4'b0110 : 4'b0011;
																assign node5095 = (inp[1]) ? 4'b0011 : 4'b0110;
														assign node5098 = (inp[1]) ? node5104 : node5099;
															assign node5099 = (inp[13]) ? 4'b0100 : node5100;
																assign node5100 = (inp[15]) ? 4'b0100 : 4'b0000;
															assign node5104 = (inp[13]) ? node5108 : node5105;
																assign node5105 = (inp[15]) ? 4'b0101 : 4'b0001;
																assign node5108 = (inp[15]) ? 4'b0001 : 4'b0101;
										assign node5111 = (inp[7]) ? node5195 : node5112;
											assign node5112 = (inp[12]) ? node5150 : node5113;
												assign node5113 = (inp[15]) ? node5127 : node5114;
													assign node5114 = (inp[13]) ? node5122 : node5115;
														assign node5115 = (inp[1]) ? 4'b0001 : node5116;
															assign node5116 = (inp[0]) ? node5118 : 4'b0100;
																assign node5118 = (inp[2]) ? 4'b0101 : 4'b0001;
														assign node5122 = (inp[1]) ? 4'b0101 : node5123;
															assign node5123 = (inp[2]) ? 4'b0001 : 4'b0101;
													assign node5127 = (inp[1]) ? node5137 : node5128;
														assign node5128 = (inp[2]) ? node5134 : node5129;
															assign node5129 = (inp[13]) ? node5131 : 4'b0000;
																assign node5131 = (inp[0]) ? 4'b0100 : 4'b0101;
															assign node5134 = (inp[13]) ? 4'b0000 : 4'b0100;
														assign node5137 = (inp[13]) ? node5143 : node5138;
															assign node5138 = (inp[2]) ? node5140 : 4'b0101;
																assign node5140 = (inp[0]) ? 4'b0000 : 4'b0001;
															assign node5143 = (inp[0]) ? node5147 : node5144;
																assign node5144 = (inp[2]) ? 4'b0100 : 4'b0000;
																assign node5147 = (inp[2]) ? 4'b0101 : 4'b0001;
												assign node5150 = (inp[1]) ? node5174 : node5151;
													assign node5151 = (inp[0]) ? node5163 : node5152;
														assign node5152 = (inp[13]) ? node5156 : node5153;
															assign node5153 = (inp[2]) ? 4'b0110 : 4'b0010;
															assign node5156 = (inp[2]) ? node5160 : node5157;
																assign node5157 = (inp[15]) ? 4'b0111 : 4'b0110;
																assign node5160 = (inp[15]) ? 4'b0010 : 4'b0011;
														assign node5163 = (inp[13]) ? node5167 : node5164;
															assign node5164 = (inp[2]) ? 4'b0111 : 4'b0011;
															assign node5167 = (inp[15]) ? node5171 : node5168;
																assign node5168 = (inp[2]) ? 4'b0011 : 4'b0111;
																assign node5171 = (inp[2]) ? 4'b0010 : 4'b0110;
													assign node5174 = (inp[15]) ? node5182 : node5175;
														assign node5175 = (inp[2]) ? node5179 : node5176;
															assign node5176 = (inp[13]) ? 4'b0010 : 4'b0110;
															assign node5179 = (inp[13]) ? 4'b0110 : 4'b0010;
														assign node5182 = (inp[13]) ? node5188 : node5183;
															assign node5183 = (inp[2]) ? node5185 : 4'b0110;
																assign node5185 = (inp[0]) ? 4'b0011 : 4'b0010;
															assign node5188 = (inp[0]) ? node5192 : node5189;
																assign node5189 = (inp[2]) ? 4'b0111 : 4'b0011;
																assign node5192 = (inp[2]) ? 4'b0110 : 4'b0010;
											assign node5195 = (inp[12]) ? node5251 : node5196;
												assign node5196 = (inp[0]) ? node5224 : node5197;
													assign node5197 = (inp[2]) ? node5209 : node5198;
														assign node5198 = (inp[13]) ? node5204 : node5199;
															assign node5199 = (inp[15]) ? 4'b0111 : node5200;
																assign node5200 = (inp[1]) ? 4'b0111 : 4'b0011;
															assign node5204 = (inp[15]) ? node5206 : 4'b0010;
																assign node5206 = (inp[1]) ? 4'b0111 : 4'b0011;
														assign node5209 = (inp[1]) ? node5217 : node5210;
															assign node5210 = (inp[13]) ? node5214 : node5211;
																assign node5211 = (inp[15]) ? 4'b0010 : 4'b0111;
																assign node5214 = (inp[15]) ? 4'b0111 : 4'b0010;
															assign node5217 = (inp[13]) ? node5221 : node5218;
																assign node5218 = (inp[15]) ? 4'b0110 : 4'b0010;
																assign node5221 = (inp[15]) ? 4'b0010 : 4'b0110;
													assign node5224 = (inp[15]) ? node5238 : node5225;
														assign node5225 = (inp[13]) ? node5231 : node5226;
															assign node5226 = (inp[1]) ? node5228 : 4'b0110;
																assign node5228 = (inp[2]) ? 4'b0010 : 4'b0110;
															assign node5231 = (inp[2]) ? node5235 : node5232;
																assign node5232 = (inp[1]) ? 4'b0010 : 4'b0110;
																assign node5235 = (inp[1]) ? 4'b0110 : 4'b0010;
														assign node5238 = (inp[1]) ? node5244 : node5239;
															assign node5239 = (inp[13]) ? 4'b0111 : node5240;
																assign node5240 = (inp[2]) ? 4'b0010 : 4'b0110;
															assign node5244 = (inp[13]) ? node5248 : node5245;
																assign node5245 = (inp[2]) ? 4'b0111 : 4'b0011;
																assign node5248 = (inp[2]) ? 4'b0010 : 4'b0110;
												assign node5251 = (inp[1]) ? node5279 : node5252;
													assign node5252 = (inp[0]) ? node5266 : node5253;
														assign node5253 = (inp[15]) ? node5261 : node5254;
															assign node5254 = (inp[13]) ? node5258 : node5255;
																assign node5255 = (inp[2]) ? 4'b0000 : 4'b0100;
																assign node5258 = (inp[2]) ? 4'b0100 : 4'b0000;
															assign node5261 = (inp[13]) ? 4'b0000 : node5262;
																assign node5262 = (inp[2]) ? 4'b0100 : 4'b0000;
														assign node5266 = (inp[2]) ? node5274 : node5267;
															assign node5267 = (inp[15]) ? node5271 : node5268;
																assign node5268 = (inp[13]) ? 4'b0001 : 4'b0100;
																assign node5271 = (inp[13]) ? 4'b0100 : 4'b0001;
															assign node5274 = (inp[13]) ? node5276 : 4'b0101;
																assign node5276 = (inp[15]) ? 4'b0000 : 4'b0101;
													assign node5279 = (inp[0]) ? node5295 : node5280;
														assign node5280 = (inp[13]) ? node5288 : node5281;
															assign node5281 = (inp[15]) ? node5285 : node5282;
																assign node5282 = (inp[2]) ? 4'b0001 : 4'b0101;
																assign node5285 = (inp[2]) ? 4'b0100 : 4'b0000;
															assign node5288 = (inp[15]) ? node5292 : node5289;
																assign node5289 = (inp[2]) ? 4'b0101 : 4'b0001;
																assign node5292 = (inp[2]) ? 4'b0001 : 4'b0101;
														assign node5295 = (inp[2]) ? node5303 : node5296;
															assign node5296 = (inp[13]) ? node5300 : node5297;
																assign node5297 = (inp[15]) ? 4'b0000 : 4'b0101;
																assign node5300 = (inp[15]) ? 4'b0101 : 4'b0000;
															assign node5303 = (inp[13]) ? node5307 : node5304;
																assign node5304 = (inp[15]) ? 4'b0100 : 4'b0000;
																assign node5307 = (inp[15]) ? 4'b0000 : 4'b0100;
									assign node5310 = (inp[9]) ? node5490 : node5311;
										assign node5311 = (inp[13]) ? node5393 : node5312;
											assign node5312 = (inp[7]) ? node5354 : node5313;
												assign node5313 = (inp[2]) ? node5335 : node5314;
													assign node5314 = (inp[12]) ? node5324 : node5315;
														assign node5315 = (inp[15]) ? node5319 : node5316;
															assign node5316 = (inp[1]) ? 4'b0100 : 4'b0000;
															assign node5319 = (inp[0]) ? node5321 : 4'b0110;
																assign node5321 = (inp[1]) ? 4'b0111 : 4'b0110;
														assign node5324 = (inp[15]) ? node5330 : node5325;
															assign node5325 = (inp[1]) ? node5327 : 4'b0110;
																assign node5327 = (inp[0]) ? 4'b0010 : 4'b0011;
															assign node5330 = (inp[1]) ? 4'b0100 : node5331;
																assign node5331 = (inp[0]) ? 4'b0001 : 4'b0000;
													assign node5335 = (inp[15]) ? node5347 : node5336;
														assign node5336 = (inp[12]) ? node5340 : node5337;
															assign node5337 = (inp[1]) ? 4'b0001 : 4'b0101;
															assign node5340 = (inp[1]) ? node5344 : node5341;
																assign node5341 = (inp[0]) ? 4'b0010 : 4'b0011;
																assign node5344 = (inp[0]) ? 4'b0111 : 4'b0110;
														assign node5347 = (inp[12]) ? node5349 : 4'b0010;
															assign node5349 = (inp[1]) ? 4'b0000 : node5350;
																assign node5350 = (inp[0]) ? 4'b0100 : 4'b0101;
												assign node5354 = (inp[2]) ? node5370 : node5355;
													assign node5355 = (inp[15]) ? node5363 : node5356;
														assign node5356 = (inp[12]) ? node5360 : node5357;
															assign node5357 = (inp[1]) ? 4'b0111 : 4'b0011;
															assign node5360 = (inp[1]) ? 4'b0001 : 4'b0000;
														assign node5363 = (inp[12]) ? node5367 : node5364;
															assign node5364 = (inp[0]) ? 4'b0000 : 4'b0001;
															assign node5367 = (inp[1]) ? 4'b0010 : 4'b0110;
													assign node5370 = (inp[15]) ? node5380 : node5371;
														assign node5371 = (inp[12]) ? node5377 : node5372;
															assign node5372 = (inp[1]) ? node5374 : 4'b0110;
																assign node5374 = (inp[0]) ? 4'b0011 : 4'b0010;
															assign node5377 = (inp[1]) ? 4'b0100 : 4'b0101;
														assign node5380 = (inp[12]) ? node5388 : node5381;
															assign node5381 = (inp[1]) ? node5385 : node5382;
																assign node5382 = (inp[0]) ? 4'b0101 : 4'b0100;
																assign node5385 = (inp[0]) ? 4'b0000 : 4'b0001;
															assign node5388 = (inp[1]) ? 4'b0111 : node5389;
																assign node5389 = (inp[0]) ? 4'b0010 : 4'b0011;
											assign node5393 = (inp[2]) ? node5435 : node5394;
												assign node5394 = (inp[7]) ? node5414 : node5395;
													assign node5395 = (inp[15]) ? node5409 : node5396;
														assign node5396 = (inp[12]) ? node5402 : node5397;
															assign node5397 = (inp[1]) ? node5399 : 4'b0100;
																assign node5399 = (inp[0]) ? 4'b0001 : 4'b0000;
															assign node5402 = (inp[1]) ? node5406 : node5403;
																assign node5403 = (inp[0]) ? 4'b0011 : 4'b0010;
																assign node5406 = (inp[0]) ? 4'b0110 : 4'b0111;
														assign node5409 = (inp[1]) ? node5411 : 4'b0011;
															assign node5411 = (inp[12]) ? 4'b0000 : 4'b0010;
													assign node5414 = (inp[1]) ? node5426 : node5415;
														assign node5415 = (inp[12]) ? node5421 : node5416;
															assign node5416 = (inp[15]) ? node5418 : 4'b0111;
																assign node5418 = (inp[0]) ? 4'b0101 : 4'b0100;
															assign node5421 = (inp[15]) ? node5423 : 4'b0100;
																assign node5423 = (inp[0]) ? 4'b0010 : 4'b0011;
														assign node5426 = (inp[12]) ? node5432 : node5427;
															assign node5427 = (inp[15]) ? 4'b0001 : node5428;
																assign node5428 = (inp[0]) ? 4'b0010 : 4'b0011;
															assign node5432 = (inp[15]) ? 4'b0111 : 4'b0101;
												assign node5435 = (inp[7]) ? node5461 : node5436;
													assign node5436 = (inp[1]) ? node5450 : node5437;
														assign node5437 = (inp[0]) ? node5443 : node5438;
															assign node5438 = (inp[12]) ? node5440 : 4'b0001;
																assign node5440 = (inp[15]) ? 4'b0001 : 4'b0111;
															assign node5443 = (inp[15]) ? node5447 : node5444;
																assign node5444 = (inp[12]) ? 4'b0110 : 4'b0000;
																assign node5447 = (inp[12]) ? 4'b0001 : 4'b0111;
														assign node5450 = (inp[12]) ? node5456 : node5451;
															assign node5451 = (inp[15]) ? 4'b0111 : node5452;
																assign node5452 = (inp[0]) ? 4'b0100 : 4'b0101;
															assign node5456 = (inp[15]) ? node5458 : 4'b0011;
																assign node5458 = (inp[0]) ? 4'b0101 : 4'b0100;
													assign node5461 = (inp[0]) ? node5475 : node5462;
														assign node5462 = (inp[1]) ? node5468 : node5463;
															assign node5463 = (inp[12]) ? 4'b0001 : node5464;
																assign node5464 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node5468 = (inp[12]) ? node5472 : node5469;
																assign node5469 = (inp[15]) ? 4'b0100 : 4'b0110;
																assign node5472 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node5475 = (inp[1]) ? node5483 : node5476;
															assign node5476 = (inp[12]) ? node5480 : node5477;
																assign node5477 = (inp[15]) ? 4'b0000 : 4'b0011;
																assign node5480 = (inp[15]) ? 4'b0111 : 4'b0000;
															assign node5483 = (inp[12]) ? node5487 : node5484;
																assign node5484 = (inp[15]) ? 4'b0101 : 4'b0111;
																assign node5487 = (inp[15]) ? 4'b0011 : 4'b0001;
										assign node5490 = (inp[13]) ? node5578 : node5491;
											assign node5491 = (inp[15]) ? node5531 : node5492;
												assign node5492 = (inp[2]) ? node5510 : node5493;
													assign node5493 = (inp[7]) ? node5503 : node5494;
														assign node5494 = (inp[12]) ? node5498 : node5495;
															assign node5495 = (inp[1]) ? 4'b0101 : 4'b0001;
															assign node5498 = (inp[1]) ? node5500 : 4'b0111;
																assign node5500 = (inp[0]) ? 4'b0011 : 4'b0010;
														assign node5503 = (inp[12]) ? node5507 : node5504;
															assign node5504 = (inp[1]) ? 4'b0110 : 4'b0010;
															assign node5507 = (inp[1]) ? 4'b0000 : 4'b0001;
													assign node5510 = (inp[1]) ? node5518 : node5511;
														assign node5511 = (inp[12]) ? node5515 : node5512;
															assign node5512 = (inp[7]) ? 4'b0111 : 4'b0100;
															assign node5515 = (inp[7]) ? 4'b0100 : 4'b0010;
														assign node5518 = (inp[12]) ? node5526 : node5519;
															assign node5519 = (inp[7]) ? node5523 : node5520;
																assign node5520 = (inp[0]) ? 4'b0001 : 4'b0000;
																assign node5523 = (inp[0]) ? 4'b0010 : 4'b0011;
															assign node5526 = (inp[7]) ? 4'b0101 : node5527;
																assign node5527 = (inp[0]) ? 4'b0110 : 4'b0111;
												assign node5531 = (inp[2]) ? node5551 : node5532;
													assign node5532 = (inp[7]) ? node5542 : node5533;
														assign node5533 = (inp[12]) ? node5539 : node5534;
															assign node5534 = (inp[1]) ? node5536 : 4'b0111;
																assign node5536 = (inp[0]) ? 4'b0110 : 4'b0111;
															assign node5539 = (inp[1]) ? 4'b0101 : 4'b0001;
														assign node5542 = (inp[12]) ? node5548 : node5543;
															assign node5543 = (inp[1]) ? 4'b0101 : node5544;
																assign node5544 = (inp[0]) ? 4'b0001 : 4'b0000;
															assign node5548 = (inp[1]) ? 4'b0011 : 4'b0111;
													assign node5551 = (inp[0]) ? node5567 : node5552;
														assign node5552 = (inp[12]) ? node5560 : node5553;
															assign node5553 = (inp[7]) ? node5557 : node5554;
																assign node5554 = (inp[1]) ? 4'b0011 : 4'b0010;
																assign node5557 = (inp[1]) ? 4'b0000 : 4'b0101;
															assign node5560 = (inp[7]) ? node5564 : node5561;
																assign node5561 = (inp[1]) ? 4'b0000 : 4'b0100;
																assign node5564 = (inp[1]) ? 4'b0110 : 4'b0010;
														assign node5567 = (inp[12]) ? node5571 : node5568;
															assign node5568 = (inp[7]) ? 4'b0001 : 4'b0011;
															assign node5571 = (inp[7]) ? node5575 : node5572;
																assign node5572 = (inp[1]) ? 4'b0001 : 4'b0101;
																assign node5575 = (inp[1]) ? 4'b0110 : 4'b0011;
											assign node5578 = (inp[12]) ? node5628 : node5579;
												assign node5579 = (inp[0]) ? node5609 : node5580;
													assign node5580 = (inp[2]) ? node5596 : node5581;
														assign node5581 = (inp[1]) ? node5589 : node5582;
															assign node5582 = (inp[7]) ? node5586 : node5583;
																assign node5583 = (inp[15]) ? 4'b0010 : 4'b0101;
																assign node5586 = (inp[15]) ? 4'b0101 : 4'b0110;
															assign node5589 = (inp[7]) ? node5593 : node5590;
																assign node5590 = (inp[15]) ? 4'b0011 : 4'b0001;
																assign node5593 = (inp[15]) ? 4'b0000 : 4'b0010;
														assign node5596 = (inp[1]) ? node5604 : node5597;
															assign node5597 = (inp[7]) ? node5601 : node5598;
																assign node5598 = (inp[15]) ? 4'b0111 : 4'b0000;
																assign node5601 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node5604 = (inp[7]) ? node5606 : 4'b0110;
																assign node5606 = (inp[15]) ? 4'b0101 : 4'b0111;
													assign node5609 = (inp[7]) ? node5617 : node5610;
														assign node5610 = (inp[15]) ? node5614 : node5611;
															assign node5611 = (inp[2]) ? 4'b0001 : 4'b0000;
															assign node5614 = (inp[2]) ? 4'b0110 : 4'b0011;
														assign node5617 = (inp[15]) ? node5625 : node5618;
															assign node5618 = (inp[2]) ? node5622 : node5619;
																assign node5619 = (inp[1]) ? 4'b0011 : 4'b0110;
																assign node5622 = (inp[1]) ? 4'b0110 : 4'b0010;
															assign node5625 = (inp[2]) ? 4'b0001 : 4'b0100;
												assign node5628 = (inp[2]) ? node5658 : node5629;
													assign node5629 = (inp[0]) ? node5643 : node5630;
														assign node5630 = (inp[1]) ? node5636 : node5631;
															assign node5631 = (inp[15]) ? node5633 : 4'b0011;
																assign node5633 = (inp[7]) ? 4'b0010 : 4'b0100;
															assign node5636 = (inp[15]) ? node5640 : node5637;
																assign node5637 = (inp[7]) ? 4'b0100 : 4'b0110;
																assign node5640 = (inp[7]) ? 4'b0110 : 4'b0000;
														assign node5643 = (inp[1]) ? node5651 : node5644;
															assign node5644 = (inp[15]) ? node5648 : node5645;
																assign node5645 = (inp[7]) ? 4'b0101 : 4'b0010;
																assign node5648 = (inp[7]) ? 4'b0011 : 4'b0101;
															assign node5651 = (inp[7]) ? node5655 : node5652;
																assign node5652 = (inp[15]) ? 4'b0001 : 4'b0111;
																assign node5655 = (inp[15]) ? 4'b0110 : 4'b0100;
													assign node5658 = (inp[7]) ? node5670 : node5659;
														assign node5659 = (inp[15]) ? node5665 : node5660;
															assign node5660 = (inp[1]) ? 4'b0010 : node5661;
																assign node5661 = (inp[0]) ? 4'b0111 : 4'b0110;
															assign node5665 = (inp[1]) ? node5667 : 4'b0000;
																assign node5667 = (inp[0]) ? 4'b0100 : 4'b0101;
														assign node5670 = (inp[15]) ? node5678 : node5671;
															assign node5671 = (inp[0]) ? node5675 : node5672;
																assign node5672 = (inp[1]) ? 4'b0001 : 4'b0000;
																assign node5675 = (inp[1]) ? 4'b0000 : 4'b0001;
															assign node5678 = (inp[1]) ? node5680 : 4'b0111;
																assign node5680 = (inp[0]) ? 4'b0010 : 4'b0011;
					assign node5683 = (inp[11]) ? node7133 : node5684;
						assign node5684 = (inp[9]) ? node6394 : node5685;
							assign node5685 = (inp[12]) ? node5965 : node5686;
								assign node5686 = (inp[2]) ? node5802 : node5687;
									assign node5687 = (inp[5]) ? node5731 : node5688;
										assign node5688 = (inp[13]) ? node5710 : node5689;
											assign node5689 = (inp[15]) ? node5693 : node5690;
												assign node5690 = (inp[7]) ? 4'b1010 : 4'b1000;
												assign node5693 = (inp[7]) ? node5703 : node5694;
													assign node5694 = (inp[1]) ? node5696 : 4'b1010;
														assign node5696 = (inp[4]) ? node5700 : node5697;
															assign node5697 = (inp[0]) ? 4'b1011 : 4'b1010;
															assign node5700 = (inp[0]) ? 4'b1111 : 4'b1110;
													assign node5703 = (inp[1]) ? 4'b1001 : node5704;
														assign node5704 = (inp[4]) ? node5706 : 4'b1100;
															assign node5706 = (inp[0]) ? 4'b1001 : 4'b1000;
											assign node5710 = (inp[15]) ? node5714 : node5711;
												assign node5711 = (inp[7]) ? 4'b1110 : 4'b1100;
												assign node5714 = (inp[7]) ? node5722 : node5715;
													assign node5715 = (inp[1]) ? node5717 : 4'b1111;
														assign node5717 = (inp[4]) ? 4'b1010 : node5718;
															assign node5718 = (inp[0]) ? 4'b1110 : 4'b1111;
													assign node5722 = (inp[1]) ? 4'b1100 : node5723;
														assign node5723 = (inp[4]) ? node5727 : node5724;
															assign node5724 = (inp[0]) ? 4'b1000 : 4'b1001;
															assign node5727 = (inp[0]) ? 4'b1100 : 4'b1101;
										assign node5731 = (inp[13]) ? node5765 : node5732;
											assign node5732 = (inp[15]) ? node5744 : node5733;
												assign node5733 = (inp[7]) ? node5739 : node5734;
													assign node5734 = (inp[4]) ? node5736 : 4'b1100;
														assign node5736 = (inp[0]) ? 4'b1101 : 4'b1100;
													assign node5739 = (inp[0]) ? node5741 : 4'b1111;
														assign node5741 = (inp[4]) ? 4'b1110 : 4'b1111;
												assign node5744 = (inp[7]) ? node5754 : node5745;
													assign node5745 = (inp[1]) ? node5747 : 4'b1110;
														assign node5747 = (inp[4]) ? node5751 : node5748;
															assign node5748 = (inp[0]) ? 4'b1111 : 4'b1110;
															assign node5751 = (inp[0]) ? 4'b1010 : 4'b1011;
													assign node5754 = (inp[1]) ? node5760 : node5755;
														assign node5755 = (inp[4]) ? 4'b1100 : node5756;
															assign node5756 = (inp[0]) ? 4'b1000 : 4'b1001;
														assign node5760 = (inp[0]) ? node5762 : 4'b1100;
															assign node5762 = (inp[4]) ? 4'b1101 : 4'b1100;
											assign node5765 = (inp[15]) ? node5777 : node5766;
												assign node5766 = (inp[7]) ? node5772 : node5767;
													assign node5767 = (inp[0]) ? 4'b1001 : node5768;
														assign node5768 = (inp[4]) ? 4'b1001 : 4'b1000;
													assign node5772 = (inp[4]) ? 4'b1010 : node5773;
														assign node5773 = (inp[0]) ? 4'b1010 : 4'b1011;
												assign node5777 = (inp[7]) ? node5789 : node5778;
													assign node5778 = (inp[1]) ? node5784 : node5779;
														assign node5779 = (inp[4]) ? 4'b1010 : node5780;
															assign node5780 = (inp[0]) ? 4'b1010 : 4'b1011;
														assign node5784 = (inp[4]) ? node5786 : 4'b1010;
															assign node5786 = (inp[0]) ? 4'b1111 : 4'b1110;
													assign node5789 = (inp[4]) ? node5797 : node5790;
														assign node5790 = (inp[1]) ? node5794 : node5791;
															assign node5791 = (inp[0]) ? 4'b1101 : 4'b1100;
															assign node5794 = (inp[0]) ? 4'b1000 : 4'b1001;
														assign node5797 = (inp[1]) ? 4'b1000 : node5798;
															assign node5798 = (inp[0]) ? 4'b1000 : 4'b1001;
									assign node5802 = (inp[15]) ? node5870 : node5803;
										assign node5803 = (inp[7]) ? node5835 : node5804;
											assign node5804 = (inp[4]) ? node5820 : node5805;
												assign node5805 = (inp[0]) ? node5813 : node5806;
													assign node5806 = (inp[5]) ? node5810 : node5807;
														assign node5807 = (inp[13]) ? 4'b1100 : 4'b1000;
														assign node5810 = (inp[13]) ? 4'b1001 : 4'b1100;
													assign node5813 = (inp[5]) ? node5817 : node5814;
														assign node5814 = (inp[13]) ? 4'b1101 : 4'b1001;
														assign node5817 = (inp[13]) ? 4'b1001 : 4'b1101;
												assign node5820 = (inp[0]) ? node5828 : node5821;
													assign node5821 = (inp[5]) ? node5825 : node5822;
														assign node5822 = (inp[13]) ? 4'b1101 : 4'b1001;
														assign node5825 = (inp[13]) ? 4'b1000 : 4'b1100;
													assign node5828 = (inp[5]) ? node5832 : node5829;
														assign node5829 = (inp[13]) ? 4'b1100 : 4'b1000;
														assign node5832 = (inp[13]) ? 4'b1001 : 4'b1100;
											assign node5835 = (inp[13]) ? node5849 : node5836;
												assign node5836 = (inp[5]) ? node5844 : node5837;
													assign node5837 = (inp[4]) ? node5841 : node5838;
														assign node5838 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node5841 = (inp[0]) ? 4'b1010 : 4'b1011;
													assign node5844 = (inp[4]) ? 4'b1111 : node5845;
														assign node5845 = (inp[0]) ? 4'b1110 : 4'b1111;
												assign node5849 = (inp[5]) ? node5865 : node5850;
													assign node5850 = (inp[1]) ? node5858 : node5851;
														assign node5851 = (inp[4]) ? node5855 : node5852;
															assign node5852 = (inp[0]) ? 4'b1111 : 4'b1110;
															assign node5855 = (inp[0]) ? 4'b1110 : 4'b1111;
														assign node5858 = (inp[4]) ? node5862 : node5859;
															assign node5859 = (inp[0]) ? 4'b1111 : 4'b1110;
															assign node5862 = (inp[0]) ? 4'b1110 : 4'b1111;
													assign node5865 = (inp[0]) ? 4'b1010 : node5866;
														assign node5866 = (inp[4]) ? 4'b1011 : 4'b1010;
										assign node5870 = (inp[7]) ? node5922 : node5871;
											assign node5871 = (inp[13]) ? node5893 : node5872;
												assign node5872 = (inp[5]) ? node5884 : node5873;
													assign node5873 = (inp[4]) ? node5879 : node5874;
														assign node5874 = (inp[1]) ? 4'b1011 : node5875;
															assign node5875 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node5879 = (inp[1]) ? 4'b1110 : node5880;
															assign node5880 = (inp[0]) ? 4'b1010 : 4'b1011;
													assign node5884 = (inp[1]) ? node5890 : node5885;
														assign node5885 = (inp[4]) ? 4'b1110 : node5886;
															assign node5886 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node5890 = (inp[4]) ? 4'b1011 : 4'b1111;
												assign node5893 = (inp[5]) ? node5913 : node5894;
													assign node5894 = (inp[1]) ? node5908 : node5895;
														assign node5895 = (inp[10]) ? node5903 : node5896;
															assign node5896 = (inp[0]) ? node5900 : node5897;
																assign node5897 = (inp[4]) ? 4'b1110 : 4'b1111;
																assign node5900 = (inp[4]) ? 4'b1111 : 4'b1110;
															assign node5903 = (inp[0]) ? node5905 : 4'b1110;
																assign node5905 = (inp[4]) ? 4'b1111 : 4'b1110;
														assign node5908 = (inp[4]) ? node5910 : 4'b1110;
															assign node5910 = (inp[0]) ? 4'b1010 : 4'b1011;
													assign node5913 = (inp[4]) ? node5919 : node5914;
														assign node5914 = (inp[1]) ? node5916 : 4'b1010;
															assign node5916 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node5919 = (inp[1]) ? 4'b1110 : 4'b1010;
											assign node5922 = (inp[13]) ? node5948 : node5923;
												assign node5923 = (inp[5]) ? node5937 : node5924;
													assign node5924 = (inp[1]) ? node5930 : node5925;
														assign node5925 = (inp[4]) ? 4'b1000 : node5926;
															assign node5926 = (inp[0]) ? 4'b1101 : 4'b1100;
														assign node5930 = (inp[4]) ? node5934 : node5931;
															assign node5931 = (inp[0]) ? 4'b1000 : 4'b1001;
															assign node5934 = (inp[0]) ? 4'b1001 : 4'b1000;
													assign node5937 = (inp[4]) ? node5943 : node5938;
														assign node5938 = (inp[1]) ? node5940 : 4'b1000;
															assign node5940 = (inp[0]) ? 4'b1101 : 4'b1100;
														assign node5943 = (inp[1]) ? 4'b1100 : node5944;
															assign node5944 = (inp[0]) ? 4'b1100 : 4'b1101;
												assign node5948 = (inp[1]) ? node5956 : node5949;
													assign node5949 = (inp[5]) ? node5953 : node5950;
														assign node5950 = (inp[4]) ? 4'b1101 : 4'b1000;
														assign node5953 = (inp[4]) ? 4'b1001 : 4'b1101;
													assign node5956 = (inp[5]) ? 4'b1000 : node5957;
														assign node5957 = (inp[0]) ? node5961 : node5958;
															assign node5958 = (inp[4]) ? 4'b1101 : 4'b1100;
															assign node5961 = (inp[4]) ? 4'b1100 : 4'b1101;
								assign node5965 = (inp[2]) ? node6169 : node5966;
									assign node5966 = (inp[7]) ? node6062 : node5967;
										assign node5967 = (inp[15]) ? node6019 : node5968;
											assign node5968 = (inp[1]) ? node5988 : node5969;
												assign node5969 = (inp[5]) ? node5979 : node5970;
													assign node5970 = (inp[13]) ? node5974 : node5971;
														assign node5971 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node5974 = (inp[4]) ? node5976 : 4'b1100;
															assign node5976 = (inp[0]) ? 4'b1001 : 4'b1000;
													assign node5979 = (inp[4]) ? node5985 : node5980;
														assign node5980 = (inp[13]) ? node5982 : 4'b1100;
															assign node5982 = (inp[0]) ? 4'b1001 : 4'b1000;
														assign node5985 = (inp[13]) ? 4'b1101 : 4'b1001;
												assign node5988 = (inp[0]) ? node6004 : node5989;
													assign node5989 = (inp[4]) ? node5997 : node5990;
														assign node5990 = (inp[5]) ? node5994 : node5991;
															assign node5991 = (inp[13]) ? 4'b1001 : 4'b1101;
															assign node5994 = (inp[13]) ? 4'b1101 : 4'b1001;
														assign node5997 = (inp[5]) ? node6001 : node5998;
															assign node5998 = (inp[13]) ? 4'b1101 : 4'b1001;
															assign node6001 = (inp[13]) ? 4'b1000 : 4'b1100;
													assign node6004 = (inp[13]) ? node6012 : node6005;
														assign node6005 = (inp[4]) ? node6009 : node6006;
															assign node6006 = (inp[5]) ? 4'b1000 : 4'b1101;
															assign node6009 = (inp[5]) ? 4'b1100 : 4'b1000;
														assign node6012 = (inp[5]) ? node6016 : node6013;
															assign node6013 = (inp[4]) ? 4'b1100 : 4'b1000;
															assign node6016 = (inp[4]) ? 4'b1001 : 4'b1100;
											assign node6019 = (inp[13]) ? node6041 : node6020;
												assign node6020 = (inp[5]) ? node6032 : node6021;
													assign node6021 = (inp[1]) ? node6027 : node6022;
														assign node6022 = (inp[4]) ? node6024 : 4'b1010;
															assign node6024 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node6027 = (inp[4]) ? 4'b1010 : node6028;
															assign node6028 = (inp[0]) ? 4'b1110 : 4'b1111;
													assign node6032 = (inp[4]) ? node6036 : node6033;
														assign node6033 = (inp[1]) ? 4'b1010 : 4'b1110;
														assign node6036 = (inp[1]) ? node6038 : 4'b1111;
															assign node6038 = (inp[0]) ? 4'b1111 : 4'b1110;
												assign node6041 = (inp[5]) ? node6051 : node6042;
													assign node6042 = (inp[4]) ? node6046 : node6043;
														assign node6043 = (inp[1]) ? 4'b1011 : 4'b1111;
														assign node6046 = (inp[1]) ? 4'b1111 : node6047;
															assign node6047 = (inp[0]) ? 4'b1110 : 4'b1111;
													assign node6051 = (inp[4]) ? node6057 : node6052;
														assign node6052 = (inp[1]) ? 4'b1111 : node6053;
															assign node6053 = (inp[0]) ? 4'b1010 : 4'b1011;
														assign node6057 = (inp[0]) ? node6059 : 4'b1010;
															assign node6059 = (inp[1]) ? 4'b1010 : 4'b1011;
										assign node6062 = (inp[15]) ? node6126 : node6063;
											assign node6063 = (inp[0]) ? node6095 : node6064;
												assign node6064 = (inp[13]) ? node6080 : node6065;
													assign node6065 = (inp[1]) ? node6073 : node6066;
														assign node6066 = (inp[5]) ? node6070 : node6067;
															assign node6067 = (inp[4]) ? 4'b1110 : 4'b1010;
															assign node6070 = (inp[4]) ? 4'b1010 : 4'b1111;
														assign node6073 = (inp[5]) ? node6077 : node6074;
															assign node6074 = (inp[4]) ? 4'b1010 : 4'b1111;
															assign node6077 = (inp[4]) ? 4'b1111 : 4'b1011;
													assign node6080 = (inp[4]) ? node6088 : node6081;
														assign node6081 = (inp[1]) ? node6085 : node6082;
															assign node6082 = (inp[5]) ? 4'b1010 : 4'b1110;
															assign node6085 = (inp[5]) ? 4'b1111 : 4'b1010;
														assign node6088 = (inp[5]) ? node6092 : node6089;
															assign node6089 = (inp[1]) ? 4'b1110 : 4'b1011;
															assign node6092 = (inp[1]) ? 4'b1010 : 4'b1110;
												assign node6095 = (inp[1]) ? node6111 : node6096;
													assign node6096 = (inp[5]) ? node6104 : node6097;
														assign node6097 = (inp[4]) ? node6101 : node6098;
															assign node6098 = (inp[13]) ? 4'b1111 : 4'b1011;
															assign node6101 = (inp[13]) ? 4'b1011 : 4'b1111;
														assign node6104 = (inp[4]) ? node6108 : node6105;
															assign node6105 = (inp[13]) ? 4'b1010 : 4'b1110;
															assign node6108 = (inp[13]) ? 4'b1111 : 4'b1011;
													assign node6111 = (inp[4]) ? node6119 : node6112;
														assign node6112 = (inp[5]) ? node6116 : node6113;
															assign node6113 = (inp[13]) ? 4'b1010 : 4'b1110;
															assign node6116 = (inp[13]) ? 4'b1111 : 4'b1011;
														assign node6119 = (inp[13]) ? node6123 : node6120;
															assign node6120 = (inp[5]) ? 4'b1110 : 4'b1010;
															assign node6123 = (inp[5]) ? 4'b1010 : 4'b1110;
											assign node6126 = (inp[13]) ? node6148 : node6127;
												assign node6127 = (inp[5]) ? node6137 : node6128;
													assign node6128 = (inp[4]) ? node6134 : node6129;
														assign node6129 = (inp[1]) ? node6131 : 4'b1001;
															assign node6131 = (inp[0]) ? 4'b1001 : 4'b1000;
														assign node6134 = (inp[1]) ? 4'b1001 : 4'b1101;
													assign node6137 = (inp[4]) ? node6143 : node6138;
														assign node6138 = (inp[1]) ? node6140 : 4'b1100;
															assign node6140 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node6143 = (inp[1]) ? node6145 : 4'b1001;
															assign node6145 = (inp[0]) ? 4'b1101 : 4'b1100;
												assign node6148 = (inp[5]) ? node6160 : node6149;
													assign node6149 = (inp[1]) ? node6155 : node6150;
														assign node6150 = (inp[4]) ? node6152 : 4'b1100;
															assign node6152 = (inp[0]) ? 4'b1001 : 4'b1000;
														assign node6155 = (inp[4]) ? 4'b1100 : node6156;
															assign node6156 = (inp[0]) ? 4'b1100 : 4'b1101;
													assign node6160 = (inp[4]) ? node6166 : node6161;
														assign node6161 = (inp[0]) ? node6163 : 4'b1001;
															assign node6163 = (inp[1]) ? 4'b1001 : 4'b1000;
														assign node6166 = (inp[1]) ? 4'b1000 : 4'b1100;
									assign node6169 = (inp[5]) ? node6275 : node6170;
										assign node6170 = (inp[13]) ? node6220 : node6171;
											assign node6171 = (inp[15]) ? node6195 : node6172;
												assign node6172 = (inp[7]) ? node6186 : node6173;
													assign node6173 = (inp[4]) ? node6181 : node6174;
														assign node6174 = (inp[1]) ? node6178 : node6175;
															assign node6175 = (inp[0]) ? 4'b1001 : 4'b1000;
															assign node6178 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node6181 = (inp[1]) ? 4'b1001 : node6182;
															assign node6182 = (inp[0]) ? 4'b1100 : 4'b1101;
													assign node6186 = (inp[4]) ? node6190 : node6187;
														assign node6187 = (inp[1]) ? 4'b1110 : 4'b1011;
														assign node6190 = (inp[1]) ? node6192 : 4'b1110;
															assign node6192 = (inp[0]) ? 4'b1010 : 4'b1011;
												assign node6195 = (inp[7]) ? node6207 : node6196;
													assign node6196 = (inp[1]) ? node6202 : node6197;
														assign node6197 = (inp[4]) ? 4'b1010 : node6198;
															assign node6198 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node6202 = (inp[4]) ? node6204 : 4'b1110;
															assign node6204 = (inp[0]) ? 4'b1010 : 4'b1011;
													assign node6207 = (inp[1]) ? node6215 : node6208;
														assign node6208 = (inp[4]) ? node6212 : node6209;
															assign node6209 = (inp[0]) ? 4'b1000 : 4'b1001;
															assign node6212 = (inp[0]) ? 4'b1101 : 4'b1100;
														assign node6215 = (inp[0]) ? 4'b1001 : node6216;
															assign node6216 = (inp[4]) ? 4'b1000 : 4'b1001;
											assign node6220 = (inp[15]) ? node6252 : node6221;
												assign node6221 = (inp[7]) ? node6237 : node6222;
													assign node6222 = (inp[0]) ? node6230 : node6223;
														assign node6223 = (inp[4]) ? node6227 : node6224;
															assign node6224 = (inp[1]) ? 4'b1000 : 4'b1100;
															assign node6227 = (inp[1]) ? 4'b1101 : 4'b1000;
														assign node6230 = (inp[4]) ? node6234 : node6231;
															assign node6231 = (inp[1]) ? 4'b1000 : 4'b1101;
															assign node6234 = (inp[1]) ? 4'b1101 : 4'b1000;
													assign node6237 = (inp[0]) ? node6245 : node6238;
														assign node6238 = (inp[1]) ? node6242 : node6239;
															assign node6239 = (inp[4]) ? 4'b1010 : 4'b1111;
															assign node6242 = (inp[4]) ? 4'b1111 : 4'b1010;
														assign node6245 = (inp[1]) ? node6249 : node6246;
															assign node6246 = (inp[4]) ? 4'b1011 : 4'b1111;
															assign node6249 = (inp[4]) ? 4'b1110 : 4'b1011;
												assign node6252 = (inp[7]) ? node6266 : node6253;
													assign node6253 = (inp[1]) ? node6259 : node6254;
														assign node6254 = (inp[0]) ? node6256 : 4'b1111;
															assign node6256 = (inp[10]) ? 4'b1111 : 4'b1110;
														assign node6259 = (inp[4]) ? node6263 : node6260;
															assign node6260 = (inp[0]) ? 4'b1010 : 4'b1011;
															assign node6263 = (inp[0]) ? 4'b1111 : 4'b1110;
													assign node6266 = (inp[1]) ? node6270 : node6267;
														assign node6267 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node6270 = (inp[0]) ? 4'b1100 : node6271;
															assign node6271 = (inp[4]) ? 4'b1101 : 4'b1100;
										assign node6275 = (inp[13]) ? node6337 : node6276;
											assign node6276 = (inp[0]) ? node6306 : node6277;
												assign node6277 = (inp[1]) ? node6293 : node6278;
													assign node6278 = (inp[4]) ? node6286 : node6279;
														assign node6279 = (inp[15]) ? node6283 : node6280;
															assign node6280 = (inp[7]) ? 4'b1110 : 4'b1100;
															assign node6283 = (inp[7]) ? 4'b1100 : 4'b1110;
														assign node6286 = (inp[7]) ? node6290 : node6287;
															assign node6287 = (inp[15]) ? 4'b1110 : 4'b1000;
															assign node6290 = (inp[15]) ? 4'b1000 : 4'b1010;
													assign node6293 = (inp[15]) ? node6301 : node6294;
														assign node6294 = (inp[7]) ? node6298 : node6295;
															assign node6295 = (inp[4]) ? 4'b1101 : 4'b1000;
															assign node6298 = (inp[4]) ? 4'b1111 : 4'b1011;
														assign node6301 = (inp[7]) ? 4'b1100 : node6302;
															assign node6302 = (inp[4]) ? 4'b1110 : 4'b1010;
												assign node6306 = (inp[1]) ? node6322 : node6307;
													assign node6307 = (inp[4]) ? node6315 : node6308;
														assign node6308 = (inp[7]) ? node6312 : node6309;
															assign node6309 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node6312 = (inp[15]) ? 4'b1101 : 4'b1110;
														assign node6315 = (inp[15]) ? node6319 : node6316;
															assign node6316 = (inp[7]) ? 4'b1010 : 4'b1001;
															assign node6319 = (inp[7]) ? 4'b1001 : 4'b1111;
													assign node6322 = (inp[4]) ? node6330 : node6323;
														assign node6323 = (inp[15]) ? node6327 : node6324;
															assign node6324 = (inp[7]) ? 4'b1010 : 4'b1000;
															assign node6327 = (inp[7]) ? 4'b1100 : 4'b1011;
														assign node6330 = (inp[7]) ? node6334 : node6331;
															assign node6331 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node6334 = (inp[15]) ? 4'b1100 : 4'b1111;
											assign node6337 = (inp[0]) ? node6367 : node6338;
												assign node6338 = (inp[1]) ? node6352 : node6339;
													assign node6339 = (inp[4]) ? node6345 : node6340;
														assign node6340 = (inp[7]) ? node6342 : 4'b1001;
															assign node6342 = (inp[15]) ? 4'b1000 : 4'b1010;
														assign node6345 = (inp[7]) ? node6349 : node6346;
															assign node6346 = (inp[15]) ? 4'b1010 : 4'b1100;
															assign node6349 = (inp[15]) ? 4'b1101 : 4'b1110;
													assign node6352 = (inp[4]) ? node6360 : node6353;
														assign node6353 = (inp[7]) ? node6357 : node6354;
															assign node6354 = (inp[15]) ? 4'b1111 : 4'b1100;
															assign node6357 = (inp[15]) ? 4'b1001 : 4'b1111;
														assign node6360 = (inp[7]) ? node6364 : node6361;
															assign node6361 = (inp[15]) ? 4'b1011 : 4'b1000;
															assign node6364 = (inp[15]) ? 4'b1001 : 4'b1011;
												assign node6367 = (inp[15]) ? node6383 : node6368;
													assign node6368 = (inp[7]) ? node6376 : node6369;
														assign node6369 = (inp[1]) ? node6373 : node6370;
															assign node6370 = (inp[4]) ? 4'b1101 : 4'b1001;
															assign node6373 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node6376 = (inp[4]) ? node6380 : node6377;
															assign node6377 = (inp[1]) ? 4'b1110 : 4'b1011;
															assign node6380 = (inp[1]) ? 4'b1010 : 4'b1110;
													assign node6383 = (inp[7]) ? node6389 : node6384;
														assign node6384 = (inp[1]) ? node6386 : 4'b1010;
															assign node6386 = (inp[4]) ? 4'b1010 : 4'b1110;
														assign node6389 = (inp[1]) ? 4'b1000 : node6390;
															assign node6390 = (inp[4]) ? 4'b1100 : 4'b1000;
							assign node6394 = (inp[12]) ? node6680 : node6395;
								assign node6395 = (inp[2]) ? node6513 : node6396;
									assign node6396 = (inp[5]) ? node6438 : node6397;
										assign node6397 = (inp[13]) ? node6417 : node6398;
											assign node6398 = (inp[15]) ? node6402 : node6399;
												assign node6399 = (inp[7]) ? 4'b1011 : 4'b1001;
												assign node6402 = (inp[7]) ? node6412 : node6403;
													assign node6403 = (inp[1]) ? node6405 : 4'b1011;
														assign node6405 = (inp[0]) ? node6409 : node6406;
															assign node6406 = (inp[4]) ? 4'b1111 : 4'b1011;
															assign node6409 = (inp[4]) ? 4'b1110 : 4'b1010;
													assign node6412 = (inp[1]) ? 4'b1000 : node6413;
														assign node6413 = (inp[4]) ? 4'b1001 : 4'b1101;
											assign node6417 = (inp[15]) ? node6421 : node6418;
												assign node6418 = (inp[7]) ? 4'b1111 : 4'b1101;
												assign node6421 = (inp[7]) ? node6429 : node6422;
													assign node6422 = (inp[1]) ? node6424 : 4'b1110;
														assign node6424 = (inp[4]) ? 4'b1011 : node6425;
															assign node6425 = (inp[0]) ? 4'b1111 : 4'b1110;
													assign node6429 = (inp[1]) ? 4'b1101 : node6430;
														assign node6430 = (inp[4]) ? node6434 : node6431;
															assign node6431 = (inp[0]) ? 4'b1001 : 4'b1000;
															assign node6434 = (inp[0]) ? 4'b1101 : 4'b1100;
										assign node6438 = (inp[13]) ? node6476 : node6439;
											assign node6439 = (inp[15]) ? node6451 : node6440;
												assign node6440 = (inp[7]) ? node6446 : node6441;
													assign node6441 = (inp[4]) ? node6443 : 4'b1101;
														assign node6443 = (inp[0]) ? 4'b1100 : 4'b1101;
													assign node6446 = (inp[0]) ? node6448 : 4'b1110;
														assign node6448 = (inp[4]) ? 4'b1111 : 4'b1110;
												assign node6451 = (inp[7]) ? node6465 : node6452;
													assign node6452 = (inp[1]) ? node6458 : node6453;
														assign node6453 = (inp[4]) ? node6455 : 4'b1111;
															assign node6455 = (inp[0]) ? 4'b1110 : 4'b1111;
														assign node6458 = (inp[4]) ? node6462 : node6459;
															assign node6459 = (inp[0]) ? 4'b1110 : 4'b1111;
															assign node6462 = (inp[0]) ? 4'b1011 : 4'b1010;
													assign node6465 = (inp[1]) ? node6471 : node6466;
														assign node6466 = (inp[4]) ? 4'b1101 : node6467;
															assign node6467 = (inp[0]) ? 4'b1001 : 4'b1000;
														assign node6471 = (inp[4]) ? node6473 : 4'b1101;
															assign node6473 = (inp[0]) ? 4'b1100 : 4'b1101;
											assign node6476 = (inp[15]) ? node6488 : node6477;
												assign node6477 = (inp[7]) ? node6483 : node6478;
													assign node6478 = (inp[0]) ? 4'b1000 : node6479;
														assign node6479 = (inp[4]) ? 4'b1000 : 4'b1001;
													assign node6483 = (inp[4]) ? 4'b1011 : node6484;
														assign node6484 = (inp[0]) ? 4'b1011 : 4'b1010;
												assign node6488 = (inp[7]) ? node6500 : node6489;
													assign node6489 = (inp[4]) ? node6495 : node6490;
														assign node6490 = (inp[1]) ? 4'b1011 : node6491;
															assign node6491 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node6495 = (inp[1]) ? node6497 : 4'b1011;
															assign node6497 = (inp[0]) ? 4'b1110 : 4'b1111;
													assign node6500 = (inp[4]) ? node6508 : node6501;
														assign node6501 = (inp[1]) ? node6505 : node6502;
															assign node6502 = (inp[0]) ? 4'b1100 : 4'b1101;
															assign node6505 = (inp[0]) ? 4'b1001 : 4'b1000;
														assign node6508 = (inp[0]) ? 4'b1001 : node6509;
															assign node6509 = (inp[1]) ? 4'b1001 : 4'b1000;
									assign node6513 = (inp[15]) ? node6589 : node6514;
										assign node6514 = (inp[7]) ? node6560 : node6515;
											assign node6515 = (inp[4]) ? node6545 : node6516;
												assign node6516 = (inp[0]) ? node6524 : node6517;
													assign node6517 = (inp[5]) ? node6521 : node6518;
														assign node6518 = (inp[13]) ? 4'b1101 : 4'b1001;
														assign node6521 = (inp[13]) ? 4'b1000 : 4'b1101;
													assign node6524 = (inp[10]) ? node6538 : node6525;
														assign node6525 = (inp[1]) ? node6533 : node6526;
															assign node6526 = (inp[13]) ? node6530 : node6527;
																assign node6527 = (inp[5]) ? 4'b1100 : 4'b1000;
																assign node6530 = (inp[5]) ? 4'b1000 : 4'b1100;
															assign node6533 = (inp[5]) ? 4'b1100 : node6534;
																assign node6534 = (inp[13]) ? 4'b1100 : 4'b1000;
														assign node6538 = (inp[13]) ? node6542 : node6539;
															assign node6539 = (inp[5]) ? 4'b1100 : 4'b1000;
															assign node6542 = (inp[5]) ? 4'b1000 : 4'b1100;
												assign node6545 = (inp[0]) ? node6553 : node6546;
													assign node6546 = (inp[5]) ? node6550 : node6547;
														assign node6547 = (inp[13]) ? 4'b1100 : 4'b1000;
														assign node6550 = (inp[13]) ? 4'b1001 : 4'b1101;
													assign node6553 = (inp[5]) ? node6557 : node6554;
														assign node6554 = (inp[13]) ? 4'b1101 : 4'b1001;
														assign node6557 = (inp[13]) ? 4'b1000 : 4'b1101;
											assign node6560 = (inp[0]) ? node6576 : node6561;
												assign node6561 = (inp[4]) ? node6569 : node6562;
													assign node6562 = (inp[5]) ? node6566 : node6563;
														assign node6563 = (inp[13]) ? 4'b1111 : 4'b1011;
														assign node6566 = (inp[13]) ? 4'b1011 : 4'b1110;
													assign node6569 = (inp[5]) ? node6573 : node6570;
														assign node6570 = (inp[13]) ? 4'b1110 : 4'b1010;
														assign node6573 = (inp[13]) ? 4'b1010 : 4'b1110;
												assign node6576 = (inp[13]) ? node6584 : node6577;
													assign node6577 = (inp[5]) ? node6581 : node6578;
														assign node6578 = (inp[4]) ? 4'b1011 : 4'b1010;
														assign node6581 = (inp[4]) ? 4'b1110 : 4'b1111;
													assign node6584 = (inp[5]) ? 4'b1011 : node6585;
														assign node6585 = (inp[4]) ? 4'b1111 : 4'b1110;
										assign node6589 = (inp[7]) ? node6633 : node6590;
											assign node6590 = (inp[13]) ? node6612 : node6591;
												assign node6591 = (inp[5]) ? node6603 : node6592;
													assign node6592 = (inp[4]) ? node6598 : node6593;
														assign node6593 = (inp[1]) ? 4'b1010 : node6594;
															assign node6594 = (inp[0]) ? 4'b1010 : 4'b1011;
														assign node6598 = (inp[1]) ? 4'b1111 : node6599;
															assign node6599 = (inp[0]) ? 4'b1011 : 4'b1010;
													assign node6603 = (inp[1]) ? node6609 : node6604;
														assign node6604 = (inp[0]) ? node6606 : 4'b1111;
															assign node6606 = (inp[4]) ? 4'b1111 : 4'b1110;
														assign node6609 = (inp[4]) ? 4'b1010 : 4'b1110;
												assign node6612 = (inp[5]) ? node6626 : node6613;
													assign node6613 = (inp[4]) ? node6619 : node6614;
														assign node6614 = (inp[0]) ? 4'b1111 : node6615;
															assign node6615 = (inp[1]) ? 4'b1111 : 4'b1110;
														assign node6619 = (inp[1]) ? node6623 : node6620;
															assign node6620 = (inp[0]) ? 4'b1110 : 4'b1111;
															assign node6623 = (inp[0]) ? 4'b1011 : 4'b1010;
													assign node6626 = (inp[1]) ? node6628 : 4'b1011;
														assign node6628 = (inp[4]) ? 4'b1111 : node6629;
															assign node6629 = (inp[10]) ? 4'b1011 : 4'b1010;
											assign node6633 = (inp[13]) ? node6659 : node6634;
												assign node6634 = (inp[5]) ? node6648 : node6635;
													assign node6635 = (inp[1]) ? node6641 : node6636;
														assign node6636 = (inp[4]) ? 4'b1001 : node6637;
															assign node6637 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node6641 = (inp[4]) ? node6645 : node6642;
															assign node6642 = (inp[0]) ? 4'b1001 : 4'b1000;
															assign node6645 = (inp[0]) ? 4'b1000 : 4'b1001;
													assign node6648 = (inp[4]) ? node6654 : node6649;
														assign node6649 = (inp[1]) ? node6651 : 4'b1001;
															assign node6651 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node6654 = (inp[1]) ? 4'b1101 : node6655;
															assign node6655 = (inp[0]) ? 4'b1101 : 4'b1100;
												assign node6659 = (inp[5]) ? node6671 : node6660;
													assign node6660 = (inp[4]) ? node6666 : node6661;
														assign node6661 = (inp[1]) ? node6663 : 4'b1001;
															assign node6663 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node6666 = (inp[0]) ? node6668 : 4'b1100;
															assign node6668 = (inp[1]) ? 4'b1101 : 4'b1100;
													assign node6671 = (inp[1]) ? node6675 : node6672;
														assign node6672 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node6675 = (inp[4]) ? node6677 : 4'b1001;
															assign node6677 = (inp[0]) ? 4'b1001 : 4'b1000;
								assign node6680 = (inp[2]) ? node6906 : node6681;
									assign node6681 = (inp[15]) ? node6819 : node6682;
										assign node6682 = (inp[7]) ? node6768 : node6683;
											assign node6683 = (inp[0]) ? node6723 : node6684;
												assign node6684 = (inp[1]) ? node6700 : node6685;
													assign node6685 = (inp[5]) ? node6693 : node6686;
														assign node6686 = (inp[4]) ? node6690 : node6687;
															assign node6687 = (inp[13]) ? 4'b1101 : 4'b1001;
															assign node6690 = (inp[13]) ? 4'b1001 : 4'b1101;
														assign node6693 = (inp[4]) ? node6697 : node6694;
															assign node6694 = (inp[13]) ? 4'b1001 : 4'b1101;
															assign node6697 = (inp[13]) ? 4'b1100 : 4'b1000;
													assign node6700 = (inp[5]) ? node6716 : node6701;
														assign node6701 = (inp[10]) ? node6709 : node6702;
															assign node6702 = (inp[13]) ? node6706 : node6703;
																assign node6703 = (inp[4]) ? 4'b1000 : 4'b1100;
																assign node6706 = (inp[4]) ? 4'b1100 : 4'b1000;
															assign node6709 = (inp[4]) ? node6713 : node6710;
																assign node6710 = (inp[13]) ? 4'b1000 : 4'b1100;
																assign node6713 = (inp[13]) ? 4'b1100 : 4'b1000;
														assign node6716 = (inp[4]) ? node6720 : node6717;
															assign node6717 = (inp[13]) ? 4'b1100 : 4'b1000;
															assign node6720 = (inp[13]) ? 4'b1001 : 4'b1101;
												assign node6723 = (inp[1]) ? node6739 : node6724;
													assign node6724 = (inp[5]) ? node6732 : node6725;
														assign node6725 = (inp[13]) ? node6729 : node6726;
															assign node6726 = (inp[4]) ? 4'b1101 : 4'b1001;
															assign node6729 = (inp[4]) ? 4'b1000 : 4'b1101;
														assign node6732 = (inp[13]) ? node6736 : node6733;
															assign node6733 = (inp[4]) ? 4'b1000 : 4'b1101;
															assign node6736 = (inp[4]) ? 4'b1100 : 4'b1000;
													assign node6739 = (inp[10]) ? node6753 : node6740;
														assign node6740 = (inp[4]) ? node6748 : node6741;
															assign node6741 = (inp[5]) ? node6745 : node6742;
																assign node6742 = (inp[13]) ? 4'b1001 : 4'b1100;
																assign node6745 = (inp[13]) ? 4'b1101 : 4'b1001;
															assign node6748 = (inp[13]) ? 4'b1101 : node6749;
																assign node6749 = (inp[5]) ? 4'b1101 : 4'b1001;
														assign node6753 = (inp[13]) ? node6761 : node6754;
															assign node6754 = (inp[5]) ? node6758 : node6755;
																assign node6755 = (inp[4]) ? 4'b1001 : 4'b1100;
																assign node6758 = (inp[4]) ? 4'b1101 : 4'b1001;
															assign node6761 = (inp[4]) ? node6765 : node6762;
																assign node6762 = (inp[5]) ? 4'b1101 : 4'b1001;
																assign node6765 = (inp[5]) ? 4'b1000 : 4'b1101;
											assign node6768 = (inp[5]) ? node6794 : node6769;
												assign node6769 = (inp[1]) ? node6785 : node6770;
													assign node6770 = (inp[0]) ? node6778 : node6771;
														assign node6771 = (inp[4]) ? node6775 : node6772;
															assign node6772 = (inp[13]) ? 4'b1111 : 4'b1011;
															assign node6775 = (inp[13]) ? 4'b1010 : 4'b1111;
														assign node6778 = (inp[4]) ? node6782 : node6779;
															assign node6779 = (inp[13]) ? 4'b1110 : 4'b1010;
															assign node6782 = (inp[13]) ? 4'b1010 : 4'b1110;
													assign node6785 = (inp[4]) ? node6791 : node6786;
														assign node6786 = (inp[13]) ? 4'b1011 : node6787;
															assign node6787 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node6791 = (inp[13]) ? 4'b1111 : 4'b1011;
												assign node6794 = (inp[1]) ? node6810 : node6795;
													assign node6795 = (inp[0]) ? node6803 : node6796;
														assign node6796 = (inp[4]) ? node6800 : node6797;
															assign node6797 = (inp[13]) ? 4'b1011 : 4'b1110;
															assign node6800 = (inp[13]) ? 4'b1111 : 4'b1011;
														assign node6803 = (inp[4]) ? node6807 : node6804;
															assign node6804 = (inp[13]) ? 4'b1011 : 4'b1111;
															assign node6807 = (inp[13]) ? 4'b1110 : 4'b1010;
													assign node6810 = (inp[4]) ? node6814 : node6811;
														assign node6811 = (inp[13]) ? 4'b1110 : 4'b1010;
														assign node6814 = (inp[0]) ? node6816 : 4'b1110;
															assign node6816 = (inp[13]) ? 4'b1011 : 4'b1111;
										assign node6819 = (inp[7]) ? node6863 : node6820;
											assign node6820 = (inp[13]) ? node6842 : node6821;
												assign node6821 = (inp[5]) ? node6833 : node6822;
													assign node6822 = (inp[4]) ? node6828 : node6823;
														assign node6823 = (inp[1]) ? node6825 : 4'b1011;
															assign node6825 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node6828 = (inp[1]) ? 4'b1011 : node6829;
															assign node6829 = (inp[0]) ? 4'b1010 : 4'b1011;
													assign node6833 = (inp[4]) ? node6837 : node6834;
														assign node6834 = (inp[1]) ? 4'b1011 : 4'b1111;
														assign node6837 = (inp[1]) ? node6839 : 4'b1110;
															assign node6839 = (inp[0]) ? 4'b1110 : 4'b1111;
												assign node6842 = (inp[5]) ? node6852 : node6843;
													assign node6843 = (inp[1]) ? node6849 : node6844;
														assign node6844 = (inp[0]) ? node6846 : 4'b1110;
															assign node6846 = (inp[4]) ? 4'b1111 : 4'b1110;
														assign node6849 = (inp[4]) ? 4'b1110 : 4'b1010;
													assign node6852 = (inp[4]) ? node6858 : node6853;
														assign node6853 = (inp[1]) ? 4'b1110 : node6854;
															assign node6854 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node6858 = (inp[1]) ? 4'b1011 : node6859;
															assign node6859 = (inp[0]) ? 4'b1010 : 4'b1011;
											assign node6863 = (inp[13]) ? node6885 : node6864;
												assign node6864 = (inp[5]) ? node6874 : node6865;
													assign node6865 = (inp[4]) ? node6871 : node6866;
														assign node6866 = (inp[0]) ? 4'b1000 : node6867;
															assign node6867 = (inp[1]) ? 4'b1001 : 4'b1000;
														assign node6871 = (inp[1]) ? 4'b1000 : 4'b1100;
													assign node6874 = (inp[4]) ? node6880 : node6875;
														assign node6875 = (inp[1]) ? node6877 : 4'b1101;
															assign node6877 = (inp[0]) ? 4'b1101 : 4'b1100;
														assign node6880 = (inp[1]) ? node6882 : 4'b1000;
															assign node6882 = (inp[0]) ? 4'b1100 : 4'b1101;
												assign node6885 = (inp[5]) ? node6897 : node6886;
													assign node6886 = (inp[4]) ? node6892 : node6887;
														assign node6887 = (inp[0]) ? 4'b1101 : node6888;
															assign node6888 = (inp[1]) ? 4'b1100 : 4'b1101;
														assign node6892 = (inp[1]) ? 4'b1101 : node6893;
															assign node6893 = (inp[0]) ? 4'b1000 : 4'b1001;
													assign node6897 = (inp[4]) ? node6903 : node6898;
														assign node6898 = (inp[1]) ? 4'b1000 : node6899;
															assign node6899 = (inp[0]) ? 4'b1001 : 4'b1000;
														assign node6903 = (inp[1]) ? 4'b1001 : 4'b1101;
									assign node6906 = (inp[5]) ? node7014 : node6907;
										assign node6907 = (inp[13]) ? node6965 : node6908;
											assign node6908 = (inp[15]) ? node6940 : node6909;
												assign node6909 = (inp[7]) ? node6923 : node6910;
													assign node6910 = (inp[4]) ? node6918 : node6911;
														assign node6911 = (inp[1]) ? node6915 : node6912;
															assign node6912 = (inp[0]) ? 4'b1000 : 4'b1001;
															assign node6915 = (inp[0]) ? 4'b1101 : 4'b1100;
														assign node6918 = (inp[1]) ? 4'b1000 : node6919;
															assign node6919 = (inp[0]) ? 4'b1101 : 4'b1100;
													assign node6923 = (inp[0]) ? node6933 : node6924;
														assign node6924 = (inp[10]) ? node6926 : 4'b1111;
															assign node6926 = (inp[1]) ? node6930 : node6927;
																assign node6927 = (inp[4]) ? 4'b1111 : 4'b1010;
																assign node6930 = (inp[4]) ? 4'b1010 : 4'b1111;
														assign node6933 = (inp[4]) ? node6937 : node6934;
															assign node6934 = (inp[1]) ? 4'b1111 : 4'b1010;
															assign node6937 = (inp[1]) ? 4'b1011 : 4'b1111;
												assign node6940 = (inp[7]) ? node6952 : node6941;
													assign node6941 = (inp[4]) ? node6947 : node6942;
														assign node6942 = (inp[1]) ? 4'b1111 : node6943;
															assign node6943 = (inp[0]) ? 4'b1010 : 4'b1011;
														assign node6947 = (inp[1]) ? node6949 : 4'b1011;
															assign node6949 = (inp[0]) ? 4'b1011 : 4'b1010;
													assign node6952 = (inp[1]) ? node6960 : node6953;
														assign node6953 = (inp[4]) ? node6957 : node6954;
															assign node6954 = (inp[0]) ? 4'b1001 : 4'b1000;
															assign node6957 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node6960 = (inp[0]) ? 4'b1000 : node6961;
															assign node6961 = (inp[4]) ? 4'b1001 : 4'b1000;
											assign node6965 = (inp[15]) ? node6989 : node6966;
												assign node6966 = (inp[7]) ? node6976 : node6967;
													assign node6967 = (inp[4]) ? node6973 : node6968;
														assign node6968 = (inp[1]) ? 4'b1001 : node6969;
															assign node6969 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node6973 = (inp[1]) ? 4'b1100 : 4'b1001;
													assign node6976 = (inp[4]) ? node6982 : node6977;
														assign node6977 = (inp[1]) ? node6979 : 4'b1110;
															assign node6979 = (inp[0]) ? 4'b1010 : 4'b1011;
														assign node6982 = (inp[1]) ? node6986 : node6983;
															assign node6983 = (inp[0]) ? 4'b1010 : 4'b1011;
															assign node6986 = (inp[0]) ? 4'b1111 : 4'b1110;
												assign node6989 = (inp[7]) ? node7003 : node6990;
													assign node6990 = (inp[4]) ? node6998 : node6991;
														assign node6991 = (inp[1]) ? node6995 : node6992;
															assign node6992 = (inp[0]) ? 4'b1111 : 4'b1110;
															assign node6995 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node6998 = (inp[1]) ? node7000 : 4'b1110;
															assign node7000 = (inp[0]) ? 4'b1110 : 4'b1111;
													assign node7003 = (inp[1]) ? node7009 : node7004;
														assign node7004 = (inp[4]) ? 4'b1001 : node7005;
															assign node7005 = (inp[10]) ? 4'b1100 : 4'b1101;
														assign node7009 = (inp[4]) ? node7011 : 4'b1101;
															assign node7011 = (inp[0]) ? 4'b1101 : 4'b1100;
										assign node7014 = (inp[13]) ? node7076 : node7015;
											assign node7015 = (inp[0]) ? node7045 : node7016;
												assign node7016 = (inp[1]) ? node7032 : node7017;
													assign node7017 = (inp[4]) ? node7025 : node7018;
														assign node7018 = (inp[7]) ? node7022 : node7019;
															assign node7019 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node7022 = (inp[15]) ? 4'b1101 : 4'b1111;
														assign node7025 = (inp[7]) ? node7029 : node7026;
															assign node7026 = (inp[15]) ? 4'b1111 : 4'b1001;
															assign node7029 = (inp[15]) ? 4'b1001 : 4'b1011;
													assign node7032 = (inp[15]) ? node7040 : node7033;
														assign node7033 = (inp[7]) ? node7037 : node7034;
															assign node7034 = (inp[4]) ? 4'b1100 : 4'b1001;
															assign node7037 = (inp[4]) ? 4'b1110 : 4'b1010;
														assign node7040 = (inp[7]) ? 4'b1101 : node7041;
															assign node7041 = (inp[4]) ? 4'b1111 : 4'b1011;
												assign node7045 = (inp[1]) ? node7061 : node7046;
													assign node7046 = (inp[4]) ? node7054 : node7047;
														assign node7047 = (inp[7]) ? node7051 : node7048;
															assign node7048 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node7051 = (inp[15]) ? 4'b1100 : 4'b1111;
														assign node7054 = (inp[7]) ? node7058 : node7055;
															assign node7055 = (inp[15]) ? 4'b1110 : 4'b1000;
															assign node7058 = (inp[15]) ? 4'b1000 : 4'b1011;
													assign node7061 = (inp[4]) ? node7069 : node7062;
														assign node7062 = (inp[7]) ? node7066 : node7063;
															assign node7063 = (inp[15]) ? 4'b1010 : 4'b1001;
															assign node7066 = (inp[15]) ? 4'b1101 : 4'b1011;
														assign node7069 = (inp[15]) ? node7073 : node7070;
															assign node7070 = (inp[7]) ? 4'b1110 : 4'b1101;
															assign node7073 = (inp[7]) ? 4'b1101 : 4'b1111;
											assign node7076 = (inp[0]) ? node7106 : node7077;
												assign node7077 = (inp[1]) ? node7091 : node7078;
													assign node7078 = (inp[4]) ? node7084 : node7079;
														assign node7079 = (inp[15]) ? 4'b1011 : node7080;
															assign node7080 = (inp[7]) ? 4'b1011 : 4'b1000;
														assign node7084 = (inp[15]) ? node7088 : node7085;
															assign node7085 = (inp[7]) ? 4'b1111 : 4'b1101;
															assign node7088 = (inp[7]) ? 4'b1100 : 4'b1011;
													assign node7091 = (inp[4]) ? node7099 : node7092;
														assign node7092 = (inp[15]) ? node7096 : node7093;
															assign node7093 = (inp[7]) ? 4'b1110 : 4'b1101;
															assign node7096 = (inp[7]) ? 4'b1000 : 4'b1110;
														assign node7099 = (inp[7]) ? node7103 : node7100;
															assign node7100 = (inp[15]) ? 4'b1010 : 4'b1001;
															assign node7103 = (inp[15]) ? 4'b1000 : 4'b1010;
												assign node7106 = (inp[15]) ? node7122 : node7107;
													assign node7107 = (inp[7]) ? node7115 : node7108;
														assign node7108 = (inp[1]) ? node7112 : node7109;
															assign node7109 = (inp[4]) ? 4'b1100 : 4'b1000;
															assign node7112 = (inp[4]) ? 4'b1001 : 4'b1101;
														assign node7115 = (inp[1]) ? node7119 : node7116;
															assign node7116 = (inp[4]) ? 4'b1111 : 4'b1010;
															assign node7119 = (inp[4]) ? 4'b1011 : 4'b1111;
													assign node7122 = (inp[7]) ? node7128 : node7123;
														assign node7123 = (inp[4]) ? 4'b1011 : node7124;
															assign node7124 = (inp[1]) ? 4'b1111 : 4'b1011;
														assign node7128 = (inp[1]) ? 4'b1001 : node7129;
															assign node7129 = (inp[4]) ? 4'b1101 : 4'b1001;
						assign node7133 = (inp[9]) ? node7819 : node7134;
							assign node7134 = (inp[12]) ? node7436 : node7135;
								assign node7135 = (inp[2]) ? node7255 : node7136;
									assign node7136 = (inp[5]) ? node7180 : node7137;
										assign node7137 = (inp[13]) ? node7159 : node7138;
											assign node7138 = (inp[15]) ? node7142 : node7139;
												assign node7139 = (inp[7]) ? 4'b1011 : 4'b1001;
												assign node7142 = (inp[7]) ? node7152 : node7143;
													assign node7143 = (inp[1]) ? node7145 : 4'b1011;
														assign node7145 = (inp[0]) ? node7149 : node7146;
															assign node7146 = (inp[4]) ? 4'b1111 : 4'b1011;
															assign node7149 = (inp[4]) ? 4'b1110 : 4'b1010;
													assign node7152 = (inp[1]) ? 4'b1000 : node7153;
														assign node7153 = (inp[4]) ? node7155 : 4'b1101;
															assign node7155 = (inp[0]) ? 4'b1000 : 4'b1001;
											assign node7159 = (inp[15]) ? node7163 : node7160;
												assign node7160 = (inp[7]) ? 4'b1111 : 4'b1101;
												assign node7163 = (inp[7]) ? node7171 : node7164;
													assign node7164 = (inp[1]) ? node7166 : 4'b1110;
														assign node7166 = (inp[4]) ? 4'b1011 : node7167;
															assign node7167 = (inp[0]) ? 4'b1111 : 4'b1110;
													assign node7171 = (inp[1]) ? 4'b1101 : node7172;
														assign node7172 = (inp[0]) ? node7176 : node7173;
															assign node7173 = (inp[4]) ? 4'b1100 : 4'b1000;
															assign node7176 = (inp[4]) ? 4'b1101 : 4'b1001;
										assign node7180 = (inp[13]) ? node7218 : node7181;
											assign node7181 = (inp[15]) ? node7193 : node7182;
												assign node7182 = (inp[7]) ? node7188 : node7183;
													assign node7183 = (inp[4]) ? node7185 : 4'b1101;
														assign node7185 = (inp[0]) ? 4'b1100 : 4'b1101;
													assign node7188 = (inp[4]) ? node7190 : 4'b1110;
														assign node7190 = (inp[0]) ? 4'b1111 : 4'b1110;
												assign node7193 = (inp[7]) ? node7207 : node7194;
													assign node7194 = (inp[4]) ? node7200 : node7195;
														assign node7195 = (inp[1]) ? node7197 : 4'b1111;
															assign node7197 = (inp[0]) ? 4'b1110 : 4'b1111;
														assign node7200 = (inp[1]) ? node7204 : node7201;
															assign node7201 = (inp[0]) ? 4'b1110 : 4'b1111;
															assign node7204 = (inp[0]) ? 4'b1011 : 4'b1010;
													assign node7207 = (inp[4]) ? node7213 : node7208;
														assign node7208 = (inp[1]) ? 4'b1101 : node7209;
															assign node7209 = (inp[0]) ? 4'b1001 : 4'b1000;
														assign node7213 = (inp[0]) ? node7215 : 4'b1101;
															assign node7215 = (inp[1]) ? 4'b1100 : 4'b1101;
											assign node7218 = (inp[15]) ? node7230 : node7219;
												assign node7219 = (inp[7]) ? node7225 : node7220;
													assign node7220 = (inp[4]) ? 4'b1000 : node7221;
														assign node7221 = (inp[0]) ? 4'b1000 : 4'b1001;
													assign node7225 = (inp[4]) ? 4'b1011 : node7226;
														assign node7226 = (inp[0]) ? 4'b1011 : 4'b1010;
												assign node7230 = (inp[7]) ? node7242 : node7231;
													assign node7231 = (inp[4]) ? node7237 : node7232;
														assign node7232 = (inp[1]) ? 4'b1011 : node7233;
															assign node7233 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node7237 = (inp[1]) ? node7239 : 4'b1011;
															assign node7239 = (inp[0]) ? 4'b1110 : 4'b1111;
													assign node7242 = (inp[4]) ? node7250 : node7243;
														assign node7243 = (inp[1]) ? node7247 : node7244;
															assign node7244 = (inp[0]) ? 4'b1100 : 4'b1101;
															assign node7247 = (inp[0]) ? 4'b1001 : 4'b1000;
														assign node7250 = (inp[0]) ? 4'b1001 : node7251;
															assign node7251 = (inp[1]) ? 4'b1001 : 4'b1000;
									assign node7255 = (inp[15]) ? node7345 : node7256;
										assign node7256 = (inp[7]) ? node7314 : node7257;
											assign node7257 = (inp[13]) ? node7285 : node7258;
												assign node7258 = (inp[5]) ? node7280 : node7259;
													assign node7259 = (inp[10]) ? node7267 : node7260;
														assign node7260 = (inp[0]) ? node7264 : node7261;
															assign node7261 = (inp[4]) ? 4'b1000 : 4'b1001;
															assign node7264 = (inp[4]) ? 4'b1001 : 4'b1000;
														assign node7267 = (inp[1]) ? node7275 : node7268;
															assign node7268 = (inp[0]) ? node7272 : node7269;
																assign node7269 = (inp[4]) ? 4'b1000 : 4'b1001;
																assign node7272 = (inp[4]) ? 4'b1001 : 4'b1000;
															assign node7275 = (inp[0]) ? node7277 : 4'b1001;
																assign node7277 = (inp[4]) ? 4'b1001 : 4'b1000;
													assign node7280 = (inp[0]) ? node7282 : 4'b1101;
														assign node7282 = (inp[4]) ? 4'b1101 : 4'b1100;
												assign node7285 = (inp[5]) ? node7309 : node7286;
													assign node7286 = (inp[1]) ? node7294 : node7287;
														assign node7287 = (inp[0]) ? node7291 : node7288;
															assign node7288 = (inp[4]) ? 4'b1100 : 4'b1101;
															assign node7291 = (inp[4]) ? 4'b1101 : 4'b1100;
														assign node7294 = (inp[10]) ? node7302 : node7295;
															assign node7295 = (inp[0]) ? node7299 : node7296;
																assign node7296 = (inp[4]) ? 4'b1100 : 4'b1101;
																assign node7299 = (inp[4]) ? 4'b1101 : 4'b1100;
															assign node7302 = (inp[0]) ? node7306 : node7303;
																assign node7303 = (inp[4]) ? 4'b1100 : 4'b1101;
																assign node7306 = (inp[4]) ? 4'b1101 : 4'b1100;
													assign node7309 = (inp[4]) ? node7311 : 4'b1000;
														assign node7311 = (inp[0]) ? 4'b1000 : 4'b1001;
											assign node7314 = (inp[4]) ? node7330 : node7315;
												assign node7315 = (inp[0]) ? node7323 : node7316;
													assign node7316 = (inp[13]) ? node7320 : node7317;
														assign node7317 = (inp[5]) ? 4'b1110 : 4'b1011;
														assign node7320 = (inp[5]) ? 4'b1011 : 4'b1111;
													assign node7323 = (inp[5]) ? node7327 : node7324;
														assign node7324 = (inp[13]) ? 4'b1110 : 4'b1010;
														assign node7327 = (inp[13]) ? 4'b1011 : 4'b1111;
												assign node7330 = (inp[0]) ? node7338 : node7331;
													assign node7331 = (inp[13]) ? node7335 : node7332;
														assign node7332 = (inp[5]) ? 4'b1110 : 4'b1010;
														assign node7335 = (inp[5]) ? 4'b1010 : 4'b1110;
													assign node7338 = (inp[5]) ? node7342 : node7339;
														assign node7339 = (inp[13]) ? 4'b1111 : 4'b1011;
														assign node7342 = (inp[13]) ? 4'b1011 : 4'b1110;
										assign node7345 = (inp[7]) ? node7391 : node7346;
											assign node7346 = (inp[13]) ? node7368 : node7347;
												assign node7347 = (inp[5]) ? node7359 : node7348;
													assign node7348 = (inp[4]) ? node7354 : node7349;
														assign node7349 = (inp[1]) ? 4'b1010 : node7350;
															assign node7350 = (inp[0]) ? 4'b1010 : 4'b1011;
														assign node7354 = (inp[1]) ? 4'b1111 : node7355;
															assign node7355 = (inp[0]) ? 4'b1011 : 4'b1010;
													assign node7359 = (inp[1]) ? node7365 : node7360;
														assign node7360 = (inp[4]) ? 4'b1111 : node7361;
															assign node7361 = (inp[10]) ? 4'b1110 : 4'b1111;
														assign node7365 = (inp[4]) ? 4'b1010 : 4'b1110;
												assign node7368 = (inp[5]) ? node7380 : node7369;
													assign node7369 = (inp[4]) ? node7375 : node7370;
														assign node7370 = (inp[1]) ? 4'b1111 : node7371;
															assign node7371 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node7375 = (inp[1]) ? node7377 : 4'b1111;
															assign node7377 = (inp[0]) ? 4'b1011 : 4'b1010;
													assign node7380 = (inp[4]) ? node7386 : node7381;
														assign node7381 = (inp[0]) ? node7383 : 4'b1011;
															assign node7383 = (inp[1]) ? 4'b1010 : 4'b1011;
														assign node7386 = (inp[1]) ? 4'b1111 : node7387;
															assign node7387 = (inp[0]) ? 4'b1011 : 4'b1010;
											assign node7391 = (inp[13]) ? node7417 : node7392;
												assign node7392 = (inp[5]) ? node7406 : node7393;
													assign node7393 = (inp[4]) ? node7401 : node7394;
														assign node7394 = (inp[1]) ? node7398 : node7395;
															assign node7395 = (inp[0]) ? 4'b1100 : 4'b1101;
															assign node7398 = (inp[0]) ? 4'b1001 : 4'b1000;
														assign node7401 = (inp[1]) ? node7403 : 4'b1001;
															assign node7403 = (inp[0]) ? 4'b1000 : 4'b1001;
													assign node7406 = (inp[1]) ? node7412 : node7407;
														assign node7407 = (inp[4]) ? node7409 : 4'b1001;
															assign node7409 = (inp[0]) ? 4'b1101 : 4'b1100;
														assign node7412 = (inp[0]) ? node7414 : 4'b1101;
															assign node7414 = (inp[4]) ? 4'b1101 : 4'b1100;
												assign node7417 = (inp[5]) ? node7427 : node7418;
													assign node7418 = (inp[4]) ? node7422 : node7419;
														assign node7419 = (inp[1]) ? 4'b1100 : 4'b1001;
														assign node7422 = (inp[1]) ? node7424 : 4'b1100;
															assign node7424 = (inp[0]) ? 4'b1101 : 4'b1100;
													assign node7427 = (inp[1]) ? node7431 : node7428;
														assign node7428 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node7431 = (inp[0]) ? 4'b1001 : node7432;
															assign node7432 = (inp[4]) ? 4'b1000 : 4'b1001;
								assign node7436 = (inp[5]) ? node7634 : node7437;
									assign node7437 = (inp[13]) ? node7539 : node7438;
										assign node7438 = (inp[15]) ? node7486 : node7439;
											assign node7439 = (inp[7]) ? node7463 : node7440;
												assign node7440 = (inp[1]) ? node7452 : node7441;
													assign node7441 = (inp[4]) ? node7447 : node7442;
														assign node7442 = (inp[2]) ? node7444 : 4'b1001;
															assign node7444 = (inp[0]) ? 4'b1000 : 4'b1001;
														assign node7447 = (inp[2]) ? node7449 : 4'b1101;
															assign node7449 = (inp[0]) ? 4'b1101 : 4'b1100;
													assign node7452 = (inp[4]) ? node7458 : node7453;
														assign node7453 = (inp[2]) ? node7455 : 4'b1100;
															assign node7455 = (inp[0]) ? 4'b1101 : 4'b1100;
														assign node7458 = (inp[0]) ? node7460 : 4'b1000;
															assign node7460 = (inp[2]) ? 4'b1000 : 4'b1001;
												assign node7463 = (inp[1]) ? node7475 : node7464;
													assign node7464 = (inp[4]) ? node7470 : node7465;
														assign node7465 = (inp[0]) ? 4'b1010 : node7466;
															assign node7466 = (inp[10]) ? 4'b1010 : 4'b1011;
														assign node7470 = (inp[0]) ? node7472 : 4'b1111;
															assign node7472 = (inp[2]) ? 4'b1111 : 4'b1110;
													assign node7475 = (inp[4]) ? node7481 : node7476;
														assign node7476 = (inp[0]) ? 4'b1111 : node7477;
															assign node7477 = (inp[2]) ? 4'b1111 : 4'b1110;
														assign node7481 = (inp[2]) ? node7483 : 4'b1011;
															assign node7483 = (inp[0]) ? 4'b1011 : 4'b1010;
											assign node7486 = (inp[7]) ? node7516 : node7487;
												assign node7487 = (inp[1]) ? node7505 : node7488;
													assign node7488 = (inp[0]) ? node7490 : 4'b1011;
														assign node7490 = (inp[10]) ? node7498 : node7491;
															assign node7491 = (inp[4]) ? node7495 : node7492;
																assign node7492 = (inp[2]) ? 4'b1010 : 4'b1011;
																assign node7495 = (inp[2]) ? 4'b1011 : 4'b1010;
															assign node7498 = (inp[4]) ? node7502 : node7499;
																assign node7499 = (inp[2]) ? 4'b1010 : 4'b1011;
																assign node7502 = (inp[2]) ? 4'b1011 : 4'b1010;
													assign node7505 = (inp[4]) ? node7511 : node7506;
														assign node7506 = (inp[2]) ? 4'b1111 : node7507;
															assign node7507 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node7511 = (inp[0]) ? 4'b1011 : node7512;
															assign node7512 = (inp[2]) ? 4'b1010 : 4'b1011;
												assign node7516 = (inp[4]) ? node7528 : node7517;
													assign node7517 = (inp[1]) ? node7523 : node7518;
														assign node7518 = (inp[2]) ? node7520 : 4'b1000;
															assign node7520 = (inp[0]) ? 4'b1001 : 4'b1000;
														assign node7523 = (inp[2]) ? 4'b1000 : node7524;
															assign node7524 = (inp[0]) ? 4'b1000 : 4'b1001;
													assign node7528 = (inp[1]) ? node7534 : node7529;
														assign node7529 = (inp[0]) ? 4'b1100 : node7530;
															assign node7530 = (inp[2]) ? 4'b1101 : 4'b1100;
														assign node7534 = (inp[0]) ? 4'b1000 : node7535;
															assign node7535 = (inp[2]) ? 4'b1001 : 4'b1000;
										assign node7539 = (inp[15]) ? node7587 : node7540;
											assign node7540 = (inp[7]) ? node7564 : node7541;
												assign node7541 = (inp[1]) ? node7553 : node7542;
													assign node7542 = (inp[4]) ? node7548 : node7543;
														assign node7543 = (inp[0]) ? node7545 : 4'b1101;
															assign node7545 = (inp[2]) ? 4'b1100 : 4'b1101;
														assign node7548 = (inp[0]) ? node7550 : 4'b1001;
															assign node7550 = (inp[2]) ? 4'b1001 : 4'b1000;
													assign node7553 = (inp[4]) ? node7559 : node7554;
														assign node7554 = (inp[2]) ? 4'b1001 : node7555;
															assign node7555 = (inp[0]) ? 4'b1001 : 4'b1000;
														assign node7559 = (inp[10]) ? 4'b1100 : node7560;
															assign node7560 = (inp[2]) ? 4'b1100 : 4'b1101;
												assign node7564 = (inp[1]) ? node7576 : node7565;
													assign node7565 = (inp[4]) ? node7571 : node7566;
														assign node7566 = (inp[0]) ? 4'b1110 : node7567;
															assign node7567 = (inp[2]) ? 4'b1110 : 4'b1111;
														assign node7571 = (inp[2]) ? node7573 : 4'b1010;
															assign node7573 = (inp[0]) ? 4'b1010 : 4'b1011;
													assign node7576 = (inp[4]) ? node7582 : node7577;
														assign node7577 = (inp[0]) ? node7579 : 4'b1011;
															assign node7579 = (inp[2]) ? 4'b1010 : 4'b1011;
														assign node7582 = (inp[0]) ? 4'b1111 : node7583;
															assign node7583 = (inp[2]) ? 4'b1110 : 4'b1111;
											assign node7587 = (inp[7]) ? node7609 : node7588;
												assign node7588 = (inp[1]) ? node7598 : node7589;
													assign node7589 = (inp[0]) ? node7591 : 4'b1110;
														assign node7591 = (inp[4]) ? node7595 : node7592;
															assign node7592 = (inp[2]) ? 4'b1111 : 4'b1110;
															assign node7595 = (inp[2]) ? 4'b1110 : 4'b1111;
													assign node7598 = (inp[4]) ? node7604 : node7599;
														assign node7599 = (inp[0]) ? node7601 : 4'b1010;
															assign node7601 = (inp[2]) ? 4'b1011 : 4'b1010;
														assign node7604 = (inp[2]) ? node7606 : 4'b1110;
															assign node7606 = (inp[0]) ? 4'b1110 : 4'b1111;
												assign node7609 = (inp[4]) ? node7623 : node7610;
													assign node7610 = (inp[10]) ? 4'b1101 : node7611;
														assign node7611 = (inp[2]) ? node7617 : node7612;
															assign node7612 = (inp[1]) ? node7614 : 4'b1101;
																assign node7614 = (inp[0]) ? 4'b1101 : 4'b1100;
															assign node7617 = (inp[1]) ? 4'b1101 : node7618;
																assign node7618 = (inp[0]) ? 4'b1100 : 4'b1101;
													assign node7623 = (inp[1]) ? node7629 : node7624;
														assign node7624 = (inp[0]) ? node7626 : 4'b1001;
															assign node7626 = (inp[2]) ? 4'b1001 : 4'b1000;
														assign node7629 = (inp[2]) ? node7631 : 4'b1101;
															assign node7631 = (inp[0]) ? 4'b1101 : 4'b1100;
									assign node7634 = (inp[13]) ? node7730 : node7635;
										assign node7635 = (inp[15]) ? node7683 : node7636;
											assign node7636 = (inp[7]) ? node7660 : node7637;
												assign node7637 = (inp[1]) ? node7649 : node7638;
													assign node7638 = (inp[4]) ? node7644 : node7639;
														assign node7639 = (inp[2]) ? node7641 : 4'b1101;
															assign node7641 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node7644 = (inp[0]) ? 4'b1000 : node7645;
															assign node7645 = (inp[2]) ? 4'b1001 : 4'b1000;
													assign node7649 = (inp[4]) ? node7655 : node7650;
														assign node7650 = (inp[0]) ? 4'b1001 : node7651;
															assign node7651 = (inp[2]) ? 4'b1001 : 4'b1000;
														assign node7655 = (inp[2]) ? node7657 : 4'b1101;
															assign node7657 = (inp[0]) ? 4'b1101 : 4'b1100;
												assign node7660 = (inp[1]) ? node7672 : node7661;
													assign node7661 = (inp[4]) ? node7667 : node7662;
														assign node7662 = (inp[0]) ? 4'b1111 : node7663;
															assign node7663 = (inp[2]) ? 4'b1111 : 4'b1110;
														assign node7667 = (inp[2]) ? 4'b1011 : node7668;
															assign node7668 = (inp[0]) ? 4'b1010 : 4'b1011;
													assign node7672 = (inp[4]) ? node7678 : node7673;
														assign node7673 = (inp[0]) ? node7675 : 4'b1010;
															assign node7675 = (inp[2]) ? 4'b1011 : 4'b1010;
														assign node7678 = (inp[0]) ? node7680 : 4'b1110;
															assign node7680 = (inp[2]) ? 4'b1110 : 4'b1111;
											assign node7683 = (inp[7]) ? node7707 : node7684;
												assign node7684 = (inp[4]) ? node7696 : node7685;
													assign node7685 = (inp[1]) ? node7691 : node7686;
														assign node7686 = (inp[0]) ? node7688 : 4'b1111;
															assign node7688 = (inp[2]) ? 4'b1110 : 4'b1111;
														assign node7691 = (inp[0]) ? node7693 : 4'b1011;
															assign node7693 = (inp[2]) ? 4'b1010 : 4'b1011;
													assign node7696 = (inp[2]) ? node7702 : node7697;
														assign node7697 = (inp[0]) ? 4'b1110 : node7698;
															assign node7698 = (inp[1]) ? 4'b1111 : 4'b1110;
														assign node7702 = (inp[0]) ? node7704 : 4'b1111;
															assign node7704 = (inp[10]) ? 4'b1111 : 4'b1110;
												assign node7707 = (inp[4]) ? node7719 : node7708;
													assign node7708 = (inp[2]) ? node7714 : node7709;
														assign node7709 = (inp[1]) ? node7711 : 4'b1101;
															assign node7711 = (inp[0]) ? 4'b1101 : 4'b1100;
														assign node7714 = (inp[0]) ? node7716 : 4'b1101;
															assign node7716 = (inp[1]) ? 4'b1101 : 4'b1100;
													assign node7719 = (inp[1]) ? node7725 : node7720;
														assign node7720 = (inp[2]) ? node7722 : 4'b1000;
															assign node7722 = (inp[10]) ? 4'b1000 : 4'b1001;
														assign node7725 = (inp[0]) ? node7727 : 4'b1101;
															assign node7727 = (inp[2]) ? 4'b1101 : 4'b1100;
										assign node7730 = (inp[15]) ? node7778 : node7731;
											assign node7731 = (inp[7]) ? node7755 : node7732;
												assign node7732 = (inp[1]) ? node7744 : node7733;
													assign node7733 = (inp[4]) ? node7739 : node7734;
														assign node7734 = (inp[2]) ? 4'b1000 : node7735;
															assign node7735 = (inp[0]) ? 4'b1000 : 4'b1001;
														assign node7739 = (inp[0]) ? 4'b1100 : node7740;
															assign node7740 = (inp[2]) ? 4'b1101 : 4'b1100;
													assign node7744 = (inp[4]) ? node7750 : node7745;
														assign node7745 = (inp[2]) ? 4'b1101 : node7746;
															assign node7746 = (inp[0]) ? 4'b1101 : 4'b1100;
														assign node7750 = (inp[0]) ? node7752 : 4'b1001;
															assign node7752 = (inp[2]) ? 4'b1001 : 4'b1000;
												assign node7755 = (inp[1]) ? node7767 : node7756;
													assign node7756 = (inp[4]) ? node7762 : node7757;
														assign node7757 = (inp[2]) ? node7759 : 4'b1011;
															assign node7759 = (inp[0]) ? 4'b1010 : 4'b1011;
														assign node7762 = (inp[2]) ? 4'b1111 : node7763;
															assign node7763 = (inp[0]) ? 4'b1110 : 4'b1111;
													assign node7767 = (inp[4]) ? node7773 : node7768;
														assign node7768 = (inp[2]) ? node7770 : 4'b1110;
															assign node7770 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node7773 = (inp[0]) ? 4'b1011 : node7774;
															assign node7774 = (inp[2]) ? 4'b1010 : 4'b1011;
											assign node7778 = (inp[7]) ? node7800 : node7779;
												assign node7779 = (inp[1]) ? node7789 : node7780;
													assign node7780 = (inp[2]) ? 4'b1011 : node7781;
														assign node7781 = (inp[0]) ? node7785 : node7782;
															assign node7782 = (inp[4]) ? 4'b1011 : 4'b1010;
															assign node7785 = (inp[4]) ? 4'b1010 : 4'b1011;
													assign node7789 = (inp[4]) ? node7795 : node7790;
														assign node7790 = (inp[2]) ? node7792 : 4'b1110;
															assign node7792 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node7795 = (inp[2]) ? node7797 : 4'b1011;
															assign node7797 = (inp[0]) ? 4'b1011 : 4'b1010;
												assign node7800 = (inp[1]) ? node7812 : node7801;
													assign node7801 = (inp[4]) ? node7807 : node7802;
														assign node7802 = (inp[0]) ? 4'b1001 : node7803;
															assign node7803 = (inp[2]) ? 4'b1001 : 4'b1000;
														assign node7807 = (inp[0]) ? 4'b1101 : node7808;
															assign node7808 = (inp[2]) ? 4'b1100 : 4'b1101;
													assign node7812 = (inp[4]) ? node7814 : 4'b1000;
														assign node7814 = (inp[2]) ? node7816 : 4'b1001;
															assign node7816 = (inp[0]) ? 4'b1001 : 4'b1000;
							assign node7819 = (inp[5]) ? node8169 : node7820;
								assign node7820 = (inp[13]) ? node8002 : node7821;
									assign node7821 = (inp[12]) ? node7907 : node7822;
										assign node7822 = (inp[15]) ? node7856 : node7823;
											assign node7823 = (inp[7]) ? node7847 : node7824;
												assign node7824 = (inp[2]) ? node7826 : 4'b1000;
													assign node7826 = (inp[1]) ? node7840 : node7827;
														assign node7827 = (inp[10]) ? node7835 : node7828;
															assign node7828 = (inp[0]) ? node7832 : node7829;
																assign node7829 = (inp[4]) ? 4'b1001 : 4'b1000;
																assign node7832 = (inp[4]) ? 4'b1000 : 4'b1001;
															assign node7835 = (inp[0]) ? node7837 : 4'b1001;
																assign node7837 = (inp[4]) ? 4'b1000 : 4'b1001;
														assign node7840 = (inp[4]) ? node7844 : node7841;
															assign node7841 = (inp[0]) ? 4'b1001 : 4'b1000;
															assign node7844 = (inp[0]) ? 4'b1000 : 4'b1001;
												assign node7847 = (inp[2]) ? node7849 : 4'b1010;
													assign node7849 = (inp[4]) ? node7853 : node7850;
														assign node7850 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node7853 = (inp[0]) ? 4'b1010 : 4'b1011;
											assign node7856 = (inp[7]) ? node7880 : node7857;
												assign node7857 = (inp[4]) ? node7869 : node7858;
													assign node7858 = (inp[0]) ? node7864 : node7859;
														assign node7859 = (inp[1]) ? node7861 : 4'b1010;
															assign node7861 = (inp[2]) ? 4'b1011 : 4'b1010;
														assign node7864 = (inp[1]) ? 4'b1011 : node7865;
															assign node7865 = (inp[2]) ? 4'b1011 : 4'b1010;
													assign node7869 = (inp[1]) ? node7875 : node7870;
														assign node7870 = (inp[0]) ? 4'b1010 : node7871;
															assign node7871 = (inp[2]) ? 4'b1011 : 4'b1010;
														assign node7875 = (inp[2]) ? 4'b1110 : node7876;
															assign node7876 = (inp[0]) ? 4'b1111 : 4'b1110;
												assign node7880 = (inp[1]) ? node7892 : node7881;
													assign node7881 = (inp[4]) ? node7887 : node7882;
														assign node7882 = (inp[2]) ? node7884 : 4'b1100;
															assign node7884 = (inp[0]) ? 4'b1101 : 4'b1100;
														assign node7887 = (inp[0]) ? node7889 : 4'b1000;
															assign node7889 = (inp[2]) ? 4'b1000 : 4'b1001;
													assign node7892 = (inp[2]) ? node7894 : 4'b1001;
														assign node7894 = (inp[10]) ? node7900 : node7895;
															assign node7895 = (inp[0]) ? node7897 : 4'b1000;
																assign node7897 = (inp[4]) ? 4'b1001 : 4'b1000;
															assign node7900 = (inp[0]) ? node7904 : node7901;
																assign node7901 = (inp[4]) ? 4'b1000 : 4'b1001;
																assign node7904 = (inp[4]) ? 4'b1001 : 4'b1000;
										assign node7907 = (inp[15]) ? node7953 : node7908;
											assign node7908 = (inp[7]) ? node7930 : node7909;
												assign node7909 = (inp[1]) ? node7921 : node7910;
													assign node7910 = (inp[4]) ? node7916 : node7911;
														assign node7911 = (inp[0]) ? node7913 : 4'b1000;
															assign node7913 = (inp[2]) ? 4'b1001 : 4'b1000;
														assign node7916 = (inp[0]) ? 4'b1100 : node7917;
															assign node7917 = (inp[10]) ? 4'b1101 : 4'b1100;
													assign node7921 = (inp[4]) ? node7925 : node7922;
														assign node7922 = (inp[10]) ? 4'b1100 : 4'b1101;
														assign node7925 = (inp[0]) ? node7927 : 4'b1001;
															assign node7927 = (inp[2]) ? 4'b1001 : 4'b1000;
												assign node7930 = (inp[1]) ? node7942 : node7931;
													assign node7931 = (inp[4]) ? node7937 : node7932;
														assign node7932 = (inp[0]) ? 4'b1011 : node7933;
															assign node7933 = (inp[2]) ? 4'b1011 : 4'b1010;
														assign node7937 = (inp[2]) ? 4'b1110 : node7938;
															assign node7938 = (inp[0]) ? 4'b1111 : 4'b1110;
													assign node7942 = (inp[4]) ? node7948 : node7943;
														assign node7943 = (inp[2]) ? 4'b1110 : node7944;
															assign node7944 = (inp[0]) ? 4'b1110 : 4'b1111;
														assign node7948 = (inp[0]) ? 4'b1010 : node7949;
															assign node7949 = (inp[2]) ? 4'b1011 : 4'b1010;
											assign node7953 = (inp[7]) ? node7975 : node7954;
												assign node7954 = (inp[1]) ? node7964 : node7955;
													assign node7955 = (inp[0]) ? node7957 : 4'b1010;
														assign node7957 = (inp[2]) ? node7961 : node7958;
															assign node7958 = (inp[4]) ? 4'b1011 : 4'b1010;
															assign node7961 = (inp[4]) ? 4'b1010 : 4'b1011;
													assign node7964 = (inp[4]) ? node7970 : node7965;
														assign node7965 = (inp[2]) ? 4'b1110 : node7966;
															assign node7966 = (inp[0]) ? 4'b1110 : 4'b1111;
														assign node7970 = (inp[0]) ? 4'b1010 : node7971;
															assign node7971 = (inp[2]) ? 4'b1011 : 4'b1010;
												assign node7975 = (inp[1]) ? node7987 : node7976;
													assign node7976 = (inp[4]) ? node7982 : node7977;
														assign node7977 = (inp[2]) ? node7979 : 4'b1001;
															assign node7979 = (inp[0]) ? 4'b1000 : 4'b1001;
														assign node7982 = (inp[0]) ? 4'b1101 : node7983;
															assign node7983 = (inp[2]) ? 4'b1100 : 4'b1101;
													assign node7987 = (inp[0]) ? 4'b1001 : node7988;
														assign node7988 = (inp[10]) ? node7994 : node7989;
															assign node7989 = (inp[4]) ? node7991 : 4'b1001;
																assign node7991 = (inp[2]) ? 4'b1000 : 4'b1001;
															assign node7994 = (inp[2]) ? node7998 : node7995;
																assign node7995 = (inp[4]) ? 4'b1001 : 4'b1000;
																assign node7998 = (inp[4]) ? 4'b1000 : 4'b1001;
									assign node8002 = (inp[12]) ? node8080 : node8003;
										assign node8003 = (inp[15]) ? node8035 : node8004;
											assign node8004 = (inp[7]) ? node8026 : node8005;
												assign node8005 = (inp[2]) ? node8007 : 4'b1100;
													assign node8007 = (inp[1]) ? node8019 : node8008;
														assign node8008 = (inp[10]) ? node8014 : node8009;
															assign node8009 = (inp[4]) ? node8011 : 4'b1101;
																assign node8011 = (inp[0]) ? 4'b1100 : 4'b1101;
															assign node8014 = (inp[0]) ? 4'b1101 : node8015;
																assign node8015 = (inp[4]) ? 4'b1101 : 4'b1100;
														assign node8019 = (inp[4]) ? node8023 : node8020;
															assign node8020 = (inp[0]) ? 4'b1101 : 4'b1100;
															assign node8023 = (inp[0]) ? 4'b1100 : 4'b1101;
												assign node8026 = (inp[2]) ? node8028 : 4'b1110;
													assign node8028 = (inp[0]) ? node8032 : node8029;
														assign node8029 = (inp[4]) ? 4'b1111 : 4'b1110;
														assign node8032 = (inp[4]) ? 4'b1110 : 4'b1111;
											assign node8035 = (inp[7]) ? node8055 : node8036;
												assign node8036 = (inp[1]) ? node8046 : node8037;
													assign node8037 = (inp[2]) ? node8039 : 4'b1111;
														assign node8039 = (inp[4]) ? node8043 : node8040;
															assign node8040 = (inp[0]) ? 4'b1110 : 4'b1111;
															assign node8043 = (inp[0]) ? 4'b1111 : 4'b1110;
													assign node8046 = (inp[4]) ? node8050 : node8047;
														assign node8047 = (inp[0]) ? 4'b1110 : 4'b1111;
														assign node8050 = (inp[2]) ? node8052 : 4'b1010;
															assign node8052 = (inp[0]) ? 4'b1010 : 4'b1011;
												assign node8055 = (inp[1]) ? node8065 : node8056;
													assign node8056 = (inp[4]) ? node8062 : node8057;
														assign node8057 = (inp[2]) ? 4'b1000 : node8058;
															assign node8058 = (inp[0]) ? 4'b1000 : 4'b1001;
														assign node8062 = (inp[0]) ? 4'b1100 : 4'b1101;
													assign node8065 = (inp[2]) ? node8067 : 4'b1100;
														assign node8067 = (inp[10]) ? node8075 : node8068;
															assign node8068 = (inp[0]) ? node8072 : node8069;
																assign node8069 = (inp[4]) ? 4'b1101 : 4'b1100;
																assign node8072 = (inp[4]) ? 4'b1100 : 4'b1101;
															assign node8075 = (inp[4]) ? 4'b1100 : node8076;
																assign node8076 = (inp[0]) ? 4'b1101 : 4'b1100;
										assign node8080 = (inp[15]) ? node8124 : node8081;
											assign node8081 = (inp[7]) ? node8101 : node8082;
												assign node8082 = (inp[1]) ? node8094 : node8083;
													assign node8083 = (inp[4]) ? node8089 : node8084;
														assign node8084 = (inp[2]) ? node8086 : 4'b1100;
															assign node8086 = (inp[0]) ? 4'b1101 : 4'b1100;
														assign node8089 = (inp[0]) ? node8091 : 4'b1000;
															assign node8091 = (inp[2]) ? 4'b1000 : 4'b1001;
													assign node8094 = (inp[4]) ? 4'b1101 : node8095;
														assign node8095 = (inp[2]) ? 4'b1000 : node8096;
															assign node8096 = (inp[0]) ? 4'b1000 : 4'b1001;
												assign node8101 = (inp[1]) ? node8113 : node8102;
													assign node8102 = (inp[4]) ? node8108 : node8103;
														assign node8103 = (inp[2]) ? 4'b1111 : node8104;
															assign node8104 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node8108 = (inp[2]) ? node8110 : 4'b1011;
															assign node8110 = (inp[0]) ? 4'b1011 : 4'b1010;
													assign node8113 = (inp[4]) ? node8119 : node8114;
														assign node8114 = (inp[0]) ? node8116 : 4'b1010;
															assign node8116 = (inp[2]) ? 4'b1011 : 4'b1010;
														assign node8119 = (inp[0]) ? 4'b1110 : node8120;
															assign node8120 = (inp[10]) ? 4'b1111 : 4'b1110;
											assign node8124 = (inp[7]) ? node8148 : node8125;
												assign node8125 = (inp[4]) ? node8137 : node8126;
													assign node8126 = (inp[1]) ? node8132 : node8127;
														assign node8127 = (inp[2]) ? node8129 : 4'b1111;
															assign node8129 = (inp[0]) ? 4'b1110 : 4'b1111;
														assign node8132 = (inp[2]) ? node8134 : 4'b1011;
															assign node8134 = (inp[0]) ? 4'b1010 : 4'b1011;
													assign node8137 = (inp[1]) ? node8143 : node8138;
														assign node8138 = (inp[2]) ? 4'b1111 : node8139;
															assign node8139 = (inp[0]) ? 4'b1110 : 4'b1111;
														assign node8143 = (inp[0]) ? 4'b1111 : node8144;
															assign node8144 = (inp[2]) ? 4'b1110 : 4'b1111;
												assign node8148 = (inp[1]) ? node8160 : node8149;
													assign node8149 = (inp[4]) ? node8155 : node8150;
														assign node8150 = (inp[0]) ? node8152 : 4'b1100;
															assign node8152 = (inp[2]) ? 4'b1101 : 4'b1100;
														assign node8155 = (inp[0]) ? node8157 : 4'b1000;
															assign node8157 = (inp[2]) ? 4'b1000 : 4'b1001;
													assign node8160 = (inp[0]) ? 4'b1100 : node8161;
														assign node8161 = (inp[4]) ? node8165 : node8162;
															assign node8162 = (inp[2]) ? 4'b1100 : 4'b1101;
															assign node8165 = (inp[2]) ? 4'b1101 : 4'b1100;
								assign node8169 = (inp[13]) ? node8345 : node8170;
									assign node8170 = (inp[12]) ? node8252 : node8171;
										assign node8171 = (inp[15]) ? node8207 : node8172;
											assign node8172 = (inp[7]) ? node8182 : node8173;
												assign node8173 = (inp[0]) ? node8175 : 4'b1100;
													assign node8175 = (inp[4]) ? node8179 : node8176;
														assign node8176 = (inp[2]) ? 4'b1101 : 4'b1100;
														assign node8179 = (inp[2]) ? 4'b1100 : 4'b1101;
												assign node8182 = (inp[0]) ? node8184 : 4'b1111;
													assign node8184 = (inp[1]) ? node8200 : node8185;
														assign node8185 = (inp[10]) ? node8193 : node8186;
															assign node8186 = (inp[4]) ? node8190 : node8187;
																assign node8187 = (inp[2]) ? 4'b1110 : 4'b1111;
																assign node8190 = (inp[2]) ? 4'b1111 : 4'b1110;
															assign node8193 = (inp[2]) ? node8197 : node8194;
																assign node8194 = (inp[4]) ? 4'b1110 : 4'b1111;
																assign node8197 = (inp[4]) ? 4'b1111 : 4'b1110;
														assign node8200 = (inp[4]) ? node8204 : node8201;
															assign node8201 = (inp[2]) ? 4'b1110 : 4'b1111;
															assign node8204 = (inp[2]) ? 4'b1111 : 4'b1110;
											assign node8207 = (inp[7]) ? node8231 : node8208;
												assign node8208 = (inp[1]) ? node8220 : node8209;
													assign node8209 = (inp[0]) ? node8211 : 4'b1110;
														assign node8211 = (inp[10]) ? node8217 : node8212;
															assign node8212 = (inp[2]) ? node8214 : 4'b1111;
																assign node8214 = (inp[4]) ? 4'b1110 : 4'b1111;
															assign node8217 = (inp[4]) ? 4'b1111 : 4'b1110;
													assign node8220 = (inp[4]) ? node8226 : node8221;
														assign node8221 = (inp[2]) ? 4'b1111 : node8222;
															assign node8222 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node8226 = (inp[2]) ? 4'b1011 : node8227;
															assign node8227 = (inp[0]) ? 4'b1010 : 4'b1011;
												assign node8231 = (inp[1]) ? node8243 : node8232;
													assign node8232 = (inp[4]) ? node8238 : node8233;
														assign node8233 = (inp[2]) ? 4'b1000 : node8234;
															assign node8234 = (inp[0]) ? 4'b1000 : 4'b1001;
														assign node8238 = (inp[0]) ? 4'b1100 : node8239;
															assign node8239 = (inp[2]) ? 4'b1101 : 4'b1100;
													assign node8243 = (inp[0]) ? node8245 : 4'b1100;
														assign node8245 = (inp[4]) ? node8249 : node8246;
															assign node8246 = (inp[2]) ? 4'b1101 : 4'b1100;
															assign node8249 = (inp[2]) ? 4'b1100 : 4'b1101;
										assign node8252 = (inp[15]) ? node8300 : node8253;
											assign node8253 = (inp[7]) ? node8277 : node8254;
												assign node8254 = (inp[4]) ? node8266 : node8255;
													assign node8255 = (inp[1]) ? node8261 : node8256;
														assign node8256 = (inp[0]) ? node8258 : 4'b1100;
															assign node8258 = (inp[2]) ? 4'b1101 : 4'b1100;
														assign node8261 = (inp[0]) ? 4'b1000 : node8262;
															assign node8262 = (inp[2]) ? 4'b1000 : 4'b1001;
													assign node8266 = (inp[1]) ? node8272 : node8267;
														assign node8267 = (inp[0]) ? 4'b1001 : node8268;
															assign node8268 = (inp[2]) ? 4'b1000 : 4'b1001;
														assign node8272 = (inp[2]) ? node8274 : 4'b1100;
															assign node8274 = (inp[0]) ? 4'b1100 : 4'b1101;
												assign node8277 = (inp[1]) ? node8289 : node8278;
													assign node8278 = (inp[4]) ? node8284 : node8279;
														assign node8279 = (inp[2]) ? 4'b1110 : node8280;
															assign node8280 = (inp[0]) ? 4'b1110 : 4'b1111;
														assign node8284 = (inp[0]) ? node8286 : 4'b1010;
															assign node8286 = (inp[2]) ? 4'b1010 : 4'b1011;
													assign node8289 = (inp[4]) ? node8295 : node8290;
														assign node8290 = (inp[0]) ? node8292 : 4'b1011;
															assign node8292 = (inp[2]) ? 4'b1010 : 4'b1011;
														assign node8295 = (inp[2]) ? 4'b1111 : node8296;
															assign node8296 = (inp[0]) ? 4'b1110 : 4'b1111;
											assign node8300 = (inp[7]) ? node8324 : node8301;
												assign node8301 = (inp[1]) ? node8313 : node8302;
													assign node8302 = (inp[0]) ? node8308 : node8303;
														assign node8303 = (inp[2]) ? 4'b1110 : node8304;
															assign node8304 = (inp[4]) ? 4'b1111 : 4'b1110;
														assign node8308 = (inp[2]) ? 4'b1111 : node8309;
															assign node8309 = (inp[4]) ? 4'b1111 : 4'b1110;
													assign node8313 = (inp[4]) ? node8319 : node8314;
														assign node8314 = (inp[2]) ? node8316 : 4'b1010;
															assign node8316 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node8319 = (inp[0]) ? node8321 : 4'b1110;
															assign node8321 = (inp[2]) ? 4'b1110 : 4'b1111;
												assign node8324 = (inp[4]) ? node8336 : node8325;
													assign node8325 = (inp[2]) ? node8331 : node8326;
														assign node8326 = (inp[1]) ? node8328 : 4'b1100;
															assign node8328 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node8331 = (inp[0]) ? node8333 : 4'b1100;
															assign node8333 = (inp[1]) ? 4'b1100 : 4'b1101;
													assign node8336 = (inp[1]) ? node8342 : node8337;
														assign node8337 = (inp[2]) ? node8339 : 4'b1001;
															assign node8339 = (inp[0]) ? 4'b1001 : 4'b1000;
														assign node8342 = (inp[0]) ? 4'b1101 : 4'b1100;
									assign node8345 = (inp[12]) ? node8429 : node8346;
										assign node8346 = (inp[15]) ? node8382 : node8347;
											assign node8347 = (inp[7]) ? node8357 : node8348;
												assign node8348 = (inp[0]) ? 4'b1001 : node8349;
													assign node8349 = (inp[2]) ? node8353 : node8350;
														assign node8350 = (inp[4]) ? 4'b1001 : 4'b1000;
														assign node8353 = (inp[4]) ? 4'b1000 : 4'b1001;
												assign node8357 = (inp[0]) ? 4'b1010 : node8358;
													assign node8358 = (inp[10]) ? node8374 : node8359;
														assign node8359 = (inp[1]) ? node8367 : node8360;
															assign node8360 = (inp[2]) ? node8364 : node8361;
																assign node8361 = (inp[4]) ? 4'b1010 : 4'b1011;
																assign node8364 = (inp[4]) ? 4'b1011 : 4'b1010;
															assign node8367 = (inp[4]) ? node8371 : node8368;
																assign node8368 = (inp[2]) ? 4'b1010 : 4'b1011;
																assign node8371 = (inp[2]) ? 4'b1011 : 4'b1010;
														assign node8374 = (inp[2]) ? node8378 : node8375;
															assign node8375 = (inp[4]) ? 4'b1010 : 4'b1011;
															assign node8378 = (inp[4]) ? 4'b1011 : 4'b1010;
											assign node8382 = (inp[7]) ? node8402 : node8383;
												assign node8383 = (inp[1]) ? node8391 : node8384;
													assign node8384 = (inp[0]) ? 4'b1010 : node8385;
														assign node8385 = (inp[2]) ? node8387 : 4'b1010;
															assign node8387 = (inp[4]) ? 4'b1011 : 4'b1010;
													assign node8391 = (inp[4]) ? node8397 : node8392;
														assign node8392 = (inp[0]) ? node8394 : 4'b1010;
															assign node8394 = (inp[2]) ? 4'b1011 : 4'b1010;
														assign node8397 = (inp[0]) ? node8399 : 4'b1110;
															assign node8399 = (inp[2]) ? 4'b1110 : 4'b1111;
												assign node8402 = (inp[1]) ? node8414 : node8403;
													assign node8403 = (inp[4]) ? node8409 : node8404;
														assign node8404 = (inp[0]) ? 4'b1101 : node8405;
															assign node8405 = (inp[2]) ? 4'b1101 : 4'b1100;
														assign node8409 = (inp[0]) ? node8411 : 4'b1001;
															assign node8411 = (inp[2]) ? 4'b1001 : 4'b1000;
													assign node8414 = (inp[0]) ? 4'b1000 : node8415;
														assign node8415 = (inp[10]) ? node8423 : node8416;
															assign node8416 = (inp[4]) ? node8420 : node8417;
																assign node8417 = (inp[2]) ? 4'b1000 : 4'b1001;
																assign node8420 = (inp[2]) ? 4'b1001 : 4'b1000;
															assign node8423 = (inp[4]) ? 4'b1000 : node8424;
																assign node8424 = (inp[2]) ? 4'b1000 : 4'b1001;
										assign node8429 = (inp[15]) ? node8477 : node8430;
											assign node8430 = (inp[7]) ? node8454 : node8431;
												assign node8431 = (inp[1]) ? node8443 : node8432;
													assign node8432 = (inp[4]) ? node8438 : node8433;
														assign node8433 = (inp[0]) ? 4'b1001 : node8434;
															assign node8434 = (inp[2]) ? 4'b1001 : 4'b1000;
														assign node8438 = (inp[0]) ? 4'b1101 : node8439;
															assign node8439 = (inp[2]) ? 4'b1100 : 4'b1101;
													assign node8443 = (inp[4]) ? node8449 : node8444;
														assign node8444 = (inp[0]) ? 4'b1100 : node8445;
															assign node8445 = (inp[2]) ? 4'b1100 : 4'b1101;
														assign node8449 = (inp[2]) ? 4'b1000 : node8450;
															assign node8450 = (inp[0]) ? 4'b1001 : 4'b1000;
												assign node8454 = (inp[4]) ? node8466 : node8455;
													assign node8455 = (inp[1]) ? node8461 : node8456;
														assign node8456 = (inp[2]) ? node8458 : 4'b1010;
															assign node8458 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node8461 = (inp[2]) ? node8463 : 4'b1111;
															assign node8463 = (inp[0]) ? 4'b1110 : 4'b1111;
													assign node8466 = (inp[1]) ? node8472 : node8467;
														assign node8467 = (inp[2]) ? 4'b1110 : node8468;
															assign node8468 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node8472 = (inp[2]) ? node8474 : 4'b1010;
															assign node8474 = (inp[0]) ? 4'b1010 : 4'b1011;
											assign node8477 = (inp[7]) ? node8507 : node8478;
												assign node8478 = (inp[1]) ? node8496 : node8479;
													assign node8479 = (inp[2]) ? 4'b1010 : node8480;
														assign node8480 = (inp[10]) ? node8488 : node8481;
															assign node8481 = (inp[4]) ? node8485 : node8482;
																assign node8482 = (inp[0]) ? 4'b1010 : 4'b1011;
																assign node8485 = (inp[0]) ? 4'b1011 : 4'b1010;
															assign node8488 = (inp[4]) ? node8492 : node8489;
																assign node8489 = (inp[0]) ? 4'b1010 : 4'b1011;
																assign node8492 = (inp[0]) ? 4'b1011 : 4'b1010;
													assign node8496 = (inp[4]) ? node8502 : node8497;
														assign node8497 = (inp[0]) ? node8499 : 4'b1111;
															assign node8499 = (inp[2]) ? 4'b1110 : 4'b1111;
														assign node8502 = (inp[2]) ? node8504 : 4'b1010;
															assign node8504 = (inp[0]) ? 4'b1010 : 4'b1011;
												assign node8507 = (inp[4]) ? node8519 : node8508;
													assign node8508 = (inp[1]) ? node8514 : node8509;
														assign node8509 = (inp[2]) ? 4'b1000 : node8510;
															assign node8510 = (inp[0]) ? 4'b1000 : 4'b1001;
														assign node8514 = (inp[2]) ? node8516 : 4'b1001;
															assign node8516 = (inp[0]) ? 4'b1000 : 4'b1001;
													assign node8519 = (inp[1]) ? node8525 : node8520;
														assign node8520 = (inp[0]) ? 4'b1100 : node8521;
															assign node8521 = (inp[2]) ? 4'b1101 : 4'b1100;
														assign node8525 = (inp[2]) ? node8527 : 4'b1000;
															assign node8527 = (inp[0]) ? 4'b1000 : 4'b1001;
				assign node8530 = (inp[13]) ? node13134 : node8531;
					assign node8531 = (inp[5]) ? node10819 : node8532;
						assign node8532 = (inp[6]) ? node9940 : node8533;
							assign node8533 = (inp[7]) ? node9191 : node8534;
								assign node8534 = (inp[12]) ? node8866 : node8535;
									assign node8535 = (inp[4]) ? node8683 : node8536;
										assign node8536 = (inp[1]) ? node8596 : node8537;
											assign node8537 = (inp[2]) ? node8561 : node8538;
												assign node8538 = (inp[10]) ? node8550 : node8539;
													assign node8539 = (inp[9]) ? node8545 : node8540;
														assign node8540 = (inp[0]) ? node8542 : 4'b1000;
															assign node8542 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node8545 = (inp[0]) ? node8547 : 4'b1001;
															assign node8547 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node8550 = (inp[9]) ? node8556 : node8551;
														assign node8551 = (inp[11]) ? 4'b1001 : node8552;
															assign node8552 = (inp[0]) ? 4'b1000 : 4'b1001;
														assign node8556 = (inp[11]) ? 4'b1000 : node8557;
															assign node8557 = (inp[0]) ? 4'b1001 : 4'b1000;
												assign node8561 = (inp[11]) ? node8583 : node8562;
													assign node8562 = (inp[15]) ? node8570 : node8563;
														assign node8563 = (inp[10]) ? 4'b1100 : node8564;
															assign node8564 = (inp[9]) ? node8566 : 4'b1100;
																assign node8566 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node8570 = (inp[9]) ? node8578 : node8571;
															assign node8571 = (inp[0]) ? node8575 : node8572;
																assign node8572 = (inp[10]) ? 4'b1101 : 4'b1100;
																assign node8575 = (inp[10]) ? 4'b1100 : 4'b1101;
															assign node8578 = (inp[0]) ? node8580 : 4'b1100;
																assign node8580 = (inp[10]) ? 4'b1101 : 4'b1100;
													assign node8583 = (inp[15]) ? node8591 : node8584;
														assign node8584 = (inp[10]) ? node8588 : node8585;
															assign node8585 = (inp[9]) ? 4'b1101 : 4'b1100;
															assign node8588 = (inp[9]) ? 4'b1100 : 4'b1101;
														assign node8591 = (inp[9]) ? 4'b1100 : node8592;
															assign node8592 = (inp[10]) ? 4'b1101 : 4'b1100;
											assign node8596 = (inp[2]) ? node8638 : node8597;
												assign node8597 = (inp[10]) ? node8619 : node8598;
													assign node8598 = (inp[9]) ? node8610 : node8599;
														assign node8599 = (inp[0]) ? node8605 : node8600;
															assign node8600 = (inp[11]) ? node8602 : 4'b1100;
																assign node8602 = (inp[15]) ? 4'b1101 : 4'b1100;
															assign node8605 = (inp[11]) ? 4'b1100 : node8606;
																assign node8606 = (inp[15]) ? 4'b1100 : 4'b1101;
														assign node8610 = (inp[11]) ? node8614 : node8611;
															assign node8611 = (inp[0]) ? 4'b1100 : 4'b1101;
															assign node8614 = (inp[15]) ? node8616 : 4'b1101;
																assign node8616 = (inp[0]) ? 4'b1101 : 4'b1100;
													assign node8619 = (inp[9]) ? node8631 : node8620;
														assign node8620 = (inp[15]) ? node8626 : node8621;
															assign node8621 = (inp[11]) ? 4'b1101 : node8622;
																assign node8622 = (inp[0]) ? 4'b1100 : 4'b1101;
															assign node8626 = (inp[0]) ? 4'b1101 : node8627;
																assign node8627 = (inp[11]) ? 4'b1100 : 4'b1101;
														assign node8631 = (inp[15]) ? 4'b1101 : node8632;
															assign node8632 = (inp[11]) ? 4'b1100 : node8633;
																assign node8633 = (inp[0]) ? 4'b1101 : 4'b1100;
												assign node8638 = (inp[15]) ? node8654 : node8639;
													assign node8639 = (inp[9]) ? node8651 : node8640;
														assign node8640 = (inp[10]) ? node8646 : node8641;
															assign node8641 = (inp[0]) ? 4'b1000 : node8642;
																assign node8642 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node8646 = (inp[0]) ? 4'b1001 : node8647;
																assign node8647 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node8651 = (inp[10]) ? 4'b1000 : 4'b1001;
													assign node8654 = (inp[11]) ? node8668 : node8655;
														assign node8655 = (inp[10]) ? node8663 : node8656;
															assign node8656 = (inp[9]) ? node8660 : node8657;
																assign node8657 = (inp[0]) ? 4'b1000 : 4'b1001;
																assign node8660 = (inp[0]) ? 4'b1001 : 4'b1000;
															assign node8663 = (inp[9]) ? node8665 : 4'b1000;
																assign node8665 = (inp[0]) ? 4'b1000 : 4'b1001;
														assign node8668 = (inp[0]) ? node8676 : node8669;
															assign node8669 = (inp[10]) ? node8673 : node8670;
																assign node8670 = (inp[9]) ? 4'b1000 : 4'b1001;
																assign node8673 = (inp[9]) ? 4'b1001 : 4'b1000;
															assign node8676 = (inp[10]) ? node8680 : node8677;
																assign node8677 = (inp[9]) ? 4'b1000 : 4'b1001;
																assign node8680 = (inp[9]) ? 4'b1001 : 4'b1000;
										assign node8683 = (inp[15]) ? node8779 : node8684;
											assign node8684 = (inp[0]) ? node8730 : node8685;
												assign node8685 = (inp[9]) ? node8711 : node8686;
													assign node8686 = (inp[11]) ? node8698 : node8687;
														assign node8687 = (inp[1]) ? node8693 : node8688;
															assign node8688 = (inp[2]) ? node8690 : 4'b1011;
																assign node8690 = (inp[10]) ? 4'b1110 : 4'b1111;
															assign node8693 = (inp[2]) ? 4'b1011 : node8694;
																assign node8694 = (inp[10]) ? 4'b1111 : 4'b1110;
														assign node8698 = (inp[10]) ? node8704 : node8699;
															assign node8699 = (inp[1]) ? 4'b1010 : node8700;
																assign node8700 = (inp[2]) ? 4'b1111 : 4'b1010;
															assign node8704 = (inp[2]) ? node8708 : node8705;
																assign node8705 = (inp[1]) ? 4'b1111 : 4'b1011;
																assign node8708 = (inp[1]) ? 4'b1011 : 4'b1110;
													assign node8711 = (inp[10]) ? node8721 : node8712;
														assign node8712 = (inp[2]) ? node8716 : node8713;
															assign node8713 = (inp[1]) ? 4'b1111 : 4'b1011;
															assign node8716 = (inp[1]) ? node8718 : 4'b1110;
																assign node8718 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node8721 = (inp[2]) ? node8725 : node8722;
															assign node8722 = (inp[1]) ? 4'b1110 : 4'b1010;
															assign node8725 = (inp[1]) ? node8727 : 4'b1111;
																assign node8727 = (inp[11]) ? 4'b1010 : 4'b1011;
												assign node8730 = (inp[1]) ? node8752 : node8731;
													assign node8731 = (inp[2]) ? node8745 : node8732;
														assign node8732 = (inp[11]) ? node8740 : node8733;
															assign node8733 = (inp[9]) ? node8737 : node8734;
																assign node8734 = (inp[10]) ? 4'b1010 : 4'b1011;
																assign node8737 = (inp[10]) ? 4'b1011 : 4'b1010;
															assign node8740 = (inp[9]) ? node8742 : 4'b1010;
																assign node8742 = (inp[10]) ? 4'b1010 : 4'b1011;
														assign node8745 = (inp[10]) ? node8747 : 4'b1110;
															assign node8747 = (inp[9]) ? 4'b1110 : node8748;
																assign node8748 = (inp[11]) ? 4'b1110 : 4'b1111;
													assign node8752 = (inp[2]) ? node8764 : node8753;
														assign node8753 = (inp[10]) ? node8759 : node8754;
															assign node8754 = (inp[9]) ? node8756 : 4'b1110;
																assign node8756 = (inp[11]) ? 4'b1111 : 4'b1110;
															assign node8759 = (inp[11]) ? node8761 : 4'b1111;
																assign node8761 = (inp[9]) ? 4'b1110 : 4'b1111;
														assign node8764 = (inp[11]) ? node8772 : node8765;
															assign node8765 = (inp[9]) ? node8769 : node8766;
																assign node8766 = (inp[10]) ? 4'b1010 : 4'b1011;
																assign node8769 = (inp[10]) ? 4'b1011 : 4'b1010;
															assign node8772 = (inp[10]) ? node8776 : node8773;
																assign node8773 = (inp[9]) ? 4'b1010 : 4'b1011;
																assign node8776 = (inp[9]) ? 4'b1011 : 4'b1010;
											assign node8779 = (inp[2]) ? node8823 : node8780;
												assign node8780 = (inp[1]) ? node8802 : node8781;
													assign node8781 = (inp[10]) ? node8791 : node8782;
														assign node8782 = (inp[9]) ? node8788 : node8783;
															assign node8783 = (inp[0]) ? node8785 : 4'b1100;
																assign node8785 = (inp[11]) ? 4'b1100 : 4'b1101;
															assign node8788 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node8791 = (inp[9]) ? node8797 : node8792;
															assign node8792 = (inp[0]) ? node8794 : 4'b1101;
																assign node8794 = (inp[11]) ? 4'b1101 : 4'b1100;
															assign node8797 = (inp[0]) ? node8799 : 4'b1100;
																assign node8799 = (inp[11]) ? 4'b1100 : 4'b1101;
													assign node8802 = (inp[9]) ? node8814 : node8803;
														assign node8803 = (inp[10]) ? node8809 : node8804;
															assign node8804 = (inp[0]) ? node8806 : 4'b1001;
																assign node8806 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node8809 = (inp[0]) ? node8811 : 4'b1000;
																assign node8811 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node8814 = (inp[10]) ? node8820 : node8815;
															assign node8815 = (inp[11]) ? 4'b1000 : node8816;
																assign node8816 = (inp[0]) ? 4'b1001 : 4'b1000;
															assign node8820 = (inp[11]) ? 4'b1001 : 4'b1000;
												assign node8823 = (inp[1]) ? node8845 : node8824;
													assign node8824 = (inp[0]) ? node8840 : node8825;
														assign node8825 = (inp[9]) ? node8833 : node8826;
															assign node8826 = (inp[10]) ? node8830 : node8827;
																assign node8827 = (inp[11]) ? 4'b1000 : 4'b1001;
																assign node8830 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node8833 = (inp[11]) ? node8837 : node8834;
																assign node8834 = (inp[10]) ? 4'b1001 : 4'b1000;
																assign node8837 = (inp[10]) ? 4'b1000 : 4'b1001;
														assign node8840 = (inp[9]) ? 4'b1001 : node8841;
															assign node8841 = (inp[10]) ? 4'b1000 : 4'b1001;
													assign node8845 = (inp[10]) ? node8855 : node8846;
														assign node8846 = (inp[0]) ? node8848 : 4'b1101;
															assign node8848 = (inp[9]) ? node8852 : node8849;
																assign node8849 = (inp[11]) ? 4'b1100 : 4'b1101;
																assign node8852 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node8855 = (inp[9]) ? node8861 : node8856;
															assign node8856 = (inp[0]) ? node8858 : 4'b1101;
																assign node8858 = (inp[11]) ? 4'b1101 : 4'b1100;
															assign node8861 = (inp[0]) ? node8863 : 4'b1100;
																assign node8863 = (inp[11]) ? 4'b1100 : 4'b1101;
									assign node8866 = (inp[4]) ? node9032 : node8867;
										assign node8867 = (inp[0]) ? node8921 : node8868;
											assign node8868 = (inp[9]) ? node8892 : node8869;
												assign node8869 = (inp[10]) ? node8881 : node8870;
													assign node8870 = (inp[1]) ? node8874 : node8871;
														assign node8871 = (inp[2]) ? 4'b1110 : 4'b1010;
														assign node8874 = (inp[2]) ? 4'b1010 : node8875;
															assign node8875 = (inp[11]) ? node8877 : 4'b1111;
																assign node8877 = (inp[15]) ? 4'b1110 : 4'b1111;
													assign node8881 = (inp[1]) ? node8885 : node8882;
														assign node8882 = (inp[2]) ? 4'b1111 : 4'b1011;
														assign node8885 = (inp[11]) ? node8889 : node8886;
															assign node8886 = (inp[2]) ? 4'b1010 : 4'b1110;
															assign node8889 = (inp[2]) ? 4'b1011 : 4'b1111;
												assign node8892 = (inp[10]) ? node8906 : node8893;
													assign node8893 = (inp[1]) ? node8897 : node8894;
														assign node8894 = (inp[2]) ? 4'b1111 : 4'b1011;
														assign node8897 = (inp[2]) ? node8901 : node8898;
															assign node8898 = (inp[11]) ? 4'b1111 : 4'b1110;
															assign node8901 = (inp[15]) ? 4'b1011 : node8902;
																assign node8902 = (inp[11]) ? 4'b1011 : 4'b1010;
													assign node8906 = (inp[1]) ? node8910 : node8907;
														assign node8907 = (inp[2]) ? 4'b1110 : 4'b1010;
														assign node8910 = (inp[2]) ? node8916 : node8911;
															assign node8911 = (inp[11]) ? node8913 : 4'b1111;
																assign node8913 = (inp[15]) ? 4'b1110 : 4'b1111;
															assign node8916 = (inp[15]) ? 4'b1010 : node8917;
																assign node8917 = (inp[11]) ? 4'b1010 : 4'b1011;
											assign node8921 = (inp[15]) ? node8979 : node8922;
												assign node8922 = (inp[10]) ? node8952 : node8923;
													assign node8923 = (inp[9]) ? node8937 : node8924;
														assign node8924 = (inp[11]) ? node8930 : node8925;
															assign node8925 = (inp[1]) ? 4'b1110 : node8926;
																assign node8926 = (inp[2]) ? 4'b1111 : 4'b1011;
															assign node8930 = (inp[1]) ? node8934 : node8931;
																assign node8931 = (inp[2]) ? 4'b1110 : 4'b1010;
																assign node8934 = (inp[2]) ? 4'b1011 : 4'b1111;
														assign node8937 = (inp[11]) ? node8945 : node8938;
															assign node8938 = (inp[1]) ? node8942 : node8939;
																assign node8939 = (inp[2]) ? 4'b1110 : 4'b1010;
																assign node8942 = (inp[2]) ? 4'b1010 : 4'b1111;
															assign node8945 = (inp[1]) ? node8949 : node8946;
																assign node8946 = (inp[2]) ? 4'b1111 : 4'b1011;
																assign node8949 = (inp[2]) ? 4'b1010 : 4'b1110;
													assign node8952 = (inp[11]) ? node8964 : node8953;
														assign node8953 = (inp[1]) ? node8957 : node8954;
															assign node8954 = (inp[9]) ? 4'b1011 : 4'b1010;
															assign node8957 = (inp[2]) ? node8961 : node8958;
																assign node8958 = (inp[9]) ? 4'b1110 : 4'b1111;
																assign node8961 = (inp[9]) ? 4'b1011 : 4'b1010;
														assign node8964 = (inp[1]) ? node8972 : node8965;
															assign node8965 = (inp[9]) ? node8969 : node8966;
																assign node8966 = (inp[2]) ? 4'b1111 : 4'b1011;
																assign node8969 = (inp[2]) ? 4'b1110 : 4'b1010;
															assign node8972 = (inp[9]) ? node8976 : node8973;
																assign node8973 = (inp[2]) ? 4'b1010 : 4'b1110;
																assign node8976 = (inp[2]) ? 4'b1011 : 4'b1111;
												assign node8979 = (inp[11]) ? node9009 : node8980;
													assign node8980 = (inp[10]) ? node8994 : node8981;
														assign node8981 = (inp[9]) ? node8987 : node8982;
															assign node8982 = (inp[1]) ? 4'b1011 : node8983;
																assign node8983 = (inp[2]) ? 4'b1111 : 4'b1011;
															assign node8987 = (inp[1]) ? node8991 : node8988;
																assign node8988 = (inp[2]) ? 4'b1110 : 4'b1010;
																assign node8991 = (inp[2]) ? 4'b1010 : 4'b1110;
														assign node8994 = (inp[9]) ? node9002 : node8995;
															assign node8995 = (inp[2]) ? node8999 : node8996;
																assign node8996 = (inp[1]) ? 4'b1110 : 4'b1010;
																assign node8999 = (inp[1]) ? 4'b1010 : 4'b1110;
															assign node9002 = (inp[2]) ? node9006 : node9003;
																assign node9003 = (inp[1]) ? 4'b1111 : 4'b1011;
																assign node9006 = (inp[1]) ? 4'b1011 : 4'b1111;
													assign node9009 = (inp[9]) ? node9025 : node9010;
														assign node9010 = (inp[10]) ? node9018 : node9011;
															assign node9011 = (inp[1]) ? node9015 : node9012;
																assign node9012 = (inp[2]) ? 4'b1110 : 4'b1010;
																assign node9015 = (inp[2]) ? 4'b1010 : 4'b1111;
															assign node9018 = (inp[2]) ? node9022 : node9019;
																assign node9019 = (inp[1]) ? 4'b1110 : 4'b1011;
																assign node9022 = (inp[1]) ? 4'b1011 : 4'b1111;
														assign node9025 = (inp[10]) ? 4'b1010 : node9026;
															assign node9026 = (inp[2]) ? node9028 : 4'b1011;
																assign node9028 = (inp[1]) ? 4'b1011 : 4'b1111;
										assign node9032 = (inp[15]) ? node9114 : node9033;
											assign node9033 = (inp[2]) ? node9071 : node9034;
												assign node9034 = (inp[10]) ? node9054 : node9035;
													assign node9035 = (inp[0]) ? node9045 : node9036;
														assign node9036 = (inp[9]) ? node9040 : node9037;
															assign node9037 = (inp[1]) ? 4'b1101 : 4'b1100;
															assign node9040 = (inp[11]) ? 4'b1101 : node9041;
																assign node9041 = (inp[1]) ? 4'b1100 : 4'b1101;
														assign node9045 = (inp[9]) ? node9051 : node9046;
															assign node9046 = (inp[1]) ? 4'b1101 : node9047;
																assign node9047 = (inp[11]) ? 4'b1100 : 4'b1101;
															assign node9051 = (inp[11]) ? 4'b1101 : 4'b1100;
													assign node9054 = (inp[0]) ? node9064 : node9055;
														assign node9055 = (inp[11]) ? 4'b1100 : node9056;
															assign node9056 = (inp[1]) ? node9060 : node9057;
																assign node9057 = (inp[9]) ? 4'b1100 : 4'b1101;
																assign node9060 = (inp[9]) ? 4'b1101 : 4'b1100;
														assign node9064 = (inp[9]) ? node9068 : node9065;
															assign node9065 = (inp[1]) ? 4'b1100 : 4'b1101;
															assign node9068 = (inp[1]) ? 4'b1101 : 4'b1100;
												assign node9071 = (inp[0]) ? node9095 : node9072;
													assign node9072 = (inp[11]) ? node9080 : node9073;
														assign node9073 = (inp[9]) ? node9077 : node9074;
															assign node9074 = (inp[10]) ? 4'b1000 : 4'b1001;
															assign node9077 = (inp[10]) ? 4'b1001 : 4'b1000;
														assign node9080 = (inp[1]) ? node9088 : node9081;
															assign node9081 = (inp[9]) ? node9085 : node9082;
																assign node9082 = (inp[10]) ? 4'b1001 : 4'b1000;
																assign node9085 = (inp[10]) ? 4'b1000 : 4'b1001;
															assign node9088 = (inp[9]) ? node9092 : node9089;
																assign node9089 = (inp[10]) ? 4'b1000 : 4'b1001;
																assign node9092 = (inp[10]) ? 4'b1001 : 4'b1000;
													assign node9095 = (inp[9]) ? node9103 : node9096;
														assign node9096 = (inp[10]) ? node9098 : 4'b1001;
															assign node9098 = (inp[11]) ? 4'b1000 : node9099;
																assign node9099 = (inp[1]) ? 4'b1001 : 4'b1000;
														assign node9103 = (inp[10]) ? node9109 : node9104;
															assign node9104 = (inp[1]) ? node9106 : 4'b1000;
																assign node9106 = (inp[11]) ? 4'b1000 : 4'b1001;
															assign node9109 = (inp[1]) ? node9111 : 4'b1001;
																assign node9111 = (inp[11]) ? 4'b1001 : 4'b1000;
											assign node9114 = (inp[11]) ? node9146 : node9115;
												assign node9115 = (inp[2]) ? node9131 : node9116;
													assign node9116 = (inp[1]) ? node9124 : node9117;
														assign node9117 = (inp[10]) ? node9121 : node9118;
															assign node9118 = (inp[9]) ? 4'b1011 : 4'b1010;
															assign node9121 = (inp[9]) ? 4'b1010 : 4'b1011;
														assign node9124 = (inp[0]) ? 4'b1111 : node9125;
															assign node9125 = (inp[9]) ? 4'b1110 : node9126;
																assign node9126 = (inp[10]) ? 4'b1111 : 4'b1110;
													assign node9131 = (inp[1]) ? node9139 : node9132;
														assign node9132 = (inp[9]) ? node9136 : node9133;
															assign node9133 = (inp[10]) ? 4'b1110 : 4'b1111;
															assign node9136 = (inp[10]) ? 4'b1111 : 4'b1110;
														assign node9139 = (inp[10]) ? node9143 : node9140;
															assign node9140 = (inp[9]) ? 4'b1010 : 4'b1011;
															assign node9143 = (inp[9]) ? 4'b1011 : 4'b1010;
												assign node9146 = (inp[1]) ? node9170 : node9147;
													assign node9147 = (inp[2]) ? node9157 : node9148;
														assign node9148 = (inp[0]) ? node9150 : 4'b1011;
															assign node9150 = (inp[10]) ? node9154 : node9151;
																assign node9151 = (inp[9]) ? 4'b1011 : 4'b1010;
																assign node9154 = (inp[9]) ? 4'b1010 : 4'b1011;
														assign node9157 = (inp[0]) ? node9165 : node9158;
															assign node9158 = (inp[9]) ? node9162 : node9159;
																assign node9159 = (inp[10]) ? 4'b1111 : 4'b1110;
																assign node9162 = (inp[10]) ? 4'b1110 : 4'b1111;
															assign node9165 = (inp[10]) ? node9167 : 4'b1111;
																assign node9167 = (inp[9]) ? 4'b1111 : 4'b1110;
													assign node9170 = (inp[2]) ? node9178 : node9171;
														assign node9171 = (inp[10]) ? node9175 : node9172;
															assign node9172 = (inp[9]) ? 4'b1111 : 4'b1110;
															assign node9175 = (inp[9]) ? 4'b1110 : 4'b1111;
														assign node9178 = (inp[9]) ? node9184 : node9179;
															assign node9179 = (inp[10]) ? 4'b1011 : node9180;
																assign node9180 = (inp[0]) ? 4'b1011 : 4'b1010;
															assign node9184 = (inp[10]) ? node9188 : node9185;
																assign node9185 = (inp[0]) ? 4'b1010 : 4'b1011;
																assign node9188 = (inp[0]) ? 4'b1011 : 4'b1010;
								assign node9191 = (inp[12]) ? node9569 : node9192;
									assign node9192 = (inp[15]) ? node9374 : node9193;
										assign node9193 = (inp[4]) ? node9283 : node9194;
											assign node9194 = (inp[2]) ? node9232 : node9195;
												assign node9195 = (inp[11]) ? node9211 : node9196;
													assign node9196 = (inp[10]) ? node9202 : node9197;
														assign node9197 = (inp[9]) ? 4'b1011 : node9198;
															assign node9198 = (inp[1]) ? 4'b1010 : 4'b1011;
														assign node9202 = (inp[9]) ? node9208 : node9203;
															assign node9203 = (inp[1]) ? 4'b1011 : node9204;
																assign node9204 = (inp[0]) ? 4'b1010 : 4'b1011;
															assign node9208 = (inp[0]) ? 4'b1011 : 4'b1010;
													assign node9211 = (inp[10]) ? node9223 : node9212;
														assign node9212 = (inp[9]) ? node9218 : node9213;
															assign node9213 = (inp[1]) ? node9215 : 4'b1010;
																assign node9215 = (inp[0]) ? 4'b1010 : 4'b1011;
															assign node9218 = (inp[0]) ? 4'b1011 : node9219;
																assign node9219 = (inp[1]) ? 4'b1010 : 4'b1011;
														assign node9223 = (inp[9]) ? node9227 : node9224;
															assign node9224 = (inp[0]) ? 4'b1011 : 4'b1010;
															assign node9227 = (inp[1]) ? node9229 : 4'b1010;
																assign node9229 = (inp[0]) ? 4'b1010 : 4'b1011;
												assign node9232 = (inp[0]) ? node9260 : node9233;
													assign node9233 = (inp[11]) ? node9245 : node9234;
														assign node9234 = (inp[1]) ? node9240 : node9235;
															assign node9235 = (inp[10]) ? node9237 : 4'b1110;
																assign node9237 = (inp[9]) ? 4'b1110 : 4'b1111;
															assign node9240 = (inp[9]) ? node9242 : 4'b1110;
																assign node9242 = (inp[10]) ? 4'b1110 : 4'b1111;
														assign node9245 = (inp[9]) ? node9253 : node9246;
															assign node9246 = (inp[10]) ? node9250 : node9247;
																assign node9247 = (inp[1]) ? 4'b1111 : 4'b1110;
																assign node9250 = (inp[1]) ? 4'b1110 : 4'b1111;
															assign node9253 = (inp[1]) ? node9257 : node9254;
																assign node9254 = (inp[10]) ? 4'b1110 : 4'b1111;
																assign node9257 = (inp[10]) ? 4'b1111 : 4'b1110;
													assign node9260 = (inp[10]) ? node9272 : node9261;
														assign node9261 = (inp[9]) ? node9267 : node9262;
															assign node9262 = (inp[1]) ? 4'b1110 : node9263;
																assign node9263 = (inp[11]) ? 4'b1110 : 4'b1111;
															assign node9267 = (inp[11]) ? 4'b1111 : node9268;
																assign node9268 = (inp[1]) ? 4'b1111 : 4'b1110;
														assign node9272 = (inp[9]) ? node9278 : node9273;
															assign node9273 = (inp[1]) ? 4'b1111 : node9274;
																assign node9274 = (inp[11]) ? 4'b1111 : 4'b1110;
															assign node9278 = (inp[1]) ? 4'b1110 : node9279;
																assign node9279 = (inp[11]) ? 4'b1110 : 4'b1111;
											assign node9283 = (inp[11]) ? node9321 : node9284;
												assign node9284 = (inp[9]) ? node9304 : node9285;
													assign node9285 = (inp[10]) ? node9295 : node9286;
														assign node9286 = (inp[2]) ? node9292 : node9287;
															assign node9287 = (inp[1]) ? 4'b1000 : node9288;
																assign node9288 = (inp[0]) ? 4'b1101 : 4'b1100;
															assign node9292 = (inp[1]) ? 4'b1101 : 4'b1001;
														assign node9295 = (inp[2]) ? node9301 : node9296;
															assign node9296 = (inp[1]) ? 4'b1001 : node9297;
																assign node9297 = (inp[0]) ? 4'b1100 : 4'b1101;
															assign node9301 = (inp[1]) ? 4'b1100 : 4'b1000;
													assign node9304 = (inp[10]) ? node9312 : node9305;
														assign node9305 = (inp[2]) ? node9309 : node9306;
															assign node9306 = (inp[1]) ? 4'b1001 : 4'b1100;
															assign node9309 = (inp[1]) ? 4'b1100 : 4'b1000;
														assign node9312 = (inp[2]) ? node9318 : node9313;
															assign node9313 = (inp[1]) ? 4'b1000 : node9314;
																assign node9314 = (inp[0]) ? 4'b1101 : 4'b1100;
															assign node9318 = (inp[1]) ? 4'b1101 : 4'b1001;
												assign node9321 = (inp[0]) ? node9345 : node9322;
													assign node9322 = (inp[1]) ? node9332 : node9323;
														assign node9323 = (inp[2]) ? 4'b1000 : node9324;
															assign node9324 = (inp[10]) ? node9328 : node9325;
																assign node9325 = (inp[9]) ? 4'b1101 : 4'b1100;
																assign node9328 = (inp[9]) ? 4'b1100 : 4'b1101;
														assign node9332 = (inp[2]) ? node9338 : node9333;
															assign node9333 = (inp[10]) ? node9335 : 4'b1000;
																assign node9335 = (inp[9]) ? 4'b1001 : 4'b1000;
															assign node9338 = (inp[10]) ? node9342 : node9339;
																assign node9339 = (inp[9]) ? 4'b1101 : 4'b1100;
																assign node9342 = (inp[9]) ? 4'b1100 : 4'b1101;
													assign node9345 = (inp[1]) ? node9361 : node9346;
														assign node9346 = (inp[2]) ? node9354 : node9347;
															assign node9347 = (inp[10]) ? node9351 : node9348;
																assign node9348 = (inp[9]) ? 4'b1101 : 4'b1100;
																assign node9351 = (inp[9]) ? 4'b1100 : 4'b1101;
															assign node9354 = (inp[10]) ? node9358 : node9355;
																assign node9355 = (inp[9]) ? 4'b1000 : 4'b1001;
																assign node9358 = (inp[9]) ? 4'b1001 : 4'b1000;
														assign node9361 = (inp[2]) ? node9367 : node9362;
															assign node9362 = (inp[10]) ? 4'b1000 : node9363;
																assign node9363 = (inp[9]) ? 4'b1001 : 4'b1000;
															assign node9367 = (inp[10]) ? node9371 : node9368;
																assign node9368 = (inp[9]) ? 4'b1100 : 4'b1101;
																assign node9371 = (inp[9]) ? 4'b1101 : 4'b1100;
										assign node9374 = (inp[9]) ? node9470 : node9375;
											assign node9375 = (inp[2]) ? node9419 : node9376;
												assign node9376 = (inp[4]) ? node9396 : node9377;
													assign node9377 = (inp[1]) ? node9389 : node9378;
														assign node9378 = (inp[10]) ? node9384 : node9379;
															assign node9379 = (inp[0]) ? node9381 : 4'b1110;
																assign node9381 = (inp[11]) ? 4'b1110 : 4'b1111;
															assign node9384 = (inp[11]) ? 4'b1111 : node9385;
																assign node9385 = (inp[0]) ? 4'b1110 : 4'b1111;
														assign node9389 = (inp[10]) ? node9391 : 4'b1111;
															assign node9391 = (inp[11]) ? 4'b1110 : node9392;
																assign node9392 = (inp[0]) ? 4'b1111 : 4'b1110;
													assign node9396 = (inp[10]) ? node9408 : node9397;
														assign node9397 = (inp[1]) ? node9403 : node9398;
															assign node9398 = (inp[11]) ? node9400 : 4'b1010;
																assign node9400 = (inp[0]) ? 4'b1010 : 4'b1011;
															assign node9403 = (inp[11]) ? node9405 : 4'b1011;
																assign node9405 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node9408 = (inp[1]) ? node9414 : node9409;
															assign node9409 = (inp[0]) ? 4'b1011 : node9410;
																assign node9410 = (inp[11]) ? 4'b1010 : 4'b1011;
															assign node9414 = (inp[11]) ? node9416 : 4'b1010;
																assign node9416 = (inp[0]) ? 4'b1010 : 4'b1011;
												assign node9419 = (inp[4]) ? node9441 : node9420;
													assign node9420 = (inp[0]) ? node9434 : node9421;
														assign node9421 = (inp[10]) ? node9427 : node9422;
															assign node9422 = (inp[11]) ? node9424 : 4'b1010;
																assign node9424 = (inp[1]) ? 4'b1010 : 4'b1011;
															assign node9427 = (inp[11]) ? node9431 : node9428;
																assign node9428 = (inp[1]) ? 4'b1010 : 4'b1011;
																assign node9431 = (inp[1]) ? 4'b1011 : 4'b1010;
														assign node9434 = (inp[10]) ? node9438 : node9435;
															assign node9435 = (inp[1]) ? 4'b1011 : 4'b1010;
															assign node9438 = (inp[1]) ? 4'b1010 : 4'b1011;
													assign node9441 = (inp[11]) ? node9457 : node9442;
														assign node9442 = (inp[0]) ? node9450 : node9443;
															assign node9443 = (inp[1]) ? node9447 : node9444;
																assign node9444 = (inp[10]) ? 4'b1110 : 4'b1111;
																assign node9447 = (inp[10]) ? 4'b1111 : 4'b1110;
															assign node9450 = (inp[1]) ? node9454 : node9451;
																assign node9451 = (inp[10]) ? 4'b1110 : 4'b1111;
																assign node9454 = (inp[10]) ? 4'b1111 : 4'b1110;
														assign node9457 = (inp[1]) ? node9463 : node9458;
															assign node9458 = (inp[10]) ? node9460 : 4'b1111;
																assign node9460 = (inp[0]) ? 4'b1110 : 4'b1111;
															assign node9463 = (inp[10]) ? node9467 : node9464;
																assign node9464 = (inp[0]) ? 4'b1110 : 4'b1111;
																assign node9467 = (inp[0]) ? 4'b1111 : 4'b1110;
											assign node9470 = (inp[0]) ? node9530 : node9471;
												assign node9471 = (inp[11]) ? node9501 : node9472;
													assign node9472 = (inp[2]) ? node9488 : node9473;
														assign node9473 = (inp[4]) ? node9481 : node9474;
															assign node9474 = (inp[1]) ? node9478 : node9475;
																assign node9475 = (inp[10]) ? 4'b1110 : 4'b1111;
																assign node9478 = (inp[10]) ? 4'b1111 : 4'b1110;
															assign node9481 = (inp[10]) ? node9485 : node9482;
																assign node9482 = (inp[1]) ? 4'b1010 : 4'b1011;
																assign node9485 = (inp[1]) ? 4'b1011 : 4'b1010;
														assign node9488 = (inp[4]) ? node9494 : node9489;
															assign node9489 = (inp[1]) ? node9491 : 4'b1011;
																assign node9491 = (inp[10]) ? 4'b1011 : 4'b1010;
															assign node9494 = (inp[1]) ? node9498 : node9495;
																assign node9495 = (inp[10]) ? 4'b1111 : 4'b1110;
																assign node9498 = (inp[10]) ? 4'b1110 : 4'b1111;
													assign node9501 = (inp[10]) ? node9517 : node9502;
														assign node9502 = (inp[1]) ? node9510 : node9503;
															assign node9503 = (inp[4]) ? node9507 : node9504;
																assign node9504 = (inp[2]) ? 4'b1010 : 4'b1111;
																assign node9507 = (inp[2]) ? 4'b1111 : 4'b1010;
															assign node9510 = (inp[4]) ? node9514 : node9511;
																assign node9511 = (inp[2]) ? 4'b1011 : 4'b1110;
																assign node9514 = (inp[2]) ? 4'b1110 : 4'b1011;
														assign node9517 = (inp[2]) ? node9525 : node9518;
															assign node9518 = (inp[4]) ? node9522 : node9519;
																assign node9519 = (inp[1]) ? 4'b1111 : 4'b1110;
																assign node9522 = (inp[1]) ? 4'b1010 : 4'b1011;
															assign node9525 = (inp[4]) ? 4'b1110 : node9526;
																assign node9526 = (inp[1]) ? 4'b1010 : 4'b1011;
												assign node9530 = (inp[4]) ? node9554 : node9531;
													assign node9531 = (inp[2]) ? node9547 : node9532;
														assign node9532 = (inp[11]) ? node9540 : node9533;
															assign node9533 = (inp[10]) ? node9537 : node9534;
																assign node9534 = (inp[1]) ? 4'b1111 : 4'b1110;
																assign node9537 = (inp[1]) ? 4'b1110 : 4'b1111;
															assign node9540 = (inp[10]) ? node9544 : node9541;
																assign node9541 = (inp[1]) ? 4'b1110 : 4'b1111;
																assign node9544 = (inp[1]) ? 4'b1111 : 4'b1110;
														assign node9547 = (inp[1]) ? node9551 : node9548;
															assign node9548 = (inp[10]) ? 4'b1010 : 4'b1011;
															assign node9551 = (inp[10]) ? 4'b1011 : 4'b1010;
													assign node9554 = (inp[2]) ? node9562 : node9555;
														assign node9555 = (inp[10]) ? node9559 : node9556;
															assign node9556 = (inp[1]) ? 4'b1010 : 4'b1011;
															assign node9559 = (inp[1]) ? 4'b1011 : 4'b1010;
														assign node9562 = (inp[1]) ? node9566 : node9563;
															assign node9563 = (inp[10]) ? 4'b1111 : 4'b1110;
															assign node9566 = (inp[10]) ? 4'b1110 : 4'b1111;
									assign node9569 = (inp[4]) ? node9739 : node9570;
										assign node9570 = (inp[0]) ? node9648 : node9571;
											assign node9571 = (inp[9]) ? node9609 : node9572;
												assign node9572 = (inp[10]) ? node9590 : node9573;
													assign node9573 = (inp[15]) ? node9583 : node9574;
														assign node9574 = (inp[1]) ? node9580 : node9575;
															assign node9575 = (inp[2]) ? 4'b1001 : node9576;
																assign node9576 = (inp[11]) ? 4'b1101 : 4'b1100;
															assign node9580 = (inp[2]) ? 4'b1100 : 4'b1000;
														assign node9583 = (inp[2]) ? node9587 : node9584;
															assign node9584 = (inp[1]) ? 4'b1101 : 4'b1001;
															assign node9587 = (inp[1]) ? 4'b1001 : 4'b1101;
													assign node9590 = (inp[2]) ? node9602 : node9591;
														assign node9591 = (inp[11]) ? node9597 : node9592;
															assign node9592 = (inp[15]) ? 4'b1101 : node9593;
																assign node9593 = (inp[1]) ? 4'b1001 : 4'b1101;
															assign node9597 = (inp[15]) ? 4'b1100 : node9598;
																assign node9598 = (inp[1]) ? 4'b1001 : 4'b1100;
														assign node9602 = (inp[15]) ? node9606 : node9603;
															assign node9603 = (inp[1]) ? 4'b1101 : 4'b1000;
															assign node9606 = (inp[1]) ? 4'b1000 : 4'b1100;
												assign node9609 = (inp[10]) ? node9633 : node9610;
													assign node9610 = (inp[15]) ? node9620 : node9611;
														assign node9611 = (inp[1]) ? node9617 : node9612;
															assign node9612 = (inp[2]) ? 4'b1000 : node9613;
																assign node9613 = (inp[11]) ? 4'b1100 : 4'b1101;
															assign node9617 = (inp[2]) ? 4'b1101 : 4'b1001;
														assign node9620 = (inp[11]) ? node9626 : node9621;
															assign node9621 = (inp[2]) ? node9623 : 4'b1101;
																assign node9623 = (inp[1]) ? 4'b1000 : 4'b1100;
															assign node9626 = (inp[1]) ? node9630 : node9627;
																assign node9627 = (inp[2]) ? 4'b1100 : 4'b1000;
																assign node9630 = (inp[2]) ? 4'b1000 : 4'b1100;
													assign node9633 = (inp[1]) ? node9641 : node9634;
														assign node9634 = (inp[15]) ? node9638 : node9635;
															assign node9635 = (inp[2]) ? 4'b1001 : 4'b1100;
															assign node9638 = (inp[2]) ? 4'b1101 : 4'b1001;
														assign node9641 = (inp[15]) ? node9645 : node9642;
															assign node9642 = (inp[2]) ? 4'b1100 : 4'b1000;
															assign node9645 = (inp[2]) ? 4'b1001 : 4'b1100;
											assign node9648 = (inp[15]) ? node9690 : node9649;
												assign node9649 = (inp[10]) ? node9665 : node9650;
													assign node9650 = (inp[1]) ? node9656 : node9651;
														assign node9651 = (inp[2]) ? 4'b1000 : node9652;
															assign node9652 = (inp[9]) ? 4'b1101 : 4'b1100;
														assign node9656 = (inp[2]) ? node9658 : 4'b1001;
															assign node9658 = (inp[9]) ? node9662 : node9659;
																assign node9659 = (inp[11]) ? 4'b1100 : 4'b1101;
																assign node9662 = (inp[11]) ? 4'b1101 : 4'b1100;
													assign node9665 = (inp[9]) ? node9679 : node9666;
														assign node9666 = (inp[11]) ? node9672 : node9667;
															assign node9667 = (inp[1]) ? node9669 : 4'b1001;
																assign node9669 = (inp[2]) ? 4'b1100 : 4'b1000;
															assign node9672 = (inp[2]) ? node9676 : node9673;
																assign node9673 = (inp[1]) ? 4'b1001 : 4'b1101;
																assign node9676 = (inp[1]) ? 4'b1101 : 4'b1000;
														assign node9679 = (inp[2]) ? node9683 : node9680;
															assign node9680 = (inp[1]) ? 4'b1000 : 4'b1100;
															assign node9683 = (inp[1]) ? node9687 : node9684;
																assign node9684 = (inp[11]) ? 4'b1001 : 4'b1000;
																assign node9687 = (inp[11]) ? 4'b1100 : 4'b1101;
												assign node9690 = (inp[10]) ? node9716 : node9691;
													assign node9691 = (inp[1]) ? node9707 : node9692;
														assign node9692 = (inp[2]) ? node9700 : node9693;
															assign node9693 = (inp[9]) ? node9697 : node9694;
																assign node9694 = (inp[11]) ? 4'b1001 : 4'b1000;
																assign node9697 = (inp[11]) ? 4'b1000 : 4'b1001;
															assign node9700 = (inp[9]) ? node9704 : node9701;
																assign node9701 = (inp[11]) ? 4'b1101 : 4'b1100;
																assign node9704 = (inp[11]) ? 4'b1100 : 4'b1101;
														assign node9707 = (inp[2]) ? node9709 : 4'b1100;
															assign node9709 = (inp[9]) ? node9713 : node9710;
																assign node9710 = (inp[11]) ? 4'b1001 : 4'b1000;
																assign node9713 = (inp[11]) ? 4'b1000 : 4'b1001;
													assign node9716 = (inp[11]) ? node9726 : node9717;
														assign node9717 = (inp[9]) ? 4'b1100 : node9718;
															assign node9718 = (inp[1]) ? node9722 : node9719;
																assign node9719 = (inp[2]) ? 4'b1101 : 4'b1001;
																assign node9722 = (inp[2]) ? 4'b1001 : 4'b1101;
														assign node9726 = (inp[9]) ? node9734 : node9727;
															assign node9727 = (inp[2]) ? node9731 : node9728;
																assign node9728 = (inp[1]) ? 4'b1101 : 4'b1000;
																assign node9731 = (inp[1]) ? 4'b1000 : 4'b1100;
															assign node9734 = (inp[2]) ? node9736 : 4'b1100;
																assign node9736 = (inp[1]) ? 4'b1001 : 4'b1101;
										assign node9739 = (inp[15]) ? node9851 : node9740;
											assign node9740 = (inp[0]) ? node9794 : node9741;
												assign node9741 = (inp[11]) ? node9763 : node9742;
													assign node9742 = (inp[2]) ? node9756 : node9743;
														assign node9743 = (inp[1]) ? node9749 : node9744;
															assign node9744 = (inp[9]) ? node9746 : 4'b1011;
																assign node9746 = (inp[10]) ? 4'b1011 : 4'b1010;
															assign node9749 = (inp[9]) ? node9753 : node9750;
																assign node9750 = (inp[10]) ? 4'b1111 : 4'b1110;
																assign node9753 = (inp[10]) ? 4'b1110 : 4'b1111;
														assign node9756 = (inp[1]) ? node9758 : 4'b1111;
															assign node9758 = (inp[10]) ? node9760 : 4'b1011;
																assign node9760 = (inp[9]) ? 4'b1011 : 4'b1010;
													assign node9763 = (inp[1]) ? node9779 : node9764;
														assign node9764 = (inp[2]) ? node9772 : node9765;
															assign node9765 = (inp[9]) ? node9769 : node9766;
																assign node9766 = (inp[10]) ? 4'b1010 : 4'b1011;
																assign node9769 = (inp[10]) ? 4'b1011 : 4'b1010;
															assign node9772 = (inp[10]) ? node9776 : node9773;
																assign node9773 = (inp[9]) ? 4'b1111 : 4'b1110;
																assign node9776 = (inp[9]) ? 4'b1110 : 4'b1111;
														assign node9779 = (inp[2]) ? node9787 : node9780;
															assign node9780 = (inp[9]) ? node9784 : node9781;
																assign node9781 = (inp[10]) ? 4'b1111 : 4'b1110;
																assign node9784 = (inp[10]) ? 4'b1110 : 4'b1111;
															assign node9787 = (inp[9]) ? node9791 : node9788;
																assign node9788 = (inp[10]) ? 4'b1011 : 4'b1010;
																assign node9791 = (inp[10]) ? 4'b1010 : 4'b1011;
												assign node9794 = (inp[11]) ? node9820 : node9795;
													assign node9795 = (inp[9]) ? node9807 : node9796;
														assign node9796 = (inp[10]) ? node9802 : node9797;
															assign node9797 = (inp[2]) ? 4'b1111 : node9798;
																assign node9798 = (inp[1]) ? 4'b1111 : 4'b1010;
															assign node9802 = (inp[2]) ? node9804 : 4'b1110;
																assign node9804 = (inp[1]) ? 4'b1010 : 4'b1110;
														assign node9807 = (inp[10]) ? node9815 : node9808;
															assign node9808 = (inp[2]) ? node9812 : node9809;
																assign node9809 = (inp[1]) ? 4'b1110 : 4'b1011;
																assign node9812 = (inp[1]) ? 4'b1010 : 4'b1110;
															assign node9815 = (inp[2]) ? node9817 : 4'b1111;
																assign node9817 = (inp[1]) ? 4'b1011 : 4'b1111;
													assign node9820 = (inp[1]) ? node9836 : node9821;
														assign node9821 = (inp[2]) ? node9829 : node9822;
															assign node9822 = (inp[10]) ? node9826 : node9823;
																assign node9823 = (inp[9]) ? 4'b1010 : 4'b1011;
																assign node9826 = (inp[9]) ? 4'b1011 : 4'b1010;
															assign node9829 = (inp[9]) ? node9833 : node9830;
																assign node9830 = (inp[10]) ? 4'b1111 : 4'b1110;
																assign node9833 = (inp[10]) ? 4'b1110 : 4'b1111;
														assign node9836 = (inp[2]) ? node9844 : node9837;
															assign node9837 = (inp[9]) ? node9841 : node9838;
																assign node9838 = (inp[10]) ? 4'b1111 : 4'b1110;
																assign node9841 = (inp[10]) ? 4'b1110 : 4'b1111;
															assign node9844 = (inp[9]) ? node9848 : node9845;
																assign node9845 = (inp[10]) ? 4'b1010 : 4'b1011;
																assign node9848 = (inp[10]) ? 4'b1011 : 4'b1010;
											assign node9851 = (inp[10]) ? node9901 : node9852;
												assign node9852 = (inp[11]) ? node9878 : node9853;
													assign node9853 = (inp[0]) ? node9863 : node9854;
														assign node9854 = (inp[2]) ? node9860 : node9855;
															assign node9855 = (inp[9]) ? node9857 : 4'b1001;
																assign node9857 = (inp[1]) ? 4'b1100 : 4'b1000;
															assign node9860 = (inp[9]) ? 4'b1001 : 4'b1000;
														assign node9863 = (inp[9]) ? node9871 : node9864;
															assign node9864 = (inp[1]) ? node9868 : node9865;
																assign node9865 = (inp[2]) ? 4'b1100 : 4'b1001;
																assign node9868 = (inp[2]) ? 4'b1000 : 4'b1100;
															assign node9871 = (inp[1]) ? node9875 : node9872;
																assign node9872 = (inp[2]) ? 4'b1101 : 4'b1000;
																assign node9875 = (inp[2]) ? 4'b1001 : 4'b1101;
													assign node9878 = (inp[9]) ? node9890 : node9879;
														assign node9879 = (inp[1]) ? node9885 : node9880;
															assign node9880 = (inp[2]) ? node9882 : 4'b1000;
																assign node9882 = (inp[0]) ? 4'b1100 : 4'b1101;
															assign node9885 = (inp[2]) ? node9887 : 4'b1101;
																assign node9887 = (inp[0]) ? 4'b1000 : 4'b1001;
														assign node9890 = (inp[1]) ? node9896 : node9891;
															assign node9891 = (inp[2]) ? 4'b1100 : node9892;
																assign node9892 = (inp[0]) ? 4'b1000 : 4'b1001;
															assign node9896 = (inp[2]) ? node9898 : 4'b1100;
																assign node9898 = (inp[0]) ? 4'b1001 : 4'b1000;
												assign node9901 = (inp[0]) ? node9921 : node9902;
													assign node9902 = (inp[2]) ? node9908 : node9903;
														assign node9903 = (inp[1]) ? node9905 : 4'b1001;
															assign node9905 = (inp[9]) ? 4'b1101 : 4'b1100;
														assign node9908 = (inp[1]) ? node9916 : node9909;
															assign node9909 = (inp[11]) ? node9913 : node9910;
																assign node9910 = (inp[9]) ? 4'b1100 : 4'b1101;
																assign node9913 = (inp[9]) ? 4'b1101 : 4'b1100;
															assign node9916 = (inp[9]) ? node9918 : 4'b1001;
																assign node9918 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node9921 = (inp[9]) ? node9931 : node9922;
														assign node9922 = (inp[2]) ? node9928 : node9923;
															assign node9923 = (inp[1]) ? node9925 : 4'b1000;
																assign node9925 = (inp[11]) ? 4'b1100 : 4'b1101;
															assign node9928 = (inp[1]) ? 4'b1001 : 4'b1101;
														assign node9931 = (inp[2]) ? node9937 : node9932;
															assign node9932 = (inp[1]) ? node9934 : 4'b1001;
																assign node9934 = (inp[11]) ? 4'b1101 : 4'b1100;
															assign node9937 = (inp[1]) ? 4'b1000 : 4'b1100;
							assign node9940 = (inp[12]) ? node10412 : node9941;
								assign node9941 = (inp[15]) ? node10219 : node9942;
									assign node9942 = (inp[7]) ? node10096 : node9943;
										assign node9943 = (inp[1]) ? node10021 : node9944;
											assign node9944 = (inp[2]) ? node9976 : node9945;
												assign node9945 = (inp[10]) ? node9961 : node9946;
													assign node9946 = (inp[0]) ? node9954 : node9947;
														assign node9947 = (inp[11]) ? node9951 : node9948;
															assign node9948 = (inp[9]) ? 4'b1001 : 4'b1000;
															assign node9951 = (inp[9]) ? 4'b1000 : 4'b1001;
														assign node9954 = (inp[9]) ? node9958 : node9955;
															assign node9955 = (inp[11]) ? 4'b1000 : 4'b1001;
															assign node9958 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node9961 = (inp[9]) ? node9969 : node9962;
														assign node9962 = (inp[11]) ? node9966 : node9963;
															assign node9963 = (inp[0]) ? 4'b1001 : 4'b1000;
															assign node9966 = (inp[0]) ? 4'b1000 : 4'b1001;
														assign node9969 = (inp[11]) ? node9973 : node9970;
															assign node9970 = (inp[0]) ? 4'b1000 : 4'b1001;
															assign node9973 = (inp[0]) ? 4'b1001 : 4'b1000;
												assign node9976 = (inp[0]) ? node10000 : node9977;
													assign node9977 = (inp[10]) ? node9991 : node9978;
														assign node9978 = (inp[11]) ? node9986 : node9979;
															assign node9979 = (inp[4]) ? node9983 : node9980;
																assign node9980 = (inp[9]) ? 4'b1001 : 4'b1000;
																assign node9983 = (inp[9]) ? 4'b1000 : 4'b1001;
															assign node9986 = (inp[9]) ? 4'b1000 : node9987;
																assign node9987 = (inp[4]) ? 4'b1000 : 4'b1001;
														assign node9991 = (inp[9]) ? node9993 : 4'b1001;
															assign node9993 = (inp[11]) ? node9997 : node9994;
																assign node9994 = (inp[4]) ? 4'b1000 : 4'b1001;
																assign node9997 = (inp[4]) ? 4'b1001 : 4'b1000;
													assign node10000 = (inp[10]) ? node10008 : node10001;
														assign node10001 = (inp[11]) ? node10003 : 4'b1001;
															assign node10003 = (inp[4]) ? 4'b1001 : node10004;
																assign node10004 = (inp[9]) ? 4'b1000 : 4'b1001;
														assign node10008 = (inp[9]) ? node10016 : node10009;
															assign node10009 = (inp[11]) ? node10013 : node10010;
																assign node10010 = (inp[4]) ? 4'b1001 : 4'b1000;
																assign node10013 = (inp[4]) ? 4'b1000 : 4'b1001;
															assign node10016 = (inp[11]) ? 4'b1001 : node10017;
																assign node10017 = (inp[4]) ? 4'b1000 : 4'b1001;
											assign node10021 = (inp[4]) ? node10067 : node10022;
												assign node10022 = (inp[10]) ? node10046 : node10023;
													assign node10023 = (inp[9]) ? node10035 : node10024;
														assign node10024 = (inp[11]) ? node10030 : node10025;
															assign node10025 = (inp[0]) ? node10027 : 4'b1100;
																assign node10027 = (inp[2]) ? 4'b1100 : 4'b1101;
															assign node10030 = (inp[2]) ? 4'b1101 : node10031;
																assign node10031 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node10035 = (inp[11]) ? node10041 : node10036;
															assign node10036 = (inp[0]) ? node10038 : 4'b1101;
																assign node10038 = (inp[2]) ? 4'b1101 : 4'b1100;
															assign node10041 = (inp[0]) ? node10043 : 4'b1100;
																assign node10043 = (inp[2]) ? 4'b1100 : 4'b1101;
													assign node10046 = (inp[0]) ? node10056 : node10047;
														assign node10047 = (inp[2]) ? 4'b1100 : node10048;
															assign node10048 = (inp[11]) ? node10052 : node10049;
																assign node10049 = (inp[9]) ? 4'b1101 : 4'b1100;
																assign node10052 = (inp[9]) ? 4'b1100 : 4'b1101;
														assign node10056 = (inp[9]) ? node10062 : node10057;
															assign node10057 = (inp[2]) ? node10059 : 4'b1100;
																assign node10059 = (inp[11]) ? 4'b1101 : 4'b1100;
															assign node10062 = (inp[11]) ? 4'b1101 : node10063;
																assign node10063 = (inp[2]) ? 4'b1101 : 4'b1100;
												assign node10067 = (inp[2]) ? node10075 : node10068;
													assign node10068 = (inp[11]) ? node10072 : node10069;
														assign node10069 = (inp[9]) ? 4'b1001 : 4'b1000;
														assign node10072 = (inp[9]) ? 4'b1000 : 4'b1001;
													assign node10075 = (inp[9]) ? node10089 : node10076;
														assign node10076 = (inp[10]) ? node10082 : node10077;
															assign node10077 = (inp[11]) ? 4'b1000 : node10078;
																assign node10078 = (inp[0]) ? 4'b1001 : 4'b1000;
															assign node10082 = (inp[0]) ? node10086 : node10083;
																assign node10083 = (inp[11]) ? 4'b1001 : 4'b1000;
																assign node10086 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node10089 = (inp[0]) ? node10093 : node10090;
															assign node10090 = (inp[11]) ? 4'b1000 : 4'b1001;
															assign node10093 = (inp[11]) ? 4'b1001 : 4'b1000;
										assign node10096 = (inp[4]) ? node10146 : node10097;
											assign node10097 = (inp[9]) ? node10121 : node10098;
												assign node10098 = (inp[11]) ? node10110 : node10099;
													assign node10099 = (inp[0]) ? node10105 : node10100;
														assign node10100 = (inp[2]) ? node10102 : 4'b1010;
															assign node10102 = (inp[1]) ? 4'b1011 : 4'b1010;
														assign node10105 = (inp[2]) ? 4'b1010 : node10106;
															assign node10106 = (inp[1]) ? 4'b1010 : 4'b1011;
													assign node10110 = (inp[2]) ? node10116 : node10111;
														assign node10111 = (inp[1]) ? 4'b1011 : node10112;
															assign node10112 = (inp[0]) ? 4'b1010 : 4'b1011;
														assign node10116 = (inp[1]) ? node10118 : 4'b1011;
															assign node10118 = (inp[0]) ? 4'b1011 : 4'b1010;
												assign node10121 = (inp[11]) ? node10133 : node10122;
													assign node10122 = (inp[2]) ? node10128 : node10123;
														assign node10123 = (inp[1]) ? 4'b1011 : node10124;
															assign node10124 = (inp[0]) ? 4'b1010 : 4'b1011;
														assign node10128 = (inp[0]) ? 4'b1011 : node10129;
															assign node10129 = (inp[1]) ? 4'b1010 : 4'b1011;
													assign node10133 = (inp[10]) ? 4'b1010 : node10134;
														assign node10134 = (inp[2]) ? node10140 : node10135;
															assign node10135 = (inp[1]) ? 4'b1010 : node10136;
																assign node10136 = (inp[0]) ? 4'b1011 : 4'b1010;
															assign node10140 = (inp[1]) ? node10142 : 4'b1010;
																assign node10142 = (inp[0]) ? 4'b1010 : 4'b1011;
											assign node10146 = (inp[1]) ? node10170 : node10147;
												assign node10147 = (inp[0]) ? node10163 : node10148;
													assign node10148 = (inp[2]) ? node10156 : node10149;
														assign node10149 = (inp[9]) ? node10153 : node10150;
															assign node10150 = (inp[11]) ? 4'b1111 : 4'b1110;
															assign node10153 = (inp[11]) ? 4'b1110 : 4'b1111;
														assign node10156 = (inp[9]) ? node10160 : node10157;
															assign node10157 = (inp[11]) ? 4'b1110 : 4'b1111;
															assign node10160 = (inp[11]) ? 4'b1111 : 4'b1110;
													assign node10163 = (inp[9]) ? node10167 : node10164;
														assign node10164 = (inp[11]) ? 4'b1110 : 4'b1111;
														assign node10167 = (inp[11]) ? 4'b1111 : 4'b1110;
												assign node10170 = (inp[2]) ? node10196 : node10171;
													assign node10171 = (inp[10]) ? node10185 : node10172;
														assign node10172 = (inp[0]) ? node10180 : node10173;
															assign node10173 = (inp[11]) ? node10177 : node10174;
																assign node10174 = (inp[9]) ? 4'b1011 : 4'b1010;
																assign node10177 = (inp[9]) ? 4'b1010 : 4'b1011;
															assign node10180 = (inp[9]) ? 4'b1010 : node10181;
																assign node10181 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node10185 = (inp[0]) ? node10191 : node10186;
															assign node10186 = (inp[9]) ? 4'b1010 : node10187;
																assign node10187 = (inp[11]) ? 4'b1011 : 4'b1010;
															assign node10191 = (inp[9]) ? node10193 : 4'b1010;
																assign node10193 = (inp[11]) ? 4'b1010 : 4'b1011;
													assign node10196 = (inp[10]) ? node10206 : node10197;
														assign node10197 = (inp[0]) ? 4'b1011 : node10198;
															assign node10198 = (inp[9]) ? node10202 : node10199;
																assign node10199 = (inp[11]) ? 4'b1011 : 4'b1010;
																assign node10202 = (inp[11]) ? 4'b1010 : 4'b1011;
														assign node10206 = (inp[0]) ? node10214 : node10207;
															assign node10207 = (inp[9]) ? node10211 : node10208;
																assign node10208 = (inp[11]) ? 4'b1011 : 4'b1010;
																assign node10211 = (inp[11]) ? 4'b1010 : 4'b1011;
															assign node10214 = (inp[11]) ? node10216 : 4'b1010;
																assign node10216 = (inp[9]) ? 4'b1011 : 4'b1010;
									assign node10219 = (inp[7]) ? node10315 : node10220;
										assign node10220 = (inp[9]) ? node10268 : node10221;
											assign node10221 = (inp[11]) ? node10245 : node10222;
												assign node10222 = (inp[1]) ? node10234 : node10223;
													assign node10223 = (inp[4]) ? node10229 : node10224;
														assign node10224 = (inp[2]) ? 4'b1010 : node10225;
															assign node10225 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node10229 = (inp[0]) ? 4'b1111 : node10230;
															assign node10230 = (inp[2]) ? 4'b1111 : 4'b1110;
													assign node10234 = (inp[4]) ? node10240 : node10235;
														assign node10235 = (inp[0]) ? 4'b1110 : node10236;
															assign node10236 = (inp[2]) ? 4'b1111 : 4'b1110;
														assign node10240 = (inp[0]) ? 4'b1010 : node10241;
															assign node10241 = (inp[2]) ? 4'b1010 : 4'b1011;
												assign node10245 = (inp[4]) ? node10257 : node10246;
													assign node10246 = (inp[1]) ? node10252 : node10247;
														assign node10247 = (inp[2]) ? 4'b1011 : node10248;
															assign node10248 = (inp[0]) ? 4'b1010 : 4'b1011;
														assign node10252 = (inp[0]) ? 4'b1111 : node10253;
															assign node10253 = (inp[2]) ? 4'b1110 : 4'b1111;
													assign node10257 = (inp[1]) ? node10263 : node10258;
														assign node10258 = (inp[2]) ? 4'b1110 : node10259;
															assign node10259 = (inp[0]) ? 4'b1110 : 4'b1111;
														assign node10263 = (inp[0]) ? 4'b1011 : node10264;
															assign node10264 = (inp[2]) ? 4'b1011 : 4'b1010;
											assign node10268 = (inp[11]) ? node10292 : node10269;
												assign node10269 = (inp[4]) ? node10281 : node10270;
													assign node10270 = (inp[1]) ? node10276 : node10271;
														assign node10271 = (inp[0]) ? node10273 : 4'b1011;
															assign node10273 = (inp[2]) ? 4'b1011 : 4'b1010;
														assign node10276 = (inp[2]) ? node10278 : 4'b1111;
															assign node10278 = (inp[0]) ? 4'b1111 : 4'b1110;
													assign node10281 = (inp[1]) ? node10287 : node10282;
														assign node10282 = (inp[0]) ? 4'b1110 : node10283;
															assign node10283 = (inp[2]) ? 4'b1110 : 4'b1111;
														assign node10287 = (inp[0]) ? 4'b1011 : node10288;
															assign node10288 = (inp[2]) ? 4'b1011 : 4'b1010;
												assign node10292 = (inp[4]) ? node10304 : node10293;
													assign node10293 = (inp[1]) ? node10299 : node10294;
														assign node10294 = (inp[2]) ? 4'b1010 : node10295;
															assign node10295 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node10299 = (inp[2]) ? node10301 : 4'b1110;
															assign node10301 = (inp[0]) ? 4'b1110 : 4'b1111;
													assign node10304 = (inp[1]) ? node10310 : node10305;
														assign node10305 = (inp[0]) ? 4'b1111 : node10306;
															assign node10306 = (inp[2]) ? 4'b1111 : 4'b1110;
														assign node10310 = (inp[0]) ? 4'b1010 : node10311;
															assign node10311 = (inp[2]) ? 4'b1010 : 4'b1011;
										assign node10315 = (inp[9]) ? node10365 : node10316;
											assign node10316 = (inp[2]) ? node10336 : node10317;
												assign node10317 = (inp[11]) ? node10327 : node10318;
													assign node10318 = (inp[1]) ? node10322 : node10319;
														assign node10319 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node10322 = (inp[4]) ? 4'b1001 : node10323;
															assign node10323 = (inp[0]) ? 4'b1100 : 4'b1101;
													assign node10327 = (inp[1]) ? node10331 : node10328;
														assign node10328 = (inp[4]) ? 4'b1101 : 4'b1001;
														assign node10331 = (inp[4]) ? 4'b1000 : node10332;
															assign node10332 = (inp[0]) ? 4'b1101 : 4'b1100;
												assign node10336 = (inp[11]) ? node10352 : node10337;
													assign node10337 = (inp[0]) ? node10345 : node10338;
														assign node10338 = (inp[4]) ? node10342 : node10339;
															assign node10339 = (inp[1]) ? 4'b1101 : 4'b1001;
															assign node10342 = (inp[1]) ? 4'b1001 : 4'b1100;
														assign node10345 = (inp[1]) ? node10349 : node10346;
															assign node10346 = (inp[4]) ? 4'b1101 : 4'b1000;
															assign node10349 = (inp[4]) ? 4'b1000 : 4'b1101;
													assign node10352 = (inp[1]) ? node10360 : node10353;
														assign node10353 = (inp[4]) ? node10357 : node10354;
															assign node10354 = (inp[0]) ? 4'b1001 : 4'b1000;
															assign node10357 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node10360 = (inp[4]) ? node10362 : 4'b1100;
															assign node10362 = (inp[0]) ? 4'b1001 : 4'b1000;
											assign node10365 = (inp[1]) ? node10389 : node10366;
												assign node10366 = (inp[4]) ? node10378 : node10367;
													assign node10367 = (inp[11]) ? node10373 : node10368;
														assign node10368 = (inp[2]) ? node10370 : 4'b1001;
															assign node10370 = (inp[0]) ? 4'b1001 : 4'b1000;
														assign node10373 = (inp[0]) ? 4'b1000 : node10374;
															assign node10374 = (inp[2]) ? 4'b1001 : 4'b1000;
													assign node10378 = (inp[11]) ? node10384 : node10379;
														assign node10379 = (inp[0]) ? node10381 : 4'b1101;
															assign node10381 = (inp[2]) ? 4'b1100 : 4'b1101;
														assign node10384 = (inp[0]) ? node10386 : 4'b1100;
															assign node10386 = (inp[2]) ? 4'b1101 : 4'b1100;
												assign node10389 = (inp[4]) ? node10401 : node10390;
													assign node10390 = (inp[11]) ? node10396 : node10391;
														assign node10391 = (inp[2]) ? 4'b1100 : node10392;
															assign node10392 = (inp[0]) ? 4'b1101 : 4'b1100;
														assign node10396 = (inp[2]) ? 4'b1101 : node10397;
															assign node10397 = (inp[0]) ? 4'b1100 : 4'b1101;
													assign node10401 = (inp[11]) ? node10407 : node10402;
														assign node10402 = (inp[0]) ? node10404 : 4'b1000;
															assign node10404 = (inp[2]) ? 4'b1001 : 4'b1000;
														assign node10407 = (inp[0]) ? node10409 : 4'b1001;
															assign node10409 = (inp[2]) ? 4'b1000 : 4'b1001;
								assign node10412 = (inp[15]) ? node10616 : node10413;
									assign node10413 = (inp[7]) ? node10519 : node10414;
										assign node10414 = (inp[4]) ? node10462 : node10415;
											assign node10415 = (inp[9]) ? node10439 : node10416;
												assign node10416 = (inp[1]) ? node10428 : node10417;
													assign node10417 = (inp[11]) ? node10423 : node10418;
														assign node10418 = (inp[0]) ? node10420 : 4'b1000;
															assign node10420 = (inp[2]) ? 4'b1000 : 4'b1001;
														assign node10423 = (inp[0]) ? node10425 : 4'b1001;
															assign node10425 = (inp[2]) ? 4'b1001 : 4'b1000;
													assign node10428 = (inp[11]) ? node10434 : node10429;
														assign node10429 = (inp[0]) ? 4'b1001 : node10430;
															assign node10430 = (inp[2]) ? 4'b1000 : 4'b1001;
														assign node10434 = (inp[2]) ? node10436 : 4'b1000;
															assign node10436 = (inp[0]) ? 4'b1000 : 4'b1001;
												assign node10439 = (inp[0]) ? node10451 : node10440;
													assign node10440 = (inp[11]) ? node10446 : node10441;
														assign node10441 = (inp[2]) ? 4'b1001 : node10442;
															assign node10442 = (inp[1]) ? 4'b1000 : 4'b1001;
														assign node10446 = (inp[1]) ? node10448 : 4'b1000;
															assign node10448 = (inp[2]) ? 4'b1000 : 4'b1001;
													assign node10451 = (inp[11]) ? node10457 : node10452;
														assign node10452 = (inp[1]) ? 4'b1000 : node10453;
															assign node10453 = (inp[2]) ? 4'b1001 : 4'b1000;
														assign node10457 = (inp[2]) ? node10459 : 4'b1001;
															assign node10459 = (inp[1]) ? 4'b1001 : 4'b1000;
											assign node10462 = (inp[1]) ? node10482 : node10463;
												assign node10463 = (inp[9]) ? node10475 : node10464;
													assign node10464 = (inp[11]) ? node10470 : node10465;
														assign node10465 = (inp[0]) ? node10467 : 4'b1000;
															assign node10467 = (inp[2]) ? 4'b1001 : 4'b1000;
														assign node10470 = (inp[0]) ? node10472 : 4'b1001;
															assign node10472 = (inp[2]) ? 4'b1000 : 4'b1001;
													assign node10475 = (inp[11]) ? 4'b1000 : node10476;
														assign node10476 = (inp[2]) ? node10478 : 4'b1001;
															assign node10478 = (inp[0]) ? 4'b1000 : 4'b1001;
												assign node10482 = (inp[2]) ? node10490 : node10483;
													assign node10483 = (inp[9]) ? node10487 : node10484;
														assign node10484 = (inp[11]) ? 4'b1100 : 4'b1101;
														assign node10487 = (inp[11]) ? 4'b1101 : 4'b1100;
													assign node10490 = (inp[9]) ? node10504 : node10491;
														assign node10491 = (inp[10]) ? node10497 : node10492;
															assign node10492 = (inp[11]) ? 4'b1100 : node10493;
																assign node10493 = (inp[0]) ? 4'b1100 : 4'b1101;
															assign node10497 = (inp[11]) ? node10501 : node10498;
																assign node10498 = (inp[0]) ? 4'b1100 : 4'b1101;
																assign node10501 = (inp[0]) ? 4'b1101 : 4'b1100;
														assign node10504 = (inp[10]) ? node10512 : node10505;
															assign node10505 = (inp[0]) ? node10509 : node10506;
																assign node10506 = (inp[11]) ? 4'b1101 : 4'b1100;
																assign node10509 = (inp[11]) ? 4'b1100 : 4'b1101;
															assign node10512 = (inp[0]) ? node10516 : node10513;
																assign node10513 = (inp[11]) ? 4'b1101 : 4'b1100;
																assign node10516 = (inp[11]) ? 4'b1100 : 4'b1101;
										assign node10519 = (inp[1]) ? node10563 : node10520;
											assign node10520 = (inp[4]) ? node10544 : node10521;
												assign node10521 = (inp[9]) ? node10533 : node10522;
													assign node10522 = (inp[11]) ? node10528 : node10523;
														assign node10523 = (inp[0]) ? 4'b1110 : node10524;
															assign node10524 = (inp[2]) ? 4'b1111 : 4'b1110;
														assign node10528 = (inp[0]) ? 4'b1111 : node10529;
															assign node10529 = (inp[2]) ? 4'b1110 : 4'b1111;
													assign node10533 = (inp[11]) ? node10539 : node10534;
														assign node10534 = (inp[0]) ? 4'b1111 : node10535;
															assign node10535 = (inp[2]) ? 4'b1110 : 4'b1111;
														assign node10539 = (inp[2]) ? node10541 : 4'b1110;
															assign node10541 = (inp[0]) ? 4'b1110 : 4'b1111;
												assign node10544 = (inp[11]) ? node10552 : node10545;
													assign node10545 = (inp[9]) ? node10547 : 4'b1010;
														assign node10547 = (inp[2]) ? 4'b1011 : node10548;
															assign node10548 = (inp[0]) ? 4'b1011 : 4'b1010;
													assign node10552 = (inp[9]) ? node10558 : node10553;
														assign node10553 = (inp[0]) ? 4'b1011 : node10554;
															assign node10554 = (inp[2]) ? 4'b1011 : 4'b1010;
														assign node10558 = (inp[0]) ? 4'b1010 : node10559;
															assign node10559 = (inp[2]) ? 4'b1010 : 4'b1011;
											assign node10563 = (inp[11]) ? node10589 : node10564;
												assign node10564 = (inp[9]) ? node10580 : node10565;
													assign node10565 = (inp[0]) ? node10567 : 4'b1010;
														assign node10567 = (inp[10]) ? node10575 : node10568;
															assign node10568 = (inp[2]) ? node10572 : node10569;
																assign node10569 = (inp[4]) ? 4'b1010 : 4'b1011;
																assign node10572 = (inp[4]) ? 4'b1011 : 4'b1010;
															assign node10575 = (inp[2]) ? 4'b1010 : node10576;
																assign node10576 = (inp[4]) ? 4'b1010 : 4'b1011;
													assign node10580 = (inp[0]) ? node10582 : 4'b1011;
														assign node10582 = (inp[2]) ? node10586 : node10583;
															assign node10583 = (inp[4]) ? 4'b1011 : 4'b1010;
															assign node10586 = (inp[4]) ? 4'b1010 : 4'b1011;
												assign node10589 = (inp[9]) ? node10599 : node10590;
													assign node10590 = (inp[0]) ? node10592 : 4'b1011;
														assign node10592 = (inp[2]) ? node10596 : node10593;
															assign node10593 = (inp[4]) ? 4'b1011 : 4'b1010;
															assign node10596 = (inp[4]) ? 4'b1010 : 4'b1011;
													assign node10599 = (inp[0]) ? node10601 : 4'b1010;
														assign node10601 = (inp[10]) ? node10609 : node10602;
															assign node10602 = (inp[4]) ? node10606 : node10603;
																assign node10603 = (inp[2]) ? 4'b1010 : 4'b1011;
																assign node10606 = (inp[2]) ? 4'b1011 : 4'b1010;
															assign node10609 = (inp[4]) ? node10613 : node10610;
																assign node10610 = (inp[2]) ? 4'b1010 : 4'b1011;
																assign node10613 = (inp[2]) ? 4'b1011 : 4'b1010;
									assign node10616 = (inp[7]) ? node10758 : node10617;
										assign node10617 = (inp[4]) ? node10699 : node10618;
											assign node10618 = (inp[10]) ? node10676 : node10619;
												assign node10619 = (inp[1]) ? node10649 : node10620;
													assign node10620 = (inp[0]) ? node10636 : node10621;
														assign node10621 = (inp[2]) ? node10629 : node10622;
															assign node10622 = (inp[11]) ? node10626 : node10623;
																assign node10623 = (inp[9]) ? 4'b1011 : 4'b1010;
																assign node10626 = (inp[9]) ? 4'b1010 : 4'b1011;
															assign node10629 = (inp[9]) ? node10633 : node10630;
																assign node10630 = (inp[11]) ? 4'b1011 : 4'b1010;
																assign node10633 = (inp[11]) ? 4'b1010 : 4'b1011;
														assign node10636 = (inp[11]) ? node10642 : node10637;
															assign node10637 = (inp[2]) ? node10639 : 4'b1010;
																assign node10639 = (inp[9]) ? 4'b1011 : 4'b1010;
															assign node10642 = (inp[2]) ? node10646 : node10643;
																assign node10643 = (inp[9]) ? 4'b1011 : 4'b1010;
																assign node10646 = (inp[9]) ? 4'b1010 : 4'b1011;
													assign node10649 = (inp[0]) ? node10661 : node10650;
														assign node10650 = (inp[2]) ? node10656 : node10651;
															assign node10651 = (inp[9]) ? node10653 : 4'b1010;
																assign node10653 = (inp[11]) ? 4'b1010 : 4'b1011;
															assign node10656 = (inp[9]) ? 4'b1010 : node10657;
																assign node10657 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node10661 = (inp[2]) ? node10669 : node10662;
															assign node10662 = (inp[11]) ? node10666 : node10663;
																assign node10663 = (inp[9]) ? 4'b1010 : 4'b1011;
																assign node10666 = (inp[9]) ? 4'b1011 : 4'b1010;
															assign node10669 = (inp[11]) ? node10673 : node10670;
																assign node10670 = (inp[9]) ? 4'b1011 : 4'b1010;
																assign node10673 = (inp[9]) ? 4'b1010 : 4'b1011;
												assign node10676 = (inp[11]) ? node10688 : node10677;
													assign node10677 = (inp[9]) ? node10683 : node10678;
														assign node10678 = (inp[0]) ? node10680 : 4'b1010;
															assign node10680 = (inp[2]) ? 4'b1010 : 4'b1011;
														assign node10683 = (inp[0]) ? node10685 : 4'b1011;
															assign node10685 = (inp[2]) ? 4'b1011 : 4'b1010;
													assign node10688 = (inp[9]) ? node10694 : node10689;
														assign node10689 = (inp[2]) ? 4'b1011 : node10690;
															assign node10690 = (inp[0]) ? 4'b1010 : 4'b1011;
														assign node10694 = (inp[0]) ? node10696 : 4'b1010;
															assign node10696 = (inp[2]) ? 4'b1010 : 4'b1011;
											assign node10699 = (inp[0]) ? node10707 : node10700;
												assign node10700 = (inp[11]) ? node10704 : node10701;
													assign node10701 = (inp[9]) ? 4'b1011 : 4'b1010;
													assign node10704 = (inp[9]) ? 4'b1010 : 4'b1011;
												assign node10707 = (inp[1]) ? node10729 : node10708;
													assign node10708 = (inp[10]) ? node10720 : node10709;
														assign node10709 = (inp[11]) ? node10715 : node10710;
															assign node10710 = (inp[9]) ? node10712 : 4'b1010;
																assign node10712 = (inp[2]) ? 4'b1010 : 4'b1011;
															assign node10715 = (inp[9]) ? node10717 : 4'b1011;
																assign node10717 = (inp[2]) ? 4'b1011 : 4'b1010;
														assign node10720 = (inp[11]) ? node10722 : 4'b1011;
															assign node10722 = (inp[2]) ? node10726 : node10723;
																assign node10723 = (inp[9]) ? 4'b1010 : 4'b1011;
																assign node10726 = (inp[9]) ? 4'b1011 : 4'b1010;
													assign node10729 = (inp[2]) ? node10743 : node10730;
														assign node10730 = (inp[10]) ? node10736 : node10731;
															assign node10731 = (inp[9]) ? 4'b1011 : node10732;
																assign node10732 = (inp[11]) ? 4'b1011 : 4'b1010;
															assign node10736 = (inp[9]) ? node10740 : node10737;
																assign node10737 = (inp[11]) ? 4'b1011 : 4'b1010;
																assign node10740 = (inp[11]) ? 4'b1010 : 4'b1011;
														assign node10743 = (inp[10]) ? node10751 : node10744;
															assign node10744 = (inp[9]) ? node10748 : node10745;
																assign node10745 = (inp[11]) ? 4'b1010 : 4'b1011;
																assign node10748 = (inp[11]) ? 4'b1011 : 4'b1010;
															assign node10751 = (inp[9]) ? node10755 : node10752;
																assign node10752 = (inp[11]) ? 4'b1010 : 4'b1011;
																assign node10755 = (inp[11]) ? 4'b1011 : 4'b1010;
										assign node10758 = (inp[4]) ? node10782 : node10759;
											assign node10759 = (inp[9]) ? node10771 : node10760;
												assign node10760 = (inp[11]) ? node10766 : node10761;
													assign node10761 = (inp[0]) ? node10763 : 4'b1001;
														assign node10763 = (inp[2]) ? 4'b1001 : 4'b1000;
													assign node10766 = (inp[0]) ? node10768 : 4'b1000;
														assign node10768 = (inp[2]) ? 4'b1000 : 4'b1001;
												assign node10771 = (inp[11]) ? node10777 : node10772;
													assign node10772 = (inp[2]) ? 4'b1000 : node10773;
														assign node10773 = (inp[0]) ? 4'b1001 : 4'b1000;
													assign node10777 = (inp[2]) ? 4'b1001 : node10778;
														assign node10778 = (inp[0]) ? 4'b1000 : 4'b1001;
											assign node10782 = (inp[0]) ? node10790 : node10783;
												assign node10783 = (inp[11]) ? node10787 : node10784;
													assign node10784 = (inp[9]) ? 4'b1000 : 4'b1001;
													assign node10787 = (inp[9]) ? 4'b1001 : 4'b1000;
												assign node10790 = (inp[9]) ? node10800 : node10791;
													assign node10791 = (inp[1]) ? 4'b1001 : node10792;
														assign node10792 = (inp[2]) ? node10796 : node10793;
															assign node10793 = (inp[11]) ? 4'b1000 : 4'b1001;
															assign node10796 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node10800 = (inp[1]) ? node10812 : node10801;
														assign node10801 = (inp[10]) ? node10807 : node10802;
															assign node10802 = (inp[2]) ? node10804 : 4'b1001;
																assign node10804 = (inp[11]) ? 4'b1000 : 4'b1001;
															assign node10807 = (inp[2]) ? 4'b1001 : node10808;
																assign node10808 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node10812 = (inp[2]) ? node10816 : node10813;
															assign node10813 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node10816 = (inp[11]) ? 4'b1000 : 4'b1001;
						assign node10819 = (inp[6]) ? node12065 : node10820;
							assign node10820 = (inp[2]) ? node11438 : node10821;
								assign node10821 = (inp[12]) ? node11157 : node10822;
									assign node10822 = (inp[7]) ? node10986 : node10823;
										assign node10823 = (inp[4]) ? node10913 : node10824;
											assign node10824 = (inp[11]) ? node10864 : node10825;
												assign node10825 = (inp[1]) ? node10843 : node10826;
													assign node10826 = (inp[10]) ? 4'b1001 : node10827;
														assign node10827 = (inp[15]) ? node10835 : node10828;
															assign node10828 = (inp[0]) ? node10832 : node10829;
																assign node10829 = (inp[9]) ? 4'b1001 : 4'b1000;
																assign node10832 = (inp[9]) ? 4'b1000 : 4'b1001;
															assign node10835 = (inp[0]) ? node10839 : node10836;
																assign node10836 = (inp[9]) ? 4'b1001 : 4'b1000;
																assign node10839 = (inp[9]) ? 4'b1000 : 4'b1001;
													assign node10843 = (inp[10]) ? node10853 : node10844;
														assign node10844 = (inp[15]) ? node10846 : 4'b1001;
															assign node10846 = (inp[9]) ? node10850 : node10847;
																assign node10847 = (inp[0]) ? 4'b1000 : 4'b1001;
																assign node10850 = (inp[0]) ? 4'b1001 : 4'b1000;
														assign node10853 = (inp[9]) ? node10859 : node10854;
															assign node10854 = (inp[0]) ? 4'b1001 : node10855;
																assign node10855 = (inp[15]) ? 4'b1000 : 4'b1001;
															assign node10859 = (inp[15]) ? node10861 : 4'b1000;
																assign node10861 = (inp[0]) ? 4'b1000 : 4'b1001;
												assign node10864 = (inp[0]) ? node10892 : node10865;
													assign node10865 = (inp[15]) ? node10879 : node10866;
														assign node10866 = (inp[10]) ? node10874 : node10867;
															assign node10867 = (inp[9]) ? node10871 : node10868;
																assign node10868 = (inp[1]) ? 4'b1001 : 4'b1000;
																assign node10871 = (inp[1]) ? 4'b1000 : 4'b1001;
															assign node10874 = (inp[9]) ? 4'b1001 : node10875;
																assign node10875 = (inp[1]) ? 4'b1000 : 4'b1001;
														assign node10879 = (inp[9]) ? node10885 : node10880;
															assign node10880 = (inp[1]) ? node10882 : 4'b1000;
																assign node10882 = (inp[10]) ? 4'b1000 : 4'b1001;
															assign node10885 = (inp[10]) ? node10889 : node10886;
																assign node10886 = (inp[1]) ? 4'b1000 : 4'b1001;
																assign node10889 = (inp[1]) ? 4'b1001 : 4'b1000;
													assign node10892 = (inp[9]) ? node10904 : node10893;
														assign node10893 = (inp[10]) ? node10899 : node10894;
															assign node10894 = (inp[1]) ? node10896 : 4'b1000;
																assign node10896 = (inp[15]) ? 4'b1001 : 4'b1000;
															assign node10899 = (inp[15]) ? node10901 : 4'b1001;
																assign node10901 = (inp[1]) ? 4'b1000 : 4'b1001;
														assign node10904 = (inp[10]) ? node10908 : node10905;
															assign node10905 = (inp[1]) ? 4'b1000 : 4'b1001;
															assign node10908 = (inp[1]) ? node10910 : 4'b1000;
																assign node10910 = (inp[15]) ? 4'b1001 : 4'b1000;
											assign node10913 = (inp[15]) ? node10945 : node10914;
												assign node10914 = (inp[9]) ? node10932 : node10915;
													assign node10915 = (inp[11]) ? node10921 : node10916;
														assign node10916 = (inp[10]) ? node10918 : 4'b1010;
															assign node10918 = (inp[1]) ? 4'b1010 : 4'b1011;
														assign node10921 = (inp[10]) ? node10927 : node10922;
															assign node10922 = (inp[1]) ? 4'b1011 : node10923;
																assign node10923 = (inp[0]) ? 4'b1010 : 4'b1011;
															assign node10927 = (inp[0]) ? node10929 : 4'b1010;
																assign node10929 = (inp[1]) ? 4'b1010 : 4'b1011;
													assign node10932 = (inp[11]) ? node10940 : node10933;
														assign node10933 = (inp[10]) ? node10937 : node10934;
															assign node10934 = (inp[1]) ? 4'b1010 : 4'b1011;
															assign node10937 = (inp[1]) ? 4'b1011 : 4'b1010;
														assign node10940 = (inp[10]) ? 4'b1011 : node10941;
															assign node10941 = (inp[1]) ? 4'b1010 : 4'b1011;
												assign node10945 = (inp[10]) ? node10963 : node10946;
													assign node10946 = (inp[11]) ? node10954 : node10947;
														assign node10947 = (inp[9]) ? node10951 : node10948;
															assign node10948 = (inp[1]) ? 4'b1101 : 4'b1100;
															assign node10951 = (inp[1]) ? 4'b1100 : 4'b1101;
														assign node10954 = (inp[9]) ? node10956 : 4'b1100;
															assign node10956 = (inp[0]) ? node10960 : node10957;
																assign node10957 = (inp[1]) ? 4'b1101 : 4'b1100;
																assign node10960 = (inp[1]) ? 4'b1100 : 4'b1101;
													assign node10963 = (inp[0]) ? node10975 : node10964;
														assign node10964 = (inp[9]) ? node10970 : node10965;
															assign node10965 = (inp[1]) ? node10967 : 4'b1101;
																assign node10967 = (inp[11]) ? 4'b1101 : 4'b1100;
															assign node10970 = (inp[1]) ? node10972 : 4'b1100;
																assign node10972 = (inp[11]) ? 4'b1100 : 4'b1101;
														assign node10975 = (inp[11]) ? node10981 : node10976;
															assign node10976 = (inp[1]) ? node10978 : 4'b1101;
																assign node10978 = (inp[9]) ? 4'b1101 : 4'b1100;
															assign node10981 = (inp[9]) ? node10983 : 4'b1101;
																assign node10983 = (inp[1]) ? 4'b1101 : 4'b1100;
										assign node10986 = (inp[15]) ? node11076 : node10987;
											assign node10987 = (inp[4]) ? node11023 : node10988;
												assign node10988 = (inp[1]) ? node11008 : node10989;
													assign node10989 = (inp[9]) ? node10999 : node10990;
														assign node10990 = (inp[10]) ? node10996 : node10991;
															assign node10991 = (inp[11]) ? 4'b1111 : node10992;
																assign node10992 = (inp[0]) ? 4'b1110 : 4'b1111;
															assign node10996 = (inp[11]) ? 4'b1110 : 4'b1111;
														assign node10999 = (inp[10]) ? node11003 : node11000;
															assign node11000 = (inp[0]) ? 4'b1111 : 4'b1110;
															assign node11003 = (inp[11]) ? 4'b1111 : node11004;
																assign node11004 = (inp[0]) ? 4'b1110 : 4'b1111;
													assign node11008 = (inp[10]) ? node11018 : node11009;
														assign node11009 = (inp[9]) ? node11013 : node11010;
															assign node11010 = (inp[11]) ? 4'b1010 : 4'b1011;
															assign node11013 = (inp[0]) ? 4'b1010 : node11014;
																assign node11014 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node11018 = (inp[9]) ? node11020 : 4'b1010;
															assign node11020 = (inp[0]) ? 4'b1011 : 4'b1010;
												assign node11023 = (inp[11]) ? node11045 : node11024;
													assign node11024 = (inp[10]) ? node11036 : node11025;
														assign node11025 = (inp[9]) ? node11031 : node11026;
															assign node11026 = (inp[1]) ? node11028 : 4'b1101;
																assign node11028 = (inp[0]) ? 4'b1101 : 4'b1100;
															assign node11031 = (inp[1]) ? node11033 : 4'b1100;
																assign node11033 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node11036 = (inp[9]) ? node11040 : node11037;
															assign node11037 = (inp[1]) ? 4'b1101 : 4'b1100;
															assign node11040 = (inp[1]) ? node11042 : 4'b1101;
																assign node11042 = (inp[0]) ? 4'b1101 : 4'b1100;
													assign node11045 = (inp[0]) ? node11061 : node11046;
														assign node11046 = (inp[1]) ? node11054 : node11047;
															assign node11047 = (inp[9]) ? node11051 : node11048;
																assign node11048 = (inp[10]) ? 4'b1101 : 4'b1100;
																assign node11051 = (inp[10]) ? 4'b1100 : 4'b1101;
															assign node11054 = (inp[10]) ? node11058 : node11055;
																assign node11055 = (inp[9]) ? 4'b1101 : 4'b1100;
																assign node11058 = (inp[9]) ? 4'b1100 : 4'b1101;
														assign node11061 = (inp[1]) ? node11069 : node11062;
															assign node11062 = (inp[9]) ? node11066 : node11063;
																assign node11063 = (inp[10]) ? 4'b1100 : 4'b1101;
																assign node11066 = (inp[10]) ? 4'b1101 : 4'b1100;
															assign node11069 = (inp[10]) ? node11073 : node11070;
																assign node11070 = (inp[9]) ? 4'b1101 : 4'b1100;
																assign node11073 = (inp[9]) ? 4'b1100 : 4'b1101;
											assign node11076 = (inp[10]) ? node11120 : node11077;
												assign node11077 = (inp[4]) ? node11101 : node11078;
													assign node11078 = (inp[1]) ? node11090 : node11079;
														assign node11079 = (inp[9]) ? node11085 : node11080;
															assign node11080 = (inp[0]) ? 4'b1011 : node11081;
																assign node11081 = (inp[11]) ? 4'b1010 : 4'b1011;
															assign node11085 = (inp[11]) ? node11087 : 4'b1010;
																assign node11087 = (inp[0]) ? 4'b1010 : 4'b1011;
														assign node11090 = (inp[9]) ? node11096 : node11091;
															assign node11091 = (inp[11]) ? 4'b1110 : node11092;
																assign node11092 = (inp[0]) ? 4'b1111 : 4'b1110;
															assign node11096 = (inp[11]) ? 4'b1111 : node11097;
																assign node11097 = (inp[0]) ? 4'b1110 : 4'b1111;
													assign node11101 = (inp[1]) ? node11111 : node11102;
														assign node11102 = (inp[9]) ? node11108 : node11103;
															assign node11103 = (inp[0]) ? node11105 : 4'b1110;
																assign node11105 = (inp[11]) ? 4'b1110 : 4'b1111;
															assign node11108 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node11111 = (inp[9]) ? node11115 : node11112;
															assign node11112 = (inp[11]) ? 4'b1011 : 4'b1010;
															assign node11115 = (inp[0]) ? node11117 : 4'b1010;
																assign node11117 = (inp[11]) ? 4'b1010 : 4'b1011;
												assign node11120 = (inp[11]) ? node11146 : node11121;
													assign node11121 = (inp[9]) ? node11135 : node11122;
														assign node11122 = (inp[4]) ? node11128 : node11123;
															assign node11123 = (inp[1]) ? node11125 : 4'b1010;
																assign node11125 = (inp[0]) ? 4'b1110 : 4'b1111;
															assign node11128 = (inp[1]) ? node11132 : node11129;
																assign node11129 = (inp[0]) ? 4'b1110 : 4'b1111;
																assign node11132 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node11135 = (inp[4]) ? node11139 : node11136;
															assign node11136 = (inp[1]) ? 4'b1111 : 4'b1011;
															assign node11139 = (inp[1]) ? node11143 : node11140;
																assign node11140 = (inp[0]) ? 4'b1111 : 4'b1110;
																assign node11143 = (inp[0]) ? 4'b1010 : 4'b1011;
													assign node11146 = (inp[1]) ? node11150 : node11147;
														assign node11147 = (inp[4]) ? 4'b1111 : 4'b1011;
														assign node11150 = (inp[4]) ? node11154 : node11151;
															assign node11151 = (inp[9]) ? 4'b1110 : 4'b1111;
															assign node11154 = (inp[9]) ? 4'b1011 : 4'b1010;
									assign node11157 = (inp[7]) ? node11293 : node11158;
										assign node11158 = (inp[15]) ? node11240 : node11159;
											assign node11159 = (inp[4]) ? node11197 : node11160;
												assign node11160 = (inp[1]) ? node11184 : node11161;
													assign node11161 = (inp[11]) ? node11177 : node11162;
														assign node11162 = (inp[10]) ? node11170 : node11163;
															assign node11163 = (inp[9]) ? node11167 : node11164;
																assign node11164 = (inp[0]) ? 4'b1011 : 4'b1010;
																assign node11167 = (inp[0]) ? 4'b1010 : 4'b1011;
															assign node11170 = (inp[9]) ? node11174 : node11171;
																assign node11171 = (inp[0]) ? 4'b1010 : 4'b1011;
																assign node11174 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node11177 = (inp[10]) ? node11181 : node11178;
															assign node11178 = (inp[9]) ? 4'b1011 : 4'b1010;
															assign node11181 = (inp[9]) ? 4'b1010 : 4'b1011;
													assign node11184 = (inp[9]) ? node11192 : node11185;
														assign node11185 = (inp[10]) ? 4'b1010 : node11186;
															assign node11186 = (inp[0]) ? 4'b1011 : node11187;
																assign node11187 = (inp[11]) ? 4'b1010 : 4'b1011;
														assign node11192 = (inp[10]) ? 4'b1011 : node11193;
															assign node11193 = (inp[11]) ? 4'b1011 : 4'b1010;
												assign node11197 = (inp[1]) ? node11221 : node11198;
													assign node11198 = (inp[10]) ? node11210 : node11199;
														assign node11199 = (inp[9]) ? node11205 : node11200;
															assign node11200 = (inp[11]) ? 4'b1001 : node11201;
																assign node11201 = (inp[0]) ? 4'b1000 : 4'b1001;
															assign node11205 = (inp[0]) ? node11207 : 4'b1000;
																assign node11207 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node11210 = (inp[9]) ? node11216 : node11211;
															assign node11211 = (inp[0]) ? node11213 : 4'b1000;
																assign node11213 = (inp[11]) ? 4'b1000 : 4'b1001;
															assign node11216 = (inp[11]) ? 4'b1001 : node11217;
																assign node11217 = (inp[0]) ? 4'b1000 : 4'b1001;
													assign node11221 = (inp[9]) ? node11233 : node11222;
														assign node11222 = (inp[10]) ? node11228 : node11223;
															assign node11223 = (inp[11]) ? 4'b1100 : node11224;
																assign node11224 = (inp[0]) ? 4'b1101 : 4'b1100;
															assign node11228 = (inp[0]) ? node11230 : 4'b1101;
																assign node11230 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node11233 = (inp[10]) ? 4'b1100 : node11234;
															assign node11234 = (inp[11]) ? 4'b1101 : node11235;
																assign node11235 = (inp[0]) ? 4'b1100 : 4'b1101;
											assign node11240 = (inp[10]) ? node11264 : node11241;
												assign node11241 = (inp[4]) ? node11253 : node11242;
													assign node11242 = (inp[9]) ? node11248 : node11243;
														assign node11243 = (inp[11]) ? 4'b1010 : node11244;
															assign node11244 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node11248 = (inp[11]) ? 4'b1011 : node11249;
															assign node11249 = (inp[0]) ? 4'b1010 : 4'b1011;
													assign node11253 = (inp[9]) ? node11259 : node11254;
														assign node11254 = (inp[0]) ? node11256 : 4'b1011;
															assign node11256 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node11259 = (inp[0]) ? node11261 : 4'b1010;
															assign node11261 = (inp[11]) ? 4'b1010 : 4'b1011;
												assign node11264 = (inp[0]) ? node11272 : node11265;
													assign node11265 = (inp[4]) ? node11269 : node11266;
														assign node11266 = (inp[9]) ? 4'b1010 : 4'b1011;
														assign node11269 = (inp[9]) ? 4'b1011 : 4'b1010;
													assign node11272 = (inp[4]) ? node11280 : node11273;
														assign node11273 = (inp[11]) ? node11277 : node11274;
															assign node11274 = (inp[9]) ? 4'b1011 : 4'b1010;
															assign node11277 = (inp[9]) ? 4'b1010 : 4'b1011;
														assign node11280 = (inp[1]) ? node11288 : node11281;
															assign node11281 = (inp[9]) ? node11285 : node11282;
																assign node11282 = (inp[11]) ? 4'b1010 : 4'b1011;
																assign node11285 = (inp[11]) ? 4'b1011 : 4'b1010;
															assign node11288 = (inp[11]) ? 4'b1010 : node11289;
																assign node11289 = (inp[9]) ? 4'b1010 : 4'b1011;
										assign node11293 = (inp[15]) ? node11367 : node11294;
											assign node11294 = (inp[4]) ? node11336 : node11295;
												assign node11295 = (inp[0]) ? node11317 : node11296;
													assign node11296 = (inp[11]) ? node11304 : node11297;
														assign node11297 = (inp[9]) ? node11301 : node11298;
															assign node11298 = (inp[10]) ? 4'b1100 : 4'b1101;
															assign node11301 = (inp[10]) ? 4'b1101 : 4'b1100;
														assign node11304 = (inp[9]) ? node11312 : node11305;
															assign node11305 = (inp[1]) ? node11309 : node11306;
																assign node11306 = (inp[10]) ? 4'b1101 : 4'b1100;
																assign node11309 = (inp[10]) ? 4'b1100 : 4'b1101;
															assign node11312 = (inp[1]) ? node11314 : 4'b1101;
																assign node11314 = (inp[10]) ? 4'b1101 : 4'b1100;
													assign node11317 = (inp[9]) ? node11327 : node11318;
														assign node11318 = (inp[11]) ? node11324 : node11319;
															assign node11319 = (inp[10]) ? node11321 : 4'b1100;
																assign node11321 = (inp[1]) ? 4'b1101 : 4'b1100;
															assign node11324 = (inp[10]) ? 4'b1100 : 4'b1101;
														assign node11327 = (inp[10]) ? node11333 : node11328;
															assign node11328 = (inp[11]) ? 4'b1100 : node11329;
																assign node11329 = (inp[1]) ? 4'b1101 : 4'b1100;
															assign node11333 = (inp[11]) ? 4'b1101 : 4'b1100;
												assign node11336 = (inp[10]) ? node11356 : node11337;
													assign node11337 = (inp[9]) ? node11345 : node11338;
														assign node11338 = (inp[0]) ? node11340 : 4'b1010;
															assign node11340 = (inp[11]) ? 4'b1010 : node11341;
																assign node11341 = (inp[1]) ? 4'b1011 : 4'b1010;
														assign node11345 = (inp[0]) ? node11351 : node11346;
															assign node11346 = (inp[11]) ? node11348 : 4'b1011;
																assign node11348 = (inp[1]) ? 4'b1011 : 4'b1010;
															assign node11351 = (inp[11]) ? 4'b1011 : node11352;
																assign node11352 = (inp[1]) ? 4'b1010 : 4'b1011;
													assign node11356 = (inp[9]) ? node11358 : 4'b1011;
														assign node11358 = (inp[11]) ? node11364 : node11359;
															assign node11359 = (inp[0]) ? node11361 : 4'b1010;
																assign node11361 = (inp[1]) ? 4'b1011 : 4'b1010;
															assign node11364 = (inp[0]) ? 4'b1010 : 4'b1011;
											assign node11367 = (inp[9]) ? node11399 : node11368;
												assign node11368 = (inp[0]) ? node11376 : node11369;
													assign node11369 = (inp[4]) ? node11373 : node11370;
														assign node11370 = (inp[10]) ? 4'b1001 : 4'b1000;
														assign node11373 = (inp[10]) ? 4'b1000 : 4'b1001;
													assign node11376 = (inp[11]) ? node11384 : node11377;
														assign node11377 = (inp[10]) ? node11381 : node11378;
															assign node11378 = (inp[4]) ? 4'b1000 : 4'b1001;
															assign node11381 = (inp[4]) ? 4'b1001 : 4'b1000;
														assign node11384 = (inp[1]) ? node11392 : node11385;
															assign node11385 = (inp[10]) ? node11389 : node11386;
																assign node11386 = (inp[4]) ? 4'b1001 : 4'b1000;
																assign node11389 = (inp[4]) ? 4'b1000 : 4'b1001;
															assign node11392 = (inp[10]) ? node11396 : node11393;
																assign node11393 = (inp[4]) ? 4'b1001 : 4'b1000;
																assign node11396 = (inp[4]) ? 4'b1000 : 4'b1001;
												assign node11399 = (inp[1]) ? node11417 : node11400;
													assign node11400 = (inp[0]) ? node11408 : node11401;
														assign node11401 = (inp[10]) ? node11405 : node11402;
															assign node11402 = (inp[4]) ? 4'b1000 : 4'b1001;
															assign node11405 = (inp[4]) ? 4'b1001 : 4'b1000;
														assign node11408 = (inp[4]) ? node11410 : 4'b1000;
															assign node11410 = (inp[10]) ? node11414 : node11411;
																assign node11411 = (inp[11]) ? 4'b1000 : 4'b1001;
																assign node11414 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node11417 = (inp[11]) ? node11431 : node11418;
														assign node11418 = (inp[10]) ? node11426 : node11419;
															assign node11419 = (inp[0]) ? node11423 : node11420;
																assign node11420 = (inp[4]) ? 4'b1000 : 4'b1001;
																assign node11423 = (inp[4]) ? 4'b1001 : 4'b1000;
															assign node11426 = (inp[0]) ? 4'b1001 : node11427;
																assign node11427 = (inp[4]) ? 4'b1001 : 4'b1000;
														assign node11431 = (inp[4]) ? node11435 : node11432;
															assign node11432 = (inp[10]) ? 4'b1000 : 4'b1001;
															assign node11435 = (inp[10]) ? 4'b1001 : 4'b1000;
								assign node11438 = (inp[7]) ? node11776 : node11439;
									assign node11439 = (inp[12]) ? node11615 : node11440;
										assign node11440 = (inp[15]) ? node11534 : node11441;
											assign node11441 = (inp[4]) ? node11489 : node11442;
												assign node11442 = (inp[10]) ? node11466 : node11443;
													assign node11443 = (inp[9]) ? node11455 : node11444;
														assign node11444 = (inp[0]) ? node11450 : node11445;
															assign node11445 = (inp[11]) ? node11447 : 4'b1100;
																assign node11447 = (inp[1]) ? 4'b1101 : 4'b1100;
															assign node11450 = (inp[1]) ? 4'b1100 : node11451;
																assign node11451 = (inp[11]) ? 4'b1100 : 4'b1101;
														assign node11455 = (inp[11]) ? node11461 : node11456;
															assign node11456 = (inp[0]) ? node11458 : 4'b1101;
																assign node11458 = (inp[1]) ? 4'b1101 : 4'b1100;
															assign node11461 = (inp[1]) ? node11463 : 4'b1101;
																assign node11463 = (inp[0]) ? 4'b1101 : 4'b1100;
													assign node11466 = (inp[9]) ? node11478 : node11467;
														assign node11467 = (inp[0]) ? node11473 : node11468;
															assign node11468 = (inp[1]) ? node11470 : 4'b1101;
																assign node11470 = (inp[11]) ? 4'b1100 : 4'b1101;
															assign node11473 = (inp[11]) ? 4'b1101 : node11474;
																assign node11474 = (inp[1]) ? 4'b1101 : 4'b1100;
														assign node11478 = (inp[11]) ? node11484 : node11479;
															assign node11479 = (inp[0]) ? node11481 : 4'b1100;
																assign node11481 = (inp[1]) ? 4'b1100 : 4'b1101;
															assign node11484 = (inp[1]) ? node11486 : 4'b1100;
																assign node11486 = (inp[0]) ? 4'b1100 : 4'b1101;
												assign node11489 = (inp[11]) ? node11511 : node11490;
													assign node11490 = (inp[10]) ? node11502 : node11491;
														assign node11491 = (inp[9]) ? node11497 : node11492;
															assign node11492 = (inp[0]) ? 4'b1111 : node11493;
																assign node11493 = (inp[1]) ? 4'b1110 : 4'b1111;
															assign node11497 = (inp[0]) ? 4'b1110 : node11498;
																assign node11498 = (inp[1]) ? 4'b1111 : 4'b1110;
														assign node11502 = (inp[9]) ? node11506 : node11503;
															assign node11503 = (inp[1]) ? 4'b1111 : 4'b1110;
															assign node11506 = (inp[0]) ? 4'b1111 : node11507;
																assign node11507 = (inp[1]) ? 4'b1110 : 4'b1111;
													assign node11511 = (inp[0]) ? node11519 : node11512;
														assign node11512 = (inp[10]) ? node11516 : node11513;
															assign node11513 = (inp[9]) ? 4'b1111 : 4'b1110;
															assign node11516 = (inp[9]) ? 4'b1110 : 4'b1111;
														assign node11519 = (inp[10]) ? node11527 : node11520;
															assign node11520 = (inp[1]) ? node11524 : node11521;
																assign node11521 = (inp[9]) ? 4'b1110 : 4'b1111;
																assign node11524 = (inp[9]) ? 4'b1111 : 4'b1110;
															assign node11527 = (inp[1]) ? node11531 : node11528;
																assign node11528 = (inp[9]) ? 4'b1111 : 4'b1110;
																assign node11531 = (inp[9]) ? 4'b1110 : 4'b1111;
											assign node11534 = (inp[4]) ? node11578 : node11535;
												assign node11535 = (inp[9]) ? node11557 : node11536;
													assign node11536 = (inp[0]) ? node11544 : node11537;
														assign node11537 = (inp[1]) ? node11541 : node11538;
															assign node11538 = (inp[10]) ? 4'b1101 : 4'b1100;
															assign node11541 = (inp[10]) ? 4'b1100 : 4'b1101;
														assign node11544 = (inp[1]) ? node11552 : node11545;
															assign node11545 = (inp[10]) ? node11549 : node11546;
																assign node11546 = (inp[11]) ? 4'b1100 : 4'b1101;
																assign node11549 = (inp[11]) ? 4'b1101 : 4'b1100;
															assign node11552 = (inp[10]) ? 4'b1100 : node11553;
																assign node11553 = (inp[11]) ? 4'b1101 : 4'b1100;
													assign node11557 = (inp[11]) ? node11571 : node11558;
														assign node11558 = (inp[10]) ? node11564 : node11559;
															assign node11559 = (inp[0]) ? 4'b1100 : node11560;
																assign node11560 = (inp[1]) ? 4'b1100 : 4'b1101;
															assign node11564 = (inp[1]) ? node11568 : node11565;
																assign node11565 = (inp[0]) ? 4'b1101 : 4'b1100;
																assign node11568 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node11571 = (inp[1]) ? node11575 : node11572;
															assign node11572 = (inp[10]) ? 4'b1100 : 4'b1101;
															assign node11575 = (inp[10]) ? 4'b1101 : 4'b1100;
												assign node11578 = (inp[1]) ? node11600 : node11579;
													assign node11579 = (inp[0]) ? node11587 : node11580;
														assign node11580 = (inp[10]) ? node11584 : node11581;
															assign node11581 = (inp[9]) ? 4'b1001 : 4'b1000;
															assign node11584 = (inp[9]) ? 4'b1000 : 4'b1001;
														assign node11587 = (inp[10]) ? node11595 : node11588;
															assign node11588 = (inp[9]) ? node11592 : node11589;
																assign node11589 = (inp[11]) ? 4'b1000 : 4'b1001;
																assign node11592 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node11595 = (inp[9]) ? node11597 : 4'b1000;
																assign node11597 = (inp[11]) ? 4'b1000 : 4'b1001;
													assign node11600 = (inp[11]) ? node11608 : node11601;
														assign node11601 = (inp[10]) ? node11603 : 4'b1000;
															assign node11603 = (inp[9]) ? node11605 : 4'b1000;
																assign node11605 = (inp[0]) ? 4'b1000 : 4'b1001;
														assign node11608 = (inp[10]) ? node11612 : node11609;
															assign node11609 = (inp[9]) ? 4'b1000 : 4'b1001;
															assign node11612 = (inp[9]) ? 4'b1001 : 4'b1000;
										assign node11615 = (inp[4]) ? node11707 : node11616;
											assign node11616 = (inp[11]) ? node11666 : node11617;
												assign node11617 = (inp[1]) ? node11645 : node11618;
													assign node11618 = (inp[15]) ? node11632 : node11619;
														assign node11619 = (inp[0]) ? node11625 : node11620;
															assign node11620 = (inp[10]) ? node11622 : 4'b1111;
																assign node11622 = (inp[9]) ? 4'b1110 : 4'b1111;
															assign node11625 = (inp[9]) ? node11629 : node11626;
																assign node11626 = (inp[10]) ? 4'b1110 : 4'b1111;
																assign node11629 = (inp[10]) ? 4'b1111 : 4'b1110;
														assign node11632 = (inp[0]) ? node11638 : node11633;
															assign node11633 = (inp[9]) ? node11635 : 4'b1110;
																assign node11635 = (inp[10]) ? 4'b1110 : 4'b1111;
															assign node11638 = (inp[10]) ? node11642 : node11639;
																assign node11639 = (inp[9]) ? 4'b1110 : 4'b1111;
																assign node11642 = (inp[9]) ? 4'b1111 : 4'b1110;
													assign node11645 = (inp[15]) ? node11653 : node11646;
														assign node11646 = (inp[10]) ? node11650 : node11647;
															assign node11647 = (inp[9]) ? 4'b1110 : 4'b1111;
															assign node11650 = (inp[9]) ? 4'b1111 : 4'b1110;
														assign node11653 = (inp[10]) ? node11659 : node11654;
															assign node11654 = (inp[9]) ? 4'b1110 : node11655;
																assign node11655 = (inp[0]) ? 4'b1111 : 4'b1110;
															assign node11659 = (inp[9]) ? node11663 : node11660;
																assign node11660 = (inp[0]) ? 4'b1110 : 4'b1111;
																assign node11663 = (inp[0]) ? 4'b1111 : 4'b1110;
												assign node11666 = (inp[1]) ? node11690 : node11667;
													assign node11667 = (inp[0]) ? node11683 : node11668;
														assign node11668 = (inp[15]) ? node11676 : node11669;
															assign node11669 = (inp[9]) ? node11673 : node11670;
																assign node11670 = (inp[10]) ? 4'b1111 : 4'b1110;
																assign node11673 = (inp[10]) ? 4'b1110 : 4'b1111;
															assign node11676 = (inp[10]) ? node11680 : node11677;
																assign node11677 = (inp[9]) ? 4'b1111 : 4'b1110;
																assign node11680 = (inp[9]) ? 4'b1110 : 4'b1111;
														assign node11683 = (inp[9]) ? node11687 : node11684;
															assign node11684 = (inp[10]) ? 4'b1111 : 4'b1110;
															assign node11687 = (inp[10]) ? 4'b1110 : 4'b1111;
													assign node11690 = (inp[10]) ? node11702 : node11691;
														assign node11691 = (inp[9]) ? node11697 : node11692;
															assign node11692 = (inp[15]) ? 4'b1110 : node11693;
																assign node11693 = (inp[0]) ? 4'b1111 : 4'b1110;
															assign node11697 = (inp[15]) ? 4'b1111 : node11698;
																assign node11698 = (inp[0]) ? 4'b1110 : 4'b1111;
														assign node11702 = (inp[9]) ? node11704 : 4'b1111;
															assign node11704 = (inp[0]) ? 4'b1111 : 4'b1110;
											assign node11707 = (inp[15]) ? node11755 : node11708;
												assign node11708 = (inp[1]) ? node11732 : node11709;
													assign node11709 = (inp[11]) ? node11725 : node11710;
														assign node11710 = (inp[0]) ? node11718 : node11711;
															assign node11711 = (inp[10]) ? node11715 : node11712;
																assign node11712 = (inp[9]) ? 4'b1101 : 4'b1100;
																assign node11715 = (inp[9]) ? 4'b1100 : 4'b1101;
															assign node11718 = (inp[9]) ? node11722 : node11719;
																assign node11719 = (inp[10]) ? 4'b1100 : 4'b1101;
																assign node11722 = (inp[10]) ? 4'b1101 : 4'b1100;
														assign node11725 = (inp[10]) ? node11729 : node11726;
															assign node11726 = (inp[9]) ? 4'b1101 : 4'b1100;
															assign node11729 = (inp[9]) ? 4'b1100 : 4'b1101;
													assign node11732 = (inp[0]) ? node11748 : node11733;
														assign node11733 = (inp[10]) ? node11741 : node11734;
															assign node11734 = (inp[9]) ? node11738 : node11735;
																assign node11735 = (inp[11]) ? 4'b1000 : 4'b1001;
																assign node11738 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node11741 = (inp[11]) ? node11745 : node11742;
																assign node11742 = (inp[9]) ? 4'b1001 : 4'b1000;
																assign node11745 = (inp[9]) ? 4'b1000 : 4'b1001;
														assign node11748 = (inp[9]) ? node11752 : node11749;
															assign node11749 = (inp[10]) ? 4'b1000 : 4'b1001;
															assign node11752 = (inp[10]) ? 4'b1001 : 4'b1000;
												assign node11755 = (inp[10]) ? node11765 : node11756;
													assign node11756 = (inp[9]) ? node11762 : node11757;
														assign node11757 = (inp[11]) ? 4'b1110 : node11758;
															assign node11758 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node11762 = (inp[11]) ? 4'b1111 : 4'b1110;
													assign node11765 = (inp[9]) ? node11771 : node11766;
														assign node11766 = (inp[0]) ? node11768 : 4'b1111;
															assign node11768 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node11771 = (inp[0]) ? node11773 : 4'b1110;
															assign node11773 = (inp[11]) ? 4'b1110 : 4'b1111;
									assign node11776 = (inp[12]) ? node11970 : node11777;
										assign node11777 = (inp[15]) ? node11861 : node11778;
											assign node11778 = (inp[4]) ? node11814 : node11779;
												assign node11779 = (inp[1]) ? node11801 : node11780;
													assign node11780 = (inp[0]) ? node11794 : node11781;
														assign node11781 = (inp[10]) ? node11787 : node11782;
															assign node11782 = (inp[9]) ? node11784 : 4'b1011;
																assign node11784 = (inp[11]) ? 4'b1011 : 4'b1010;
															assign node11787 = (inp[11]) ? node11791 : node11788;
																assign node11788 = (inp[9]) ? 4'b1011 : 4'b1010;
																assign node11791 = (inp[9]) ? 4'b1010 : 4'b1011;
														assign node11794 = (inp[9]) ? node11798 : node11795;
															assign node11795 = (inp[10]) ? 4'b1010 : 4'b1011;
															assign node11798 = (inp[10]) ? 4'b1011 : 4'b1010;
													assign node11801 = (inp[9]) ? node11809 : node11802;
														assign node11802 = (inp[10]) ? 4'b1110 : node11803;
															assign node11803 = (inp[0]) ? 4'b1111 : node11804;
																assign node11804 = (inp[11]) ? 4'b1110 : 4'b1111;
														assign node11809 = (inp[10]) ? 4'b1111 : node11810;
															assign node11810 = (inp[11]) ? 4'b1111 : 4'b1110;
												assign node11814 = (inp[10]) ? node11838 : node11815;
													assign node11815 = (inp[9]) ? node11827 : node11816;
														assign node11816 = (inp[1]) ? node11822 : node11817;
															assign node11817 = (inp[11]) ? 4'b1001 : node11818;
																assign node11818 = (inp[0]) ? 4'b1000 : 4'b1001;
															assign node11822 = (inp[11]) ? node11824 : 4'b1001;
																assign node11824 = (inp[0]) ? 4'b1001 : 4'b1000;
														assign node11827 = (inp[0]) ? node11833 : node11828;
															assign node11828 = (inp[1]) ? node11830 : 4'b1000;
																assign node11830 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node11833 = (inp[1]) ? 4'b1000 : node11834;
																assign node11834 = (inp[11]) ? 4'b1000 : 4'b1001;
													assign node11838 = (inp[9]) ? node11850 : node11839;
														assign node11839 = (inp[0]) ? node11845 : node11840;
															assign node11840 = (inp[11]) ? node11842 : 4'b1000;
																assign node11842 = (inp[1]) ? 4'b1001 : 4'b1000;
															assign node11845 = (inp[11]) ? 4'b1000 : node11846;
																assign node11846 = (inp[1]) ? 4'b1000 : 4'b1001;
														assign node11850 = (inp[11]) ? node11856 : node11851;
															assign node11851 = (inp[1]) ? 4'b1001 : node11852;
																assign node11852 = (inp[0]) ? 4'b1000 : 4'b1001;
															assign node11856 = (inp[0]) ? 4'b1001 : node11857;
																assign node11857 = (inp[1]) ? 4'b1000 : 4'b1001;
											assign node11861 = (inp[11]) ? node11921 : node11862;
												assign node11862 = (inp[0]) ? node11890 : node11863;
													assign node11863 = (inp[9]) ? node11877 : node11864;
														assign node11864 = (inp[1]) ? node11870 : node11865;
															assign node11865 = (inp[10]) ? node11867 : 4'b1011;
																assign node11867 = (inp[4]) ? 4'b1010 : 4'b1110;
															assign node11870 = (inp[10]) ? node11874 : node11871;
																assign node11871 = (inp[4]) ? 4'b1110 : 4'b1010;
																assign node11874 = (inp[4]) ? 4'b1111 : 4'b1011;
														assign node11877 = (inp[10]) ? node11885 : node11878;
															assign node11878 = (inp[1]) ? node11882 : node11879;
																assign node11879 = (inp[4]) ? 4'b1010 : 4'b1110;
																assign node11882 = (inp[4]) ? 4'b1111 : 4'b1011;
															assign node11885 = (inp[1]) ? 4'b1010 : node11886;
																assign node11886 = (inp[4]) ? 4'b1011 : 4'b1111;
													assign node11890 = (inp[10]) ? node11906 : node11891;
														assign node11891 = (inp[9]) ? node11899 : node11892;
															assign node11892 = (inp[1]) ? node11896 : node11893;
																assign node11893 = (inp[4]) ? 4'b1011 : 4'b1111;
																assign node11896 = (inp[4]) ? 4'b1111 : 4'b1010;
															assign node11899 = (inp[4]) ? node11903 : node11900;
																assign node11900 = (inp[1]) ? 4'b1011 : 4'b1110;
																assign node11903 = (inp[1]) ? 4'b1110 : 4'b1010;
														assign node11906 = (inp[9]) ? node11914 : node11907;
															assign node11907 = (inp[4]) ? node11911 : node11908;
																assign node11908 = (inp[1]) ? 4'b1011 : 4'b1110;
																assign node11911 = (inp[1]) ? 4'b1110 : 4'b1010;
															assign node11914 = (inp[4]) ? node11918 : node11915;
																assign node11915 = (inp[1]) ? 4'b1010 : 4'b1111;
																assign node11918 = (inp[1]) ? 4'b1111 : 4'b1011;
												assign node11921 = (inp[4]) ? node11945 : node11922;
													assign node11922 = (inp[1]) ? node11938 : node11923;
														assign node11923 = (inp[10]) ? node11931 : node11924;
															assign node11924 = (inp[0]) ? node11928 : node11925;
																assign node11925 = (inp[9]) ? 4'b1111 : 4'b1110;
																assign node11928 = (inp[9]) ? 4'b1110 : 4'b1111;
															assign node11931 = (inp[0]) ? node11935 : node11932;
																assign node11932 = (inp[9]) ? 4'b1110 : 4'b1111;
																assign node11935 = (inp[9]) ? 4'b1111 : 4'b1110;
														assign node11938 = (inp[9]) ? node11940 : 4'b1011;
															assign node11940 = (inp[10]) ? node11942 : 4'b1011;
																assign node11942 = (inp[0]) ? 4'b1010 : 4'b1011;
													assign node11945 = (inp[1]) ? node11957 : node11946;
														assign node11946 = (inp[10]) ? node11952 : node11947;
															assign node11947 = (inp[9]) ? 4'b1010 : node11948;
																assign node11948 = (inp[0]) ? 4'b1011 : 4'b1010;
															assign node11952 = (inp[0]) ? 4'b1011 : node11953;
																assign node11953 = (inp[9]) ? 4'b1010 : 4'b1011;
														assign node11957 = (inp[0]) ? node11963 : node11958;
															assign node11958 = (inp[9]) ? node11960 : 4'b1110;
																assign node11960 = (inp[10]) ? 4'b1110 : 4'b1111;
															assign node11963 = (inp[9]) ? node11967 : node11964;
																assign node11964 = (inp[10]) ? 4'b1111 : 4'b1110;
																assign node11967 = (inp[10]) ? 4'b1110 : 4'b1111;
										assign node11970 = (inp[15]) ? node12042 : node11971;
											assign node11971 = (inp[4]) ? node12009 : node11972;
												assign node11972 = (inp[9]) ? node11990 : node11973;
													assign node11973 = (inp[0]) ? node11983 : node11974;
														assign node11974 = (inp[10]) ? node11980 : node11975;
															assign node11975 = (inp[11]) ? 4'b1000 : node11976;
																assign node11976 = (inp[1]) ? 4'b1001 : 4'b1000;
															assign node11980 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node11983 = (inp[10]) ? 4'b1000 : node11984;
															assign node11984 = (inp[1]) ? 4'b1001 : node11985;
																assign node11985 = (inp[11]) ? 4'b1000 : 4'b1001;
													assign node11990 = (inp[10]) ? node11998 : node11991;
														assign node11991 = (inp[0]) ? node11993 : 4'b1001;
															assign node11993 = (inp[1]) ? 4'b1000 : node11994;
																assign node11994 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node11998 = (inp[0]) ? node12004 : node11999;
															assign node11999 = (inp[11]) ? 4'b1000 : node12000;
																assign node12000 = (inp[1]) ? 4'b1001 : 4'b1000;
															assign node12004 = (inp[11]) ? node12006 : 4'b1001;
																assign node12006 = (inp[1]) ? 4'b1001 : 4'b1000;
												assign node12009 = (inp[10]) ? node12027 : node12010;
													assign node12010 = (inp[9]) ? node12016 : node12011;
														assign node12011 = (inp[1]) ? node12013 : 4'b1111;
															assign node12013 = (inp[0]) ? 4'b1110 : 4'b1111;
														assign node12016 = (inp[11]) ? node12022 : node12017;
															assign node12017 = (inp[0]) ? node12019 : 4'b1110;
																assign node12019 = (inp[1]) ? 4'b1111 : 4'b1110;
															assign node12022 = (inp[1]) ? 4'b1110 : node12023;
																assign node12023 = (inp[0]) ? 4'b1110 : 4'b1111;
													assign node12027 = (inp[9]) ? node12035 : node12028;
														assign node12028 = (inp[0]) ? node12032 : node12029;
															assign node12029 = (inp[11]) ? 4'b1111 : 4'b1110;
															assign node12032 = (inp[11]) ? 4'b1110 : 4'b1111;
														assign node12035 = (inp[0]) ? 4'b1111 : node12036;
															assign node12036 = (inp[1]) ? 4'b1111 : node12037;
																assign node12037 = (inp[11]) ? 4'b1110 : 4'b1111;
											assign node12042 = (inp[10]) ? node12054 : node12043;
												assign node12043 = (inp[9]) ? node12049 : node12044;
													assign node12044 = (inp[11]) ? 4'b1100 : node12045;
														assign node12045 = (inp[0]) ? 4'b1101 : 4'b1100;
													assign node12049 = (inp[0]) ? node12051 : 4'b1101;
														assign node12051 = (inp[11]) ? 4'b1101 : 4'b1100;
												assign node12054 = (inp[9]) ? node12060 : node12055;
													assign node12055 = (inp[0]) ? node12057 : 4'b1101;
														assign node12057 = (inp[11]) ? 4'b1101 : 4'b1100;
													assign node12060 = (inp[11]) ? 4'b1100 : node12061;
														assign node12061 = (inp[0]) ? 4'b1101 : 4'b1100;
							assign node12065 = (inp[12]) ? node12575 : node12066;
								assign node12066 = (inp[15]) ? node12282 : node12067;
									assign node12067 = (inp[7]) ? node12187 : node12068;
										assign node12068 = (inp[4]) ? node12122 : node12069;
											assign node12069 = (inp[1]) ? node12101 : node12070;
												assign node12070 = (inp[2]) ? node12094 : node12071;
													assign node12071 = (inp[11]) ? node12081 : node12072;
														assign node12072 = (inp[10]) ? node12074 : 4'b1101;
															assign node12074 = (inp[0]) ? node12078 : node12075;
																assign node12075 = (inp[9]) ? 4'b1101 : 4'b1100;
																assign node12078 = (inp[9]) ? 4'b1100 : 4'b1101;
														assign node12081 = (inp[10]) ? node12087 : node12082;
															assign node12082 = (inp[0]) ? node12084 : 4'b1100;
																assign node12084 = (inp[9]) ? 4'b1101 : 4'b1100;
															assign node12087 = (inp[9]) ? node12091 : node12088;
																assign node12088 = (inp[0]) ? 4'b1100 : 4'b1101;
																assign node12091 = (inp[0]) ? 4'b1101 : 4'b1100;
													assign node12094 = (inp[11]) ? node12098 : node12095;
														assign node12095 = (inp[9]) ? 4'b1101 : 4'b1100;
														assign node12098 = (inp[9]) ? 4'b1100 : 4'b1101;
												assign node12101 = (inp[9]) ? node12111 : node12102;
													assign node12102 = (inp[11]) ? node12108 : node12103;
														assign node12103 = (inp[0]) ? 4'b1000 : node12104;
															assign node12104 = (inp[2]) ? 4'b1001 : 4'b1000;
														assign node12108 = (inp[2]) ? 4'b1000 : 4'b1001;
													assign node12111 = (inp[11]) ? node12117 : node12112;
														assign node12112 = (inp[0]) ? 4'b1001 : node12113;
															assign node12113 = (inp[2]) ? 4'b1000 : 4'b1001;
														assign node12117 = (inp[0]) ? 4'b1000 : node12118;
															assign node12118 = (inp[2]) ? 4'b1001 : 4'b1000;
											assign node12122 = (inp[2]) ? node12146 : node12123;
												assign node12123 = (inp[9]) ? node12135 : node12124;
													assign node12124 = (inp[11]) ? node12130 : node12125;
														assign node12125 = (inp[0]) ? 4'b1100 : node12126;
															assign node12126 = (inp[1]) ? 4'b1101 : 4'b1100;
														assign node12130 = (inp[1]) ? node12132 : 4'b1101;
															assign node12132 = (inp[0]) ? 4'b1101 : 4'b1100;
													assign node12135 = (inp[11]) ? node12141 : node12136;
														assign node12136 = (inp[1]) ? node12138 : 4'b1101;
															assign node12138 = (inp[0]) ? 4'b1101 : 4'b1100;
														assign node12141 = (inp[1]) ? node12143 : 4'b1100;
															assign node12143 = (inp[0]) ? 4'b1100 : 4'b1101;
												assign node12146 = (inp[10]) ? node12164 : node12147;
													assign node12147 = (inp[11]) ? node12159 : node12148;
														assign node12148 = (inp[9]) ? node12154 : node12149;
															assign node12149 = (inp[0]) ? node12151 : 4'b1100;
																assign node12151 = (inp[1]) ? 4'b1100 : 4'b1101;
															assign node12154 = (inp[1]) ? 4'b1101 : node12155;
																assign node12155 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node12159 = (inp[9]) ? 4'b1100 : node12160;
															assign node12160 = (inp[0]) ? 4'b1100 : 4'b1101;
													assign node12164 = (inp[11]) ? node12176 : node12165;
														assign node12165 = (inp[9]) ? node12171 : node12166;
															assign node12166 = (inp[1]) ? 4'b1100 : node12167;
																assign node12167 = (inp[0]) ? 4'b1101 : 4'b1100;
															assign node12171 = (inp[0]) ? node12173 : 4'b1101;
																assign node12173 = (inp[1]) ? 4'b1101 : 4'b1100;
														assign node12176 = (inp[9]) ? node12182 : node12177;
															assign node12177 = (inp[0]) ? node12179 : 4'b1101;
																assign node12179 = (inp[1]) ? 4'b1101 : 4'b1100;
															assign node12182 = (inp[1]) ? 4'b1100 : node12183;
																assign node12183 = (inp[0]) ? 4'b1101 : 4'b1100;
										assign node12187 = (inp[4]) ? node12235 : node12188;
											assign node12188 = (inp[0]) ? node12212 : node12189;
												assign node12189 = (inp[11]) ? node12201 : node12190;
													assign node12190 = (inp[9]) ? node12196 : node12191;
														assign node12191 = (inp[1]) ? node12193 : 4'b1111;
															assign node12193 = (inp[2]) ? 4'b1110 : 4'b1111;
														assign node12196 = (inp[2]) ? node12198 : 4'b1110;
															assign node12198 = (inp[1]) ? 4'b1111 : 4'b1110;
													assign node12201 = (inp[9]) ? node12207 : node12202;
														assign node12202 = (inp[1]) ? node12204 : 4'b1110;
															assign node12204 = (inp[2]) ? 4'b1111 : 4'b1110;
														assign node12207 = (inp[2]) ? node12209 : 4'b1111;
															assign node12209 = (inp[1]) ? 4'b1110 : 4'b1111;
												assign node12212 = (inp[9]) ? node12224 : node12213;
													assign node12213 = (inp[11]) ? node12219 : node12214;
														assign node12214 = (inp[2]) ? 4'b1111 : node12215;
															assign node12215 = (inp[1]) ? 4'b1111 : 4'b1110;
														assign node12219 = (inp[1]) ? 4'b1110 : node12220;
															assign node12220 = (inp[2]) ? 4'b1110 : 4'b1111;
													assign node12224 = (inp[11]) ? node12230 : node12225;
														assign node12225 = (inp[2]) ? 4'b1110 : node12226;
															assign node12226 = (inp[1]) ? 4'b1110 : 4'b1111;
														assign node12230 = (inp[2]) ? 4'b1111 : node12231;
															assign node12231 = (inp[1]) ? 4'b1111 : 4'b1110;
											assign node12235 = (inp[1]) ? node12259 : node12236;
												assign node12236 = (inp[9]) ? node12248 : node12237;
													assign node12237 = (inp[11]) ? node12243 : node12238;
														assign node12238 = (inp[0]) ? 4'b1011 : node12239;
															assign node12239 = (inp[2]) ? 4'b1011 : 4'b1010;
														assign node12243 = (inp[0]) ? 4'b1010 : node12244;
															assign node12244 = (inp[2]) ? 4'b1010 : 4'b1011;
													assign node12248 = (inp[11]) ? node12254 : node12249;
														assign node12249 = (inp[2]) ? 4'b1010 : node12250;
															assign node12250 = (inp[0]) ? 4'b1010 : 4'b1011;
														assign node12254 = (inp[0]) ? 4'b1011 : node12255;
															assign node12255 = (inp[2]) ? 4'b1011 : 4'b1010;
												assign node12259 = (inp[0]) ? node12275 : node12260;
													assign node12260 = (inp[9]) ? node12268 : node12261;
														assign node12261 = (inp[10]) ? 4'b1111 : node12262;
															assign node12262 = (inp[2]) ? node12264 : 4'b1111;
																assign node12264 = (inp[11]) ? 4'b1110 : 4'b1111;
														assign node12268 = (inp[11]) ? node12272 : node12269;
															assign node12269 = (inp[2]) ? 4'b1110 : 4'b1111;
															assign node12272 = (inp[2]) ? 4'b1111 : 4'b1110;
													assign node12275 = (inp[9]) ? node12279 : node12276;
														assign node12276 = (inp[11]) ? 4'b1110 : 4'b1111;
														assign node12279 = (inp[11]) ? 4'b1111 : 4'b1110;
									assign node12282 = (inp[7]) ? node12484 : node12283;
										assign node12283 = (inp[0]) ? node12381 : node12284;
											assign node12284 = (inp[2]) ? node12332 : node12285;
												assign node12285 = (inp[10]) ? node12307 : node12286;
													assign node12286 = (inp[4]) ? node12298 : node12287;
														assign node12287 = (inp[1]) ? node12293 : node12288;
															assign node12288 = (inp[9]) ? 4'b1111 : node12289;
																assign node12289 = (inp[11]) ? 4'b1111 : 4'b1110;
															assign node12293 = (inp[9]) ? 4'b1010 : node12294;
																assign node12294 = (inp[11]) ? 4'b1010 : 4'b1011;
														assign node12298 = (inp[1]) ? 4'b1111 : node12299;
															assign node12299 = (inp[11]) ? node12303 : node12300;
																assign node12300 = (inp[9]) ? 4'b1010 : 4'b1011;
																assign node12303 = (inp[9]) ? 4'b1011 : 4'b1010;
													assign node12307 = (inp[1]) ? node12321 : node12308;
														assign node12308 = (inp[4]) ? node12314 : node12309;
															assign node12309 = (inp[9]) ? node12311 : 4'b1111;
																assign node12311 = (inp[11]) ? 4'b1110 : 4'b1111;
															assign node12314 = (inp[9]) ? node12318 : node12315;
																assign node12315 = (inp[11]) ? 4'b1010 : 4'b1011;
																assign node12318 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node12321 = (inp[4]) ? node12325 : node12322;
															assign node12322 = (inp[9]) ? 4'b1011 : 4'b1010;
															assign node12325 = (inp[9]) ? node12329 : node12326;
																assign node12326 = (inp[11]) ? 4'b1110 : 4'b1111;
																assign node12329 = (inp[11]) ? 4'b1111 : 4'b1110;
												assign node12332 = (inp[10]) ? node12362 : node12333;
													assign node12333 = (inp[11]) ? node12347 : node12334;
														assign node12334 = (inp[1]) ? node12340 : node12335;
															assign node12335 = (inp[4]) ? node12337 : 4'b1110;
																assign node12337 = (inp[9]) ? 4'b1011 : 4'b1010;
															assign node12340 = (inp[4]) ? node12344 : node12341;
																assign node12341 = (inp[9]) ? 4'b1010 : 4'b1011;
																assign node12344 = (inp[9]) ? 4'b1110 : 4'b1111;
														assign node12347 = (inp[4]) ? node12355 : node12348;
															assign node12348 = (inp[1]) ? node12352 : node12349;
																assign node12349 = (inp[9]) ? 4'b1110 : 4'b1111;
																assign node12352 = (inp[9]) ? 4'b1011 : 4'b1010;
															assign node12355 = (inp[1]) ? node12359 : node12356;
																assign node12356 = (inp[9]) ? 4'b1010 : 4'b1011;
																assign node12359 = (inp[9]) ? 4'b1111 : 4'b1110;
													assign node12362 = (inp[9]) ? node12376 : node12363;
														assign node12363 = (inp[4]) ? node12371 : node12364;
															assign node12364 = (inp[1]) ? node12368 : node12365;
																assign node12365 = (inp[11]) ? 4'b1111 : 4'b1110;
																assign node12368 = (inp[11]) ? 4'b1010 : 4'b1011;
															assign node12371 = (inp[1]) ? 4'b1111 : node12372;
																assign node12372 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node12376 = (inp[4]) ? 4'b1011 : node12377;
															assign node12377 = (inp[11]) ? 4'b1011 : 4'b1010;
											assign node12381 = (inp[10]) ? node12429 : node12382;
												assign node12382 = (inp[11]) ? node12404 : node12383;
													assign node12383 = (inp[2]) ? node12397 : node12384;
														assign node12384 = (inp[4]) ? node12390 : node12385;
															assign node12385 = (inp[1]) ? 4'b1011 : node12386;
																assign node12386 = (inp[9]) ? 4'b1110 : 4'b1111;
															assign node12390 = (inp[1]) ? node12394 : node12391;
																assign node12391 = (inp[9]) ? 4'b1011 : 4'b1010;
																assign node12394 = (inp[9]) ? 4'b1110 : 4'b1111;
														assign node12397 = (inp[9]) ? node12399 : 4'b1110;
															assign node12399 = (inp[1]) ? node12401 : 4'b1111;
																assign node12401 = (inp[4]) ? 4'b1111 : 4'b1010;
													assign node12404 = (inp[9]) ? node12418 : node12405;
														assign node12405 = (inp[1]) ? node12411 : node12406;
															assign node12406 = (inp[4]) ? 4'b1011 : node12407;
																assign node12407 = (inp[2]) ? 4'b1111 : 4'b1110;
															assign node12411 = (inp[4]) ? node12415 : node12412;
																assign node12412 = (inp[2]) ? 4'b1010 : 4'b1011;
																assign node12415 = (inp[2]) ? 4'b1111 : 4'b1110;
														assign node12418 = (inp[1]) ? node12424 : node12419;
															assign node12419 = (inp[4]) ? 4'b1010 : node12420;
																assign node12420 = (inp[2]) ? 4'b1110 : 4'b1111;
															assign node12424 = (inp[4]) ? node12426 : 4'b1011;
																assign node12426 = (inp[2]) ? 4'b1110 : 4'b1111;
												assign node12429 = (inp[1]) ? node12453 : node12430;
													assign node12430 = (inp[4]) ? node12446 : node12431;
														assign node12431 = (inp[11]) ? node12439 : node12432;
															assign node12432 = (inp[9]) ? node12436 : node12433;
																assign node12433 = (inp[2]) ? 4'b1110 : 4'b1111;
																assign node12436 = (inp[2]) ? 4'b1111 : 4'b1110;
															assign node12439 = (inp[9]) ? node12443 : node12440;
																assign node12440 = (inp[2]) ? 4'b1111 : 4'b1110;
																assign node12443 = (inp[2]) ? 4'b1110 : 4'b1111;
														assign node12446 = (inp[11]) ? node12450 : node12447;
															assign node12447 = (inp[9]) ? 4'b1011 : 4'b1010;
															assign node12450 = (inp[9]) ? 4'b1010 : 4'b1011;
													assign node12453 = (inp[4]) ? node12469 : node12454;
														assign node12454 = (inp[9]) ? node12462 : node12455;
															assign node12455 = (inp[2]) ? node12459 : node12456;
																assign node12456 = (inp[11]) ? 4'b1011 : 4'b1010;
																assign node12459 = (inp[11]) ? 4'b1010 : 4'b1011;
															assign node12462 = (inp[2]) ? node12466 : node12463;
																assign node12463 = (inp[11]) ? 4'b1010 : 4'b1011;
																assign node12466 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node12469 = (inp[11]) ? node12477 : node12470;
															assign node12470 = (inp[9]) ? node12474 : node12471;
																assign node12471 = (inp[2]) ? 4'b1110 : 4'b1111;
																assign node12474 = (inp[2]) ? 4'b1111 : 4'b1110;
															assign node12477 = (inp[9]) ? node12481 : node12478;
																assign node12478 = (inp[2]) ? 4'b1111 : 4'b1110;
																assign node12481 = (inp[2]) ? 4'b1110 : 4'b1111;
										assign node12484 = (inp[0]) ? node12538 : node12485;
											assign node12485 = (inp[11]) ? node12511 : node12486;
												assign node12486 = (inp[9]) ? node12500 : node12487;
													assign node12487 = (inp[1]) ? node12493 : node12488;
														assign node12488 = (inp[4]) ? 4'b1000 : node12489;
															assign node12489 = (inp[2]) ? 4'b1100 : 4'b1101;
														assign node12493 = (inp[4]) ? node12497 : node12494;
															assign node12494 = (inp[2]) ? 4'b1001 : 4'b1000;
															assign node12497 = (inp[2]) ? 4'b1100 : 4'b1101;
													assign node12500 = (inp[2]) ? node12506 : node12501;
														assign node12501 = (inp[1]) ? 4'b1100 : node12502;
															assign node12502 = (inp[4]) ? 4'b1001 : 4'b1100;
														assign node12506 = (inp[4]) ? node12508 : 4'b1101;
															assign node12508 = (inp[1]) ? 4'b1101 : 4'b1001;
												assign node12511 = (inp[9]) ? node12525 : node12512;
													assign node12512 = (inp[2]) ? node12518 : node12513;
														assign node12513 = (inp[4]) ? 4'b1100 : node12514;
															assign node12514 = (inp[1]) ? 4'b1001 : 4'b1100;
														assign node12518 = (inp[4]) ? node12522 : node12519;
															assign node12519 = (inp[1]) ? 4'b1000 : 4'b1101;
															assign node12522 = (inp[1]) ? 4'b1101 : 4'b1001;
													assign node12525 = (inp[4]) ? node12533 : node12526;
														assign node12526 = (inp[1]) ? node12530 : node12527;
															assign node12527 = (inp[2]) ? 4'b1100 : 4'b1101;
															assign node12530 = (inp[2]) ? 4'b1001 : 4'b1000;
														assign node12533 = (inp[1]) ? node12535 : 4'b1000;
															assign node12535 = (inp[2]) ? 4'b1100 : 4'b1101;
											assign node12538 = (inp[9]) ? node12556 : node12539;
												assign node12539 = (inp[11]) ? node12549 : node12540;
													assign node12540 = (inp[1]) ? node12546 : node12541;
														assign node12541 = (inp[4]) ? node12543 : 4'b1101;
															assign node12543 = (inp[2]) ? 4'b1001 : 4'b1000;
														assign node12546 = (inp[4]) ? 4'b1100 : 4'b1000;
													assign node12549 = (inp[1]) ? node12553 : node12550;
														assign node12550 = (inp[4]) ? 4'b1001 : 4'b1100;
														assign node12553 = (inp[4]) ? 4'b1101 : 4'b1001;
												assign node12556 = (inp[11]) ? node12566 : node12557;
													assign node12557 = (inp[1]) ? node12563 : node12558;
														assign node12558 = (inp[4]) ? node12560 : 4'b1100;
															assign node12560 = (inp[2]) ? 4'b1000 : 4'b1001;
														assign node12563 = (inp[4]) ? 4'b1101 : 4'b1001;
													assign node12566 = (inp[1]) ? node12572 : node12567;
														assign node12567 = (inp[4]) ? node12569 : 4'b1101;
															assign node12569 = (inp[2]) ? 4'b1001 : 4'b1000;
														assign node12572 = (inp[4]) ? 4'b1100 : 4'b1000;
								assign node12575 = (inp[15]) ? node12839 : node12576;
									assign node12576 = (inp[7]) ? node12708 : node12577;
										assign node12577 = (inp[1]) ? node12633 : node12578;
											assign node12578 = (inp[9]) ? node12614 : node12579;
												assign node12579 = (inp[11]) ? node12597 : node12580;
													assign node12580 = (inp[2]) ? 4'b1100 : node12581;
														assign node12581 = (inp[10]) ? node12589 : node12582;
															assign node12582 = (inp[4]) ? node12586 : node12583;
																assign node12583 = (inp[0]) ? 4'b1101 : 4'b1100;
																assign node12586 = (inp[0]) ? 4'b1100 : 4'b1101;
															assign node12589 = (inp[0]) ? node12593 : node12590;
																assign node12590 = (inp[4]) ? 4'b1101 : 4'b1100;
																assign node12593 = (inp[4]) ? 4'b1100 : 4'b1101;
													assign node12597 = (inp[2]) ? 4'b1101 : node12598;
														assign node12598 = (inp[10]) ? node12606 : node12599;
															assign node12599 = (inp[4]) ? node12603 : node12600;
																assign node12600 = (inp[0]) ? 4'b1100 : 4'b1101;
																assign node12603 = (inp[0]) ? 4'b1101 : 4'b1100;
															assign node12606 = (inp[4]) ? node12610 : node12607;
																assign node12607 = (inp[0]) ? 4'b1100 : 4'b1101;
																assign node12610 = (inp[0]) ? 4'b1101 : 4'b1100;
												assign node12614 = (inp[11]) ? node12624 : node12615;
													assign node12615 = (inp[2]) ? 4'b1101 : node12616;
														assign node12616 = (inp[4]) ? node12620 : node12617;
															assign node12617 = (inp[0]) ? 4'b1100 : 4'b1101;
															assign node12620 = (inp[0]) ? 4'b1101 : 4'b1100;
													assign node12624 = (inp[2]) ? 4'b1100 : node12625;
														assign node12625 = (inp[4]) ? node12629 : node12626;
															assign node12626 = (inp[0]) ? 4'b1101 : 4'b1100;
															assign node12629 = (inp[0]) ? 4'b1100 : 4'b1101;
											assign node12633 = (inp[4]) ? node12657 : node12634;
												assign node12634 = (inp[11]) ? node12646 : node12635;
													assign node12635 = (inp[9]) ? node12641 : node12636;
														assign node12636 = (inp[2]) ? node12638 : 4'b1101;
															assign node12638 = (inp[0]) ? 4'b1101 : 4'b1100;
														assign node12641 = (inp[2]) ? node12643 : 4'b1100;
															assign node12643 = (inp[0]) ? 4'b1100 : 4'b1101;
													assign node12646 = (inp[9]) ? node12652 : node12647;
														assign node12647 = (inp[2]) ? node12649 : 4'b1100;
															assign node12649 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node12652 = (inp[0]) ? 4'b1101 : node12653;
															assign node12653 = (inp[2]) ? 4'b1100 : 4'b1101;
												assign node12657 = (inp[10]) ? node12687 : node12658;
													assign node12658 = (inp[0]) ? node12672 : node12659;
														assign node12659 = (inp[2]) ? node12665 : node12660;
															assign node12660 = (inp[11]) ? 4'b1000 : node12661;
																assign node12661 = (inp[9]) ? 4'b1001 : 4'b1000;
															assign node12665 = (inp[11]) ? node12669 : node12666;
																assign node12666 = (inp[9]) ? 4'b1001 : 4'b1000;
																assign node12669 = (inp[9]) ? 4'b1000 : 4'b1001;
														assign node12672 = (inp[9]) ? node12680 : node12673;
															assign node12673 = (inp[11]) ? node12677 : node12674;
																assign node12674 = (inp[2]) ? 4'b1001 : 4'b1000;
																assign node12677 = (inp[2]) ? 4'b1000 : 4'b1001;
															assign node12680 = (inp[2]) ? node12684 : node12681;
																assign node12681 = (inp[11]) ? 4'b1000 : 4'b1001;
																assign node12684 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node12687 = (inp[11]) ? node12697 : node12688;
														assign node12688 = (inp[2]) ? node12690 : 4'b1001;
															assign node12690 = (inp[0]) ? node12694 : node12691;
																assign node12691 = (inp[9]) ? 4'b1001 : 4'b1000;
																assign node12694 = (inp[9]) ? 4'b1000 : 4'b1001;
														assign node12697 = (inp[9]) ? node12703 : node12698;
															assign node12698 = (inp[2]) ? node12700 : 4'b1001;
																assign node12700 = (inp[0]) ? 4'b1000 : 4'b1001;
															assign node12703 = (inp[0]) ? node12705 : 4'b1000;
																assign node12705 = (inp[2]) ? 4'b1001 : 4'b1000;
										assign node12708 = (inp[1]) ? node12782 : node12709;
											assign node12709 = (inp[4]) ? node12745 : node12710;
												assign node12710 = (inp[2]) ? node12738 : node12711;
													assign node12711 = (inp[11]) ? node12727 : node12712;
														assign node12712 = (inp[10]) ? node12720 : node12713;
															assign node12713 = (inp[9]) ? node12717 : node12714;
																assign node12714 = (inp[0]) ? 4'b1011 : 4'b1010;
																assign node12717 = (inp[0]) ? 4'b1010 : 4'b1011;
															assign node12720 = (inp[0]) ? node12724 : node12721;
																assign node12721 = (inp[9]) ? 4'b1011 : 4'b1010;
																assign node12724 = (inp[9]) ? 4'b1010 : 4'b1011;
														assign node12727 = (inp[10]) ? node12733 : node12728;
															assign node12728 = (inp[0]) ? node12730 : 4'b1010;
																assign node12730 = (inp[9]) ? 4'b1011 : 4'b1010;
															assign node12733 = (inp[0]) ? 4'b1010 : node12734;
																assign node12734 = (inp[9]) ? 4'b1010 : 4'b1011;
													assign node12738 = (inp[11]) ? node12742 : node12739;
														assign node12739 = (inp[9]) ? 4'b1011 : 4'b1010;
														assign node12742 = (inp[9]) ? 4'b1010 : 4'b1011;
												assign node12745 = (inp[2]) ? node12753 : node12746;
													assign node12746 = (inp[9]) ? node12750 : node12747;
														assign node12747 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node12750 = (inp[11]) ? 4'b1110 : 4'b1111;
													assign node12753 = (inp[10]) ? node12769 : node12754;
														assign node12754 = (inp[0]) ? node12762 : node12755;
															assign node12755 = (inp[11]) ? node12759 : node12756;
																assign node12756 = (inp[9]) ? 4'b1111 : 4'b1110;
																assign node12759 = (inp[9]) ? 4'b1110 : 4'b1111;
															assign node12762 = (inp[11]) ? node12766 : node12763;
																assign node12763 = (inp[9]) ? 4'b1110 : 4'b1111;
																assign node12766 = (inp[9]) ? 4'b1111 : 4'b1110;
														assign node12769 = (inp[9]) ? node12777 : node12770;
															assign node12770 = (inp[0]) ? node12774 : node12771;
																assign node12771 = (inp[11]) ? 4'b1111 : 4'b1110;
																assign node12774 = (inp[11]) ? 4'b1110 : 4'b1111;
															assign node12777 = (inp[11]) ? 4'b1111 : node12778;
																assign node12778 = (inp[0]) ? 4'b1110 : 4'b1111;
											assign node12782 = (inp[0]) ? node12818 : node12783;
												assign node12783 = (inp[10]) ? node12803 : node12784;
													assign node12784 = (inp[11]) ? node12794 : node12785;
														assign node12785 = (inp[2]) ? 4'b1111 : node12786;
															assign node12786 = (inp[9]) ? node12790 : node12787;
																assign node12787 = (inp[4]) ? 4'b1110 : 4'b1111;
																assign node12790 = (inp[4]) ? 4'b1111 : 4'b1110;
														assign node12794 = (inp[9]) ? node12800 : node12795;
															assign node12795 = (inp[4]) ? node12797 : 4'b1110;
																assign node12797 = (inp[2]) ? 4'b1110 : 4'b1111;
															assign node12800 = (inp[4]) ? 4'b1110 : 4'b1111;
													assign node12803 = (inp[4]) ? node12811 : node12804;
														assign node12804 = (inp[11]) ? node12808 : node12805;
															assign node12805 = (inp[9]) ? 4'b1110 : 4'b1111;
															assign node12808 = (inp[9]) ? 4'b1111 : 4'b1110;
														assign node12811 = (inp[11]) ? node12813 : 4'b1110;
															assign node12813 = (inp[2]) ? node12815 : 4'b1110;
																assign node12815 = (inp[9]) ? 4'b1111 : 4'b1110;
												assign node12818 = (inp[9]) ? node12830 : node12819;
													assign node12819 = (inp[11]) ? node12825 : node12820;
														assign node12820 = (inp[4]) ? 4'b1111 : node12821;
															assign node12821 = (inp[2]) ? 4'b1111 : 4'b1110;
														assign node12825 = (inp[2]) ? 4'b1110 : node12826;
															assign node12826 = (inp[4]) ? 4'b1110 : 4'b1111;
													assign node12830 = (inp[11]) ? node12834 : node12831;
														assign node12831 = (inp[2]) ? 4'b1110 : 4'b1111;
														assign node12834 = (inp[2]) ? 4'b1111 : node12835;
															assign node12835 = (inp[4]) ? 4'b1111 : 4'b1110;
									assign node12839 = (inp[7]) ? node12981 : node12840;
										assign node12840 = (inp[1]) ? node12894 : node12841;
											assign node12841 = (inp[2]) ? node12887 : node12842;
												assign node12842 = (inp[9]) ? node12866 : node12843;
													assign node12843 = (inp[4]) ? node12851 : node12844;
														assign node12844 = (inp[0]) ? node12848 : node12845;
															assign node12845 = (inp[11]) ? 4'b1111 : 4'b1110;
															assign node12848 = (inp[11]) ? 4'b1110 : 4'b1111;
														assign node12851 = (inp[10]) ? node12859 : node12852;
															assign node12852 = (inp[0]) ? node12856 : node12853;
																assign node12853 = (inp[11]) ? 4'b1110 : 4'b1111;
																assign node12856 = (inp[11]) ? 4'b1111 : 4'b1110;
															assign node12859 = (inp[11]) ? node12863 : node12860;
																assign node12860 = (inp[0]) ? 4'b1110 : 4'b1111;
																assign node12863 = (inp[0]) ? 4'b1111 : 4'b1110;
													assign node12866 = (inp[10]) ? node12876 : node12867;
														assign node12867 = (inp[0]) ? node12869 : 4'b1111;
															assign node12869 = (inp[4]) ? node12873 : node12870;
																assign node12870 = (inp[11]) ? 4'b1111 : 4'b1110;
																assign node12873 = (inp[11]) ? 4'b1110 : 4'b1111;
														assign node12876 = (inp[0]) ? node12882 : node12877;
															assign node12877 = (inp[11]) ? node12879 : 4'b1110;
																assign node12879 = (inp[4]) ? 4'b1111 : 4'b1110;
															assign node12882 = (inp[4]) ? node12884 : 4'b1111;
																assign node12884 = (inp[11]) ? 4'b1110 : 4'b1111;
												assign node12887 = (inp[11]) ? node12891 : node12888;
													assign node12888 = (inp[9]) ? 4'b1111 : 4'b1110;
													assign node12891 = (inp[9]) ? 4'b1110 : 4'b1111;
											assign node12894 = (inp[0]) ? node12942 : node12895;
												assign node12895 = (inp[2]) ? node12927 : node12896;
													assign node12896 = (inp[10]) ? node12912 : node12897;
														assign node12897 = (inp[11]) ? node12905 : node12898;
															assign node12898 = (inp[9]) ? node12902 : node12899;
																assign node12899 = (inp[4]) ? 4'b1111 : 4'b1110;
																assign node12902 = (inp[4]) ? 4'b1110 : 4'b1111;
															assign node12905 = (inp[4]) ? node12909 : node12906;
																assign node12906 = (inp[9]) ? 4'b1110 : 4'b1111;
																assign node12909 = (inp[9]) ? 4'b1111 : 4'b1110;
														assign node12912 = (inp[4]) ? node12920 : node12913;
															assign node12913 = (inp[9]) ? node12917 : node12914;
																assign node12914 = (inp[11]) ? 4'b1111 : 4'b1110;
																assign node12917 = (inp[11]) ? 4'b1110 : 4'b1111;
															assign node12920 = (inp[11]) ? node12924 : node12921;
																assign node12921 = (inp[9]) ? 4'b1110 : 4'b1111;
																assign node12924 = (inp[9]) ? 4'b1111 : 4'b1110;
													assign node12927 = (inp[10]) ? node12935 : node12928;
														assign node12928 = (inp[9]) ? node12932 : node12929;
															assign node12929 = (inp[11]) ? 4'b1111 : 4'b1110;
															assign node12932 = (inp[11]) ? 4'b1110 : 4'b1111;
														assign node12935 = (inp[11]) ? node12939 : node12936;
															assign node12936 = (inp[9]) ? 4'b1111 : 4'b1110;
															assign node12939 = (inp[9]) ? 4'b1110 : 4'b1111;
												assign node12942 = (inp[2]) ? node12958 : node12943;
													assign node12943 = (inp[9]) ? node12951 : node12944;
														assign node12944 = (inp[11]) ? node12948 : node12945;
															assign node12945 = (inp[4]) ? 4'b1110 : 4'b1111;
															assign node12948 = (inp[4]) ? 4'b1111 : 4'b1110;
														assign node12951 = (inp[4]) ? node12955 : node12952;
															assign node12952 = (inp[11]) ? 4'b1111 : 4'b1110;
															assign node12955 = (inp[11]) ? 4'b1110 : 4'b1111;
													assign node12958 = (inp[4]) ? node12972 : node12959;
														assign node12959 = (inp[10]) ? node12965 : node12960;
															assign node12960 = (inp[11]) ? 4'b1110 : node12961;
																assign node12961 = (inp[9]) ? 4'b1111 : 4'b1110;
															assign node12965 = (inp[11]) ? node12969 : node12966;
																assign node12966 = (inp[9]) ? 4'b1111 : 4'b1110;
																assign node12969 = (inp[9]) ? 4'b1110 : 4'b1111;
														assign node12972 = (inp[10]) ? 4'b1110 : node12973;
															assign node12973 = (inp[11]) ? node12977 : node12974;
																assign node12974 = (inp[9]) ? 4'b1111 : 4'b1110;
																assign node12977 = (inp[9]) ? 4'b1110 : 4'b1111;
										assign node12981 = (inp[4]) ? node13051 : node12982;
											assign node12982 = (inp[2]) ? node13044 : node12983;
												assign node12983 = (inp[1]) ? node13015 : node12984;
													assign node12984 = (inp[9]) ? node13000 : node12985;
														assign node12985 = (inp[10]) ? node12993 : node12986;
															assign node12986 = (inp[0]) ? node12990 : node12987;
																assign node12987 = (inp[11]) ? 4'b1101 : 4'b1100;
																assign node12990 = (inp[11]) ? 4'b1100 : 4'b1101;
															assign node12993 = (inp[11]) ? node12997 : node12994;
																assign node12994 = (inp[0]) ? 4'b1101 : 4'b1100;
																assign node12997 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node13000 = (inp[10]) ? node13008 : node13001;
															assign node13001 = (inp[0]) ? node13005 : node13002;
																assign node13002 = (inp[11]) ? 4'b1100 : 4'b1101;
																assign node13005 = (inp[11]) ? 4'b1101 : 4'b1100;
															assign node13008 = (inp[0]) ? node13012 : node13009;
																assign node13009 = (inp[11]) ? 4'b1100 : 4'b1101;
																assign node13012 = (inp[11]) ? 4'b1101 : 4'b1100;
													assign node13015 = (inp[10]) ? node13031 : node13016;
														assign node13016 = (inp[9]) ? node13024 : node13017;
															assign node13017 = (inp[11]) ? node13021 : node13018;
																assign node13018 = (inp[0]) ? 4'b1101 : 4'b1100;
																assign node13021 = (inp[0]) ? 4'b1100 : 4'b1101;
															assign node13024 = (inp[0]) ? node13028 : node13025;
																assign node13025 = (inp[11]) ? 4'b1100 : 4'b1101;
																assign node13028 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node13031 = (inp[9]) ? node13039 : node13032;
															assign node13032 = (inp[0]) ? node13036 : node13033;
																assign node13033 = (inp[11]) ? 4'b1101 : 4'b1100;
																assign node13036 = (inp[11]) ? 4'b1100 : 4'b1101;
															assign node13039 = (inp[0]) ? 4'b1100 : node13040;
																assign node13040 = (inp[11]) ? 4'b1100 : 4'b1101;
												assign node13044 = (inp[9]) ? node13048 : node13045;
													assign node13045 = (inp[11]) ? 4'b1101 : 4'b1100;
													assign node13048 = (inp[11]) ? 4'b1100 : 4'b1101;
											assign node13051 = (inp[2]) ? node13103 : node13052;
												assign node13052 = (inp[1]) ? node13076 : node13053;
													assign node13053 = (inp[0]) ? node13061 : node13054;
														assign node13054 = (inp[9]) ? node13058 : node13055;
															assign node13055 = (inp[11]) ? 4'b1100 : 4'b1101;
															assign node13058 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node13061 = (inp[10]) ? node13069 : node13062;
															assign node13062 = (inp[11]) ? node13066 : node13063;
																assign node13063 = (inp[9]) ? 4'b1101 : 4'b1100;
																assign node13066 = (inp[9]) ? 4'b1100 : 4'b1101;
															assign node13069 = (inp[9]) ? node13073 : node13070;
																assign node13070 = (inp[11]) ? 4'b1101 : 4'b1100;
																assign node13073 = (inp[11]) ? 4'b1100 : 4'b1101;
													assign node13076 = (inp[0]) ? node13088 : node13077;
														assign node13077 = (inp[10]) ? node13083 : node13078;
															assign node13078 = (inp[9]) ? 4'b1100 : node13079;
																assign node13079 = (inp[11]) ? 4'b1100 : 4'b1101;
															assign node13083 = (inp[9]) ? node13085 : 4'b1100;
																assign node13085 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node13088 = (inp[10]) ? node13096 : node13089;
															assign node13089 = (inp[9]) ? node13093 : node13090;
																assign node13090 = (inp[11]) ? 4'b1101 : 4'b1100;
																assign node13093 = (inp[11]) ? 4'b1100 : 4'b1101;
															assign node13096 = (inp[11]) ? node13100 : node13097;
																assign node13097 = (inp[9]) ? 4'b1101 : 4'b1100;
																assign node13100 = (inp[9]) ? 4'b1100 : 4'b1101;
												assign node13103 = (inp[0]) ? node13111 : node13104;
													assign node13104 = (inp[11]) ? node13108 : node13105;
														assign node13105 = (inp[9]) ? 4'b1101 : 4'b1100;
														assign node13108 = (inp[9]) ? 4'b1100 : 4'b1101;
													assign node13111 = (inp[10]) ? node13121 : node13112;
														assign node13112 = (inp[1]) ? 4'b1100 : node13113;
															assign node13113 = (inp[9]) ? node13117 : node13114;
																assign node13114 = (inp[11]) ? 4'b1101 : 4'b1100;
																assign node13117 = (inp[11]) ? 4'b1100 : 4'b1101;
														assign node13121 = (inp[1]) ? node13127 : node13122;
															assign node13122 = (inp[9]) ? node13124 : 4'b1100;
																assign node13124 = (inp[11]) ? 4'b1100 : 4'b1101;
															assign node13127 = (inp[11]) ? node13131 : node13128;
																assign node13128 = (inp[9]) ? 4'b1101 : 4'b1100;
																assign node13131 = (inp[9]) ? 4'b1100 : 4'b1101;
					assign node13134 = (inp[5]) ? node15688 : node13135;
						assign node13135 = (inp[6]) ? node14695 : node13136;
							assign node13136 = (inp[0]) ? node13890 : node13137;
								assign node13137 = (inp[7]) ? node13501 : node13138;
									assign node13138 = (inp[12]) ? node13336 : node13139;
										assign node13139 = (inp[15]) ? node13227 : node13140;
											assign node13140 = (inp[4]) ? node13192 : node13141;
												assign node13141 = (inp[9]) ? node13169 : node13142;
													assign node13142 = (inp[10]) ? node13154 : node13143;
														assign node13143 = (inp[11]) ? node13149 : node13144;
															assign node13144 = (inp[1]) ? 4'b1001 : node13145;
																assign node13145 = (inp[2]) ? 4'b1001 : 4'b1100;
															assign node13149 = (inp[1]) ? 4'b1101 : node13150;
																assign node13150 = (inp[2]) ? 4'b1001 : 4'b1101;
														assign node13154 = (inp[11]) ? node13162 : node13155;
															assign node13155 = (inp[2]) ? node13159 : node13156;
																assign node13156 = (inp[1]) ? 4'b1000 : 4'b1101;
																assign node13159 = (inp[1]) ? 4'b1100 : 4'b1000;
															assign node13162 = (inp[1]) ? node13166 : node13163;
																assign node13163 = (inp[2]) ? 4'b1000 : 4'b1100;
																assign node13166 = (inp[2]) ? 4'b1100 : 4'b1000;
													assign node13169 = (inp[10]) ? node13183 : node13170;
														assign node13170 = (inp[11]) ? node13176 : node13171;
															assign node13171 = (inp[1]) ? node13173 : 4'b1101;
																assign node13173 = (inp[2]) ? 4'b1100 : 4'b1000;
															assign node13176 = (inp[2]) ? node13180 : node13177;
																assign node13177 = (inp[1]) ? 4'b1000 : 4'b1100;
																assign node13180 = (inp[1]) ? 4'b1100 : 4'b1000;
														assign node13183 = (inp[1]) ? node13189 : node13184;
															assign node13184 = (inp[2]) ? 4'b1001 : node13185;
																assign node13185 = (inp[11]) ? 4'b1101 : 4'b1100;
															assign node13189 = (inp[2]) ? 4'b1101 : 4'b1001;
												assign node13192 = (inp[9]) ? node13210 : node13193;
													assign node13193 = (inp[10]) ? node13201 : node13194;
														assign node13194 = (inp[2]) ? 4'b1110 : node13195;
															assign node13195 = (inp[1]) ? 4'b1011 : node13196;
																assign node13196 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node13201 = (inp[2]) ? node13207 : node13202;
															assign node13202 = (inp[1]) ? 4'b1010 : node13203;
																assign node13203 = (inp[11]) ? 4'b1110 : 4'b1111;
															assign node13207 = (inp[1]) ? 4'b1111 : 4'b1011;
													assign node13210 = (inp[1]) ? node13220 : node13211;
														assign node13211 = (inp[2]) ? node13217 : node13212;
															assign node13212 = (inp[11]) ? node13214 : 4'b1110;
																assign node13214 = (inp[10]) ? 4'b1111 : 4'b1110;
															assign node13217 = (inp[10]) ? 4'b1010 : 4'b1011;
														assign node13220 = (inp[2]) ? node13224 : node13221;
															assign node13221 = (inp[10]) ? 4'b1011 : 4'b1010;
															assign node13224 = (inp[10]) ? 4'b1110 : 4'b1111;
											assign node13227 = (inp[1]) ? node13275 : node13228;
												assign node13228 = (inp[2]) ? node13252 : node13229;
													assign node13229 = (inp[4]) ? node13245 : node13230;
														assign node13230 = (inp[10]) ? node13238 : node13231;
															assign node13231 = (inp[9]) ? node13235 : node13232;
																assign node13232 = (inp[11]) ? 4'b1100 : 4'b1101;
																assign node13235 = (inp[11]) ? 4'b1101 : 4'b1100;
															assign node13238 = (inp[9]) ? node13242 : node13239;
																assign node13239 = (inp[11]) ? 4'b1101 : 4'b1100;
																assign node13242 = (inp[11]) ? 4'b1100 : 4'b1101;
														assign node13245 = (inp[9]) ? node13249 : node13246;
															assign node13246 = (inp[10]) ? 4'b1001 : 4'b1000;
															assign node13249 = (inp[10]) ? 4'b1000 : 4'b1001;
													assign node13252 = (inp[4]) ? node13268 : node13253;
														assign node13253 = (inp[11]) ? node13261 : node13254;
															assign node13254 = (inp[9]) ? node13258 : node13255;
																assign node13255 = (inp[10]) ? 4'b1001 : 4'b1000;
																assign node13258 = (inp[10]) ? 4'b1000 : 4'b1001;
															assign node13261 = (inp[10]) ? node13265 : node13262;
																assign node13262 = (inp[9]) ? 4'b1001 : 4'b1000;
																assign node13265 = (inp[9]) ? 4'b1000 : 4'b1001;
														assign node13268 = (inp[10]) ? node13272 : node13269;
															assign node13269 = (inp[9]) ? 4'b1100 : 4'b1101;
															assign node13272 = (inp[9]) ? 4'b1101 : 4'b1100;
												assign node13275 = (inp[2]) ? node13307 : node13276;
													assign node13276 = (inp[4]) ? node13292 : node13277;
														assign node13277 = (inp[9]) ? node13285 : node13278;
															assign node13278 = (inp[11]) ? node13282 : node13279;
																assign node13279 = (inp[10]) ? 4'b1001 : 4'b1000;
																assign node13282 = (inp[10]) ? 4'b1000 : 4'b1001;
															assign node13285 = (inp[11]) ? node13289 : node13286;
																assign node13286 = (inp[10]) ? 4'b1000 : 4'b1001;
																assign node13289 = (inp[10]) ? 4'b1001 : 4'b1000;
														assign node13292 = (inp[10]) ? node13300 : node13293;
															assign node13293 = (inp[9]) ? node13297 : node13294;
																assign node13294 = (inp[11]) ? 4'b1101 : 4'b1100;
																assign node13297 = (inp[11]) ? 4'b1100 : 4'b1101;
															assign node13300 = (inp[11]) ? node13304 : node13301;
																assign node13301 = (inp[9]) ? 4'b1100 : 4'b1101;
																assign node13304 = (inp[9]) ? 4'b1101 : 4'b1100;
													assign node13307 = (inp[4]) ? node13323 : node13308;
														assign node13308 = (inp[11]) ? node13316 : node13309;
															assign node13309 = (inp[9]) ? node13313 : node13310;
																assign node13310 = (inp[10]) ? 4'b1101 : 4'b1100;
																assign node13313 = (inp[10]) ? 4'b1100 : 4'b1101;
															assign node13316 = (inp[10]) ? node13320 : node13317;
																assign node13317 = (inp[9]) ? 4'b1100 : 4'b1101;
																assign node13320 = (inp[9]) ? 4'b1101 : 4'b1100;
														assign node13323 = (inp[11]) ? node13331 : node13324;
															assign node13324 = (inp[9]) ? node13328 : node13325;
																assign node13325 = (inp[10]) ? 4'b1001 : 4'b1000;
																assign node13328 = (inp[10]) ? 4'b1000 : 4'b1001;
															assign node13331 = (inp[10]) ? node13333 : 4'b1000;
																assign node13333 = (inp[9]) ? 4'b1000 : 4'b1001;
										assign node13336 = (inp[15]) ? node13412 : node13337;
											assign node13337 = (inp[4]) ? node13369 : node13338;
												assign node13338 = (inp[1]) ? node13356 : node13339;
													assign node13339 = (inp[2]) ? node13349 : node13340;
														assign node13340 = (inp[10]) ? 4'b1110 : node13341;
															assign node13341 = (inp[11]) ? node13345 : node13342;
																assign node13342 = (inp[9]) ? 4'b1111 : 4'b1110;
																assign node13345 = (inp[9]) ? 4'b1110 : 4'b1111;
														assign node13349 = (inp[9]) ? node13353 : node13350;
															assign node13350 = (inp[10]) ? 4'b1010 : 4'b1011;
															assign node13353 = (inp[10]) ? 4'b1011 : 4'b1010;
													assign node13356 = (inp[2]) ? node13362 : node13357;
														assign node13357 = (inp[10]) ? 4'b1011 : node13358;
															assign node13358 = (inp[9]) ? 4'b1011 : 4'b1010;
														assign node13362 = (inp[10]) ? node13366 : node13363;
															assign node13363 = (inp[9]) ? 4'b1111 : 4'b1110;
															assign node13366 = (inp[9]) ? 4'b1110 : 4'b1111;
												assign node13369 = (inp[2]) ? node13393 : node13370;
													assign node13370 = (inp[11]) ? node13386 : node13371;
														assign node13371 = (inp[1]) ? node13379 : node13372;
															assign node13372 = (inp[9]) ? node13376 : node13373;
																assign node13373 = (inp[10]) ? 4'b1000 : 4'b1001;
																assign node13376 = (inp[10]) ? 4'b1001 : 4'b1000;
															assign node13379 = (inp[9]) ? node13383 : node13380;
																assign node13380 = (inp[10]) ? 4'b1001 : 4'b1000;
																assign node13383 = (inp[10]) ? 4'b1000 : 4'b1001;
														assign node13386 = (inp[9]) ? node13390 : node13387;
															assign node13387 = (inp[10]) ? 4'b1000 : 4'b1001;
															assign node13390 = (inp[10]) ? 4'b1001 : 4'b1000;
													assign node13393 = (inp[10]) ? node13403 : node13394;
														assign node13394 = (inp[9]) ? node13398 : node13395;
															assign node13395 = (inp[1]) ? 4'b1101 : 4'b1100;
															assign node13398 = (inp[1]) ? node13400 : 4'b1101;
																assign node13400 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node13403 = (inp[9]) ? node13407 : node13404;
															assign node13404 = (inp[1]) ? 4'b1100 : 4'b1101;
															assign node13407 = (inp[11]) ? 4'b1100 : node13408;
																assign node13408 = (inp[1]) ? 4'b1101 : 4'b1100;
											assign node13412 = (inp[10]) ? node13460 : node13413;
												assign node13413 = (inp[9]) ? node13435 : node13414;
													assign node13414 = (inp[11]) ? node13426 : node13415;
														assign node13415 = (inp[1]) ? node13421 : node13416;
															assign node13416 = (inp[2]) ? 4'b1010 : node13417;
																assign node13417 = (inp[4]) ? 4'b1110 : 4'b1111;
															assign node13421 = (inp[2]) ? 4'b1111 : node13422;
																assign node13422 = (inp[4]) ? 4'b1010 : 4'b1011;
														assign node13426 = (inp[1]) ? node13430 : node13427;
															assign node13427 = (inp[2]) ? 4'b1010 : 4'b1110;
															assign node13430 = (inp[2]) ? node13432 : 4'b1010;
																assign node13432 = (inp[4]) ? 4'b1111 : 4'b1110;
													assign node13435 = (inp[11]) ? node13451 : node13436;
														assign node13436 = (inp[4]) ? node13444 : node13437;
															assign node13437 = (inp[2]) ? node13441 : node13438;
																assign node13438 = (inp[1]) ? 4'b1010 : 4'b1110;
																assign node13441 = (inp[1]) ? 4'b1110 : 4'b1011;
															assign node13444 = (inp[2]) ? node13448 : node13445;
																assign node13445 = (inp[1]) ? 4'b1011 : 4'b1111;
																assign node13448 = (inp[1]) ? 4'b1110 : 4'b1010;
														assign node13451 = (inp[1]) ? node13455 : node13452;
															assign node13452 = (inp[2]) ? 4'b1011 : 4'b1111;
															assign node13455 = (inp[2]) ? node13457 : 4'b1011;
																assign node13457 = (inp[4]) ? 4'b1110 : 4'b1111;
												assign node13460 = (inp[9]) ? node13482 : node13461;
													assign node13461 = (inp[11]) ? node13467 : node13462;
														assign node13462 = (inp[1]) ? node13464 : 4'b1111;
															assign node13464 = (inp[2]) ? 4'b1110 : 4'b1010;
														assign node13467 = (inp[4]) ? node13475 : node13468;
															assign node13468 = (inp[2]) ? node13472 : node13469;
																assign node13469 = (inp[1]) ? 4'b1011 : 4'b1111;
																assign node13472 = (inp[1]) ? 4'b1111 : 4'b1011;
															assign node13475 = (inp[2]) ? node13479 : node13476;
																assign node13476 = (inp[1]) ? 4'b1011 : 4'b1111;
																assign node13479 = (inp[1]) ? 4'b1110 : 4'b1011;
													assign node13482 = (inp[11]) ? node13492 : node13483;
														assign node13483 = (inp[1]) ? 4'b1111 : node13484;
															assign node13484 = (inp[2]) ? node13488 : node13485;
																assign node13485 = (inp[4]) ? 4'b1110 : 4'b1111;
																assign node13488 = (inp[4]) ? 4'b1011 : 4'b1010;
														assign node13492 = (inp[1]) ? node13496 : node13493;
															assign node13493 = (inp[2]) ? 4'b1010 : 4'b1110;
															assign node13496 = (inp[2]) ? node13498 : 4'b1010;
																assign node13498 = (inp[4]) ? 4'b1111 : 4'b1110;
									assign node13501 = (inp[12]) ? node13679 : node13502;
										assign node13502 = (inp[4]) ? node13586 : node13503;
											assign node13503 = (inp[10]) ? node13541 : node13504;
												assign node13504 = (inp[9]) ? node13524 : node13505;
													assign node13505 = (inp[1]) ? node13515 : node13506;
														assign node13506 = (inp[15]) ? node13512 : node13507;
															assign node13507 = (inp[2]) ? 4'b1011 : node13508;
																assign node13508 = (inp[11]) ? 4'b1111 : 4'b1110;
															assign node13512 = (inp[2]) ? 4'b1110 : 4'b1010;
														assign node13515 = (inp[2]) ? node13519 : node13516;
															assign node13516 = (inp[15]) ? 4'b1011 : 4'b1111;
															assign node13519 = (inp[15]) ? 4'b1111 : node13520;
																assign node13520 = (inp[11]) ? 4'b1010 : 4'b1011;
													assign node13524 = (inp[1]) ? node13534 : node13525;
														assign node13525 = (inp[15]) ? node13531 : node13526;
															assign node13526 = (inp[2]) ? 4'b1010 : node13527;
																assign node13527 = (inp[11]) ? 4'b1110 : 4'b1111;
															assign node13531 = (inp[2]) ? 4'b1111 : 4'b1011;
														assign node13534 = (inp[15]) ? node13538 : node13535;
															assign node13535 = (inp[2]) ? 4'b1011 : 4'b1110;
															assign node13538 = (inp[2]) ? 4'b1110 : 4'b1010;
												assign node13541 = (inp[9]) ? node13567 : node13542;
													assign node13542 = (inp[1]) ? node13552 : node13543;
														assign node13543 = (inp[15]) ? node13549 : node13544;
															assign node13544 = (inp[2]) ? 4'b1010 : node13545;
																assign node13545 = (inp[11]) ? 4'b1110 : 4'b1111;
															assign node13549 = (inp[11]) ? 4'b1011 : 4'b1111;
														assign node13552 = (inp[11]) ? node13560 : node13553;
															assign node13553 = (inp[2]) ? node13557 : node13554;
																assign node13554 = (inp[15]) ? 4'b1010 : 4'b1110;
																assign node13557 = (inp[15]) ? 4'b1110 : 4'b1010;
															assign node13560 = (inp[15]) ? node13564 : node13561;
																assign node13561 = (inp[2]) ? 4'b1011 : 4'b1110;
																assign node13564 = (inp[2]) ? 4'b1110 : 4'b1010;
													assign node13567 = (inp[1]) ? node13577 : node13568;
														assign node13568 = (inp[15]) ? node13574 : node13569;
															assign node13569 = (inp[2]) ? 4'b1011 : node13570;
																assign node13570 = (inp[11]) ? 4'b1111 : 4'b1110;
															assign node13574 = (inp[2]) ? 4'b1110 : 4'b1010;
														assign node13577 = (inp[2]) ? node13581 : node13578;
															assign node13578 = (inp[15]) ? 4'b1011 : 4'b1111;
															assign node13581 = (inp[15]) ? 4'b1111 : node13582;
																assign node13582 = (inp[11]) ? 4'b1010 : 4'b1011;
											assign node13586 = (inp[15]) ? node13626 : node13587;
												assign node13587 = (inp[1]) ? node13603 : node13588;
													assign node13588 = (inp[2]) ? node13596 : node13589;
														assign node13589 = (inp[9]) ? node13593 : node13590;
															assign node13590 = (inp[10]) ? 4'b1000 : 4'b1001;
															assign node13593 = (inp[10]) ? 4'b1001 : 4'b1000;
														assign node13596 = (inp[9]) ? node13600 : node13597;
															assign node13597 = (inp[10]) ? 4'b1101 : 4'b1100;
															assign node13600 = (inp[10]) ? 4'b1100 : 4'b1101;
													assign node13603 = (inp[2]) ? node13611 : node13604;
														assign node13604 = (inp[9]) ? node13608 : node13605;
															assign node13605 = (inp[10]) ? 4'b1100 : 4'b1101;
															assign node13608 = (inp[10]) ? 4'b1101 : 4'b1100;
														assign node13611 = (inp[9]) ? node13619 : node13612;
															assign node13612 = (inp[10]) ? node13616 : node13613;
																assign node13613 = (inp[11]) ? 4'b1001 : 4'b1000;
																assign node13616 = (inp[11]) ? 4'b1000 : 4'b1001;
															assign node13619 = (inp[10]) ? node13623 : node13620;
																assign node13620 = (inp[11]) ? 4'b1000 : 4'b1001;
																assign node13623 = (inp[11]) ? 4'b1001 : 4'b1000;
												assign node13626 = (inp[2]) ? node13648 : node13627;
													assign node13627 = (inp[9]) ? node13635 : node13628;
														assign node13628 = (inp[1]) ? node13632 : node13629;
															assign node13629 = (inp[10]) ? 4'b1111 : 4'b1110;
															assign node13632 = (inp[10]) ? 4'b1110 : 4'b1111;
														assign node13635 = (inp[11]) ? node13643 : node13636;
															assign node13636 = (inp[1]) ? node13640 : node13637;
																assign node13637 = (inp[10]) ? 4'b1110 : 4'b1111;
																assign node13640 = (inp[10]) ? 4'b1111 : 4'b1110;
															assign node13643 = (inp[1]) ? 4'b1111 : node13644;
																assign node13644 = (inp[10]) ? 4'b1110 : 4'b1111;
													assign node13648 = (inp[11]) ? node13664 : node13649;
														assign node13649 = (inp[10]) ? node13657 : node13650;
															assign node13650 = (inp[1]) ? node13654 : node13651;
																assign node13651 = (inp[9]) ? 4'b1010 : 4'b1011;
																assign node13654 = (inp[9]) ? 4'b1011 : 4'b1010;
															assign node13657 = (inp[9]) ? node13661 : node13658;
																assign node13658 = (inp[1]) ? 4'b1011 : 4'b1010;
																assign node13661 = (inp[1]) ? 4'b1010 : 4'b1011;
														assign node13664 = (inp[1]) ? node13672 : node13665;
															assign node13665 = (inp[9]) ? node13669 : node13666;
																assign node13666 = (inp[10]) ? 4'b1011 : 4'b1010;
																assign node13669 = (inp[10]) ? 4'b1010 : 4'b1011;
															assign node13672 = (inp[9]) ? node13676 : node13673;
																assign node13673 = (inp[10]) ? 4'b1010 : 4'b1011;
																assign node13676 = (inp[10]) ? 4'b1011 : 4'b1010;
										assign node13679 = (inp[4]) ? node13789 : node13680;
											assign node13680 = (inp[15]) ? node13732 : node13681;
												assign node13681 = (inp[9]) ? node13707 : node13682;
													assign node13682 = (inp[10]) ? node13696 : node13683;
														assign node13683 = (inp[2]) ? node13691 : node13684;
															assign node13684 = (inp[1]) ? node13688 : node13685;
																assign node13685 = (inp[11]) ? 4'b1000 : 4'b1001;
																assign node13688 = (inp[11]) ? 4'b1101 : 4'b1100;
															assign node13691 = (inp[1]) ? 4'b1001 : node13692;
																assign node13692 = (inp[11]) ? 4'b1100 : 4'b1101;
														assign node13696 = (inp[2]) ? node13702 : node13697;
															assign node13697 = (inp[1]) ? node13699 : 4'b1001;
																assign node13699 = (inp[11]) ? 4'b1100 : 4'b1101;
															assign node13702 = (inp[1]) ? 4'b1000 : node13703;
																assign node13703 = (inp[11]) ? 4'b1101 : 4'b1100;
													assign node13707 = (inp[2]) ? node13721 : node13708;
														assign node13708 = (inp[1]) ? node13716 : node13709;
															assign node13709 = (inp[11]) ? node13713 : node13710;
																assign node13710 = (inp[10]) ? 4'b1001 : 4'b1000;
																assign node13713 = (inp[10]) ? 4'b1000 : 4'b1001;
															assign node13716 = (inp[10]) ? 4'b1100 : node13717;
																assign node13717 = (inp[11]) ? 4'b1100 : 4'b1101;
														assign node13721 = (inp[1]) ? node13729 : node13722;
															assign node13722 = (inp[11]) ? node13726 : node13723;
																assign node13723 = (inp[10]) ? 4'b1101 : 4'b1100;
																assign node13726 = (inp[10]) ? 4'b1100 : 4'b1101;
															assign node13729 = (inp[11]) ? 4'b1001 : 4'b1000;
												assign node13732 = (inp[11]) ? node13760 : node13733;
													assign node13733 = (inp[9]) ? node13747 : node13734;
														assign node13734 = (inp[10]) ? node13742 : node13735;
															assign node13735 = (inp[2]) ? node13739 : node13736;
																assign node13736 = (inp[1]) ? 4'b1000 : 4'b1100;
																assign node13739 = (inp[1]) ? 4'b1100 : 4'b1001;
															assign node13742 = (inp[1]) ? node13744 : 4'b1000;
																assign node13744 = (inp[2]) ? 4'b1101 : 4'b1001;
														assign node13747 = (inp[10]) ? node13753 : node13748;
															assign node13748 = (inp[2]) ? 4'b1000 : node13749;
																assign node13749 = (inp[1]) ? 4'b1001 : 4'b1101;
															assign node13753 = (inp[2]) ? node13757 : node13754;
																assign node13754 = (inp[1]) ? 4'b1000 : 4'b1100;
																assign node13757 = (inp[1]) ? 4'b1100 : 4'b1001;
													assign node13760 = (inp[10]) ? node13776 : node13761;
														assign node13761 = (inp[9]) ? node13769 : node13762;
															assign node13762 = (inp[2]) ? node13766 : node13763;
																assign node13763 = (inp[1]) ? 4'b1001 : 4'b1101;
																assign node13766 = (inp[1]) ? 4'b1101 : 4'b1001;
															assign node13769 = (inp[2]) ? node13773 : node13770;
																assign node13770 = (inp[1]) ? 4'b1000 : 4'b1100;
																assign node13773 = (inp[1]) ? 4'b1100 : 4'b1000;
														assign node13776 = (inp[9]) ? node13782 : node13777;
															assign node13777 = (inp[1]) ? node13779 : 4'b1000;
																assign node13779 = (inp[2]) ? 4'b1100 : 4'b1000;
															assign node13782 = (inp[1]) ? node13786 : node13783;
																assign node13783 = (inp[2]) ? 4'b1001 : 4'b1101;
																assign node13786 = (inp[2]) ? 4'b1101 : 4'b1001;
											assign node13789 = (inp[15]) ? node13835 : node13790;
												assign node13790 = (inp[9]) ? node13810 : node13791;
													assign node13791 = (inp[10]) ? node13801 : node13792;
														assign node13792 = (inp[1]) ? node13798 : node13793;
															assign node13793 = (inp[2]) ? 4'b1011 : node13794;
																assign node13794 = (inp[11]) ? 4'b1110 : 4'b1111;
															assign node13798 = (inp[2]) ? 4'b1110 : 4'b1011;
														assign node13801 = (inp[1]) ? node13807 : node13802;
															assign node13802 = (inp[2]) ? 4'b1010 : node13803;
																assign node13803 = (inp[11]) ? 4'b1111 : 4'b1110;
															assign node13807 = (inp[2]) ? 4'b1111 : 4'b1010;
													assign node13810 = (inp[10]) ? node13826 : node13811;
														assign node13811 = (inp[11]) ? node13819 : node13812;
															assign node13812 = (inp[2]) ? node13816 : node13813;
																assign node13813 = (inp[1]) ? 4'b1010 : 4'b1110;
																assign node13816 = (inp[1]) ? 4'b1111 : 4'b1010;
															assign node13819 = (inp[1]) ? node13823 : node13820;
																assign node13820 = (inp[2]) ? 4'b1010 : 4'b1111;
																assign node13823 = (inp[2]) ? 4'b1111 : 4'b1010;
														assign node13826 = (inp[2]) ? node13832 : node13827;
															assign node13827 = (inp[1]) ? 4'b1011 : node13828;
																assign node13828 = (inp[11]) ? 4'b1110 : 4'b1111;
															assign node13832 = (inp[1]) ? 4'b1110 : 4'b1011;
												assign node13835 = (inp[11]) ? node13865 : node13836;
													assign node13836 = (inp[9]) ? node13852 : node13837;
														assign node13837 = (inp[2]) ? node13845 : node13838;
															assign node13838 = (inp[10]) ? node13842 : node13839;
																assign node13839 = (inp[1]) ? 4'b1001 : 4'b1101;
																assign node13842 = (inp[1]) ? 4'b1000 : 4'b1100;
															assign node13845 = (inp[1]) ? node13849 : node13846;
																assign node13846 = (inp[10]) ? 4'b1001 : 4'b1000;
																assign node13849 = (inp[10]) ? 4'b1101 : 4'b1100;
														assign node13852 = (inp[1]) ? node13858 : node13853;
															assign node13853 = (inp[2]) ? 4'b1001 : node13854;
																assign node13854 = (inp[10]) ? 4'b1101 : 4'b1100;
															assign node13858 = (inp[2]) ? node13862 : node13859;
																assign node13859 = (inp[10]) ? 4'b1001 : 4'b1000;
																assign node13862 = (inp[10]) ? 4'b1100 : 4'b1101;
													assign node13865 = (inp[9]) ? node13879 : node13866;
														assign node13866 = (inp[10]) ? node13872 : node13867;
															assign node13867 = (inp[1]) ? 4'b1100 : node13868;
																assign node13868 = (inp[2]) ? 4'b1001 : 4'b1101;
															assign node13872 = (inp[2]) ? node13876 : node13873;
																assign node13873 = (inp[1]) ? 4'b1000 : 4'b1100;
																assign node13876 = (inp[1]) ? 4'b1101 : 4'b1000;
														assign node13879 = (inp[10]) ? node13887 : node13880;
															assign node13880 = (inp[1]) ? node13884 : node13881;
																assign node13881 = (inp[2]) ? 4'b1000 : 4'b1100;
																assign node13884 = (inp[2]) ? 4'b1101 : 4'b1000;
															assign node13887 = (inp[2]) ? 4'b1100 : 4'b1101;
								assign node13890 = (inp[15]) ? node14328 : node13891;
									assign node13891 = (inp[11]) ? node14095 : node13892;
										assign node13892 = (inp[2]) ? node13996 : node13893;
											assign node13893 = (inp[12]) ? node13951 : node13894;
												assign node13894 = (inp[1]) ? node13924 : node13895;
													assign node13895 = (inp[7]) ? node13911 : node13896;
														assign node13896 = (inp[4]) ? node13904 : node13897;
															assign node13897 = (inp[9]) ? node13901 : node13898;
																assign node13898 = (inp[10]) ? 4'b1101 : 4'b1100;
																assign node13901 = (inp[10]) ? 4'b1100 : 4'b1101;
															assign node13904 = (inp[9]) ? node13908 : node13905;
																assign node13905 = (inp[10]) ? 4'b1111 : 4'b1110;
																assign node13908 = (inp[10]) ? 4'b1110 : 4'b1111;
														assign node13911 = (inp[4]) ? node13919 : node13912;
															assign node13912 = (inp[10]) ? node13916 : node13913;
																assign node13913 = (inp[9]) ? 4'b1111 : 4'b1110;
																assign node13916 = (inp[9]) ? 4'b1110 : 4'b1111;
															assign node13919 = (inp[9]) ? 4'b1001 : node13920;
																assign node13920 = (inp[10]) ? 4'b1001 : 4'b1000;
													assign node13924 = (inp[7]) ? node13940 : node13925;
														assign node13925 = (inp[4]) ? node13933 : node13926;
															assign node13926 = (inp[9]) ? node13930 : node13927;
																assign node13927 = (inp[10]) ? 4'b1001 : 4'b1000;
																assign node13930 = (inp[10]) ? 4'b1000 : 4'b1001;
															assign node13933 = (inp[10]) ? node13937 : node13934;
																assign node13934 = (inp[9]) ? 4'b1011 : 4'b1010;
																assign node13937 = (inp[9]) ? 4'b1010 : 4'b1011;
														assign node13940 = (inp[4]) ? node13946 : node13941;
															assign node13941 = (inp[10]) ? node13943 : 4'b1110;
																assign node13943 = (inp[9]) ? 4'b1110 : 4'b1111;
															assign node13946 = (inp[9]) ? 4'b1101 : node13947;
																assign node13947 = (inp[10]) ? 4'b1101 : 4'b1100;
												assign node13951 = (inp[7]) ? node13967 : node13952;
													assign node13952 = (inp[4]) ? node13960 : node13953;
														assign node13953 = (inp[1]) ? node13955 : 4'b1111;
															assign node13955 = (inp[9]) ? node13957 : 4'b1011;
																assign node13957 = (inp[10]) ? 4'b1011 : 4'b1010;
														assign node13960 = (inp[10]) ? node13964 : node13961;
															assign node13961 = (inp[9]) ? 4'b1001 : 4'b1000;
															assign node13964 = (inp[9]) ? 4'b1000 : 4'b1001;
													assign node13967 = (inp[4]) ? node13983 : node13968;
														assign node13968 = (inp[1]) ? node13976 : node13969;
															assign node13969 = (inp[9]) ? node13973 : node13970;
																assign node13970 = (inp[10]) ? 4'b1000 : 4'b1001;
																assign node13973 = (inp[10]) ? 4'b1001 : 4'b1000;
															assign node13976 = (inp[9]) ? node13980 : node13977;
																assign node13977 = (inp[10]) ? 4'b1101 : 4'b1100;
																assign node13980 = (inp[10]) ? 4'b1100 : 4'b1101;
														assign node13983 = (inp[1]) ? node13989 : node13984;
															assign node13984 = (inp[9]) ? 4'b1111 : node13985;
																assign node13985 = (inp[10]) ? 4'b1110 : 4'b1111;
															assign node13989 = (inp[10]) ? node13993 : node13990;
																assign node13990 = (inp[9]) ? 4'b1011 : 4'b1010;
																assign node13993 = (inp[9]) ? 4'b1010 : 4'b1011;
											assign node13996 = (inp[7]) ? node14050 : node13997;
												assign node13997 = (inp[1]) ? node14021 : node13998;
													assign node13998 = (inp[4]) ? node14012 : node13999;
														assign node13999 = (inp[12]) ? node14007 : node14000;
															assign node14000 = (inp[9]) ? node14004 : node14001;
																assign node14001 = (inp[10]) ? 4'b1001 : 4'b1000;
																assign node14004 = (inp[10]) ? 4'b1000 : 4'b1001;
															assign node14007 = (inp[10]) ? 4'b1010 : node14008;
																assign node14008 = (inp[9]) ? 4'b1011 : 4'b1010;
														assign node14012 = (inp[12]) ? node14016 : node14013;
															assign node14013 = (inp[10]) ? 4'b1010 : 4'b1011;
															assign node14016 = (inp[9]) ? node14018 : 4'b1100;
																assign node14018 = (inp[10]) ? 4'b1101 : 4'b1100;
													assign node14021 = (inp[4]) ? node14037 : node14022;
														assign node14022 = (inp[12]) ? node14030 : node14023;
															assign node14023 = (inp[10]) ? node14027 : node14024;
																assign node14024 = (inp[9]) ? 4'b1101 : 4'b1100;
																assign node14027 = (inp[9]) ? 4'b1100 : 4'b1101;
															assign node14030 = (inp[9]) ? node14034 : node14031;
																assign node14031 = (inp[10]) ? 4'b1110 : 4'b1111;
																assign node14034 = (inp[10]) ? 4'b1111 : 4'b1110;
														assign node14037 = (inp[12]) ? node14043 : node14038;
															assign node14038 = (inp[9]) ? 4'b1110 : node14039;
																assign node14039 = (inp[10]) ? 4'b1110 : 4'b1111;
															assign node14043 = (inp[9]) ? node14047 : node14044;
																assign node14044 = (inp[10]) ? 4'b1100 : 4'b1101;
																assign node14047 = (inp[10]) ? 4'b1101 : 4'b1100;
												assign node14050 = (inp[1]) ? node14074 : node14051;
													assign node14051 = (inp[10]) ? node14065 : node14052;
														assign node14052 = (inp[4]) ? node14058 : node14053;
															assign node14053 = (inp[12]) ? 4'b1100 : node14054;
																assign node14054 = (inp[9]) ? 4'b1011 : 4'b1010;
															assign node14058 = (inp[12]) ? node14062 : node14059;
																assign node14059 = (inp[9]) ? 4'b1100 : 4'b1101;
																assign node14062 = (inp[9]) ? 4'b1011 : 4'b1010;
														assign node14065 = (inp[9]) ? node14067 : 4'b1100;
															assign node14067 = (inp[12]) ? node14071 : node14068;
																assign node14068 = (inp[4]) ? 4'b1101 : 4'b1010;
																assign node14071 = (inp[4]) ? 4'b1010 : 4'b1101;
													assign node14074 = (inp[4]) ? node14086 : node14075;
														assign node14075 = (inp[12]) ? node14079 : node14076;
															assign node14076 = (inp[10]) ? 4'b1010 : 4'b1011;
															assign node14079 = (inp[10]) ? node14083 : node14080;
																assign node14080 = (inp[9]) ? 4'b1001 : 4'b1000;
																assign node14083 = (inp[9]) ? 4'b1000 : 4'b1001;
														assign node14086 = (inp[12]) ? 4'b1111 : node14087;
															assign node14087 = (inp[9]) ? node14091 : node14088;
																assign node14088 = (inp[10]) ? 4'b1001 : 4'b1000;
																assign node14091 = (inp[10]) ? 4'b1000 : 4'b1001;
										assign node14095 = (inp[1]) ? node14211 : node14096;
											assign node14096 = (inp[2]) ? node14158 : node14097;
												assign node14097 = (inp[12]) ? node14129 : node14098;
													assign node14098 = (inp[4]) ? node14114 : node14099;
														assign node14099 = (inp[7]) ? node14107 : node14100;
															assign node14100 = (inp[10]) ? node14104 : node14101;
																assign node14101 = (inp[9]) ? 4'b1101 : 4'b1100;
																assign node14104 = (inp[9]) ? 4'b1100 : 4'b1101;
															assign node14107 = (inp[9]) ? node14111 : node14108;
																assign node14108 = (inp[10]) ? 4'b1111 : 4'b1110;
																assign node14111 = (inp[10]) ? 4'b1110 : 4'b1111;
														assign node14114 = (inp[7]) ? node14122 : node14115;
															assign node14115 = (inp[10]) ? node14119 : node14116;
																assign node14116 = (inp[9]) ? 4'b1111 : 4'b1110;
																assign node14119 = (inp[9]) ? 4'b1110 : 4'b1111;
															assign node14122 = (inp[10]) ? node14126 : node14123;
																assign node14123 = (inp[9]) ? 4'b1000 : 4'b1001;
																assign node14126 = (inp[9]) ? 4'b1001 : 4'b1000;
													assign node14129 = (inp[7]) ? node14143 : node14130;
														assign node14130 = (inp[4]) ? node14136 : node14131;
															assign node14131 = (inp[9]) ? node14133 : 4'b1111;
																assign node14133 = (inp[10]) ? 4'b1110 : 4'b1111;
															assign node14136 = (inp[9]) ? node14140 : node14137;
																assign node14137 = (inp[10]) ? 4'b1000 : 4'b1001;
																assign node14140 = (inp[10]) ? 4'b1001 : 4'b1000;
														assign node14143 = (inp[4]) ? node14151 : node14144;
															assign node14144 = (inp[9]) ? node14148 : node14145;
																assign node14145 = (inp[10]) ? 4'b1000 : 4'b1001;
																assign node14148 = (inp[10]) ? 4'b1001 : 4'b1000;
															assign node14151 = (inp[10]) ? node14155 : node14152;
																assign node14152 = (inp[9]) ? 4'b1110 : 4'b1111;
																assign node14155 = (inp[9]) ? 4'b1111 : 4'b1110;
												assign node14158 = (inp[7]) ? node14184 : node14159;
													assign node14159 = (inp[4]) ? node14175 : node14160;
														assign node14160 = (inp[12]) ? node14168 : node14161;
															assign node14161 = (inp[9]) ? node14165 : node14162;
																assign node14162 = (inp[10]) ? 4'b1000 : 4'b1001;
																assign node14165 = (inp[10]) ? 4'b1001 : 4'b1000;
															assign node14168 = (inp[9]) ? node14172 : node14169;
																assign node14169 = (inp[10]) ? 4'b1010 : 4'b1011;
																assign node14172 = (inp[10]) ? 4'b1011 : 4'b1010;
														assign node14175 = (inp[12]) ? 4'b1101 : node14176;
															assign node14176 = (inp[9]) ? node14180 : node14177;
																assign node14177 = (inp[10]) ? 4'b1011 : 4'b1010;
																assign node14180 = (inp[10]) ? 4'b1010 : 4'b1011;
													assign node14184 = (inp[4]) ? node14198 : node14185;
														assign node14185 = (inp[12]) ? node14193 : node14186;
															assign node14186 = (inp[10]) ? node14190 : node14187;
																assign node14187 = (inp[9]) ? 4'b1010 : 4'b1011;
																assign node14190 = (inp[9]) ? 4'b1011 : 4'b1010;
															assign node14193 = (inp[10]) ? 4'b1101 : node14194;
																assign node14194 = (inp[9]) ? 4'b1100 : 4'b1101;
														assign node14198 = (inp[12]) ? node14206 : node14199;
															assign node14199 = (inp[9]) ? node14203 : node14200;
																assign node14200 = (inp[10]) ? 4'b1101 : 4'b1100;
																assign node14203 = (inp[10]) ? 4'b1100 : 4'b1101;
															assign node14206 = (inp[10]) ? 4'b1011 : node14207;
																assign node14207 = (inp[9]) ? 4'b1010 : 4'b1011;
											assign node14211 = (inp[2]) ? node14265 : node14212;
												assign node14212 = (inp[7]) ? node14236 : node14213;
													assign node14213 = (inp[12]) ? node14223 : node14214;
														assign node14214 = (inp[4]) ? node14216 : 4'b1001;
															assign node14216 = (inp[10]) ? node14220 : node14217;
																assign node14217 = (inp[9]) ? 4'b1010 : 4'b1011;
																assign node14220 = (inp[9]) ? 4'b1011 : 4'b1010;
														assign node14223 = (inp[4]) ? node14229 : node14224;
															assign node14224 = (inp[9]) ? node14226 : 4'b1010;
																assign node14226 = (inp[10]) ? 4'b1010 : 4'b1011;
															assign node14229 = (inp[10]) ? node14233 : node14230;
																assign node14230 = (inp[9]) ? 4'b1001 : 4'b1000;
																assign node14233 = (inp[9]) ? 4'b1000 : 4'b1001;
													assign node14236 = (inp[4]) ? node14252 : node14237;
														assign node14237 = (inp[12]) ? node14245 : node14238;
															assign node14238 = (inp[9]) ? node14242 : node14239;
																assign node14239 = (inp[10]) ? 4'b1110 : 4'b1111;
																assign node14242 = (inp[10]) ? 4'b1111 : 4'b1110;
															assign node14245 = (inp[9]) ? node14249 : node14246;
																assign node14246 = (inp[10]) ? 4'b1101 : 4'b1100;
																assign node14249 = (inp[10]) ? 4'b1100 : 4'b1101;
														assign node14252 = (inp[12]) ? node14260 : node14253;
															assign node14253 = (inp[10]) ? node14257 : node14254;
																assign node14254 = (inp[9]) ? 4'b1100 : 4'b1101;
																assign node14257 = (inp[9]) ? 4'b1101 : 4'b1100;
															assign node14260 = (inp[10]) ? 4'b1011 : node14261;
																assign node14261 = (inp[9]) ? 4'b1010 : 4'b1011;
												assign node14265 = (inp[7]) ? node14297 : node14266;
													assign node14266 = (inp[10]) ? node14282 : node14267;
														assign node14267 = (inp[12]) ? node14275 : node14268;
															assign node14268 = (inp[4]) ? node14272 : node14269;
																assign node14269 = (inp[9]) ? 4'b1100 : 4'b1101;
																assign node14272 = (inp[9]) ? 4'b1111 : 4'b1110;
															assign node14275 = (inp[4]) ? node14279 : node14276;
																assign node14276 = (inp[9]) ? 4'b1111 : 4'b1110;
																assign node14279 = (inp[9]) ? 4'b1100 : 4'b1101;
														assign node14282 = (inp[12]) ? node14290 : node14283;
															assign node14283 = (inp[4]) ? node14287 : node14284;
																assign node14284 = (inp[9]) ? 4'b1101 : 4'b1100;
																assign node14287 = (inp[9]) ? 4'b1110 : 4'b1111;
															assign node14290 = (inp[4]) ? node14294 : node14291;
																assign node14291 = (inp[9]) ? 4'b1110 : 4'b1111;
																assign node14294 = (inp[9]) ? 4'b1101 : 4'b1100;
													assign node14297 = (inp[4]) ? node14313 : node14298;
														assign node14298 = (inp[12]) ? node14306 : node14299;
															assign node14299 = (inp[10]) ? node14303 : node14300;
																assign node14300 = (inp[9]) ? 4'b1010 : 4'b1011;
																assign node14303 = (inp[9]) ? 4'b1011 : 4'b1010;
															assign node14306 = (inp[10]) ? node14310 : node14307;
																assign node14307 = (inp[9]) ? 4'b1000 : 4'b1001;
																assign node14310 = (inp[9]) ? 4'b1001 : 4'b1000;
														assign node14313 = (inp[12]) ? node14321 : node14314;
															assign node14314 = (inp[9]) ? node14318 : node14315;
																assign node14315 = (inp[10]) ? 4'b1001 : 4'b1000;
																assign node14318 = (inp[10]) ? 4'b1000 : 4'b1001;
															assign node14321 = (inp[10]) ? node14325 : node14322;
																assign node14322 = (inp[9]) ? 4'b1111 : 4'b1110;
																assign node14325 = (inp[9]) ? 4'b1110 : 4'b1111;
									assign node14328 = (inp[12]) ? node14504 : node14329;
										assign node14329 = (inp[7]) ? node14417 : node14330;
											assign node14330 = (inp[10]) ? node14368 : node14331;
												assign node14331 = (inp[4]) ? node14351 : node14332;
													assign node14332 = (inp[1]) ? node14344 : node14333;
														assign node14333 = (inp[2]) ? node14337 : node14334;
															assign node14334 = (inp[9]) ? 4'b1100 : 4'b1101;
															assign node14337 = (inp[11]) ? node14341 : node14338;
																assign node14338 = (inp[9]) ? 4'b1000 : 4'b1001;
																assign node14341 = (inp[9]) ? 4'b1001 : 4'b1000;
														assign node14344 = (inp[2]) ? node14348 : node14345;
															assign node14345 = (inp[9]) ? 4'b1001 : 4'b1000;
															assign node14348 = (inp[9]) ? 4'b1101 : 4'b1100;
													assign node14351 = (inp[1]) ? node14359 : node14352;
														assign node14352 = (inp[2]) ? node14354 : 4'b1000;
															assign node14354 = (inp[9]) ? 4'b1100 : node14355;
																assign node14355 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node14359 = (inp[2]) ? node14363 : node14360;
															assign node14360 = (inp[9]) ? 4'b1101 : 4'b1100;
															assign node14363 = (inp[11]) ? 4'b1000 : node14364;
																assign node14364 = (inp[9]) ? 4'b1000 : 4'b1001;
												assign node14368 = (inp[9]) ? node14398 : node14369;
													assign node14369 = (inp[1]) ? node14383 : node14370;
														assign node14370 = (inp[4]) ? node14376 : node14371;
															assign node14371 = (inp[2]) ? node14373 : 4'b1100;
																assign node14373 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node14376 = (inp[2]) ? node14380 : node14377;
																assign node14377 = (inp[11]) ? 4'b1001 : 4'b1000;
																assign node14380 = (inp[11]) ? 4'b1100 : 4'b1101;
														assign node14383 = (inp[11]) ? node14391 : node14384;
															assign node14384 = (inp[4]) ? node14388 : node14385;
																assign node14385 = (inp[2]) ? 4'b1101 : 4'b1001;
																assign node14388 = (inp[2]) ? 4'b1000 : 4'b1101;
															assign node14391 = (inp[2]) ? node14395 : node14392;
																assign node14392 = (inp[4]) ? 4'b1101 : 4'b1001;
																assign node14395 = (inp[4]) ? 4'b1001 : 4'b1101;
													assign node14398 = (inp[1]) ? node14408 : node14399;
														assign node14399 = (inp[11]) ? node14401 : 4'b1001;
															assign node14401 = (inp[4]) ? node14405 : node14402;
																assign node14402 = (inp[2]) ? 4'b1000 : 4'b1101;
																assign node14405 = (inp[2]) ? 4'b1101 : 4'b1000;
														assign node14408 = (inp[2]) ? node14412 : node14409;
															assign node14409 = (inp[4]) ? 4'b1100 : 4'b1000;
															assign node14412 = (inp[4]) ? node14414 : 4'b1100;
																assign node14414 = (inp[11]) ? 4'b1000 : 4'b1001;
											assign node14417 = (inp[10]) ? node14449 : node14418;
												assign node14418 = (inp[4]) ? node14438 : node14419;
													assign node14419 = (inp[2]) ? node14429 : node14420;
														assign node14420 = (inp[9]) ? 4'b1010 : node14421;
															assign node14421 = (inp[11]) ? node14425 : node14422;
																assign node14422 = (inp[1]) ? 4'b1010 : 4'b1011;
																assign node14425 = (inp[1]) ? 4'b1011 : 4'b1010;
														assign node14429 = (inp[11]) ? node14431 : 4'b1110;
															assign node14431 = (inp[1]) ? node14435 : node14432;
																assign node14432 = (inp[9]) ? 4'b1111 : 4'b1110;
																assign node14435 = (inp[9]) ? 4'b1110 : 4'b1111;
													assign node14438 = (inp[2]) ? node14442 : node14439;
														assign node14439 = (inp[9]) ? 4'b1111 : 4'b1110;
														assign node14442 = (inp[9]) ? node14446 : node14443;
															assign node14443 = (inp[1]) ? 4'b1010 : 4'b1011;
															assign node14446 = (inp[1]) ? 4'b1011 : 4'b1010;
												assign node14449 = (inp[11]) ? node14475 : node14450;
													assign node14450 = (inp[9]) ? node14460 : node14451;
														assign node14451 = (inp[1]) ? node14453 : 4'b1010;
															assign node14453 = (inp[4]) ? node14457 : node14454;
																assign node14454 = (inp[2]) ? 4'b1111 : 4'b1011;
																assign node14457 = (inp[2]) ? 4'b1011 : 4'b1111;
														assign node14460 = (inp[1]) ? node14468 : node14461;
															assign node14461 = (inp[2]) ? node14465 : node14462;
																assign node14462 = (inp[4]) ? 4'b1111 : 4'b1011;
																assign node14465 = (inp[4]) ? 4'b1011 : 4'b1111;
															assign node14468 = (inp[2]) ? node14472 : node14469;
																assign node14469 = (inp[4]) ? 4'b1110 : 4'b1010;
																assign node14472 = (inp[4]) ? 4'b1010 : 4'b1110;
													assign node14475 = (inp[2]) ? node14491 : node14476;
														assign node14476 = (inp[4]) ? node14484 : node14477;
															assign node14477 = (inp[9]) ? node14481 : node14478;
																assign node14478 = (inp[1]) ? 4'b1010 : 4'b1011;
																assign node14481 = (inp[1]) ? 4'b1011 : 4'b1010;
															assign node14484 = (inp[1]) ? node14488 : node14485;
																assign node14485 = (inp[9]) ? 4'b1110 : 4'b1111;
																assign node14488 = (inp[9]) ? 4'b1111 : 4'b1110;
														assign node14491 = (inp[4]) ? node14499 : node14492;
															assign node14492 = (inp[1]) ? node14496 : node14493;
																assign node14493 = (inp[9]) ? 4'b1110 : 4'b1111;
																assign node14496 = (inp[9]) ? 4'b1111 : 4'b1110;
															assign node14499 = (inp[1]) ? node14501 : 4'b1010;
																assign node14501 = (inp[9]) ? 4'b1010 : 4'b1011;
										assign node14504 = (inp[7]) ? node14610 : node14505;
											assign node14505 = (inp[11]) ? node14561 : node14506;
												assign node14506 = (inp[2]) ? node14530 : node14507;
													assign node14507 = (inp[1]) ? node14523 : node14508;
														assign node14508 = (inp[4]) ? node14516 : node14509;
															assign node14509 = (inp[10]) ? node14513 : node14510;
																assign node14510 = (inp[9]) ? 4'b1110 : 4'b1111;
																assign node14513 = (inp[9]) ? 4'b1111 : 4'b1110;
															assign node14516 = (inp[10]) ? node14520 : node14517;
																assign node14517 = (inp[9]) ? 4'b1110 : 4'b1111;
																assign node14520 = (inp[9]) ? 4'b1111 : 4'b1110;
														assign node14523 = (inp[9]) ? node14527 : node14524;
															assign node14524 = (inp[10]) ? 4'b1010 : 4'b1011;
															assign node14527 = (inp[10]) ? 4'b1011 : 4'b1010;
													assign node14530 = (inp[1]) ? node14546 : node14531;
														assign node14531 = (inp[4]) ? node14539 : node14532;
															assign node14532 = (inp[9]) ? node14536 : node14533;
																assign node14533 = (inp[10]) ? 4'b1010 : 4'b1011;
																assign node14536 = (inp[10]) ? 4'b1011 : 4'b1010;
															assign node14539 = (inp[10]) ? node14543 : node14540;
																assign node14540 = (inp[9]) ? 4'b1010 : 4'b1011;
																assign node14543 = (inp[9]) ? 4'b1011 : 4'b1010;
														assign node14546 = (inp[10]) ? node14554 : node14547;
															assign node14547 = (inp[9]) ? node14551 : node14548;
																assign node14548 = (inp[4]) ? 4'b1110 : 4'b1111;
																assign node14551 = (inp[4]) ? 4'b1111 : 4'b1110;
															assign node14554 = (inp[4]) ? node14558 : node14555;
																assign node14555 = (inp[9]) ? 4'b1111 : 4'b1110;
																assign node14558 = (inp[9]) ? 4'b1110 : 4'b1111;
												assign node14561 = (inp[9]) ? node14587 : node14562;
													assign node14562 = (inp[10]) ? node14574 : node14563;
														assign node14563 = (inp[2]) ? node14569 : node14564;
															assign node14564 = (inp[1]) ? 4'b1010 : node14565;
																assign node14565 = (inp[4]) ? 4'b1110 : 4'b1111;
															assign node14569 = (inp[1]) ? 4'b1111 : node14570;
																assign node14570 = (inp[4]) ? 4'b1011 : 4'b1010;
														assign node14574 = (inp[2]) ? node14582 : node14575;
															assign node14575 = (inp[4]) ? node14579 : node14576;
																assign node14576 = (inp[1]) ? 4'b1010 : 4'b1110;
																assign node14579 = (inp[1]) ? 4'b1011 : 4'b1111;
															assign node14582 = (inp[1]) ? 4'b1110 : node14583;
																assign node14583 = (inp[4]) ? 4'b1010 : 4'b1011;
													assign node14587 = (inp[4]) ? node14599 : node14588;
														assign node14588 = (inp[10]) ? node14596 : node14589;
															assign node14589 = (inp[2]) ? node14593 : node14590;
																assign node14590 = (inp[1]) ? 4'b1010 : 4'b1110;
																assign node14593 = (inp[1]) ? 4'b1110 : 4'b1011;
															assign node14596 = (inp[2]) ? 4'b1010 : 4'b1011;
														assign node14599 = (inp[1]) ? node14605 : node14600;
															assign node14600 = (inp[2]) ? 4'b1010 : node14601;
																assign node14601 = (inp[10]) ? 4'b1110 : 4'b1111;
															assign node14605 = (inp[2]) ? 4'b1111 : node14606;
																assign node14606 = (inp[10]) ? 4'b1010 : 4'b1011;
											assign node14610 = (inp[4]) ? node14652 : node14611;
												assign node14611 = (inp[2]) ? node14627 : node14612;
													assign node14612 = (inp[1]) ? node14620 : node14613;
														assign node14613 = (inp[10]) ? node14617 : node14614;
															assign node14614 = (inp[9]) ? 4'b1101 : 4'b1100;
															assign node14617 = (inp[9]) ? 4'b1100 : 4'b1101;
														assign node14620 = (inp[10]) ? node14624 : node14621;
															assign node14621 = (inp[9]) ? 4'b1001 : 4'b1000;
															assign node14624 = (inp[9]) ? 4'b1000 : 4'b1001;
													assign node14627 = (inp[1]) ? node14639 : node14628;
														assign node14628 = (inp[10]) ? node14634 : node14629;
															assign node14629 = (inp[9]) ? 4'b1000 : node14630;
																assign node14630 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node14634 = (inp[9]) ? 4'b1001 : node14635;
																assign node14635 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node14639 = (inp[11]) ? node14647 : node14640;
															assign node14640 = (inp[10]) ? node14644 : node14641;
																assign node14641 = (inp[9]) ? 4'b1101 : 4'b1100;
																assign node14644 = (inp[9]) ? 4'b1100 : 4'b1101;
															assign node14647 = (inp[10]) ? 4'b1100 : node14648;
																assign node14648 = (inp[9]) ? 4'b1101 : 4'b1100;
												assign node14652 = (inp[10]) ? node14678 : node14653;
													assign node14653 = (inp[2]) ? node14667 : node14654;
														assign node14654 = (inp[1]) ? node14660 : node14655;
															assign node14655 = (inp[11]) ? node14657 : 4'b1101;
																assign node14657 = (inp[9]) ? 4'b1100 : 4'b1101;
															assign node14660 = (inp[11]) ? node14664 : node14661;
																assign node14661 = (inp[9]) ? 4'b1001 : 4'b1000;
																assign node14664 = (inp[9]) ? 4'b1000 : 4'b1001;
														assign node14667 = (inp[1]) ? node14671 : node14668;
															assign node14668 = (inp[9]) ? 4'b1001 : 4'b1000;
															assign node14671 = (inp[11]) ? node14675 : node14672;
																assign node14672 = (inp[9]) ? 4'b1100 : 4'b1101;
																assign node14675 = (inp[9]) ? 4'b1101 : 4'b1100;
													assign node14678 = (inp[11]) ? node14686 : node14679;
														assign node14679 = (inp[9]) ? node14681 : 4'b1001;
															assign node14681 = (inp[1]) ? node14683 : 4'b1000;
																assign node14683 = (inp[2]) ? 4'b1101 : 4'b1000;
														assign node14686 = (inp[2]) ? node14692 : node14687;
															assign node14687 = (inp[1]) ? 4'b1001 : node14688;
																assign node14688 = (inp[9]) ? 4'b1101 : 4'b1100;
															assign node14692 = (inp[1]) ? 4'b1101 : 4'b1001;
							assign node14695 = (inp[12]) ? node15191 : node14696;
								assign node14696 = (inp[15]) ? node14940 : node14697;
									assign node14697 = (inp[7]) ? node14839 : node14698;
										assign node14698 = (inp[1]) ? node14776 : node14699;
											assign node14699 = (inp[0]) ? node14739 : node14700;
												assign node14700 = (inp[10]) ? node14720 : node14701;
													assign node14701 = (inp[9]) ? node14713 : node14702;
														assign node14702 = (inp[11]) ? node14708 : node14703;
															assign node14703 = (inp[2]) ? node14705 : 4'b1100;
																assign node14705 = (inp[4]) ? 4'b1100 : 4'b1101;
															assign node14708 = (inp[4]) ? 4'b1101 : node14709;
																assign node14709 = (inp[2]) ? 4'b1100 : 4'b1101;
														assign node14713 = (inp[11]) ? node14715 : 4'b1101;
															assign node14715 = (inp[2]) ? node14717 : 4'b1100;
																assign node14717 = (inp[4]) ? 4'b1100 : 4'b1101;
													assign node14720 = (inp[9]) ? node14728 : node14721;
														assign node14721 = (inp[11]) ? 4'b1101 : node14722;
															assign node14722 = (inp[4]) ? 4'b1100 : node14723;
																assign node14723 = (inp[2]) ? 4'b1101 : 4'b1100;
														assign node14728 = (inp[11]) ? node14734 : node14729;
															assign node14729 = (inp[4]) ? 4'b1101 : node14730;
																assign node14730 = (inp[2]) ? 4'b1100 : 4'b1101;
															assign node14734 = (inp[4]) ? 4'b1100 : node14735;
																assign node14735 = (inp[2]) ? 4'b1101 : 4'b1100;
												assign node14739 = (inp[10]) ? node14763 : node14740;
													assign node14740 = (inp[9]) ? node14752 : node14741;
														assign node14741 = (inp[11]) ? node14747 : node14742;
															assign node14742 = (inp[4]) ? node14744 : 4'b1100;
																assign node14744 = (inp[2]) ? 4'b1101 : 4'b1100;
															assign node14747 = (inp[2]) ? node14749 : 4'b1101;
																assign node14749 = (inp[4]) ? 4'b1100 : 4'b1101;
														assign node14752 = (inp[11]) ? node14758 : node14753;
															assign node14753 = (inp[4]) ? node14755 : 4'b1101;
																assign node14755 = (inp[2]) ? 4'b1100 : 4'b1101;
															assign node14758 = (inp[2]) ? node14760 : 4'b1100;
																assign node14760 = (inp[4]) ? 4'b1101 : 4'b1100;
													assign node14763 = (inp[11]) ? node14769 : node14764;
														assign node14764 = (inp[9]) ? node14766 : 4'b1100;
															assign node14766 = (inp[4]) ? 4'b1100 : 4'b1101;
														assign node14769 = (inp[9]) ? node14771 : 4'b1101;
															assign node14771 = (inp[4]) ? node14773 : 4'b1100;
																assign node14773 = (inp[2]) ? 4'b1101 : 4'b1100;
											assign node14776 = (inp[4]) ? node14800 : node14777;
												assign node14777 = (inp[9]) ? node14789 : node14778;
													assign node14778 = (inp[11]) ? node14784 : node14779;
														assign node14779 = (inp[2]) ? 4'b1001 : node14780;
															assign node14780 = (inp[0]) ? 4'b1000 : 4'b1001;
														assign node14784 = (inp[2]) ? 4'b1000 : node14785;
															assign node14785 = (inp[0]) ? 4'b1001 : 4'b1000;
													assign node14789 = (inp[11]) ? node14795 : node14790;
														assign node14790 = (inp[2]) ? 4'b1000 : node14791;
															assign node14791 = (inp[0]) ? 4'b1001 : 4'b1000;
														assign node14795 = (inp[2]) ? 4'b1001 : node14796;
															assign node14796 = (inp[0]) ? 4'b1000 : 4'b1001;
												assign node14800 = (inp[10]) ? node14818 : node14801;
													assign node14801 = (inp[2]) ? node14811 : node14802;
														assign node14802 = (inp[11]) ? node14804 : 4'b1101;
															assign node14804 = (inp[0]) ? node14808 : node14805;
																assign node14805 = (inp[9]) ? 4'b1101 : 4'b1100;
																assign node14808 = (inp[9]) ? 4'b1100 : 4'b1101;
														assign node14811 = (inp[11]) ? node14815 : node14812;
															assign node14812 = (inp[9]) ? 4'b1101 : 4'b1100;
															assign node14815 = (inp[9]) ? 4'b1100 : 4'b1101;
													assign node14818 = (inp[0]) ? node14834 : node14819;
														assign node14819 = (inp[9]) ? node14827 : node14820;
															assign node14820 = (inp[2]) ? node14824 : node14821;
																assign node14821 = (inp[11]) ? 4'b1100 : 4'b1101;
																assign node14824 = (inp[11]) ? 4'b1101 : 4'b1100;
															assign node14827 = (inp[11]) ? node14831 : node14828;
																assign node14828 = (inp[2]) ? 4'b1101 : 4'b1100;
																assign node14831 = (inp[2]) ? 4'b1100 : 4'b1101;
														assign node14834 = (inp[9]) ? 4'b1100 : node14835;
															assign node14835 = (inp[11]) ? 4'b1101 : 4'b1100;
										assign node14839 = (inp[1]) ? node14893 : node14840;
											assign node14840 = (inp[4]) ? node14862 : node14841;
												assign node14841 = (inp[9]) ? node14851 : node14842;
													assign node14842 = (inp[11]) ? node14848 : node14843;
														assign node14843 = (inp[0]) ? 4'b1110 : node14844;
															assign node14844 = (inp[2]) ? 4'b1111 : 4'b1110;
														assign node14848 = (inp[2]) ? 4'b1110 : 4'b1111;
													assign node14851 = (inp[11]) ? node14857 : node14852;
														assign node14852 = (inp[0]) ? 4'b1111 : node14853;
															assign node14853 = (inp[2]) ? 4'b1110 : 4'b1111;
														assign node14857 = (inp[0]) ? 4'b1110 : node14858;
															assign node14858 = (inp[2]) ? 4'b1111 : 4'b1110;
												assign node14862 = (inp[2]) ? node14886 : node14863;
													assign node14863 = (inp[0]) ? node14879 : node14864;
														assign node14864 = (inp[10]) ? node14872 : node14865;
															assign node14865 = (inp[11]) ? node14869 : node14866;
																assign node14866 = (inp[9]) ? 4'b1010 : 4'b1011;
																assign node14869 = (inp[9]) ? 4'b1011 : 4'b1010;
															assign node14872 = (inp[9]) ? node14876 : node14873;
																assign node14873 = (inp[11]) ? 4'b1010 : 4'b1011;
																assign node14876 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node14879 = (inp[9]) ? node14883 : node14880;
															assign node14880 = (inp[11]) ? 4'b1011 : 4'b1010;
															assign node14883 = (inp[11]) ? 4'b1010 : 4'b1011;
													assign node14886 = (inp[9]) ? node14890 : node14887;
														assign node14887 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node14890 = (inp[11]) ? 4'b1010 : 4'b1011;
											assign node14893 = (inp[9]) ? node14917 : node14894;
												assign node14894 = (inp[0]) ? node14906 : node14895;
													assign node14895 = (inp[11]) ? node14901 : node14896;
														assign node14896 = (inp[2]) ? node14898 : 4'b1111;
															assign node14898 = (inp[4]) ? 4'b1110 : 4'b1111;
														assign node14901 = (inp[4]) ? node14903 : 4'b1110;
															assign node14903 = (inp[2]) ? 4'b1111 : 4'b1110;
													assign node14906 = (inp[11]) ? node14912 : node14907;
														assign node14907 = (inp[2]) ? node14909 : 4'b1110;
															assign node14909 = (inp[4]) ? 4'b1110 : 4'b1111;
														assign node14912 = (inp[2]) ? node14914 : 4'b1111;
															assign node14914 = (inp[4]) ? 4'b1111 : 4'b1110;
												assign node14917 = (inp[2]) ? node14925 : node14918;
													assign node14918 = (inp[11]) ? node14922 : node14919;
														assign node14919 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node14922 = (inp[0]) ? 4'b1110 : 4'b1111;
													assign node14925 = (inp[0]) ? node14933 : node14926;
														assign node14926 = (inp[11]) ? node14930 : node14927;
															assign node14927 = (inp[4]) ? 4'b1111 : 4'b1110;
															assign node14930 = (inp[4]) ? 4'b1110 : 4'b1111;
														assign node14933 = (inp[4]) ? node14937 : node14934;
															assign node14934 = (inp[11]) ? 4'b1111 : 4'b1110;
															assign node14937 = (inp[11]) ? 4'b1110 : 4'b1111;
									assign node14940 = (inp[7]) ? node15074 : node14941;
										assign node14941 = (inp[1]) ? node14989 : node14942;
											assign node14942 = (inp[4]) ? node14966 : node14943;
												assign node14943 = (inp[11]) ? node14955 : node14944;
													assign node14944 = (inp[9]) ? node14950 : node14945;
														assign node14945 = (inp[0]) ? 4'b1111 : node14946;
															assign node14946 = (inp[2]) ? 4'b1110 : 4'b1111;
														assign node14950 = (inp[0]) ? 4'b1110 : node14951;
															assign node14951 = (inp[2]) ? 4'b1111 : 4'b1110;
													assign node14955 = (inp[9]) ? node14961 : node14956;
														assign node14956 = (inp[0]) ? 4'b1110 : node14957;
															assign node14957 = (inp[2]) ? 4'b1111 : 4'b1110;
														assign node14961 = (inp[0]) ? 4'b1111 : node14962;
															assign node14962 = (inp[2]) ? 4'b1110 : 4'b1111;
												assign node14966 = (inp[9]) ? node14978 : node14967;
													assign node14967 = (inp[11]) ? node14973 : node14968;
														assign node14968 = (inp[0]) ? 4'b1011 : node14969;
															assign node14969 = (inp[2]) ? 4'b1011 : 4'b1010;
														assign node14973 = (inp[2]) ? 4'b1010 : node14974;
															assign node14974 = (inp[0]) ? 4'b1010 : 4'b1011;
													assign node14978 = (inp[11]) ? node14984 : node14979;
														assign node14979 = (inp[0]) ? 4'b1010 : node14980;
															assign node14980 = (inp[2]) ? 4'b1010 : 4'b1011;
														assign node14984 = (inp[0]) ? 4'b1011 : node14985;
															assign node14985 = (inp[2]) ? 4'b1011 : 4'b1010;
											assign node14989 = (inp[4]) ? node15029 : node14990;
												assign node14990 = (inp[0]) ? node15014 : node14991;
													assign node14991 = (inp[9]) ? node15007 : node14992;
														assign node14992 = (inp[10]) ? node15000 : node14993;
															assign node14993 = (inp[2]) ? node14997 : node14994;
																assign node14994 = (inp[11]) ? 4'b1011 : 4'b1010;
																assign node14997 = (inp[11]) ? 4'b1010 : 4'b1011;
															assign node15000 = (inp[11]) ? node15004 : node15001;
																assign node15001 = (inp[2]) ? 4'b1011 : 4'b1010;
																assign node15004 = (inp[2]) ? 4'b1010 : 4'b1011;
														assign node15007 = (inp[11]) ? node15011 : node15008;
															assign node15008 = (inp[2]) ? 4'b1010 : 4'b1011;
															assign node15011 = (inp[2]) ? 4'b1011 : 4'b1010;
													assign node15014 = (inp[2]) ? node15022 : node15015;
														assign node15015 = (inp[11]) ? node15019 : node15016;
															assign node15016 = (inp[9]) ? 4'b1011 : 4'b1010;
															assign node15019 = (inp[9]) ? 4'b1010 : 4'b1011;
														assign node15022 = (inp[9]) ? node15026 : node15023;
															assign node15023 = (inp[11]) ? 4'b1011 : 4'b1010;
															assign node15026 = (inp[11]) ? 4'b1010 : 4'b1011;
												assign node15029 = (inp[2]) ? node15053 : node15030;
													assign node15030 = (inp[10]) ? node15038 : node15031;
														assign node15031 = (inp[11]) ? node15035 : node15032;
															assign node15032 = (inp[9]) ? 4'b1111 : 4'b1110;
															assign node15035 = (inp[9]) ? 4'b1110 : 4'b1111;
														assign node15038 = (inp[0]) ? node15046 : node15039;
															assign node15039 = (inp[9]) ? node15043 : node15040;
																assign node15040 = (inp[11]) ? 4'b1111 : 4'b1110;
																assign node15043 = (inp[11]) ? 4'b1110 : 4'b1111;
															assign node15046 = (inp[11]) ? node15050 : node15047;
																assign node15047 = (inp[9]) ? 4'b1111 : 4'b1110;
																assign node15050 = (inp[9]) ? 4'b1110 : 4'b1111;
													assign node15053 = (inp[11]) ? node15067 : node15054;
														assign node15054 = (inp[10]) ? node15060 : node15055;
															assign node15055 = (inp[9]) ? node15057 : 4'b1110;
																assign node15057 = (inp[0]) ? 4'b1110 : 4'b1111;
															assign node15060 = (inp[9]) ? node15064 : node15061;
																assign node15061 = (inp[0]) ? 4'b1111 : 4'b1110;
																assign node15064 = (inp[0]) ? 4'b1110 : 4'b1111;
														assign node15067 = (inp[0]) ? node15071 : node15068;
															assign node15068 = (inp[9]) ? 4'b1110 : 4'b1111;
															assign node15071 = (inp[9]) ? 4'b1111 : 4'b1110;
										assign node15074 = (inp[4]) ? node15122 : node15075;
											assign node15075 = (inp[1]) ? node15101 : node15076;
												assign node15076 = (inp[2]) ? node15094 : node15077;
													assign node15077 = (inp[9]) ? node15087 : node15078;
														assign node15078 = (inp[10]) ? 4'b1101 : node15079;
															assign node15079 = (inp[11]) ? node15083 : node15080;
																assign node15080 = (inp[0]) ? 4'b1101 : 4'b1100;
																assign node15083 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node15087 = (inp[0]) ? node15091 : node15088;
															assign node15088 = (inp[11]) ? 4'b1100 : 4'b1101;
															assign node15091 = (inp[11]) ? 4'b1101 : 4'b1100;
													assign node15094 = (inp[11]) ? node15098 : node15095;
														assign node15095 = (inp[9]) ? 4'b1101 : 4'b1100;
														assign node15098 = (inp[9]) ? 4'b1100 : 4'b1101;
												assign node15101 = (inp[11]) ? node15113 : node15102;
													assign node15102 = (inp[9]) ? node15108 : node15103;
														assign node15103 = (inp[2]) ? 4'b1001 : node15104;
															assign node15104 = (inp[0]) ? 4'b1000 : 4'b1001;
														assign node15108 = (inp[2]) ? 4'b1000 : node15109;
															assign node15109 = (inp[0]) ? 4'b1001 : 4'b1000;
													assign node15113 = (inp[9]) ? node15117 : node15114;
														assign node15114 = (inp[2]) ? 4'b1000 : 4'b1001;
														assign node15117 = (inp[0]) ? node15119 : 4'b1001;
															assign node15119 = (inp[2]) ? 4'b1001 : 4'b1000;
											assign node15122 = (inp[1]) ? node15168 : node15123;
												assign node15123 = (inp[10]) ? node15145 : node15124;
													assign node15124 = (inp[11]) ? node15134 : node15125;
														assign node15125 = (inp[9]) ? node15131 : node15126;
															assign node15126 = (inp[0]) ? node15128 : 4'b1000;
																assign node15128 = (inp[2]) ? 4'b1001 : 4'b1000;
															assign node15131 = (inp[2]) ? 4'b1000 : 4'b1001;
														assign node15134 = (inp[9]) ? node15140 : node15135;
															assign node15135 = (inp[0]) ? node15137 : 4'b1001;
																assign node15137 = (inp[2]) ? 4'b1000 : 4'b1001;
															assign node15140 = (inp[2]) ? node15142 : 4'b1000;
																assign node15142 = (inp[0]) ? 4'b1001 : 4'b1000;
													assign node15145 = (inp[2]) ? node15153 : node15146;
														assign node15146 = (inp[11]) ? node15150 : node15147;
															assign node15147 = (inp[9]) ? 4'b1001 : 4'b1000;
															assign node15150 = (inp[9]) ? 4'b1000 : 4'b1001;
														assign node15153 = (inp[0]) ? node15161 : node15154;
															assign node15154 = (inp[9]) ? node15158 : node15155;
																assign node15155 = (inp[11]) ? 4'b1001 : 4'b1000;
																assign node15158 = (inp[11]) ? 4'b1000 : 4'b1001;
															assign node15161 = (inp[9]) ? node15165 : node15162;
																assign node15162 = (inp[11]) ? 4'b1000 : 4'b1001;
																assign node15165 = (inp[11]) ? 4'b1001 : 4'b1000;
												assign node15168 = (inp[9]) ? node15180 : node15169;
													assign node15169 = (inp[11]) ? node15175 : node15170;
														assign node15170 = (inp[2]) ? 4'b1100 : node15171;
															assign node15171 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node15175 = (inp[2]) ? 4'b1101 : node15176;
															assign node15176 = (inp[0]) ? 4'b1101 : 4'b1100;
													assign node15180 = (inp[11]) ? node15186 : node15181;
														assign node15181 = (inp[0]) ? 4'b1101 : node15182;
															assign node15182 = (inp[2]) ? 4'b1101 : 4'b1100;
														assign node15186 = (inp[0]) ? 4'b1100 : node15187;
															assign node15187 = (inp[2]) ? 4'b1100 : 4'b1101;
								assign node15191 = (inp[15]) ? node15453 : node15192;
									assign node15192 = (inp[7]) ? node15300 : node15193;
										assign node15193 = (inp[4]) ? node15241 : node15194;
											assign node15194 = (inp[9]) ? node15218 : node15195;
												assign node15195 = (inp[11]) ? node15207 : node15196;
													assign node15196 = (inp[1]) ? node15202 : node15197;
														assign node15197 = (inp[0]) ? 4'b1100 : node15198;
															assign node15198 = (inp[2]) ? 4'b1101 : 4'b1100;
														assign node15202 = (inp[2]) ? 4'b1100 : node15203;
															assign node15203 = (inp[0]) ? 4'b1101 : 4'b1100;
													assign node15207 = (inp[2]) ? node15213 : node15208;
														assign node15208 = (inp[0]) ? node15210 : 4'b1101;
															assign node15210 = (inp[1]) ? 4'b1100 : 4'b1101;
														assign node15213 = (inp[0]) ? 4'b1101 : node15214;
															assign node15214 = (inp[1]) ? 4'b1101 : 4'b1100;
												assign node15218 = (inp[11]) ? node15230 : node15219;
													assign node15219 = (inp[2]) ? node15225 : node15220;
														assign node15220 = (inp[0]) ? node15222 : 4'b1101;
															assign node15222 = (inp[1]) ? 4'b1100 : 4'b1101;
														assign node15225 = (inp[0]) ? 4'b1101 : node15226;
															assign node15226 = (inp[1]) ? 4'b1101 : 4'b1100;
													assign node15230 = (inp[1]) ? node15236 : node15231;
														assign node15231 = (inp[0]) ? 4'b1100 : node15232;
															assign node15232 = (inp[2]) ? 4'b1101 : 4'b1100;
														assign node15236 = (inp[0]) ? node15238 : 4'b1100;
															assign node15238 = (inp[2]) ? 4'b1100 : 4'b1101;
											assign node15241 = (inp[1]) ? node15263 : node15242;
												assign node15242 = (inp[11]) ? node15252 : node15243;
													assign node15243 = (inp[9]) ? node15247 : node15244;
														assign node15244 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node15247 = (inp[0]) ? 4'b1101 : node15248;
															assign node15248 = (inp[2]) ? 4'b1101 : 4'b1100;
													assign node15252 = (inp[9]) ? node15258 : node15253;
														assign node15253 = (inp[0]) ? 4'b1101 : node15254;
															assign node15254 = (inp[2]) ? 4'b1101 : 4'b1100;
														assign node15258 = (inp[0]) ? 4'b1100 : node15259;
															assign node15259 = (inp[2]) ? 4'b1100 : 4'b1101;
												assign node15263 = (inp[2]) ? node15271 : node15264;
													assign node15264 = (inp[11]) ? node15268 : node15265;
														assign node15265 = (inp[9]) ? 4'b1001 : 4'b1000;
														assign node15268 = (inp[9]) ? 4'b1000 : 4'b1001;
													assign node15271 = (inp[10]) ? node15285 : node15272;
														assign node15272 = (inp[0]) ? node15280 : node15273;
															assign node15273 = (inp[9]) ? node15277 : node15274;
																assign node15274 = (inp[11]) ? 4'b1001 : 4'b1000;
																assign node15277 = (inp[11]) ? 4'b1000 : 4'b1001;
															assign node15280 = (inp[9]) ? node15282 : 4'b1000;
																assign node15282 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node15285 = (inp[9]) ? node15293 : node15286;
															assign node15286 = (inp[11]) ? node15290 : node15287;
																assign node15287 = (inp[0]) ? 4'b1001 : 4'b1000;
																assign node15290 = (inp[0]) ? 4'b1000 : 4'b1001;
															assign node15293 = (inp[0]) ? node15297 : node15294;
																assign node15294 = (inp[11]) ? 4'b1000 : 4'b1001;
																assign node15297 = (inp[11]) ? 4'b1001 : 4'b1000;
										assign node15300 = (inp[4]) ? node15366 : node15301;
											assign node15301 = (inp[1]) ? node15343 : node15302;
												assign node15302 = (inp[0]) ? node15320 : node15303;
													assign node15303 = (inp[10]) ? node15311 : node15304;
														assign node15304 = (inp[2]) ? 4'b1011 : node15305;
															assign node15305 = (inp[11]) ? 4'b1010 : node15306;
																assign node15306 = (inp[9]) ? 4'b1010 : 4'b1011;
														assign node15311 = (inp[2]) ? node15313 : 4'b1011;
															assign node15313 = (inp[9]) ? node15317 : node15314;
																assign node15314 = (inp[11]) ? 4'b1011 : 4'b1010;
																assign node15317 = (inp[11]) ? 4'b1010 : 4'b1011;
													assign node15320 = (inp[2]) ? node15330 : node15321;
														assign node15321 = (inp[10]) ? 4'b1011 : node15322;
															assign node15322 = (inp[11]) ? node15326 : node15323;
																assign node15323 = (inp[9]) ? 4'b1010 : 4'b1011;
																assign node15326 = (inp[9]) ? 4'b1011 : 4'b1010;
														assign node15330 = (inp[10]) ? node15338 : node15331;
															assign node15331 = (inp[11]) ? node15335 : node15332;
																assign node15332 = (inp[9]) ? 4'b1010 : 4'b1011;
																assign node15335 = (inp[9]) ? 4'b1011 : 4'b1010;
															assign node15338 = (inp[9]) ? node15340 : 4'b1010;
																assign node15340 = (inp[11]) ? 4'b1011 : 4'b1010;
												assign node15343 = (inp[11]) ? node15355 : node15344;
													assign node15344 = (inp[9]) ? node15350 : node15345;
														assign node15345 = (inp[2]) ? node15347 : 4'b1110;
															assign node15347 = (inp[0]) ? 4'b1110 : 4'b1111;
														assign node15350 = (inp[0]) ? 4'b1111 : node15351;
															assign node15351 = (inp[2]) ? 4'b1110 : 4'b1111;
													assign node15355 = (inp[9]) ? node15361 : node15356;
														assign node15356 = (inp[0]) ? 4'b1111 : node15357;
															assign node15357 = (inp[2]) ? 4'b1110 : 4'b1111;
														assign node15361 = (inp[0]) ? 4'b1110 : node15362;
															assign node15362 = (inp[2]) ? 4'b1111 : 4'b1110;
											assign node15366 = (inp[10]) ? node15410 : node15367;
												assign node15367 = (inp[1]) ? node15391 : node15368;
													assign node15368 = (inp[2]) ? node15376 : node15369;
														assign node15369 = (inp[11]) ? node15373 : node15370;
															assign node15370 = (inp[9]) ? 4'b1110 : 4'b1111;
															assign node15373 = (inp[9]) ? 4'b1111 : 4'b1110;
														assign node15376 = (inp[9]) ? node15384 : node15377;
															assign node15377 = (inp[0]) ? node15381 : node15378;
																assign node15378 = (inp[11]) ? 4'b1110 : 4'b1111;
																assign node15381 = (inp[11]) ? 4'b1111 : 4'b1110;
															assign node15384 = (inp[11]) ? node15388 : node15385;
																assign node15385 = (inp[0]) ? 4'b1111 : 4'b1110;
																assign node15388 = (inp[0]) ? 4'b1110 : 4'b1111;
													assign node15391 = (inp[9]) ? node15403 : node15392;
														assign node15392 = (inp[11]) ? node15398 : node15393;
															assign node15393 = (inp[2]) ? 4'b1110 : node15394;
																assign node15394 = (inp[0]) ? 4'b1110 : 4'b1111;
															assign node15398 = (inp[2]) ? 4'b1111 : node15399;
																assign node15399 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node15403 = (inp[11]) ? 4'b1110 : node15404;
															assign node15404 = (inp[2]) ? 4'b1111 : node15405;
																assign node15405 = (inp[0]) ? 4'b1111 : 4'b1110;
												assign node15410 = (inp[0]) ? node15434 : node15411;
													assign node15411 = (inp[1]) ? node15419 : node15412;
														assign node15412 = (inp[9]) ? node15416 : node15413;
															assign node15413 = (inp[11]) ? 4'b1110 : 4'b1111;
															assign node15416 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node15419 = (inp[9]) ? node15427 : node15420;
															assign node15420 = (inp[2]) ? node15424 : node15421;
																assign node15421 = (inp[11]) ? 4'b1110 : 4'b1111;
																assign node15424 = (inp[11]) ? 4'b1111 : 4'b1110;
															assign node15427 = (inp[11]) ? node15431 : node15428;
																assign node15428 = (inp[2]) ? 4'b1111 : 4'b1110;
																assign node15431 = (inp[2]) ? 4'b1110 : 4'b1111;
													assign node15434 = (inp[9]) ? node15442 : node15435;
														assign node15435 = (inp[11]) ? node15437 : 4'b1110;
															assign node15437 = (inp[1]) ? 4'b1111 : node15438;
																assign node15438 = (inp[2]) ? 4'b1111 : 4'b1110;
														assign node15442 = (inp[11]) ? node15448 : node15443;
															assign node15443 = (inp[2]) ? 4'b1111 : node15444;
																assign node15444 = (inp[1]) ? 4'b1111 : 4'b1110;
															assign node15448 = (inp[2]) ? 4'b1110 : node15449;
																assign node15449 = (inp[1]) ? 4'b1110 : 4'b1111;
									assign node15453 = (inp[7]) ? node15613 : node15454;
										assign node15454 = (inp[0]) ? node15556 : node15455;
											assign node15455 = (inp[10]) ? node15503 : node15456;
												assign node15456 = (inp[2]) ? node15486 : node15457;
													assign node15457 = (inp[1]) ? node15473 : node15458;
														assign node15458 = (inp[9]) ? node15466 : node15459;
															assign node15459 = (inp[11]) ? node15463 : node15460;
																assign node15460 = (inp[4]) ? 4'b1110 : 4'b1111;
																assign node15463 = (inp[4]) ? 4'b1111 : 4'b1110;
															assign node15466 = (inp[11]) ? node15470 : node15467;
																assign node15467 = (inp[4]) ? 4'b1111 : 4'b1110;
																assign node15470 = (inp[4]) ? 4'b1110 : 4'b1111;
														assign node15473 = (inp[4]) ? node15479 : node15474;
															assign node15474 = (inp[9]) ? node15476 : 4'b1110;
																assign node15476 = (inp[11]) ? 4'b1111 : 4'b1110;
															assign node15479 = (inp[9]) ? node15483 : node15480;
																assign node15480 = (inp[11]) ? 4'b1111 : 4'b1110;
																assign node15483 = (inp[11]) ? 4'b1110 : 4'b1111;
													assign node15486 = (inp[4]) ? node15494 : node15487;
														assign node15487 = (inp[11]) ? node15491 : node15488;
															assign node15488 = (inp[9]) ? 4'b1111 : 4'b1110;
															assign node15491 = (inp[9]) ? 4'b1110 : 4'b1111;
														assign node15494 = (inp[1]) ? node15496 : 4'b1110;
															assign node15496 = (inp[11]) ? node15500 : node15497;
																assign node15497 = (inp[9]) ? 4'b1110 : 4'b1111;
																assign node15500 = (inp[9]) ? 4'b1111 : 4'b1110;
												assign node15503 = (inp[1]) ? node15529 : node15504;
													assign node15504 = (inp[11]) ? node15514 : node15505;
														assign node15505 = (inp[9]) ? node15507 : 4'b1111;
															assign node15507 = (inp[2]) ? node15511 : node15508;
																assign node15508 = (inp[4]) ? 4'b1111 : 4'b1110;
																assign node15511 = (inp[4]) ? 4'b1110 : 4'b1111;
														assign node15514 = (inp[2]) ? node15522 : node15515;
															assign node15515 = (inp[4]) ? node15519 : node15516;
																assign node15516 = (inp[9]) ? 4'b1111 : 4'b1110;
																assign node15519 = (inp[9]) ? 4'b1110 : 4'b1111;
															assign node15522 = (inp[9]) ? node15526 : node15523;
																assign node15523 = (inp[4]) ? 4'b1110 : 4'b1111;
																assign node15526 = (inp[4]) ? 4'b1111 : 4'b1110;
													assign node15529 = (inp[4]) ? node15543 : node15530;
														assign node15530 = (inp[9]) ? node15538 : node15531;
															assign node15531 = (inp[11]) ? node15535 : node15532;
																assign node15532 = (inp[2]) ? 4'b1110 : 4'b1111;
																assign node15535 = (inp[2]) ? 4'b1111 : 4'b1110;
															assign node15538 = (inp[2]) ? node15540 : 4'b1110;
																assign node15540 = (inp[11]) ? 4'b1110 : 4'b1111;
														assign node15543 = (inp[11]) ? node15549 : node15544;
															assign node15544 = (inp[9]) ? node15546 : 4'b1110;
																assign node15546 = (inp[2]) ? 4'b1110 : 4'b1111;
															assign node15549 = (inp[2]) ? node15553 : node15550;
																assign node15550 = (inp[9]) ? 4'b1110 : 4'b1111;
																assign node15553 = (inp[9]) ? 4'b1111 : 4'b1110;
											assign node15556 = (inp[1]) ? node15580 : node15557;
												assign node15557 = (inp[2]) ? node15565 : node15558;
													assign node15558 = (inp[11]) ? node15562 : node15559;
														assign node15559 = (inp[9]) ? 4'b1110 : 4'b1111;
														assign node15562 = (inp[9]) ? 4'b1111 : 4'b1110;
													assign node15565 = (inp[4]) ? node15573 : node15566;
														assign node15566 = (inp[9]) ? node15570 : node15567;
															assign node15567 = (inp[11]) ? 4'b1110 : 4'b1111;
															assign node15570 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node15573 = (inp[10]) ? 4'b1110 : node15574;
															assign node15574 = (inp[9]) ? 4'b1110 : node15575;
																assign node15575 = (inp[11]) ? 4'b1110 : 4'b1111;
												assign node15580 = (inp[2]) ? node15590 : node15581;
													assign node15581 = (inp[10]) ? node15583 : 4'b1111;
														assign node15583 = (inp[11]) ? node15587 : node15584;
															assign node15584 = (inp[9]) ? 4'b1110 : 4'b1111;
															assign node15587 = (inp[9]) ? 4'b1111 : 4'b1110;
													assign node15590 = (inp[10]) ? node15606 : node15591;
														assign node15591 = (inp[4]) ? node15599 : node15592;
															assign node15592 = (inp[11]) ? node15596 : node15593;
																assign node15593 = (inp[9]) ? 4'b1110 : 4'b1111;
																assign node15596 = (inp[9]) ? 4'b1111 : 4'b1110;
															assign node15599 = (inp[11]) ? node15603 : node15600;
																assign node15600 = (inp[9]) ? 4'b1110 : 4'b1111;
																assign node15603 = (inp[9]) ? 4'b1111 : 4'b1110;
														assign node15606 = (inp[11]) ? node15610 : node15607;
															assign node15607 = (inp[9]) ? 4'b1110 : 4'b1111;
															assign node15610 = (inp[9]) ? 4'b1111 : 4'b1110;
										assign node15613 = (inp[9]) ? node15639 : node15614;
											assign node15614 = (inp[11]) ? node15624 : node15615;
												assign node15615 = (inp[0]) ? 4'b1100 : node15616;
													assign node15616 = (inp[2]) ? node15620 : node15617;
														assign node15617 = (inp[4]) ? 4'b1101 : 4'b1100;
														assign node15620 = (inp[4]) ? 4'b1100 : 4'b1101;
												assign node15624 = (inp[0]) ? 4'b1101 : node15625;
													assign node15625 = (inp[1]) ? node15633 : node15626;
														assign node15626 = (inp[2]) ? node15630 : node15627;
															assign node15627 = (inp[4]) ? 4'b1100 : 4'b1101;
															assign node15630 = (inp[4]) ? 4'b1101 : 4'b1100;
														assign node15633 = (inp[4]) ? 4'b1100 : node15634;
															assign node15634 = (inp[2]) ? 4'b1100 : 4'b1101;
											assign node15639 = (inp[11]) ? node15657 : node15640;
												assign node15640 = (inp[0]) ? 4'b1101 : node15641;
													assign node15641 = (inp[1]) ? node15649 : node15642;
														assign node15642 = (inp[2]) ? node15646 : node15643;
															assign node15643 = (inp[4]) ? 4'b1100 : 4'b1101;
															assign node15646 = (inp[4]) ? 4'b1101 : 4'b1100;
														assign node15649 = (inp[4]) ? node15653 : node15650;
															assign node15650 = (inp[2]) ? 4'b1100 : 4'b1101;
															assign node15653 = (inp[2]) ? 4'b1101 : 4'b1100;
												assign node15657 = (inp[0]) ? 4'b1100 : node15658;
													assign node15658 = (inp[1]) ? node15672 : node15659;
														assign node15659 = (inp[10]) ? node15665 : node15660;
															assign node15660 = (inp[4]) ? node15662 : 4'b1101;
																assign node15662 = (inp[2]) ? 4'b1100 : 4'b1101;
															assign node15665 = (inp[4]) ? node15669 : node15666;
																assign node15666 = (inp[2]) ? 4'b1101 : 4'b1100;
																assign node15669 = (inp[2]) ? 4'b1100 : 4'b1101;
														assign node15672 = (inp[10]) ? node15680 : node15673;
															assign node15673 = (inp[4]) ? node15677 : node15674;
																assign node15674 = (inp[2]) ? 4'b1101 : 4'b1100;
																assign node15677 = (inp[2]) ? 4'b1100 : 4'b1101;
															assign node15680 = (inp[4]) ? node15684 : node15681;
																assign node15681 = (inp[2]) ? 4'b1101 : 4'b1100;
																assign node15684 = (inp[2]) ? 4'b1100 : 4'b1101;
						assign node15688 = (inp[6]) ? node17004 : node15689;
							assign node15689 = (inp[2]) ? node16333 : node15690;
								assign node15690 = (inp[7]) ? node16042 : node15691;
									assign node15691 = (inp[12]) ? node15869 : node15692;
										assign node15692 = (inp[15]) ? node15784 : node15693;
											assign node15693 = (inp[4]) ? node15737 : node15694;
												assign node15694 = (inp[9]) ? node15718 : node15695;
													assign node15695 = (inp[10]) ? node15707 : node15696;
														assign node15696 = (inp[11]) ? node15702 : node15697;
															assign node15697 = (inp[0]) ? 4'b1100 : node15698;
																assign node15698 = (inp[1]) ? 4'b1101 : 4'b1100;
															assign node15702 = (inp[1]) ? 4'b1101 : node15703;
																assign node15703 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node15707 = (inp[0]) ? node15713 : node15708;
															assign node15708 = (inp[11]) ? 4'b1100 : node15709;
																assign node15709 = (inp[1]) ? 4'b1100 : 4'b1101;
															assign node15713 = (inp[11]) ? node15715 : 4'b1101;
																assign node15715 = (inp[1]) ? 4'b1100 : 4'b1101;
													assign node15718 = (inp[0]) ? node15728 : node15719;
														assign node15719 = (inp[11]) ? 4'b1100 : node15720;
															assign node15720 = (inp[1]) ? node15724 : node15721;
																assign node15721 = (inp[10]) ? 4'b1100 : 4'b1101;
																assign node15724 = (inp[10]) ? 4'b1101 : 4'b1100;
														assign node15728 = (inp[10]) ? node15732 : node15729;
															assign node15729 = (inp[1]) ? 4'b1100 : 4'b1101;
															assign node15732 = (inp[11]) ? node15734 : 4'b1100;
																assign node15734 = (inp[1]) ? 4'b1101 : 4'b1100;
												assign node15737 = (inp[10]) ? node15761 : node15738;
													assign node15738 = (inp[9]) ? node15750 : node15739;
														assign node15739 = (inp[1]) ? node15745 : node15740;
															assign node15740 = (inp[0]) ? node15742 : 4'b1111;
																assign node15742 = (inp[11]) ? 4'b1111 : 4'b1110;
															assign node15745 = (inp[11]) ? node15747 : 4'b1111;
																assign node15747 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node15750 = (inp[0]) ? node15756 : node15751;
															assign node15751 = (inp[11]) ? node15753 : 4'b1110;
																assign node15753 = (inp[1]) ? 4'b1111 : 4'b1110;
															assign node15756 = (inp[11]) ? 4'b1110 : node15757;
																assign node15757 = (inp[1]) ? 4'b1110 : 4'b1111;
													assign node15761 = (inp[9]) ? node15773 : node15762;
														assign node15762 = (inp[1]) ? node15768 : node15763;
															assign node15763 = (inp[11]) ? 4'b1110 : node15764;
																assign node15764 = (inp[0]) ? 4'b1111 : 4'b1110;
															assign node15768 = (inp[0]) ? 4'b1110 : node15769;
																assign node15769 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node15773 = (inp[11]) ? node15779 : node15774;
															assign node15774 = (inp[0]) ? node15776 : 4'b1111;
																assign node15776 = (inp[1]) ? 4'b1111 : 4'b1110;
															assign node15779 = (inp[0]) ? 4'b1111 : node15780;
																assign node15780 = (inp[1]) ? 4'b1110 : 4'b1111;
											assign node15784 = (inp[4]) ? node15826 : node15785;
												assign node15785 = (inp[11]) ? node15801 : node15786;
													assign node15786 = (inp[9]) ? node15794 : node15787;
														assign node15787 = (inp[10]) ? node15791 : node15788;
															assign node15788 = (inp[1]) ? 4'b1100 : 4'b1101;
															assign node15791 = (inp[1]) ? 4'b1101 : 4'b1100;
														assign node15794 = (inp[1]) ? node15798 : node15795;
															assign node15795 = (inp[10]) ? 4'b1101 : 4'b1100;
															assign node15798 = (inp[10]) ? 4'b1100 : 4'b1101;
													assign node15801 = (inp[1]) ? node15817 : node15802;
														assign node15802 = (inp[10]) ? node15810 : node15803;
															assign node15803 = (inp[0]) ? node15807 : node15804;
																assign node15804 = (inp[9]) ? 4'b1101 : 4'b1100;
																assign node15807 = (inp[9]) ? 4'b1100 : 4'b1101;
															assign node15810 = (inp[0]) ? node15814 : node15811;
																assign node15811 = (inp[9]) ? 4'b1100 : 4'b1101;
																assign node15814 = (inp[9]) ? 4'b1101 : 4'b1100;
														assign node15817 = (inp[9]) ? node15819 : 4'b1101;
															assign node15819 = (inp[0]) ? node15823 : node15820;
																assign node15820 = (inp[10]) ? 4'b1101 : 4'b1100;
																assign node15823 = (inp[10]) ? 4'b1100 : 4'b1101;
												assign node15826 = (inp[1]) ? node15848 : node15827;
													assign node15827 = (inp[9]) ? node15839 : node15828;
														assign node15828 = (inp[10]) ? node15834 : node15829;
															assign node15829 = (inp[0]) ? 4'b1000 : node15830;
																assign node15830 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node15834 = (inp[0]) ? 4'b1001 : node15835;
																assign node15835 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node15839 = (inp[10]) ? node15845 : node15840;
															assign node15840 = (inp[11]) ? node15842 : 4'b1001;
																assign node15842 = (inp[0]) ? 4'b1001 : 4'b1000;
															assign node15845 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node15848 = (inp[0]) ? node15862 : node15849;
														assign node15849 = (inp[10]) ? node15857 : node15850;
															assign node15850 = (inp[11]) ? node15854 : node15851;
																assign node15851 = (inp[9]) ? 4'b1000 : 4'b1001;
																assign node15854 = (inp[9]) ? 4'b1001 : 4'b1000;
															assign node15857 = (inp[9]) ? 4'b1000 : node15858;
																assign node15858 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node15862 = (inp[10]) ? node15866 : node15863;
															assign node15863 = (inp[9]) ? 4'b1000 : 4'b1001;
															assign node15866 = (inp[9]) ? 4'b1001 : 4'b1000;
										assign node15869 = (inp[15]) ? node15963 : node15870;
											assign node15870 = (inp[4]) ? node15908 : node15871;
												assign node15871 = (inp[11]) ? node15887 : node15872;
													assign node15872 = (inp[0]) ? node15880 : node15873;
														assign node15873 = (inp[10]) ? node15877 : node15874;
															assign node15874 = (inp[9]) ? 4'b1111 : 4'b1110;
															assign node15877 = (inp[9]) ? 4'b1110 : 4'b1111;
														assign node15880 = (inp[1]) ? node15882 : 4'b1111;
															assign node15882 = (inp[9]) ? node15884 : 4'b1111;
																assign node15884 = (inp[10]) ? 4'b1111 : 4'b1110;
													assign node15887 = (inp[1]) ? node15901 : node15888;
														assign node15888 = (inp[0]) ? node15894 : node15889;
															assign node15889 = (inp[10]) ? node15891 : 4'b1110;
																assign node15891 = (inp[9]) ? 4'b1111 : 4'b1110;
															assign node15894 = (inp[10]) ? node15898 : node15895;
																assign node15895 = (inp[9]) ? 4'b1111 : 4'b1110;
																assign node15898 = (inp[9]) ? 4'b1110 : 4'b1111;
														assign node15901 = (inp[9]) ? node15905 : node15902;
															assign node15902 = (inp[10]) ? 4'b1111 : 4'b1110;
															assign node15905 = (inp[10]) ? 4'b1110 : 4'b1111;
												assign node15908 = (inp[1]) ? node15940 : node15909;
													assign node15909 = (inp[11]) ? node15925 : node15910;
														assign node15910 = (inp[0]) ? node15918 : node15911;
															assign node15911 = (inp[10]) ? node15915 : node15912;
																assign node15912 = (inp[9]) ? 4'b1100 : 4'b1101;
																assign node15915 = (inp[9]) ? 4'b1101 : 4'b1100;
															assign node15918 = (inp[10]) ? node15922 : node15919;
																assign node15919 = (inp[9]) ? 4'b1100 : 4'b1101;
																assign node15922 = (inp[9]) ? 4'b1101 : 4'b1100;
														assign node15925 = (inp[10]) ? node15933 : node15926;
															assign node15926 = (inp[0]) ? node15930 : node15927;
																assign node15927 = (inp[9]) ? 4'b1101 : 4'b1100;
																assign node15930 = (inp[9]) ? 4'b1100 : 4'b1101;
															assign node15933 = (inp[9]) ? node15937 : node15934;
																assign node15934 = (inp[0]) ? 4'b1100 : 4'b1101;
																assign node15937 = (inp[0]) ? 4'b1101 : 4'b1100;
													assign node15940 = (inp[11]) ? node15956 : node15941;
														assign node15941 = (inp[10]) ? node15949 : node15942;
															assign node15942 = (inp[9]) ? node15946 : node15943;
																assign node15943 = (inp[0]) ? 4'b1000 : 4'b1001;
																assign node15946 = (inp[0]) ? 4'b1001 : 4'b1000;
															assign node15949 = (inp[0]) ? node15953 : node15950;
																assign node15950 = (inp[9]) ? 4'b1001 : 4'b1000;
																assign node15953 = (inp[9]) ? 4'b1000 : 4'b1001;
														assign node15956 = (inp[9]) ? node15960 : node15957;
															assign node15957 = (inp[10]) ? 4'b1000 : 4'b1001;
															assign node15960 = (inp[10]) ? 4'b1001 : 4'b1000;
											assign node15963 = (inp[4]) ? node16017 : node15964;
												assign node15964 = (inp[0]) ? node15994 : node15965;
													assign node15965 = (inp[1]) ? node15981 : node15966;
														assign node15966 = (inp[9]) ? node15974 : node15967;
															assign node15967 = (inp[10]) ? node15971 : node15968;
																assign node15968 = (inp[11]) ? 4'b1110 : 4'b1111;
																assign node15971 = (inp[11]) ? 4'b1111 : 4'b1110;
															assign node15974 = (inp[11]) ? node15978 : node15975;
																assign node15975 = (inp[10]) ? 4'b1111 : 4'b1110;
																assign node15978 = (inp[10]) ? 4'b1110 : 4'b1111;
														assign node15981 = (inp[10]) ? node15989 : node15982;
															assign node15982 = (inp[11]) ? node15986 : node15983;
																assign node15983 = (inp[9]) ? 4'b1110 : 4'b1111;
																assign node15986 = (inp[9]) ? 4'b1111 : 4'b1110;
															assign node15989 = (inp[9]) ? node15991 : 4'b1110;
																assign node15991 = (inp[11]) ? 4'b1110 : 4'b1111;
													assign node15994 = (inp[11]) ? node16010 : node15995;
														assign node15995 = (inp[1]) ? node16003 : node15996;
															assign node15996 = (inp[10]) ? node16000 : node15997;
																assign node15997 = (inp[9]) ? 4'b1110 : 4'b1111;
																assign node16000 = (inp[9]) ? 4'b1111 : 4'b1110;
															assign node16003 = (inp[10]) ? node16007 : node16004;
																assign node16004 = (inp[9]) ? 4'b1110 : 4'b1111;
																assign node16007 = (inp[9]) ? 4'b1111 : 4'b1110;
														assign node16010 = (inp[9]) ? node16014 : node16011;
															assign node16011 = (inp[10]) ? 4'b1110 : 4'b1111;
															assign node16014 = (inp[10]) ? 4'b1111 : 4'b1110;
												assign node16017 = (inp[11]) ? node16025 : node16018;
													assign node16018 = (inp[9]) ? node16022 : node16019;
														assign node16019 = (inp[10]) ? 4'b1111 : 4'b1110;
														assign node16022 = (inp[10]) ? 4'b1110 : 4'b1111;
													assign node16025 = (inp[0]) ? node16035 : node16026;
														assign node16026 = (inp[1]) ? node16032 : node16027;
															assign node16027 = (inp[9]) ? node16029 : 4'b1111;
																assign node16029 = (inp[10]) ? 4'b1111 : 4'b1110;
															assign node16032 = (inp[9]) ? 4'b1111 : 4'b1110;
														assign node16035 = (inp[10]) ? node16039 : node16036;
															assign node16036 = (inp[9]) ? 4'b1111 : 4'b1110;
															assign node16039 = (inp[9]) ? 4'b1110 : 4'b1111;
									assign node16042 = (inp[12]) ? node16202 : node16043;
										assign node16043 = (inp[4]) ? node16131 : node16044;
											assign node16044 = (inp[0]) ? node16076 : node16045;
												assign node16045 = (inp[10]) ? node16061 : node16046;
													assign node16046 = (inp[9]) ? node16054 : node16047;
														assign node16047 = (inp[1]) ? node16051 : node16048;
															assign node16048 = (inp[15]) ? 4'b1111 : 4'b1010;
															assign node16051 = (inp[15]) ? 4'b1010 : 4'b1110;
														assign node16054 = (inp[15]) ? node16058 : node16055;
															assign node16055 = (inp[1]) ? 4'b1111 : 4'b1011;
															assign node16058 = (inp[1]) ? 4'b1011 : 4'b1110;
													assign node16061 = (inp[9]) ? node16069 : node16062;
														assign node16062 = (inp[1]) ? node16066 : node16063;
															assign node16063 = (inp[15]) ? 4'b1110 : 4'b1011;
															assign node16066 = (inp[15]) ? 4'b1011 : 4'b1111;
														assign node16069 = (inp[15]) ? node16073 : node16070;
															assign node16070 = (inp[1]) ? 4'b1110 : 4'b1010;
															assign node16073 = (inp[1]) ? 4'b1010 : 4'b1111;
												assign node16076 = (inp[1]) ? node16106 : node16077;
													assign node16077 = (inp[15]) ? node16091 : node16078;
														assign node16078 = (inp[9]) ? node16086 : node16079;
															assign node16079 = (inp[10]) ? node16083 : node16080;
																assign node16080 = (inp[11]) ? 4'b1010 : 4'b1011;
																assign node16083 = (inp[11]) ? 4'b1011 : 4'b1010;
															assign node16086 = (inp[10]) ? node16088 : 4'b1010;
																assign node16088 = (inp[11]) ? 4'b1010 : 4'b1011;
														assign node16091 = (inp[11]) ? node16099 : node16092;
															assign node16092 = (inp[10]) ? node16096 : node16093;
																assign node16093 = (inp[9]) ? 4'b1111 : 4'b1110;
																assign node16096 = (inp[9]) ? 4'b1110 : 4'b1111;
															assign node16099 = (inp[9]) ? node16103 : node16100;
																assign node16100 = (inp[10]) ? 4'b1110 : 4'b1111;
																assign node16103 = (inp[10]) ? 4'b1111 : 4'b1110;
													assign node16106 = (inp[15]) ? node16122 : node16107;
														assign node16107 = (inp[9]) ? node16115 : node16108;
															assign node16108 = (inp[11]) ? node16112 : node16109;
																assign node16109 = (inp[10]) ? 4'b1110 : 4'b1111;
																assign node16112 = (inp[10]) ? 4'b1111 : 4'b1110;
															assign node16115 = (inp[10]) ? node16119 : node16116;
																assign node16116 = (inp[11]) ? 4'b1111 : 4'b1110;
																assign node16119 = (inp[11]) ? 4'b1110 : 4'b1111;
														assign node16122 = (inp[9]) ? node16124 : 4'b1010;
															assign node16124 = (inp[11]) ? node16128 : node16125;
																assign node16125 = (inp[10]) ? 4'b1011 : 4'b1010;
																assign node16128 = (inp[10]) ? 4'b1010 : 4'b1011;
											assign node16131 = (inp[15]) ? node16169 : node16132;
												assign node16132 = (inp[9]) ? node16150 : node16133;
													assign node16133 = (inp[0]) ? node16145 : node16134;
														assign node16134 = (inp[10]) ? node16140 : node16135;
															assign node16135 = (inp[1]) ? 4'b1001 : node16136;
																assign node16136 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node16140 = (inp[11]) ? 4'b1000 : node16141;
																assign node16141 = (inp[1]) ? 4'b1000 : 4'b1001;
														assign node16145 = (inp[10]) ? node16147 : 4'b1000;
															assign node16147 = (inp[11]) ? 4'b1000 : 4'b1001;
													assign node16150 = (inp[0]) ? node16158 : node16151;
														assign node16151 = (inp[10]) ? node16153 : 4'b1000;
															assign node16153 = (inp[1]) ? 4'b1001 : node16154;
																assign node16154 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node16158 = (inp[10]) ? node16164 : node16159;
															assign node16159 = (inp[11]) ? node16161 : 4'b1001;
																assign node16161 = (inp[1]) ? 4'b1000 : 4'b1001;
															assign node16164 = (inp[11]) ? node16166 : 4'b1000;
																assign node16166 = (inp[1]) ? 4'b1001 : 4'b1000;
												assign node16169 = (inp[1]) ? node16185 : node16170;
													assign node16170 = (inp[11]) ? node16178 : node16171;
														assign node16171 = (inp[0]) ? 4'b1011 : node16172;
															assign node16172 = (inp[10]) ? 4'b1011 : node16173;
																assign node16173 = (inp[9]) ? 4'b1011 : 4'b1010;
														assign node16178 = (inp[9]) ? node16182 : node16179;
															assign node16179 = (inp[10]) ? 4'b1011 : 4'b1010;
															assign node16182 = (inp[10]) ? 4'b1010 : 4'b1011;
													assign node16185 = (inp[10]) ? node16195 : node16186;
														assign node16186 = (inp[9]) ? node16190 : node16187;
															assign node16187 = (inp[11]) ? 4'b1111 : 4'b1110;
															assign node16190 = (inp[0]) ? 4'b1111 : node16191;
																assign node16191 = (inp[11]) ? 4'b1110 : 4'b1111;
														assign node16195 = (inp[9]) ? 4'b1110 : node16196;
															assign node16196 = (inp[11]) ? node16198 : 4'b1111;
																assign node16198 = (inp[0]) ? 4'b1111 : 4'b1110;
										assign node16202 = (inp[4]) ? node16270 : node16203;
											assign node16203 = (inp[15]) ? node16241 : node16204;
												assign node16204 = (inp[10]) ? node16222 : node16205;
													assign node16205 = (inp[9]) ? node16217 : node16206;
														assign node16206 = (inp[1]) ? node16212 : node16207;
															assign node16207 = (inp[0]) ? 4'b1000 : node16208;
																assign node16208 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node16212 = (inp[11]) ? 4'b1000 : node16213;
																assign node16213 = (inp[0]) ? 4'b1001 : 4'b1000;
														assign node16217 = (inp[1]) ? node16219 : 4'b1001;
															assign node16219 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node16222 = (inp[9]) ? node16230 : node16223;
														assign node16223 = (inp[0]) ? 4'b1001 : node16224;
															assign node16224 = (inp[1]) ? 4'b1001 : node16225;
																assign node16225 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node16230 = (inp[0]) ? node16236 : node16231;
															assign node16231 = (inp[11]) ? node16233 : 4'b1000;
																assign node16233 = (inp[1]) ? 4'b1000 : 4'b1001;
															assign node16236 = (inp[11]) ? 4'b1000 : node16237;
																assign node16237 = (inp[1]) ? 4'b1001 : 4'b1000;
												assign node16241 = (inp[0]) ? node16263 : node16242;
													assign node16242 = (inp[9]) ? node16250 : node16243;
														assign node16243 = (inp[10]) ? node16247 : node16244;
															assign node16244 = (inp[11]) ? 4'b1100 : 4'b1101;
															assign node16247 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node16250 = (inp[1]) ? node16258 : node16251;
															assign node16251 = (inp[11]) ? node16255 : node16252;
																assign node16252 = (inp[10]) ? 4'b1101 : 4'b1100;
																assign node16255 = (inp[10]) ? 4'b1100 : 4'b1101;
															assign node16258 = (inp[10]) ? node16260 : 4'b1101;
																assign node16260 = (inp[11]) ? 4'b1100 : 4'b1101;
													assign node16263 = (inp[9]) ? node16267 : node16264;
														assign node16264 = (inp[10]) ? 4'b1100 : 4'b1101;
														assign node16267 = (inp[10]) ? 4'b1101 : 4'b1100;
											assign node16270 = (inp[15]) ? node16310 : node16271;
												assign node16271 = (inp[10]) ? node16291 : node16272;
													assign node16272 = (inp[1]) ? node16280 : node16273;
														assign node16273 = (inp[0]) ? node16275 : 4'b1111;
															assign node16275 = (inp[11]) ? 4'b1111 : node16276;
																assign node16276 = (inp[9]) ? 4'b1111 : 4'b1110;
														assign node16280 = (inp[9]) ? node16286 : node16281;
															assign node16281 = (inp[0]) ? 4'b1110 : node16282;
																assign node16282 = (inp[11]) ? 4'b1111 : 4'b1110;
															assign node16286 = (inp[11]) ? node16288 : 4'b1111;
																assign node16288 = (inp[0]) ? 4'b1111 : 4'b1110;
													assign node16291 = (inp[9]) ? node16303 : node16292;
														assign node16292 = (inp[1]) ? node16298 : node16293;
															assign node16293 = (inp[11]) ? 4'b1110 : node16294;
																assign node16294 = (inp[0]) ? 4'b1111 : 4'b1110;
															assign node16298 = (inp[0]) ? 4'b1111 : node16299;
																assign node16299 = (inp[11]) ? 4'b1110 : 4'b1111;
														assign node16303 = (inp[11]) ? node16305 : 4'b1110;
															assign node16305 = (inp[0]) ? node16307 : 4'b1111;
																assign node16307 = (inp[1]) ? 4'b1110 : 4'b1111;
												assign node16310 = (inp[9]) ? node16322 : node16311;
													assign node16311 = (inp[10]) ? node16317 : node16312;
														assign node16312 = (inp[0]) ? 4'b1100 : node16313;
															assign node16313 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node16317 = (inp[11]) ? node16319 : 4'b1101;
															assign node16319 = (inp[0]) ? 4'b1101 : 4'b1100;
													assign node16322 = (inp[10]) ? node16328 : node16323;
														assign node16323 = (inp[11]) ? node16325 : 4'b1101;
															assign node16325 = (inp[0]) ? 4'b1101 : 4'b1100;
														assign node16328 = (inp[0]) ? 4'b1100 : node16329;
															assign node16329 = (inp[11]) ? 4'b1101 : 4'b1100;
								assign node16333 = (inp[12]) ? node16683 : node16334;
									assign node16334 = (inp[7]) ? node16520 : node16335;
										assign node16335 = (inp[15]) ? node16431 : node16336;
											assign node16336 = (inp[4]) ? node16384 : node16337;
												assign node16337 = (inp[0]) ? node16361 : node16338;
													assign node16338 = (inp[1]) ? node16346 : node16339;
														assign node16339 = (inp[9]) ? node16343 : node16340;
															assign node16340 = (inp[10]) ? 4'b1000 : 4'b1001;
															assign node16343 = (inp[10]) ? 4'b1001 : 4'b1000;
														assign node16346 = (inp[10]) ? node16354 : node16347;
															assign node16347 = (inp[11]) ? node16351 : node16348;
																assign node16348 = (inp[9]) ? 4'b1000 : 4'b1001;
																assign node16351 = (inp[9]) ? 4'b1001 : 4'b1000;
															assign node16354 = (inp[11]) ? node16358 : node16355;
																assign node16355 = (inp[9]) ? 4'b1001 : 4'b1000;
																assign node16358 = (inp[9]) ? 4'b1000 : 4'b1001;
													assign node16361 = (inp[10]) ? node16373 : node16362;
														assign node16362 = (inp[9]) ? node16368 : node16363;
															assign node16363 = (inp[1]) ? 4'b1001 : node16364;
																assign node16364 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node16368 = (inp[11]) ? 4'b1000 : node16369;
																assign node16369 = (inp[1]) ? 4'b1000 : 4'b1001;
														assign node16373 = (inp[9]) ? node16379 : node16374;
															assign node16374 = (inp[1]) ? 4'b1000 : node16375;
																assign node16375 = (inp[11]) ? 4'b1000 : 4'b1001;
															assign node16379 = (inp[1]) ? 4'b1001 : node16380;
																assign node16380 = (inp[11]) ? 4'b1001 : 4'b1000;
												assign node16384 = (inp[11]) ? node16410 : node16385;
													assign node16385 = (inp[1]) ? node16401 : node16386;
														assign node16386 = (inp[0]) ? node16394 : node16387;
															assign node16387 = (inp[9]) ? node16391 : node16388;
																assign node16388 = (inp[10]) ? 4'b1011 : 4'b1010;
																assign node16391 = (inp[10]) ? 4'b1010 : 4'b1011;
															assign node16394 = (inp[10]) ? node16398 : node16395;
																assign node16395 = (inp[9]) ? 4'b1011 : 4'b1010;
																assign node16398 = (inp[9]) ? 4'b1010 : 4'b1011;
														assign node16401 = (inp[9]) ? 4'b1011 : node16402;
															assign node16402 = (inp[0]) ? node16406 : node16403;
																assign node16403 = (inp[10]) ? 4'b1010 : 4'b1011;
																assign node16406 = (inp[10]) ? 4'b1011 : 4'b1010;
													assign node16410 = (inp[10]) ? node16422 : node16411;
														assign node16411 = (inp[9]) ? node16417 : node16412;
															assign node16412 = (inp[0]) ? node16414 : 4'b1011;
																assign node16414 = (inp[1]) ? 4'b1011 : 4'b1010;
															assign node16417 = (inp[0]) ? node16419 : 4'b1010;
																assign node16419 = (inp[1]) ? 4'b1010 : 4'b1011;
														assign node16422 = (inp[9]) ? node16428 : node16423;
															assign node16423 = (inp[0]) ? node16425 : 4'b1010;
																assign node16425 = (inp[1]) ? 4'b1010 : 4'b1011;
															assign node16428 = (inp[1]) ? 4'b1011 : 4'b1010;
											assign node16431 = (inp[4]) ? node16473 : node16432;
												assign node16432 = (inp[10]) ? node16452 : node16433;
													assign node16433 = (inp[0]) ? node16439 : node16434;
														assign node16434 = (inp[1]) ? 4'b1000 : node16435;
															assign node16435 = (inp[9]) ? 4'b1001 : 4'b1000;
														assign node16439 = (inp[11]) ? node16447 : node16440;
															assign node16440 = (inp[9]) ? node16444 : node16441;
																assign node16441 = (inp[1]) ? 4'b1000 : 4'b1001;
																assign node16444 = (inp[1]) ? 4'b1001 : 4'b1000;
															assign node16447 = (inp[9]) ? 4'b1000 : node16448;
																assign node16448 = (inp[1]) ? 4'b1001 : 4'b1000;
													assign node16452 = (inp[1]) ? node16464 : node16453;
														assign node16453 = (inp[9]) ? node16459 : node16454;
															assign node16454 = (inp[0]) ? node16456 : 4'b1001;
																assign node16456 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node16459 = (inp[11]) ? 4'b1000 : node16460;
																assign node16460 = (inp[0]) ? 4'b1001 : 4'b1000;
														assign node16464 = (inp[9]) ? node16468 : node16465;
															assign node16465 = (inp[11]) ? 4'b1000 : 4'b1001;
															assign node16468 = (inp[11]) ? 4'b1001 : node16469;
																assign node16469 = (inp[0]) ? 4'b1000 : 4'b1001;
												assign node16473 = (inp[11]) ? node16495 : node16474;
													assign node16474 = (inp[10]) ? node16482 : node16475;
														assign node16475 = (inp[1]) ? node16479 : node16476;
															assign node16476 = (inp[9]) ? 4'b1100 : 4'b1101;
															assign node16479 = (inp[9]) ? 4'b1101 : 4'b1100;
														assign node16482 = (inp[0]) ? node16488 : node16483;
															assign node16483 = (inp[9]) ? node16485 : 4'b1101;
																assign node16485 = (inp[1]) ? 4'b1100 : 4'b1101;
															assign node16488 = (inp[1]) ? node16492 : node16489;
																assign node16489 = (inp[9]) ? 4'b1101 : 4'b1100;
																assign node16492 = (inp[9]) ? 4'b1100 : 4'b1101;
													assign node16495 = (inp[1]) ? node16505 : node16496;
														assign node16496 = (inp[0]) ? node16498 : 4'b1100;
															assign node16498 = (inp[9]) ? node16502 : node16499;
																assign node16499 = (inp[10]) ? 4'b1100 : 4'b1101;
																assign node16502 = (inp[10]) ? 4'b1101 : 4'b1100;
														assign node16505 = (inp[9]) ? node16513 : node16506;
															assign node16506 = (inp[0]) ? node16510 : node16507;
																assign node16507 = (inp[10]) ? 4'b1100 : 4'b1101;
																assign node16510 = (inp[10]) ? 4'b1101 : 4'b1100;
															assign node16513 = (inp[10]) ? node16517 : node16514;
																assign node16514 = (inp[0]) ? 4'b1101 : 4'b1100;
																assign node16517 = (inp[0]) ? 4'b1100 : 4'b1101;
										assign node16520 = (inp[4]) ? node16600 : node16521;
											assign node16521 = (inp[10]) ? node16559 : node16522;
												assign node16522 = (inp[9]) ? node16542 : node16523;
													assign node16523 = (inp[15]) ? node16533 : node16524;
														assign node16524 = (inp[1]) ? node16528 : node16525;
															assign node16525 = (inp[0]) ? 4'b1111 : 4'b1110;
															assign node16528 = (inp[0]) ? 4'b1010 : node16529;
																assign node16529 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node16533 = (inp[1]) ? node16539 : node16534;
															assign node16534 = (inp[0]) ? 4'b1011 : node16535;
																assign node16535 = (inp[11]) ? 4'b1010 : 4'b1011;
															assign node16539 = (inp[11]) ? 4'b1110 : 4'b1111;
													assign node16542 = (inp[1]) ? node16552 : node16543;
														assign node16543 = (inp[15]) ? node16547 : node16544;
															assign node16544 = (inp[0]) ? 4'b1110 : 4'b1111;
															assign node16547 = (inp[11]) ? node16549 : 4'b1010;
																assign node16549 = (inp[0]) ? 4'b1010 : 4'b1011;
														assign node16552 = (inp[15]) ? node16554 : 4'b1011;
															assign node16554 = (inp[0]) ? node16556 : 4'b1111;
																assign node16556 = (inp[11]) ? 4'b1111 : 4'b1110;
												assign node16559 = (inp[9]) ? node16583 : node16560;
													assign node16560 = (inp[11]) ? node16572 : node16561;
														assign node16561 = (inp[1]) ? node16567 : node16562;
															assign node16562 = (inp[15]) ? 4'b1010 : node16563;
																assign node16563 = (inp[0]) ? 4'b1110 : 4'b1111;
															assign node16567 = (inp[15]) ? node16569 : 4'b1011;
																assign node16569 = (inp[0]) ? 4'b1110 : 4'b1111;
														assign node16572 = (inp[15]) ? node16578 : node16573;
															assign node16573 = (inp[1]) ? node16575 : 4'b1111;
																assign node16575 = (inp[0]) ? 4'b1011 : 4'b1010;
															assign node16578 = (inp[1]) ? 4'b1111 : node16579;
																assign node16579 = (inp[0]) ? 4'b1010 : 4'b1011;
													assign node16583 = (inp[1]) ? node16593 : node16584;
														assign node16584 = (inp[15]) ? node16590 : node16585;
															assign node16585 = (inp[11]) ? 4'b1110 : node16586;
																assign node16586 = (inp[0]) ? 4'b1111 : 4'b1110;
															assign node16590 = (inp[11]) ? 4'b1010 : 4'b1011;
														assign node16593 = (inp[15]) ? 4'b1110 : node16594;
															assign node16594 = (inp[0]) ? 4'b1010 : node16595;
																assign node16595 = (inp[11]) ? 4'b1011 : 4'b1010;
											assign node16600 = (inp[15]) ? node16640 : node16601;
												assign node16601 = (inp[9]) ? node16621 : node16602;
													assign node16602 = (inp[10]) ? node16610 : node16603;
														assign node16603 = (inp[11]) ? 4'b1100 : node16604;
															assign node16604 = (inp[0]) ? 4'b1101 : node16605;
																assign node16605 = (inp[1]) ? 4'b1100 : 4'b1101;
														assign node16610 = (inp[11]) ? node16616 : node16611;
															assign node16611 = (inp[1]) ? node16613 : 4'b1100;
																assign node16613 = (inp[0]) ? 4'b1100 : 4'b1101;
															assign node16616 = (inp[1]) ? 4'b1101 : node16617;
																assign node16617 = (inp[0]) ? 4'b1100 : 4'b1101;
													assign node16621 = (inp[10]) ? node16629 : node16622;
														assign node16622 = (inp[1]) ? 4'b1101 : node16623;
															assign node16623 = (inp[11]) ? node16625 : 4'b1100;
																assign node16625 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node16629 = (inp[11]) ? node16635 : node16630;
															assign node16630 = (inp[0]) ? 4'b1101 : node16631;
																assign node16631 = (inp[1]) ? 4'b1100 : 4'b1101;
															assign node16635 = (inp[0]) ? node16637 : 4'b1100;
																assign node16637 = (inp[1]) ? 4'b1100 : 4'b1101;
												assign node16640 = (inp[1]) ? node16658 : node16641;
													assign node16641 = (inp[9]) ? node16651 : node16642;
														assign node16642 = (inp[10]) ? node16648 : node16643;
															assign node16643 = (inp[11]) ? 4'b1111 : node16644;
																assign node16644 = (inp[0]) ? 4'b1110 : 4'b1111;
															assign node16648 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node16651 = (inp[10]) ? node16653 : 4'b1110;
															assign node16653 = (inp[11]) ? 4'b1111 : node16654;
																assign node16654 = (inp[0]) ? 4'b1110 : 4'b1111;
													assign node16658 = (inp[11]) ? node16674 : node16659;
														assign node16659 = (inp[0]) ? node16667 : node16660;
															assign node16660 = (inp[9]) ? node16664 : node16661;
																assign node16661 = (inp[10]) ? 4'b1011 : 4'b1010;
																assign node16664 = (inp[10]) ? 4'b1010 : 4'b1011;
															assign node16667 = (inp[10]) ? node16671 : node16668;
																assign node16668 = (inp[9]) ? 4'b1010 : 4'b1011;
																assign node16671 = (inp[9]) ? 4'b1011 : 4'b1010;
														assign node16674 = (inp[0]) ? node16676 : 4'b1011;
															assign node16676 = (inp[9]) ? node16680 : node16677;
																assign node16677 = (inp[10]) ? 4'b1011 : 4'b1010;
																assign node16680 = (inp[10]) ? 4'b1010 : 4'b1011;
									assign node16683 = (inp[7]) ? node16849 : node16684;
										assign node16684 = (inp[4]) ? node16778 : node16685;
											assign node16685 = (inp[11]) ? node16733 : node16686;
												assign node16686 = (inp[1]) ? node16716 : node16687;
													assign node16687 = (inp[0]) ? node16701 : node16688;
														assign node16688 = (inp[10]) ? node16696 : node16689;
															assign node16689 = (inp[15]) ? node16693 : node16690;
																assign node16690 = (inp[9]) ? 4'b1010 : 4'b1011;
																assign node16693 = (inp[9]) ? 4'b1011 : 4'b1010;
															assign node16696 = (inp[15]) ? 4'b1010 : node16697;
																assign node16697 = (inp[9]) ? 4'b1011 : 4'b1010;
														assign node16701 = (inp[15]) ? node16709 : node16702;
															assign node16702 = (inp[10]) ? node16706 : node16703;
																assign node16703 = (inp[9]) ? 4'b1011 : 4'b1010;
																assign node16706 = (inp[9]) ? 4'b1010 : 4'b1011;
															assign node16709 = (inp[9]) ? node16713 : node16710;
																assign node16710 = (inp[10]) ? 4'b1010 : 4'b1011;
																assign node16713 = (inp[10]) ? 4'b1011 : 4'b1010;
													assign node16716 = (inp[10]) ? node16728 : node16717;
														assign node16717 = (inp[9]) ? node16723 : node16718;
															assign node16718 = (inp[0]) ? node16720 : 4'b1010;
																assign node16720 = (inp[15]) ? 4'b1011 : 4'b1010;
															assign node16723 = (inp[15]) ? node16725 : 4'b1011;
																assign node16725 = (inp[0]) ? 4'b1010 : 4'b1011;
														assign node16728 = (inp[9]) ? node16730 : 4'b1011;
															assign node16730 = (inp[15]) ? 4'b1011 : 4'b1010;
												assign node16733 = (inp[15]) ? node16763 : node16734;
													assign node16734 = (inp[1]) ? node16750 : node16735;
														assign node16735 = (inp[0]) ? node16743 : node16736;
															assign node16736 = (inp[10]) ? node16740 : node16737;
																assign node16737 = (inp[9]) ? 4'b1010 : 4'b1011;
																assign node16740 = (inp[9]) ? 4'b1011 : 4'b1010;
															assign node16743 = (inp[10]) ? node16747 : node16744;
																assign node16744 = (inp[9]) ? 4'b1010 : 4'b1011;
																assign node16747 = (inp[9]) ? 4'b1011 : 4'b1010;
														assign node16750 = (inp[0]) ? node16756 : node16751;
															assign node16751 = (inp[10]) ? 4'b1010 : node16752;
																assign node16752 = (inp[9]) ? 4'b1010 : 4'b1011;
															assign node16756 = (inp[9]) ? node16760 : node16757;
																assign node16757 = (inp[10]) ? 4'b1011 : 4'b1010;
																assign node16760 = (inp[10]) ? 4'b1010 : 4'b1011;
													assign node16763 = (inp[1]) ? node16771 : node16764;
														assign node16764 = (inp[10]) ? node16768 : node16765;
															assign node16765 = (inp[9]) ? 4'b1011 : 4'b1010;
															assign node16768 = (inp[9]) ? 4'b1010 : 4'b1011;
														assign node16771 = (inp[10]) ? node16775 : node16772;
															assign node16772 = (inp[9]) ? 4'b1011 : 4'b1010;
															assign node16775 = (inp[9]) ? 4'b1010 : 4'b1011;
											assign node16778 = (inp[15]) ? node16826 : node16779;
												assign node16779 = (inp[1]) ? node16801 : node16780;
													assign node16780 = (inp[9]) ? node16792 : node16781;
														assign node16781 = (inp[10]) ? node16787 : node16782;
															assign node16782 = (inp[0]) ? node16784 : 4'b1001;
																assign node16784 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node16787 = (inp[0]) ? node16789 : 4'b1000;
																assign node16789 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node16792 = (inp[10]) ? node16796 : node16793;
															assign node16793 = (inp[0]) ? 4'b1001 : 4'b1000;
															assign node16796 = (inp[0]) ? node16798 : 4'b1001;
																assign node16798 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node16801 = (inp[0]) ? node16817 : node16802;
														assign node16802 = (inp[11]) ? node16810 : node16803;
															assign node16803 = (inp[10]) ? node16807 : node16804;
																assign node16804 = (inp[9]) ? 4'b1101 : 4'b1100;
																assign node16807 = (inp[9]) ? 4'b1100 : 4'b1101;
															assign node16810 = (inp[10]) ? node16814 : node16811;
																assign node16811 = (inp[9]) ? 4'b1101 : 4'b1100;
																assign node16814 = (inp[9]) ? 4'b1100 : 4'b1101;
														assign node16817 = (inp[9]) ? node16819 : 4'b1100;
															assign node16819 = (inp[11]) ? node16823 : node16820;
																assign node16820 = (inp[10]) ? 4'b1101 : 4'b1100;
																assign node16823 = (inp[10]) ? 4'b1100 : 4'b1101;
												assign node16826 = (inp[10]) ? node16838 : node16827;
													assign node16827 = (inp[9]) ? node16833 : node16828;
														assign node16828 = (inp[0]) ? node16830 : 4'b1010;
															assign node16830 = (inp[11]) ? 4'b1010 : 4'b1011;
														assign node16833 = (inp[0]) ? node16835 : 4'b1011;
															assign node16835 = (inp[11]) ? 4'b1011 : 4'b1010;
													assign node16838 = (inp[9]) ? node16844 : node16839;
														assign node16839 = (inp[0]) ? node16841 : 4'b1011;
															assign node16841 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node16844 = (inp[11]) ? 4'b1010 : node16845;
															assign node16845 = (inp[0]) ? 4'b1011 : 4'b1010;
										assign node16849 = (inp[15]) ? node16941 : node16850;
											assign node16850 = (inp[4]) ? node16890 : node16851;
												assign node16851 = (inp[9]) ? node16873 : node16852;
													assign node16852 = (inp[10]) ? node16864 : node16853;
														assign node16853 = (inp[11]) ? node16859 : node16854;
															assign node16854 = (inp[0]) ? node16856 : 4'b1100;
																assign node16856 = (inp[1]) ? 4'b1101 : 4'b1100;
															assign node16859 = (inp[0]) ? 4'b1100 : node16860;
																assign node16860 = (inp[1]) ? 4'b1100 : 4'b1101;
														assign node16864 = (inp[0]) ? node16868 : node16865;
															assign node16865 = (inp[11]) ? 4'b1100 : 4'b1101;
															assign node16868 = (inp[11]) ? 4'b1101 : node16869;
																assign node16869 = (inp[1]) ? 4'b1100 : 4'b1101;
													assign node16873 = (inp[10]) ? node16881 : node16874;
														assign node16874 = (inp[0]) ? node16876 : 4'b1101;
															assign node16876 = (inp[11]) ? 4'b1101 : node16877;
																assign node16877 = (inp[1]) ? 4'b1100 : 4'b1101;
														assign node16881 = (inp[11]) ? node16885 : node16882;
															assign node16882 = (inp[1]) ? 4'b1101 : 4'b1100;
															assign node16885 = (inp[0]) ? 4'b1100 : node16886;
																assign node16886 = (inp[1]) ? 4'b1100 : 4'b1101;
												assign node16890 = (inp[11]) ? node16918 : node16891;
													assign node16891 = (inp[0]) ? node16905 : node16892;
														assign node16892 = (inp[1]) ? node16900 : node16893;
															assign node16893 = (inp[9]) ? node16897 : node16894;
																assign node16894 = (inp[10]) ? 4'b1011 : 4'b1010;
																assign node16897 = (inp[10]) ? 4'b1010 : 4'b1011;
															assign node16900 = (inp[10]) ? node16902 : 4'b1011;
																assign node16902 = (inp[9]) ? 4'b1010 : 4'b1011;
														assign node16905 = (inp[10]) ? node16913 : node16906;
															assign node16906 = (inp[9]) ? node16910 : node16907;
																assign node16907 = (inp[1]) ? 4'b1011 : 4'b1010;
																assign node16910 = (inp[1]) ? 4'b1010 : 4'b1011;
															assign node16913 = (inp[1]) ? node16915 : 4'b1011;
																assign node16915 = (inp[9]) ? 4'b1011 : 4'b1010;
													assign node16918 = (inp[9]) ? node16930 : node16919;
														assign node16919 = (inp[10]) ? node16925 : node16920;
															assign node16920 = (inp[1]) ? 4'b1010 : node16921;
																assign node16921 = (inp[0]) ? 4'b1010 : 4'b1011;
															assign node16925 = (inp[1]) ? 4'b1011 : node16926;
																assign node16926 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node16930 = (inp[10]) ? node16936 : node16931;
															assign node16931 = (inp[1]) ? 4'b1011 : node16932;
																assign node16932 = (inp[0]) ? 4'b1011 : 4'b1010;
															assign node16936 = (inp[0]) ? 4'b1010 : node16937;
																assign node16937 = (inp[1]) ? 4'b1010 : 4'b1011;
											assign node16941 = (inp[11]) ? node16973 : node16942;
												assign node16942 = (inp[10]) ? node16958 : node16943;
													assign node16943 = (inp[4]) ? node16951 : node16944;
														assign node16944 = (inp[9]) ? node16948 : node16945;
															assign node16945 = (inp[0]) ? 4'b1001 : 4'b1000;
															assign node16948 = (inp[0]) ? 4'b1000 : 4'b1001;
														assign node16951 = (inp[0]) ? node16955 : node16952;
															assign node16952 = (inp[9]) ? 4'b1001 : 4'b1000;
															assign node16955 = (inp[9]) ? 4'b1000 : 4'b1001;
													assign node16958 = (inp[1]) ? node16966 : node16959;
														assign node16959 = (inp[0]) ? node16963 : node16960;
															assign node16960 = (inp[9]) ? 4'b1000 : 4'b1001;
															assign node16963 = (inp[9]) ? 4'b1001 : 4'b1000;
														assign node16966 = (inp[9]) ? node16970 : node16967;
															assign node16967 = (inp[0]) ? 4'b1000 : 4'b1001;
															assign node16970 = (inp[0]) ? 4'b1001 : 4'b1000;
												assign node16973 = (inp[1]) ? node16981 : node16974;
													assign node16974 = (inp[9]) ? node16978 : node16975;
														assign node16975 = (inp[10]) ? 4'b1001 : 4'b1000;
														assign node16978 = (inp[10]) ? 4'b1000 : 4'b1001;
													assign node16981 = (inp[4]) ? node16997 : node16982;
														assign node16982 = (inp[0]) ? node16990 : node16983;
															assign node16983 = (inp[10]) ? node16987 : node16984;
																assign node16984 = (inp[9]) ? 4'b1001 : 4'b1000;
																assign node16987 = (inp[9]) ? 4'b1000 : 4'b1001;
															assign node16990 = (inp[9]) ? node16994 : node16991;
																assign node16991 = (inp[10]) ? 4'b1001 : 4'b1000;
																assign node16994 = (inp[10]) ? 4'b1000 : 4'b1001;
														assign node16997 = (inp[9]) ? node17001 : node16998;
															assign node16998 = (inp[10]) ? 4'b1001 : 4'b1000;
															assign node17001 = (inp[10]) ? 4'b1000 : 4'b1001;
							assign node17004 = (inp[12]) ? node17576 : node17005;
								assign node17005 = (inp[15]) ? node17281 : node17006;
									assign node17006 = (inp[7]) ? node17164 : node17007;
										assign node17007 = (inp[4]) ? node17099 : node17008;
											assign node17008 = (inp[1]) ? node17052 : node17009;
												assign node17009 = (inp[2]) ? node17039 : node17010;
													assign node17010 = (inp[10]) ? node17024 : node17011;
														assign node17011 = (inp[0]) ? node17017 : node17012;
															assign node17012 = (inp[11]) ? 4'b1001 : node17013;
																assign node17013 = (inp[9]) ? 4'b1000 : 4'b1001;
															assign node17017 = (inp[9]) ? node17021 : node17018;
																assign node17018 = (inp[11]) ? 4'b1001 : 4'b1000;
																assign node17021 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node17024 = (inp[0]) ? node17032 : node17025;
															assign node17025 = (inp[11]) ? node17029 : node17026;
																assign node17026 = (inp[9]) ? 4'b1000 : 4'b1001;
																assign node17029 = (inp[9]) ? 4'b1001 : 4'b1000;
															assign node17032 = (inp[9]) ? node17036 : node17033;
																assign node17033 = (inp[11]) ? 4'b1001 : 4'b1000;
																assign node17036 = (inp[11]) ? 4'b1000 : 4'b1001;
													assign node17039 = (inp[10]) ? node17047 : node17040;
														assign node17040 = (inp[11]) ? node17044 : node17041;
															assign node17041 = (inp[9]) ? 4'b1000 : 4'b1001;
															assign node17044 = (inp[9]) ? 4'b1001 : 4'b1000;
														assign node17047 = (inp[11]) ? node17049 : 4'b1000;
															assign node17049 = (inp[9]) ? 4'b1001 : 4'b1000;
												assign node17052 = (inp[10]) ? node17074 : node17053;
													assign node17053 = (inp[9]) ? node17063 : node17054;
														assign node17054 = (inp[11]) ? node17060 : node17055;
															assign node17055 = (inp[2]) ? 4'b1101 : node17056;
																assign node17056 = (inp[0]) ? 4'b1100 : 4'b1101;
															assign node17060 = (inp[2]) ? 4'b1100 : 4'b1101;
														assign node17063 = (inp[11]) ? node17069 : node17064;
															assign node17064 = (inp[2]) ? 4'b1100 : node17065;
																assign node17065 = (inp[0]) ? 4'b1101 : 4'b1100;
															assign node17069 = (inp[0]) ? node17071 : 4'b1101;
																assign node17071 = (inp[2]) ? 4'b1101 : 4'b1100;
													assign node17074 = (inp[0]) ? node17090 : node17075;
														assign node17075 = (inp[2]) ? node17083 : node17076;
															assign node17076 = (inp[11]) ? node17080 : node17077;
																assign node17077 = (inp[9]) ? 4'b1100 : 4'b1101;
																assign node17080 = (inp[9]) ? 4'b1101 : 4'b1100;
															assign node17083 = (inp[9]) ? node17087 : node17084;
																assign node17084 = (inp[11]) ? 4'b1100 : 4'b1101;
																assign node17087 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node17090 = (inp[2]) ? 4'b1100 : node17091;
															assign node17091 = (inp[9]) ? node17095 : node17092;
																assign node17092 = (inp[11]) ? 4'b1101 : 4'b1100;
																assign node17095 = (inp[11]) ? 4'b1100 : 4'b1101;
											assign node17099 = (inp[0]) ? node17123 : node17100;
												assign node17100 = (inp[9]) ? node17112 : node17101;
													assign node17101 = (inp[11]) ? node17107 : node17102;
														assign node17102 = (inp[1]) ? node17104 : 4'b1001;
															assign node17104 = (inp[2]) ? 4'b1001 : 4'b1000;
														assign node17107 = (inp[2]) ? 4'b1000 : node17108;
															assign node17108 = (inp[1]) ? 4'b1001 : 4'b1000;
													assign node17112 = (inp[11]) ? node17118 : node17113;
														assign node17113 = (inp[2]) ? 4'b1000 : node17114;
															assign node17114 = (inp[1]) ? 4'b1001 : 4'b1000;
														assign node17118 = (inp[2]) ? 4'b1001 : node17119;
															assign node17119 = (inp[1]) ? 4'b1000 : 4'b1001;
												assign node17123 = (inp[1]) ? node17141 : node17124;
													assign node17124 = (inp[11]) ? node17132 : node17125;
														assign node17125 = (inp[2]) ? node17129 : node17126;
															assign node17126 = (inp[9]) ? 4'b1000 : 4'b1001;
															assign node17129 = (inp[9]) ? 4'b1001 : 4'b1000;
														assign node17132 = (inp[10]) ? 4'b1001 : node17133;
															assign node17133 = (inp[9]) ? node17137 : node17134;
																assign node17134 = (inp[2]) ? 4'b1001 : 4'b1000;
																assign node17137 = (inp[2]) ? 4'b1000 : 4'b1001;
													assign node17141 = (inp[10]) ? node17149 : node17142;
														assign node17142 = (inp[9]) ? node17146 : node17143;
															assign node17143 = (inp[11]) ? 4'b1000 : 4'b1001;
															assign node17146 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node17149 = (inp[2]) ? node17157 : node17150;
															assign node17150 = (inp[11]) ? node17154 : node17151;
																assign node17151 = (inp[9]) ? 4'b1000 : 4'b1001;
																assign node17154 = (inp[9]) ? 4'b1001 : 4'b1000;
															assign node17157 = (inp[11]) ? node17161 : node17158;
																assign node17158 = (inp[9]) ? 4'b1000 : 4'b1001;
																assign node17161 = (inp[9]) ? 4'b1001 : 4'b1000;
										assign node17164 = (inp[4]) ? node17214 : node17165;
											assign node17165 = (inp[2]) ? node17191 : node17166;
												assign node17166 = (inp[0]) ? node17174 : node17167;
													assign node17167 = (inp[9]) ? node17171 : node17168;
														assign node17168 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node17171 = (inp[11]) ? 4'b1010 : 4'b1011;
													assign node17174 = (inp[11]) ? node17182 : node17175;
														assign node17175 = (inp[9]) ? node17179 : node17176;
															assign node17176 = (inp[1]) ? 4'b1010 : 4'b1011;
															assign node17179 = (inp[1]) ? 4'b1011 : 4'b1010;
														assign node17182 = (inp[10]) ? node17184 : 4'b1011;
															assign node17184 = (inp[9]) ? node17188 : node17185;
																assign node17185 = (inp[1]) ? 4'b1011 : 4'b1010;
																assign node17188 = (inp[1]) ? 4'b1010 : 4'b1011;
												assign node17191 = (inp[11]) ? node17203 : node17192;
													assign node17192 = (inp[9]) ? node17198 : node17193;
														assign node17193 = (inp[1]) ? node17195 : 4'b1010;
															assign node17195 = (inp[0]) ? 4'b1010 : 4'b1011;
														assign node17198 = (inp[0]) ? 4'b1011 : node17199;
															assign node17199 = (inp[1]) ? 4'b1010 : 4'b1011;
													assign node17203 = (inp[9]) ? node17209 : node17204;
														assign node17204 = (inp[0]) ? 4'b1011 : node17205;
															assign node17205 = (inp[1]) ? 4'b1010 : 4'b1011;
														assign node17209 = (inp[1]) ? node17211 : 4'b1010;
															assign node17211 = (inp[0]) ? 4'b1010 : 4'b1011;
											assign node17214 = (inp[1]) ? node17258 : node17215;
												assign node17215 = (inp[0]) ? node17237 : node17216;
													assign node17216 = (inp[2]) ? node17230 : node17217;
														assign node17217 = (inp[10]) ? node17225 : node17218;
															assign node17218 = (inp[9]) ? node17222 : node17219;
																assign node17219 = (inp[11]) ? 4'b1111 : 4'b1110;
																assign node17222 = (inp[11]) ? 4'b1110 : 4'b1111;
															assign node17225 = (inp[9]) ? 4'b1110 : node17226;
																assign node17226 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node17230 = (inp[9]) ? node17234 : node17231;
															assign node17231 = (inp[11]) ? 4'b1111 : 4'b1110;
															assign node17234 = (inp[11]) ? 4'b1110 : 4'b1111;
													assign node17237 = (inp[10]) ? node17245 : node17238;
														assign node17238 = (inp[11]) ? 4'b1110 : node17239;
															assign node17239 = (inp[2]) ? node17241 : 4'b1110;
																assign node17241 = (inp[9]) ? 4'b1110 : 4'b1111;
														assign node17245 = (inp[9]) ? node17251 : node17246;
															assign node17246 = (inp[2]) ? 4'b1110 : node17247;
																assign node17247 = (inp[11]) ? 4'b1111 : 4'b1110;
															assign node17251 = (inp[2]) ? node17255 : node17252;
																assign node17252 = (inp[11]) ? 4'b1110 : 4'b1111;
																assign node17255 = (inp[11]) ? 4'b1111 : 4'b1110;
												assign node17258 = (inp[11]) ? node17270 : node17259;
													assign node17259 = (inp[9]) ? node17265 : node17260;
														assign node17260 = (inp[2]) ? 4'b1010 : node17261;
															assign node17261 = (inp[0]) ? 4'b1010 : 4'b1011;
														assign node17265 = (inp[2]) ? 4'b1011 : node17266;
															assign node17266 = (inp[0]) ? 4'b1011 : 4'b1010;
													assign node17270 = (inp[9]) ? node17276 : node17271;
														assign node17271 = (inp[2]) ? 4'b1011 : node17272;
															assign node17272 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node17276 = (inp[2]) ? 4'b1010 : node17277;
															assign node17277 = (inp[0]) ? 4'b1010 : 4'b1011;
									assign node17281 = (inp[7]) ? node17437 : node17282;
										assign node17282 = (inp[2]) ? node17378 : node17283;
											assign node17283 = (inp[10]) ? node17327 : node17284;
												assign node17284 = (inp[1]) ? node17312 : node17285;
													assign node17285 = (inp[4]) ? node17299 : node17286;
														assign node17286 = (inp[9]) ? node17292 : node17287;
															assign node17287 = (inp[11]) ? node17289 : 4'b1011;
																assign node17289 = (inp[0]) ? 4'b1010 : 4'b1011;
															assign node17292 = (inp[0]) ? node17296 : node17293;
																assign node17293 = (inp[11]) ? 4'b1010 : 4'b1011;
																assign node17296 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node17299 = (inp[0]) ? node17305 : node17300;
															assign node17300 = (inp[11]) ? node17302 : 4'b1111;
																assign node17302 = (inp[9]) ? 4'b1110 : 4'b1111;
															assign node17305 = (inp[11]) ? node17309 : node17306;
																assign node17306 = (inp[9]) ? 4'b1111 : 4'b1110;
																assign node17309 = (inp[9]) ? 4'b1110 : 4'b1111;
													assign node17312 = (inp[4]) ? node17320 : node17313;
														assign node17313 = (inp[9]) ? node17317 : node17314;
															assign node17314 = (inp[11]) ? 4'b1111 : 4'b1110;
															assign node17317 = (inp[11]) ? 4'b1110 : 4'b1111;
														assign node17320 = (inp[9]) ? node17324 : node17321;
															assign node17321 = (inp[11]) ? 4'b1010 : 4'b1011;
															assign node17324 = (inp[11]) ? 4'b1011 : 4'b1010;
												assign node17327 = (inp[0]) ? node17355 : node17328;
													assign node17328 = (inp[9]) ? node17344 : node17329;
														assign node17329 = (inp[11]) ? node17337 : node17330;
															assign node17330 = (inp[1]) ? node17334 : node17331;
																assign node17331 = (inp[4]) ? 4'b1110 : 4'b1010;
																assign node17334 = (inp[4]) ? 4'b1011 : 4'b1110;
															assign node17337 = (inp[4]) ? node17341 : node17338;
																assign node17338 = (inp[1]) ? 4'b1111 : 4'b1011;
																assign node17341 = (inp[1]) ? 4'b1010 : 4'b1111;
														assign node17344 = (inp[11]) ? node17350 : node17345;
															assign node17345 = (inp[1]) ? 4'b1010 : node17346;
																assign node17346 = (inp[4]) ? 4'b1111 : 4'b1011;
															assign node17350 = (inp[4]) ? 4'b1011 : node17351;
																assign node17351 = (inp[1]) ? 4'b1110 : 4'b1010;
													assign node17355 = (inp[11]) ? node17363 : node17356;
														assign node17356 = (inp[9]) ? 4'b1111 : node17357;
															assign node17357 = (inp[1]) ? 4'b1011 : node17358;
																assign node17358 = (inp[4]) ? 4'b1110 : 4'b1011;
														assign node17363 = (inp[1]) ? node17371 : node17364;
															assign node17364 = (inp[4]) ? node17368 : node17365;
																assign node17365 = (inp[9]) ? 4'b1011 : 4'b1010;
																assign node17368 = (inp[9]) ? 4'b1110 : 4'b1111;
															assign node17371 = (inp[4]) ? node17375 : node17372;
																assign node17372 = (inp[9]) ? 4'b1110 : 4'b1111;
																assign node17375 = (inp[9]) ? 4'b1011 : 4'b1010;
											assign node17378 = (inp[9]) ? node17408 : node17379;
												assign node17379 = (inp[11]) ? node17393 : node17380;
													assign node17380 = (inp[1]) ? node17386 : node17381;
														assign node17381 = (inp[4]) ? node17383 : 4'b1010;
															assign node17383 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node17386 = (inp[4]) ? node17390 : node17387;
															assign node17387 = (inp[0]) ? 4'b1110 : 4'b1111;
															assign node17390 = (inp[0]) ? 4'b1010 : 4'b1011;
													assign node17393 = (inp[0]) ? node17401 : node17394;
														assign node17394 = (inp[1]) ? node17398 : node17395;
															assign node17395 = (inp[4]) ? 4'b1111 : 4'b1011;
															assign node17398 = (inp[4]) ? 4'b1010 : 4'b1110;
														assign node17401 = (inp[1]) ? node17405 : node17402;
															assign node17402 = (inp[4]) ? 4'b1110 : 4'b1011;
															assign node17405 = (inp[4]) ? 4'b1011 : 4'b1111;
												assign node17408 = (inp[11]) ? node17424 : node17409;
													assign node17409 = (inp[0]) ? node17417 : node17410;
														assign node17410 = (inp[1]) ? node17414 : node17411;
															assign node17411 = (inp[4]) ? 4'b1111 : 4'b1011;
															assign node17414 = (inp[4]) ? 4'b1010 : 4'b1110;
														assign node17417 = (inp[1]) ? node17421 : node17418;
															assign node17418 = (inp[4]) ? 4'b1110 : 4'b1011;
															assign node17421 = (inp[4]) ? 4'b1011 : 4'b1111;
													assign node17424 = (inp[1]) ? node17430 : node17425;
														assign node17425 = (inp[4]) ? node17427 : 4'b1010;
															assign node17427 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node17430 = (inp[0]) ? node17434 : node17431;
															assign node17431 = (inp[4]) ? 4'b1011 : 4'b1111;
															assign node17434 = (inp[4]) ? 4'b1010 : 4'b1110;
										assign node17437 = (inp[1]) ? node17515 : node17438;
											assign node17438 = (inp[4]) ? node17472 : node17439;
												assign node17439 = (inp[2]) ? node17457 : node17440;
													assign node17440 = (inp[0]) ? node17450 : node17441;
														assign node17441 = (inp[10]) ? 4'b1001 : node17442;
															assign node17442 = (inp[11]) ? node17446 : node17443;
																assign node17443 = (inp[9]) ? 4'b1000 : 4'b1001;
																assign node17446 = (inp[9]) ? 4'b1001 : 4'b1000;
														assign node17450 = (inp[11]) ? node17454 : node17451;
															assign node17451 = (inp[9]) ? 4'b1000 : 4'b1001;
															assign node17454 = (inp[9]) ? 4'b1001 : 4'b1000;
													assign node17457 = (inp[11]) ? node17465 : node17458;
														assign node17458 = (inp[0]) ? node17462 : node17459;
															assign node17459 = (inp[9]) ? 4'b1001 : 4'b1000;
															assign node17462 = (inp[9]) ? 4'b1000 : 4'b1001;
														assign node17465 = (inp[9]) ? node17469 : node17466;
															assign node17466 = (inp[0]) ? 4'b1000 : 4'b1001;
															assign node17469 = (inp[0]) ? 4'b1001 : 4'b1000;
												assign node17472 = (inp[0]) ? node17502 : node17473;
													assign node17473 = (inp[2]) ? node17487 : node17474;
														assign node17474 = (inp[10]) ? node17480 : node17475;
															assign node17475 = (inp[11]) ? 4'b1101 : node17476;
																assign node17476 = (inp[9]) ? 4'b1101 : 4'b1100;
															assign node17480 = (inp[11]) ? node17484 : node17481;
																assign node17481 = (inp[9]) ? 4'b1101 : 4'b1100;
																assign node17484 = (inp[9]) ? 4'b1100 : 4'b1101;
														assign node17487 = (inp[10]) ? node17495 : node17488;
															assign node17488 = (inp[9]) ? node17492 : node17489;
																assign node17489 = (inp[11]) ? 4'b1100 : 4'b1101;
																assign node17492 = (inp[11]) ? 4'b1101 : 4'b1100;
															assign node17495 = (inp[9]) ? node17499 : node17496;
																assign node17496 = (inp[11]) ? 4'b1100 : 4'b1101;
																assign node17499 = (inp[11]) ? 4'b1101 : 4'b1100;
													assign node17502 = (inp[10]) ? node17510 : node17503;
														assign node17503 = (inp[11]) ? node17507 : node17504;
															assign node17504 = (inp[9]) ? 4'b1100 : 4'b1101;
															assign node17507 = (inp[9]) ? 4'b1101 : 4'b1100;
														assign node17510 = (inp[11]) ? node17512 : 4'b1101;
															assign node17512 = (inp[9]) ? 4'b1101 : 4'b1100;
											assign node17515 = (inp[4]) ? node17535 : node17516;
												assign node17516 = (inp[11]) ? node17526 : node17517;
													assign node17517 = (inp[9]) ? node17523 : node17518;
														assign node17518 = (inp[0]) ? node17520 : 4'b1100;
															assign node17520 = (inp[2]) ? 4'b1100 : 4'b1101;
														assign node17523 = (inp[2]) ? 4'b1101 : 4'b1100;
													assign node17526 = (inp[9]) ? node17532 : node17527;
														assign node17527 = (inp[2]) ? 4'b1101 : node17528;
															assign node17528 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node17532 = (inp[0]) ? 4'b1101 : 4'b1100;
												assign node17535 = (inp[10]) ? node17555 : node17536;
													assign node17536 = (inp[11]) ? node17544 : node17537;
														assign node17537 = (inp[9]) ? 4'b1001 : node17538;
															assign node17538 = (inp[0]) ? 4'b1000 : node17539;
																assign node17539 = (inp[2]) ? 4'b1000 : 4'b1001;
														assign node17544 = (inp[9]) ? node17550 : node17545;
															assign node17545 = (inp[2]) ? 4'b1001 : node17546;
																assign node17546 = (inp[0]) ? 4'b1001 : 4'b1000;
															assign node17550 = (inp[0]) ? 4'b1000 : node17551;
																assign node17551 = (inp[2]) ? 4'b1000 : 4'b1001;
													assign node17555 = (inp[2]) ? node17569 : node17556;
														assign node17556 = (inp[0]) ? node17564 : node17557;
															assign node17557 = (inp[11]) ? node17561 : node17558;
																assign node17558 = (inp[9]) ? 4'b1000 : 4'b1001;
																assign node17561 = (inp[9]) ? 4'b1001 : 4'b1000;
															assign node17564 = (inp[11]) ? 4'b1000 : node17565;
																assign node17565 = (inp[9]) ? 4'b1001 : 4'b1000;
														assign node17569 = (inp[11]) ? node17573 : node17570;
															assign node17570 = (inp[9]) ? 4'b1001 : 4'b1000;
															assign node17573 = (inp[9]) ? 4'b1000 : 4'b1001;
								assign node17576 = (inp[15]) ? node17902 : node17577;
									assign node17577 = (inp[7]) ? node17721 : node17578;
										assign node17578 = (inp[1]) ? node17674 : node17579;
											assign node17579 = (inp[10]) ? node17629 : node17580;
												assign node17580 = (inp[2]) ? node17610 : node17581;
													assign node17581 = (inp[11]) ? node17597 : node17582;
														assign node17582 = (inp[0]) ? node17590 : node17583;
															assign node17583 = (inp[9]) ? node17587 : node17584;
																assign node17584 = (inp[4]) ? 4'b1000 : 4'b1001;
																assign node17587 = (inp[4]) ? 4'b1001 : 4'b1000;
															assign node17590 = (inp[4]) ? node17594 : node17591;
																assign node17591 = (inp[9]) ? 4'b1001 : 4'b1000;
																assign node17594 = (inp[9]) ? 4'b1000 : 4'b1001;
														assign node17597 = (inp[9]) ? node17605 : node17598;
															assign node17598 = (inp[4]) ? node17602 : node17599;
																assign node17599 = (inp[0]) ? 4'b1001 : 4'b1000;
																assign node17602 = (inp[0]) ? 4'b1000 : 4'b1001;
															assign node17605 = (inp[0]) ? node17607 : 4'b1000;
																assign node17607 = (inp[4]) ? 4'b1001 : 4'b1000;
													assign node17610 = (inp[4]) ? node17622 : node17611;
														assign node17611 = (inp[0]) ? node17617 : node17612;
															assign node17612 = (inp[9]) ? node17614 : 4'b1000;
																assign node17614 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node17617 = (inp[9]) ? 4'b1001 : node17618;
																assign node17618 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node17622 = (inp[0]) ? 4'b1000 : node17623;
															assign node17623 = (inp[11]) ? 4'b1001 : node17624;
																assign node17624 = (inp[9]) ? 4'b1000 : 4'b1001;
												assign node17629 = (inp[4]) ? node17651 : node17630;
													assign node17630 = (inp[9]) ? node17640 : node17631;
														assign node17631 = (inp[11]) ? node17637 : node17632;
															assign node17632 = (inp[2]) ? 4'b1001 : node17633;
																assign node17633 = (inp[0]) ? 4'b1000 : 4'b1001;
															assign node17637 = (inp[0]) ? 4'b1001 : 4'b1000;
														assign node17640 = (inp[11]) ? node17646 : node17641;
															assign node17641 = (inp[2]) ? 4'b1000 : node17642;
																assign node17642 = (inp[0]) ? 4'b1001 : 4'b1000;
															assign node17646 = (inp[0]) ? node17648 : 4'b1001;
																assign node17648 = (inp[2]) ? 4'b1001 : 4'b1000;
													assign node17651 = (inp[9]) ? node17663 : node17652;
														assign node17652 = (inp[11]) ? node17658 : node17653;
															assign node17653 = (inp[2]) ? 4'b1001 : node17654;
																assign node17654 = (inp[0]) ? 4'b1001 : 4'b1000;
															assign node17658 = (inp[2]) ? 4'b1000 : node17659;
																assign node17659 = (inp[0]) ? 4'b1000 : 4'b1001;
														assign node17663 = (inp[11]) ? node17669 : node17664;
															assign node17664 = (inp[0]) ? 4'b1000 : node17665;
																assign node17665 = (inp[2]) ? 4'b1000 : 4'b1001;
															assign node17669 = (inp[2]) ? 4'b1001 : node17670;
																assign node17670 = (inp[0]) ? 4'b1001 : 4'b1000;
											assign node17674 = (inp[4]) ? node17698 : node17675;
												assign node17675 = (inp[0]) ? node17691 : node17676;
													assign node17676 = (inp[2]) ? node17684 : node17677;
														assign node17677 = (inp[9]) ? node17681 : node17678;
															assign node17678 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node17681 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node17684 = (inp[11]) ? node17688 : node17685;
															assign node17685 = (inp[9]) ? 4'b1000 : 4'b1001;
															assign node17688 = (inp[9]) ? 4'b1001 : 4'b1000;
													assign node17691 = (inp[11]) ? node17695 : node17692;
														assign node17692 = (inp[9]) ? 4'b1001 : 4'b1000;
														assign node17695 = (inp[9]) ? 4'b1000 : 4'b1001;
												assign node17698 = (inp[9]) ? node17710 : node17699;
													assign node17699 = (inp[11]) ? node17705 : node17700;
														assign node17700 = (inp[2]) ? 4'b1100 : node17701;
															assign node17701 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node17705 = (inp[2]) ? 4'b1101 : node17706;
															assign node17706 = (inp[0]) ? 4'b1101 : 4'b1100;
													assign node17710 = (inp[11]) ? node17716 : node17711;
														assign node17711 = (inp[2]) ? 4'b1101 : node17712;
															assign node17712 = (inp[0]) ? 4'b1101 : 4'b1100;
														assign node17716 = (inp[0]) ? 4'b1100 : node17717;
															assign node17717 = (inp[2]) ? 4'b1100 : 4'b1101;
										assign node17721 = (inp[1]) ? node17811 : node17722;
											assign node17722 = (inp[4]) ? node17762 : node17723;
												assign node17723 = (inp[2]) ? node17747 : node17724;
													assign node17724 = (inp[0]) ? node17732 : node17725;
														assign node17725 = (inp[9]) ? node17729 : node17726;
															assign node17726 = (inp[11]) ? 4'b1111 : 4'b1110;
															assign node17729 = (inp[11]) ? 4'b1110 : 4'b1111;
														assign node17732 = (inp[10]) ? node17740 : node17733;
															assign node17733 = (inp[9]) ? node17737 : node17734;
																assign node17734 = (inp[11]) ? 4'b1111 : 4'b1110;
																assign node17737 = (inp[11]) ? 4'b1110 : 4'b1111;
															assign node17740 = (inp[11]) ? node17744 : node17741;
																assign node17741 = (inp[9]) ? 4'b1111 : 4'b1110;
																assign node17744 = (inp[9]) ? 4'b1110 : 4'b1111;
													assign node17747 = (inp[11]) ? node17755 : node17748;
														assign node17748 = (inp[9]) ? node17752 : node17749;
															assign node17749 = (inp[0]) ? 4'b1110 : 4'b1111;
															assign node17752 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node17755 = (inp[0]) ? node17759 : node17756;
															assign node17756 = (inp[9]) ? 4'b1111 : 4'b1110;
															assign node17759 = (inp[9]) ? 4'b1110 : 4'b1111;
												assign node17762 = (inp[10]) ? node17790 : node17763;
													assign node17763 = (inp[2]) ? node17777 : node17764;
														assign node17764 = (inp[0]) ? node17772 : node17765;
															assign node17765 = (inp[9]) ? node17769 : node17766;
																assign node17766 = (inp[11]) ? 4'b1010 : 4'b1011;
																assign node17769 = (inp[11]) ? 4'b1011 : 4'b1010;
															assign node17772 = (inp[11]) ? node17774 : 4'b1011;
																assign node17774 = (inp[9]) ? 4'b1011 : 4'b1010;
														assign node17777 = (inp[0]) ? node17785 : node17778;
															assign node17778 = (inp[9]) ? node17782 : node17779;
																assign node17779 = (inp[11]) ? 4'b1010 : 4'b1011;
																assign node17782 = (inp[11]) ? 4'b1011 : 4'b1010;
															assign node17785 = (inp[11]) ? 4'b1010 : node17786;
																assign node17786 = (inp[9]) ? 4'b1011 : 4'b1010;
													assign node17790 = (inp[0]) ? node17798 : node17791;
														assign node17791 = (inp[9]) ? node17795 : node17792;
															assign node17792 = (inp[11]) ? 4'b1010 : 4'b1011;
															assign node17795 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node17798 = (inp[9]) ? node17804 : node17799;
															assign node17799 = (inp[2]) ? 4'b1010 : node17800;
																assign node17800 = (inp[11]) ? 4'b1010 : 4'b1011;
															assign node17804 = (inp[2]) ? node17808 : node17805;
																assign node17805 = (inp[11]) ? 4'b1011 : 4'b1010;
																assign node17808 = (inp[11]) ? 4'b1010 : 4'b1011;
											assign node17811 = (inp[10]) ? node17859 : node17812;
												assign node17812 = (inp[4]) ? node17838 : node17813;
													assign node17813 = (inp[2]) ? node17827 : node17814;
														assign node17814 = (inp[11]) ? node17822 : node17815;
															assign node17815 = (inp[9]) ? node17819 : node17816;
																assign node17816 = (inp[0]) ? 4'b1011 : 4'b1010;
																assign node17819 = (inp[0]) ? 4'b1010 : 4'b1011;
															assign node17822 = (inp[9]) ? 4'b1010 : node17823;
																assign node17823 = (inp[0]) ? 4'b1010 : 4'b1011;
														assign node17827 = (inp[0]) ? node17833 : node17828;
															assign node17828 = (inp[11]) ? 4'b1010 : node17829;
																assign node17829 = (inp[9]) ? 4'b1011 : 4'b1010;
															assign node17833 = (inp[9]) ? 4'b1010 : node17834;
																assign node17834 = (inp[11]) ? 4'b1011 : 4'b1010;
													assign node17838 = (inp[9]) ? node17848 : node17839;
														assign node17839 = (inp[11]) ? node17843 : node17840;
															assign node17840 = (inp[2]) ? 4'b1010 : 4'b1011;
															assign node17843 = (inp[0]) ? 4'b1011 : node17844;
																assign node17844 = (inp[2]) ? 4'b1011 : 4'b1010;
														assign node17848 = (inp[11]) ? node17854 : node17849;
															assign node17849 = (inp[2]) ? 4'b1011 : node17850;
																assign node17850 = (inp[0]) ? 4'b1011 : 4'b1010;
															assign node17854 = (inp[2]) ? 4'b1010 : node17855;
																assign node17855 = (inp[0]) ? 4'b1010 : 4'b1011;
												assign node17859 = (inp[0]) ? node17879 : node17860;
													assign node17860 = (inp[9]) ? node17870 : node17861;
														assign node17861 = (inp[11]) ? node17865 : node17862;
															assign node17862 = (inp[4]) ? 4'b1011 : 4'b1010;
															assign node17865 = (inp[4]) ? node17867 : 4'b1011;
																assign node17867 = (inp[2]) ? 4'b1011 : 4'b1010;
														assign node17870 = (inp[11]) ? node17876 : node17871;
															assign node17871 = (inp[4]) ? node17873 : 4'b1011;
																assign node17873 = (inp[2]) ? 4'b1011 : 4'b1010;
															assign node17876 = (inp[2]) ? 4'b1010 : 4'b1011;
													assign node17879 = (inp[9]) ? node17891 : node17880;
														assign node17880 = (inp[11]) ? node17886 : node17881;
															assign node17881 = (inp[4]) ? 4'b1010 : node17882;
																assign node17882 = (inp[2]) ? 4'b1010 : 4'b1011;
															assign node17886 = (inp[2]) ? 4'b1011 : node17887;
																assign node17887 = (inp[4]) ? 4'b1011 : 4'b1010;
														assign node17891 = (inp[11]) ? node17897 : node17892;
															assign node17892 = (inp[4]) ? 4'b1011 : node17893;
																assign node17893 = (inp[2]) ? 4'b1011 : 4'b1010;
															assign node17897 = (inp[4]) ? 4'b1010 : node17898;
																assign node17898 = (inp[2]) ? 4'b1010 : 4'b1011;
									assign node17902 = (inp[7]) ? node18036 : node17903;
										assign node17903 = (inp[4]) ? node17973 : node17904;
											assign node17904 = (inp[2]) ? node17942 : node17905;
												assign node17905 = (inp[11]) ? node17935 : node17906;
													assign node17906 = (inp[10]) ? node17922 : node17907;
														assign node17907 = (inp[1]) ? node17915 : node17908;
															assign node17908 = (inp[9]) ? node17912 : node17909;
																assign node17909 = (inp[0]) ? 4'b1011 : 4'b1010;
																assign node17912 = (inp[0]) ? 4'b1010 : 4'b1011;
															assign node17915 = (inp[9]) ? node17919 : node17916;
																assign node17916 = (inp[0]) ? 4'b1011 : 4'b1010;
																assign node17919 = (inp[0]) ? 4'b1010 : 4'b1011;
														assign node17922 = (inp[1]) ? node17928 : node17923;
															assign node17923 = (inp[0]) ? node17925 : 4'b1011;
																assign node17925 = (inp[9]) ? 4'b1010 : 4'b1011;
															assign node17928 = (inp[0]) ? node17932 : node17929;
																assign node17929 = (inp[9]) ? 4'b1011 : 4'b1010;
																assign node17932 = (inp[9]) ? 4'b1010 : 4'b1011;
													assign node17935 = (inp[0]) ? node17939 : node17936;
														assign node17936 = (inp[9]) ? 4'b1010 : 4'b1011;
														assign node17939 = (inp[9]) ? 4'b1011 : 4'b1010;
												assign node17942 = (inp[10]) ? node17966 : node17943;
													assign node17943 = (inp[1]) ? node17959 : node17944;
														assign node17944 = (inp[0]) ? node17952 : node17945;
															assign node17945 = (inp[9]) ? node17949 : node17946;
																assign node17946 = (inp[11]) ? 4'b1011 : 4'b1010;
																assign node17949 = (inp[11]) ? 4'b1010 : 4'b1011;
															assign node17952 = (inp[9]) ? node17956 : node17953;
																assign node17953 = (inp[11]) ? 4'b1011 : 4'b1010;
																assign node17956 = (inp[11]) ? 4'b1010 : 4'b1011;
														assign node17959 = (inp[11]) ? node17963 : node17960;
															assign node17960 = (inp[9]) ? 4'b1011 : 4'b1010;
															assign node17963 = (inp[9]) ? 4'b1010 : 4'b1011;
													assign node17966 = (inp[9]) ? node17970 : node17967;
														assign node17967 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node17970 = (inp[11]) ? 4'b1010 : 4'b1011;
											assign node17973 = (inp[10]) ? node18013 : node17974;
												assign node17974 = (inp[1]) ? node17990 : node17975;
													assign node17975 = (inp[0]) ? node17983 : node17976;
														assign node17976 = (inp[2]) ? 4'b1011 : node17977;
															assign node17977 = (inp[9]) ? node17979 : 4'b1011;
																assign node17979 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node17983 = (inp[9]) ? node17987 : node17984;
															assign node17984 = (inp[11]) ? 4'b1011 : 4'b1010;
															assign node17987 = (inp[11]) ? 4'b1010 : 4'b1011;
													assign node17990 = (inp[2]) ? node18006 : node17991;
														assign node17991 = (inp[9]) ? node17999 : node17992;
															assign node17992 = (inp[11]) ? node17996 : node17993;
																assign node17993 = (inp[0]) ? 4'b1010 : 4'b1011;
																assign node17996 = (inp[0]) ? 4'b1011 : 4'b1010;
															assign node17999 = (inp[0]) ? node18003 : node18000;
																assign node18000 = (inp[11]) ? 4'b1011 : 4'b1010;
																assign node18003 = (inp[11]) ? 4'b1010 : 4'b1011;
														assign node18006 = (inp[11]) ? node18010 : node18007;
															assign node18007 = (inp[9]) ? 4'b1011 : 4'b1010;
															assign node18010 = (inp[9]) ? 4'b1010 : 4'b1011;
												assign node18013 = (inp[9]) ? node18025 : node18014;
													assign node18014 = (inp[11]) ? node18020 : node18015;
														assign node18015 = (inp[0]) ? 4'b1010 : node18016;
															assign node18016 = (inp[2]) ? 4'b1010 : 4'b1011;
														assign node18020 = (inp[0]) ? 4'b1011 : node18021;
															assign node18021 = (inp[2]) ? 4'b1011 : 4'b1010;
													assign node18025 = (inp[11]) ? node18031 : node18026;
														assign node18026 = (inp[2]) ? 4'b1011 : node18027;
															assign node18027 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node18031 = (inp[0]) ? 4'b1010 : node18032;
															assign node18032 = (inp[2]) ? 4'b1010 : 4'b1011;
										assign node18036 = (inp[11]) ? node18064 : node18037;
											assign node18037 = (inp[9]) ? node18055 : node18038;
												assign node18038 = (inp[2]) ? 4'b1000 : node18039;
													assign node18039 = (inp[1]) ? node18047 : node18040;
														assign node18040 = (inp[4]) ? node18044 : node18041;
															assign node18041 = (inp[0]) ? 4'b1001 : 4'b1000;
															assign node18044 = (inp[0]) ? 4'b1000 : 4'b1001;
														assign node18047 = (inp[0]) ? node18051 : node18048;
															assign node18048 = (inp[4]) ? 4'b1001 : 4'b1000;
															assign node18051 = (inp[4]) ? 4'b1000 : 4'b1001;
												assign node18055 = (inp[2]) ? 4'b1001 : node18056;
													assign node18056 = (inp[4]) ? node18060 : node18057;
														assign node18057 = (inp[0]) ? 4'b1000 : 4'b1001;
														assign node18060 = (inp[0]) ? 4'b1001 : 4'b1000;
											assign node18064 = (inp[9]) ? node18080 : node18065;
												assign node18065 = (inp[2]) ? 4'b1001 : node18066;
													assign node18066 = (inp[1]) ? node18072 : node18067;
														assign node18067 = (inp[4]) ? node18069 : 4'b1000;
															assign node18069 = (inp[0]) ? 4'b1001 : 4'b1000;
														assign node18072 = (inp[0]) ? node18076 : node18073;
															assign node18073 = (inp[4]) ? 4'b1000 : 4'b1001;
															assign node18076 = (inp[4]) ? 4'b1001 : 4'b1000;
												assign node18080 = (inp[2]) ? 4'b1000 : node18081;
													assign node18081 = (inp[10]) ? node18089 : node18082;
														assign node18082 = (inp[0]) ? node18086 : node18083;
															assign node18083 = (inp[4]) ? 4'b1001 : 4'b1000;
															assign node18086 = (inp[4]) ? 4'b1000 : 4'b1001;
														assign node18089 = (inp[1]) ? node18097 : node18090;
															assign node18090 = (inp[4]) ? node18094 : node18091;
																assign node18091 = (inp[0]) ? 4'b1001 : 4'b1000;
																assign node18094 = (inp[0]) ? 4'b1000 : 4'b1001;
															assign node18097 = (inp[0]) ? node18099 : 4'b1001;
																assign node18099 = (inp[4]) ? 4'b1000 : 4'b1001;
			assign node18103 = (inp[3]) ? node24273 : node18104;
				assign node18104 = (inp[6]) ? node21056 : node18105;
					assign node18105 = (inp[10]) ? node19593 : node18106;
						assign node18106 = (inp[0]) ? node18926 : node18107;
							assign node18107 = (inp[7]) ? node18441 : node18108;
								assign node18108 = (inp[13]) ? node18230 : node18109;
									assign node18109 = (inp[1]) ? node18153 : node18110;
										assign node18110 = (inp[2]) ? node18132 : node18111;
											assign node18111 = (inp[4]) ? node18115 : node18112;
												assign node18112 = (inp[12]) ? 4'b1010 : 4'b1000;
												assign node18115 = (inp[12]) ? node18125 : node18116;
													assign node18116 = (inp[5]) ? node18118 : 4'b1010;
														assign node18118 = (inp[11]) ? node18122 : node18119;
															assign node18119 = (inp[15]) ? 4'b1110 : 4'b1010;
															assign node18122 = (inp[15]) ? 4'b1111 : 4'b1011;
													assign node18125 = (inp[5]) ? 4'b1001 : node18126;
														assign node18126 = (inp[15]) ? node18128 : 4'b1100;
															assign node18128 = (inp[11]) ? 4'b1001 : 4'b1000;
											assign node18132 = (inp[4]) ? node18136 : node18133;
												assign node18133 = (inp[12]) ? 4'b1110 : 4'b1100;
												assign node18136 = (inp[12]) ? node18144 : node18137;
													assign node18137 = (inp[5]) ? node18139 : 4'b1111;
														assign node18139 = (inp[15]) ? 4'b1010 : node18140;
															assign node18140 = (inp[11]) ? 4'b1110 : 4'b1111;
													assign node18144 = (inp[5]) ? 4'b1100 : node18145;
														assign node18145 = (inp[15]) ? node18149 : node18146;
															assign node18146 = (inp[11]) ? 4'b1000 : 4'b1001;
															assign node18149 = (inp[11]) ? 4'b1100 : 4'b1101;
										assign node18153 = (inp[2]) ? node18193 : node18154;
											assign node18154 = (inp[4]) ? node18166 : node18155;
												assign node18155 = (inp[12]) ? node18161 : node18156;
													assign node18156 = (inp[11]) ? node18158 : 4'b1100;
														assign node18158 = (inp[15]) ? 4'b1101 : 4'b1100;
													assign node18161 = (inp[15]) ? node18163 : 4'b1111;
														assign node18163 = (inp[11]) ? 4'b1110 : 4'b1111;
												assign node18166 = (inp[12]) ? node18182 : node18167;
													assign node18167 = (inp[5]) ? node18175 : node18168;
														assign node18168 = (inp[9]) ? 4'b1110 : node18169;
															assign node18169 = (inp[11]) ? node18171 : 4'b1110;
																assign node18171 = (inp[15]) ? 4'b1111 : 4'b1110;
														assign node18175 = (inp[15]) ? node18179 : node18176;
															assign node18176 = (inp[11]) ? 4'b1111 : 4'b1110;
															assign node18179 = (inp[11]) ? 4'b1010 : 4'b1011;
													assign node18182 = (inp[5]) ? node18188 : node18183;
														assign node18183 = (inp[15]) ? 4'b1100 : node18184;
															assign node18184 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node18188 = (inp[11]) ? node18190 : 4'b1100;
															assign node18190 = (inp[15]) ? 4'b1101 : 4'b1100;
											assign node18193 = (inp[4]) ? node18205 : node18194;
												assign node18194 = (inp[12]) ? node18200 : node18195;
													assign node18195 = (inp[11]) ? 4'b1001 : node18196;
														assign node18196 = (inp[15]) ? 4'b1001 : 4'b1000;
													assign node18200 = (inp[11]) ? 4'b1010 : node18201;
														assign node18201 = (inp[15]) ? 4'b1010 : 4'b1011;
												assign node18205 = (inp[12]) ? node18217 : node18206;
													assign node18206 = (inp[5]) ? node18212 : node18207;
														assign node18207 = (inp[11]) ? 4'b1010 : node18208;
															assign node18208 = (inp[15]) ? 4'b1010 : 4'b1011;
														assign node18212 = (inp[15]) ? node18214 : 4'b1010;
															assign node18214 = (inp[11]) ? 4'b1111 : 4'b1110;
													assign node18217 = (inp[15]) ? node18225 : node18218;
														assign node18218 = (inp[5]) ? node18222 : node18219;
															assign node18219 = (inp[11]) ? 4'b1101 : 4'b1100;
															assign node18222 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node18225 = (inp[5]) ? 4'b1000 : node18226;
															assign node18226 = (inp[11]) ? 4'b1000 : 4'b1001;
									assign node18230 = (inp[5]) ? node18336 : node18231;
										assign node18231 = (inp[2]) ? node18287 : node18232;
											assign node18232 = (inp[1]) ? node18264 : node18233;
												assign node18233 = (inp[15]) ? node18249 : node18234;
													assign node18234 = (inp[11]) ? node18242 : node18235;
														assign node18235 = (inp[4]) ? node18239 : node18236;
															assign node18236 = (inp[12]) ? 4'b1010 : 4'b1000;
															assign node18239 = (inp[12]) ? 4'b1100 : 4'b1010;
														assign node18242 = (inp[12]) ? node18246 : node18243;
															assign node18243 = (inp[4]) ? 4'b1011 : 4'b1001;
															assign node18246 = (inp[4]) ? 4'b1101 : 4'b1011;
													assign node18249 = (inp[11]) ? node18257 : node18250;
														assign node18250 = (inp[12]) ? node18254 : node18251;
															assign node18251 = (inp[4]) ? 4'b1011 : 4'b1001;
															assign node18254 = (inp[4]) ? 4'b1000 : 4'b1011;
														assign node18257 = (inp[12]) ? node18261 : node18258;
															assign node18258 = (inp[4]) ? 4'b1010 : 4'b1000;
															assign node18261 = (inp[4]) ? 4'b1000 : 4'b1010;
												assign node18264 = (inp[12]) ? node18276 : node18265;
													assign node18265 = (inp[4]) ? node18271 : node18266;
														assign node18266 = (inp[11]) ? node18268 : 4'b1100;
															assign node18268 = (inp[15]) ? 4'b1100 : 4'b1101;
														assign node18271 = (inp[11]) ? node18273 : 4'b1110;
															assign node18273 = (inp[15]) ? 4'b1110 : 4'b1111;
													assign node18276 = (inp[4]) ? node18282 : node18277;
														assign node18277 = (inp[15]) ? 4'b1111 : node18278;
															assign node18278 = (inp[11]) ? 4'b1110 : 4'b1111;
														assign node18282 = (inp[15]) ? node18284 : 4'b1000;
															assign node18284 = (inp[11]) ? 4'b1100 : 4'b1101;
											assign node18287 = (inp[1]) ? node18315 : node18288;
												assign node18288 = (inp[15]) ? node18302 : node18289;
													assign node18289 = (inp[4]) ? node18297 : node18290;
														assign node18290 = (inp[11]) ? node18294 : node18291;
															assign node18291 = (inp[12]) ? 4'b1110 : 4'b1100;
															assign node18294 = (inp[12]) ? 4'b1111 : 4'b1101;
														assign node18297 = (inp[12]) ? 4'b1000 : node18298;
															assign node18298 = (inp[11]) ? 4'b1110 : 4'b1111;
													assign node18302 = (inp[11]) ? node18310 : node18303;
														assign node18303 = (inp[4]) ? node18307 : node18304;
															assign node18304 = (inp[12]) ? 4'b1111 : 4'b1101;
															assign node18307 = (inp[12]) ? 4'b1101 : 4'b1110;
														assign node18310 = (inp[4]) ? node18312 : 4'b1110;
															assign node18312 = (inp[12]) ? 4'b1101 : 4'b1111;
												assign node18315 = (inp[15]) ? node18323 : node18316;
													assign node18316 = (inp[4]) ? node18320 : node18317;
														assign node18317 = (inp[12]) ? 4'b1010 : 4'b1001;
														assign node18320 = (inp[12]) ? 4'b1101 : 4'b1010;
													assign node18323 = (inp[12]) ? node18331 : node18324;
														assign node18324 = (inp[4]) ? node18328 : node18325;
															assign node18325 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node18328 = (inp[11]) ? 4'b1010 : 4'b1011;
														assign node18331 = (inp[4]) ? 4'b1001 : node18332;
															assign node18332 = (inp[11]) ? 4'b1010 : 4'b1011;
										assign node18336 = (inp[2]) ? node18386 : node18337;
											assign node18337 = (inp[1]) ? node18365 : node18338;
												assign node18338 = (inp[15]) ? node18352 : node18339;
													assign node18339 = (inp[4]) ? node18347 : node18340;
														assign node18340 = (inp[11]) ? node18344 : node18341;
															assign node18341 = (inp[12]) ? 4'b1010 : 4'b1000;
															assign node18344 = (inp[12]) ? 4'b1011 : 4'b1001;
														assign node18347 = (inp[12]) ? node18349 : 4'b1011;
															assign node18349 = (inp[11]) ? 4'b1000 : 4'b1001;
													assign node18352 = (inp[4]) ? node18360 : node18353;
														assign node18353 = (inp[11]) ? node18357 : node18354;
															assign node18354 = (inp[12]) ? 4'b1011 : 4'b1001;
															assign node18357 = (inp[12]) ? 4'b1010 : 4'b1000;
														assign node18360 = (inp[12]) ? node18362 : 4'b1110;
															assign node18362 = (inp[11]) ? 4'b1001 : 4'b1000;
												assign node18365 = (inp[15]) ? node18379 : node18366;
													assign node18366 = (inp[12]) ? node18372 : node18367;
														assign node18367 = (inp[4]) ? 4'b1111 : node18368;
															assign node18368 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node18372 = (inp[4]) ? node18376 : node18373;
															assign node18373 = (inp[11]) ? 4'b1110 : 4'b1111;
															assign node18376 = (inp[11]) ? 4'b1101 : 4'b1100;
													assign node18379 = (inp[12]) ? node18383 : node18380;
														assign node18380 = (inp[4]) ? 4'b1011 : 4'b1100;
														assign node18383 = (inp[4]) ? 4'b1100 : 4'b1111;
											assign node18386 = (inp[1]) ? node18418 : node18387;
												assign node18387 = (inp[15]) ? node18403 : node18388;
													assign node18388 = (inp[11]) ? node18396 : node18389;
														assign node18389 = (inp[12]) ? node18393 : node18390;
															assign node18390 = (inp[4]) ? 4'b1110 : 4'b1100;
															assign node18393 = (inp[4]) ? 4'b1100 : 4'b1110;
														assign node18396 = (inp[12]) ? node18400 : node18397;
															assign node18397 = (inp[4]) ? 4'b1110 : 4'b1101;
															assign node18400 = (inp[4]) ? 4'b1101 : 4'b1111;
													assign node18403 = (inp[11]) ? node18411 : node18404;
														assign node18404 = (inp[4]) ? node18408 : node18405;
															assign node18405 = (inp[12]) ? 4'b1111 : 4'b1101;
															assign node18408 = (inp[12]) ? 4'b1101 : 4'b1011;
														assign node18411 = (inp[12]) ? node18415 : node18412;
															assign node18412 = (inp[4]) ? 4'b1010 : 4'b1100;
															assign node18415 = (inp[4]) ? 4'b1100 : 4'b1110;
												assign node18418 = (inp[12]) ? node18430 : node18419;
													assign node18419 = (inp[4]) ? node18425 : node18420;
														assign node18420 = (inp[15]) ? node18422 : 4'b1001;
															assign node18422 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node18425 = (inp[15]) ? 4'b1110 : node18426;
															assign node18426 = (inp[11]) ? 4'b1011 : 4'b1010;
													assign node18430 = (inp[4]) ? node18436 : node18431;
														assign node18431 = (inp[15]) ? node18433 : 4'b1010;
															assign node18433 = (inp[11]) ? 4'b1010 : 4'b1011;
														assign node18436 = (inp[15]) ? node18438 : 4'b1000;
															assign node18438 = (inp[11]) ? 4'b1000 : 4'b1001;
								assign node18441 = (inp[13]) ? node18693 : node18442;
									assign node18442 = (inp[15]) ? node18570 : node18443;
										assign node18443 = (inp[5]) ? node18493 : node18444;
											assign node18444 = (inp[12]) ? node18470 : node18445;
												assign node18445 = (inp[4]) ? node18461 : node18446;
													assign node18446 = (inp[11]) ? node18454 : node18447;
														assign node18447 = (inp[2]) ? node18451 : node18448;
															assign node18448 = (inp[1]) ? 4'b1100 : 4'b1000;
															assign node18451 = (inp[1]) ? 4'b1000 : 4'b1100;
														assign node18454 = (inp[1]) ? node18458 : node18455;
															assign node18455 = (inp[2]) ? 4'b1100 : 4'b1000;
															assign node18458 = (inp[2]) ? 4'b1001 : 4'b1100;
													assign node18461 = (inp[2]) ? node18465 : node18462;
														assign node18462 = (inp[1]) ? 4'b1110 : 4'b1010;
														assign node18465 = (inp[1]) ? node18467 : 4'b1111;
															assign node18467 = (inp[11]) ? 4'b1010 : 4'b1011;
												assign node18470 = (inp[4]) ? node18484 : node18471;
													assign node18471 = (inp[2]) ? node18479 : node18472;
														assign node18472 = (inp[1]) ? node18476 : node18473;
															assign node18473 = (inp[11]) ? 4'b1011 : 4'b1010;
															assign node18476 = (inp[11]) ? 4'b1110 : 4'b1111;
														assign node18479 = (inp[1]) ? 4'b1010 : node18480;
															assign node18480 = (inp[11]) ? 4'b1111 : 4'b1110;
													assign node18484 = (inp[1]) ? node18488 : node18485;
														assign node18485 = (inp[2]) ? 4'b1100 : 4'b1001;
														assign node18488 = (inp[2]) ? node18490 : 4'b1100;
															assign node18490 = (inp[11]) ? 4'b1000 : 4'b1001;
											assign node18493 = (inp[11]) ? node18533 : node18494;
												assign node18494 = (inp[4]) ? node18518 : node18495;
													assign node18495 = (inp[12]) ? node18511 : node18496;
														assign node18496 = (inp[9]) ? node18504 : node18497;
															assign node18497 = (inp[1]) ? node18501 : node18498;
																assign node18498 = (inp[2]) ? 4'b1001 : 4'b1101;
																assign node18501 = (inp[2]) ? 4'b1101 : 4'b1001;
															assign node18504 = (inp[1]) ? node18508 : node18505;
																assign node18505 = (inp[2]) ? 4'b1001 : 4'b1101;
																assign node18508 = (inp[2]) ? 4'b1101 : 4'b1001;
														assign node18511 = (inp[2]) ? node18515 : node18512;
															assign node18512 = (inp[1]) ? 4'b1011 : 4'b1111;
															assign node18515 = (inp[1]) ? 4'b1111 : 4'b1010;
													assign node18518 = (inp[12]) ? node18526 : node18519;
														assign node18519 = (inp[2]) ? node18523 : node18520;
															assign node18520 = (inp[1]) ? 4'b1010 : 4'b1111;
															assign node18523 = (inp[1]) ? 4'b1111 : 4'b1011;
														assign node18526 = (inp[1]) ? node18530 : node18527;
															assign node18527 = (inp[2]) ? 4'b1101 : 4'b1000;
															assign node18530 = (inp[2]) ? 4'b1001 : 4'b1101;
												assign node18533 = (inp[12]) ? node18549 : node18534;
													assign node18534 = (inp[4]) ? node18542 : node18535;
														assign node18535 = (inp[1]) ? node18539 : node18536;
															assign node18536 = (inp[2]) ? 4'b1000 : 4'b1101;
															assign node18539 = (inp[2]) ? 4'b1100 : 4'b1000;
														assign node18542 = (inp[2]) ? node18546 : node18543;
															assign node18543 = (inp[1]) ? 4'b1010 : 4'b1110;
															assign node18546 = (inp[1]) ? 4'b1111 : 4'b1011;
													assign node18549 = (inp[4]) ? node18557 : node18550;
														assign node18550 = (inp[1]) ? node18554 : node18551;
															assign node18551 = (inp[2]) ? 4'b1010 : 4'b1110;
															assign node18554 = (inp[2]) ? 4'b1111 : 4'b1011;
														assign node18557 = (inp[9]) ? node18565 : node18558;
															assign node18558 = (inp[1]) ? node18562 : node18559;
																assign node18559 = (inp[2]) ? 4'b1100 : 4'b1001;
																assign node18562 = (inp[2]) ? 4'b1001 : 4'b1100;
															assign node18565 = (inp[2]) ? 4'b1100 : node18566;
																assign node18566 = (inp[1]) ? 4'b1100 : 4'b1001;
										assign node18570 = (inp[5]) ? node18642 : node18571;
											assign node18571 = (inp[11]) ? node18603 : node18572;
												assign node18572 = (inp[1]) ? node18588 : node18573;
													assign node18573 = (inp[2]) ? node18581 : node18574;
														assign node18574 = (inp[12]) ? node18578 : node18575;
															assign node18575 = (inp[4]) ? 4'b1010 : 4'b1100;
															assign node18578 = (inp[4]) ? 4'b1101 : 4'b1110;
														assign node18581 = (inp[12]) ? node18585 : node18582;
															assign node18582 = (inp[4]) ? 4'b1111 : 4'b1000;
															assign node18585 = (inp[4]) ? 4'b1000 : 4'b1011;
													assign node18588 = (inp[2]) ? node18596 : node18589;
														assign node18589 = (inp[4]) ? node18593 : node18590;
															assign node18590 = (inp[12]) ? 4'b1010 : 4'b1001;
															assign node18593 = (inp[12]) ? 4'b1001 : 4'b1111;
														assign node18596 = (inp[4]) ? node18600 : node18597;
															assign node18597 = (inp[12]) ? 4'b1110 : 4'b1101;
															assign node18600 = (inp[12]) ? 4'b1100 : 4'b1010;
												assign node18603 = (inp[12]) ? node18619 : node18604;
													assign node18604 = (inp[4]) ? node18612 : node18605;
														assign node18605 = (inp[1]) ? node18609 : node18606;
															assign node18606 = (inp[2]) ? 4'b1001 : 4'b1100;
															assign node18609 = (inp[2]) ? 4'b1101 : 4'b1001;
														assign node18612 = (inp[1]) ? node18616 : node18613;
															assign node18613 = (inp[2]) ? 4'b1110 : 4'b1011;
															assign node18616 = (inp[2]) ? 4'b1011 : 4'b1111;
													assign node18619 = (inp[4]) ? node18635 : node18620;
														assign node18620 = (inp[9]) ? node18628 : node18621;
															assign node18621 = (inp[1]) ? node18625 : node18622;
																assign node18622 = (inp[2]) ? 4'b1011 : 4'b1111;
																assign node18625 = (inp[2]) ? 4'b1111 : 4'b1011;
															assign node18628 = (inp[1]) ? node18632 : node18629;
																assign node18629 = (inp[2]) ? 4'b1011 : 4'b1111;
																assign node18632 = (inp[2]) ? 4'b1111 : 4'b1011;
														assign node18635 = (inp[1]) ? node18639 : node18636;
															assign node18636 = (inp[2]) ? 4'b1001 : 4'b1101;
															assign node18639 = (inp[2]) ? 4'b1100 : 4'b1001;
											assign node18642 = (inp[2]) ? node18674 : node18643;
												assign node18643 = (inp[1]) ? node18659 : node18644;
													assign node18644 = (inp[11]) ? node18652 : node18645;
														assign node18645 = (inp[12]) ? node18649 : node18646;
															assign node18646 = (inp[4]) ? 4'b1010 : 4'b1001;
															assign node18649 = (inp[4]) ? 4'b1001 : 4'b1010;
														assign node18652 = (inp[12]) ? node18656 : node18653;
															assign node18653 = (inp[4]) ? 4'b1010 : 4'b1000;
															assign node18656 = (inp[4]) ? 4'b1001 : 4'b1010;
													assign node18659 = (inp[11]) ? node18667 : node18660;
														assign node18660 = (inp[12]) ? node18664 : node18661;
															assign node18661 = (inp[4]) ? 4'b1110 : 4'b1100;
															assign node18664 = (inp[4]) ? 4'b1100 : 4'b1111;
														assign node18667 = (inp[4]) ? node18671 : node18668;
															assign node18668 = (inp[12]) ? 4'b1110 : 4'b1100;
															assign node18671 = (inp[12]) ? 4'b1101 : 4'b1111;
												assign node18674 = (inp[1]) ? node18684 : node18675;
													assign node18675 = (inp[12]) ? node18681 : node18676;
														assign node18676 = (inp[4]) ? 4'b1111 : node18677;
															assign node18677 = (inp[11]) ? 4'b1100 : 4'b1101;
														assign node18681 = (inp[4]) ? 4'b1100 : 4'b1110;
													assign node18684 = (inp[4]) ? node18690 : node18685;
														assign node18685 = (inp[12]) ? 4'b1010 : node18686;
															assign node18686 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node18690 = (inp[12]) ? 4'b1000 : 4'b1010;
									assign node18693 = (inp[1]) ? node18807 : node18694;
										assign node18694 = (inp[2]) ? node18744 : node18695;
											assign node18695 = (inp[4]) ? node18719 : node18696;
												assign node18696 = (inp[12]) ? node18710 : node18697;
													assign node18697 = (inp[5]) ? node18705 : node18698;
														assign node18698 = (inp[15]) ? node18702 : node18699;
															assign node18699 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node18702 = (inp[11]) ? 4'b1100 : 4'b1101;
														assign node18705 = (inp[15]) ? 4'b1001 : node18706;
															assign node18706 = (inp[11]) ? 4'b1100 : 4'b1101;
													assign node18710 = (inp[15]) ? node18714 : node18711;
														assign node18711 = (inp[5]) ? 4'b1110 : 4'b1011;
														assign node18714 = (inp[5]) ? node18716 : 4'b1110;
															assign node18716 = (inp[11]) ? 4'b1010 : 4'b1011;
												assign node18719 = (inp[12]) ? node18731 : node18720;
													assign node18720 = (inp[5]) ? node18726 : node18721;
														assign node18721 = (inp[15]) ? 4'b1010 : node18722;
															assign node18722 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node18726 = (inp[15]) ? node18728 : 4'b1110;
															assign node18728 = (inp[11]) ? 4'b1010 : 4'b1011;
													assign node18731 = (inp[15]) ? node18737 : node18732;
														assign node18732 = (inp[11]) ? node18734 : 4'b1001;
															assign node18734 = (inp[5]) ? 4'b1001 : 4'b1000;
														assign node18737 = (inp[11]) ? node18741 : node18738;
															assign node18738 = (inp[5]) ? 4'b1000 : 4'b1100;
															assign node18741 = (inp[5]) ? 4'b1001 : 4'b1101;
											assign node18744 = (inp[4]) ? node18782 : node18745;
												assign node18745 = (inp[12]) ? node18769 : node18746;
													assign node18746 = (inp[11]) ? node18754 : node18747;
														assign node18747 = (inp[5]) ? node18751 : node18748;
															assign node18748 = (inp[15]) ? 4'b1000 : 4'b1100;
															assign node18751 = (inp[15]) ? 4'b1101 : 4'b1000;
														assign node18754 = (inp[9]) ? node18762 : node18755;
															assign node18755 = (inp[15]) ? node18759 : node18756;
																assign node18756 = (inp[5]) ? 4'b1000 : 4'b1101;
																assign node18759 = (inp[5]) ? 4'b1101 : 4'b1000;
															assign node18762 = (inp[5]) ? node18766 : node18763;
																assign node18763 = (inp[15]) ? 4'b1000 : 4'b1101;
																assign node18766 = (inp[15]) ? 4'b1101 : 4'b1000;
													assign node18769 = (inp[15]) ? node18775 : node18770;
														assign node18770 = (inp[5]) ? node18772 : 4'b1111;
															assign node18772 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node18775 = (inp[5]) ? node18779 : node18776;
															assign node18776 = (inp[11]) ? 4'b1011 : 4'b1010;
															assign node18779 = (inp[11]) ? 4'b1110 : 4'b1111;
												assign node18782 = (inp[12]) ? node18796 : node18783;
													assign node18783 = (inp[5]) ? node18789 : node18784;
														assign node18784 = (inp[15]) ? 4'b1111 : node18785;
															assign node18785 = (inp[11]) ? 4'b1110 : 4'b1111;
														assign node18789 = (inp[15]) ? node18793 : node18790;
															assign node18790 = (inp[11]) ? 4'b1010 : 4'b1011;
															assign node18793 = (inp[11]) ? 4'b1111 : 4'b1110;
													assign node18796 = (inp[15]) ? node18802 : node18797;
														assign node18797 = (inp[11]) ? node18799 : 4'b1100;
															assign node18799 = (inp[5]) ? 4'b1100 : 4'b1101;
														assign node18802 = (inp[5]) ? node18804 : 4'b1000;
															assign node18804 = (inp[11]) ? 4'b1100 : 4'b1101;
										assign node18807 = (inp[2]) ? node18867 : node18808;
											assign node18808 = (inp[11]) ? node18836 : node18809;
												assign node18809 = (inp[4]) ? node18825 : node18810;
													assign node18810 = (inp[12]) ? node18818 : node18811;
														assign node18811 = (inp[5]) ? node18815 : node18812;
															assign node18812 = (inp[15]) ? 4'b1000 : 4'b1100;
															assign node18815 = (inp[15]) ? 4'b1101 : 4'b1000;
														assign node18818 = (inp[5]) ? node18822 : node18819;
															assign node18819 = (inp[15]) ? 4'b1010 : 4'b1110;
															assign node18822 = (inp[15]) ? 4'b1111 : 4'b1011;
													assign node18825 = (inp[12]) ? node18831 : node18826;
														assign node18826 = (inp[5]) ? node18828 : 4'b1110;
															assign node18828 = (inp[15]) ? 4'b1110 : 4'b1010;
														assign node18831 = (inp[5]) ? 4'b1100 : node18832;
															assign node18832 = (inp[15]) ? 4'b1000 : 4'b1100;
												assign node18836 = (inp[5]) ? node18852 : node18837;
													assign node18837 = (inp[15]) ? node18845 : node18838;
														assign node18838 = (inp[4]) ? node18842 : node18839;
															assign node18839 = (inp[12]) ? 4'b1110 : 4'b1101;
															assign node18842 = (inp[12]) ? 4'b1101 : 4'b1111;
														assign node18845 = (inp[12]) ? node18849 : node18846;
															assign node18846 = (inp[4]) ? 4'b1111 : 4'b1001;
															assign node18849 = (inp[4]) ? 4'b1001 : 4'b1010;
													assign node18852 = (inp[15]) ? node18860 : node18853;
														assign node18853 = (inp[4]) ? node18857 : node18854;
															assign node18854 = (inp[12]) ? 4'b1010 : 4'b1000;
															assign node18857 = (inp[12]) ? 4'b1100 : 4'b1011;
														assign node18860 = (inp[4]) ? node18864 : node18861;
															assign node18861 = (inp[12]) ? 4'b1111 : 4'b1100;
															assign node18864 = (inp[12]) ? 4'b1100 : 4'b1110;
											assign node18867 = (inp[11]) ? node18899 : node18868;
												assign node18868 = (inp[5]) ? node18884 : node18869;
													assign node18869 = (inp[15]) ? node18877 : node18870;
														assign node18870 = (inp[4]) ? node18874 : node18871;
															assign node18871 = (inp[12]) ? 4'b1010 : 4'b1001;
															assign node18874 = (inp[12]) ? 4'b1000 : 4'b1010;
														assign node18877 = (inp[12]) ? node18881 : node18878;
															assign node18878 = (inp[4]) ? 4'b1010 : 4'b1100;
															assign node18881 = (inp[4]) ? 4'b1101 : 4'b1110;
													assign node18884 = (inp[15]) ? node18892 : node18885;
														assign node18885 = (inp[4]) ? node18889 : node18886;
															assign node18886 = (inp[12]) ? 4'b1111 : 4'b1100;
															assign node18889 = (inp[12]) ? 4'b1001 : 4'b1111;
														assign node18892 = (inp[12]) ? node18896 : node18893;
															assign node18893 = (inp[4]) ? 4'b1011 : 4'b1000;
															assign node18896 = (inp[4]) ? 4'b1001 : 4'b1011;
												assign node18899 = (inp[4]) ? node18915 : node18900;
													assign node18900 = (inp[12]) ? node18908 : node18901;
														assign node18901 = (inp[5]) ? node18905 : node18902;
															assign node18902 = (inp[15]) ? 4'b1101 : 4'b1001;
															assign node18905 = (inp[15]) ? 4'b1000 : 4'b1100;
														assign node18908 = (inp[5]) ? node18912 : node18909;
															assign node18909 = (inp[15]) ? 4'b1110 : 4'b1011;
															assign node18912 = (inp[15]) ? 4'b1010 : 4'b1110;
													assign node18915 = (inp[12]) ? node18921 : node18916;
														assign node18916 = (inp[15]) ? 4'b1010 : node18917;
															assign node18917 = (inp[5]) ? 4'b1110 : 4'b1010;
														assign node18921 = (inp[15]) ? node18923 : 4'b1000;
															assign node18923 = (inp[5]) ? 4'b1000 : 4'b1100;
							assign node18926 = (inp[7]) ? node19212 : node18927;
								assign node18927 = (inp[13]) ? node19047 : node18928;
									assign node18928 = (inp[1]) ? node18972 : node18929;
										assign node18929 = (inp[2]) ? node18951 : node18930;
											assign node18930 = (inp[4]) ? node18934 : node18931;
												assign node18931 = (inp[12]) ? 4'b1011 : 4'b1001;
												assign node18934 = (inp[12]) ? node18944 : node18935;
													assign node18935 = (inp[5]) ? node18937 : 4'b1011;
														assign node18937 = (inp[15]) ? node18941 : node18938;
															assign node18938 = (inp[11]) ? 4'b1010 : 4'b1011;
															assign node18941 = (inp[11]) ? 4'b1110 : 4'b1111;
													assign node18944 = (inp[5]) ? 4'b1000 : node18945;
														assign node18945 = (inp[15]) ? node18947 : 4'b1101;
															assign node18947 = (inp[11]) ? 4'b1000 : 4'b1001;
											assign node18951 = (inp[4]) ? node18955 : node18952;
												assign node18952 = (inp[12]) ? 4'b1111 : 4'b1101;
												assign node18955 = (inp[12]) ? node18963 : node18956;
													assign node18956 = (inp[5]) ? node18958 : 4'b1110;
														assign node18958 = (inp[15]) ? 4'b1011 : node18959;
															assign node18959 = (inp[11]) ? 4'b1111 : 4'b1110;
													assign node18963 = (inp[5]) ? 4'b1101 : node18964;
														assign node18964 = (inp[15]) ? node18968 : node18965;
															assign node18965 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node18968 = (inp[11]) ? 4'b1101 : 4'b1100;
										assign node18972 = (inp[2]) ? node19010 : node18973;
											assign node18973 = (inp[4]) ? node18985 : node18974;
												assign node18974 = (inp[12]) ? node18980 : node18975;
													assign node18975 = (inp[15]) ? node18977 : 4'b1101;
														assign node18977 = (inp[11]) ? 4'b1100 : 4'b1101;
													assign node18980 = (inp[11]) ? node18982 : 4'b1110;
														assign node18982 = (inp[15]) ? 4'b1111 : 4'b1110;
												assign node18985 = (inp[12]) ? node18999 : node18986;
													assign node18986 = (inp[5]) ? node18992 : node18987;
														assign node18987 = (inp[15]) ? node18989 : 4'b1111;
															assign node18989 = (inp[11]) ? 4'b1110 : 4'b1111;
														assign node18992 = (inp[15]) ? node18996 : node18993;
															assign node18993 = (inp[11]) ? 4'b1110 : 4'b1111;
															assign node18996 = (inp[11]) ? 4'b1011 : 4'b1010;
													assign node18999 = (inp[5]) ? node19005 : node19000;
														assign node19000 = (inp[15]) ? 4'b1101 : node19001;
															assign node19001 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node19005 = (inp[11]) ? node19007 : 4'b1101;
															assign node19007 = (inp[15]) ? 4'b1100 : 4'b1101;
											assign node19010 = (inp[4]) ? node19022 : node19011;
												assign node19011 = (inp[12]) ? node19017 : node19012;
													assign node19012 = (inp[11]) ? 4'b1000 : node19013;
														assign node19013 = (inp[15]) ? 4'b1000 : 4'b1001;
													assign node19017 = (inp[15]) ? 4'b1011 : node19018;
														assign node19018 = (inp[11]) ? 4'b1011 : 4'b1010;
												assign node19022 = (inp[12]) ? node19034 : node19023;
													assign node19023 = (inp[5]) ? node19029 : node19024;
														assign node19024 = (inp[15]) ? 4'b1011 : node19025;
															assign node19025 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node19029 = (inp[15]) ? node19031 : 4'b1011;
															assign node19031 = (inp[11]) ? 4'b1110 : 4'b1111;
													assign node19034 = (inp[5]) ? node19042 : node19035;
														assign node19035 = (inp[15]) ? node19039 : node19036;
															assign node19036 = (inp[11]) ? 4'b1100 : 4'b1101;
															assign node19039 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node19042 = (inp[11]) ? 4'b1001 : node19043;
															assign node19043 = (inp[15]) ? 4'b1001 : 4'b1000;
									assign node19047 = (inp[4]) ? node19117 : node19048;
										assign node19048 = (inp[12]) ? node19088 : node19049;
											assign node19049 = (inp[15]) ? node19073 : node19050;
												assign node19050 = (inp[11]) ? node19058 : node19051;
													assign node19051 = (inp[1]) ? node19055 : node19052;
														assign node19052 = (inp[2]) ? 4'b1101 : 4'b1001;
														assign node19055 = (inp[2]) ? 4'b1000 : 4'b1101;
													assign node19058 = (inp[5]) ? node19066 : node19059;
														assign node19059 = (inp[2]) ? node19063 : node19060;
															assign node19060 = (inp[1]) ? 4'b1100 : 4'b1000;
															assign node19063 = (inp[1]) ? 4'b1000 : 4'b1100;
														assign node19066 = (inp[1]) ? node19070 : node19067;
															assign node19067 = (inp[2]) ? 4'b1100 : 4'b1000;
															assign node19070 = (inp[2]) ? 4'b1000 : 4'b1100;
												assign node19073 = (inp[11]) ? node19081 : node19074;
													assign node19074 = (inp[1]) ? node19078 : node19075;
														assign node19075 = (inp[2]) ? 4'b1100 : 4'b1000;
														assign node19078 = (inp[2]) ? 4'b1001 : 4'b1101;
													assign node19081 = (inp[2]) ? node19085 : node19082;
														assign node19082 = (inp[1]) ? 4'b1101 : 4'b1001;
														assign node19085 = (inp[1]) ? 4'b1000 : 4'b1101;
											assign node19088 = (inp[15]) ? node19102 : node19089;
												assign node19089 = (inp[1]) ? node19097 : node19090;
													assign node19090 = (inp[11]) ? node19094 : node19091;
														assign node19091 = (inp[2]) ? 4'b1111 : 4'b1011;
														assign node19094 = (inp[2]) ? 4'b1110 : 4'b1010;
													assign node19097 = (inp[2]) ? 4'b1011 : node19098;
														assign node19098 = (inp[11]) ? 4'b1111 : 4'b1110;
												assign node19102 = (inp[11]) ? node19110 : node19103;
													assign node19103 = (inp[1]) ? node19107 : node19104;
														assign node19104 = (inp[2]) ? 4'b1110 : 4'b1010;
														assign node19107 = (inp[2]) ? 4'b1010 : 4'b1110;
													assign node19110 = (inp[2]) ? node19114 : node19111;
														assign node19111 = (inp[1]) ? 4'b1110 : 4'b1011;
														assign node19114 = (inp[1]) ? 4'b1011 : 4'b1111;
										assign node19117 = (inp[12]) ? node19159 : node19118;
											assign node19118 = (inp[2]) ? node19138 : node19119;
												assign node19119 = (inp[1]) ? node19131 : node19120;
													assign node19120 = (inp[15]) ? node19126 : node19121;
														assign node19121 = (inp[5]) ? 4'b1010 : node19122;
															assign node19122 = (inp[9]) ? 4'b1011 : 4'b1010;
														assign node19126 = (inp[5]) ? 4'b1111 : node19127;
															assign node19127 = (inp[11]) ? 4'b1011 : 4'b1010;
													assign node19131 = (inp[5]) ? node19135 : node19132;
														assign node19132 = (inp[11]) ? 4'b1110 : 4'b1111;
														assign node19135 = (inp[15]) ? 4'b1010 : 4'b1110;
												assign node19138 = (inp[1]) ? node19148 : node19139;
													assign node19139 = (inp[15]) ? node19141 : 4'b1111;
														assign node19141 = (inp[5]) ? node19145 : node19142;
															assign node19142 = (inp[11]) ? 4'b1110 : 4'b1111;
															assign node19145 = (inp[11]) ? 4'b1011 : 4'b1010;
													assign node19148 = (inp[5]) ? node19154 : node19149;
														assign node19149 = (inp[11]) ? 4'b1011 : node19150;
															assign node19150 = (inp[15]) ? 4'b1010 : 4'b1011;
														assign node19154 = (inp[15]) ? 4'b1111 : node19155;
															assign node19155 = (inp[11]) ? 4'b1010 : 4'b1011;
											assign node19159 = (inp[2]) ? node19191 : node19160;
												assign node19160 = (inp[1]) ? node19182 : node19161;
													assign node19161 = (inp[5]) ? node19167 : node19162;
														assign node19162 = (inp[15]) ? 4'b1001 : node19163;
															assign node19163 = (inp[11]) ? 4'b1100 : 4'b1101;
														assign node19167 = (inp[9]) ? node19175 : node19168;
															assign node19168 = (inp[15]) ? node19172 : node19169;
																assign node19169 = (inp[11]) ? 4'b1001 : 4'b1000;
																assign node19172 = (inp[11]) ? 4'b1000 : 4'b1001;
															assign node19175 = (inp[11]) ? node19179 : node19176;
																assign node19176 = (inp[15]) ? 4'b1001 : 4'b1000;
																assign node19179 = (inp[15]) ? 4'b1000 : 4'b1001;
													assign node19182 = (inp[15]) ? node19186 : node19183;
														assign node19183 = (inp[5]) ? 4'b1101 : 4'b1001;
														assign node19186 = (inp[5]) ? 4'b1101 : node19187;
															assign node19187 = (inp[11]) ? 4'b1101 : 4'b1100;
												assign node19191 = (inp[1]) ? node19203 : node19192;
													assign node19192 = (inp[15]) ? node19198 : node19193;
														assign node19193 = (inp[5]) ? node19195 : 4'b1001;
															assign node19195 = (inp[11]) ? 4'b1100 : 4'b1101;
														assign node19198 = (inp[11]) ? node19200 : 4'b1100;
															assign node19200 = (inp[5]) ? 4'b1101 : 4'b1100;
													assign node19203 = (inp[5]) ? node19207 : node19204;
														assign node19204 = (inp[15]) ? 4'b1000 : 4'b1100;
														assign node19207 = (inp[15]) ? node19209 : 4'b1001;
															assign node19209 = (inp[11]) ? 4'b1001 : 4'b1000;
								assign node19212 = (inp[1]) ? node19404 : node19213;
									assign node19213 = (inp[2]) ? node19309 : node19214;
										assign node19214 = (inp[4]) ? node19258 : node19215;
											assign node19215 = (inp[12]) ? node19235 : node19216;
												assign node19216 = (inp[5]) ? node19228 : node19217;
													assign node19217 = (inp[15]) ? node19223 : node19218;
														assign node19218 = (inp[13]) ? node19220 : 4'b1001;
															assign node19220 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node19223 = (inp[11]) ? 4'b1101 : node19224;
															assign node19224 = (inp[13]) ? 4'b1100 : 4'b1101;
													assign node19228 = (inp[15]) ? node19230 : 4'b1100;
														assign node19230 = (inp[11]) ? node19232 : 4'b1000;
															assign node19232 = (inp[13]) ? 4'b1000 : 4'b1001;
												assign node19235 = (inp[5]) ? node19247 : node19236;
													assign node19236 = (inp[15]) ? node19242 : node19237;
														assign node19237 = (inp[11]) ? 4'b1010 : node19238;
															assign node19238 = (inp[13]) ? 4'b1010 : 4'b1011;
														assign node19242 = (inp[11]) ? node19244 : 4'b1111;
															assign node19244 = (inp[13]) ? 4'b1111 : 4'b1110;
													assign node19247 = (inp[15]) ? node19253 : node19248;
														assign node19248 = (inp[11]) ? 4'b1111 : node19249;
															assign node19249 = (inp[13]) ? 4'b1111 : 4'b1110;
														assign node19253 = (inp[13]) ? node19255 : 4'b1011;
															assign node19255 = (inp[11]) ? 4'b1011 : 4'b1010;
											assign node19258 = (inp[12]) ? node19288 : node19259;
												assign node19259 = (inp[5]) ? node19277 : node19260;
													assign node19260 = (inp[11]) ? node19262 : 4'b1011;
														assign node19262 = (inp[9]) ? node19270 : node19263;
															assign node19263 = (inp[15]) ? node19267 : node19264;
																assign node19264 = (inp[13]) ? 4'b1010 : 4'b1011;
																assign node19267 = (inp[13]) ? 4'b1011 : 4'b1010;
															assign node19270 = (inp[15]) ? node19274 : node19271;
																assign node19271 = (inp[13]) ? 4'b1010 : 4'b1011;
																assign node19274 = (inp[13]) ? 4'b1011 : 4'b1010;
													assign node19277 = (inp[15]) ? node19283 : node19278;
														assign node19278 = (inp[13]) ? 4'b1111 : node19279;
															assign node19279 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node19283 = (inp[13]) ? node19285 : 4'b1011;
															assign node19285 = (inp[11]) ? 4'b1011 : 4'b1010;
												assign node19288 = (inp[5]) ? node19300 : node19289;
													assign node19289 = (inp[15]) ? node19295 : node19290;
														assign node19290 = (inp[11]) ? node19292 : 4'b1000;
															assign node19292 = (inp[13]) ? 4'b1001 : 4'b1000;
														assign node19295 = (inp[11]) ? 4'b1100 : node19296;
															assign node19296 = (inp[13]) ? 4'b1101 : 4'b1100;
													assign node19300 = (inp[11]) ? 4'b1000 : node19301;
														assign node19301 = (inp[15]) ? node19305 : node19302;
															assign node19302 = (inp[13]) ? 4'b1000 : 4'b1001;
															assign node19305 = (inp[13]) ? 4'b1001 : 4'b1000;
										assign node19309 = (inp[4]) ? node19357 : node19310;
											assign node19310 = (inp[12]) ? node19334 : node19311;
												assign node19311 = (inp[15]) ? node19323 : node19312;
													assign node19312 = (inp[5]) ? node19318 : node19313;
														assign node19313 = (inp[13]) ? node19315 : 4'b1101;
															assign node19315 = (inp[11]) ? 4'b1100 : 4'b1101;
														assign node19318 = (inp[11]) ? 4'b1001 : node19319;
															assign node19319 = (inp[13]) ? 4'b1001 : 4'b1000;
													assign node19323 = (inp[5]) ? node19329 : node19324;
														assign node19324 = (inp[13]) ? 4'b1001 : node19325;
															assign node19325 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node19329 = (inp[13]) ? 4'b1100 : node19330;
															assign node19330 = (inp[11]) ? 4'b1101 : 4'b1100;
												assign node19334 = (inp[5]) ? node19346 : node19335;
													assign node19335 = (inp[15]) ? node19341 : node19336;
														assign node19336 = (inp[11]) ? 4'b1110 : node19337;
															assign node19337 = (inp[13]) ? 4'b1110 : 4'b1111;
														assign node19341 = (inp[13]) ? node19343 : 4'b1010;
															assign node19343 = (inp[11]) ? 4'b1010 : 4'b1011;
													assign node19346 = (inp[15]) ? node19352 : node19347;
														assign node19347 = (inp[13]) ? node19349 : 4'b1011;
															assign node19349 = (inp[11]) ? 4'b1010 : 4'b1011;
														assign node19352 = (inp[13]) ? node19354 : 4'b1111;
															assign node19354 = (inp[11]) ? 4'b1111 : 4'b1110;
											assign node19357 = (inp[12]) ? node19385 : node19358;
												assign node19358 = (inp[5]) ? node19374 : node19359;
													assign node19359 = (inp[11]) ? node19361 : 4'b1110;
														assign node19361 = (inp[9]) ? node19369 : node19362;
															assign node19362 = (inp[15]) ? node19366 : node19363;
																assign node19363 = (inp[13]) ? 4'b1111 : 4'b1110;
																assign node19366 = (inp[13]) ? 4'b1110 : 4'b1111;
															assign node19369 = (inp[15]) ? 4'b1111 : node19370;
																assign node19370 = (inp[13]) ? 4'b1111 : 4'b1110;
													assign node19374 = (inp[15]) ? node19380 : node19375;
														assign node19375 = (inp[11]) ? node19377 : 4'b1010;
															assign node19377 = (inp[13]) ? 4'b1011 : 4'b1010;
														assign node19380 = (inp[13]) ? node19382 : 4'b1110;
															assign node19382 = (inp[11]) ? 4'b1110 : 4'b1111;
												assign node19385 = (inp[15]) ? node19393 : node19386;
													assign node19386 = (inp[13]) ? node19388 : 4'b1101;
														assign node19388 = (inp[11]) ? node19390 : 4'b1101;
															assign node19390 = (inp[5]) ? 4'b1101 : 4'b1100;
													assign node19393 = (inp[5]) ? node19399 : node19394;
														assign node19394 = (inp[13]) ? 4'b1001 : node19395;
															assign node19395 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node19399 = (inp[13]) ? node19401 : 4'b1101;
															assign node19401 = (inp[11]) ? 4'b1101 : 4'b1100;
									assign node19404 = (inp[2]) ? node19498 : node19405;
										assign node19405 = (inp[4]) ? node19451 : node19406;
											assign node19406 = (inp[12]) ? node19430 : node19407;
												assign node19407 = (inp[5]) ? node19419 : node19408;
													assign node19408 = (inp[15]) ? node19414 : node19409;
														assign node19409 = (inp[11]) ? node19411 : 4'b1101;
															assign node19411 = (inp[13]) ? 4'b1100 : 4'b1101;
														assign node19414 = (inp[11]) ? 4'b1000 : node19415;
															assign node19415 = (inp[13]) ? 4'b1001 : 4'b1000;
													assign node19419 = (inp[15]) ? node19425 : node19420;
														assign node19420 = (inp[11]) ? 4'b1001 : node19421;
															assign node19421 = (inp[13]) ? 4'b1001 : 4'b1000;
														assign node19425 = (inp[13]) ? node19427 : 4'b1101;
															assign node19427 = (inp[11]) ? 4'b1101 : 4'b1100;
												assign node19430 = (inp[5]) ? node19442 : node19431;
													assign node19431 = (inp[15]) ? node19437 : node19432;
														assign node19432 = (inp[13]) ? 4'b1111 : node19433;
															assign node19433 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node19437 = (inp[11]) ? node19439 : 4'b1011;
															assign node19439 = (inp[13]) ? 4'b1011 : 4'b1010;
													assign node19442 = (inp[15]) ? node19446 : node19443;
														assign node19443 = (inp[13]) ? 4'b1011 : 4'b1010;
														assign node19446 = (inp[13]) ? 4'b1110 : node19447;
															assign node19447 = (inp[11]) ? 4'b1111 : 4'b1110;
											assign node19451 = (inp[12]) ? node19475 : node19452;
												assign node19452 = (inp[11]) ? node19462 : node19453;
													assign node19453 = (inp[15]) ? node19457 : node19454;
														assign node19454 = (inp[5]) ? 4'b1011 : 4'b1111;
														assign node19457 = (inp[5]) ? 4'b1111 : node19458;
															assign node19458 = (inp[13]) ? 4'b1111 : 4'b1110;
													assign node19462 = (inp[15]) ? node19470 : node19463;
														assign node19463 = (inp[5]) ? node19467 : node19464;
															assign node19464 = (inp[13]) ? 4'b1110 : 4'b1111;
															assign node19467 = (inp[13]) ? 4'b1010 : 4'b1011;
														assign node19470 = (inp[5]) ? node19472 : 4'b1110;
															assign node19472 = (inp[13]) ? 4'b1111 : 4'b1110;
												assign node19475 = (inp[15]) ? node19487 : node19476;
													assign node19476 = (inp[5]) ? node19482 : node19477;
														assign node19477 = (inp[11]) ? node19479 : 4'b1101;
															assign node19479 = (inp[13]) ? 4'b1100 : 4'b1101;
														assign node19482 = (inp[11]) ? 4'b1101 : node19483;
															assign node19483 = (inp[13]) ? 4'b1101 : 4'b1100;
													assign node19487 = (inp[5]) ? node19493 : node19488;
														assign node19488 = (inp[11]) ? 4'b1000 : node19489;
															assign node19489 = (inp[13]) ? 4'b1001 : 4'b1000;
														assign node19493 = (inp[13]) ? 4'b1101 : node19494;
															assign node19494 = (inp[11]) ? 4'b1100 : 4'b1101;
										assign node19498 = (inp[15]) ? node19540 : node19499;
											assign node19499 = (inp[5]) ? node19521 : node19500;
												assign node19500 = (inp[12]) ? node19510 : node19501;
													assign node19501 = (inp[4]) ? node19507 : node19502;
														assign node19502 = (inp[11]) ? 4'b1000 : node19503;
															assign node19503 = (inp[13]) ? 4'b1000 : 4'b1001;
														assign node19507 = (inp[13]) ? 4'b1011 : 4'b1010;
													assign node19510 = (inp[4]) ? node19516 : node19511;
														assign node19511 = (inp[13]) ? node19513 : 4'b1011;
															assign node19513 = (inp[11]) ? 4'b1010 : 4'b1011;
														assign node19516 = (inp[9]) ? 4'b1001 : node19517;
															assign node19517 = (inp[13]) ? 4'b1001 : 4'b1000;
												assign node19521 = (inp[12]) ? node19533 : node19522;
													assign node19522 = (inp[4]) ? node19528 : node19523;
														assign node19523 = (inp[11]) ? 4'b1101 : node19524;
															assign node19524 = (inp[13]) ? 4'b1101 : 4'b1100;
														assign node19528 = (inp[13]) ? node19530 : 4'b1110;
															assign node19530 = (inp[11]) ? 4'b1111 : 4'b1110;
													assign node19533 = (inp[4]) ? 4'b1000 : node19534;
														assign node19534 = (inp[13]) ? node19536 : 4'b1110;
															assign node19536 = (inp[11]) ? 4'b1111 : 4'b1110;
											assign node19540 = (inp[5]) ? node19564 : node19541;
												assign node19541 = (inp[12]) ? node19553 : node19542;
													assign node19542 = (inp[4]) ? node19548 : node19543;
														assign node19543 = (inp[11]) ? 4'b1100 : node19544;
															assign node19544 = (inp[13]) ? 4'b1101 : 4'b1100;
														assign node19548 = (inp[13]) ? 4'b1011 : node19549;
															assign node19549 = (inp[11]) ? 4'b1010 : 4'b1011;
													assign node19553 = (inp[4]) ? node19559 : node19554;
														assign node19554 = (inp[13]) ? 4'b1111 : node19555;
															assign node19555 = (inp[11]) ? 4'b1110 : 4'b1111;
														assign node19559 = (inp[13]) ? node19561 : 4'b1101;
															assign node19561 = (inp[11]) ? 4'b1101 : 4'b1100;
												assign node19564 = (inp[11]) ? node19578 : node19565;
													assign node19565 = (inp[13]) ? node19571 : node19566;
														assign node19566 = (inp[4]) ? 4'b1011 : node19567;
															assign node19567 = (inp[12]) ? 4'b1011 : 4'b1001;
														assign node19571 = (inp[12]) ? node19575 : node19572;
															assign node19572 = (inp[4]) ? 4'b1010 : 4'b1001;
															assign node19575 = (inp[4]) ? 4'b1000 : 4'b1010;
													assign node19578 = (inp[13]) ? node19586 : node19579;
														assign node19579 = (inp[12]) ? node19583 : node19580;
															assign node19580 = (inp[4]) ? 4'b1011 : 4'b1000;
															assign node19583 = (inp[4]) ? 4'b1001 : 4'b1011;
														assign node19586 = (inp[12]) ? node19590 : node19587;
															assign node19587 = (inp[4]) ? 4'b1011 : 4'b1001;
															assign node19590 = (inp[4]) ? 4'b1001 : 4'b1011;
						assign node19593 = (inp[0]) ? node20343 : node19594;
							assign node19594 = (inp[13]) ? node19918 : node19595;
								assign node19595 = (inp[7]) ? node19711 : node19596;
									assign node19596 = (inp[1]) ? node19638 : node19597;
										assign node19597 = (inp[2]) ? node19619 : node19598;
											assign node19598 = (inp[4]) ? node19602 : node19599;
												assign node19599 = (inp[12]) ? 4'b1011 : 4'b1001;
												assign node19602 = (inp[12]) ? node19612 : node19603;
													assign node19603 = (inp[5]) ? node19605 : 4'b1011;
														assign node19605 = (inp[15]) ? node19609 : node19606;
															assign node19606 = (inp[11]) ? 4'b1010 : 4'b1011;
															assign node19609 = (inp[11]) ? 4'b1110 : 4'b1111;
													assign node19612 = (inp[5]) ? 4'b1000 : node19613;
														assign node19613 = (inp[15]) ? node19615 : 4'b1101;
															assign node19615 = (inp[11]) ? 4'b1000 : 4'b1001;
											assign node19619 = (inp[4]) ? node19623 : node19620;
												assign node19620 = (inp[12]) ? 4'b1111 : 4'b1101;
												assign node19623 = (inp[12]) ? node19631 : node19624;
													assign node19624 = (inp[5]) ? node19626 : 4'b1110;
														assign node19626 = (inp[15]) ? 4'b1011 : node19627;
															assign node19627 = (inp[11]) ? 4'b1111 : 4'b1110;
													assign node19631 = (inp[5]) ? 4'b1101 : node19632;
														assign node19632 = (inp[11]) ? 4'b1001 : node19633;
															assign node19633 = (inp[15]) ? 4'b1100 : 4'b1000;
										assign node19638 = (inp[2]) ? node19676 : node19639;
											assign node19639 = (inp[4]) ? node19651 : node19640;
												assign node19640 = (inp[12]) ? node19646 : node19641;
													assign node19641 = (inp[11]) ? node19643 : 4'b1101;
														assign node19643 = (inp[15]) ? 4'b1100 : 4'b1101;
													assign node19646 = (inp[15]) ? node19648 : 4'b1110;
														assign node19648 = (inp[11]) ? 4'b1111 : 4'b1110;
												assign node19651 = (inp[12]) ? node19665 : node19652;
													assign node19652 = (inp[5]) ? node19658 : node19653;
														assign node19653 = (inp[11]) ? node19655 : 4'b1111;
															assign node19655 = (inp[15]) ? 4'b1110 : 4'b1111;
														assign node19658 = (inp[15]) ? node19662 : node19659;
															assign node19659 = (inp[11]) ? 4'b1110 : 4'b1111;
															assign node19662 = (inp[11]) ? 4'b1011 : 4'b1010;
													assign node19665 = (inp[15]) ? node19671 : node19666;
														assign node19666 = (inp[5]) ? 4'b1101 : node19667;
															assign node19667 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node19671 = (inp[5]) ? node19673 : 4'b1101;
															assign node19673 = (inp[11]) ? 4'b1100 : 4'b1101;
											assign node19676 = (inp[4]) ? node19688 : node19677;
												assign node19677 = (inp[12]) ? node19683 : node19678;
													assign node19678 = (inp[11]) ? 4'b1000 : node19679;
														assign node19679 = (inp[15]) ? 4'b1000 : 4'b1001;
													assign node19683 = (inp[11]) ? 4'b1011 : node19684;
														assign node19684 = (inp[15]) ? 4'b1011 : 4'b1010;
												assign node19688 = (inp[12]) ? node19698 : node19689;
													assign node19689 = (inp[5]) ? node19695 : node19690;
														assign node19690 = (inp[15]) ? 4'b1011 : node19691;
															assign node19691 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node19695 = (inp[15]) ? 4'b1111 : 4'b1011;
													assign node19698 = (inp[5]) ? node19706 : node19699;
														assign node19699 = (inp[15]) ? node19703 : node19700;
															assign node19700 = (inp[11]) ? 4'b1100 : 4'b1101;
															assign node19703 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node19706 = (inp[11]) ? 4'b1001 : node19707;
															assign node19707 = (inp[15]) ? 4'b1001 : 4'b1000;
									assign node19711 = (inp[4]) ? node19831 : node19712;
										assign node19712 = (inp[12]) ? node19778 : node19713;
											assign node19713 = (inp[15]) ? node19745 : node19714;
												assign node19714 = (inp[5]) ? node19724 : node19715;
													assign node19715 = (inp[2]) ? node19719 : node19716;
														assign node19716 = (inp[1]) ? 4'b1101 : 4'b1001;
														assign node19719 = (inp[1]) ? node19721 : 4'b1101;
															assign node19721 = (inp[11]) ? 4'b1000 : 4'b1001;
													assign node19724 = (inp[11]) ? node19738 : node19725;
														assign node19725 = (inp[9]) ? node19731 : node19726;
															assign node19726 = (inp[2]) ? 4'b1100 : node19727;
																assign node19727 = (inp[1]) ? 4'b1000 : 4'b1100;
															assign node19731 = (inp[2]) ? node19735 : node19732;
																assign node19732 = (inp[1]) ? 4'b1000 : 4'b1100;
																assign node19735 = (inp[1]) ? 4'b1100 : 4'b1000;
														assign node19738 = (inp[1]) ? node19742 : node19739;
															assign node19739 = (inp[2]) ? 4'b1001 : 4'b1100;
															assign node19742 = (inp[2]) ? 4'b1101 : 4'b1001;
												assign node19745 = (inp[2]) ? node19755 : node19746;
													assign node19746 = (inp[1]) ? node19752 : node19747;
														assign node19747 = (inp[5]) ? node19749 : 4'b1101;
															assign node19749 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node19752 = (inp[5]) ? 4'b1101 : 4'b1000;
													assign node19755 = (inp[11]) ? node19771 : node19756;
														assign node19756 = (inp[9]) ? node19764 : node19757;
															assign node19757 = (inp[1]) ? node19761 : node19758;
																assign node19758 = (inp[5]) ? 4'b1100 : 4'b1001;
																assign node19761 = (inp[5]) ? 4'b1001 : 4'b1100;
															assign node19764 = (inp[5]) ? node19768 : node19765;
																assign node19765 = (inp[1]) ? 4'b1100 : 4'b1001;
																assign node19768 = (inp[1]) ? 4'b1001 : 4'b1100;
														assign node19771 = (inp[5]) ? node19775 : node19772;
															assign node19772 = (inp[1]) ? 4'b1100 : 4'b1000;
															assign node19775 = (inp[1]) ? 4'b1000 : 4'b1101;
											assign node19778 = (inp[15]) ? node19802 : node19779;
												assign node19779 = (inp[5]) ? node19793 : node19780;
													assign node19780 = (inp[2]) ? node19788 : node19781;
														assign node19781 = (inp[1]) ? node19785 : node19782;
															assign node19782 = (inp[11]) ? 4'b1010 : 4'b1011;
															assign node19785 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node19788 = (inp[1]) ? 4'b1011 : node19789;
															assign node19789 = (inp[11]) ? 4'b1110 : 4'b1111;
													assign node19793 = (inp[1]) ? node19799 : node19794;
														assign node19794 = (inp[2]) ? 4'b1011 : node19795;
															assign node19795 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node19799 = (inp[2]) ? 4'b1110 : 4'b1010;
												assign node19802 = (inp[5]) ? node19816 : node19803;
													assign node19803 = (inp[11]) ? node19811 : node19804;
														assign node19804 = (inp[2]) ? node19808 : node19805;
															assign node19805 = (inp[1]) ? 4'b1011 : 4'b1111;
															assign node19808 = (inp[1]) ? 4'b1111 : 4'b1010;
														assign node19811 = (inp[2]) ? 4'b1010 : node19812;
															assign node19812 = (inp[1]) ? 4'b1010 : 4'b1110;
													assign node19816 = (inp[11]) ? node19824 : node19817;
														assign node19817 = (inp[2]) ? node19821 : node19818;
															assign node19818 = (inp[1]) ? 4'b1110 : 4'b1011;
															assign node19821 = (inp[1]) ? 4'b1011 : 4'b1111;
														assign node19824 = (inp[1]) ? node19828 : node19825;
															assign node19825 = (inp[2]) ? 4'b1111 : 4'b1011;
															assign node19828 = (inp[2]) ? 4'b1011 : 4'b1111;
										assign node19831 = (inp[12]) ? node19875 : node19832;
											assign node19832 = (inp[2]) ? node19854 : node19833;
												assign node19833 = (inp[1]) ? node19845 : node19834;
													assign node19834 = (inp[15]) ? node19840 : node19835;
														assign node19835 = (inp[5]) ? node19837 : 4'b1011;
															assign node19837 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node19840 = (inp[11]) ? node19842 : 4'b1011;
															assign node19842 = (inp[5]) ? 4'b1011 : 4'b1010;
													assign node19845 = (inp[15]) ? node19849 : node19846;
														assign node19846 = (inp[5]) ? 4'b1011 : 4'b1111;
														assign node19849 = (inp[11]) ? 4'b1110 : node19850;
															assign node19850 = (inp[5]) ? 4'b1111 : 4'b1110;
												assign node19854 = (inp[1]) ? node19864 : node19855;
													assign node19855 = (inp[5]) ? node19861 : node19856;
														assign node19856 = (inp[11]) ? node19858 : 4'b1110;
															assign node19858 = (inp[15]) ? 4'b1111 : 4'b1110;
														assign node19861 = (inp[15]) ? 4'b1110 : 4'b1010;
													assign node19864 = (inp[15]) ? node19870 : node19865;
														assign node19865 = (inp[5]) ? 4'b1110 : node19866;
															assign node19866 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node19870 = (inp[5]) ? 4'b1011 : node19871;
															assign node19871 = (inp[11]) ? 4'b1010 : 4'b1011;
											assign node19875 = (inp[2]) ? node19897 : node19876;
												assign node19876 = (inp[1]) ? node19886 : node19877;
													assign node19877 = (inp[15]) ? node19883 : node19878;
														assign node19878 = (inp[11]) ? 4'b1000 : node19879;
															assign node19879 = (inp[5]) ? 4'b1001 : 4'b1000;
														assign node19883 = (inp[5]) ? 4'b1000 : 4'b1100;
													assign node19886 = (inp[15]) ? node19892 : node19887;
														assign node19887 = (inp[5]) ? node19889 : 4'b1101;
															assign node19889 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node19892 = (inp[5]) ? node19894 : 4'b1000;
															assign node19894 = (inp[11]) ? 4'b1100 : 4'b1101;
												assign node19897 = (inp[1]) ? node19909 : node19898;
													assign node19898 = (inp[5]) ? node19904 : node19899;
														assign node19899 = (inp[15]) ? node19901 : 4'b1101;
															assign node19901 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node19904 = (inp[11]) ? 4'b1101 : node19905;
															assign node19905 = (inp[15]) ? 4'b1101 : 4'b1100;
													assign node19909 = (inp[15]) ? node19915 : node19910;
														assign node19910 = (inp[5]) ? 4'b1000 : node19911;
															assign node19911 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node19915 = (inp[5]) ? 4'b1001 : 4'b1101;
								assign node19918 = (inp[1]) ? node20154 : node19919;
									assign node19919 = (inp[2]) ? node20019 : node19920;
										assign node19920 = (inp[7]) ? node19970 : node19921;
											assign node19921 = (inp[4]) ? node19945 : node19922;
												assign node19922 = (inp[12]) ? node19930 : node19923;
													assign node19923 = (inp[11]) ? node19927 : node19924;
														assign node19924 = (inp[15]) ? 4'b1000 : 4'b1001;
														assign node19927 = (inp[15]) ? 4'b1001 : 4'b1000;
													assign node19930 = (inp[9]) ? node19938 : node19931;
														assign node19931 = (inp[15]) ? node19935 : node19932;
															assign node19932 = (inp[11]) ? 4'b1010 : 4'b1011;
															assign node19935 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node19938 = (inp[15]) ? node19942 : node19939;
															assign node19939 = (inp[11]) ? 4'b1010 : 4'b1011;
															assign node19942 = (inp[11]) ? 4'b1011 : 4'b1010;
												assign node19945 = (inp[12]) ? node19957 : node19946;
													assign node19946 = (inp[15]) ? node19952 : node19947;
														assign node19947 = (inp[5]) ? 4'b1010 : node19948;
															assign node19948 = (inp[11]) ? 4'b1010 : 4'b1011;
														assign node19952 = (inp[5]) ? 4'b1111 : node19953;
															assign node19953 = (inp[11]) ? 4'b1011 : 4'b1010;
													assign node19957 = (inp[5]) ? node19963 : node19958;
														assign node19958 = (inp[15]) ? 4'b1001 : node19959;
															assign node19959 = (inp[11]) ? 4'b1100 : 4'b1101;
														assign node19963 = (inp[11]) ? node19967 : node19964;
															assign node19964 = (inp[15]) ? 4'b1001 : 4'b1000;
															assign node19967 = (inp[15]) ? 4'b1000 : 4'b1001;
											assign node19970 = (inp[4]) ? node19994 : node19971;
												assign node19971 = (inp[12]) ? node19985 : node19972;
													assign node19972 = (inp[5]) ? node19980 : node19973;
														assign node19973 = (inp[15]) ? node19977 : node19974;
															assign node19974 = (inp[11]) ? 4'b1000 : 4'b1001;
															assign node19977 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node19980 = (inp[15]) ? 4'b1000 : node19981;
															assign node19981 = (inp[11]) ? 4'b1101 : 4'b1100;
													assign node19985 = (inp[5]) ? node19989 : node19986;
														assign node19986 = (inp[15]) ? 4'b1111 : 4'b1010;
														assign node19989 = (inp[15]) ? node19991 : 4'b1111;
															assign node19991 = (inp[11]) ? 4'b1011 : 4'b1010;
												assign node19994 = (inp[12]) ? node20006 : node19995;
													assign node19995 = (inp[15]) ? node20001 : node19996;
														assign node19996 = (inp[5]) ? 4'b1111 : node19997;
															assign node19997 = (inp[11]) ? 4'b1010 : 4'b1011;
														assign node20001 = (inp[11]) ? 4'b1011 : node20002;
															assign node20002 = (inp[5]) ? 4'b1010 : 4'b1011;
													assign node20006 = (inp[5]) ? node20014 : node20007;
														assign node20007 = (inp[15]) ? node20011 : node20008;
															assign node20008 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node20011 = (inp[11]) ? 4'b1100 : 4'b1101;
														assign node20014 = (inp[11]) ? 4'b1000 : node20015;
															assign node20015 = (inp[15]) ? 4'b1001 : 4'b1000;
										assign node20019 = (inp[7]) ? node20099 : node20020;
											assign node20020 = (inp[4]) ? node20074 : node20021;
												assign node20021 = (inp[12]) ? node20043 : node20022;
													assign node20022 = (inp[9]) ? node20036 : node20023;
														assign node20023 = (inp[5]) ? node20031 : node20024;
															assign node20024 = (inp[15]) ? node20028 : node20025;
																assign node20025 = (inp[11]) ? 4'b1100 : 4'b1101;
																assign node20028 = (inp[11]) ? 4'b1101 : 4'b1100;
															assign node20031 = (inp[11]) ? 4'b1101 : node20032;
																assign node20032 = (inp[15]) ? 4'b1100 : 4'b1101;
														assign node20036 = (inp[15]) ? node20040 : node20037;
															assign node20037 = (inp[11]) ? 4'b1100 : 4'b1101;
															assign node20040 = (inp[11]) ? 4'b1101 : 4'b1100;
													assign node20043 = (inp[5]) ? node20059 : node20044;
														assign node20044 = (inp[9]) ? node20052 : node20045;
															assign node20045 = (inp[15]) ? node20049 : node20046;
																assign node20046 = (inp[11]) ? 4'b1110 : 4'b1111;
																assign node20049 = (inp[11]) ? 4'b1111 : 4'b1110;
															assign node20052 = (inp[11]) ? node20056 : node20053;
																assign node20053 = (inp[15]) ? 4'b1110 : 4'b1111;
																assign node20056 = (inp[15]) ? 4'b1111 : 4'b1110;
														assign node20059 = (inp[9]) ? node20067 : node20060;
															assign node20060 = (inp[15]) ? node20064 : node20061;
																assign node20061 = (inp[11]) ? 4'b1110 : 4'b1111;
																assign node20064 = (inp[11]) ? 4'b1111 : 4'b1110;
															assign node20067 = (inp[15]) ? node20071 : node20068;
																assign node20068 = (inp[11]) ? 4'b1110 : 4'b1111;
																assign node20071 = (inp[11]) ? 4'b1111 : 4'b1110;
												assign node20074 = (inp[12]) ? node20088 : node20075;
													assign node20075 = (inp[15]) ? node20081 : node20076;
														assign node20076 = (inp[5]) ? 4'b1111 : node20077;
															assign node20077 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node20081 = (inp[5]) ? node20085 : node20082;
															assign node20082 = (inp[11]) ? 4'b1110 : 4'b1111;
															assign node20085 = (inp[11]) ? 4'b1011 : 4'b1010;
													assign node20088 = (inp[15]) ? node20094 : node20089;
														assign node20089 = (inp[5]) ? node20091 : 4'b1001;
															assign node20091 = (inp[11]) ? 4'b1100 : 4'b1101;
														assign node20094 = (inp[11]) ? node20096 : 4'b1100;
															assign node20096 = (inp[5]) ? 4'b1101 : 4'b1100;
											assign node20099 = (inp[4]) ? node20129 : node20100;
												assign node20100 = (inp[12]) ? node20116 : node20101;
													assign node20101 = (inp[11]) ? node20109 : node20102;
														assign node20102 = (inp[15]) ? node20106 : node20103;
															assign node20103 = (inp[5]) ? 4'b1001 : 4'b1101;
															assign node20106 = (inp[5]) ? 4'b1100 : 4'b1001;
														assign node20109 = (inp[5]) ? node20113 : node20110;
															assign node20110 = (inp[15]) ? 4'b1001 : 4'b1100;
															assign node20113 = (inp[15]) ? 4'b1100 : 4'b1001;
													assign node20116 = (inp[15]) ? node20122 : node20117;
														assign node20117 = (inp[5]) ? node20119 : 4'b1110;
															assign node20119 = (inp[11]) ? 4'b1010 : 4'b1011;
														assign node20122 = (inp[5]) ? node20126 : node20123;
															assign node20123 = (inp[11]) ? 4'b1010 : 4'b1011;
															assign node20126 = (inp[11]) ? 4'b1111 : 4'b1110;
												assign node20129 = (inp[12]) ? node20143 : node20130;
													assign node20130 = (inp[15]) ? node20138 : node20131;
														assign node20131 = (inp[11]) ? node20135 : node20132;
															assign node20132 = (inp[5]) ? 4'b1010 : 4'b1110;
															assign node20135 = (inp[5]) ? 4'b1011 : 4'b1111;
														assign node20138 = (inp[5]) ? node20140 : 4'b1110;
															assign node20140 = (inp[11]) ? 4'b1110 : 4'b1111;
													assign node20143 = (inp[5]) ? node20149 : node20144;
														assign node20144 = (inp[15]) ? 4'b1001 : node20145;
															assign node20145 = (inp[11]) ? 4'b1100 : 4'b1101;
														assign node20149 = (inp[15]) ? node20151 : 4'b1101;
															assign node20151 = (inp[11]) ? 4'b1101 : 4'b1100;
									assign node20154 = (inp[2]) ? node20250 : node20155;
										assign node20155 = (inp[11]) ? node20199 : node20156;
											assign node20156 = (inp[7]) ? node20172 : node20157;
												assign node20157 = (inp[12]) ? node20165 : node20158;
													assign node20158 = (inp[4]) ? node20160 : 4'b1101;
														assign node20160 = (inp[5]) ? node20162 : 4'b1111;
															assign node20162 = (inp[15]) ? 4'b1010 : 4'b1110;
													assign node20165 = (inp[4]) ? node20167 : 4'b1110;
														assign node20167 = (inp[5]) ? 4'b1101 : node20168;
															assign node20168 = (inp[15]) ? 4'b1100 : 4'b1001;
												assign node20172 = (inp[4]) ? node20188 : node20173;
													assign node20173 = (inp[12]) ? node20181 : node20174;
														assign node20174 = (inp[15]) ? node20178 : node20175;
															assign node20175 = (inp[5]) ? 4'b1001 : 4'b1101;
															assign node20178 = (inp[5]) ? 4'b1100 : 4'b1001;
														assign node20181 = (inp[5]) ? node20185 : node20182;
															assign node20182 = (inp[15]) ? 4'b1011 : 4'b1111;
															assign node20185 = (inp[15]) ? 4'b1110 : 4'b1010;
													assign node20188 = (inp[12]) ? node20194 : node20189;
														assign node20189 = (inp[5]) ? node20191 : 4'b1111;
															assign node20191 = (inp[15]) ? 4'b1111 : 4'b1011;
														assign node20194 = (inp[5]) ? 4'b1101 : node20195;
															assign node20195 = (inp[15]) ? 4'b1001 : 4'b1101;
											assign node20199 = (inp[12]) ? node20225 : node20200;
												assign node20200 = (inp[4]) ? node20212 : node20201;
													assign node20201 = (inp[15]) ? node20207 : node20202;
														assign node20202 = (inp[7]) ? node20204 : 4'b1100;
															assign node20204 = (inp[5]) ? 4'b1001 : 4'b1100;
														assign node20207 = (inp[5]) ? 4'b1101 : node20208;
															assign node20208 = (inp[9]) ? 4'b1000 : 4'b1101;
													assign node20212 = (inp[15]) ? node20218 : node20213;
														assign node20213 = (inp[7]) ? node20215 : 4'b1110;
															assign node20215 = (inp[5]) ? 4'b1010 : 4'b1110;
														assign node20218 = (inp[7]) ? node20222 : node20219;
															assign node20219 = (inp[5]) ? 4'b1010 : 4'b1111;
															assign node20222 = (inp[5]) ? 4'b1111 : 4'b1110;
												assign node20225 = (inp[4]) ? node20237 : node20226;
													assign node20226 = (inp[15]) ? node20232 : node20227;
														assign node20227 = (inp[7]) ? node20229 : 4'b1111;
															assign node20229 = (inp[5]) ? 4'b1011 : 4'b1111;
														assign node20232 = (inp[5]) ? 4'b1110 : node20233;
															assign node20233 = (inp[7]) ? 4'b1011 : 4'b1110;
													assign node20237 = (inp[5]) ? node20245 : node20238;
														assign node20238 = (inp[7]) ? node20242 : node20239;
															assign node20239 = (inp[15]) ? 4'b1101 : 4'b1001;
															assign node20242 = (inp[15]) ? 4'b1000 : 4'b1100;
														assign node20245 = (inp[15]) ? 4'b1101 : node20246;
															assign node20246 = (inp[7]) ? 4'b1101 : 4'b1100;
										assign node20250 = (inp[7]) ? node20284 : node20251;
											assign node20251 = (inp[4]) ? node20263 : node20252;
												assign node20252 = (inp[12]) ? node20258 : node20253;
													assign node20253 = (inp[15]) ? node20255 : 4'b1000;
														assign node20255 = (inp[11]) ? 4'b1000 : 4'b1001;
													assign node20258 = (inp[11]) ? 4'b1011 : node20259;
														assign node20259 = (inp[15]) ? 4'b1010 : 4'b1011;
												assign node20263 = (inp[12]) ? node20275 : node20264;
													assign node20264 = (inp[15]) ? node20270 : node20265;
														assign node20265 = (inp[5]) ? node20267 : 4'b1011;
															assign node20267 = (inp[11]) ? 4'b1010 : 4'b1011;
														assign node20270 = (inp[5]) ? 4'b1111 : node20271;
															assign node20271 = (inp[11]) ? 4'b1011 : 4'b1010;
													assign node20275 = (inp[5]) ? node20279 : node20276;
														assign node20276 = (inp[15]) ? 4'b1000 : 4'b1100;
														assign node20279 = (inp[15]) ? node20281 : 4'b1001;
															assign node20281 = (inp[11]) ? 4'b1001 : 4'b1000;
											assign node20284 = (inp[11]) ? node20316 : node20285;
												assign node20285 = (inp[5]) ? node20301 : node20286;
													assign node20286 = (inp[15]) ? node20294 : node20287;
														assign node20287 = (inp[12]) ? node20291 : node20288;
															assign node20288 = (inp[4]) ? 4'b1011 : 4'b1000;
															assign node20291 = (inp[4]) ? 4'b1001 : 4'b1011;
														assign node20294 = (inp[12]) ? node20298 : node20295;
															assign node20295 = (inp[4]) ? 4'b1011 : 4'b1101;
															assign node20298 = (inp[4]) ? 4'b1100 : 4'b1111;
													assign node20301 = (inp[15]) ? node20309 : node20302;
														assign node20302 = (inp[4]) ? node20306 : node20303;
															assign node20303 = (inp[12]) ? 4'b1110 : 4'b1101;
															assign node20306 = (inp[12]) ? 4'b1000 : 4'b1110;
														assign node20309 = (inp[12]) ? node20313 : node20310;
															assign node20310 = (inp[4]) ? 4'b1010 : 4'b1001;
															assign node20313 = (inp[4]) ? 4'b1000 : 4'b1010;
												assign node20316 = (inp[4]) ? node20332 : node20317;
													assign node20317 = (inp[12]) ? node20325 : node20318;
														assign node20318 = (inp[5]) ? node20322 : node20319;
															assign node20319 = (inp[15]) ? 4'b1100 : 4'b1000;
															assign node20322 = (inp[15]) ? 4'b1001 : 4'b1101;
														assign node20325 = (inp[5]) ? node20329 : node20326;
															assign node20326 = (inp[15]) ? 4'b1111 : 4'b1010;
															assign node20329 = (inp[15]) ? 4'b1011 : 4'b1111;
													assign node20332 = (inp[12]) ? node20338 : node20333;
														assign node20333 = (inp[15]) ? 4'b1011 : node20334;
															assign node20334 = (inp[5]) ? 4'b1111 : 4'b1011;
														assign node20338 = (inp[5]) ? 4'b1001 : node20339;
															assign node20339 = (inp[15]) ? 4'b1101 : 4'b1001;
							assign node20343 = (inp[13]) ? node20657 : node20344;
								assign node20344 = (inp[7]) ? node20464 : node20345;
									assign node20345 = (inp[1]) ? node20389 : node20346;
										assign node20346 = (inp[2]) ? node20368 : node20347;
											assign node20347 = (inp[4]) ? node20351 : node20348;
												assign node20348 = (inp[12]) ? 4'b1010 : 4'b1000;
												assign node20351 = (inp[12]) ? node20361 : node20352;
													assign node20352 = (inp[5]) ? node20354 : 4'b1010;
														assign node20354 = (inp[11]) ? node20358 : node20355;
															assign node20355 = (inp[15]) ? 4'b1110 : 4'b1010;
															assign node20358 = (inp[15]) ? 4'b1111 : 4'b1011;
													assign node20361 = (inp[5]) ? 4'b1001 : node20362;
														assign node20362 = (inp[15]) ? node20364 : 4'b1100;
															assign node20364 = (inp[11]) ? 4'b1001 : 4'b1000;
											assign node20368 = (inp[4]) ? node20372 : node20369;
												assign node20369 = (inp[12]) ? 4'b1110 : 4'b1100;
												assign node20372 = (inp[12]) ? node20380 : node20373;
													assign node20373 = (inp[5]) ? node20375 : 4'b1111;
														assign node20375 = (inp[15]) ? 4'b1010 : node20376;
															assign node20376 = (inp[9]) ? 4'b1110 : 4'b1111;
													assign node20380 = (inp[5]) ? 4'b1100 : node20381;
														assign node20381 = (inp[15]) ? node20385 : node20382;
															assign node20382 = (inp[11]) ? 4'b1000 : 4'b1001;
															assign node20385 = (inp[11]) ? 4'b1100 : 4'b1101;
										assign node20389 = (inp[2]) ? node20427 : node20390;
											assign node20390 = (inp[4]) ? node20402 : node20391;
												assign node20391 = (inp[12]) ? node20397 : node20392;
													assign node20392 = (inp[11]) ? node20394 : 4'b1100;
														assign node20394 = (inp[15]) ? 4'b1101 : 4'b1100;
													assign node20397 = (inp[15]) ? node20399 : 4'b1111;
														assign node20399 = (inp[11]) ? 4'b1110 : 4'b1111;
												assign node20402 = (inp[12]) ? node20416 : node20403;
													assign node20403 = (inp[15]) ? node20409 : node20404;
														assign node20404 = (inp[11]) ? node20406 : 4'b1110;
															assign node20406 = (inp[5]) ? 4'b1111 : 4'b1110;
														assign node20409 = (inp[5]) ? node20413 : node20410;
															assign node20410 = (inp[11]) ? 4'b1111 : 4'b1110;
															assign node20413 = (inp[11]) ? 4'b1010 : 4'b1011;
													assign node20416 = (inp[15]) ? node20422 : node20417;
														assign node20417 = (inp[5]) ? 4'b1100 : node20418;
															assign node20418 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node20422 = (inp[5]) ? node20424 : 4'b1100;
															assign node20424 = (inp[11]) ? 4'b1101 : 4'b1100;
											assign node20427 = (inp[4]) ? node20439 : node20428;
												assign node20428 = (inp[12]) ? node20434 : node20429;
													assign node20429 = (inp[11]) ? 4'b1001 : node20430;
														assign node20430 = (inp[15]) ? 4'b1001 : 4'b1000;
													assign node20434 = (inp[11]) ? 4'b1010 : node20435;
														assign node20435 = (inp[15]) ? 4'b1010 : 4'b1011;
												assign node20439 = (inp[12]) ? node20451 : node20440;
													assign node20440 = (inp[5]) ? node20446 : node20441;
														assign node20441 = (inp[15]) ? 4'b1010 : node20442;
															assign node20442 = (inp[9]) ? 4'b1011 : 4'b1010;
														assign node20446 = (inp[15]) ? node20448 : 4'b1010;
															assign node20448 = (inp[11]) ? 4'b1111 : 4'b1110;
													assign node20451 = (inp[15]) ? node20459 : node20452;
														assign node20452 = (inp[5]) ? node20456 : node20453;
															assign node20453 = (inp[11]) ? 4'b1101 : 4'b1100;
															assign node20456 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node20459 = (inp[11]) ? 4'b1000 : node20460;
															assign node20460 = (inp[5]) ? 4'b1000 : 4'b1001;
									assign node20464 = (inp[4]) ? node20570 : node20465;
										assign node20465 = (inp[12]) ? node20521 : node20466;
											assign node20466 = (inp[15]) ? node20496 : node20467;
												assign node20467 = (inp[5]) ? node20477 : node20468;
													assign node20468 = (inp[1]) ? node20472 : node20469;
														assign node20469 = (inp[2]) ? 4'b1100 : 4'b1000;
														assign node20472 = (inp[2]) ? node20474 : 4'b1100;
															assign node20474 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node20477 = (inp[11]) ? node20489 : node20478;
														assign node20478 = (inp[9]) ? node20484 : node20479;
															assign node20479 = (inp[2]) ? node20481 : 4'b1001;
																assign node20481 = (inp[1]) ? 4'b1101 : 4'b1001;
															assign node20484 = (inp[2]) ? 4'b1001 : node20485;
																assign node20485 = (inp[1]) ? 4'b1001 : 4'b1101;
														assign node20489 = (inp[1]) ? node20493 : node20490;
															assign node20490 = (inp[2]) ? 4'b1000 : 4'b1101;
															assign node20493 = (inp[2]) ? 4'b1100 : 4'b1000;
												assign node20496 = (inp[5]) ? node20506 : node20497;
													assign node20497 = (inp[1]) ? node20503 : node20498;
														assign node20498 = (inp[2]) ? node20500 : 4'b1100;
															assign node20500 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node20503 = (inp[2]) ? 4'b1101 : 4'b1001;
													assign node20506 = (inp[11]) ? node20514 : node20507;
														assign node20507 = (inp[1]) ? node20511 : node20508;
															assign node20508 = (inp[2]) ? 4'b1101 : 4'b1001;
															assign node20511 = (inp[2]) ? 4'b1000 : 4'b1100;
														assign node20514 = (inp[2]) ? node20518 : node20515;
															assign node20515 = (inp[1]) ? 4'b1100 : 4'b1000;
															assign node20518 = (inp[1]) ? 4'b1001 : 4'b1100;
											assign node20521 = (inp[15]) ? node20545 : node20522;
												assign node20522 = (inp[5]) ? node20536 : node20523;
													assign node20523 = (inp[1]) ? node20531 : node20524;
														assign node20524 = (inp[2]) ? node20528 : node20525;
															assign node20525 = (inp[11]) ? 4'b1011 : 4'b1010;
															assign node20528 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node20531 = (inp[2]) ? 4'b1010 : node20532;
															assign node20532 = (inp[11]) ? 4'b1110 : 4'b1111;
													assign node20536 = (inp[1]) ? node20542 : node20537;
														assign node20537 = (inp[2]) ? 4'b1010 : node20538;
															assign node20538 = (inp[11]) ? 4'b1110 : 4'b1111;
														assign node20542 = (inp[2]) ? 4'b1111 : 4'b1011;
												assign node20545 = (inp[5]) ? node20561 : node20546;
													assign node20546 = (inp[11]) ? node20554 : node20547;
														assign node20547 = (inp[9]) ? 4'b1110 : node20548;
															assign node20548 = (inp[2]) ? 4'b1110 : node20549;
																assign node20549 = (inp[1]) ? 4'b1010 : 4'b1110;
														assign node20554 = (inp[2]) ? node20558 : node20555;
															assign node20555 = (inp[1]) ? 4'b1011 : 4'b1111;
															assign node20558 = (inp[1]) ? 4'b1111 : 4'b1011;
													assign node20561 = (inp[2]) ? node20567 : node20562;
														assign node20562 = (inp[1]) ? node20564 : 4'b1010;
															assign node20564 = (inp[11]) ? 4'b1110 : 4'b1111;
														assign node20567 = (inp[1]) ? 4'b1010 : 4'b1110;
										assign node20570 = (inp[12]) ? node20614 : node20571;
											assign node20571 = (inp[2]) ? node20593 : node20572;
												assign node20572 = (inp[1]) ? node20584 : node20573;
													assign node20573 = (inp[15]) ? node20579 : node20574;
														assign node20574 = (inp[5]) ? node20576 : 4'b1010;
															assign node20576 = (inp[11]) ? 4'b1110 : 4'b1111;
														assign node20579 = (inp[11]) ? node20581 : 4'b1010;
															assign node20581 = (inp[5]) ? 4'b1010 : 4'b1011;
													assign node20584 = (inp[15]) ? node20588 : node20585;
														assign node20585 = (inp[5]) ? 4'b1010 : 4'b1110;
														assign node20588 = (inp[5]) ? node20590 : 4'b1111;
															assign node20590 = (inp[11]) ? 4'b1111 : 4'b1110;
												assign node20593 = (inp[1]) ? node20603 : node20594;
													assign node20594 = (inp[15]) ? node20598 : node20595;
														assign node20595 = (inp[5]) ? 4'b1011 : 4'b1111;
														assign node20598 = (inp[5]) ? 4'b1111 : node20599;
															assign node20599 = (inp[11]) ? 4'b1110 : 4'b1111;
													assign node20603 = (inp[15]) ? node20609 : node20604;
														assign node20604 = (inp[5]) ? 4'b1111 : node20605;
															assign node20605 = (inp[11]) ? 4'b1010 : 4'b1011;
														assign node20609 = (inp[5]) ? 4'b1010 : node20610;
															assign node20610 = (inp[11]) ? 4'b1011 : 4'b1010;
											assign node20614 = (inp[2]) ? node20636 : node20615;
												assign node20615 = (inp[1]) ? node20625 : node20616;
													assign node20616 = (inp[5]) ? node20620 : node20617;
														assign node20617 = (inp[15]) ? 4'b1101 : 4'b1001;
														assign node20620 = (inp[15]) ? 4'b1001 : node20621;
															assign node20621 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node20625 = (inp[15]) ? node20631 : node20626;
														assign node20626 = (inp[5]) ? node20628 : 4'b1100;
															assign node20628 = (inp[11]) ? 4'b1100 : 4'b1101;
														assign node20631 = (inp[5]) ? node20633 : 4'b1001;
															assign node20633 = (inp[11]) ? 4'b1101 : 4'b1100;
												assign node20636 = (inp[1]) ? node20648 : node20637;
													assign node20637 = (inp[5]) ? node20643 : node20638;
														assign node20638 = (inp[15]) ? node20640 : 4'b1100;
															assign node20640 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node20643 = (inp[15]) ? 4'b1100 : node20644;
															assign node20644 = (inp[11]) ? 4'b1100 : 4'b1101;
													assign node20648 = (inp[15]) ? node20654 : node20649;
														assign node20649 = (inp[5]) ? 4'b1001 : node20650;
															assign node20650 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node20654 = (inp[5]) ? 4'b1000 : 4'b1100;
								assign node20657 = (inp[1]) ? node20869 : node20658;
									assign node20658 = (inp[2]) ? node20762 : node20659;
										assign node20659 = (inp[7]) ? node20711 : node20660;
											assign node20660 = (inp[4]) ? node20686 : node20661;
												assign node20661 = (inp[12]) ? node20679 : node20662;
													assign node20662 = (inp[5]) ? node20668 : node20663;
														assign node20663 = (inp[11]) ? 4'b1001 : node20664;
															assign node20664 = (inp[15]) ? 4'b1001 : 4'b1000;
														assign node20668 = (inp[9]) ? node20674 : node20669;
															assign node20669 = (inp[11]) ? node20671 : 4'b1000;
																assign node20671 = (inp[15]) ? 4'b1000 : 4'b1001;
															assign node20674 = (inp[15]) ? node20676 : 4'b1001;
																assign node20676 = (inp[11]) ? 4'b1000 : 4'b1001;
													assign node20679 = (inp[11]) ? node20683 : node20680;
														assign node20680 = (inp[15]) ? 4'b1011 : 4'b1010;
														assign node20683 = (inp[15]) ? 4'b1010 : 4'b1011;
												assign node20686 = (inp[12]) ? node20698 : node20687;
													assign node20687 = (inp[15]) ? node20693 : node20688;
														assign node20688 = (inp[5]) ? 4'b1011 : node20689;
															assign node20689 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node20693 = (inp[5]) ? 4'b1110 : node20694;
															assign node20694 = (inp[11]) ? 4'b1010 : 4'b1011;
													assign node20698 = (inp[5]) ? node20704 : node20699;
														assign node20699 = (inp[15]) ? 4'b1000 : node20700;
															assign node20700 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node20704 = (inp[11]) ? node20708 : node20705;
															assign node20705 = (inp[15]) ? 4'b1000 : 4'b1001;
															assign node20708 = (inp[15]) ? 4'b1001 : 4'b1000;
											assign node20711 = (inp[4]) ? node20737 : node20712;
												assign node20712 = (inp[12]) ? node20728 : node20713;
													assign node20713 = (inp[11]) ? node20721 : node20714;
														assign node20714 = (inp[9]) ? 4'b1101 : node20715;
															assign node20715 = (inp[15]) ? node20717 : 4'b1000;
																assign node20717 = (inp[5]) ? 4'b1001 : 4'b1101;
														assign node20721 = (inp[15]) ? node20725 : node20722;
															assign node20722 = (inp[5]) ? 4'b1100 : 4'b1001;
															assign node20725 = (inp[5]) ? 4'b1001 : 4'b1100;
													assign node20728 = (inp[15]) ? node20732 : node20729;
														assign node20729 = (inp[5]) ? 4'b1110 : 4'b1011;
														assign node20732 = (inp[5]) ? node20734 : 4'b1110;
															assign node20734 = (inp[11]) ? 4'b1010 : 4'b1011;
												assign node20737 = (inp[12]) ? node20749 : node20738;
													assign node20738 = (inp[15]) ? node20744 : node20739;
														assign node20739 = (inp[5]) ? 4'b1110 : node20740;
															assign node20740 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node20744 = (inp[5]) ? node20746 : 4'b1010;
															assign node20746 = (inp[11]) ? 4'b1010 : 4'b1011;
													assign node20749 = (inp[15]) ? node20755 : node20750;
														assign node20750 = (inp[11]) ? node20752 : 4'b1001;
															assign node20752 = (inp[5]) ? 4'b1001 : 4'b1000;
														assign node20755 = (inp[5]) ? node20759 : node20756;
															assign node20756 = (inp[11]) ? 4'b1101 : 4'b1100;
															assign node20759 = (inp[11]) ? 4'b1001 : 4'b1000;
										assign node20762 = (inp[7]) ? node20804 : node20763;
											assign node20763 = (inp[4]) ? node20779 : node20764;
												assign node20764 = (inp[12]) ? node20772 : node20765;
													assign node20765 = (inp[15]) ? node20769 : node20766;
														assign node20766 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node20769 = (inp[11]) ? 4'b1100 : 4'b1101;
													assign node20772 = (inp[15]) ? node20776 : node20773;
														assign node20773 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node20776 = (inp[11]) ? 4'b1110 : 4'b1111;
												assign node20779 = (inp[12]) ? node20793 : node20780;
													assign node20780 = (inp[5]) ? node20788 : node20781;
														assign node20781 = (inp[11]) ? node20785 : node20782;
															assign node20782 = (inp[15]) ? 4'b1110 : 4'b1111;
															assign node20785 = (inp[15]) ? 4'b1111 : 4'b1110;
														assign node20788 = (inp[15]) ? node20790 : 4'b1110;
															assign node20790 = (inp[11]) ? 4'b1010 : 4'b1011;
													assign node20793 = (inp[15]) ? node20799 : node20794;
														assign node20794 = (inp[5]) ? node20796 : 4'b1000;
															assign node20796 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node20799 = (inp[5]) ? node20801 : 4'b1101;
															assign node20801 = (inp[11]) ? 4'b1100 : 4'b1101;
											assign node20804 = (inp[4]) ? node20844 : node20805;
												assign node20805 = (inp[12]) ? node20821 : node20806;
													assign node20806 = (inp[11]) ? node20814 : node20807;
														assign node20807 = (inp[5]) ? node20811 : node20808;
															assign node20808 = (inp[15]) ? 4'b1000 : 4'b1100;
															assign node20811 = (inp[15]) ? 4'b1101 : 4'b1000;
														assign node20814 = (inp[15]) ? node20818 : node20815;
															assign node20815 = (inp[5]) ? 4'b1000 : 4'b1101;
															assign node20818 = (inp[5]) ? 4'b1101 : 4'b1000;
													assign node20821 = (inp[11]) ? node20837 : node20822;
														assign node20822 = (inp[9]) ? node20830 : node20823;
															assign node20823 = (inp[15]) ? node20827 : node20824;
																assign node20824 = (inp[5]) ? 4'b1010 : 4'b1111;
																assign node20827 = (inp[5]) ? 4'b1111 : 4'b1010;
															assign node20830 = (inp[15]) ? node20834 : node20831;
																assign node20831 = (inp[5]) ? 4'b1010 : 4'b1111;
																assign node20834 = (inp[5]) ? 4'b1111 : 4'b1010;
														assign node20837 = (inp[5]) ? node20841 : node20838;
															assign node20838 = (inp[15]) ? 4'b1011 : 4'b1111;
															assign node20841 = (inp[9]) ? 4'b1110 : 4'b1011;
												assign node20844 = (inp[12]) ? node20858 : node20845;
													assign node20845 = (inp[5]) ? node20851 : node20846;
														assign node20846 = (inp[11]) ? node20848 : 4'b1111;
															assign node20848 = (inp[15]) ? 4'b1111 : 4'b1110;
														assign node20851 = (inp[15]) ? node20855 : node20852;
															assign node20852 = (inp[11]) ? 4'b1010 : 4'b1011;
															assign node20855 = (inp[11]) ? 4'b1111 : 4'b1110;
													assign node20858 = (inp[5]) ? node20864 : node20859;
														assign node20859 = (inp[15]) ? 4'b1000 : node20860;
															assign node20860 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node20864 = (inp[11]) ? 4'b1100 : node20865;
															assign node20865 = (inp[15]) ? 4'b1101 : 4'b1100;
									assign node20869 = (inp[2]) ? node20963 : node20870;
										assign node20870 = (inp[7]) ? node20904 : node20871;
											assign node20871 = (inp[4]) ? node20883 : node20872;
												assign node20872 = (inp[12]) ? node20878 : node20873;
													assign node20873 = (inp[15]) ? 4'b1100 : node20874;
														assign node20874 = (inp[11]) ? 4'b1101 : 4'b1100;
													assign node20878 = (inp[11]) ? node20880 : 4'b1111;
														assign node20880 = (inp[15]) ? 4'b1111 : 4'b1110;
												assign node20883 = (inp[12]) ? node20893 : node20884;
													assign node20884 = (inp[5]) ? node20890 : node20885;
														assign node20885 = (inp[15]) ? 4'b1110 : node20886;
															assign node20886 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node20890 = (inp[15]) ? 4'b1011 : 4'b1111;
													assign node20893 = (inp[5]) ? node20899 : node20894;
														assign node20894 = (inp[15]) ? node20896 : 4'b1000;
															assign node20896 = (inp[11]) ? 4'b1100 : 4'b1101;
														assign node20899 = (inp[15]) ? 4'b1100 : node20900;
															assign node20900 = (inp[11]) ? 4'b1101 : 4'b1100;
											assign node20904 = (inp[11]) ? node20932 : node20905;
												assign node20905 = (inp[4]) ? node20921 : node20906;
													assign node20906 = (inp[12]) ? node20914 : node20907;
														assign node20907 = (inp[15]) ? node20911 : node20908;
															assign node20908 = (inp[5]) ? 4'b1000 : 4'b1100;
															assign node20911 = (inp[5]) ? 4'b1101 : 4'b1000;
														assign node20914 = (inp[5]) ? node20918 : node20915;
															assign node20915 = (inp[15]) ? 4'b1010 : 4'b1110;
															assign node20918 = (inp[15]) ? 4'b1111 : 4'b1011;
													assign node20921 = (inp[12]) ? node20927 : node20922;
														assign node20922 = (inp[15]) ? 4'b1110 : node20923;
															assign node20923 = (inp[5]) ? 4'b1010 : 4'b1110;
														assign node20927 = (inp[5]) ? 4'b1100 : node20928;
															assign node20928 = (inp[15]) ? 4'b1000 : 4'b1100;
												assign node20932 = (inp[5]) ? node20948 : node20933;
													assign node20933 = (inp[15]) ? node20941 : node20934;
														assign node20934 = (inp[12]) ? node20938 : node20935;
															assign node20935 = (inp[4]) ? 4'b1111 : 4'b1101;
															assign node20938 = (inp[4]) ? 4'b1101 : 4'b1110;
														assign node20941 = (inp[4]) ? node20945 : node20942;
															assign node20942 = (inp[12]) ? 4'b1010 : 4'b1001;
															assign node20945 = (inp[12]) ? 4'b1001 : 4'b1111;
													assign node20948 = (inp[15]) ? node20956 : node20949;
														assign node20949 = (inp[4]) ? node20953 : node20950;
															assign node20950 = (inp[12]) ? 4'b1010 : 4'b1000;
															assign node20953 = (inp[12]) ? 4'b1100 : 4'b1011;
														assign node20956 = (inp[4]) ? node20960 : node20957;
															assign node20957 = (inp[12]) ? 4'b1111 : 4'b1100;
															assign node20960 = (inp[12]) ? 4'b1100 : 4'b1110;
										assign node20963 = (inp[7]) ? node20997 : node20964;
											assign node20964 = (inp[4]) ? node20976 : node20965;
												assign node20965 = (inp[12]) ? node20971 : node20966;
													assign node20966 = (inp[15]) ? node20968 : 4'b1001;
														assign node20968 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node20971 = (inp[15]) ? node20973 : 4'b1010;
														assign node20973 = (inp[11]) ? 4'b1010 : 4'b1011;
												assign node20976 = (inp[12]) ? node20988 : node20977;
													assign node20977 = (inp[15]) ? node20983 : node20978;
														assign node20978 = (inp[11]) ? node20980 : 4'b1010;
															assign node20980 = (inp[5]) ? 4'b1011 : 4'b1010;
														assign node20983 = (inp[5]) ? 4'b1110 : node20984;
															assign node20984 = (inp[11]) ? 4'b1010 : 4'b1011;
													assign node20988 = (inp[5]) ? node20992 : node20989;
														assign node20989 = (inp[15]) ? 4'b1001 : 4'b1101;
														assign node20992 = (inp[11]) ? 4'b1000 : node20993;
															assign node20993 = (inp[15]) ? 4'b1001 : 4'b1000;
											assign node20997 = (inp[11]) ? node21029 : node20998;
												assign node20998 = (inp[5]) ? node21014 : node20999;
													assign node20999 = (inp[15]) ? node21007 : node21000;
														assign node21000 = (inp[12]) ? node21004 : node21001;
															assign node21001 = (inp[4]) ? 4'b1010 : 4'b1001;
															assign node21004 = (inp[4]) ? 4'b1000 : 4'b1010;
														assign node21007 = (inp[12]) ? node21011 : node21008;
															assign node21008 = (inp[4]) ? 4'b1010 : 4'b1100;
															assign node21011 = (inp[4]) ? 4'b1101 : 4'b1110;
													assign node21014 = (inp[15]) ? node21022 : node21015;
														assign node21015 = (inp[12]) ? node21019 : node21016;
															assign node21016 = (inp[4]) ? 4'b1111 : 4'b1100;
															assign node21019 = (inp[4]) ? 4'b1001 : 4'b1111;
														assign node21022 = (inp[12]) ? node21026 : node21023;
															assign node21023 = (inp[4]) ? 4'b1011 : 4'b1000;
															assign node21026 = (inp[4]) ? 4'b1001 : 4'b1011;
												assign node21029 = (inp[4]) ? node21045 : node21030;
													assign node21030 = (inp[12]) ? node21038 : node21031;
														assign node21031 = (inp[5]) ? node21035 : node21032;
															assign node21032 = (inp[15]) ? 4'b1101 : 4'b1001;
															assign node21035 = (inp[15]) ? 4'b1000 : 4'b1100;
														assign node21038 = (inp[5]) ? node21042 : node21039;
															assign node21039 = (inp[15]) ? 4'b1110 : 4'b1011;
															assign node21042 = (inp[15]) ? 4'b1010 : 4'b1110;
													assign node21045 = (inp[12]) ? node21051 : node21046;
														assign node21046 = (inp[15]) ? 4'b1010 : node21047;
															assign node21047 = (inp[5]) ? 4'b1110 : 4'b1010;
														assign node21051 = (inp[5]) ? 4'b1000 : node21052;
															assign node21052 = (inp[15]) ? 4'b1100 : 4'b1000;
					assign node21056 = (inp[10]) ? node22484 : node21057;
						assign node21057 = (inp[11]) ? node21767 : node21058;
							assign node21058 = (inp[0]) ? node21442 : node21059;
								assign node21059 = (inp[13]) ? node21247 : node21060;
									assign node21060 = (inp[4]) ? node21136 : node21061;
										assign node21061 = (inp[15]) ? node21099 : node21062;
											assign node21062 = (inp[1]) ? node21076 : node21063;
												assign node21063 = (inp[5]) ? node21071 : node21064;
													assign node21064 = (inp[12]) ? node21066 : 4'b0000;
														assign node21066 = (inp[7]) ? node21068 : 4'b0000;
															assign node21068 = (inp[2]) ? 4'b0101 : 4'b0100;
													assign node21071 = (inp[7]) ? node21073 : 4'b0100;
														assign node21073 = (inp[12]) ? 4'b0000 : 4'b0101;
												assign node21076 = (inp[5]) ? node21084 : node21077;
													assign node21077 = (inp[7]) ? node21081 : node21078;
														assign node21078 = (inp[12]) ? 4'b0101 : 4'b0100;
														assign node21081 = (inp[12]) ? 4'b0000 : 4'b0100;
													assign node21084 = (inp[12]) ? node21094 : node21085;
														assign node21085 = (inp[9]) ? node21087 : 4'b0001;
															assign node21087 = (inp[2]) ? node21091 : node21088;
																assign node21088 = (inp[7]) ? 4'b0001 : 4'b0000;
																assign node21091 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node21094 = (inp[7]) ? 4'b0101 : node21095;
															assign node21095 = (inp[2]) ? 4'b0000 : 4'b0001;
											assign node21099 = (inp[5]) ? node21121 : node21100;
												assign node21100 = (inp[1]) ? node21108 : node21101;
													assign node21101 = (inp[12]) ? node21105 : node21102;
														assign node21102 = (inp[7]) ? 4'b0110 : 4'b0010;
														assign node21105 = (inp[7]) ? 4'b0011 : 4'b0010;
													assign node21108 = (inp[7]) ? node21116 : node21109;
														assign node21109 = (inp[2]) ? node21113 : node21110;
															assign node21110 = (inp[12]) ? 4'b0111 : 4'b0110;
															assign node21113 = (inp[12]) ? 4'b0110 : 4'b0111;
														assign node21116 = (inp[12]) ? node21118 : 4'b0011;
															assign node21118 = (inp[2]) ? 4'b0111 : 4'b0110;
												assign node21121 = (inp[1]) ? node21129 : node21122;
													assign node21122 = (inp[12]) ? 4'b0110 : node21123;
														assign node21123 = (inp[7]) ? node21125 : 4'b0110;
															assign node21125 = (inp[2]) ? 4'b0010 : 4'b0011;
													assign node21129 = (inp[7]) ? node21133 : node21130;
														assign node21130 = (inp[12]) ? 4'b0010 : 4'b0011;
														assign node21133 = (inp[12]) ? 4'b0010 : 4'b0110;
										assign node21136 = (inp[15]) ? node21194 : node21137;
											assign node21137 = (inp[2]) ? node21171 : node21138;
												assign node21138 = (inp[5]) ? node21158 : node21139;
													assign node21139 = (inp[12]) ? node21143 : node21140;
														assign node21140 = (inp[1]) ? 4'b0110 : 4'b0010;
														assign node21143 = (inp[9]) ? node21151 : node21144;
															assign node21144 = (inp[7]) ? node21148 : node21145;
																assign node21145 = (inp[1]) ? 4'b0011 : 4'b0110;
																assign node21148 = (inp[1]) ? 4'b0110 : 4'b0011;
															assign node21151 = (inp[7]) ? node21155 : node21152;
																assign node21152 = (inp[1]) ? 4'b0011 : 4'b0110;
																assign node21155 = (inp[1]) ? 4'b0110 : 4'b0011;
													assign node21158 = (inp[1]) ? node21166 : node21159;
														assign node21159 = (inp[12]) ? node21163 : node21160;
															assign node21160 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node21163 = (inp[7]) ? 4'b0110 : 4'b0011;
														assign node21166 = (inp[12]) ? 4'b0110 : node21167;
															assign node21167 = (inp[7]) ? 4'b0010 : 4'b0011;
												assign node21171 = (inp[5]) ? node21181 : node21172;
													assign node21172 = (inp[1]) ? node21176 : node21173;
														assign node21173 = (inp[12]) ? 4'b0111 : 4'b0011;
														assign node21176 = (inp[7]) ? 4'b0111 : node21177;
															assign node21177 = (inp[12]) ? 4'b0011 : 4'b0111;
													assign node21181 = (inp[1]) ? node21189 : node21182;
														assign node21182 = (inp[7]) ? node21186 : node21183;
															assign node21183 = (inp[12]) ? 4'b0010 : 4'b0110;
															assign node21186 = (inp[12]) ? 4'b0110 : 4'b0111;
														assign node21189 = (inp[7]) ? 4'b0011 : node21190;
															assign node21190 = (inp[12]) ? 4'b0111 : 4'b0010;
											assign node21194 = (inp[2]) ? node21220 : node21195;
												assign node21195 = (inp[5]) ? node21209 : node21196;
													assign node21196 = (inp[1]) ? node21204 : node21197;
														assign node21197 = (inp[7]) ? node21201 : node21198;
															assign node21198 = (inp[12]) ? 4'b0000 : 4'b0100;
															assign node21201 = (inp[12]) ? 4'b0001 : 4'b0000;
														assign node21204 = (inp[12]) ? node21206 : 4'b0001;
															assign node21206 = (inp[9]) ? 4'b0101 : 4'b0100;
													assign node21209 = (inp[1]) ? node21215 : node21210;
														assign node21210 = (inp[12]) ? 4'b0101 : node21211;
															assign node21211 = (inp[7]) ? 4'b0100 : 4'b0001;
														assign node21215 = (inp[7]) ? 4'b0001 : node21216;
															assign node21216 = (inp[12]) ? 4'b0001 : 4'b0101;
												assign node21220 = (inp[1]) ? node21236 : node21221;
													assign node21221 = (inp[5]) ? node21229 : node21222;
														assign node21222 = (inp[7]) ? node21226 : node21223;
															assign node21223 = (inp[12]) ? 4'b0000 : 4'b0101;
															assign node21226 = (inp[12]) ? 4'b0001 : 4'b0000;
														assign node21229 = (inp[7]) ? node21233 : node21230;
															assign node21230 = (inp[12]) ? 4'b0100 : 4'b0000;
															assign node21233 = (inp[12]) ? 4'b0100 : 4'b0101;
													assign node21236 = (inp[5]) ? node21242 : node21237;
														assign node21237 = (inp[7]) ? 4'b0100 : node21238;
															assign node21238 = (inp[12]) ? 4'b0101 : 4'b0000;
														assign node21242 = (inp[7]) ? 4'b0000 : node21243;
															assign node21243 = (inp[12]) ? 4'b0000 : 4'b0101;
									assign node21247 = (inp[4]) ? node21357 : node21248;
										assign node21248 = (inp[15]) ? node21304 : node21249;
											assign node21249 = (inp[2]) ? node21277 : node21250;
												assign node21250 = (inp[12]) ? node21262 : node21251;
													assign node21251 = (inp[5]) ? node21255 : node21252;
														assign node21252 = (inp[1]) ? 4'b0100 : 4'b0000;
														assign node21255 = (inp[1]) ? node21259 : node21256;
															assign node21256 = (inp[9]) ? 4'b0101 : 4'b0100;
															assign node21259 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node21262 = (inp[7]) ? node21270 : node21263;
														assign node21263 = (inp[1]) ? node21267 : node21264;
															assign node21264 = (inp[5]) ? 4'b0100 : 4'b0000;
															assign node21267 = (inp[5]) ? 4'b0000 : 4'b0101;
														assign node21270 = (inp[5]) ? node21274 : node21271;
															assign node21271 = (inp[1]) ? 4'b0000 : 4'b0101;
															assign node21274 = (inp[1]) ? 4'b0101 : 4'b0000;
												assign node21277 = (inp[1]) ? node21289 : node21278;
													assign node21278 = (inp[5]) ? node21284 : node21279;
														assign node21279 = (inp[12]) ? node21281 : 4'b0001;
															assign node21281 = (inp[7]) ? 4'b0101 : 4'b0001;
														assign node21284 = (inp[7]) ? node21286 : 4'b0101;
															assign node21286 = (inp[12]) ? 4'b0001 : 4'b0100;
													assign node21289 = (inp[5]) ? node21297 : node21290;
														assign node21290 = (inp[7]) ? node21294 : node21291;
															assign node21291 = (inp[12]) ? 4'b0100 : 4'b0101;
															assign node21294 = (inp[12]) ? 4'b0001 : 4'b0101;
														assign node21297 = (inp[12]) ? node21301 : node21298;
															assign node21298 = (inp[7]) ? 4'b0000 : 4'b0001;
															assign node21301 = (inp[7]) ? 4'b0100 : 4'b0000;
											assign node21304 = (inp[2]) ? node21332 : node21305;
												assign node21305 = (inp[1]) ? node21319 : node21306;
													assign node21306 = (inp[5]) ? node21314 : node21307;
														assign node21307 = (inp[12]) ? node21311 : node21308;
															assign node21308 = (inp[7]) ? 4'b0111 : 4'b0011;
															assign node21311 = (inp[7]) ? 4'b0010 : 4'b0011;
														assign node21314 = (inp[7]) ? node21316 : 4'b0111;
															assign node21316 = (inp[12]) ? 4'b0111 : 4'b0011;
													assign node21319 = (inp[5]) ? node21327 : node21320;
														assign node21320 = (inp[12]) ? node21324 : node21321;
															assign node21321 = (inp[7]) ? 4'b0010 : 4'b0110;
															assign node21324 = (inp[7]) ? 4'b0110 : 4'b0111;
														assign node21327 = (inp[12]) ? 4'b0011 : node21328;
															assign node21328 = (inp[7]) ? 4'b0111 : 4'b0010;
												assign node21332 = (inp[12]) ? node21346 : node21333;
													assign node21333 = (inp[7]) ? node21341 : node21334;
														assign node21334 = (inp[5]) ? node21338 : node21335;
															assign node21335 = (inp[1]) ? 4'b0110 : 4'b0010;
															assign node21338 = (inp[1]) ? 4'b0011 : 4'b0110;
														assign node21341 = (inp[1]) ? 4'b0011 : node21342;
															assign node21342 = (inp[5]) ? 4'b0011 : 4'b0110;
													assign node21346 = (inp[5]) ? node21354 : node21347;
														assign node21347 = (inp[1]) ? node21351 : node21348;
															assign node21348 = (inp[7]) ? 4'b0011 : 4'b0010;
															assign node21351 = (inp[7]) ? 4'b0110 : 4'b0111;
														assign node21354 = (inp[1]) ? 4'b0010 : 4'b0110;
										assign node21357 = (inp[15]) ? node21403 : node21358;
											assign node21358 = (inp[1]) ? node21388 : node21359;
												assign node21359 = (inp[5]) ? node21367 : node21360;
													assign node21360 = (inp[7]) ? node21364 : node21361;
														assign node21361 = (inp[12]) ? 4'b0110 : 4'b0010;
														assign node21364 = (inp[12]) ? 4'b0011 : 4'b0010;
													assign node21367 = (inp[7]) ? node21373 : node21368;
														assign node21368 = (inp[12]) ? 4'b0011 : node21369;
															assign node21369 = (inp[2]) ? 4'b0110 : 4'b0111;
														assign node21373 = (inp[9]) ? node21381 : node21374;
															assign node21374 = (inp[12]) ? node21378 : node21375;
																assign node21375 = (inp[2]) ? 4'b0111 : 4'b0110;
																assign node21378 = (inp[2]) ? 4'b0110 : 4'b0111;
															assign node21381 = (inp[12]) ? node21385 : node21382;
																assign node21382 = (inp[2]) ? 4'b0111 : 4'b0110;
																assign node21385 = (inp[2]) ? 4'b0110 : 4'b0111;
												assign node21388 = (inp[5]) ? node21396 : node21389;
													assign node21389 = (inp[7]) ? 4'b0110 : node21390;
														assign node21390 = (inp[12]) ? node21392 : 4'b0110;
															assign node21392 = (inp[2]) ? 4'b0011 : 4'b0010;
													assign node21396 = (inp[12]) ? node21400 : node21397;
														assign node21397 = (inp[7]) ? 4'b0010 : 4'b0011;
														assign node21400 = (inp[7]) ? 4'b0010 : 4'b0110;
											assign node21403 = (inp[7]) ? node21429 : node21404;
												assign node21404 = (inp[5]) ? node21420 : node21405;
													assign node21405 = (inp[2]) ? node21413 : node21406;
														assign node21406 = (inp[1]) ? node21410 : node21407;
															assign node21407 = (inp[12]) ? 4'b0000 : 4'b0101;
															assign node21410 = (inp[12]) ? 4'b0101 : 4'b0000;
														assign node21413 = (inp[12]) ? node21417 : node21414;
															assign node21414 = (inp[1]) ? 4'b0000 : 4'b0101;
															assign node21417 = (inp[1]) ? 4'b0101 : 4'b0001;
													assign node21420 = (inp[1]) ? node21424 : node21421;
														assign node21421 = (inp[12]) ? 4'b0100 : 4'b0000;
														assign node21424 = (inp[12]) ? 4'b0000 : node21425;
															assign node21425 = (inp[2]) ? 4'b0100 : 4'b0101;
												assign node21429 = (inp[1]) ? node21439 : node21430;
													assign node21430 = (inp[5]) ? node21436 : node21431;
														assign node21431 = (inp[2]) ? 4'b0000 : node21432;
															assign node21432 = (inp[12]) ? 4'b0001 : 4'b0000;
														assign node21436 = (inp[12]) ? 4'b0100 : 4'b0101;
													assign node21439 = (inp[5]) ? 4'b0000 : 4'b0100;
								assign node21442 = (inp[7]) ? node21608 : node21443;
									assign node21443 = (inp[1]) ? node21513 : node21444;
										assign node21444 = (inp[5]) ? node21478 : node21445;
											assign node21445 = (inp[4]) ? node21457 : node21446;
												assign node21446 = (inp[15]) ? node21452 : node21447;
													assign node21447 = (inp[2]) ? node21449 : 4'b0001;
														assign node21449 = (inp[13]) ? 4'b0000 : 4'b0001;
													assign node21452 = (inp[13]) ? node21454 : 4'b0011;
														assign node21454 = (inp[2]) ? 4'b0011 : 4'b0010;
												assign node21457 = (inp[15]) ? node21469 : node21458;
													assign node21458 = (inp[12]) ? node21464 : node21459;
														assign node21459 = (inp[13]) ? 4'b0011 : node21460;
															assign node21460 = (inp[2]) ? 4'b0010 : 4'b0011;
														assign node21464 = (inp[13]) ? 4'b0111 : node21465;
															assign node21465 = (inp[2]) ? 4'b0110 : 4'b0111;
													assign node21469 = (inp[12]) ? node21475 : node21470;
														assign node21470 = (inp[2]) ? 4'b0100 : node21471;
															assign node21471 = (inp[9]) ? 4'b0101 : 4'b0100;
														assign node21475 = (inp[2]) ? 4'b0000 : 4'b0001;
											assign node21478 = (inp[4]) ? node21490 : node21479;
												assign node21479 = (inp[15]) ? node21485 : node21480;
													assign node21480 = (inp[2]) ? node21482 : 4'b0101;
														assign node21482 = (inp[13]) ? 4'b0100 : 4'b0101;
													assign node21485 = (inp[13]) ? node21487 : 4'b0111;
														assign node21487 = (inp[2]) ? 4'b0111 : 4'b0110;
												assign node21490 = (inp[15]) ? node21502 : node21491;
													assign node21491 = (inp[12]) ? node21497 : node21492;
														assign node21492 = (inp[13]) ? node21494 : 4'b0111;
															assign node21494 = (inp[2]) ? 4'b0111 : 4'b0110;
														assign node21497 = (inp[13]) ? 4'b0010 : node21498;
															assign node21498 = (inp[2]) ? 4'b0011 : 4'b0010;
													assign node21502 = (inp[12]) ? node21508 : node21503;
														assign node21503 = (inp[2]) ? 4'b0001 : node21504;
															assign node21504 = (inp[13]) ? 4'b0001 : 4'b0000;
														assign node21508 = (inp[13]) ? 4'b0101 : node21509;
															assign node21509 = (inp[2]) ? 4'b0101 : 4'b0100;
										assign node21513 = (inp[5]) ? node21561 : node21514;
											assign node21514 = (inp[12]) ? node21538 : node21515;
												assign node21515 = (inp[15]) ? node21527 : node21516;
													assign node21516 = (inp[4]) ? node21522 : node21517;
														assign node21517 = (inp[2]) ? node21519 : 4'b0101;
															assign node21519 = (inp[9]) ? 4'b0101 : 4'b0100;
														assign node21522 = (inp[13]) ? 4'b0111 : node21523;
															assign node21523 = (inp[2]) ? 4'b0110 : 4'b0111;
													assign node21527 = (inp[4]) ? node21533 : node21528;
														assign node21528 = (inp[13]) ? 4'b0111 : node21529;
															assign node21529 = (inp[2]) ? 4'b0110 : 4'b0111;
														assign node21533 = (inp[13]) ? 4'b0001 : node21534;
															assign node21534 = (inp[2]) ? 4'b0001 : 4'b0000;
												assign node21538 = (inp[15]) ? node21550 : node21539;
													assign node21539 = (inp[4]) ? node21545 : node21540;
														assign node21540 = (inp[2]) ? node21542 : 4'b0100;
															assign node21542 = (inp[13]) ? 4'b0101 : 4'b0100;
														assign node21545 = (inp[13]) ? node21547 : 4'b0010;
															assign node21547 = (inp[2]) ? 4'b0010 : 4'b0011;
													assign node21550 = (inp[4]) ? node21556 : node21551;
														assign node21551 = (inp[2]) ? node21553 : 4'b0110;
															assign node21553 = (inp[13]) ? 4'b0110 : 4'b0111;
														assign node21556 = (inp[2]) ? 4'b0100 : node21557;
															assign node21557 = (inp[13]) ? 4'b0100 : 4'b0101;
											assign node21561 = (inp[4]) ? node21585 : node21562;
												assign node21562 = (inp[15]) ? node21574 : node21563;
													assign node21563 = (inp[12]) ? node21569 : node21564;
														assign node21564 = (inp[13]) ? 4'b0000 : node21565;
															assign node21565 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node21569 = (inp[13]) ? 4'b0001 : node21570;
															assign node21570 = (inp[2]) ? 4'b0001 : 4'b0000;
													assign node21574 = (inp[12]) ? node21580 : node21575;
														assign node21575 = (inp[2]) ? 4'b0010 : node21576;
															assign node21576 = (inp[13]) ? 4'b0011 : 4'b0010;
														assign node21580 = (inp[2]) ? 4'b0011 : node21581;
															assign node21581 = (inp[13]) ? 4'b0010 : 4'b0011;
												assign node21585 = (inp[15]) ? node21597 : node21586;
													assign node21586 = (inp[12]) ? node21592 : node21587;
														assign node21587 = (inp[13]) ? 4'b0010 : node21588;
															assign node21588 = (inp[2]) ? 4'b0011 : 4'b0010;
														assign node21592 = (inp[2]) ? node21594 : 4'b0111;
															assign node21594 = (inp[13]) ? 4'b0111 : 4'b0110;
													assign node21597 = (inp[12]) ? node21603 : node21598;
														assign node21598 = (inp[13]) ? node21600 : 4'b0100;
															assign node21600 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node21603 = (inp[2]) ? 4'b0001 : node21604;
															assign node21604 = (inp[13]) ? 4'b0001 : 4'b0000;
									assign node21608 = (inp[1]) ? node21696 : node21609;
										assign node21609 = (inp[5]) ? node21655 : node21610;
											assign node21610 = (inp[12]) ? node21634 : node21611;
												assign node21611 = (inp[4]) ? node21623 : node21612;
													assign node21612 = (inp[15]) ? node21618 : node21613;
														assign node21613 = (inp[2]) ? node21615 : 4'b0001;
															assign node21615 = (inp[13]) ? 4'b0000 : 4'b0001;
														assign node21618 = (inp[2]) ? 4'b0111 : node21619;
															assign node21619 = (inp[13]) ? 4'b0110 : 4'b0111;
													assign node21623 = (inp[15]) ? node21629 : node21624;
														assign node21624 = (inp[13]) ? 4'b0011 : node21625;
															assign node21625 = (inp[2]) ? 4'b0010 : 4'b0011;
														assign node21629 = (inp[2]) ? node21631 : 4'b0001;
															assign node21631 = (inp[13]) ? 4'b0000 : 4'b0001;
												assign node21634 = (inp[15]) ? node21644 : node21635;
													assign node21635 = (inp[4]) ? node21641 : node21636;
														assign node21636 = (inp[2]) ? 4'b0100 : node21637;
															assign node21637 = (inp[13]) ? 4'b0100 : 4'b0101;
														assign node21641 = (inp[13]) ? 4'b0010 : 4'b0011;
													assign node21644 = (inp[4]) ? node21650 : node21645;
														assign node21645 = (inp[13]) ? node21647 : 4'b0010;
															assign node21647 = (inp[2]) ? 4'b0010 : 4'b0011;
														assign node21650 = (inp[2]) ? node21652 : 4'b0000;
															assign node21652 = (inp[13]) ? 4'b0001 : 4'b0000;
											assign node21655 = (inp[4]) ? node21679 : node21656;
												assign node21656 = (inp[15]) ? node21668 : node21657;
													assign node21657 = (inp[12]) ? node21663 : node21658;
														assign node21658 = (inp[2]) ? node21660 : 4'b0100;
															assign node21660 = (inp[13]) ? 4'b0101 : 4'b0100;
														assign node21663 = (inp[13]) ? node21665 : 4'b0001;
															assign node21665 = (inp[2]) ? 4'b0000 : 4'b0001;
													assign node21668 = (inp[12]) ? node21674 : node21669;
														assign node21669 = (inp[13]) ? 4'b0010 : node21670;
															assign node21670 = (inp[2]) ? 4'b0011 : 4'b0010;
														assign node21674 = (inp[13]) ? node21676 : 4'b0111;
															assign node21676 = (inp[2]) ? 4'b0111 : 4'b0110;
												assign node21679 = (inp[15]) ? node21691 : node21680;
													assign node21680 = (inp[12]) ? node21686 : node21681;
														assign node21681 = (inp[2]) ? 4'b0110 : node21682;
															assign node21682 = (inp[13]) ? 4'b0111 : 4'b0110;
														assign node21686 = (inp[2]) ? 4'b0111 : node21687;
															assign node21687 = (inp[13]) ? 4'b0110 : 4'b0111;
													assign node21691 = (inp[12]) ? 4'b0101 : node21692;
														assign node21692 = (inp[2]) ? 4'b0100 : 4'b0101;
										assign node21696 = (inp[5]) ? node21732 : node21697;
											assign node21697 = (inp[4]) ? node21721 : node21698;
												assign node21698 = (inp[15]) ? node21710 : node21699;
													assign node21699 = (inp[12]) ? node21705 : node21700;
														assign node21700 = (inp[13]) ? node21702 : 4'b0101;
															assign node21702 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node21705 = (inp[2]) ? node21707 : 4'b0001;
															assign node21707 = (inp[13]) ? 4'b0000 : 4'b0001;
													assign node21710 = (inp[12]) ? node21716 : node21711;
														assign node21711 = (inp[2]) ? 4'b0010 : node21712;
															assign node21712 = (inp[13]) ? 4'b0011 : 4'b0010;
														assign node21716 = (inp[13]) ? 4'b0111 : node21717;
															assign node21717 = (inp[2]) ? 4'b0110 : 4'b0111;
												assign node21721 = (inp[15]) ? node21727 : node21722;
													assign node21722 = (inp[2]) ? node21724 : 4'b0111;
														assign node21724 = (inp[13]) ? 4'b0111 : 4'b0110;
													assign node21727 = (inp[13]) ? 4'b0101 : node21728;
														assign node21728 = (inp[2]) ? 4'b0101 : 4'b0100;
											assign node21732 = (inp[4]) ? node21756 : node21733;
												assign node21733 = (inp[15]) ? node21745 : node21734;
													assign node21734 = (inp[12]) ? node21740 : node21735;
														assign node21735 = (inp[2]) ? 4'b0001 : node21736;
															assign node21736 = (inp[13]) ? 4'b0001 : 4'b0000;
														assign node21740 = (inp[13]) ? node21742 : 4'b0100;
															assign node21742 = (inp[2]) ? 4'b0101 : 4'b0100;
													assign node21745 = (inp[12]) ? node21751 : node21746;
														assign node21746 = (inp[13]) ? node21748 : 4'b0111;
															assign node21748 = (inp[2]) ? 4'b0111 : 4'b0110;
														assign node21751 = (inp[13]) ? node21753 : 4'b0011;
															assign node21753 = (inp[2]) ? 4'b0011 : 4'b0010;
												assign node21756 = (inp[15]) ? node21762 : node21757;
													assign node21757 = (inp[2]) ? node21759 : 4'b0011;
														assign node21759 = (inp[13]) ? 4'b0011 : 4'b0010;
													assign node21762 = (inp[2]) ? 4'b0001 : node21763;
														assign node21763 = (inp[13]) ? 4'b0001 : 4'b0000;
							assign node21767 = (inp[0]) ? node22147 : node21768;
								assign node21768 = (inp[2]) ? node21956 : node21769;
									assign node21769 = (inp[15]) ? node21839 : node21770;
										assign node21770 = (inp[4]) ? node21804 : node21771;
											assign node21771 = (inp[1]) ? node21785 : node21772;
												assign node21772 = (inp[5]) ? node21780 : node21773;
													assign node21773 = (inp[12]) ? node21775 : 4'b0001;
														assign node21775 = (inp[7]) ? node21777 : 4'b0001;
															assign node21777 = (inp[13]) ? 4'b0100 : 4'b0101;
													assign node21780 = (inp[7]) ? node21782 : 4'b0101;
														assign node21782 = (inp[12]) ? 4'b0001 : 4'b0100;
												assign node21785 = (inp[5]) ? node21791 : node21786;
													assign node21786 = (inp[12]) ? node21788 : 4'b0101;
														assign node21788 = (inp[7]) ? 4'b0001 : 4'b0100;
													assign node21791 = (inp[12]) ? node21799 : node21792;
														assign node21792 = (inp[13]) ? node21796 : node21793;
															assign node21793 = (inp[7]) ? 4'b0000 : 4'b0001;
															assign node21796 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node21799 = (inp[7]) ? 4'b0100 : node21800;
															assign node21800 = (inp[13]) ? 4'b0001 : 4'b0000;
											assign node21804 = (inp[1]) ? node21826 : node21805;
												assign node21805 = (inp[5]) ? node21811 : node21806;
													assign node21806 = (inp[12]) ? node21808 : 4'b0011;
														assign node21808 = (inp[7]) ? 4'b0010 : 4'b0111;
													assign node21811 = (inp[12]) ? node21821 : node21812;
														assign node21812 = (inp[9]) ? node21814 : 4'b0111;
															assign node21814 = (inp[7]) ? node21818 : node21815;
																assign node21815 = (inp[13]) ? 4'b0110 : 4'b0111;
																assign node21818 = (inp[13]) ? 4'b0111 : 4'b0110;
														assign node21821 = (inp[7]) ? node21823 : 4'b0010;
															assign node21823 = (inp[13]) ? 4'b0110 : 4'b0111;
												assign node21826 = (inp[5]) ? node21834 : node21827;
													assign node21827 = (inp[7]) ? 4'b0111 : node21828;
														assign node21828 = (inp[12]) ? node21830 : 4'b0111;
															assign node21830 = (inp[13]) ? 4'b0011 : 4'b0010;
													assign node21834 = (inp[7]) ? 4'b0011 : node21835;
														assign node21835 = (inp[12]) ? 4'b0111 : 4'b0010;
										assign node21839 = (inp[4]) ? node21891 : node21840;
											assign node21840 = (inp[13]) ? node21868 : node21841;
												assign node21841 = (inp[7]) ? node21853 : node21842;
													assign node21842 = (inp[1]) ? node21846 : node21843;
														assign node21843 = (inp[5]) ? 4'b0111 : 4'b0011;
														assign node21846 = (inp[5]) ? node21850 : node21847;
															assign node21847 = (inp[12]) ? 4'b0110 : 4'b0111;
															assign node21850 = (inp[12]) ? 4'b0011 : 4'b0010;
													assign node21853 = (inp[12]) ? node21861 : node21854;
														assign node21854 = (inp[5]) ? node21858 : node21855;
															assign node21855 = (inp[1]) ? 4'b0010 : 4'b0111;
															assign node21858 = (inp[1]) ? 4'b0111 : 4'b0010;
														assign node21861 = (inp[1]) ? node21865 : node21862;
															assign node21862 = (inp[5]) ? 4'b0111 : 4'b0010;
															assign node21865 = (inp[5]) ? 4'b0011 : 4'b0111;
												assign node21868 = (inp[5]) ? node21880 : node21869;
													assign node21869 = (inp[1]) ? node21873 : node21870;
														assign node21870 = (inp[7]) ? 4'b0011 : 4'b0010;
														assign node21873 = (inp[7]) ? node21877 : node21874;
															assign node21874 = (inp[12]) ? 4'b0110 : 4'b0111;
															assign node21877 = (inp[12]) ? 4'b0111 : 4'b0011;
													assign node21880 = (inp[1]) ? node21886 : node21881;
														assign node21881 = (inp[7]) ? node21883 : 4'b0110;
															assign node21883 = (inp[12]) ? 4'b0110 : 4'b0010;
														assign node21886 = (inp[12]) ? 4'b0010 : node21887;
															assign node21887 = (inp[7]) ? 4'b0110 : 4'b0011;
											assign node21891 = (inp[13]) ? node21921 : node21892;
												assign node21892 = (inp[1]) ? node21908 : node21893;
													assign node21893 = (inp[5]) ? node21901 : node21894;
														assign node21894 = (inp[12]) ? node21898 : node21895;
															assign node21895 = (inp[7]) ? 4'b0001 : 4'b0101;
															assign node21898 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node21901 = (inp[7]) ? node21905 : node21902;
															assign node21902 = (inp[12]) ? 4'b0100 : 4'b0000;
															assign node21905 = (inp[12]) ? 4'b0100 : 4'b0101;
													assign node21908 = (inp[5]) ? node21916 : node21909;
														assign node21909 = (inp[12]) ? node21913 : node21910;
															assign node21910 = (inp[7]) ? 4'b0100 : 4'b0000;
															assign node21913 = (inp[7]) ? 4'b0100 : 4'b0101;
														assign node21916 = (inp[7]) ? 4'b0000 : node21917;
															assign node21917 = (inp[12]) ? 4'b0000 : 4'b0100;
												assign node21921 = (inp[5]) ? node21937 : node21922;
													assign node21922 = (inp[1]) ? node21930 : node21923;
														assign node21923 = (inp[7]) ? node21927 : node21924;
															assign node21924 = (inp[12]) ? 4'b0001 : 4'b0100;
															assign node21927 = (inp[12]) ? 4'b0000 : 4'b0001;
														assign node21930 = (inp[12]) ? node21934 : node21931;
															assign node21931 = (inp[7]) ? 4'b0101 : 4'b0001;
															assign node21934 = (inp[7]) ? 4'b0101 : 4'b0100;
													assign node21937 = (inp[12]) ? node21953 : node21938;
														assign node21938 = (inp[9]) ? node21946 : node21939;
															assign node21939 = (inp[1]) ? node21943 : node21940;
																assign node21940 = (inp[7]) ? 4'b0100 : 4'b0001;
																assign node21943 = (inp[7]) ? 4'b0001 : 4'b0100;
															assign node21946 = (inp[7]) ? node21950 : node21947;
																assign node21947 = (inp[1]) ? 4'b0100 : 4'b0001;
																assign node21950 = (inp[1]) ? 4'b0001 : 4'b0100;
														assign node21953 = (inp[1]) ? 4'b0001 : 4'b0101;
									assign node21956 = (inp[15]) ? node22066 : node21957;
										assign node21957 = (inp[4]) ? node22011 : node21958;
											assign node21958 = (inp[13]) ? node21986 : node21959;
												assign node21959 = (inp[5]) ? node21973 : node21960;
													assign node21960 = (inp[1]) ? node21966 : node21961;
														assign node21961 = (inp[12]) ? node21963 : 4'b0001;
															assign node21963 = (inp[7]) ? 4'b0100 : 4'b0001;
														assign node21966 = (inp[7]) ? node21970 : node21967;
															assign node21967 = (inp[12]) ? 4'b0100 : 4'b0101;
															assign node21970 = (inp[12]) ? 4'b0001 : 4'b0101;
													assign node21973 = (inp[1]) ? node21979 : node21974;
														assign node21974 = (inp[12]) ? node21976 : 4'b0100;
															assign node21976 = (inp[7]) ? 4'b0001 : 4'b0101;
														assign node21979 = (inp[12]) ? node21983 : node21980;
															assign node21980 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node21983 = (inp[7]) ? 4'b0100 : 4'b0001;
												assign node21986 = (inp[1]) ? node21998 : node21987;
													assign node21987 = (inp[5]) ? node21993 : node21988;
														assign node21988 = (inp[12]) ? node21990 : 4'b0000;
															assign node21990 = (inp[7]) ? 4'b0100 : 4'b0000;
														assign node21993 = (inp[7]) ? node21995 : 4'b0100;
															assign node21995 = (inp[12]) ? 4'b0000 : 4'b0101;
													assign node21998 = (inp[5]) ? node22004 : node21999;
														assign node21999 = (inp[12]) ? node22001 : 4'b0100;
															assign node22001 = (inp[7]) ? 4'b0000 : 4'b0101;
														assign node22004 = (inp[12]) ? node22008 : node22005;
															assign node22005 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node22008 = (inp[7]) ? 4'b0101 : 4'b0001;
											assign node22011 = (inp[13]) ? node22041 : node22012;
												assign node22012 = (inp[5]) ? node22026 : node22013;
													assign node22013 = (inp[1]) ? node22021 : node22014;
														assign node22014 = (inp[7]) ? node22018 : node22015;
															assign node22015 = (inp[12]) ? 4'b0110 : 4'b0010;
															assign node22018 = (inp[12]) ? 4'b0011 : 4'b0010;
														assign node22021 = (inp[12]) ? node22023 : 4'b0110;
															assign node22023 = (inp[7]) ? 4'b0110 : 4'b0010;
													assign node22026 = (inp[1]) ? node22034 : node22027;
														assign node22027 = (inp[7]) ? node22031 : node22028;
															assign node22028 = (inp[12]) ? 4'b0011 : 4'b0111;
															assign node22031 = (inp[12]) ? 4'b0111 : 4'b0110;
														assign node22034 = (inp[12]) ? node22038 : node22035;
															assign node22035 = (inp[7]) ? 4'b0010 : 4'b0011;
															assign node22038 = (inp[7]) ? 4'b0010 : 4'b0110;
												assign node22041 = (inp[5]) ? node22053 : node22042;
													assign node22042 = (inp[1]) ? node22048 : node22043;
														assign node22043 = (inp[12]) ? node22045 : 4'b0011;
															assign node22045 = (inp[7]) ? 4'b0010 : 4'b0111;
														assign node22048 = (inp[7]) ? 4'b0111 : node22049;
															assign node22049 = (inp[12]) ? 4'b0010 : 4'b0111;
													assign node22053 = (inp[1]) ? node22061 : node22054;
														assign node22054 = (inp[12]) ? node22058 : node22055;
															assign node22055 = (inp[7]) ? 4'b0110 : 4'b0111;
															assign node22058 = (inp[7]) ? 4'b0111 : 4'b0010;
														assign node22061 = (inp[7]) ? 4'b0011 : node22062;
															assign node22062 = (inp[12]) ? 4'b0111 : 4'b0010;
										assign node22066 = (inp[4]) ? node22104 : node22067;
											assign node22067 = (inp[5]) ? node22089 : node22068;
												assign node22068 = (inp[1]) ? node22076 : node22069;
													assign node22069 = (inp[12]) ? node22073 : node22070;
														assign node22070 = (inp[7]) ? 4'b0111 : 4'b0011;
														assign node22073 = (inp[7]) ? 4'b0010 : 4'b0011;
													assign node22076 = (inp[7]) ? node22084 : node22077;
														assign node22077 = (inp[12]) ? node22081 : node22078;
															assign node22078 = (inp[13]) ? 4'b0111 : 4'b0110;
															assign node22081 = (inp[13]) ? 4'b0110 : 4'b0111;
														assign node22084 = (inp[12]) ? node22086 : 4'b0010;
															assign node22086 = (inp[13]) ? 4'b0111 : 4'b0110;
												assign node22089 = (inp[1]) ? node22097 : node22090;
													assign node22090 = (inp[12]) ? 4'b0111 : node22091;
														assign node22091 = (inp[7]) ? node22093 : 4'b0111;
															assign node22093 = (inp[13]) ? 4'b0010 : 4'b0011;
													assign node22097 = (inp[7]) ? node22101 : node22098;
														assign node22098 = (inp[12]) ? 4'b0011 : 4'b0010;
														assign node22101 = (inp[12]) ? 4'b0011 : 4'b0111;
											assign node22104 = (inp[1]) ? node22132 : node22105;
												assign node22105 = (inp[5]) ? node22125 : node22106;
													assign node22106 = (inp[12]) ? node22112 : node22107;
														assign node22107 = (inp[7]) ? node22109 : 4'b0100;
															assign node22109 = (inp[13]) ? 4'b0000 : 4'b0001;
														assign node22112 = (inp[9]) ? node22118 : node22113;
															assign node22113 = (inp[7]) ? 4'b0000 : node22114;
																assign node22114 = (inp[13]) ? 4'b0000 : 4'b0001;
															assign node22118 = (inp[13]) ? node22122 : node22119;
																assign node22119 = (inp[7]) ? 4'b0000 : 4'b0001;
																assign node22122 = (inp[7]) ? 4'b0001 : 4'b0000;
													assign node22125 = (inp[7]) ? node22129 : node22126;
														assign node22126 = (inp[12]) ? 4'b0101 : 4'b0001;
														assign node22129 = (inp[12]) ? 4'b0101 : 4'b0100;
												assign node22132 = (inp[5]) ? node22140 : node22133;
													assign node22133 = (inp[12]) ? node22137 : node22134;
														assign node22134 = (inp[7]) ? 4'b0101 : 4'b0001;
														assign node22137 = (inp[7]) ? 4'b0101 : 4'b0100;
													assign node22140 = (inp[12]) ? 4'b0001 : node22141;
														assign node22141 = (inp[7]) ? 4'b0001 : node22142;
															assign node22142 = (inp[13]) ? 4'b0101 : 4'b0100;
								assign node22147 = (inp[1]) ? node22311 : node22148;
									assign node22148 = (inp[5]) ? node22228 : node22149;
										assign node22149 = (inp[13]) ? node22185 : node22150;
											assign node22150 = (inp[12]) ? node22164 : node22151;
												assign node22151 = (inp[15]) ? node22157 : node22152;
													assign node22152 = (inp[4]) ? node22154 : 4'b0000;
														assign node22154 = (inp[2]) ? 4'b0011 : 4'b0010;
													assign node22157 = (inp[4]) ? node22161 : node22158;
														assign node22158 = (inp[7]) ? 4'b0110 : 4'b0010;
														assign node22161 = (inp[7]) ? 4'b0000 : 4'b0100;
												assign node22164 = (inp[7]) ? node22174 : node22165;
													assign node22165 = (inp[4]) ? node22169 : node22166;
														assign node22166 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node22169 = (inp[15]) ? 4'b0000 : node22170;
															assign node22170 = (inp[2]) ? 4'b0111 : 4'b0110;
													assign node22174 = (inp[15]) ? node22182 : node22175;
														assign node22175 = (inp[4]) ? node22179 : node22176;
															assign node22176 = (inp[2]) ? 4'b0101 : 4'b0100;
															assign node22179 = (inp[2]) ? 4'b0010 : 4'b0011;
														assign node22182 = (inp[4]) ? 4'b0001 : 4'b0011;
											assign node22185 = (inp[4]) ? node22209 : node22186;
												assign node22186 = (inp[15]) ? node22198 : node22187;
													assign node22187 = (inp[2]) ? node22193 : node22188;
														assign node22188 = (inp[7]) ? node22190 : 4'b0000;
															assign node22190 = (inp[12]) ? 4'b0101 : 4'b0000;
														assign node22193 = (inp[7]) ? node22195 : 4'b0001;
															assign node22195 = (inp[12]) ? 4'b0101 : 4'b0001;
													assign node22198 = (inp[2]) ? node22204 : node22199;
														assign node22199 = (inp[7]) ? node22201 : 4'b0011;
															assign node22201 = (inp[12]) ? 4'b0010 : 4'b0111;
														assign node22204 = (inp[7]) ? node22206 : 4'b0010;
															assign node22206 = (inp[12]) ? 4'b0011 : 4'b0110;
												assign node22209 = (inp[15]) ? node22215 : node22210;
													assign node22210 = (inp[12]) ? node22212 : 4'b0010;
														assign node22212 = (inp[7]) ? 4'b0011 : 4'b0110;
													assign node22215 = (inp[12]) ? node22221 : node22216;
														assign node22216 = (inp[7]) ? node22218 : 4'b0101;
															assign node22218 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node22221 = (inp[7]) ? node22225 : node22222;
															assign node22222 = (inp[2]) ? 4'b0001 : 4'b0000;
															assign node22225 = (inp[2]) ? 4'b0000 : 4'b0001;
										assign node22228 = (inp[7]) ? node22264 : node22229;
											assign node22229 = (inp[4]) ? node22241 : node22230;
												assign node22230 = (inp[15]) ? node22236 : node22231;
													assign node22231 = (inp[2]) ? node22233 : 4'b0100;
														assign node22233 = (inp[13]) ? 4'b0101 : 4'b0100;
													assign node22236 = (inp[2]) ? 4'b0110 : node22237;
														assign node22237 = (inp[13]) ? 4'b0111 : 4'b0110;
												assign node22241 = (inp[15]) ? node22253 : node22242;
													assign node22242 = (inp[12]) ? node22248 : node22243;
														assign node22243 = (inp[13]) ? node22245 : 4'b0110;
															assign node22245 = (inp[2]) ? 4'b0110 : 4'b0111;
														assign node22248 = (inp[13]) ? 4'b0011 : node22249;
															assign node22249 = (inp[2]) ? 4'b0010 : 4'b0011;
													assign node22253 = (inp[12]) ? node22259 : node22254;
														assign node22254 = (inp[2]) ? 4'b0000 : node22255;
															assign node22255 = (inp[13]) ? 4'b0000 : 4'b0001;
														assign node22259 = (inp[2]) ? 4'b0100 : node22260;
															assign node22260 = (inp[13]) ? 4'b0100 : 4'b0101;
											assign node22264 = (inp[12]) ? node22288 : node22265;
												assign node22265 = (inp[15]) ? node22277 : node22266;
													assign node22266 = (inp[4]) ? node22272 : node22267;
														assign node22267 = (inp[2]) ? node22269 : 4'b0101;
															assign node22269 = (inp[13]) ? 4'b0100 : 4'b0101;
														assign node22272 = (inp[2]) ? 4'b0111 : node22273;
															assign node22273 = (inp[13]) ? 4'b0110 : 4'b0111;
													assign node22277 = (inp[4]) ? node22283 : node22278;
														assign node22278 = (inp[13]) ? 4'b0011 : node22279;
															assign node22279 = (inp[2]) ? 4'b0010 : 4'b0011;
														assign node22283 = (inp[13]) ? 4'b0101 : node22284;
															assign node22284 = (inp[2]) ? 4'b0101 : 4'b0100;
												assign node22288 = (inp[15]) ? node22300 : node22289;
													assign node22289 = (inp[4]) ? node22295 : node22290;
														assign node22290 = (inp[2]) ? node22292 : 4'b0000;
															assign node22292 = (inp[13]) ? 4'b0001 : 4'b0000;
														assign node22295 = (inp[13]) ? node22297 : 4'b0110;
															assign node22297 = (inp[2]) ? 4'b0110 : 4'b0111;
													assign node22300 = (inp[4]) ? node22306 : node22301;
														assign node22301 = (inp[13]) ? node22303 : 4'b0110;
															assign node22303 = (inp[2]) ? 4'b0110 : 4'b0111;
														assign node22306 = (inp[13]) ? 4'b0100 : node22307;
															assign node22307 = (inp[2]) ? 4'b0100 : 4'b0101;
									assign node22311 = (inp[5]) ? node22391 : node22312;
										assign node22312 = (inp[12]) ? node22344 : node22313;
											assign node22313 = (inp[15]) ? node22325 : node22314;
												assign node22314 = (inp[4]) ? node22320 : node22315;
													assign node22315 = (inp[2]) ? node22317 : 4'b0100;
														assign node22317 = (inp[13]) ? 4'b0101 : 4'b0100;
													assign node22320 = (inp[2]) ? node22322 : 4'b0110;
														assign node22322 = (inp[13]) ? 4'b0110 : 4'b0111;
												assign node22325 = (inp[4]) ? node22337 : node22326;
													assign node22326 = (inp[7]) ? node22332 : node22327;
														assign node22327 = (inp[2]) ? node22329 : 4'b0110;
															assign node22329 = (inp[13]) ? 4'b0110 : 4'b0111;
														assign node22332 = (inp[13]) ? node22334 : 4'b0011;
															assign node22334 = (inp[2]) ? 4'b0011 : 4'b0010;
													assign node22337 = (inp[7]) ? node22339 : 4'b0000;
														assign node22339 = (inp[13]) ? 4'b0100 : node22340;
															assign node22340 = (inp[2]) ? 4'b0100 : 4'b0101;
											assign node22344 = (inp[7]) ? node22368 : node22345;
												assign node22345 = (inp[15]) ? node22357 : node22346;
													assign node22346 = (inp[4]) ? node22352 : node22347;
														assign node22347 = (inp[2]) ? node22349 : 4'b0101;
															assign node22349 = (inp[13]) ? 4'b0100 : 4'b0101;
														assign node22352 = (inp[2]) ? 4'b0011 : node22353;
															assign node22353 = (inp[13]) ? 4'b0010 : 4'b0011;
													assign node22357 = (inp[4]) ? node22363 : node22358;
														assign node22358 = (inp[13]) ? 4'b0111 : node22359;
															assign node22359 = (inp[2]) ? 4'b0110 : 4'b0111;
														assign node22363 = (inp[2]) ? 4'b0101 : node22364;
															assign node22364 = (inp[13]) ? 4'b0101 : 4'b0100;
												assign node22368 = (inp[15]) ? node22380 : node22369;
													assign node22369 = (inp[4]) ? node22375 : node22370;
														assign node22370 = (inp[2]) ? node22372 : 4'b0000;
															assign node22372 = (inp[13]) ? 4'b0001 : 4'b0000;
														assign node22375 = (inp[2]) ? node22377 : 4'b0110;
															assign node22377 = (inp[13]) ? 4'b0110 : 4'b0111;
													assign node22380 = (inp[4]) ? node22386 : node22381;
														assign node22381 = (inp[13]) ? 4'b0110 : node22382;
															assign node22382 = (inp[2]) ? 4'b0111 : 4'b0110;
														assign node22386 = (inp[13]) ? 4'b0100 : node22387;
															assign node22387 = (inp[2]) ? 4'b0100 : 4'b0101;
										assign node22391 = (inp[2]) ? node22445 : node22392;
											assign node22392 = (inp[13]) ? node22418 : node22393;
												assign node22393 = (inp[4]) ? node22409 : node22394;
													assign node22394 = (inp[15]) ? node22402 : node22395;
														assign node22395 = (inp[7]) ? node22399 : node22396;
															assign node22396 = (inp[12]) ? 4'b0001 : 4'b0000;
															assign node22399 = (inp[12]) ? 4'b0101 : 4'b0001;
														assign node22402 = (inp[7]) ? node22406 : node22403;
															assign node22403 = (inp[12]) ? 4'b0010 : 4'b0011;
															assign node22406 = (inp[12]) ? 4'b0010 : 4'b0110;
													assign node22409 = (inp[15]) ? node22413 : node22410;
														assign node22410 = (inp[7]) ? 4'b0010 : 4'b0011;
														assign node22413 = (inp[12]) ? 4'b0001 : node22414;
															assign node22414 = (inp[7]) ? 4'b0001 : 4'b0101;
												assign node22418 = (inp[4]) ? node22432 : node22419;
													assign node22419 = (inp[15]) ? node22427 : node22420;
														assign node22420 = (inp[7]) ? node22424 : node22421;
															assign node22421 = (inp[12]) ? 4'b0000 : 4'b0001;
															assign node22424 = (inp[12]) ? 4'b0101 : 4'b0000;
														assign node22427 = (inp[12]) ? 4'b0011 : node22428;
															assign node22428 = (inp[7]) ? 4'b0111 : 4'b0010;
													assign node22432 = (inp[15]) ? node22440 : node22433;
														assign node22433 = (inp[12]) ? node22437 : node22434;
															assign node22434 = (inp[7]) ? 4'b0010 : 4'b0011;
															assign node22437 = (inp[7]) ? 4'b0010 : 4'b0110;
														assign node22440 = (inp[12]) ? 4'b0000 : node22441;
															assign node22441 = (inp[7]) ? 4'b0000 : 4'b0101;
											assign node22445 = (inp[15]) ? node22471 : node22446;
												assign node22446 = (inp[4]) ? node22456 : node22447;
													assign node22447 = (inp[12]) ? node22451 : node22448;
														assign node22448 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node22451 = (inp[7]) ? node22453 : 4'b0000;
															assign node22453 = (inp[13]) ? 4'b0100 : 4'b0101;
													assign node22456 = (inp[12]) ? node22464 : node22457;
														assign node22457 = (inp[7]) ? node22461 : node22458;
															assign node22458 = (inp[13]) ? 4'b0011 : 4'b0010;
															assign node22461 = (inp[13]) ? 4'b0010 : 4'b0011;
														assign node22464 = (inp[7]) ? node22468 : node22465;
															assign node22465 = (inp[13]) ? 4'b0110 : 4'b0111;
															assign node22468 = (inp[13]) ? 4'b0010 : 4'b0011;
												assign node22471 = (inp[4]) ? node22477 : node22472;
													assign node22472 = (inp[12]) ? 4'b0010 : node22473;
														assign node22473 = (inp[7]) ? 4'b0110 : 4'b0011;
													assign node22477 = (inp[12]) ? 4'b0000 : node22478;
														assign node22478 = (inp[7]) ? 4'b0000 : node22479;
															assign node22479 = (inp[13]) ? 4'b0100 : 4'b0101;
						assign node22484 = (inp[1]) ? node23486 : node22485;
							assign node22485 = (inp[5]) ? node22857 : node22486;
								assign node22486 = (inp[0]) ? node22686 : node22487;
									assign node22487 = (inp[11]) ? node22579 : node22488;
										assign node22488 = (inp[13]) ? node22526 : node22489;
											assign node22489 = (inp[12]) ? node22505 : node22490;
												assign node22490 = (inp[15]) ? node22496 : node22491;
													assign node22491 = (inp[4]) ? node22493 : 4'b0000;
														assign node22493 = (inp[2]) ? 4'b0011 : 4'b0010;
													assign node22496 = (inp[4]) ? node22500 : node22497;
														assign node22497 = (inp[7]) ? 4'b0110 : 4'b0010;
														assign node22500 = (inp[7]) ? 4'b0000 : node22501;
															assign node22501 = (inp[2]) ? 4'b0101 : 4'b0100;
												assign node22505 = (inp[7]) ? node22515 : node22506;
													assign node22506 = (inp[15]) ? node22512 : node22507;
														assign node22507 = (inp[4]) ? node22509 : 4'b0000;
															assign node22509 = (inp[2]) ? 4'b0111 : 4'b0110;
														assign node22512 = (inp[4]) ? 4'b0000 : 4'b0010;
													assign node22515 = (inp[15]) ? node22523 : node22516;
														assign node22516 = (inp[4]) ? node22520 : node22517;
															assign node22517 = (inp[2]) ? 4'b0101 : 4'b0100;
															assign node22520 = (inp[2]) ? 4'b0010 : 4'b0011;
														assign node22523 = (inp[4]) ? 4'b0001 : 4'b0011;
											assign node22526 = (inp[4]) ? node22550 : node22527;
												assign node22527 = (inp[15]) ? node22539 : node22528;
													assign node22528 = (inp[2]) ? node22534 : node22529;
														assign node22529 = (inp[12]) ? node22531 : 4'b0000;
															assign node22531 = (inp[7]) ? 4'b0101 : 4'b0000;
														assign node22534 = (inp[12]) ? node22536 : 4'b0001;
															assign node22536 = (inp[7]) ? 4'b0101 : 4'b0001;
													assign node22539 = (inp[7]) ? node22543 : node22540;
														assign node22540 = (inp[2]) ? 4'b0010 : 4'b0011;
														assign node22543 = (inp[12]) ? node22547 : node22544;
															assign node22544 = (inp[2]) ? 4'b0110 : 4'b0111;
															assign node22547 = (inp[2]) ? 4'b0011 : 4'b0010;
												assign node22550 = (inp[15]) ? node22558 : node22551;
													assign node22551 = (inp[7]) ? node22555 : node22552;
														assign node22552 = (inp[12]) ? 4'b0110 : 4'b0010;
														assign node22555 = (inp[12]) ? 4'b0011 : 4'b0010;
													assign node22558 = (inp[7]) ? node22564 : node22559;
														assign node22559 = (inp[12]) ? node22561 : 4'b0101;
															assign node22561 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node22564 = (inp[9]) ? node22572 : node22565;
															assign node22565 = (inp[2]) ? node22569 : node22566;
																assign node22566 = (inp[12]) ? 4'b0001 : 4'b0000;
																assign node22569 = (inp[12]) ? 4'b0000 : 4'b0001;
															assign node22572 = (inp[12]) ? node22576 : node22573;
																assign node22573 = (inp[2]) ? 4'b0001 : 4'b0000;
																assign node22576 = (inp[2]) ? 4'b0000 : 4'b0001;
										assign node22579 = (inp[13]) ? node22635 : node22580;
											assign node22580 = (inp[2]) ? node22608 : node22581;
												assign node22581 = (inp[7]) ? node22593 : node22582;
													assign node22582 = (inp[4]) ? node22586 : node22583;
														assign node22583 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node22586 = (inp[15]) ? node22590 : node22587;
															assign node22587 = (inp[12]) ? 4'b0111 : 4'b0011;
															assign node22590 = (inp[12]) ? 4'b0001 : 4'b0101;
													assign node22593 = (inp[4]) ? node22601 : node22594;
														assign node22594 = (inp[15]) ? node22598 : node22595;
															assign node22595 = (inp[12]) ? 4'b0101 : 4'b0001;
															assign node22598 = (inp[12]) ? 4'b0010 : 4'b0111;
														assign node22601 = (inp[12]) ? node22605 : node22602;
															assign node22602 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node22605 = (inp[15]) ? 4'b0000 : 4'b0010;
												assign node22608 = (inp[4]) ? node22620 : node22609;
													assign node22609 = (inp[15]) ? node22615 : node22610;
														assign node22610 = (inp[7]) ? node22612 : 4'b0001;
															assign node22612 = (inp[12]) ? 4'b0100 : 4'b0001;
														assign node22615 = (inp[7]) ? node22617 : 4'b0011;
															assign node22617 = (inp[12]) ? 4'b0010 : 4'b0111;
													assign node22620 = (inp[15]) ? node22628 : node22621;
														assign node22621 = (inp[7]) ? node22625 : node22622;
															assign node22622 = (inp[12]) ? 4'b0110 : 4'b0010;
															assign node22625 = (inp[12]) ? 4'b0011 : 4'b0010;
														assign node22628 = (inp[7]) ? node22632 : node22629;
															assign node22629 = (inp[12]) ? 4'b0001 : 4'b0100;
															assign node22632 = (inp[12]) ? 4'b0000 : 4'b0001;
											assign node22635 = (inp[15]) ? node22653 : node22636;
												assign node22636 = (inp[4]) ? node22648 : node22637;
													assign node22637 = (inp[2]) ? node22643 : node22638;
														assign node22638 = (inp[12]) ? node22640 : 4'b0001;
															assign node22640 = (inp[7]) ? 4'b0100 : 4'b0001;
														assign node22643 = (inp[12]) ? node22645 : 4'b0000;
															assign node22645 = (inp[7]) ? 4'b0100 : 4'b0000;
													assign node22648 = (inp[12]) ? node22650 : 4'b0011;
														assign node22650 = (inp[7]) ? 4'b0010 : 4'b0111;
												assign node22653 = (inp[4]) ? node22665 : node22654;
													assign node22654 = (inp[2]) ? node22660 : node22655;
														assign node22655 = (inp[7]) ? node22657 : 4'b0010;
															assign node22657 = (inp[12]) ? 4'b0011 : 4'b0110;
														assign node22660 = (inp[7]) ? node22662 : 4'b0011;
															assign node22662 = (inp[12]) ? 4'b0010 : 4'b0111;
													assign node22665 = (inp[12]) ? node22671 : node22666;
														assign node22666 = (inp[7]) ? node22668 : 4'b0100;
															assign node22668 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node22671 = (inp[9]) ? node22679 : node22672;
															assign node22672 = (inp[2]) ? node22676 : node22673;
																assign node22673 = (inp[7]) ? 4'b0000 : 4'b0001;
																assign node22676 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node22679 = (inp[7]) ? node22683 : node22680;
																assign node22680 = (inp[2]) ? 4'b0000 : 4'b0001;
																assign node22683 = (inp[2]) ? 4'b0001 : 4'b0000;
									assign node22686 = (inp[11]) ? node22772 : node22687;
										assign node22687 = (inp[13]) ? node22727 : node22688;
											assign node22688 = (inp[4]) ? node22702 : node22689;
												assign node22689 = (inp[15]) ? node22697 : node22690;
													assign node22690 = (inp[7]) ? node22692 : 4'b0001;
														assign node22692 = (inp[12]) ? node22694 : 4'b0001;
															assign node22694 = (inp[2]) ? 4'b0100 : 4'b0101;
													assign node22697 = (inp[7]) ? node22699 : 4'b0011;
														assign node22699 = (inp[12]) ? 4'b0010 : 4'b0111;
												assign node22702 = (inp[15]) ? node22718 : node22703;
													assign node22703 = (inp[7]) ? node22711 : node22704;
														assign node22704 = (inp[2]) ? node22708 : node22705;
															assign node22705 = (inp[12]) ? 4'b0111 : 4'b0011;
															assign node22708 = (inp[12]) ? 4'b0110 : 4'b0010;
														assign node22711 = (inp[2]) ? node22715 : node22712;
															assign node22712 = (inp[12]) ? 4'b0010 : 4'b0011;
															assign node22715 = (inp[12]) ? 4'b0011 : 4'b0010;
													assign node22718 = (inp[12]) ? node22724 : node22719;
														assign node22719 = (inp[7]) ? 4'b0001 : node22720;
															assign node22720 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node22724 = (inp[7]) ? 4'b0000 : 4'b0001;
											assign node22727 = (inp[12]) ? node22747 : node22728;
												assign node22728 = (inp[15]) ? node22734 : node22729;
													assign node22729 = (inp[4]) ? 4'b0011 : node22730;
														assign node22730 = (inp[2]) ? 4'b0000 : 4'b0001;
													assign node22734 = (inp[4]) ? node22742 : node22735;
														assign node22735 = (inp[2]) ? node22739 : node22736;
															assign node22736 = (inp[7]) ? 4'b0110 : 4'b0010;
															assign node22739 = (inp[7]) ? 4'b0111 : 4'b0011;
														assign node22742 = (inp[7]) ? node22744 : 4'b0100;
															assign node22744 = (inp[2]) ? 4'b0000 : 4'b0001;
												assign node22747 = (inp[15]) ? node22757 : node22748;
													assign node22748 = (inp[4]) ? node22754 : node22749;
														assign node22749 = (inp[7]) ? 4'b0100 : node22750;
															assign node22750 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node22754 = (inp[7]) ? 4'b0010 : 4'b0111;
													assign node22757 = (inp[4]) ? node22765 : node22758;
														assign node22758 = (inp[2]) ? node22762 : node22759;
															assign node22759 = (inp[7]) ? 4'b0011 : 4'b0010;
															assign node22762 = (inp[7]) ? 4'b0010 : 4'b0011;
														assign node22765 = (inp[7]) ? node22769 : node22766;
															assign node22766 = (inp[2]) ? 4'b0000 : 4'b0001;
															assign node22769 = (inp[2]) ? 4'b0001 : 4'b0000;
										assign node22772 = (inp[13]) ? node22808 : node22773;
											assign node22773 = (inp[12]) ? node22789 : node22774;
												assign node22774 = (inp[15]) ? node22780 : node22775;
													assign node22775 = (inp[4]) ? node22777 : 4'b0000;
														assign node22777 = (inp[2]) ? 4'b0011 : 4'b0010;
													assign node22780 = (inp[4]) ? node22784 : node22781;
														assign node22781 = (inp[7]) ? 4'b0110 : 4'b0010;
														assign node22784 = (inp[7]) ? 4'b0000 : node22785;
															assign node22785 = (inp[2]) ? 4'b0101 : 4'b0100;
												assign node22789 = (inp[7]) ? node22799 : node22790;
													assign node22790 = (inp[15]) ? node22796 : node22791;
														assign node22791 = (inp[4]) ? node22793 : 4'b0000;
															assign node22793 = (inp[2]) ? 4'b0111 : 4'b0110;
														assign node22796 = (inp[4]) ? 4'b0000 : 4'b0010;
													assign node22799 = (inp[15]) ? node22805 : node22800;
														assign node22800 = (inp[4]) ? node22802 : 4'b0100;
															assign node22802 = (inp[2]) ? 4'b0010 : 4'b0011;
														assign node22805 = (inp[4]) ? 4'b0001 : 4'b0011;
											assign node22808 = (inp[2]) ? node22834 : node22809;
												assign node22809 = (inp[15]) ? node22821 : node22810;
													assign node22810 = (inp[4]) ? node22816 : node22811;
														assign node22811 = (inp[7]) ? node22813 : 4'b0000;
															assign node22813 = (inp[12]) ? 4'b0101 : 4'b0000;
														assign node22816 = (inp[12]) ? node22818 : 4'b0010;
															assign node22818 = (inp[7]) ? 4'b0011 : 4'b0110;
													assign node22821 = (inp[4]) ? node22827 : node22822;
														assign node22822 = (inp[7]) ? node22824 : 4'b0011;
															assign node22824 = (inp[12]) ? 4'b0010 : 4'b0111;
														assign node22827 = (inp[7]) ? node22831 : node22828;
															assign node22828 = (inp[12]) ? 4'b0000 : 4'b0101;
															assign node22831 = (inp[12]) ? 4'b0001 : 4'b0000;
												assign node22834 = (inp[15]) ? node22846 : node22835;
													assign node22835 = (inp[4]) ? node22841 : node22836;
														assign node22836 = (inp[7]) ? node22838 : 4'b0001;
															assign node22838 = (inp[12]) ? 4'b0101 : 4'b0001;
														assign node22841 = (inp[7]) ? node22843 : 4'b0110;
															assign node22843 = (inp[12]) ? 4'b0011 : 4'b0010;
													assign node22846 = (inp[4]) ? node22852 : node22847;
														assign node22847 = (inp[12]) ? node22849 : 4'b0110;
															assign node22849 = (inp[7]) ? 4'b0011 : 4'b0010;
														assign node22852 = (inp[12]) ? node22854 : 4'b0001;
															assign node22854 = (inp[7]) ? 4'b0000 : 4'b0001;
								assign node22857 = (inp[13]) ? node23097 : node22858;
									assign node22858 = (inp[7]) ? node22976 : node22859;
										assign node22859 = (inp[4]) ? node22891 : node22860;
											assign node22860 = (inp[15]) ? node22884 : node22861;
												assign node22861 = (inp[12]) ? node22869 : node22862;
													assign node22862 = (inp[11]) ? node22866 : node22863;
														assign node22863 = (inp[0]) ? 4'b0101 : 4'b0100;
														assign node22866 = (inp[0]) ? 4'b0100 : 4'b0101;
													assign node22869 = (inp[9]) ? node22877 : node22870;
														assign node22870 = (inp[0]) ? node22874 : node22871;
															assign node22871 = (inp[11]) ? 4'b0101 : 4'b0100;
															assign node22874 = (inp[11]) ? 4'b0100 : 4'b0101;
														assign node22877 = (inp[0]) ? node22881 : node22878;
															assign node22878 = (inp[11]) ? 4'b0101 : 4'b0100;
															assign node22881 = (inp[11]) ? 4'b0100 : 4'b0101;
												assign node22884 = (inp[11]) ? node22888 : node22885;
													assign node22885 = (inp[0]) ? 4'b0111 : 4'b0110;
													assign node22888 = (inp[0]) ? 4'b0110 : 4'b0111;
											assign node22891 = (inp[15]) ? node22939 : node22892;
												assign node22892 = (inp[12]) ? node22916 : node22893;
													assign node22893 = (inp[2]) ? node22901 : node22894;
														assign node22894 = (inp[0]) ? node22898 : node22895;
															assign node22895 = (inp[11]) ? 4'b0111 : 4'b0110;
															assign node22898 = (inp[11]) ? 4'b0110 : 4'b0111;
														assign node22901 = (inp[9]) ? node22909 : node22902;
															assign node22902 = (inp[11]) ? node22906 : node22903;
																assign node22903 = (inp[0]) ? 4'b0111 : 4'b0110;
																assign node22906 = (inp[0]) ? 4'b0110 : 4'b0111;
															assign node22909 = (inp[11]) ? node22913 : node22910;
																assign node22910 = (inp[0]) ? 4'b0111 : 4'b0110;
																assign node22913 = (inp[0]) ? 4'b0110 : 4'b0111;
													assign node22916 = (inp[9]) ? node22926 : node22917;
														assign node22917 = (inp[0]) ? 4'b0011 : node22918;
															assign node22918 = (inp[11]) ? node22922 : node22919;
																assign node22919 = (inp[2]) ? 4'b0010 : 4'b0011;
																assign node22922 = (inp[2]) ? 4'b0011 : 4'b0010;
														assign node22926 = (inp[2]) ? node22934 : node22927;
															assign node22927 = (inp[11]) ? node22931 : node22928;
																assign node22928 = (inp[0]) ? 4'b0010 : 4'b0011;
																assign node22931 = (inp[0]) ? 4'b0011 : 4'b0010;
															assign node22934 = (inp[0]) ? 4'b0010 : node22935;
																assign node22935 = (inp[11]) ? 4'b0011 : 4'b0010;
												assign node22939 = (inp[12]) ? node22955 : node22940;
													assign node22940 = (inp[0]) ? node22948 : node22941;
														assign node22941 = (inp[11]) ? node22945 : node22942;
															assign node22942 = (inp[2]) ? 4'b0000 : 4'b0001;
															assign node22945 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node22948 = (inp[11]) ? node22952 : node22949;
															assign node22949 = (inp[2]) ? 4'b0001 : 4'b0000;
															assign node22952 = (inp[2]) ? 4'b0000 : 4'b0001;
													assign node22955 = (inp[2]) ? node22971 : node22956;
														assign node22956 = (inp[9]) ? node22964 : node22957;
															assign node22957 = (inp[11]) ? node22961 : node22958;
																assign node22958 = (inp[0]) ? 4'b0100 : 4'b0101;
																assign node22961 = (inp[0]) ? 4'b0101 : 4'b0100;
															assign node22964 = (inp[0]) ? node22968 : node22965;
																assign node22965 = (inp[11]) ? 4'b0100 : 4'b0101;
																assign node22968 = (inp[11]) ? 4'b0101 : 4'b0100;
														assign node22971 = (inp[0]) ? node22973 : 4'b0101;
															assign node22973 = (inp[11]) ? 4'b0100 : 4'b0101;
										assign node22976 = (inp[4]) ? node23018 : node22977;
											assign node22977 = (inp[15]) ? node22993 : node22978;
												assign node22978 = (inp[12]) ? node22986 : node22979;
													assign node22979 = (inp[0]) ? node22983 : node22980;
														assign node22980 = (inp[11]) ? 4'b0100 : 4'b0101;
														assign node22983 = (inp[11]) ? 4'b0101 : 4'b0100;
													assign node22986 = (inp[11]) ? node22990 : node22987;
														assign node22987 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node22990 = (inp[0]) ? 4'b0000 : 4'b0001;
												assign node22993 = (inp[12]) ? node23011 : node22994;
													assign node22994 = (inp[11]) ? node23004 : node22995;
														assign node22995 = (inp[9]) ? node23001 : node22996;
															assign node22996 = (inp[0]) ? 4'b0010 : node22997;
																assign node22997 = (inp[2]) ? 4'b0010 : 4'b0011;
															assign node23001 = (inp[2]) ? 4'b0011 : 4'b0010;
														assign node23004 = (inp[2]) ? node23008 : node23005;
															assign node23005 = (inp[0]) ? 4'b0011 : 4'b0010;
															assign node23008 = (inp[0]) ? 4'b0010 : 4'b0011;
													assign node23011 = (inp[11]) ? node23015 : node23012;
														assign node23012 = (inp[0]) ? 4'b0111 : 4'b0110;
														assign node23015 = (inp[0]) ? 4'b0110 : 4'b0111;
											assign node23018 = (inp[15]) ? node23048 : node23019;
												assign node23019 = (inp[0]) ? node23033 : node23020;
													assign node23020 = (inp[2]) ? node23028 : node23021;
														assign node23021 = (inp[11]) ? node23025 : node23022;
															assign node23022 = (inp[12]) ? 4'b0110 : 4'b0111;
															assign node23025 = (inp[9]) ? 4'b0111 : 4'b0110;
														assign node23028 = (inp[12]) ? node23030 : 4'b0110;
															assign node23030 = (inp[11]) ? 4'b0111 : 4'b0110;
													assign node23033 = (inp[9]) ? node23039 : node23034;
														assign node23034 = (inp[11]) ? 4'b0110 : node23035;
															assign node23035 = (inp[12]) ? 4'b0111 : 4'b0110;
														assign node23039 = (inp[2]) ? 4'b0111 : node23040;
															assign node23040 = (inp[11]) ? node23044 : node23041;
																assign node23041 = (inp[12]) ? 4'b0111 : 4'b0110;
																assign node23044 = (inp[12]) ? 4'b0110 : 4'b0111;
												assign node23048 = (inp[9]) ? node23070 : node23049;
													assign node23049 = (inp[11]) ? node23065 : node23050;
														assign node23050 = (inp[0]) ? node23058 : node23051;
															assign node23051 = (inp[2]) ? node23055 : node23052;
																assign node23052 = (inp[12]) ? 4'b0101 : 4'b0100;
																assign node23055 = (inp[12]) ? 4'b0100 : 4'b0101;
															assign node23058 = (inp[12]) ? node23062 : node23059;
																assign node23059 = (inp[2]) ? 4'b0100 : 4'b0101;
																assign node23062 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node23065 = (inp[2]) ? node23067 : 4'b0100;
															assign node23067 = (inp[12]) ? 4'b0101 : 4'b0100;
													assign node23070 = (inp[0]) ? node23084 : node23071;
														assign node23071 = (inp[11]) ? node23079 : node23072;
															assign node23072 = (inp[2]) ? node23076 : node23073;
																assign node23073 = (inp[12]) ? 4'b0101 : 4'b0100;
																assign node23076 = (inp[12]) ? 4'b0100 : 4'b0101;
															assign node23079 = (inp[12]) ? node23081 : 4'b0101;
																assign node23081 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node23084 = (inp[11]) ? node23090 : node23085;
															assign node23085 = (inp[12]) ? 4'b0101 : node23086;
																assign node23086 = (inp[2]) ? 4'b0100 : 4'b0101;
															assign node23090 = (inp[2]) ? node23094 : node23091;
																assign node23091 = (inp[12]) ? 4'b0101 : 4'b0100;
																assign node23094 = (inp[12]) ? 4'b0100 : 4'b0101;
									assign node23097 = (inp[9]) ? node23299 : node23098;
										assign node23098 = (inp[7]) ? node23200 : node23099;
											assign node23099 = (inp[4]) ? node23155 : node23100;
												assign node23100 = (inp[15]) ? node23130 : node23101;
													assign node23101 = (inp[12]) ? node23117 : node23102;
														assign node23102 = (inp[0]) ? node23110 : node23103;
															assign node23103 = (inp[11]) ? node23107 : node23104;
																assign node23104 = (inp[2]) ? 4'b0101 : 4'b0100;
																assign node23107 = (inp[2]) ? 4'b0100 : 4'b0101;
															assign node23110 = (inp[2]) ? node23114 : node23111;
																assign node23111 = (inp[11]) ? 4'b0100 : 4'b0101;
																assign node23114 = (inp[11]) ? 4'b0101 : 4'b0100;
														assign node23117 = (inp[11]) ? node23123 : node23118;
															assign node23118 = (inp[0]) ? 4'b0100 : node23119;
																assign node23119 = (inp[2]) ? 4'b0101 : 4'b0100;
															assign node23123 = (inp[0]) ? node23127 : node23124;
																assign node23124 = (inp[2]) ? 4'b0100 : 4'b0101;
																assign node23127 = (inp[2]) ? 4'b0101 : 4'b0100;
													assign node23130 = (inp[12]) ? node23146 : node23131;
														assign node23131 = (inp[0]) ? node23139 : node23132;
															assign node23132 = (inp[11]) ? node23136 : node23133;
																assign node23133 = (inp[2]) ? 4'b0110 : 4'b0111;
																assign node23136 = (inp[2]) ? 4'b0111 : 4'b0110;
															assign node23139 = (inp[11]) ? node23143 : node23140;
																assign node23140 = (inp[2]) ? 4'b0111 : 4'b0110;
																assign node23143 = (inp[2]) ? 4'b0110 : 4'b0111;
														assign node23146 = (inp[2]) ? node23148 : 4'b0111;
															assign node23148 = (inp[0]) ? node23152 : node23149;
																assign node23149 = (inp[11]) ? 4'b0111 : 4'b0110;
																assign node23152 = (inp[11]) ? 4'b0110 : 4'b0111;
												assign node23155 = (inp[15]) ? node23179 : node23156;
													assign node23156 = (inp[12]) ? node23172 : node23157;
														assign node23157 = (inp[11]) ? node23165 : node23158;
															assign node23158 = (inp[0]) ? node23162 : node23159;
																assign node23159 = (inp[2]) ? 4'b0110 : 4'b0111;
																assign node23162 = (inp[2]) ? 4'b0111 : 4'b0110;
															assign node23165 = (inp[2]) ? node23169 : node23166;
																assign node23166 = (inp[0]) ? 4'b0111 : 4'b0110;
																assign node23169 = (inp[0]) ? 4'b0110 : 4'b0111;
														assign node23172 = (inp[11]) ? node23176 : node23173;
															assign node23173 = (inp[0]) ? 4'b0010 : 4'b0011;
															assign node23176 = (inp[0]) ? 4'b0011 : 4'b0010;
													assign node23179 = (inp[12]) ? node23193 : node23180;
														assign node23180 = (inp[2]) ? node23188 : node23181;
															assign node23181 = (inp[0]) ? node23185 : node23182;
																assign node23182 = (inp[11]) ? 4'b0001 : 4'b0000;
																assign node23185 = (inp[11]) ? 4'b0000 : 4'b0001;
															assign node23188 = (inp[11]) ? 4'b0001 : node23189;
																assign node23189 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node23193 = (inp[0]) ? node23197 : node23194;
															assign node23194 = (inp[11]) ? 4'b0101 : 4'b0100;
															assign node23197 = (inp[11]) ? 4'b0100 : 4'b0101;
											assign node23200 = (inp[4]) ? node23254 : node23201;
												assign node23201 = (inp[15]) ? node23231 : node23202;
													assign node23202 = (inp[12]) ? node23216 : node23203;
														assign node23203 = (inp[0]) ? node23211 : node23204;
															assign node23204 = (inp[11]) ? node23208 : node23205;
																assign node23205 = (inp[2]) ? 4'b0100 : 4'b0101;
																assign node23208 = (inp[2]) ? 4'b0101 : 4'b0100;
															assign node23211 = (inp[2]) ? 4'b0101 : node23212;
																assign node23212 = (inp[11]) ? 4'b0101 : 4'b0100;
														assign node23216 = (inp[2]) ? node23224 : node23217;
															assign node23217 = (inp[0]) ? node23221 : node23218;
																assign node23218 = (inp[11]) ? 4'b0001 : 4'b0000;
																assign node23221 = (inp[11]) ? 4'b0000 : 4'b0001;
															assign node23224 = (inp[11]) ? node23228 : node23225;
																assign node23225 = (inp[0]) ? 4'b0000 : 4'b0001;
																assign node23228 = (inp[0]) ? 4'b0001 : 4'b0000;
													assign node23231 = (inp[12]) ? node23239 : node23232;
														assign node23232 = (inp[0]) ? node23236 : node23233;
															assign node23233 = (inp[11]) ? 4'b0010 : 4'b0011;
															assign node23236 = (inp[11]) ? 4'b0011 : 4'b0010;
														assign node23239 = (inp[11]) ? node23247 : node23240;
															assign node23240 = (inp[0]) ? node23244 : node23241;
																assign node23241 = (inp[2]) ? 4'b0110 : 4'b0111;
																assign node23244 = (inp[2]) ? 4'b0111 : 4'b0110;
															assign node23247 = (inp[0]) ? node23251 : node23248;
																assign node23248 = (inp[2]) ? 4'b0111 : 4'b0110;
																assign node23251 = (inp[2]) ? 4'b0110 : 4'b0111;
												assign node23254 = (inp[15]) ? node23280 : node23255;
													assign node23255 = (inp[2]) ? node23271 : node23256;
														assign node23256 = (inp[12]) ? node23264 : node23257;
															assign node23257 = (inp[11]) ? node23261 : node23258;
																assign node23258 = (inp[0]) ? 4'b0111 : 4'b0110;
																assign node23261 = (inp[0]) ? 4'b0110 : 4'b0111;
															assign node23264 = (inp[0]) ? node23268 : node23265;
																assign node23265 = (inp[11]) ? 4'b0110 : 4'b0111;
																assign node23268 = (inp[11]) ? 4'b0111 : 4'b0110;
														assign node23271 = (inp[12]) ? node23273 : 4'b0110;
															assign node23273 = (inp[0]) ? node23277 : node23274;
																assign node23274 = (inp[11]) ? 4'b0111 : 4'b0110;
																assign node23277 = (inp[11]) ? 4'b0110 : 4'b0111;
													assign node23280 = (inp[11]) ? node23292 : node23281;
														assign node23281 = (inp[2]) ? node23287 : node23282;
															assign node23282 = (inp[12]) ? node23284 : 4'b0100;
																assign node23284 = (inp[0]) ? 4'b0101 : 4'b0100;
															assign node23287 = (inp[12]) ? 4'b0100 : node23288;
																assign node23288 = (inp[0]) ? 4'b0100 : 4'b0101;
														assign node23292 = (inp[0]) ? node23296 : node23293;
															assign node23293 = (inp[12]) ? 4'b0101 : 4'b0100;
															assign node23296 = (inp[12]) ? 4'b0100 : 4'b0101;
										assign node23299 = (inp[2]) ? node23391 : node23300;
											assign node23300 = (inp[11]) ? node23348 : node23301;
												assign node23301 = (inp[0]) ? node23327 : node23302;
													assign node23302 = (inp[7]) ? node23314 : node23303;
														assign node23303 = (inp[4]) ? node23307 : node23304;
															assign node23304 = (inp[15]) ? 4'b0111 : 4'b0100;
															assign node23307 = (inp[15]) ? node23311 : node23308;
																assign node23308 = (inp[12]) ? 4'b0011 : 4'b0111;
																assign node23311 = (inp[12]) ? 4'b0100 : 4'b0000;
														assign node23314 = (inp[4]) ? node23320 : node23315;
															assign node23315 = (inp[15]) ? node23317 : 4'b0101;
																assign node23317 = (inp[12]) ? 4'b0111 : 4'b0011;
															assign node23320 = (inp[15]) ? node23324 : node23321;
																assign node23321 = (inp[12]) ? 4'b0111 : 4'b0110;
																assign node23324 = (inp[12]) ? 4'b0100 : 4'b0101;
													assign node23327 = (inp[15]) ? node23341 : node23328;
														assign node23328 = (inp[4]) ? node23336 : node23329;
															assign node23329 = (inp[12]) ? node23333 : node23330;
																assign node23330 = (inp[7]) ? 4'b0100 : 4'b0101;
																assign node23333 = (inp[7]) ? 4'b0001 : 4'b0101;
															assign node23336 = (inp[7]) ? node23338 : 4'b0110;
																assign node23338 = (inp[12]) ? 4'b0110 : 4'b0111;
														assign node23341 = (inp[4]) ? node23343 : 4'b0110;
															assign node23343 = (inp[7]) ? 4'b0100 : node23344;
																assign node23344 = (inp[12]) ? 4'b0101 : 4'b0001;
												assign node23348 = (inp[0]) ? node23368 : node23349;
													assign node23349 = (inp[4]) ? node23357 : node23350;
														assign node23350 = (inp[15]) ? node23352 : 4'b0101;
															assign node23352 = (inp[12]) ? 4'b0110 : node23353;
																assign node23353 = (inp[7]) ? 4'b0010 : 4'b0110;
														assign node23357 = (inp[15]) ? node23365 : node23358;
															assign node23358 = (inp[12]) ? node23362 : node23359;
																assign node23359 = (inp[7]) ? 4'b0111 : 4'b0110;
																assign node23362 = (inp[7]) ? 4'b0110 : 4'b0010;
															assign node23365 = (inp[12]) ? 4'b0101 : 4'b0100;
													assign node23368 = (inp[15]) ? node23382 : node23369;
														assign node23369 = (inp[4]) ? node23375 : node23370;
															assign node23370 = (inp[7]) ? node23372 : 4'b0100;
																assign node23372 = (inp[12]) ? 4'b0000 : 4'b0101;
															assign node23375 = (inp[7]) ? node23379 : node23376;
																assign node23376 = (inp[12]) ? 4'b0011 : 4'b0111;
																assign node23379 = (inp[12]) ? 4'b0111 : 4'b0110;
														assign node23382 = (inp[4]) ? node23388 : node23383;
															assign node23383 = (inp[7]) ? node23385 : 4'b0111;
																assign node23385 = (inp[12]) ? 4'b0111 : 4'b0011;
															assign node23388 = (inp[12]) ? 4'b0100 : 4'b0101;
											assign node23391 = (inp[0]) ? node23439 : node23392;
												assign node23392 = (inp[11]) ? node23418 : node23393;
													assign node23393 = (inp[15]) ? node23405 : node23394;
														assign node23394 = (inp[4]) ? node23400 : node23395;
															assign node23395 = (inp[7]) ? node23397 : 4'b0101;
																assign node23397 = (inp[12]) ? 4'b0001 : 4'b0100;
															assign node23400 = (inp[12]) ? 4'b0011 : node23401;
																assign node23401 = (inp[7]) ? 4'b0111 : 4'b0110;
														assign node23405 = (inp[4]) ? node23411 : node23406;
															assign node23406 = (inp[12]) ? 4'b0110 : node23407;
																assign node23407 = (inp[7]) ? 4'b0011 : 4'b0110;
															assign node23411 = (inp[7]) ? node23415 : node23412;
																assign node23412 = (inp[12]) ? 4'b0100 : 4'b0000;
																assign node23415 = (inp[12]) ? 4'b0100 : 4'b0101;
													assign node23418 = (inp[15]) ? node23430 : node23419;
														assign node23419 = (inp[4]) ? node23425 : node23420;
															assign node23420 = (inp[12]) ? 4'b0000 : node23421;
																assign node23421 = (inp[7]) ? 4'b0101 : 4'b0100;
															assign node23425 = (inp[12]) ? node23427 : 4'b0111;
																assign node23427 = (inp[7]) ? 4'b0111 : 4'b0010;
														assign node23430 = (inp[4]) ? node23432 : 4'b0111;
															assign node23432 = (inp[7]) ? node23436 : node23433;
																assign node23433 = (inp[12]) ? 4'b0101 : 4'b0001;
																assign node23436 = (inp[12]) ? 4'b0101 : 4'b0100;
												assign node23439 = (inp[4]) ? node23463 : node23440;
													assign node23440 = (inp[15]) ? node23452 : node23441;
														assign node23441 = (inp[12]) ? node23447 : node23442;
															assign node23442 = (inp[7]) ? 4'b0100 : node23443;
																assign node23443 = (inp[11]) ? 4'b0101 : 4'b0100;
															assign node23447 = (inp[11]) ? node23449 : 4'b0000;
																assign node23449 = (inp[7]) ? 4'b0001 : 4'b0101;
														assign node23452 = (inp[7]) ? node23456 : node23453;
															assign node23453 = (inp[11]) ? 4'b0110 : 4'b0111;
															assign node23456 = (inp[12]) ? node23460 : node23457;
																assign node23457 = (inp[11]) ? 4'b0011 : 4'b0010;
																assign node23460 = (inp[11]) ? 4'b0110 : 4'b0111;
													assign node23463 = (inp[15]) ? node23479 : node23464;
														assign node23464 = (inp[7]) ? node23472 : node23465;
															assign node23465 = (inp[12]) ? node23469 : node23466;
																assign node23466 = (inp[11]) ? 4'b0110 : 4'b0111;
																assign node23469 = (inp[11]) ? 4'b0011 : 4'b0010;
															assign node23472 = (inp[12]) ? node23476 : node23473;
																assign node23473 = (inp[11]) ? 4'b0111 : 4'b0110;
																assign node23476 = (inp[11]) ? 4'b0110 : 4'b0111;
														assign node23479 = (inp[12]) ? 4'b0101 : node23480;
															assign node23480 = (inp[7]) ? 4'b0101 : node23481;
																assign node23481 = (inp[11]) ? 4'b0000 : 4'b0001;
							assign node23486 = (inp[5]) ? node23818 : node23487;
								assign node23487 = (inp[11]) ? node23651 : node23488;
									assign node23488 = (inp[0]) ? node23568 : node23489;
										assign node23489 = (inp[7]) ? node23533 : node23490;
											assign node23490 = (inp[4]) ? node23514 : node23491;
												assign node23491 = (inp[15]) ? node23503 : node23492;
													assign node23492 = (inp[12]) ? node23498 : node23493;
														assign node23493 = (inp[13]) ? node23495 : 4'b0100;
															assign node23495 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node23498 = (inp[2]) ? node23500 : 4'b0101;
															assign node23500 = (inp[13]) ? 4'b0100 : 4'b0101;
													assign node23503 = (inp[12]) ? node23509 : node23504;
														assign node23504 = (inp[2]) ? node23506 : 4'b0110;
															assign node23506 = (inp[13]) ? 4'b0110 : 4'b0111;
														assign node23509 = (inp[13]) ? 4'b0111 : node23510;
															assign node23510 = (inp[2]) ? 4'b0110 : 4'b0111;
												assign node23514 = (inp[15]) ? node23526 : node23515;
													assign node23515 = (inp[12]) ? node23521 : node23516;
														assign node23516 = (inp[2]) ? node23518 : 4'b0110;
															assign node23518 = (inp[13]) ? 4'b0110 : 4'b0111;
														assign node23521 = (inp[2]) ? 4'b0011 : node23522;
															assign node23522 = (inp[13]) ? 4'b0010 : 4'b0011;
													assign node23526 = (inp[12]) ? 4'b0101 : node23527;
														assign node23527 = (inp[2]) ? 4'b0000 : node23528;
															assign node23528 = (inp[13]) ? 4'b0000 : 4'b0001;
											assign node23533 = (inp[4]) ? node23557 : node23534;
												assign node23534 = (inp[15]) ? node23546 : node23535;
													assign node23535 = (inp[12]) ? node23541 : node23536;
														assign node23536 = (inp[13]) ? node23538 : 4'b0100;
															assign node23538 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node23541 = (inp[13]) ? node23543 : 4'b0000;
															assign node23543 = (inp[2]) ? 4'b0001 : 4'b0000;
													assign node23546 = (inp[12]) ? node23552 : node23547;
														assign node23547 = (inp[13]) ? node23549 : 4'b0011;
															assign node23549 = (inp[2]) ? 4'b0011 : 4'b0010;
														assign node23552 = (inp[2]) ? node23554 : 4'b0110;
															assign node23554 = (inp[13]) ? 4'b0110 : 4'b0111;
												assign node23557 = (inp[15]) ? node23563 : node23558;
													assign node23558 = (inp[2]) ? node23560 : 4'b0110;
														assign node23560 = (inp[13]) ? 4'b0110 : 4'b0111;
													assign node23563 = (inp[13]) ? 4'b0100 : node23564;
														assign node23564 = (inp[2]) ? 4'b0100 : 4'b0101;
										assign node23568 = (inp[13]) ? node23612 : node23569;
											assign node23569 = (inp[12]) ? node23589 : node23570;
												assign node23570 = (inp[15]) ? node23576 : node23571;
													assign node23571 = (inp[4]) ? node23573 : 4'b0101;
														assign node23573 = (inp[2]) ? 4'b0110 : 4'b0111;
													assign node23576 = (inp[4]) ? node23582 : node23577;
														assign node23577 = (inp[7]) ? 4'b0010 : node23578;
															assign node23578 = (inp[2]) ? 4'b0110 : 4'b0111;
														assign node23582 = (inp[7]) ? node23586 : node23583;
															assign node23583 = (inp[2]) ? 4'b0001 : 4'b0000;
															assign node23586 = (inp[2]) ? 4'b0101 : 4'b0100;
												assign node23589 = (inp[15]) ? node23599 : node23590;
													assign node23590 = (inp[4]) ? node23594 : node23591;
														assign node23591 = (inp[7]) ? 4'b0001 : 4'b0100;
														assign node23594 = (inp[7]) ? node23596 : 4'b0010;
															assign node23596 = (inp[2]) ? 4'b0110 : 4'b0111;
													assign node23599 = (inp[4]) ? node23605 : node23600;
														assign node23600 = (inp[2]) ? 4'b0110 : node23601;
															assign node23601 = (inp[7]) ? 4'b0111 : 4'b0110;
														assign node23605 = (inp[2]) ? node23609 : node23606;
															assign node23606 = (inp[7]) ? 4'b0100 : 4'b0101;
															assign node23609 = (inp[7]) ? 4'b0101 : 4'b0100;
											assign node23612 = (inp[7]) ? node23634 : node23613;
												assign node23613 = (inp[12]) ? node23623 : node23614;
													assign node23614 = (inp[15]) ? node23620 : node23615;
														assign node23615 = (inp[4]) ? 4'b0111 : node23616;
															assign node23616 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node23620 = (inp[4]) ? 4'b0001 : 4'b0111;
													assign node23623 = (inp[15]) ? node23631 : node23624;
														assign node23624 = (inp[4]) ? node23628 : node23625;
															assign node23625 = (inp[2]) ? 4'b0101 : 4'b0100;
															assign node23628 = (inp[2]) ? 4'b0010 : 4'b0011;
														assign node23631 = (inp[4]) ? 4'b0100 : 4'b0110;
												assign node23634 = (inp[4]) ? node23648 : node23635;
													assign node23635 = (inp[15]) ? node23643 : node23636;
														assign node23636 = (inp[12]) ? node23640 : node23637;
															assign node23637 = (inp[2]) ? 4'b0100 : 4'b0101;
															assign node23640 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node23643 = (inp[12]) ? 4'b0111 : node23644;
															assign node23644 = (inp[2]) ? 4'b0010 : 4'b0011;
													assign node23648 = (inp[15]) ? 4'b0101 : 4'b0111;
									assign node23651 = (inp[0]) ? node23735 : node23652;
										assign node23652 = (inp[7]) ? node23700 : node23653;
											assign node23653 = (inp[4]) ? node23677 : node23654;
												assign node23654 = (inp[15]) ? node23666 : node23655;
													assign node23655 = (inp[12]) ? node23661 : node23656;
														assign node23656 = (inp[13]) ? node23658 : 4'b0101;
															assign node23658 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node23661 = (inp[2]) ? node23663 : 4'b0100;
															assign node23663 = (inp[13]) ? 4'b0101 : 4'b0100;
													assign node23666 = (inp[12]) ? node23672 : node23667;
														assign node23667 = (inp[2]) ? node23669 : 4'b0111;
															assign node23669 = (inp[13]) ? 4'b0111 : 4'b0110;
														assign node23672 = (inp[13]) ? 4'b0110 : node23673;
															assign node23673 = (inp[2]) ? 4'b0111 : 4'b0110;
												assign node23677 = (inp[15]) ? node23689 : node23678;
													assign node23678 = (inp[12]) ? node23684 : node23679;
														assign node23679 = (inp[2]) ? node23681 : 4'b0111;
															assign node23681 = (inp[13]) ? 4'b0111 : 4'b0110;
														assign node23684 = (inp[2]) ? 4'b0010 : node23685;
															assign node23685 = (inp[13]) ? 4'b0011 : 4'b0010;
													assign node23689 = (inp[12]) ? node23695 : node23690;
														assign node23690 = (inp[13]) ? 4'b0001 : node23691;
															assign node23691 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node23695 = (inp[2]) ? 4'b0100 : node23696;
															assign node23696 = (inp[13]) ? 4'b0100 : 4'b0101;
											assign node23700 = (inp[4]) ? node23724 : node23701;
												assign node23701 = (inp[15]) ? node23713 : node23702;
													assign node23702 = (inp[12]) ? node23708 : node23703;
														assign node23703 = (inp[2]) ? node23705 : 4'b0101;
															assign node23705 = (inp[13]) ? 4'b0100 : 4'b0101;
														assign node23708 = (inp[13]) ? node23710 : 4'b0001;
															assign node23710 = (inp[2]) ? 4'b0000 : 4'b0001;
													assign node23713 = (inp[12]) ? node23719 : node23714;
														assign node23714 = (inp[2]) ? 4'b0010 : node23715;
															assign node23715 = (inp[13]) ? 4'b0011 : 4'b0010;
														assign node23719 = (inp[13]) ? 4'b0111 : node23720;
															assign node23720 = (inp[2]) ? 4'b0110 : 4'b0111;
												assign node23724 = (inp[15]) ? node23730 : node23725;
													assign node23725 = (inp[2]) ? node23727 : 4'b0111;
														assign node23727 = (inp[13]) ? 4'b0111 : 4'b0110;
													assign node23730 = (inp[2]) ? 4'b0101 : node23731;
														assign node23731 = (inp[13]) ? 4'b0101 : 4'b0100;
										assign node23735 = (inp[2]) ? node23773 : node23736;
											assign node23736 = (inp[15]) ? node23752 : node23737;
												assign node23737 = (inp[4]) ? node23745 : node23738;
													assign node23738 = (inp[7]) ? node23742 : node23739;
														assign node23739 = (inp[12]) ? 4'b0101 : 4'b0100;
														assign node23742 = (inp[12]) ? 4'b0000 : 4'b0100;
													assign node23745 = (inp[12]) ? node23747 : 4'b0110;
														assign node23747 = (inp[7]) ? 4'b0110 : node23748;
															assign node23748 = (inp[13]) ? 4'b0010 : 4'b0011;
												assign node23752 = (inp[4]) ? node23762 : node23753;
													assign node23753 = (inp[12]) ? node23759 : node23754;
														assign node23754 = (inp[7]) ? node23756 : 4'b0110;
															assign node23756 = (inp[13]) ? 4'b0010 : 4'b0011;
														assign node23759 = (inp[7]) ? 4'b0110 : 4'b0111;
													assign node23762 = (inp[7]) ? node23770 : node23763;
														assign node23763 = (inp[12]) ? node23767 : node23764;
															assign node23764 = (inp[13]) ? 4'b0000 : 4'b0001;
															assign node23767 = (inp[13]) ? 4'b0101 : 4'b0100;
														assign node23770 = (inp[13]) ? 4'b0100 : 4'b0101;
											assign node23773 = (inp[15]) ? node23797 : node23774;
												assign node23774 = (inp[4]) ? node23786 : node23775;
													assign node23775 = (inp[12]) ? node23779 : node23776;
														assign node23776 = (inp[13]) ? 4'b0101 : 4'b0100;
														assign node23779 = (inp[7]) ? node23783 : node23780;
															assign node23780 = (inp[13]) ? 4'b0100 : 4'b0101;
															assign node23783 = (inp[13]) ? 4'b0001 : 4'b0000;
													assign node23786 = (inp[13]) ? node23792 : node23787;
														assign node23787 = (inp[12]) ? node23789 : 4'b0111;
															assign node23789 = (inp[7]) ? 4'b0111 : 4'b0011;
														assign node23792 = (inp[7]) ? 4'b0110 : node23793;
															assign node23793 = (inp[12]) ? 4'b0011 : 4'b0110;
												assign node23797 = (inp[4]) ? node23811 : node23798;
													assign node23798 = (inp[12]) ? node23804 : node23799;
														assign node23799 = (inp[7]) ? 4'b0011 : node23800;
															assign node23800 = (inp[13]) ? 4'b0110 : 4'b0111;
														assign node23804 = (inp[7]) ? node23808 : node23805;
															assign node23805 = (inp[13]) ? 4'b0111 : 4'b0110;
															assign node23808 = (inp[13]) ? 4'b0110 : 4'b0111;
													assign node23811 = (inp[12]) ? node23815 : node23812;
														assign node23812 = (inp[7]) ? 4'b0100 : 4'b0000;
														assign node23815 = (inp[7]) ? 4'b0100 : 4'b0101;
								assign node23818 = (inp[2]) ? node24040 : node23819;
									assign node23819 = (inp[0]) ? node23933 : node23820;
										assign node23820 = (inp[13]) ? node23878 : node23821;
											assign node23821 = (inp[11]) ? node23851 : node23822;
												assign node23822 = (inp[15]) ? node23838 : node23823;
													assign node23823 = (inp[4]) ? node23831 : node23824;
														assign node23824 = (inp[12]) ? node23828 : node23825;
															assign node23825 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node23828 = (inp[7]) ? 4'b0101 : 4'b0001;
														assign node23831 = (inp[12]) ? node23835 : node23832;
															assign node23832 = (inp[7]) ? 4'b0010 : 4'b0011;
															assign node23835 = (inp[7]) ? 4'b0010 : 4'b0110;
													assign node23838 = (inp[4]) ? node23846 : node23839;
														assign node23839 = (inp[7]) ? node23843 : node23840;
															assign node23840 = (inp[12]) ? 4'b0010 : 4'b0011;
															assign node23843 = (inp[12]) ? 4'b0010 : 4'b0110;
														assign node23846 = (inp[7]) ? 4'b0001 : node23847;
															assign node23847 = (inp[12]) ? 4'b0001 : 4'b0101;
												assign node23851 = (inp[7]) ? node23867 : node23852;
													assign node23852 = (inp[4]) ? node23860 : node23853;
														assign node23853 = (inp[15]) ? node23857 : node23854;
															assign node23854 = (inp[12]) ? 4'b0000 : 4'b0001;
															assign node23857 = (inp[12]) ? 4'b0011 : 4'b0010;
														assign node23860 = (inp[15]) ? node23864 : node23861;
															assign node23861 = (inp[12]) ? 4'b0111 : 4'b0010;
															assign node23864 = (inp[12]) ? 4'b0000 : 4'b0100;
													assign node23867 = (inp[4]) ? node23875 : node23868;
														assign node23868 = (inp[15]) ? node23872 : node23869;
															assign node23869 = (inp[12]) ? 4'b0100 : 4'b0000;
															assign node23872 = (inp[12]) ? 4'b0011 : 4'b0111;
														assign node23875 = (inp[15]) ? 4'b0000 : 4'b0011;
											assign node23878 = (inp[11]) ? node23906 : node23879;
												assign node23879 = (inp[4]) ? node23895 : node23880;
													assign node23880 = (inp[15]) ? node23888 : node23881;
														assign node23881 = (inp[7]) ? node23885 : node23882;
															assign node23882 = (inp[12]) ? 4'b0000 : 4'b0001;
															assign node23885 = (inp[12]) ? 4'b0101 : 4'b0000;
														assign node23888 = (inp[7]) ? node23892 : node23889;
															assign node23889 = (inp[12]) ? 4'b0011 : 4'b0010;
															assign node23892 = (inp[12]) ? 4'b0011 : 4'b0111;
													assign node23895 = (inp[15]) ? node23901 : node23896;
														assign node23896 = (inp[7]) ? 4'b0010 : node23897;
															assign node23897 = (inp[12]) ? 4'b0110 : 4'b0011;
														assign node23901 = (inp[7]) ? 4'b0000 : node23902;
															assign node23902 = (inp[12]) ? 4'b0000 : 4'b0101;
												assign node23906 = (inp[4]) ? node23920 : node23907;
													assign node23907 = (inp[15]) ? node23915 : node23908;
														assign node23908 = (inp[12]) ? node23912 : node23909;
															assign node23909 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node23912 = (inp[7]) ? 4'b0100 : 4'b0001;
														assign node23915 = (inp[12]) ? 4'b0010 : node23916;
															assign node23916 = (inp[7]) ? 4'b0110 : 4'b0011;
													assign node23920 = (inp[15]) ? node23928 : node23921;
														assign node23921 = (inp[12]) ? node23925 : node23922;
															assign node23922 = (inp[7]) ? 4'b0011 : 4'b0010;
															assign node23925 = (inp[7]) ? 4'b0011 : 4'b0111;
														assign node23928 = (inp[12]) ? 4'b0001 : node23929;
															assign node23929 = (inp[7]) ? 4'b0001 : 4'b0100;
										assign node23933 = (inp[11]) ? node23983 : node23934;
											assign node23934 = (inp[15]) ? node23956 : node23935;
												assign node23935 = (inp[4]) ? node23949 : node23936;
													assign node23936 = (inp[12]) ? node23944 : node23937;
														assign node23937 = (inp[13]) ? node23941 : node23938;
															assign node23938 = (inp[7]) ? 4'b0000 : 4'b0001;
															assign node23941 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node23944 = (inp[7]) ? 4'b0100 : node23945;
															assign node23945 = (inp[9]) ? 4'b0000 : 4'b0001;
													assign node23949 = (inp[12]) ? node23953 : node23950;
														assign node23950 = (inp[7]) ? 4'b0011 : 4'b0010;
														assign node23953 = (inp[7]) ? 4'b0011 : 4'b0111;
												assign node23956 = (inp[4]) ? node23972 : node23957;
													assign node23957 = (inp[7]) ? node23965 : node23958;
														assign node23958 = (inp[12]) ? node23962 : node23959;
															assign node23959 = (inp[13]) ? 4'b0011 : 4'b0010;
															assign node23962 = (inp[13]) ? 4'b0010 : 4'b0011;
														assign node23965 = (inp[12]) ? node23969 : node23966;
															assign node23966 = (inp[13]) ? 4'b0110 : 4'b0111;
															assign node23969 = (inp[13]) ? 4'b0010 : 4'b0011;
													assign node23972 = (inp[13]) ? node23978 : node23973;
														assign node23973 = (inp[12]) ? 4'b0000 : node23974;
															assign node23974 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node23978 = (inp[12]) ? 4'b0001 : node23979;
															assign node23979 = (inp[7]) ? 4'b0001 : 4'b0100;
											assign node23983 = (inp[13]) ? node24011 : node23984;
												assign node23984 = (inp[15]) ? node23998 : node23985;
													assign node23985 = (inp[4]) ? node23993 : node23986;
														assign node23986 = (inp[12]) ? node23990 : node23987;
															assign node23987 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node23990 = (inp[7]) ? 4'b0101 : 4'b0001;
														assign node23993 = (inp[12]) ? node23995 : 4'b0011;
															assign node23995 = (inp[7]) ? 4'b0010 : 4'b0110;
													assign node23998 = (inp[4]) ? node24006 : node23999;
														assign node23999 = (inp[7]) ? node24003 : node24000;
															assign node24000 = (inp[12]) ? 4'b0010 : 4'b0011;
															assign node24003 = (inp[12]) ? 4'b0010 : 4'b0110;
														assign node24006 = (inp[12]) ? 4'b0001 : node24007;
															assign node24007 = (inp[7]) ? 4'b0001 : 4'b0101;
												assign node24011 = (inp[4]) ? node24027 : node24012;
													assign node24012 = (inp[15]) ? node24020 : node24013;
														assign node24013 = (inp[12]) ? node24017 : node24014;
															assign node24014 = (inp[7]) ? 4'b0000 : 4'b0001;
															assign node24017 = (inp[7]) ? 4'b0101 : 4'b0000;
														assign node24020 = (inp[7]) ? node24024 : node24021;
															assign node24021 = (inp[12]) ? 4'b0011 : 4'b0010;
															assign node24024 = (inp[12]) ? 4'b0011 : 4'b0111;
													assign node24027 = (inp[15]) ? node24035 : node24028;
														assign node24028 = (inp[12]) ? node24032 : node24029;
															assign node24029 = (inp[7]) ? 4'b0010 : 4'b0011;
															assign node24032 = (inp[7]) ? 4'b0010 : 4'b0110;
														assign node24035 = (inp[7]) ? 4'b0000 : node24036;
															assign node24036 = (inp[12]) ? 4'b0000 : 4'b0101;
									assign node24040 = (inp[12]) ? node24168 : node24041;
										assign node24041 = (inp[15]) ? node24099 : node24042;
											assign node24042 = (inp[4]) ? node24066 : node24043;
												assign node24043 = (inp[0]) ? node24051 : node24044;
													assign node24044 = (inp[7]) ? node24048 : node24045;
														assign node24045 = (inp[11]) ? 4'b0000 : 4'b0001;
														assign node24048 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node24051 = (inp[13]) ? node24059 : node24052;
														assign node24052 = (inp[7]) ? node24056 : node24053;
															assign node24053 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node24056 = (inp[11]) ? 4'b0000 : 4'b0001;
														assign node24059 = (inp[7]) ? node24063 : node24060;
															assign node24060 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node24063 = (inp[11]) ? 4'b0000 : 4'b0001;
												assign node24066 = (inp[13]) ? node24086 : node24067;
													assign node24067 = (inp[7]) ? node24079 : node24068;
														assign node24068 = (inp[9]) ? node24074 : node24069;
															assign node24069 = (inp[0]) ? 4'b0011 : node24070;
																assign node24070 = (inp[11]) ? 4'b0011 : 4'b0010;
															assign node24074 = (inp[0]) ? node24076 : 4'b0011;
																assign node24076 = (inp[11]) ? 4'b0010 : 4'b0011;
														assign node24079 = (inp[0]) ? node24083 : node24080;
															assign node24080 = (inp[11]) ? 4'b0010 : 4'b0011;
															assign node24083 = (inp[11]) ? 4'b0011 : 4'b0010;
													assign node24086 = (inp[11]) ? node24094 : node24087;
														assign node24087 = (inp[7]) ? node24091 : node24088;
															assign node24088 = (inp[0]) ? 4'b0010 : 4'b0011;
															assign node24091 = (inp[0]) ? 4'b0011 : 4'b0010;
														assign node24094 = (inp[0]) ? node24096 : 4'b0010;
															assign node24096 = (inp[7]) ? 4'b0010 : 4'b0011;
											assign node24099 = (inp[4]) ? node24131 : node24100;
												assign node24100 = (inp[7]) ? node24114 : node24101;
													assign node24101 = (inp[13]) ? node24109 : node24102;
														assign node24102 = (inp[0]) ? node24106 : node24103;
															assign node24103 = (inp[11]) ? 4'b0010 : 4'b0011;
															assign node24106 = (inp[11]) ? 4'b0011 : 4'b0010;
														assign node24109 = (inp[0]) ? node24111 : 4'b0010;
															assign node24111 = (inp[11]) ? 4'b0011 : 4'b0010;
													assign node24114 = (inp[13]) ? node24122 : node24115;
														assign node24115 = (inp[11]) ? node24119 : node24116;
															assign node24116 = (inp[0]) ? 4'b0111 : 4'b0110;
															assign node24119 = (inp[0]) ? 4'b0110 : 4'b0111;
														assign node24122 = (inp[9]) ? node24128 : node24123;
															assign node24123 = (inp[11]) ? 4'b0110 : node24124;
																assign node24124 = (inp[0]) ? 4'b0111 : 4'b0110;
															assign node24128 = (inp[0]) ? 4'b0110 : 4'b0111;
												assign node24131 = (inp[7]) ? node24161 : node24132;
													assign node24132 = (inp[0]) ? node24148 : node24133;
														assign node24133 = (inp[9]) ? node24141 : node24134;
															assign node24134 = (inp[13]) ? node24138 : node24135;
																assign node24135 = (inp[11]) ? 4'b0100 : 4'b0101;
																assign node24138 = (inp[11]) ? 4'b0101 : 4'b0100;
															assign node24141 = (inp[11]) ? node24145 : node24142;
																assign node24142 = (inp[13]) ? 4'b0100 : 4'b0101;
																assign node24145 = (inp[13]) ? 4'b0101 : 4'b0100;
														assign node24148 = (inp[9]) ? node24156 : node24149;
															assign node24149 = (inp[11]) ? node24153 : node24150;
																assign node24150 = (inp[13]) ? 4'b0101 : 4'b0100;
																assign node24153 = (inp[13]) ? 4'b0100 : 4'b0101;
															assign node24156 = (inp[13]) ? 4'b0101 : node24157;
																assign node24157 = (inp[11]) ? 4'b0101 : 4'b0100;
													assign node24161 = (inp[11]) ? node24165 : node24162;
														assign node24162 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node24165 = (inp[0]) ? 4'b0000 : 4'b0001;
										assign node24168 = (inp[15]) ? node24218 : node24169;
											assign node24169 = (inp[4]) ? node24191 : node24170;
												assign node24170 = (inp[7]) ? node24178 : node24171;
													assign node24171 = (inp[0]) ? node24175 : node24172;
														assign node24172 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node24175 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node24178 = (inp[0]) ? 4'b0101 : node24179;
														assign node24179 = (inp[9]) ? node24185 : node24180;
															assign node24180 = (inp[13]) ? 4'b0100 : node24181;
																assign node24181 = (inp[11]) ? 4'b0100 : 4'b0101;
															assign node24185 = (inp[11]) ? node24187 : 4'b0100;
																assign node24187 = (inp[13]) ? 4'b0101 : 4'b0100;
												assign node24191 = (inp[7]) ? node24203 : node24192;
													assign node24192 = (inp[13]) ? node24198 : node24193;
														assign node24193 = (inp[0]) ? node24195 : 4'b0111;
															assign node24195 = (inp[11]) ? 4'b0111 : 4'b0110;
														assign node24198 = (inp[0]) ? node24200 : 4'b0110;
															assign node24200 = (inp[11]) ? 4'b0110 : 4'b0111;
													assign node24203 = (inp[11]) ? node24211 : node24204;
														assign node24204 = (inp[13]) ? node24208 : node24205;
															assign node24205 = (inp[0]) ? 4'b0010 : 4'b0011;
															assign node24208 = (inp[0]) ? 4'b0011 : 4'b0010;
														assign node24211 = (inp[13]) ? node24215 : node24212;
															assign node24212 = (inp[0]) ? 4'b0011 : 4'b0010;
															assign node24215 = (inp[0]) ? 4'b0010 : 4'b0011;
											assign node24218 = (inp[4]) ? node24242 : node24219;
												assign node24219 = (inp[9]) ? node24235 : node24220;
													assign node24220 = (inp[13]) ? node24228 : node24221;
														assign node24221 = (inp[0]) ? node24225 : node24222;
															assign node24222 = (inp[11]) ? 4'b0011 : 4'b0010;
															assign node24225 = (inp[11]) ? 4'b0010 : 4'b0011;
														assign node24228 = (inp[11]) ? node24232 : node24229;
															assign node24229 = (inp[0]) ? 4'b0011 : 4'b0010;
															assign node24232 = (inp[0]) ? 4'b0010 : 4'b0011;
													assign node24235 = (inp[11]) ? node24239 : node24236;
														assign node24236 = (inp[0]) ? 4'b0011 : 4'b0010;
														assign node24239 = (inp[0]) ? 4'b0010 : 4'b0011;
												assign node24242 = (inp[13]) ? node24258 : node24243;
													assign node24243 = (inp[7]) ? node24251 : node24244;
														assign node24244 = (inp[11]) ? node24248 : node24245;
															assign node24245 = (inp[0]) ? 4'b0001 : 4'b0000;
															assign node24248 = (inp[0]) ? 4'b0000 : 4'b0001;
														assign node24251 = (inp[0]) ? node24255 : node24252;
															assign node24252 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node24255 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node24258 = (inp[9]) ? node24266 : node24259;
														assign node24259 = (inp[11]) ? node24263 : node24260;
															assign node24260 = (inp[0]) ? 4'b0001 : 4'b0000;
															assign node24263 = (inp[0]) ? 4'b0000 : 4'b0001;
														assign node24266 = (inp[11]) ? node24270 : node24267;
															assign node24267 = (inp[0]) ? 4'b0001 : 4'b0000;
															assign node24270 = (inp[0]) ? 4'b0000 : 4'b0001;
				assign node24273 = (inp[15]) ? node27035 : node24274;
					assign node24274 = (inp[12]) ? node25242 : node24275;
						assign node24275 = (inp[6]) ? node24999 : node24276;
							assign node24276 = (inp[5]) ? node24774 : node24277;
								assign node24277 = (inp[0]) ? node24439 : node24278;
									assign node24278 = (inp[10]) ? node24360 : node24279;
										assign node24279 = (inp[13]) ? node24323 : node24280;
											assign node24280 = (inp[1]) ? node24296 : node24281;
												assign node24281 = (inp[2]) ? node24285 : node24282;
													assign node24282 = (inp[7]) ? 4'b0100 : 4'b0000;
													assign node24285 = (inp[7]) ? node24289 : node24286;
														assign node24286 = (inp[4]) ? 4'b0101 : 4'b0100;
														assign node24289 = (inp[4]) ? node24293 : node24290;
															assign node24290 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node24293 = (inp[11]) ? 4'b0000 : 4'b0001;
												assign node24296 = (inp[11]) ? node24308 : node24297;
													assign node24297 = (inp[2]) ? node24301 : node24298;
														assign node24298 = (inp[7]) ? 4'b0100 : 4'b0000;
														assign node24301 = (inp[7]) ? node24305 : node24302;
															assign node24302 = (inp[4]) ? 4'b0101 : 4'b0100;
															assign node24305 = (inp[4]) ? 4'b0000 : 4'b0001;
													assign node24308 = (inp[4]) ? node24316 : node24309;
														assign node24309 = (inp[7]) ? node24313 : node24310;
															assign node24310 = (inp[2]) ? 4'b0101 : 4'b0001;
															assign node24313 = (inp[2]) ? 4'b0001 : 4'b0101;
														assign node24316 = (inp[2]) ? node24320 : node24317;
															assign node24317 = (inp[7]) ? 4'b0101 : 4'b0001;
															assign node24320 = (inp[7]) ? 4'b0000 : 4'b0100;
											assign node24323 = (inp[11]) ? node24337 : node24324;
												assign node24324 = (inp[2]) ? node24328 : node24325;
													assign node24325 = (inp[7]) ? 4'b0101 : 4'b0001;
													assign node24328 = (inp[7]) ? node24332 : node24329;
														assign node24329 = (inp[4]) ? 4'b0100 : 4'b0101;
														assign node24332 = (inp[4]) ? 4'b0001 : node24333;
															assign node24333 = (inp[1]) ? 4'b0000 : 4'b0001;
												assign node24337 = (inp[1]) ? node24349 : node24338;
													assign node24338 = (inp[2]) ? node24342 : node24339;
														assign node24339 = (inp[7]) ? 4'b0101 : 4'b0001;
														assign node24342 = (inp[7]) ? node24346 : node24343;
															assign node24343 = (inp[4]) ? 4'b0100 : 4'b0101;
															assign node24346 = (inp[4]) ? 4'b0001 : 4'b0000;
													assign node24349 = (inp[2]) ? node24353 : node24350;
														assign node24350 = (inp[7]) ? 4'b0100 : 4'b0000;
														assign node24353 = (inp[4]) ? node24357 : node24354;
															assign node24354 = (inp[7]) ? 4'b0000 : 4'b0100;
															assign node24357 = (inp[7]) ? 4'b0001 : 4'b0101;
										assign node24360 = (inp[13]) ? node24404 : node24361;
											assign node24361 = (inp[1]) ? node24383 : node24362;
												assign node24362 = (inp[2]) ? node24366 : node24363;
													assign node24363 = (inp[7]) ? 4'b0101 : 4'b0001;
													assign node24366 = (inp[7]) ? node24370 : node24367;
														assign node24367 = (inp[4]) ? 4'b0100 : 4'b0101;
														assign node24370 = (inp[9]) ? node24378 : node24371;
															assign node24371 = (inp[11]) ? node24375 : node24372;
																assign node24372 = (inp[4]) ? 4'b0000 : 4'b0001;
																assign node24375 = (inp[4]) ? 4'b0001 : 4'b0000;
															assign node24378 = (inp[11]) ? 4'b0001 : node24379;
																assign node24379 = (inp[4]) ? 4'b0000 : 4'b0001;
												assign node24383 = (inp[11]) ? node24395 : node24384;
													assign node24384 = (inp[2]) ? node24388 : node24385;
														assign node24385 = (inp[7]) ? 4'b0101 : 4'b0001;
														assign node24388 = (inp[7]) ? node24392 : node24389;
															assign node24389 = (inp[4]) ? 4'b0100 : 4'b0101;
															assign node24392 = (inp[4]) ? 4'b0001 : 4'b0000;
													assign node24395 = (inp[2]) ? node24399 : node24396;
														assign node24396 = (inp[7]) ? 4'b0100 : 4'b0000;
														assign node24399 = (inp[4]) ? 4'b0101 : node24400;
															assign node24400 = (inp[7]) ? 4'b0000 : 4'b0100;
											assign node24404 = (inp[2]) ? node24416 : node24405;
												assign node24405 = (inp[7]) ? node24411 : node24406;
													assign node24406 = (inp[11]) ? node24408 : 4'b0000;
														assign node24408 = (inp[1]) ? 4'b0001 : 4'b0000;
													assign node24411 = (inp[11]) ? node24413 : 4'b0100;
														assign node24413 = (inp[1]) ? 4'b0101 : 4'b0100;
												assign node24416 = (inp[7]) ? node24428 : node24417;
													assign node24417 = (inp[4]) ? node24423 : node24418;
														assign node24418 = (inp[9]) ? 4'b0100 : node24419;
															assign node24419 = (inp[1]) ? 4'b0101 : 4'b0100;
														assign node24423 = (inp[11]) ? node24425 : 4'b0101;
															assign node24425 = (inp[1]) ? 4'b0100 : 4'b0101;
													assign node24428 = (inp[4]) ? node24434 : node24429;
														assign node24429 = (inp[11]) ? 4'b0001 : node24430;
															assign node24430 = (inp[1]) ? 4'b0001 : 4'b0000;
														assign node24434 = (inp[1]) ? 4'b0000 : node24435;
															assign node24435 = (inp[11]) ? 4'b0000 : 4'b0001;
									assign node24439 = (inp[9]) ? node24609 : node24440;
										assign node24440 = (inp[4]) ? node24544 : node24441;
											assign node24441 = (inp[13]) ? node24497 : node24442;
												assign node24442 = (inp[10]) ? node24472 : node24443;
													assign node24443 = (inp[11]) ? node24459 : node24444;
														assign node24444 = (inp[1]) ? node24452 : node24445;
															assign node24445 = (inp[7]) ? node24449 : node24446;
																assign node24446 = (inp[2]) ? 4'b0100 : 4'b0000;
																assign node24449 = (inp[2]) ? 4'b0000 : 4'b0100;
															assign node24452 = (inp[2]) ? node24456 : node24453;
																assign node24453 = (inp[7]) ? 4'b0100 : 4'b0000;
																assign node24456 = (inp[7]) ? 4'b0001 : 4'b0100;
														assign node24459 = (inp[1]) ? node24467 : node24460;
															assign node24460 = (inp[2]) ? node24464 : node24461;
																assign node24461 = (inp[7]) ? 4'b0100 : 4'b0000;
																assign node24464 = (inp[7]) ? 4'b0001 : 4'b0100;
															assign node24467 = (inp[2]) ? node24469 : 4'b0101;
																assign node24469 = (inp[7]) ? 4'b0001 : 4'b0101;
													assign node24472 = (inp[11]) ? node24482 : node24473;
														assign node24473 = (inp[7]) ? node24477 : node24474;
															assign node24474 = (inp[2]) ? 4'b0101 : 4'b0001;
															assign node24477 = (inp[2]) ? node24479 : 4'b0101;
																assign node24479 = (inp[1]) ? 4'b0000 : 4'b0001;
														assign node24482 = (inp[1]) ? node24490 : node24483;
															assign node24483 = (inp[7]) ? node24487 : node24484;
																assign node24484 = (inp[2]) ? 4'b0101 : 4'b0001;
																assign node24487 = (inp[2]) ? 4'b0000 : 4'b0101;
															assign node24490 = (inp[7]) ? node24494 : node24491;
																assign node24491 = (inp[2]) ? 4'b0100 : 4'b0000;
																assign node24494 = (inp[2]) ? 4'b0000 : 4'b0100;
												assign node24497 = (inp[1]) ? node24513 : node24498;
													assign node24498 = (inp[10]) ? node24508 : node24499;
														assign node24499 = (inp[2]) ? node24503 : node24500;
															assign node24500 = (inp[7]) ? 4'b0101 : 4'b0001;
															assign node24503 = (inp[7]) ? node24505 : 4'b0101;
																assign node24505 = (inp[11]) ? 4'b0000 : 4'b0001;
														assign node24508 = (inp[2]) ? node24510 : 4'b0100;
															assign node24510 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node24513 = (inp[10]) ? node24529 : node24514;
														assign node24514 = (inp[11]) ? node24522 : node24515;
															assign node24515 = (inp[2]) ? node24519 : node24516;
																assign node24516 = (inp[7]) ? 4'b0101 : 4'b0001;
																assign node24519 = (inp[7]) ? 4'b0000 : 4'b0101;
															assign node24522 = (inp[2]) ? node24526 : node24523;
																assign node24523 = (inp[7]) ? 4'b0100 : 4'b0000;
																assign node24526 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node24529 = (inp[11]) ? node24537 : node24530;
															assign node24530 = (inp[2]) ? node24534 : node24531;
																assign node24531 = (inp[7]) ? 4'b0100 : 4'b0000;
																assign node24534 = (inp[7]) ? 4'b0001 : 4'b0100;
															assign node24537 = (inp[2]) ? node24541 : node24538;
																assign node24538 = (inp[7]) ? 4'b0101 : 4'b0001;
																assign node24541 = (inp[7]) ? 4'b0001 : 4'b0101;
											assign node24544 = (inp[13]) ? node24572 : node24545;
												assign node24545 = (inp[10]) ? node24561 : node24546;
													assign node24546 = (inp[2]) ? node24554 : node24547;
														assign node24547 = (inp[7]) ? 4'b0101 : node24548;
															assign node24548 = (inp[1]) ? node24550 : 4'b0000;
																assign node24550 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node24554 = (inp[7]) ? node24556 : 4'b0101;
															assign node24556 = (inp[11]) ? 4'b0000 : node24557;
																assign node24557 = (inp[1]) ? 4'b0000 : 4'b0001;
													assign node24561 = (inp[7]) ? node24569 : node24562;
														assign node24562 = (inp[2]) ? node24566 : node24563;
															assign node24563 = (inp[11]) ? 4'b0000 : 4'b0001;
															assign node24566 = (inp[11]) ? 4'b0101 : 4'b0100;
														assign node24569 = (inp[2]) ? 4'b0001 : 4'b0101;
												assign node24572 = (inp[10]) ? node24590 : node24573;
													assign node24573 = (inp[2]) ? node24581 : node24574;
														assign node24574 = (inp[7]) ? 4'b0101 : node24575;
															assign node24575 = (inp[11]) ? node24577 : 4'b0001;
																assign node24577 = (inp[1]) ? 4'b0000 : 4'b0001;
														assign node24581 = (inp[7]) ? node24587 : node24582;
															assign node24582 = (inp[11]) ? node24584 : 4'b0100;
																assign node24584 = (inp[1]) ? 4'b0101 : 4'b0100;
															assign node24587 = (inp[1]) ? 4'b0001 : 4'b0000;
													assign node24590 = (inp[2]) ? node24600 : node24591;
														assign node24591 = (inp[7]) ? node24597 : node24592;
															assign node24592 = (inp[11]) ? node24594 : 4'b0000;
																assign node24594 = (inp[1]) ? 4'b0001 : 4'b0000;
															assign node24597 = (inp[11]) ? 4'b0101 : 4'b0100;
														assign node24600 = (inp[7]) ? node24604 : node24601;
															assign node24601 = (inp[1]) ? 4'b0100 : 4'b0101;
															assign node24604 = (inp[1]) ? 4'b0000 : node24605;
																assign node24605 = (inp[11]) ? 4'b0000 : 4'b0001;
										assign node24609 = (inp[2]) ? node24677 : node24610;
											assign node24610 = (inp[7]) ? node24632 : node24611;
												assign node24611 = (inp[13]) ? node24621 : node24612;
													assign node24612 = (inp[10]) ? node24618 : node24613;
														assign node24613 = (inp[1]) ? node24615 : 4'b0000;
															assign node24615 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node24618 = (inp[1]) ? 4'b0000 : 4'b0001;
													assign node24621 = (inp[10]) ? node24627 : node24622;
														assign node24622 = (inp[11]) ? node24624 : 4'b0001;
															assign node24624 = (inp[1]) ? 4'b0000 : 4'b0001;
														assign node24627 = (inp[1]) ? node24629 : 4'b0000;
															assign node24629 = (inp[11]) ? 4'b0001 : 4'b0000;
												assign node24632 = (inp[1]) ? node24646 : node24633;
													assign node24633 = (inp[11]) ? node24641 : node24634;
														assign node24634 = (inp[13]) ? node24638 : node24635;
															assign node24635 = (inp[10]) ? 4'b0101 : 4'b0100;
															assign node24638 = (inp[10]) ? 4'b0100 : 4'b0101;
														assign node24641 = (inp[10]) ? 4'b0100 : node24642;
															assign node24642 = (inp[13]) ? 4'b0101 : 4'b0100;
													assign node24646 = (inp[4]) ? node24662 : node24647;
														assign node24647 = (inp[11]) ? node24655 : node24648;
															assign node24648 = (inp[13]) ? node24652 : node24649;
																assign node24649 = (inp[10]) ? 4'b0101 : 4'b0100;
																assign node24652 = (inp[10]) ? 4'b0100 : 4'b0101;
															assign node24655 = (inp[10]) ? node24659 : node24656;
																assign node24656 = (inp[13]) ? 4'b0100 : 4'b0101;
																assign node24659 = (inp[13]) ? 4'b0101 : 4'b0100;
														assign node24662 = (inp[13]) ? node24670 : node24663;
															assign node24663 = (inp[10]) ? node24667 : node24664;
																assign node24664 = (inp[11]) ? 4'b0101 : 4'b0100;
																assign node24667 = (inp[11]) ? 4'b0100 : 4'b0101;
															assign node24670 = (inp[11]) ? node24674 : node24671;
																assign node24671 = (inp[10]) ? 4'b0100 : 4'b0101;
																assign node24674 = (inp[10]) ? 4'b0101 : 4'b0100;
											assign node24677 = (inp[7]) ? node24731 : node24678;
												assign node24678 = (inp[11]) ? node24702 : node24679;
													assign node24679 = (inp[4]) ? node24687 : node24680;
														assign node24680 = (inp[13]) ? node24684 : node24681;
															assign node24681 = (inp[10]) ? 4'b0101 : 4'b0100;
															assign node24684 = (inp[10]) ? 4'b0100 : 4'b0101;
														assign node24687 = (inp[1]) ? node24695 : node24688;
															assign node24688 = (inp[13]) ? node24692 : node24689;
																assign node24689 = (inp[10]) ? 4'b0100 : 4'b0101;
																assign node24692 = (inp[10]) ? 4'b0101 : 4'b0100;
															assign node24695 = (inp[10]) ? node24699 : node24696;
																assign node24696 = (inp[13]) ? 4'b0100 : 4'b0101;
																assign node24699 = (inp[13]) ? 4'b0101 : 4'b0100;
													assign node24702 = (inp[1]) ? node24718 : node24703;
														assign node24703 = (inp[10]) ? node24711 : node24704;
															assign node24704 = (inp[13]) ? node24708 : node24705;
																assign node24705 = (inp[4]) ? 4'b0101 : 4'b0100;
																assign node24708 = (inp[4]) ? 4'b0100 : 4'b0101;
															assign node24711 = (inp[4]) ? node24715 : node24712;
																assign node24712 = (inp[13]) ? 4'b0100 : 4'b0101;
																assign node24715 = (inp[13]) ? 4'b0101 : 4'b0100;
														assign node24718 = (inp[10]) ? node24724 : node24719;
															assign node24719 = (inp[13]) ? node24721 : 4'b0101;
																assign node24721 = (inp[4]) ? 4'b0101 : 4'b0100;
															assign node24724 = (inp[13]) ? node24728 : node24725;
																assign node24725 = (inp[4]) ? 4'b0101 : 4'b0100;
																assign node24728 = (inp[4]) ? 4'b0100 : 4'b0101;
												assign node24731 = (inp[13]) ? node24753 : node24732;
													assign node24732 = (inp[1]) ? node24746 : node24733;
														assign node24733 = (inp[11]) ? node24741 : node24734;
															assign node24734 = (inp[10]) ? node24738 : node24735;
																assign node24735 = (inp[4]) ? 4'b0001 : 4'b0000;
																assign node24738 = (inp[4]) ? 4'b0000 : 4'b0001;
															assign node24741 = (inp[10]) ? node24743 : 4'b0001;
																assign node24743 = (inp[4]) ? 4'b0001 : 4'b0000;
														assign node24746 = (inp[4]) ? node24750 : node24747;
															assign node24747 = (inp[10]) ? 4'b0000 : 4'b0001;
															assign node24750 = (inp[10]) ? 4'b0001 : 4'b0000;
													assign node24753 = (inp[11]) ? node24767 : node24754;
														assign node24754 = (inp[4]) ? node24762 : node24755;
															assign node24755 = (inp[1]) ? node24759 : node24756;
																assign node24756 = (inp[10]) ? 4'b0000 : 4'b0001;
																assign node24759 = (inp[10]) ? 4'b0001 : 4'b0000;
															assign node24762 = (inp[1]) ? 4'b0000 : node24763;
																assign node24763 = (inp[10]) ? 4'b0001 : 4'b0000;
														assign node24767 = (inp[4]) ? node24771 : node24768;
															assign node24768 = (inp[10]) ? 4'b0001 : 4'b0000;
															assign node24771 = (inp[10]) ? 4'b0000 : 4'b0001;
								assign node24774 = (inp[10]) ? node24870 : node24775;
									assign node24775 = (inp[13]) ? node24823 : node24776;
										assign node24776 = (inp[2]) ? node24800 : node24777;
											assign node24777 = (inp[11]) ? node24787 : node24778;
												assign node24778 = (inp[4]) ? node24782 : node24779;
													assign node24779 = (inp[7]) ? 4'b0101 : 4'b0000;
													assign node24782 = (inp[7]) ? 4'b0000 : node24783;
														assign node24783 = (inp[1]) ? 4'b0101 : 4'b0100;
												assign node24787 = (inp[4]) ? node24795 : node24788;
													assign node24788 = (inp[7]) ? node24792 : node24789;
														assign node24789 = (inp[1]) ? 4'b0001 : 4'b0000;
														assign node24792 = (inp[1]) ? 4'b0100 : 4'b0101;
													assign node24795 = (inp[7]) ? node24797 : 4'b0101;
														assign node24797 = (inp[1]) ? 4'b0001 : 4'b0000;
											assign node24800 = (inp[4]) ? node24812 : node24801;
												assign node24801 = (inp[7]) ? node24807 : node24802;
													assign node24802 = (inp[1]) ? node24804 : 4'b0100;
														assign node24804 = (inp[11]) ? 4'b0101 : 4'b0100;
													assign node24807 = (inp[1]) ? 4'b0000 : node24808;
														assign node24808 = (inp[11]) ? 4'b0000 : 4'b0001;
												assign node24812 = (inp[7]) ? node24818 : node24813;
													assign node24813 = (inp[1]) ? node24815 : 4'b0000;
														assign node24815 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node24818 = (inp[11]) ? node24820 : 4'b0101;
														assign node24820 = (inp[1]) ? 4'b0100 : 4'b0101;
										assign node24823 = (inp[2]) ? node24847 : node24824;
											assign node24824 = (inp[1]) ? node24834 : node24825;
												assign node24825 = (inp[4]) ? node24829 : node24826;
													assign node24826 = (inp[7]) ? 4'b0100 : 4'b0001;
													assign node24829 = (inp[7]) ? 4'b0001 : node24830;
														assign node24830 = (inp[11]) ? 4'b0100 : 4'b0101;
												assign node24834 = (inp[7]) ? node24840 : node24835;
													assign node24835 = (inp[4]) ? 4'b0100 : node24836;
														assign node24836 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node24840 = (inp[4]) ? node24844 : node24841;
														assign node24841 = (inp[11]) ? 4'b0101 : 4'b0100;
														assign node24844 = (inp[11]) ? 4'b0000 : 4'b0001;
											assign node24847 = (inp[4]) ? node24859 : node24848;
												assign node24848 = (inp[7]) ? node24854 : node24849;
													assign node24849 = (inp[1]) ? node24851 : 4'b0101;
														assign node24851 = (inp[11]) ? 4'b0100 : 4'b0101;
													assign node24854 = (inp[11]) ? 4'b0001 : node24855;
														assign node24855 = (inp[1]) ? 4'b0001 : 4'b0000;
												assign node24859 = (inp[7]) ? node24865 : node24860;
													assign node24860 = (inp[11]) ? node24862 : 4'b0001;
														assign node24862 = (inp[1]) ? 4'b0000 : 4'b0001;
													assign node24865 = (inp[1]) ? node24867 : 4'b0100;
														assign node24867 = (inp[11]) ? 4'b0101 : 4'b0100;
									assign node24870 = (inp[13]) ? node24952 : node24871;
										assign node24871 = (inp[1]) ? node24891 : node24872;
											assign node24872 = (inp[7]) ? node24882 : node24873;
												assign node24873 = (inp[2]) ? node24879 : node24874;
													assign node24874 = (inp[4]) ? node24876 : 4'b0001;
														assign node24876 = (inp[11]) ? 4'b0100 : 4'b0101;
													assign node24879 = (inp[4]) ? 4'b0001 : 4'b0101;
												assign node24882 = (inp[2]) ? node24886 : node24883;
													assign node24883 = (inp[4]) ? 4'b0001 : 4'b0100;
													assign node24886 = (inp[4]) ? 4'b0100 : node24887;
														assign node24887 = (inp[11]) ? 4'b0001 : 4'b0000;
											assign node24891 = (inp[7]) ? node24929 : node24892;
												assign node24892 = (inp[11]) ? node24906 : node24893;
													assign node24893 = (inp[9]) ? node24901 : node24894;
														assign node24894 = (inp[4]) ? node24898 : node24895;
															assign node24895 = (inp[2]) ? 4'b0101 : 4'b0001;
															assign node24898 = (inp[2]) ? 4'b0001 : 4'b0100;
														assign node24901 = (inp[4]) ? 4'b0001 : node24902;
															assign node24902 = (inp[2]) ? 4'b0101 : 4'b0001;
													assign node24906 = (inp[0]) ? node24914 : node24907;
														assign node24907 = (inp[4]) ? node24911 : node24908;
															assign node24908 = (inp[2]) ? 4'b0100 : 4'b0000;
															assign node24911 = (inp[2]) ? 4'b0000 : 4'b0100;
														assign node24914 = (inp[9]) ? node24922 : node24915;
															assign node24915 = (inp[2]) ? node24919 : node24916;
																assign node24916 = (inp[4]) ? 4'b0100 : 4'b0000;
																assign node24919 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node24922 = (inp[2]) ? node24926 : node24923;
																assign node24923 = (inp[4]) ? 4'b0100 : 4'b0000;
																assign node24926 = (inp[4]) ? 4'b0000 : 4'b0100;
												assign node24929 = (inp[11]) ? node24945 : node24930;
													assign node24930 = (inp[9]) ? node24938 : node24931;
														assign node24931 = (inp[4]) ? node24935 : node24932;
															assign node24932 = (inp[2]) ? 4'b0001 : 4'b0100;
															assign node24935 = (inp[2]) ? 4'b0100 : 4'b0001;
														assign node24938 = (inp[2]) ? node24942 : node24939;
															assign node24939 = (inp[4]) ? 4'b0001 : 4'b0100;
															assign node24942 = (inp[4]) ? 4'b0100 : 4'b0001;
													assign node24945 = (inp[2]) ? node24949 : node24946;
														assign node24946 = (inp[4]) ? 4'b0000 : 4'b0101;
														assign node24949 = (inp[4]) ? 4'b0101 : 4'b0001;
										assign node24952 = (inp[2]) ? node24976 : node24953;
											assign node24953 = (inp[11]) ? node24963 : node24954;
												assign node24954 = (inp[7]) ? node24960 : node24955;
													assign node24955 = (inp[4]) ? node24957 : 4'b0000;
														assign node24957 = (inp[1]) ? 4'b0101 : 4'b0100;
													assign node24960 = (inp[4]) ? 4'b0000 : 4'b0101;
												assign node24963 = (inp[7]) ? node24969 : node24964;
													assign node24964 = (inp[4]) ? 4'b0101 : node24965;
														assign node24965 = (inp[1]) ? 4'b0001 : 4'b0000;
													assign node24969 = (inp[4]) ? node24973 : node24970;
														assign node24970 = (inp[1]) ? 4'b0100 : 4'b0101;
														assign node24973 = (inp[1]) ? 4'b0001 : 4'b0000;
											assign node24976 = (inp[7]) ? node24988 : node24977;
												assign node24977 = (inp[4]) ? node24983 : node24978;
													assign node24978 = (inp[11]) ? node24980 : 4'b0100;
														assign node24980 = (inp[1]) ? 4'b0101 : 4'b0100;
													assign node24983 = (inp[11]) ? node24985 : 4'b0000;
														assign node24985 = (inp[1]) ? 4'b0001 : 4'b0000;
												assign node24988 = (inp[4]) ? node24994 : node24989;
													assign node24989 = (inp[1]) ? 4'b0000 : node24990;
														assign node24990 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node24994 = (inp[1]) ? node24996 : 4'b0101;
														assign node24996 = (inp[11]) ? 4'b0100 : 4'b0101;
							assign node24999 = (inp[11]) ? node25155 : node25000;
								assign node25000 = (inp[13]) ? node25112 : node25001;
									assign node25001 = (inp[2]) ? node25017 : node25002;
										assign node25002 = (inp[5]) ? node25006 : node25003;
											assign node25003 = (inp[7]) ? 4'b0110 : 4'b0010;
											assign node25006 = (inp[7]) ? node25012 : node25007;
												assign node25007 = (inp[1]) ? node25009 : 4'b0110;
													assign node25009 = (inp[4]) ? 4'b0111 : 4'b0110;
												assign node25012 = (inp[4]) ? 4'b0010 : node25013;
													assign node25013 = (inp[1]) ? 4'b0010 : 4'b0011;
										assign node25017 = (inp[5]) ? node25101 : node25018;
											assign node25018 = (inp[7]) ? node25072 : node25019;
												assign node25019 = (inp[9]) ? node25041 : node25020;
													assign node25020 = (inp[10]) ? node25034 : node25021;
														assign node25021 = (inp[0]) ? node25029 : node25022;
															assign node25022 = (inp[1]) ? node25026 : node25023;
																assign node25023 = (inp[4]) ? 4'b0011 : 4'b0010;
																assign node25026 = (inp[4]) ? 4'b0010 : 4'b0011;
															assign node25029 = (inp[1]) ? 4'b0010 : node25030;
																assign node25030 = (inp[4]) ? 4'b0011 : 4'b0010;
														assign node25034 = (inp[4]) ? node25038 : node25035;
															assign node25035 = (inp[1]) ? 4'b0011 : 4'b0010;
															assign node25038 = (inp[1]) ? 4'b0010 : 4'b0011;
													assign node25041 = (inp[10]) ? node25057 : node25042;
														assign node25042 = (inp[0]) ? node25050 : node25043;
															assign node25043 = (inp[1]) ? node25047 : node25044;
																assign node25044 = (inp[4]) ? 4'b0011 : 4'b0010;
																assign node25047 = (inp[4]) ? 4'b0010 : 4'b0011;
															assign node25050 = (inp[1]) ? node25054 : node25051;
																assign node25051 = (inp[4]) ? 4'b0011 : 4'b0010;
																assign node25054 = (inp[4]) ? 4'b0010 : 4'b0011;
														assign node25057 = (inp[0]) ? node25065 : node25058;
															assign node25058 = (inp[4]) ? node25062 : node25059;
																assign node25059 = (inp[1]) ? 4'b0011 : 4'b0010;
																assign node25062 = (inp[1]) ? 4'b0010 : 4'b0011;
															assign node25065 = (inp[4]) ? node25069 : node25066;
																assign node25066 = (inp[1]) ? 4'b0011 : 4'b0010;
																assign node25069 = (inp[1]) ? 4'b0010 : 4'b0011;
												assign node25072 = (inp[0]) ? node25094 : node25073;
													assign node25073 = (inp[10]) ? node25081 : node25074;
														assign node25074 = (inp[4]) ? node25078 : node25075;
															assign node25075 = (inp[1]) ? 4'b0111 : 4'b0110;
															assign node25078 = (inp[1]) ? 4'b0110 : 4'b0111;
														assign node25081 = (inp[9]) ? node25089 : node25082;
															assign node25082 = (inp[1]) ? node25086 : node25083;
																assign node25083 = (inp[4]) ? 4'b0111 : 4'b0110;
																assign node25086 = (inp[4]) ? 4'b0110 : 4'b0111;
															assign node25089 = (inp[4]) ? 4'b0110 : node25090;
																assign node25090 = (inp[1]) ? 4'b0111 : 4'b0110;
													assign node25094 = (inp[4]) ? node25098 : node25095;
														assign node25095 = (inp[1]) ? 4'b0111 : 4'b0110;
														assign node25098 = (inp[1]) ? 4'b0110 : 4'b0111;
											assign node25101 = (inp[7]) ? node25107 : node25102;
												assign node25102 = (inp[1]) ? node25104 : 4'b0110;
													assign node25104 = (inp[4]) ? 4'b0110 : 4'b0111;
												assign node25107 = (inp[1]) ? 4'b0010 : node25108;
													assign node25108 = (inp[4]) ? 4'b0011 : 4'b0010;
									assign node25112 = (inp[2]) ? node25128 : node25113;
										assign node25113 = (inp[5]) ? node25117 : node25114;
											assign node25114 = (inp[7]) ? 4'b0111 : 4'b0011;
											assign node25117 = (inp[7]) ? node25123 : node25118;
												assign node25118 = (inp[4]) ? node25120 : 4'b0111;
													assign node25120 = (inp[1]) ? 4'b0110 : 4'b0111;
												assign node25123 = (inp[4]) ? 4'b0011 : node25124;
													assign node25124 = (inp[1]) ? 4'b0011 : 4'b0010;
										assign node25128 = (inp[5]) ? node25144 : node25129;
											assign node25129 = (inp[7]) ? node25137 : node25130;
												assign node25130 = (inp[4]) ? node25134 : node25131;
													assign node25131 = (inp[1]) ? 4'b0010 : 4'b0011;
													assign node25134 = (inp[1]) ? 4'b0011 : 4'b0010;
												assign node25137 = (inp[1]) ? node25141 : node25138;
													assign node25138 = (inp[4]) ? 4'b0110 : 4'b0111;
													assign node25141 = (inp[4]) ? 4'b0111 : 4'b0110;
											assign node25144 = (inp[7]) ? node25150 : node25145;
												assign node25145 = (inp[1]) ? node25147 : 4'b0111;
													assign node25147 = (inp[4]) ? 4'b0111 : 4'b0110;
												assign node25150 = (inp[4]) ? node25152 : 4'b0011;
													assign node25152 = (inp[1]) ? 4'b0011 : 4'b0010;
								assign node25155 = (inp[13]) ? node25199 : node25156;
									assign node25156 = (inp[2]) ? node25172 : node25157;
										assign node25157 = (inp[5]) ? node25161 : node25158;
											assign node25158 = (inp[7]) ? 4'b0111 : 4'b0011;
											assign node25161 = (inp[7]) ? node25167 : node25162;
												assign node25162 = (inp[4]) ? node25164 : 4'b0111;
													assign node25164 = (inp[1]) ? 4'b0110 : 4'b0111;
												assign node25167 = (inp[1]) ? 4'b0011 : node25168;
													assign node25168 = (inp[4]) ? 4'b0011 : 4'b0010;
										assign node25172 = (inp[5]) ? node25188 : node25173;
											assign node25173 = (inp[7]) ? node25181 : node25174;
												assign node25174 = (inp[4]) ? node25178 : node25175;
													assign node25175 = (inp[1]) ? 4'b0010 : 4'b0011;
													assign node25178 = (inp[1]) ? 4'b0011 : 4'b0010;
												assign node25181 = (inp[4]) ? node25185 : node25182;
													assign node25182 = (inp[1]) ? 4'b0110 : 4'b0111;
													assign node25185 = (inp[1]) ? 4'b0111 : 4'b0110;
											assign node25188 = (inp[7]) ? node25194 : node25189;
												assign node25189 = (inp[4]) ? 4'b0111 : node25190;
													assign node25190 = (inp[1]) ? 4'b0110 : 4'b0111;
												assign node25194 = (inp[4]) ? node25196 : 4'b0011;
													assign node25196 = (inp[1]) ? 4'b0011 : 4'b0010;
									assign node25199 = (inp[2]) ? node25215 : node25200;
										assign node25200 = (inp[5]) ? node25204 : node25201;
											assign node25201 = (inp[7]) ? 4'b0110 : 4'b0010;
											assign node25204 = (inp[7]) ? node25210 : node25205;
												assign node25205 = (inp[1]) ? node25207 : 4'b0110;
													assign node25207 = (inp[4]) ? 4'b0111 : 4'b0110;
												assign node25210 = (inp[1]) ? 4'b0010 : node25211;
													assign node25211 = (inp[4]) ? 4'b0010 : 4'b0011;
										assign node25215 = (inp[5]) ? node25231 : node25216;
											assign node25216 = (inp[7]) ? node25224 : node25217;
												assign node25217 = (inp[1]) ? node25221 : node25218;
													assign node25218 = (inp[4]) ? 4'b0011 : 4'b0010;
													assign node25221 = (inp[4]) ? 4'b0010 : 4'b0011;
												assign node25224 = (inp[1]) ? node25228 : node25225;
													assign node25225 = (inp[4]) ? 4'b0111 : 4'b0110;
													assign node25228 = (inp[4]) ? 4'b0110 : 4'b0111;
											assign node25231 = (inp[7]) ? node25237 : node25232;
												assign node25232 = (inp[1]) ? node25234 : 4'b0110;
													assign node25234 = (inp[4]) ? 4'b0110 : 4'b0111;
												assign node25237 = (inp[4]) ? node25239 : 4'b0010;
													assign node25239 = (inp[1]) ? 4'b0010 : 4'b0011;
						assign node25242 = (inp[1]) ? node25894 : node25243;
							assign node25243 = (inp[4]) ? node25553 : node25244;
								assign node25244 = (inp[6]) ? node25340 : node25245;
									assign node25245 = (inp[13]) ? node25293 : node25246;
										assign node25246 = (inp[10]) ? node25278 : node25247;
											assign node25247 = (inp[7]) ? node25251 : node25248;
												assign node25248 = (inp[2]) ? 4'b0110 : 4'b0010;
												assign node25251 = (inp[2]) ? node25275 : node25252;
													assign node25252 = (inp[0]) ? node25260 : node25253;
														assign node25253 = (inp[11]) ? node25257 : node25254;
															assign node25254 = (inp[5]) ? 4'b0111 : 4'b0110;
															assign node25257 = (inp[5]) ? 4'b0110 : 4'b0111;
														assign node25260 = (inp[9]) ? node25268 : node25261;
															assign node25261 = (inp[11]) ? node25265 : node25262;
																assign node25262 = (inp[5]) ? 4'b0111 : 4'b0110;
																assign node25265 = (inp[5]) ? 4'b0110 : 4'b0111;
															assign node25268 = (inp[11]) ? node25272 : node25269;
																assign node25269 = (inp[5]) ? 4'b0111 : 4'b0110;
																assign node25272 = (inp[5]) ? 4'b0110 : 4'b0111;
													assign node25275 = (inp[5]) ? 4'b0010 : 4'b0011;
											assign node25278 = (inp[7]) ? node25282 : node25279;
												assign node25279 = (inp[2]) ? 4'b0111 : 4'b0011;
												assign node25282 = (inp[2]) ? node25290 : node25283;
													assign node25283 = (inp[11]) ? node25287 : node25284;
														assign node25284 = (inp[5]) ? 4'b0110 : 4'b0111;
														assign node25287 = (inp[5]) ? 4'b0111 : 4'b0110;
													assign node25290 = (inp[5]) ? 4'b0011 : 4'b0010;
										assign node25293 = (inp[10]) ? node25309 : node25294;
											assign node25294 = (inp[7]) ? node25298 : node25295;
												assign node25295 = (inp[2]) ? 4'b0111 : 4'b0011;
												assign node25298 = (inp[2]) ? node25306 : node25299;
													assign node25299 = (inp[5]) ? node25303 : node25300;
														assign node25300 = (inp[11]) ? 4'b0110 : 4'b0111;
														assign node25303 = (inp[11]) ? 4'b0111 : 4'b0110;
													assign node25306 = (inp[5]) ? 4'b0011 : 4'b0010;
											assign node25309 = (inp[7]) ? node25313 : node25310;
												assign node25310 = (inp[2]) ? 4'b0110 : 4'b0010;
												assign node25313 = (inp[2]) ? node25337 : node25314;
													assign node25314 = (inp[9]) ? node25322 : node25315;
														assign node25315 = (inp[5]) ? node25319 : node25316;
															assign node25316 = (inp[11]) ? 4'b0111 : 4'b0110;
															assign node25319 = (inp[11]) ? 4'b0110 : 4'b0111;
														assign node25322 = (inp[0]) ? node25330 : node25323;
															assign node25323 = (inp[11]) ? node25327 : node25324;
																assign node25324 = (inp[5]) ? 4'b0111 : 4'b0110;
																assign node25327 = (inp[5]) ? 4'b0110 : 4'b0111;
															assign node25330 = (inp[11]) ? node25334 : node25331;
																assign node25331 = (inp[5]) ? 4'b0111 : 4'b0110;
																assign node25334 = (inp[5]) ? 4'b0110 : 4'b0111;
													assign node25337 = (inp[5]) ? 4'b0010 : 4'b0011;
									assign node25340 = (inp[5]) ? node25428 : node25341;
										assign node25341 = (inp[7]) ? node25373 : node25342;
											assign node25342 = (inp[2]) ? node25366 : node25343;
												assign node25343 = (inp[10]) ? node25351 : node25344;
													assign node25344 = (inp[13]) ? node25348 : node25345;
														assign node25345 = (inp[11]) ? 4'b0011 : 4'b0010;
														assign node25348 = (inp[11]) ? 4'b0010 : 4'b0011;
													assign node25351 = (inp[0]) ? node25359 : node25352;
														assign node25352 = (inp[13]) ? node25356 : node25353;
															assign node25353 = (inp[11]) ? 4'b0011 : 4'b0010;
															assign node25356 = (inp[11]) ? 4'b0010 : 4'b0011;
														assign node25359 = (inp[11]) ? node25363 : node25360;
															assign node25360 = (inp[13]) ? 4'b0011 : 4'b0010;
															assign node25363 = (inp[13]) ? 4'b0010 : 4'b0011;
												assign node25366 = (inp[13]) ? node25370 : node25367;
													assign node25367 = (inp[11]) ? 4'b0011 : 4'b0010;
													assign node25370 = (inp[11]) ? 4'b0010 : 4'b0011;
											assign node25373 = (inp[11]) ? node25421 : node25374;
												assign node25374 = (inp[10]) ? node25398 : node25375;
													assign node25375 = (inp[0]) ? node25383 : node25376;
														assign node25376 = (inp[13]) ? node25380 : node25377;
															assign node25377 = (inp[2]) ? 4'b0111 : 4'b0110;
															assign node25380 = (inp[2]) ? 4'b0110 : 4'b0111;
														assign node25383 = (inp[9]) ? node25391 : node25384;
															assign node25384 = (inp[13]) ? node25388 : node25385;
																assign node25385 = (inp[2]) ? 4'b0111 : 4'b0110;
																assign node25388 = (inp[2]) ? 4'b0110 : 4'b0111;
															assign node25391 = (inp[2]) ? node25395 : node25392;
																assign node25392 = (inp[13]) ? 4'b0111 : 4'b0110;
																assign node25395 = (inp[13]) ? 4'b0110 : 4'b0111;
													assign node25398 = (inp[0]) ? node25406 : node25399;
														assign node25399 = (inp[2]) ? node25403 : node25400;
															assign node25400 = (inp[13]) ? 4'b0111 : 4'b0110;
															assign node25403 = (inp[13]) ? 4'b0110 : 4'b0111;
														assign node25406 = (inp[9]) ? node25414 : node25407;
															assign node25407 = (inp[2]) ? node25411 : node25408;
																assign node25408 = (inp[13]) ? 4'b0111 : 4'b0110;
																assign node25411 = (inp[13]) ? 4'b0110 : 4'b0111;
															assign node25414 = (inp[13]) ? node25418 : node25415;
																assign node25415 = (inp[2]) ? 4'b0111 : 4'b0110;
																assign node25418 = (inp[2]) ? 4'b0110 : 4'b0111;
												assign node25421 = (inp[2]) ? node25425 : node25422;
													assign node25422 = (inp[13]) ? 4'b0110 : 4'b0111;
													assign node25425 = (inp[13]) ? 4'b0111 : 4'b0110;
										assign node25428 = (inp[7]) ? node25522 : node25429;
											assign node25429 = (inp[2]) ? node25477 : node25430;
												assign node25430 = (inp[0]) ? node25462 : node25431;
													assign node25431 = (inp[10]) ? node25447 : node25432;
														assign node25432 = (inp[9]) ? node25440 : node25433;
															assign node25433 = (inp[11]) ? node25437 : node25434;
																assign node25434 = (inp[13]) ? 4'b0111 : 4'b0110;
																assign node25437 = (inp[13]) ? 4'b0110 : 4'b0111;
															assign node25440 = (inp[13]) ? node25444 : node25441;
																assign node25441 = (inp[11]) ? 4'b0111 : 4'b0110;
																assign node25444 = (inp[11]) ? 4'b0110 : 4'b0111;
														assign node25447 = (inp[9]) ? node25455 : node25448;
															assign node25448 = (inp[11]) ? node25452 : node25449;
																assign node25449 = (inp[13]) ? 4'b0111 : 4'b0110;
																assign node25452 = (inp[13]) ? 4'b0110 : 4'b0111;
															assign node25455 = (inp[13]) ? node25459 : node25456;
																assign node25456 = (inp[11]) ? 4'b0111 : 4'b0110;
																assign node25459 = (inp[11]) ? 4'b0110 : 4'b0111;
													assign node25462 = (inp[10]) ? node25470 : node25463;
														assign node25463 = (inp[11]) ? node25467 : node25464;
															assign node25464 = (inp[13]) ? 4'b0111 : 4'b0110;
															assign node25467 = (inp[13]) ? 4'b0110 : 4'b0111;
														assign node25470 = (inp[13]) ? node25474 : node25471;
															assign node25471 = (inp[11]) ? 4'b0111 : 4'b0110;
															assign node25474 = (inp[11]) ? 4'b0110 : 4'b0111;
												assign node25477 = (inp[0]) ? node25499 : node25478;
													assign node25478 = (inp[10]) ? node25492 : node25479;
														assign node25479 = (inp[9]) ? node25487 : node25480;
															assign node25480 = (inp[11]) ? node25484 : node25481;
																assign node25481 = (inp[13]) ? 4'b0111 : 4'b0110;
																assign node25484 = (inp[13]) ? 4'b0110 : 4'b0111;
															assign node25487 = (inp[13]) ? node25489 : 4'b0110;
																assign node25489 = (inp[11]) ? 4'b0110 : 4'b0111;
														assign node25492 = (inp[13]) ? node25496 : node25493;
															assign node25493 = (inp[11]) ? 4'b0111 : 4'b0110;
															assign node25496 = (inp[11]) ? 4'b0110 : 4'b0111;
													assign node25499 = (inp[10]) ? node25515 : node25500;
														assign node25500 = (inp[9]) ? node25508 : node25501;
															assign node25501 = (inp[13]) ? node25505 : node25502;
																assign node25502 = (inp[11]) ? 4'b0111 : 4'b0110;
																assign node25505 = (inp[11]) ? 4'b0110 : 4'b0111;
															assign node25508 = (inp[11]) ? node25512 : node25509;
																assign node25509 = (inp[13]) ? 4'b0111 : 4'b0110;
																assign node25512 = (inp[13]) ? 4'b0110 : 4'b0111;
														assign node25515 = (inp[11]) ? node25519 : node25516;
															assign node25516 = (inp[13]) ? 4'b0111 : 4'b0110;
															assign node25519 = (inp[13]) ? 4'b0110 : 4'b0111;
											assign node25522 = (inp[9]) ? node25530 : node25523;
												assign node25523 = (inp[13]) ? node25527 : node25524;
													assign node25524 = (inp[11]) ? 4'b0011 : 4'b0010;
													assign node25527 = (inp[11]) ? 4'b0010 : 4'b0011;
												assign node25530 = (inp[10]) ? node25546 : node25531;
													assign node25531 = (inp[0]) ? node25539 : node25532;
														assign node25532 = (inp[13]) ? node25536 : node25533;
															assign node25533 = (inp[11]) ? 4'b0011 : 4'b0010;
															assign node25536 = (inp[11]) ? 4'b0010 : 4'b0011;
														assign node25539 = (inp[11]) ? node25543 : node25540;
															assign node25540 = (inp[13]) ? 4'b0011 : 4'b0010;
															assign node25543 = (inp[13]) ? 4'b0010 : 4'b0011;
													assign node25546 = (inp[11]) ? node25550 : node25547;
														assign node25547 = (inp[13]) ? 4'b0011 : 4'b0010;
														assign node25550 = (inp[13]) ? 4'b0010 : 4'b0011;
								assign node25553 = (inp[7]) ? node25735 : node25554;
									assign node25554 = (inp[5]) ? node25632 : node25555;
										assign node25555 = (inp[2]) ? node25609 : node25556;
											assign node25556 = (inp[6]) ? node25594 : node25557;
												assign node25557 = (inp[0]) ? node25579 : node25558;
													assign node25558 = (inp[11]) ? node25566 : node25559;
														assign node25559 = (inp[13]) ? node25563 : node25560;
															assign node25560 = (inp[10]) ? 4'b0111 : 4'b0110;
															assign node25563 = (inp[10]) ? 4'b0110 : 4'b0111;
														assign node25566 = (inp[9]) ? node25572 : node25567;
															assign node25567 = (inp[13]) ? 4'b0110 : node25568;
																assign node25568 = (inp[10]) ? 4'b0111 : 4'b0110;
															assign node25572 = (inp[10]) ? node25576 : node25573;
																assign node25573 = (inp[13]) ? 4'b0111 : 4'b0110;
																assign node25576 = (inp[13]) ? 4'b0110 : 4'b0111;
													assign node25579 = (inp[9]) ? node25587 : node25580;
														assign node25580 = (inp[13]) ? node25584 : node25581;
															assign node25581 = (inp[10]) ? 4'b0111 : 4'b0110;
															assign node25584 = (inp[10]) ? 4'b0110 : 4'b0111;
														assign node25587 = (inp[10]) ? node25591 : node25588;
															assign node25588 = (inp[13]) ? 4'b0111 : 4'b0110;
															assign node25591 = (inp[13]) ? 4'b0110 : 4'b0111;
												assign node25594 = (inp[0]) ? node25602 : node25595;
													assign node25595 = (inp[13]) ? node25599 : node25596;
														assign node25596 = (inp[11]) ? 4'b0011 : 4'b0010;
														assign node25599 = (inp[11]) ? 4'b0010 : 4'b0011;
													assign node25602 = (inp[13]) ? node25606 : node25603;
														assign node25603 = (inp[11]) ? 4'b0011 : 4'b0010;
														assign node25606 = (inp[11]) ? 4'b0010 : 4'b0011;
											assign node25609 = (inp[11]) ? node25621 : node25610;
												assign node25610 = (inp[13]) ? node25616 : node25611;
													assign node25611 = (inp[10]) ? 4'b0010 : node25612;
														assign node25612 = (inp[6]) ? 4'b0010 : 4'b0011;
													assign node25616 = (inp[6]) ? 4'b0011 : node25617;
														assign node25617 = (inp[10]) ? 4'b0011 : 4'b0010;
												assign node25621 = (inp[13]) ? node25627 : node25622;
													assign node25622 = (inp[10]) ? 4'b0011 : node25623;
														assign node25623 = (inp[6]) ? 4'b0011 : 4'b0010;
													assign node25627 = (inp[6]) ? 4'b0010 : node25628;
														assign node25628 = (inp[10]) ? 4'b0010 : 4'b0011;
										assign node25632 = (inp[6]) ? node25688 : node25633;
											assign node25633 = (inp[2]) ? node25649 : node25634;
												assign node25634 = (inp[0]) ? node25642 : node25635;
													assign node25635 = (inp[10]) ? node25639 : node25636;
														assign node25636 = (inp[13]) ? 4'b0010 : 4'b0011;
														assign node25639 = (inp[13]) ? 4'b0011 : 4'b0010;
													assign node25642 = (inp[13]) ? node25646 : node25643;
														assign node25643 = (inp[10]) ? 4'b0010 : 4'b0011;
														assign node25646 = (inp[10]) ? 4'b0011 : 4'b0010;
												assign node25649 = (inp[0]) ? node25667 : node25650;
													assign node25650 = (inp[11]) ? node25660 : node25651;
														assign node25651 = (inp[9]) ? 4'b0110 : node25652;
															assign node25652 = (inp[13]) ? node25656 : node25653;
																assign node25653 = (inp[10]) ? 4'b0111 : 4'b0110;
																assign node25656 = (inp[10]) ? 4'b0110 : 4'b0111;
														assign node25660 = (inp[13]) ? node25664 : node25661;
															assign node25661 = (inp[10]) ? 4'b0111 : 4'b0110;
															assign node25664 = (inp[10]) ? 4'b0110 : 4'b0111;
													assign node25667 = (inp[11]) ? node25673 : node25668;
														assign node25668 = (inp[10]) ? 4'b0111 : node25669;
															assign node25669 = (inp[13]) ? 4'b0111 : 4'b0110;
														assign node25673 = (inp[9]) ? node25681 : node25674;
															assign node25674 = (inp[13]) ? node25678 : node25675;
																assign node25675 = (inp[10]) ? 4'b0111 : 4'b0110;
																assign node25678 = (inp[10]) ? 4'b0110 : 4'b0111;
															assign node25681 = (inp[13]) ? node25685 : node25682;
																assign node25682 = (inp[10]) ? 4'b0111 : 4'b0110;
																assign node25685 = (inp[10]) ? 4'b0110 : 4'b0111;
											assign node25688 = (inp[11]) ? node25696 : node25689;
												assign node25689 = (inp[13]) ? node25693 : node25690;
													assign node25690 = (inp[2]) ? 4'b0110 : 4'b0111;
													assign node25693 = (inp[2]) ? 4'b0111 : 4'b0110;
												assign node25696 = (inp[9]) ? node25720 : node25697;
													assign node25697 = (inp[0]) ? node25713 : node25698;
														assign node25698 = (inp[10]) ? node25706 : node25699;
															assign node25699 = (inp[13]) ? node25703 : node25700;
																assign node25700 = (inp[2]) ? 4'b0111 : 4'b0110;
																assign node25703 = (inp[2]) ? 4'b0110 : 4'b0111;
															assign node25706 = (inp[2]) ? node25710 : node25707;
																assign node25707 = (inp[13]) ? 4'b0111 : 4'b0110;
																assign node25710 = (inp[13]) ? 4'b0110 : 4'b0111;
														assign node25713 = (inp[2]) ? node25717 : node25714;
															assign node25714 = (inp[13]) ? 4'b0111 : 4'b0110;
															assign node25717 = (inp[13]) ? 4'b0110 : 4'b0111;
													assign node25720 = (inp[0]) ? node25728 : node25721;
														assign node25721 = (inp[13]) ? node25725 : node25722;
															assign node25722 = (inp[2]) ? 4'b0111 : 4'b0110;
															assign node25725 = (inp[2]) ? 4'b0110 : 4'b0111;
														assign node25728 = (inp[2]) ? node25732 : node25729;
															assign node25729 = (inp[13]) ? 4'b0111 : 4'b0110;
															assign node25732 = (inp[13]) ? 4'b0110 : 4'b0111;
									assign node25735 = (inp[5]) ? node25793 : node25736;
										assign node25736 = (inp[2]) ? node25770 : node25737;
											assign node25737 = (inp[6]) ? node25763 : node25738;
												assign node25738 = (inp[11]) ? node25756 : node25739;
													assign node25739 = (inp[0]) ? node25749 : node25740;
														assign node25740 = (inp[9]) ? 4'b0011 : node25741;
															assign node25741 = (inp[10]) ? node25745 : node25742;
																assign node25742 = (inp[13]) ? 4'b0010 : 4'b0011;
																assign node25745 = (inp[13]) ? 4'b0011 : 4'b0010;
														assign node25749 = (inp[13]) ? node25753 : node25750;
															assign node25750 = (inp[10]) ? 4'b0010 : 4'b0011;
															assign node25753 = (inp[10]) ? 4'b0011 : 4'b0010;
													assign node25756 = (inp[10]) ? node25760 : node25757;
														assign node25757 = (inp[13]) ? 4'b0010 : 4'b0011;
														assign node25760 = (inp[13]) ? 4'b0011 : 4'b0010;
												assign node25763 = (inp[13]) ? node25767 : node25764;
													assign node25764 = (inp[11]) ? 4'b0110 : 4'b0111;
													assign node25767 = (inp[11]) ? 4'b0111 : 4'b0110;
											assign node25770 = (inp[13]) ? node25782 : node25771;
												assign node25771 = (inp[11]) ? node25777 : node25772;
													assign node25772 = (inp[6]) ? 4'b0110 : node25773;
														assign node25773 = (inp[10]) ? 4'b0111 : 4'b0110;
													assign node25777 = (inp[6]) ? 4'b0111 : node25778;
														assign node25778 = (inp[10]) ? 4'b0111 : 4'b0110;
												assign node25782 = (inp[10]) ? node25788 : node25783;
													assign node25783 = (inp[11]) ? node25785 : 4'b0111;
														assign node25785 = (inp[6]) ? 4'b0110 : 4'b0111;
													assign node25788 = (inp[11]) ? 4'b0110 : node25789;
														assign node25789 = (inp[6]) ? 4'b0111 : 4'b0110;
										assign node25793 = (inp[6]) ? node25843 : node25794;
											assign node25794 = (inp[2]) ? node25836 : node25795;
												assign node25795 = (inp[10]) ? node25819 : node25796;
													assign node25796 = (inp[0]) ? node25804 : node25797;
														assign node25797 = (inp[11]) ? node25801 : node25798;
															assign node25798 = (inp[13]) ? 4'b0111 : 4'b0110;
															assign node25801 = (inp[13]) ? 4'b0110 : 4'b0111;
														assign node25804 = (inp[9]) ? node25812 : node25805;
															assign node25805 = (inp[13]) ? node25809 : node25806;
																assign node25806 = (inp[11]) ? 4'b0111 : 4'b0110;
																assign node25809 = (inp[11]) ? 4'b0110 : 4'b0111;
															assign node25812 = (inp[13]) ? node25816 : node25813;
																assign node25813 = (inp[11]) ? 4'b0111 : 4'b0110;
																assign node25816 = (inp[11]) ? 4'b0110 : 4'b0111;
													assign node25819 = (inp[0]) ? node25829 : node25820;
														assign node25820 = (inp[9]) ? node25822 : 4'b0111;
															assign node25822 = (inp[11]) ? node25826 : node25823;
																assign node25823 = (inp[13]) ? 4'b0110 : 4'b0111;
																assign node25826 = (inp[13]) ? 4'b0111 : 4'b0110;
														assign node25829 = (inp[13]) ? node25833 : node25830;
															assign node25830 = (inp[11]) ? 4'b0110 : 4'b0111;
															assign node25833 = (inp[11]) ? 4'b0111 : 4'b0110;
												assign node25836 = (inp[10]) ? node25840 : node25837;
													assign node25837 = (inp[13]) ? 4'b0011 : 4'b0010;
													assign node25840 = (inp[13]) ? 4'b0010 : 4'b0011;
											assign node25843 = (inp[11]) ? node25851 : node25844;
												assign node25844 = (inp[13]) ? node25848 : node25845;
													assign node25845 = (inp[2]) ? 4'b0010 : 4'b0011;
													assign node25848 = (inp[2]) ? 4'b0011 : 4'b0010;
												assign node25851 = (inp[9]) ? node25881 : node25852;
													assign node25852 = (inp[10]) ? node25866 : node25853;
														assign node25853 = (inp[0]) ? node25859 : node25854;
															assign node25854 = (inp[2]) ? node25856 : 4'b0010;
																assign node25856 = (inp[13]) ? 4'b0010 : 4'b0011;
															assign node25859 = (inp[13]) ? node25863 : node25860;
																assign node25860 = (inp[2]) ? 4'b0011 : 4'b0010;
																assign node25863 = (inp[2]) ? 4'b0010 : 4'b0011;
														assign node25866 = (inp[0]) ? node25874 : node25867;
															assign node25867 = (inp[2]) ? node25871 : node25868;
																assign node25868 = (inp[13]) ? 4'b0011 : 4'b0010;
																assign node25871 = (inp[13]) ? 4'b0010 : 4'b0011;
															assign node25874 = (inp[2]) ? node25878 : node25875;
																assign node25875 = (inp[13]) ? 4'b0011 : 4'b0010;
																assign node25878 = (inp[13]) ? 4'b0010 : 4'b0011;
													assign node25881 = (inp[0]) ? node25889 : node25882;
														assign node25882 = (inp[13]) ? node25886 : node25883;
															assign node25883 = (inp[2]) ? 4'b0011 : 4'b0010;
															assign node25886 = (inp[2]) ? 4'b0010 : 4'b0011;
														assign node25889 = (inp[13]) ? 4'b0011 : node25890;
															assign node25890 = (inp[2]) ? 4'b0011 : 4'b0010;
							assign node25894 = (inp[9]) ? node26492 : node25895;
								assign node25895 = (inp[10]) ? node26141 : node25896;
									assign node25896 = (inp[13]) ? node26020 : node25897;
										assign node25897 = (inp[2]) ? node25955 : node25898;
											assign node25898 = (inp[7]) ? node25926 : node25899;
												assign node25899 = (inp[11]) ? node25913 : node25900;
													assign node25900 = (inp[4]) ? node25906 : node25901;
														assign node25901 = (inp[6]) ? node25903 : 4'b0011;
															assign node25903 = (inp[5]) ? 4'b0111 : 4'b0011;
														assign node25906 = (inp[5]) ? node25910 : node25907;
															assign node25907 = (inp[6]) ? 4'b0010 : 4'b0111;
															assign node25910 = (inp[6]) ? 4'b0110 : 4'b0010;
													assign node25913 = (inp[4]) ? node25919 : node25914;
														assign node25914 = (inp[6]) ? node25916 : 4'b0010;
															assign node25916 = (inp[5]) ? 4'b0110 : 4'b0010;
														assign node25919 = (inp[6]) ? node25923 : node25920;
															assign node25920 = (inp[5]) ? 4'b0011 : 4'b0110;
															assign node25923 = (inp[5]) ? 4'b0111 : 4'b0011;
												assign node25926 = (inp[6]) ? node25936 : node25927;
													assign node25927 = (inp[5]) ? node25933 : node25928;
														assign node25928 = (inp[4]) ? node25930 : 4'b0110;
															assign node25930 = (inp[11]) ? 4'b0011 : 4'b0010;
														assign node25933 = (inp[4]) ? 4'b0110 : 4'b0111;
													assign node25936 = (inp[5]) ? node25940 : node25937;
														assign node25937 = (inp[11]) ? 4'b0111 : 4'b0110;
														assign node25940 = (inp[0]) ? node25948 : node25941;
															assign node25941 = (inp[11]) ? node25945 : node25942;
																assign node25942 = (inp[4]) ? 4'b0010 : 4'b0011;
																assign node25945 = (inp[4]) ? 4'b0011 : 4'b0010;
															assign node25948 = (inp[4]) ? node25952 : node25949;
																assign node25949 = (inp[11]) ? 4'b0010 : 4'b0011;
																assign node25952 = (inp[11]) ? 4'b0011 : 4'b0010;
											assign node25955 = (inp[7]) ? node25993 : node25956;
												assign node25956 = (inp[5]) ? node25978 : node25957;
													assign node25957 = (inp[6]) ? node25963 : node25958;
														assign node25958 = (inp[4]) ? 4'b0011 : node25959;
															assign node25959 = (inp[11]) ? 4'b0110 : 4'b0111;
														assign node25963 = (inp[0]) ? node25971 : node25964;
															assign node25964 = (inp[4]) ? node25968 : node25965;
																assign node25965 = (inp[11]) ? 4'b0011 : 4'b0010;
																assign node25968 = (inp[11]) ? 4'b0010 : 4'b0011;
															assign node25971 = (inp[11]) ? node25975 : node25972;
																assign node25972 = (inp[4]) ? 4'b0011 : 4'b0010;
																assign node25975 = (inp[4]) ? 4'b0010 : 4'b0011;
													assign node25978 = (inp[0]) ? node25986 : node25979;
														assign node25979 = (inp[6]) ? node25983 : node25980;
															assign node25980 = (inp[11]) ? 4'b0110 : 4'b0111;
															assign node25983 = (inp[11]) ? 4'b0111 : 4'b0110;
														assign node25986 = (inp[11]) ? node25990 : node25987;
															assign node25987 = (inp[6]) ? 4'b0110 : 4'b0111;
															assign node25990 = (inp[6]) ? 4'b0111 : 4'b0110;
												assign node25993 = (inp[5]) ? node26005 : node25994;
													assign node25994 = (inp[6]) ? node26002 : node25995;
														assign node25995 = (inp[4]) ? node25999 : node25996;
															assign node25996 = (inp[11]) ? 4'b0011 : 4'b0010;
															assign node25999 = (inp[11]) ? 4'b0110 : 4'b0111;
														assign node26002 = (inp[11]) ? 4'b0111 : 4'b0110;
													assign node26005 = (inp[0]) ? node26013 : node26006;
														assign node26006 = (inp[6]) ? node26010 : node26007;
															assign node26007 = (inp[11]) ? 4'b0010 : 4'b0011;
															assign node26010 = (inp[11]) ? 4'b0011 : 4'b0010;
														assign node26013 = (inp[6]) ? node26017 : node26014;
															assign node26014 = (inp[11]) ? 4'b0010 : 4'b0011;
															assign node26017 = (inp[11]) ? 4'b0011 : 4'b0010;
										assign node26020 = (inp[11]) ? node26076 : node26021;
											assign node26021 = (inp[6]) ? node26045 : node26022;
												assign node26022 = (inp[2]) ? node26034 : node26023;
													assign node26023 = (inp[4]) ? node26029 : node26024;
														assign node26024 = (inp[7]) ? node26026 : 4'b0010;
															assign node26026 = (inp[5]) ? 4'b0110 : 4'b0111;
														assign node26029 = (inp[7]) ? node26031 : 4'b0011;
															assign node26031 = (inp[5]) ? 4'b0111 : 4'b0011;
													assign node26034 = (inp[7]) ? node26040 : node26035;
														assign node26035 = (inp[4]) ? node26037 : 4'b0110;
															assign node26037 = (inp[5]) ? 4'b0110 : 4'b0010;
														assign node26040 = (inp[5]) ? 4'b0010 : node26041;
															assign node26041 = (inp[4]) ? 4'b0110 : 4'b0011;
												assign node26045 = (inp[4]) ? node26061 : node26046;
													assign node26046 = (inp[2]) ? node26054 : node26047;
														assign node26047 = (inp[5]) ? node26051 : node26048;
															assign node26048 = (inp[7]) ? 4'b0111 : 4'b0010;
															assign node26051 = (inp[7]) ? 4'b0010 : 4'b0110;
														assign node26054 = (inp[5]) ? node26058 : node26055;
															assign node26055 = (inp[7]) ? 4'b0111 : 4'b0011;
															assign node26058 = (inp[7]) ? 4'b0011 : 4'b0111;
													assign node26061 = (inp[2]) ? node26069 : node26062;
														assign node26062 = (inp[7]) ? node26066 : node26063;
															assign node26063 = (inp[5]) ? 4'b0111 : 4'b0011;
															assign node26066 = (inp[5]) ? 4'b0011 : 4'b0111;
														assign node26069 = (inp[5]) ? node26073 : node26070;
															assign node26070 = (inp[7]) ? 4'b0111 : 4'b0010;
															assign node26073 = (inp[7]) ? 4'b0011 : 4'b0111;
											assign node26076 = (inp[6]) ? node26104 : node26077;
												assign node26077 = (inp[7]) ? node26089 : node26078;
													assign node26078 = (inp[2]) ? node26084 : node26079;
														assign node26079 = (inp[4]) ? node26081 : 4'b0011;
															assign node26081 = (inp[5]) ? 4'b0010 : 4'b0111;
														assign node26084 = (inp[5]) ? 4'b0111 : node26085;
															assign node26085 = (inp[4]) ? 4'b0010 : 4'b0111;
													assign node26089 = (inp[2]) ? node26097 : node26090;
														assign node26090 = (inp[5]) ? node26094 : node26091;
															assign node26091 = (inp[4]) ? 4'b0010 : 4'b0111;
															assign node26094 = (inp[4]) ? 4'b0111 : 4'b0110;
														assign node26097 = (inp[4]) ? node26101 : node26098;
															assign node26098 = (inp[5]) ? 4'b0011 : 4'b0010;
															assign node26101 = (inp[5]) ? 4'b0011 : 4'b0111;
												assign node26104 = (inp[2]) ? node26126 : node26105;
													assign node26105 = (inp[4]) ? node26113 : node26106;
														assign node26106 = (inp[5]) ? node26110 : node26107;
															assign node26107 = (inp[7]) ? 4'b0110 : 4'b0011;
															assign node26110 = (inp[7]) ? 4'b0011 : 4'b0111;
														assign node26113 = (inp[0]) ? node26121 : node26114;
															assign node26114 = (inp[5]) ? node26118 : node26115;
																assign node26115 = (inp[7]) ? 4'b0110 : 4'b0010;
																assign node26118 = (inp[7]) ? 4'b0010 : 4'b0110;
															assign node26121 = (inp[5]) ? node26123 : 4'b0010;
																assign node26123 = (inp[7]) ? 4'b0010 : 4'b0110;
													assign node26126 = (inp[0]) ? node26134 : node26127;
														assign node26127 = (inp[7]) ? node26131 : node26128;
															assign node26128 = (inp[4]) ? 4'b0011 : 4'b0010;
															assign node26131 = (inp[5]) ? 4'b0010 : 4'b0110;
														assign node26134 = (inp[7]) ? node26138 : node26135;
															assign node26135 = (inp[5]) ? 4'b0110 : 4'b0010;
															assign node26138 = (inp[5]) ? 4'b0010 : 4'b0110;
									assign node26141 = (inp[0]) ? node26325 : node26142;
										assign node26142 = (inp[4]) ? node26234 : node26143;
											assign node26143 = (inp[13]) ? node26183 : node26144;
												assign node26144 = (inp[11]) ? node26170 : node26145;
													assign node26145 = (inp[2]) ? node26159 : node26146;
														assign node26146 = (inp[6]) ? node26152 : node26147;
															assign node26147 = (inp[7]) ? node26149 : 4'b0010;
																assign node26149 = (inp[5]) ? 4'b0110 : 4'b0111;
															assign node26152 = (inp[5]) ? node26156 : node26153;
																assign node26153 = (inp[7]) ? 4'b0110 : 4'b0011;
																assign node26156 = (inp[7]) ? 4'b0011 : 4'b0111;
														assign node26159 = (inp[7]) ? node26163 : node26160;
															assign node26160 = (inp[6]) ? 4'b0010 : 4'b0110;
															assign node26163 = (inp[6]) ? node26167 : node26164;
																assign node26164 = (inp[5]) ? 4'b0010 : 4'b0011;
																assign node26167 = (inp[5]) ? 4'b0010 : 4'b0110;
													assign node26170 = (inp[2]) ? node26178 : node26171;
														assign node26171 = (inp[5]) ? 4'b0110 : node26172;
															assign node26172 = (inp[7]) ? 4'b0111 : node26173;
																assign node26173 = (inp[6]) ? 4'b0010 : 4'b0011;
														assign node26178 = (inp[7]) ? node26180 : 4'b0111;
															assign node26180 = (inp[5]) ? 4'b0011 : 4'b0111;
												assign node26183 = (inp[11]) ? node26209 : node26184;
													assign node26184 = (inp[2]) ? node26198 : node26185;
														assign node26185 = (inp[6]) ? node26191 : node26186;
															assign node26186 = (inp[7]) ? node26188 : 4'b0011;
																assign node26188 = (inp[5]) ? 4'b0111 : 4'b0110;
															assign node26191 = (inp[7]) ? node26195 : node26192;
																assign node26192 = (inp[5]) ? 4'b0110 : 4'b0010;
																assign node26195 = (inp[5]) ? 4'b0010 : 4'b0111;
														assign node26198 = (inp[7]) ? node26204 : node26199;
															assign node26199 = (inp[6]) ? node26201 : 4'b0111;
																assign node26201 = (inp[5]) ? 4'b0111 : 4'b0011;
															assign node26204 = (inp[6]) ? 4'b0111 : node26205;
																assign node26205 = (inp[5]) ? 4'b0011 : 4'b0010;
													assign node26209 = (inp[2]) ? node26221 : node26210;
														assign node26210 = (inp[6]) ? node26214 : node26211;
															assign node26211 = (inp[7]) ? 4'b0110 : 4'b0010;
															assign node26214 = (inp[5]) ? node26218 : node26215;
																assign node26215 = (inp[7]) ? 4'b0110 : 4'b0011;
																assign node26218 = (inp[7]) ? 4'b0011 : 4'b0111;
														assign node26221 = (inp[7]) ? node26227 : node26222;
															assign node26222 = (inp[6]) ? node26224 : 4'b0110;
																assign node26224 = (inp[5]) ? 4'b0110 : 4'b0010;
															assign node26227 = (inp[6]) ? node26231 : node26228;
																assign node26228 = (inp[5]) ? 4'b0010 : 4'b0011;
																assign node26231 = (inp[5]) ? 4'b0010 : 4'b0110;
											assign node26234 = (inp[13]) ? node26280 : node26235;
												assign node26235 = (inp[11]) ? node26259 : node26236;
													assign node26236 = (inp[6]) ? node26250 : node26237;
														assign node26237 = (inp[2]) ? node26243 : node26238;
															assign node26238 = (inp[7]) ? node26240 : 4'b0011;
																assign node26240 = (inp[5]) ? 4'b0111 : 4'b0011;
															assign node26243 = (inp[7]) ? node26247 : node26244;
																assign node26244 = (inp[5]) ? 4'b0110 : 4'b0010;
																assign node26247 = (inp[5]) ? 4'b0010 : 4'b0110;
														assign node26250 = (inp[5]) ? node26256 : node26251;
															assign node26251 = (inp[7]) ? 4'b0110 : node26252;
																assign node26252 = (inp[2]) ? 4'b0011 : 4'b0010;
															assign node26256 = (inp[7]) ? 4'b0010 : 4'b0110;
													assign node26259 = (inp[7]) ? node26269 : node26260;
														assign node26260 = (inp[5]) ? node26264 : node26261;
															assign node26261 = (inp[2]) ? 4'b0010 : 4'b0111;
															assign node26264 = (inp[6]) ? 4'b0111 : node26265;
																assign node26265 = (inp[2]) ? 4'b0111 : 4'b0010;
														assign node26269 = (inp[5]) ? node26275 : node26270;
															assign node26270 = (inp[6]) ? 4'b0111 : node26271;
																assign node26271 = (inp[2]) ? 4'b0111 : 4'b0010;
															assign node26275 = (inp[6]) ? 4'b0011 : node26276;
																assign node26276 = (inp[2]) ? 4'b0011 : 4'b0111;
												assign node26280 = (inp[11]) ? node26304 : node26281;
													assign node26281 = (inp[6]) ? node26297 : node26282;
														assign node26282 = (inp[2]) ? node26290 : node26283;
															assign node26283 = (inp[7]) ? node26287 : node26284;
																assign node26284 = (inp[5]) ? 4'b0010 : 4'b0111;
																assign node26287 = (inp[5]) ? 4'b0110 : 4'b0010;
															assign node26290 = (inp[7]) ? node26294 : node26291;
																assign node26291 = (inp[5]) ? 4'b0111 : 4'b0011;
																assign node26294 = (inp[5]) ? 4'b0011 : 4'b0111;
														assign node26297 = (inp[5]) ? node26301 : node26298;
															assign node26298 = (inp[7]) ? 4'b0111 : 4'b0011;
															assign node26301 = (inp[7]) ? 4'b0011 : 4'b0111;
													assign node26304 = (inp[7]) ? node26314 : node26305;
														assign node26305 = (inp[5]) ? node26311 : node26306;
															assign node26306 = (inp[2]) ? 4'b0011 : node26307;
																assign node26307 = (inp[6]) ? 4'b0010 : 4'b0110;
															assign node26311 = (inp[2]) ? 4'b0110 : 4'b0011;
														assign node26314 = (inp[5]) ? node26320 : node26315;
															assign node26315 = (inp[6]) ? 4'b0110 : node26316;
																assign node26316 = (inp[2]) ? 4'b0110 : 4'b0011;
															assign node26320 = (inp[6]) ? 4'b0010 : node26321;
																assign node26321 = (inp[2]) ? 4'b0010 : 4'b0110;
										assign node26325 = (inp[11]) ? node26407 : node26326;
											assign node26326 = (inp[13]) ? node26366 : node26327;
												assign node26327 = (inp[2]) ? node26351 : node26328;
													assign node26328 = (inp[7]) ? node26338 : node26329;
														assign node26329 = (inp[6]) ? node26335 : node26330;
															assign node26330 = (inp[4]) ? node26332 : 4'b0010;
																assign node26332 = (inp[5]) ? 4'b0011 : 4'b0110;
															assign node26335 = (inp[4]) ? 4'b0010 : 4'b0011;
														assign node26338 = (inp[6]) ? node26346 : node26339;
															assign node26339 = (inp[5]) ? node26343 : node26340;
																assign node26340 = (inp[4]) ? 4'b0011 : 4'b0111;
																assign node26343 = (inp[4]) ? 4'b0111 : 4'b0110;
															assign node26346 = (inp[5]) ? node26348 : 4'b0110;
																assign node26348 = (inp[4]) ? 4'b0010 : 4'b0011;
													assign node26351 = (inp[5]) ? node26363 : node26352;
														assign node26352 = (inp[7]) ? node26358 : node26353;
															assign node26353 = (inp[6]) ? node26355 : 4'b0010;
																assign node26355 = (inp[4]) ? 4'b0011 : 4'b0010;
															assign node26358 = (inp[4]) ? 4'b0110 : node26359;
																assign node26359 = (inp[6]) ? 4'b0110 : 4'b0011;
														assign node26363 = (inp[7]) ? 4'b0010 : 4'b0110;
												assign node26366 = (inp[2]) ? node26392 : node26367;
													assign node26367 = (inp[7]) ? node26381 : node26368;
														assign node26368 = (inp[6]) ? node26374 : node26369;
															assign node26369 = (inp[4]) ? node26371 : 4'b0011;
																assign node26371 = (inp[5]) ? 4'b0010 : 4'b0111;
															assign node26374 = (inp[4]) ? node26378 : node26375;
																assign node26375 = (inp[5]) ? 4'b0110 : 4'b0010;
																assign node26378 = (inp[5]) ? 4'b0111 : 4'b0011;
														assign node26381 = (inp[6]) ? node26387 : node26382;
															assign node26382 = (inp[4]) ? node26384 : 4'b0110;
																assign node26384 = (inp[5]) ? 4'b0110 : 4'b0010;
															assign node26387 = (inp[5]) ? node26389 : 4'b0111;
																assign node26389 = (inp[4]) ? 4'b0011 : 4'b0010;
													assign node26392 = (inp[7]) ? node26402 : node26393;
														assign node26393 = (inp[5]) ? 4'b0111 : node26394;
															assign node26394 = (inp[6]) ? node26398 : node26395;
																assign node26395 = (inp[4]) ? 4'b0011 : 4'b0111;
																assign node26398 = (inp[4]) ? 4'b0010 : 4'b0011;
														assign node26402 = (inp[5]) ? 4'b0011 : node26403;
															assign node26403 = (inp[4]) ? 4'b0111 : 4'b0010;
											assign node26407 = (inp[13]) ? node26453 : node26408;
												assign node26408 = (inp[4]) ? node26430 : node26409;
													assign node26409 = (inp[2]) ? node26423 : node26410;
														assign node26410 = (inp[6]) ? node26416 : node26411;
															assign node26411 = (inp[7]) ? node26413 : 4'b0011;
																assign node26413 = (inp[5]) ? 4'b0110 : 4'b0111;
															assign node26416 = (inp[5]) ? node26420 : node26417;
																assign node26417 = (inp[7]) ? 4'b0111 : 4'b0010;
																assign node26420 = (inp[7]) ? 4'b0010 : 4'b0110;
														assign node26423 = (inp[7]) ? node26425 : 4'b0111;
															assign node26425 = (inp[6]) ? node26427 : 4'b0010;
																assign node26427 = (inp[5]) ? 4'b0011 : 4'b0111;
													assign node26430 = (inp[6]) ? node26444 : node26431;
														assign node26431 = (inp[7]) ? node26437 : node26432;
															assign node26432 = (inp[2]) ? 4'b0010 : node26433;
																assign node26433 = (inp[5]) ? 4'b0010 : 4'b0111;
															assign node26437 = (inp[2]) ? node26441 : node26438;
																assign node26438 = (inp[5]) ? 4'b0111 : 4'b0010;
																assign node26441 = (inp[5]) ? 4'b0011 : 4'b0111;
														assign node26444 = (inp[5]) ? node26450 : node26445;
															assign node26445 = (inp[2]) ? 4'b0010 : node26446;
																assign node26446 = (inp[7]) ? 4'b0111 : 4'b0011;
															assign node26450 = (inp[7]) ? 4'b0011 : 4'b0111;
												assign node26453 = (inp[2]) ? node26477 : node26454;
													assign node26454 = (inp[5]) ? node26464 : node26455;
														assign node26455 = (inp[7]) ? 4'b0110 : node26456;
															assign node26456 = (inp[6]) ? node26460 : node26457;
																assign node26457 = (inp[4]) ? 4'b0110 : 4'b0010;
																assign node26460 = (inp[4]) ? 4'b0010 : 4'b0011;
														assign node26464 = (inp[4]) ? node26472 : node26465;
															assign node26465 = (inp[6]) ? node26469 : node26466;
																assign node26466 = (inp[7]) ? 4'b0111 : 4'b0010;
																assign node26469 = (inp[7]) ? 4'b0011 : 4'b0111;
															assign node26472 = (inp[6]) ? node26474 : 4'b0011;
																assign node26474 = (inp[7]) ? 4'b0010 : 4'b0110;
													assign node26477 = (inp[5]) ? node26489 : node26478;
														assign node26478 = (inp[7]) ? node26484 : node26479;
															assign node26479 = (inp[4]) ? 4'b0011 : node26480;
																assign node26480 = (inp[6]) ? 4'b0010 : 4'b0110;
															assign node26484 = (inp[4]) ? 4'b0110 : node26485;
																assign node26485 = (inp[6]) ? 4'b0110 : 4'b0011;
														assign node26489 = (inp[7]) ? 4'b0010 : 4'b0110;
								assign node26492 = (inp[2]) ? node26796 : node26493;
									assign node26493 = (inp[7]) ? node26655 : node26494;
										assign node26494 = (inp[5]) ? node26570 : node26495;
											assign node26495 = (inp[6]) ? node26525 : node26496;
												assign node26496 = (inp[4]) ? node26512 : node26497;
													assign node26497 = (inp[13]) ? node26505 : node26498;
														assign node26498 = (inp[10]) ? node26502 : node26499;
															assign node26499 = (inp[11]) ? 4'b0010 : 4'b0011;
															assign node26502 = (inp[11]) ? 4'b0011 : 4'b0010;
														assign node26505 = (inp[11]) ? node26509 : node26506;
															assign node26506 = (inp[10]) ? 4'b0011 : 4'b0010;
															assign node26509 = (inp[10]) ? 4'b0010 : 4'b0011;
													assign node26512 = (inp[10]) ? node26520 : node26513;
														assign node26513 = (inp[13]) ? node26517 : node26514;
															assign node26514 = (inp[11]) ? 4'b0110 : 4'b0111;
															assign node26517 = (inp[11]) ? 4'b0111 : 4'b0110;
														assign node26520 = (inp[13]) ? 4'b0110 : node26521;
															assign node26521 = (inp[11]) ? 4'b0111 : 4'b0110;
												assign node26525 = (inp[0]) ? node26541 : node26526;
													assign node26526 = (inp[11]) ? node26534 : node26527;
														assign node26527 = (inp[13]) ? node26531 : node26528;
															assign node26528 = (inp[4]) ? 4'b0010 : 4'b0011;
															assign node26531 = (inp[4]) ? 4'b0011 : 4'b0010;
														assign node26534 = (inp[13]) ? node26538 : node26535;
															assign node26535 = (inp[4]) ? 4'b0011 : 4'b0010;
															assign node26538 = (inp[4]) ? 4'b0010 : 4'b0011;
													assign node26541 = (inp[10]) ? node26557 : node26542;
														assign node26542 = (inp[4]) ? node26550 : node26543;
															assign node26543 = (inp[11]) ? node26547 : node26544;
																assign node26544 = (inp[13]) ? 4'b0010 : 4'b0011;
																assign node26547 = (inp[13]) ? 4'b0011 : 4'b0010;
															assign node26550 = (inp[11]) ? node26554 : node26551;
																assign node26551 = (inp[13]) ? 4'b0011 : 4'b0010;
																assign node26554 = (inp[13]) ? 4'b0010 : 4'b0011;
														assign node26557 = (inp[4]) ? node26565 : node26558;
															assign node26558 = (inp[13]) ? node26562 : node26559;
																assign node26559 = (inp[11]) ? 4'b0010 : 4'b0011;
																assign node26562 = (inp[11]) ? 4'b0011 : 4'b0010;
															assign node26565 = (inp[13]) ? node26567 : 4'b0011;
																assign node26567 = (inp[11]) ? 4'b0010 : 4'b0011;
											assign node26570 = (inp[6]) ? node26628 : node26571;
												assign node26571 = (inp[0]) ? node26601 : node26572;
													assign node26572 = (inp[4]) ? node26586 : node26573;
														assign node26573 = (inp[13]) ? node26579 : node26574;
															assign node26574 = (inp[11]) ? 4'b0010 : node26575;
																assign node26575 = (inp[10]) ? 4'b0010 : 4'b0011;
															assign node26579 = (inp[10]) ? node26583 : node26580;
																assign node26580 = (inp[11]) ? 4'b0011 : 4'b0010;
																assign node26583 = (inp[11]) ? 4'b0010 : 4'b0011;
														assign node26586 = (inp[10]) ? node26594 : node26587;
															assign node26587 = (inp[13]) ? node26591 : node26588;
																assign node26588 = (inp[11]) ? 4'b0011 : 4'b0010;
																assign node26591 = (inp[11]) ? 4'b0010 : 4'b0011;
															assign node26594 = (inp[11]) ? node26598 : node26595;
																assign node26595 = (inp[13]) ? 4'b0010 : 4'b0011;
																assign node26598 = (inp[13]) ? 4'b0011 : 4'b0010;
													assign node26601 = (inp[4]) ? node26615 : node26602;
														assign node26602 = (inp[11]) ? node26608 : node26603;
															assign node26603 = (inp[10]) ? node26605 : 4'b0010;
																assign node26605 = (inp[13]) ? 4'b0011 : 4'b0010;
															assign node26608 = (inp[10]) ? node26612 : node26609;
																assign node26609 = (inp[13]) ? 4'b0011 : 4'b0010;
																assign node26612 = (inp[13]) ? 4'b0010 : 4'b0011;
														assign node26615 = (inp[13]) ? node26623 : node26616;
															assign node26616 = (inp[11]) ? node26620 : node26617;
																assign node26617 = (inp[10]) ? 4'b0011 : 4'b0010;
																assign node26620 = (inp[10]) ? 4'b0010 : 4'b0011;
															assign node26623 = (inp[10]) ? 4'b0010 : node26624;
																assign node26624 = (inp[11]) ? 4'b0010 : 4'b0011;
												assign node26628 = (inp[4]) ? node26636 : node26629;
													assign node26629 = (inp[11]) ? node26633 : node26630;
														assign node26630 = (inp[13]) ? 4'b0110 : 4'b0111;
														assign node26633 = (inp[13]) ? 4'b0111 : 4'b0110;
													assign node26636 = (inp[10]) ? node26650 : node26637;
														assign node26637 = (inp[0]) ? node26645 : node26638;
															assign node26638 = (inp[13]) ? node26642 : node26639;
																assign node26639 = (inp[11]) ? 4'b0111 : 4'b0110;
																assign node26642 = (inp[11]) ? 4'b0110 : 4'b0111;
															assign node26645 = (inp[13]) ? node26647 : 4'b0110;
																assign node26647 = (inp[11]) ? 4'b0110 : 4'b0111;
														assign node26650 = (inp[13]) ? 4'b0110 : node26651;
															assign node26651 = (inp[11]) ? 4'b0111 : 4'b0110;
										assign node26655 = (inp[6]) ? node26749 : node26656;
											assign node26656 = (inp[5]) ? node26700 : node26657;
												assign node26657 = (inp[4]) ? node26675 : node26658;
													assign node26658 = (inp[0]) ? node26666 : node26659;
														assign node26659 = (inp[13]) ? node26663 : node26660;
															assign node26660 = (inp[10]) ? 4'b0111 : 4'b0110;
															assign node26663 = (inp[10]) ? 4'b0110 : 4'b0111;
														assign node26666 = (inp[11]) ? node26668 : 4'b0110;
															assign node26668 = (inp[13]) ? node26672 : node26669;
																assign node26669 = (inp[10]) ? 4'b0111 : 4'b0110;
																assign node26672 = (inp[10]) ? 4'b0110 : 4'b0111;
													assign node26675 = (inp[0]) ? node26685 : node26676;
														assign node26676 = (inp[13]) ? 4'b0010 : node26677;
															assign node26677 = (inp[11]) ? node26681 : node26678;
																assign node26678 = (inp[10]) ? 4'b0011 : 4'b0010;
																assign node26681 = (inp[10]) ? 4'b0010 : 4'b0011;
														assign node26685 = (inp[10]) ? node26693 : node26686;
															assign node26686 = (inp[11]) ? node26690 : node26687;
																assign node26687 = (inp[13]) ? 4'b0011 : 4'b0010;
																assign node26690 = (inp[13]) ? 4'b0010 : 4'b0011;
															assign node26693 = (inp[13]) ? node26697 : node26694;
																assign node26694 = (inp[11]) ? 4'b0010 : 4'b0011;
																assign node26697 = (inp[11]) ? 4'b0011 : 4'b0010;
												assign node26700 = (inp[0]) ? node26724 : node26701;
													assign node26701 = (inp[10]) ? node26709 : node26702;
														assign node26702 = (inp[13]) ? node26706 : node26703;
															assign node26703 = (inp[4]) ? 4'b0110 : 4'b0111;
															assign node26706 = (inp[4]) ? 4'b0111 : 4'b0110;
														assign node26709 = (inp[11]) ? node26717 : node26710;
															assign node26710 = (inp[13]) ? node26714 : node26711;
																assign node26711 = (inp[4]) ? 4'b0111 : 4'b0110;
																assign node26714 = (inp[4]) ? 4'b0110 : 4'b0111;
															assign node26717 = (inp[13]) ? node26721 : node26718;
																assign node26718 = (inp[4]) ? 4'b0111 : 4'b0110;
																assign node26721 = (inp[4]) ? 4'b0110 : 4'b0111;
													assign node26724 = (inp[10]) ? node26740 : node26725;
														assign node26725 = (inp[11]) ? node26733 : node26726;
															assign node26726 = (inp[4]) ? node26730 : node26727;
																assign node26727 = (inp[13]) ? 4'b0110 : 4'b0111;
																assign node26730 = (inp[13]) ? 4'b0111 : 4'b0110;
															assign node26733 = (inp[4]) ? node26737 : node26734;
																assign node26734 = (inp[13]) ? 4'b0110 : 4'b0111;
																assign node26737 = (inp[13]) ? 4'b0111 : 4'b0110;
														assign node26740 = (inp[11]) ? node26742 : 4'b0110;
															assign node26742 = (inp[13]) ? node26746 : node26743;
																assign node26743 = (inp[4]) ? 4'b0111 : 4'b0110;
																assign node26746 = (inp[4]) ? 4'b0110 : 4'b0111;
											assign node26749 = (inp[5]) ? node26765 : node26750;
												assign node26750 = (inp[10]) ? node26758 : node26751;
													assign node26751 = (inp[11]) ? node26755 : node26752;
														assign node26752 = (inp[13]) ? 4'b0111 : 4'b0110;
														assign node26755 = (inp[13]) ? 4'b0110 : 4'b0111;
													assign node26758 = (inp[13]) ? node26762 : node26759;
														assign node26759 = (inp[11]) ? 4'b0111 : 4'b0110;
														assign node26762 = (inp[11]) ? 4'b0110 : 4'b0111;
												assign node26765 = (inp[11]) ? node26781 : node26766;
													assign node26766 = (inp[10]) ? node26774 : node26767;
														assign node26767 = (inp[4]) ? node26771 : node26768;
															assign node26768 = (inp[13]) ? 4'b0010 : 4'b0011;
															assign node26771 = (inp[13]) ? 4'b0011 : 4'b0010;
														assign node26774 = (inp[4]) ? node26778 : node26775;
															assign node26775 = (inp[13]) ? 4'b0010 : 4'b0011;
															assign node26778 = (inp[13]) ? 4'b0011 : 4'b0010;
													assign node26781 = (inp[10]) ? node26789 : node26782;
														assign node26782 = (inp[13]) ? node26786 : node26783;
															assign node26783 = (inp[4]) ? 4'b0011 : 4'b0010;
															assign node26786 = (inp[4]) ? 4'b0010 : 4'b0011;
														assign node26789 = (inp[13]) ? node26793 : node26790;
															assign node26790 = (inp[4]) ? 4'b0011 : 4'b0010;
															assign node26793 = (inp[4]) ? 4'b0010 : 4'b0011;
									assign node26796 = (inp[7]) ? node26922 : node26797;
										assign node26797 = (inp[5]) ? node26861 : node26798;
											assign node26798 = (inp[4]) ? node26838 : node26799;
												assign node26799 = (inp[6]) ? node26823 : node26800;
													assign node26800 = (inp[11]) ? node26812 : node26801;
														assign node26801 = (inp[0]) ? node26807 : node26802;
															assign node26802 = (inp[13]) ? node26804 : 4'b0111;
																assign node26804 = (inp[10]) ? 4'b0111 : 4'b0110;
															assign node26807 = (inp[10]) ? node26809 : 4'b0111;
																assign node26809 = (inp[13]) ? 4'b0111 : 4'b0110;
														assign node26812 = (inp[0]) ? node26818 : node26813;
															assign node26813 = (inp[13]) ? node26815 : 4'b0110;
																assign node26815 = (inp[10]) ? 4'b0110 : 4'b0111;
															assign node26818 = (inp[13]) ? 4'b0110 : node26819;
																assign node26819 = (inp[10]) ? 4'b0111 : 4'b0110;
													assign node26823 = (inp[10]) ? node26831 : node26824;
														assign node26824 = (inp[13]) ? node26828 : node26825;
															assign node26825 = (inp[11]) ? 4'b0011 : 4'b0010;
															assign node26828 = (inp[11]) ? 4'b0010 : 4'b0011;
														assign node26831 = (inp[11]) ? node26835 : node26832;
															assign node26832 = (inp[13]) ? 4'b0011 : 4'b0010;
															assign node26835 = (inp[13]) ? 4'b0010 : 4'b0011;
												assign node26838 = (inp[13]) ? node26850 : node26839;
													assign node26839 = (inp[10]) ? node26845 : node26840;
														assign node26840 = (inp[6]) ? node26842 : 4'b0011;
															assign node26842 = (inp[11]) ? 4'b0010 : 4'b0011;
														assign node26845 = (inp[11]) ? 4'b0010 : node26846;
															assign node26846 = (inp[6]) ? 4'b0011 : 4'b0010;
													assign node26850 = (inp[10]) ? node26856 : node26851;
														assign node26851 = (inp[6]) ? node26853 : 4'b0010;
															assign node26853 = (inp[11]) ? 4'b0011 : 4'b0010;
														assign node26856 = (inp[11]) ? 4'b0011 : node26857;
															assign node26857 = (inp[6]) ? 4'b0010 : 4'b0011;
											assign node26861 = (inp[0]) ? node26899 : node26862;
												assign node26862 = (inp[4]) ? node26876 : node26863;
													assign node26863 = (inp[10]) ? node26869 : node26864;
														assign node26864 = (inp[13]) ? 4'b0111 : node26865;
															assign node26865 = (inp[6]) ? 4'b0110 : 4'b0111;
														assign node26869 = (inp[13]) ? node26873 : node26870;
															assign node26870 = (inp[11]) ? 4'b0111 : 4'b0110;
															assign node26873 = (inp[11]) ? 4'b0110 : 4'b0111;
													assign node26876 = (inp[11]) ? node26888 : node26877;
														assign node26877 = (inp[13]) ? node26883 : node26878;
															assign node26878 = (inp[6]) ? 4'b0110 : node26879;
																assign node26879 = (inp[10]) ? 4'b0110 : 4'b0111;
															assign node26883 = (inp[6]) ? 4'b0111 : node26884;
																assign node26884 = (inp[10]) ? 4'b0111 : 4'b0110;
														assign node26888 = (inp[13]) ? node26894 : node26889;
															assign node26889 = (inp[6]) ? 4'b0111 : node26890;
																assign node26890 = (inp[10]) ? 4'b0111 : 4'b0110;
															assign node26894 = (inp[10]) ? 4'b0110 : node26895;
																assign node26895 = (inp[6]) ? 4'b0110 : 4'b0111;
												assign node26899 = (inp[13]) ? node26911 : node26900;
													assign node26900 = (inp[11]) ? node26906 : node26901;
														assign node26901 = (inp[10]) ? 4'b0110 : node26902;
															assign node26902 = (inp[6]) ? 4'b0110 : 4'b0111;
														assign node26906 = (inp[6]) ? 4'b0111 : node26907;
															assign node26907 = (inp[10]) ? 4'b0111 : 4'b0110;
													assign node26911 = (inp[11]) ? node26917 : node26912;
														assign node26912 = (inp[10]) ? 4'b0111 : node26913;
															assign node26913 = (inp[6]) ? 4'b0111 : 4'b0110;
														assign node26917 = (inp[10]) ? 4'b0110 : node26918;
															assign node26918 = (inp[6]) ? 4'b0110 : 4'b0111;
										assign node26922 = (inp[5]) ? node26980 : node26923;
											assign node26923 = (inp[4]) ? node26957 : node26924;
												assign node26924 = (inp[6]) ? node26940 : node26925;
													assign node26925 = (inp[13]) ? node26933 : node26926;
														assign node26926 = (inp[10]) ? node26930 : node26927;
															assign node26927 = (inp[11]) ? 4'b0011 : 4'b0010;
															assign node26930 = (inp[11]) ? 4'b0010 : 4'b0011;
														assign node26933 = (inp[11]) ? node26937 : node26934;
															assign node26934 = (inp[10]) ? 4'b0010 : 4'b0011;
															assign node26937 = (inp[10]) ? 4'b0011 : 4'b0010;
													assign node26940 = (inp[10]) ? node26950 : node26941;
														assign node26941 = (inp[0]) ? 4'b0110 : node26942;
															assign node26942 = (inp[11]) ? node26946 : node26943;
																assign node26943 = (inp[13]) ? 4'b0111 : 4'b0110;
																assign node26946 = (inp[13]) ? 4'b0110 : 4'b0111;
														assign node26950 = (inp[13]) ? node26954 : node26951;
															assign node26951 = (inp[11]) ? 4'b0111 : 4'b0110;
															assign node26954 = (inp[11]) ? 4'b0110 : 4'b0111;
												assign node26957 = (inp[11]) ? node26969 : node26958;
													assign node26958 = (inp[13]) ? node26964 : node26959;
														assign node26959 = (inp[10]) ? 4'b0110 : node26960;
															assign node26960 = (inp[6]) ? 4'b0110 : 4'b0111;
														assign node26964 = (inp[6]) ? 4'b0111 : node26965;
															assign node26965 = (inp[10]) ? 4'b0111 : 4'b0110;
													assign node26969 = (inp[13]) ? node26975 : node26970;
														assign node26970 = (inp[10]) ? 4'b0111 : node26971;
															assign node26971 = (inp[6]) ? 4'b0111 : 4'b0110;
														assign node26975 = (inp[6]) ? 4'b0110 : node26976;
															assign node26976 = (inp[0]) ? 4'b0111 : 4'b0110;
											assign node26980 = (inp[0]) ? node27004 : node26981;
												assign node26981 = (inp[11]) ? node26993 : node26982;
													assign node26982 = (inp[13]) ? node26988 : node26983;
														assign node26983 = (inp[10]) ? 4'b0010 : node26984;
															assign node26984 = (inp[6]) ? 4'b0010 : 4'b0011;
														assign node26988 = (inp[10]) ? 4'b0011 : node26989;
															assign node26989 = (inp[6]) ? 4'b0011 : 4'b0010;
													assign node26993 = (inp[13]) ? node26999 : node26994;
														assign node26994 = (inp[10]) ? 4'b0011 : node26995;
															assign node26995 = (inp[6]) ? 4'b0011 : 4'b0010;
														assign node26999 = (inp[10]) ? 4'b0010 : node27000;
															assign node27000 = (inp[6]) ? 4'b0010 : 4'b0011;
												assign node27004 = (inp[10]) ? node27028 : node27005;
													assign node27005 = (inp[6]) ? node27013 : node27006;
														assign node27006 = (inp[13]) ? node27010 : node27007;
															assign node27007 = (inp[11]) ? 4'b0010 : 4'b0011;
															assign node27010 = (inp[11]) ? 4'b0011 : 4'b0010;
														assign node27013 = (inp[4]) ? node27021 : node27014;
															assign node27014 = (inp[13]) ? node27018 : node27015;
																assign node27015 = (inp[11]) ? 4'b0011 : 4'b0010;
																assign node27018 = (inp[11]) ? 4'b0010 : 4'b0011;
															assign node27021 = (inp[13]) ? node27025 : node27022;
																assign node27022 = (inp[11]) ? 4'b0011 : 4'b0010;
																assign node27025 = (inp[11]) ? 4'b0010 : 4'b0011;
													assign node27028 = (inp[13]) ? node27032 : node27029;
														assign node27029 = (inp[11]) ? 4'b0011 : 4'b0010;
														assign node27032 = (inp[11]) ? 4'b0010 : 4'b0011;
					assign node27035 = (inp[6]) ? node27643 : node27036;
						assign node27036 = (inp[12]) ? node27256 : node27037;
							assign node27037 = (inp[10]) ? node27125 : node27038;
								assign node27038 = (inp[1]) ? node27082 : node27039;
									assign node27039 = (inp[7]) ? node27055 : node27040;
										assign node27040 = (inp[4]) ? node27044 : node27041;
											assign node27041 = (inp[2]) ? 4'b0110 : 4'b0010;
											assign node27044 = (inp[2]) ? node27050 : node27045;
												assign node27045 = (inp[11]) ? node27047 : 4'b0110;
													assign node27047 = (inp[5]) ? 4'b0111 : 4'b0110;
												assign node27050 = (inp[11]) ? 4'b0010 : node27051;
													assign node27051 = (inp[5]) ? 4'b0010 : 4'b0011;
										assign node27055 = (inp[4]) ? node27071 : node27056;
											assign node27056 = (inp[2]) ? node27064 : node27057;
												assign node27057 = (inp[5]) ? node27061 : node27058;
													assign node27058 = (inp[11]) ? 4'b0011 : 4'b0010;
													assign node27061 = (inp[11]) ? 4'b0010 : 4'b0011;
												assign node27064 = (inp[5]) ? node27068 : node27065;
													assign node27065 = (inp[11]) ? 4'b0111 : 4'b0110;
													assign node27068 = (inp[11]) ? 4'b0110 : 4'b0111;
											assign node27071 = (inp[2]) ? node27077 : node27072;
												assign node27072 = (inp[5]) ? 4'b0110 : node27073;
													assign node27073 = (inp[11]) ? 4'b0111 : 4'b0110;
												assign node27077 = (inp[5]) ? node27079 : 4'b0010;
													assign node27079 = (inp[11]) ? 4'b0010 : 4'b0011;
									assign node27082 = (inp[7]) ? node27098 : node27083;
										assign node27083 = (inp[4]) ? node27087 : node27084;
											assign node27084 = (inp[2]) ? 4'b0111 : 4'b0011;
											assign node27087 = (inp[2]) ? node27093 : node27088;
												assign node27088 = (inp[5]) ? node27090 : 4'b0111;
													assign node27090 = (inp[11]) ? 4'b0110 : 4'b0111;
												assign node27093 = (inp[5]) ? 4'b0011 : node27094;
													assign node27094 = (inp[11]) ? 4'b0011 : 4'b0010;
										assign node27098 = (inp[4]) ? node27114 : node27099;
											assign node27099 = (inp[2]) ? node27107 : node27100;
												assign node27100 = (inp[5]) ? node27104 : node27101;
													assign node27101 = (inp[11]) ? 4'b0010 : 4'b0011;
													assign node27104 = (inp[11]) ? 4'b0011 : 4'b0010;
												assign node27107 = (inp[5]) ? node27111 : node27108;
													assign node27108 = (inp[11]) ? 4'b0110 : 4'b0111;
													assign node27111 = (inp[11]) ? 4'b0111 : 4'b0110;
											assign node27114 = (inp[2]) ? node27120 : node27115;
												assign node27115 = (inp[11]) ? node27117 : 4'b0111;
													assign node27117 = (inp[5]) ? 4'b0111 : 4'b0110;
												assign node27120 = (inp[5]) ? node27122 : 4'b0011;
													assign node27122 = (inp[11]) ? 4'b0011 : 4'b0010;
								assign node27125 = (inp[1]) ? node27191 : node27126;
									assign node27126 = (inp[7]) ? node27142 : node27127;
										assign node27127 = (inp[4]) ? node27131 : node27128;
											assign node27128 = (inp[2]) ? 4'b0111 : 4'b0011;
											assign node27131 = (inp[2]) ? node27137 : node27132;
												assign node27132 = (inp[5]) ? node27134 : 4'b0111;
													assign node27134 = (inp[11]) ? 4'b0110 : 4'b0111;
												assign node27137 = (inp[11]) ? 4'b0011 : node27138;
													assign node27138 = (inp[5]) ? 4'b0011 : 4'b0010;
										assign node27142 = (inp[4]) ? node27180 : node27143;
											assign node27143 = (inp[2]) ? node27173 : node27144;
												assign node27144 = (inp[9]) ? node27152 : node27145;
													assign node27145 = (inp[5]) ? node27149 : node27146;
														assign node27146 = (inp[11]) ? 4'b0010 : 4'b0011;
														assign node27149 = (inp[11]) ? 4'b0011 : 4'b0010;
													assign node27152 = (inp[13]) ? node27160 : node27153;
														assign node27153 = (inp[11]) ? node27157 : node27154;
															assign node27154 = (inp[5]) ? 4'b0010 : 4'b0011;
															assign node27157 = (inp[5]) ? 4'b0011 : 4'b0010;
														assign node27160 = (inp[0]) ? node27168 : node27161;
															assign node27161 = (inp[5]) ? node27165 : node27162;
																assign node27162 = (inp[11]) ? 4'b0010 : 4'b0011;
																assign node27165 = (inp[11]) ? 4'b0011 : 4'b0010;
															assign node27168 = (inp[11]) ? node27170 : 4'b0010;
																assign node27170 = (inp[5]) ? 4'b0011 : 4'b0010;
												assign node27173 = (inp[11]) ? node27177 : node27174;
													assign node27174 = (inp[5]) ? 4'b0110 : 4'b0111;
													assign node27177 = (inp[5]) ? 4'b0111 : 4'b0110;
											assign node27180 = (inp[2]) ? node27186 : node27181;
												assign node27181 = (inp[11]) ? node27183 : 4'b0111;
													assign node27183 = (inp[5]) ? 4'b0111 : 4'b0110;
												assign node27186 = (inp[5]) ? node27188 : 4'b0011;
													assign node27188 = (inp[11]) ? 4'b0011 : 4'b0010;
									assign node27191 = (inp[7]) ? node27207 : node27192;
										assign node27192 = (inp[4]) ? node27196 : node27193;
											assign node27193 = (inp[2]) ? 4'b0110 : 4'b0010;
											assign node27196 = (inp[2]) ? node27202 : node27197;
												assign node27197 = (inp[11]) ? node27199 : 4'b0110;
													assign node27199 = (inp[5]) ? 4'b0111 : 4'b0110;
												assign node27202 = (inp[11]) ? 4'b0010 : node27203;
													assign node27203 = (inp[5]) ? 4'b0010 : 4'b0011;
										assign node27207 = (inp[4]) ? node27245 : node27208;
											assign node27208 = (inp[2]) ? node27216 : node27209;
												assign node27209 = (inp[5]) ? node27213 : node27210;
													assign node27210 = (inp[11]) ? 4'b0011 : 4'b0010;
													assign node27213 = (inp[11]) ? 4'b0010 : 4'b0011;
												assign node27216 = (inp[9]) ? node27230 : node27217;
													assign node27217 = (inp[0]) ? node27223 : node27218;
														assign node27218 = (inp[13]) ? node27220 : 4'b0110;
															assign node27220 = (inp[11]) ? 4'b0110 : 4'b0111;
														assign node27223 = (inp[5]) ? node27227 : node27224;
															assign node27224 = (inp[11]) ? 4'b0111 : 4'b0110;
															assign node27227 = (inp[11]) ? 4'b0110 : 4'b0111;
													assign node27230 = (inp[0]) ? node27238 : node27231;
														assign node27231 = (inp[5]) ? node27235 : node27232;
															assign node27232 = (inp[11]) ? 4'b0111 : 4'b0110;
															assign node27235 = (inp[11]) ? 4'b0110 : 4'b0111;
														assign node27238 = (inp[5]) ? node27242 : node27239;
															assign node27239 = (inp[11]) ? 4'b0111 : 4'b0110;
															assign node27242 = (inp[11]) ? 4'b0110 : 4'b0111;
											assign node27245 = (inp[2]) ? node27251 : node27246;
												assign node27246 = (inp[5]) ? 4'b0110 : node27247;
													assign node27247 = (inp[11]) ? 4'b0111 : 4'b0110;
												assign node27251 = (inp[11]) ? 4'b0010 : node27252;
													assign node27252 = (inp[5]) ? 4'b0011 : 4'b0010;
							assign node27256 = (inp[2]) ? node27404 : node27257;
								assign node27257 = (inp[5]) ? node27281 : node27258;
									assign node27258 = (inp[7]) ? node27270 : node27259;
										assign node27259 = (inp[10]) ? node27265 : node27260;
											assign node27260 = (inp[4]) ? node27262 : 4'b0000;
												assign node27262 = (inp[11]) ? 4'b0001 : 4'b0000;
											assign node27265 = (inp[4]) ? node27267 : 4'b0001;
												assign node27267 = (inp[11]) ? 4'b0000 : 4'b0001;
										assign node27270 = (inp[10]) ? node27276 : node27271;
											assign node27271 = (inp[4]) ? node27273 : 4'b0001;
												assign node27273 = (inp[11]) ? 4'b0000 : 4'b0001;
											assign node27276 = (inp[11]) ? node27278 : 4'b0000;
												assign node27278 = (inp[4]) ? 4'b0001 : 4'b0000;
									assign node27281 = (inp[7]) ? node27337 : node27282;
										assign node27282 = (inp[1]) ? node27322 : node27283;
											assign node27283 = (inp[0]) ? node27315 : node27284;
												assign node27284 = (inp[13]) ? node27292 : node27285;
													assign node27285 = (inp[10]) ? node27289 : node27286;
														assign node27286 = (inp[4]) ? 4'b0101 : 4'b0100;
														assign node27289 = (inp[4]) ? 4'b0100 : 4'b0101;
													assign node27292 = (inp[9]) ? node27300 : node27293;
														assign node27293 = (inp[4]) ? node27297 : node27294;
															assign node27294 = (inp[10]) ? 4'b0101 : 4'b0100;
															assign node27297 = (inp[10]) ? 4'b0100 : 4'b0101;
														assign node27300 = (inp[11]) ? node27308 : node27301;
															assign node27301 = (inp[10]) ? node27305 : node27302;
																assign node27302 = (inp[4]) ? 4'b0101 : 4'b0100;
																assign node27305 = (inp[4]) ? 4'b0100 : 4'b0101;
															assign node27308 = (inp[4]) ? node27312 : node27309;
																assign node27309 = (inp[10]) ? 4'b0101 : 4'b0100;
																assign node27312 = (inp[10]) ? 4'b0100 : 4'b0101;
												assign node27315 = (inp[4]) ? node27319 : node27316;
													assign node27316 = (inp[10]) ? 4'b0101 : 4'b0100;
													assign node27319 = (inp[10]) ? 4'b0100 : 4'b0101;
											assign node27322 = (inp[0]) ? node27330 : node27323;
												assign node27323 = (inp[10]) ? node27327 : node27324;
													assign node27324 = (inp[4]) ? 4'b0101 : 4'b0100;
													assign node27327 = (inp[4]) ? 4'b0100 : 4'b0101;
												assign node27330 = (inp[4]) ? node27334 : node27331;
													assign node27331 = (inp[10]) ? 4'b0101 : 4'b0100;
													assign node27334 = (inp[10]) ? 4'b0100 : 4'b0101;
										assign node27337 = (inp[1]) ? node27381 : node27338;
											assign node27338 = (inp[9]) ? node27366 : node27339;
												assign node27339 = (inp[11]) ? node27359 : node27340;
													assign node27340 = (inp[13]) ? node27354 : node27341;
														assign node27341 = (inp[0]) ? node27349 : node27342;
															assign node27342 = (inp[10]) ? node27346 : node27343;
																assign node27343 = (inp[4]) ? 4'b0101 : 4'b0100;
																assign node27346 = (inp[4]) ? 4'b0100 : 4'b0101;
															assign node27349 = (inp[4]) ? 4'b0101 : node27350;
																assign node27350 = (inp[10]) ? 4'b0101 : 4'b0100;
														assign node27354 = (inp[4]) ? node27356 : 4'b0101;
															assign node27356 = (inp[10]) ? 4'b0100 : 4'b0101;
													assign node27359 = (inp[10]) ? node27363 : node27360;
														assign node27360 = (inp[4]) ? 4'b0101 : 4'b0100;
														assign node27363 = (inp[4]) ? 4'b0100 : 4'b0101;
												assign node27366 = (inp[0]) ? node27374 : node27367;
													assign node27367 = (inp[4]) ? node27371 : node27368;
														assign node27368 = (inp[10]) ? 4'b0101 : 4'b0100;
														assign node27371 = (inp[10]) ? 4'b0100 : 4'b0101;
													assign node27374 = (inp[4]) ? node27378 : node27375;
														assign node27375 = (inp[10]) ? 4'b0101 : 4'b0100;
														assign node27378 = (inp[10]) ? 4'b0100 : 4'b0101;
											assign node27381 = (inp[13]) ? node27397 : node27382;
												assign node27382 = (inp[9]) ? node27390 : node27383;
													assign node27383 = (inp[4]) ? node27387 : node27384;
														assign node27384 = (inp[10]) ? 4'b0101 : 4'b0100;
														assign node27387 = (inp[10]) ? 4'b0100 : 4'b0101;
													assign node27390 = (inp[10]) ? node27394 : node27391;
														assign node27391 = (inp[4]) ? 4'b0101 : 4'b0100;
														assign node27394 = (inp[4]) ? 4'b0100 : 4'b0101;
												assign node27397 = (inp[10]) ? node27401 : node27398;
													assign node27398 = (inp[4]) ? 4'b0101 : 4'b0100;
													assign node27401 = (inp[4]) ? 4'b0100 : 4'b0101;
								assign node27404 = (inp[5]) ? node27490 : node27405;
									assign node27405 = (inp[0]) ? node27467 : node27406;
										assign node27406 = (inp[11]) ? node27430 : node27407;
											assign node27407 = (inp[4]) ? node27415 : node27408;
												assign node27408 = (inp[7]) ? node27412 : node27409;
													assign node27409 = (inp[10]) ? 4'b0101 : 4'b0100;
													assign node27412 = (inp[10]) ? 4'b0100 : 4'b0101;
												assign node27415 = (inp[9]) ? node27423 : node27416;
													assign node27416 = (inp[7]) ? node27420 : node27417;
														assign node27417 = (inp[10]) ? 4'b0100 : 4'b0101;
														assign node27420 = (inp[10]) ? 4'b0101 : 4'b0100;
													assign node27423 = (inp[7]) ? node27427 : node27424;
														assign node27424 = (inp[10]) ? 4'b0100 : 4'b0101;
														assign node27427 = (inp[10]) ? 4'b0101 : 4'b0100;
											assign node27430 = (inp[1]) ? node27438 : node27431;
												assign node27431 = (inp[7]) ? node27435 : node27432;
													assign node27432 = (inp[10]) ? 4'b0101 : 4'b0100;
													assign node27435 = (inp[10]) ? 4'b0100 : 4'b0101;
												assign node27438 = (inp[13]) ? node27460 : node27439;
													assign node27439 = (inp[4]) ? node27453 : node27440;
														assign node27440 = (inp[9]) ? node27446 : node27441;
															assign node27441 = (inp[10]) ? 4'b0100 : node27442;
																assign node27442 = (inp[7]) ? 4'b0101 : 4'b0100;
															assign node27446 = (inp[7]) ? node27450 : node27447;
																assign node27447 = (inp[10]) ? 4'b0101 : 4'b0100;
																assign node27450 = (inp[10]) ? 4'b0100 : 4'b0101;
														assign node27453 = (inp[10]) ? node27457 : node27454;
															assign node27454 = (inp[7]) ? 4'b0101 : 4'b0100;
															assign node27457 = (inp[7]) ? 4'b0100 : 4'b0101;
													assign node27460 = (inp[7]) ? node27464 : node27461;
														assign node27461 = (inp[10]) ? 4'b0101 : 4'b0100;
														assign node27464 = (inp[10]) ? 4'b0100 : 4'b0101;
										assign node27467 = (inp[10]) ? node27479 : node27468;
											assign node27468 = (inp[7]) ? node27474 : node27469;
												assign node27469 = (inp[11]) ? 4'b0100 : node27470;
													assign node27470 = (inp[4]) ? 4'b0101 : 4'b0100;
												assign node27474 = (inp[4]) ? node27476 : 4'b0101;
													assign node27476 = (inp[11]) ? 4'b0101 : 4'b0100;
											assign node27479 = (inp[7]) ? node27485 : node27480;
												assign node27480 = (inp[4]) ? node27482 : 4'b0101;
													assign node27482 = (inp[11]) ? 4'b0101 : 4'b0100;
												assign node27485 = (inp[11]) ? 4'b0100 : node27486;
													assign node27486 = (inp[4]) ? 4'b0101 : 4'b0100;
									assign node27490 = (inp[7]) ? node27564 : node27491;
										assign node27491 = (inp[9]) ? node27541 : node27492;
											assign node27492 = (inp[1]) ? node27518 : node27493;
												assign node27493 = (inp[13]) ? node27501 : node27494;
													assign node27494 = (inp[11]) ? node27498 : node27495;
														assign node27495 = (inp[10]) ? 4'b0001 : 4'b0000;
														assign node27498 = (inp[10]) ? 4'b0000 : 4'b0001;
													assign node27501 = (inp[0]) ? node27511 : node27502;
														assign node27502 = (inp[4]) ? node27508 : node27503;
															assign node27503 = (inp[10]) ? 4'b0000 : node27504;
																assign node27504 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node27508 = (inp[11]) ? 4'b0000 : 4'b0001;
														assign node27511 = (inp[11]) ? node27515 : node27512;
															assign node27512 = (inp[10]) ? 4'b0001 : 4'b0000;
															assign node27515 = (inp[10]) ? 4'b0000 : 4'b0001;
												assign node27518 = (inp[13]) ? node27526 : node27519;
													assign node27519 = (inp[10]) ? node27523 : node27520;
														assign node27520 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node27523 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node27526 = (inp[4]) ? node27534 : node27527;
														assign node27527 = (inp[10]) ? node27531 : node27528;
															assign node27528 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node27531 = (inp[11]) ? 4'b0000 : 4'b0001;
														assign node27534 = (inp[11]) ? node27538 : node27535;
															assign node27535 = (inp[10]) ? 4'b0001 : 4'b0000;
															assign node27538 = (inp[10]) ? 4'b0000 : 4'b0001;
											assign node27541 = (inp[1]) ? node27557 : node27542;
												assign node27542 = (inp[13]) ? node27550 : node27543;
													assign node27543 = (inp[11]) ? node27547 : node27544;
														assign node27544 = (inp[10]) ? 4'b0001 : 4'b0000;
														assign node27547 = (inp[10]) ? 4'b0000 : 4'b0001;
													assign node27550 = (inp[11]) ? node27554 : node27551;
														assign node27551 = (inp[10]) ? 4'b0001 : 4'b0000;
														assign node27554 = (inp[10]) ? 4'b0000 : 4'b0001;
												assign node27557 = (inp[10]) ? node27561 : node27558;
													assign node27558 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node27561 = (inp[11]) ? 4'b0000 : 4'b0001;
										assign node27564 = (inp[4]) ? node27588 : node27565;
											assign node27565 = (inp[9]) ? node27573 : node27566;
												assign node27566 = (inp[10]) ? node27570 : node27567;
													assign node27567 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node27570 = (inp[11]) ? 4'b0000 : 4'b0001;
												assign node27573 = (inp[1]) ? node27581 : node27574;
													assign node27574 = (inp[11]) ? node27578 : node27575;
														assign node27575 = (inp[10]) ? 4'b0001 : 4'b0000;
														assign node27578 = (inp[10]) ? 4'b0000 : 4'b0001;
													assign node27581 = (inp[11]) ? node27585 : node27582;
														assign node27582 = (inp[10]) ? 4'b0001 : 4'b0000;
														assign node27585 = (inp[10]) ? 4'b0000 : 4'b0001;
											assign node27588 = (inp[0]) ? node27628 : node27589;
												assign node27589 = (inp[13]) ? node27605 : node27590;
													assign node27590 = (inp[9]) ? node27598 : node27591;
														assign node27591 = (inp[10]) ? node27595 : node27592;
															assign node27592 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node27595 = (inp[11]) ? 4'b0000 : 4'b0001;
														assign node27598 = (inp[10]) ? node27602 : node27599;
															assign node27599 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node27602 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node27605 = (inp[1]) ? node27613 : node27606;
														assign node27606 = (inp[10]) ? node27610 : node27607;
															assign node27607 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node27610 = (inp[11]) ? 4'b0000 : 4'b0001;
														assign node27613 = (inp[9]) ? node27621 : node27614;
															assign node27614 = (inp[11]) ? node27618 : node27615;
																assign node27615 = (inp[10]) ? 4'b0001 : 4'b0000;
																assign node27618 = (inp[10]) ? 4'b0000 : 4'b0001;
															assign node27621 = (inp[10]) ? node27625 : node27622;
																assign node27622 = (inp[11]) ? 4'b0001 : 4'b0000;
																assign node27625 = (inp[11]) ? 4'b0000 : 4'b0001;
												assign node27628 = (inp[9]) ? node27636 : node27629;
													assign node27629 = (inp[10]) ? node27633 : node27630;
														assign node27630 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node27633 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node27636 = (inp[11]) ? node27640 : node27637;
														assign node27637 = (inp[10]) ? 4'b0001 : 4'b0000;
														assign node27640 = (inp[10]) ? 4'b0000 : 4'b0001;
						assign node27643 = (inp[5]) ? node28055 : node27644;
							assign node27644 = (inp[12]) ? node27904 : node27645;
								assign node27645 = (inp[4]) ? node27881 : node27646;
									assign node27646 = (inp[7]) ? node27748 : node27647;
										assign node27647 = (inp[0]) ? node27711 : node27648;
											assign node27648 = (inp[13]) ? node27696 : node27649;
												assign node27649 = (inp[2]) ? node27673 : node27650;
													assign node27650 = (inp[9]) ? node27666 : node27651;
														assign node27651 = (inp[10]) ? node27659 : node27652;
															assign node27652 = (inp[1]) ? node27656 : node27653;
																assign node27653 = (inp[11]) ? 4'b0001 : 4'b0000;
																assign node27656 = (inp[11]) ? 4'b0000 : 4'b0001;
															assign node27659 = (inp[11]) ? node27663 : node27660;
																assign node27660 = (inp[1]) ? 4'b0001 : 4'b0000;
																assign node27663 = (inp[1]) ? 4'b0000 : 4'b0001;
														assign node27666 = (inp[1]) ? node27670 : node27667;
															assign node27667 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node27670 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node27673 = (inp[9]) ? node27689 : node27674;
														assign node27674 = (inp[10]) ? node27682 : node27675;
															assign node27675 = (inp[11]) ? node27679 : node27676;
																assign node27676 = (inp[1]) ? 4'b0001 : 4'b0000;
																assign node27679 = (inp[1]) ? 4'b0000 : 4'b0001;
															assign node27682 = (inp[1]) ? node27686 : node27683;
																assign node27683 = (inp[11]) ? 4'b0001 : 4'b0000;
																assign node27686 = (inp[11]) ? 4'b0000 : 4'b0001;
														assign node27689 = (inp[1]) ? node27693 : node27690;
															assign node27690 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node27693 = (inp[11]) ? 4'b0000 : 4'b0001;
												assign node27696 = (inp[2]) ? node27704 : node27697;
													assign node27697 = (inp[1]) ? node27701 : node27698;
														assign node27698 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node27701 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node27704 = (inp[1]) ? node27708 : node27705;
														assign node27705 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node27708 = (inp[11]) ? 4'b0000 : 4'b0001;
											assign node27711 = (inp[2]) ? node27727 : node27712;
												assign node27712 = (inp[13]) ? node27720 : node27713;
													assign node27713 = (inp[1]) ? node27717 : node27714;
														assign node27714 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node27717 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node27720 = (inp[1]) ? node27724 : node27721;
														assign node27721 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node27724 = (inp[11]) ? 4'b0000 : 4'b0001;
												assign node27727 = (inp[9]) ? node27735 : node27728;
													assign node27728 = (inp[11]) ? node27732 : node27729;
														assign node27729 = (inp[1]) ? 4'b0001 : 4'b0000;
														assign node27732 = (inp[1]) ? 4'b0000 : 4'b0001;
													assign node27735 = (inp[10]) ? node27743 : node27736;
														assign node27736 = (inp[11]) ? node27740 : node27737;
															assign node27737 = (inp[1]) ? 4'b0001 : 4'b0000;
															assign node27740 = (inp[13]) ? 4'b0001 : 4'b0000;
														assign node27743 = (inp[1]) ? node27745 : 4'b0001;
															assign node27745 = (inp[11]) ? 4'b0000 : 4'b0001;
										assign node27748 = (inp[0]) ? node27812 : node27749;
											assign node27749 = (inp[13]) ? node27789 : node27750;
												assign node27750 = (inp[1]) ? node27766 : node27751;
													assign node27751 = (inp[9]) ? node27759 : node27752;
														assign node27752 = (inp[11]) ? node27756 : node27753;
															assign node27753 = (inp[2]) ? 4'b0001 : 4'b0000;
															assign node27756 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node27759 = (inp[11]) ? node27763 : node27760;
															assign node27760 = (inp[2]) ? 4'b0001 : 4'b0000;
															assign node27763 = (inp[2]) ? 4'b0000 : 4'b0001;
													assign node27766 = (inp[9]) ? node27774 : node27767;
														assign node27767 = (inp[11]) ? node27771 : node27768;
															assign node27768 = (inp[2]) ? 4'b0000 : 4'b0001;
															assign node27771 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node27774 = (inp[10]) ? node27782 : node27775;
															assign node27775 = (inp[11]) ? node27779 : node27776;
																assign node27776 = (inp[2]) ? 4'b0000 : 4'b0001;
																assign node27779 = (inp[2]) ? 4'b0001 : 4'b0000;
															assign node27782 = (inp[11]) ? node27786 : node27783;
																assign node27783 = (inp[2]) ? 4'b0000 : 4'b0001;
																assign node27786 = (inp[2]) ? 4'b0001 : 4'b0000;
												assign node27789 = (inp[2]) ? node27805 : node27790;
													assign node27790 = (inp[9]) ? node27798 : node27791;
														assign node27791 = (inp[1]) ? node27795 : node27792;
															assign node27792 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node27795 = (inp[11]) ? 4'b0000 : 4'b0001;
														assign node27798 = (inp[11]) ? node27802 : node27799;
															assign node27799 = (inp[1]) ? 4'b0001 : 4'b0000;
															assign node27802 = (inp[1]) ? 4'b0000 : 4'b0001;
													assign node27805 = (inp[11]) ? node27809 : node27806;
														assign node27806 = (inp[1]) ? 4'b0000 : 4'b0001;
														assign node27809 = (inp[1]) ? 4'b0001 : 4'b0000;
											assign node27812 = (inp[13]) ? node27852 : node27813;
												assign node27813 = (inp[10]) ? node27829 : node27814;
													assign node27814 = (inp[11]) ? node27822 : node27815;
														assign node27815 = (inp[2]) ? node27819 : node27816;
															assign node27816 = (inp[1]) ? 4'b0001 : 4'b0000;
															assign node27819 = (inp[1]) ? 4'b0000 : 4'b0001;
														assign node27822 = (inp[2]) ? node27826 : node27823;
															assign node27823 = (inp[1]) ? 4'b0000 : 4'b0001;
															assign node27826 = (inp[1]) ? 4'b0001 : 4'b0000;
													assign node27829 = (inp[2]) ? node27845 : node27830;
														assign node27830 = (inp[9]) ? node27838 : node27831;
															assign node27831 = (inp[11]) ? node27835 : node27832;
																assign node27832 = (inp[1]) ? 4'b0001 : 4'b0000;
																assign node27835 = (inp[1]) ? 4'b0000 : 4'b0001;
															assign node27838 = (inp[1]) ? node27842 : node27839;
																assign node27839 = (inp[11]) ? 4'b0001 : 4'b0000;
																assign node27842 = (inp[11]) ? 4'b0000 : 4'b0001;
														assign node27845 = (inp[11]) ? node27849 : node27846;
															assign node27846 = (inp[1]) ? 4'b0000 : 4'b0001;
															assign node27849 = (inp[1]) ? 4'b0001 : 4'b0000;
												assign node27852 = (inp[9]) ? node27868 : node27853;
													assign node27853 = (inp[2]) ? node27861 : node27854;
														assign node27854 = (inp[1]) ? node27858 : node27855;
															assign node27855 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node27858 = (inp[11]) ? 4'b0000 : 4'b0001;
														assign node27861 = (inp[11]) ? node27865 : node27862;
															assign node27862 = (inp[1]) ? 4'b0000 : 4'b0001;
															assign node27865 = (inp[1]) ? 4'b0001 : 4'b0000;
													assign node27868 = (inp[2]) ? node27874 : node27869;
														assign node27869 = (inp[11]) ? 4'b0000 : node27870;
															assign node27870 = (inp[1]) ? 4'b0001 : 4'b0000;
														assign node27874 = (inp[11]) ? node27878 : node27875;
															assign node27875 = (inp[1]) ? 4'b0000 : 4'b0001;
															assign node27878 = (inp[1]) ? 4'b0001 : 4'b0000;
									assign node27881 = (inp[11]) ? node27893 : node27882;
										assign node27882 = (inp[1]) ? node27888 : node27883;
											assign node27883 = (inp[7]) ? 4'b0100 : node27884;
												assign node27884 = (inp[2]) ? 4'b0101 : 4'b0100;
											assign node27888 = (inp[2]) ? node27890 : 4'b0101;
												assign node27890 = (inp[7]) ? 4'b0101 : 4'b0100;
										assign node27893 = (inp[1]) ? node27899 : node27894;
											assign node27894 = (inp[2]) ? node27896 : 4'b0101;
												assign node27896 = (inp[7]) ? 4'b0101 : 4'b0100;
											assign node27899 = (inp[2]) ? node27901 : 4'b0100;
												assign node27901 = (inp[7]) ? 4'b0100 : 4'b0101;
								assign node27904 = (inp[13]) ? node27912 : node27905;
									assign node27905 = (inp[7]) ? node27909 : node27906;
										assign node27906 = (inp[11]) ? 4'b0101 : 4'b0100;
										assign node27909 = (inp[11]) ? 4'b0100 : 4'b0101;
									assign node27912 = (inp[10]) ? node27994 : node27913;
										assign node27913 = (inp[1]) ? node27953 : node27914;
											assign node27914 = (inp[4]) ? node27930 : node27915;
												assign node27915 = (inp[0]) ? node27923 : node27916;
													assign node27916 = (inp[7]) ? node27920 : node27917;
														assign node27917 = (inp[11]) ? 4'b0101 : 4'b0100;
														assign node27920 = (inp[11]) ? 4'b0100 : 4'b0101;
													assign node27923 = (inp[11]) ? node27927 : node27924;
														assign node27924 = (inp[7]) ? 4'b0101 : 4'b0100;
														assign node27927 = (inp[7]) ? 4'b0100 : 4'b0101;
												assign node27930 = (inp[0]) ? node27946 : node27931;
													assign node27931 = (inp[9]) ? node27939 : node27932;
														assign node27932 = (inp[7]) ? node27936 : node27933;
															assign node27933 = (inp[11]) ? 4'b0101 : 4'b0100;
															assign node27936 = (inp[11]) ? 4'b0100 : 4'b0101;
														assign node27939 = (inp[11]) ? node27943 : node27940;
															assign node27940 = (inp[7]) ? 4'b0101 : 4'b0100;
															assign node27943 = (inp[7]) ? 4'b0100 : 4'b0101;
													assign node27946 = (inp[11]) ? node27950 : node27947;
														assign node27947 = (inp[7]) ? 4'b0101 : 4'b0100;
														assign node27950 = (inp[7]) ? 4'b0100 : 4'b0101;
											assign node27953 = (inp[9]) ? node27979 : node27954;
												assign node27954 = (inp[4]) ? node27962 : node27955;
													assign node27955 = (inp[7]) ? node27959 : node27956;
														assign node27956 = (inp[11]) ? 4'b0101 : 4'b0100;
														assign node27959 = (inp[11]) ? 4'b0100 : 4'b0101;
													assign node27962 = (inp[0]) ? node27970 : node27963;
														assign node27963 = (inp[2]) ? 4'b0100 : node27964;
															assign node27964 = (inp[7]) ? node27966 : 4'b0100;
																assign node27966 = (inp[11]) ? 4'b0100 : 4'b0101;
														assign node27970 = (inp[2]) ? node27972 : 4'b0100;
															assign node27972 = (inp[11]) ? node27976 : node27973;
																assign node27973 = (inp[7]) ? 4'b0101 : 4'b0100;
																assign node27976 = (inp[7]) ? 4'b0100 : 4'b0101;
												assign node27979 = (inp[2]) ? node27987 : node27980;
													assign node27980 = (inp[11]) ? node27984 : node27981;
														assign node27981 = (inp[7]) ? 4'b0101 : 4'b0100;
														assign node27984 = (inp[7]) ? 4'b0100 : 4'b0101;
													assign node27987 = (inp[11]) ? node27991 : node27988;
														assign node27988 = (inp[7]) ? 4'b0101 : 4'b0100;
														assign node27991 = (inp[7]) ? 4'b0100 : 4'b0101;
										assign node27994 = (inp[4]) ? node28048 : node27995;
											assign node27995 = (inp[9]) ? node28041 : node27996;
												assign node27996 = (inp[1]) ? node28028 : node27997;
													assign node27997 = (inp[2]) ? node28013 : node27998;
														assign node27998 = (inp[0]) ? node28006 : node27999;
															assign node27999 = (inp[7]) ? node28003 : node28000;
																assign node28000 = (inp[11]) ? 4'b0101 : 4'b0100;
																assign node28003 = (inp[11]) ? 4'b0100 : 4'b0101;
															assign node28006 = (inp[11]) ? node28010 : node28007;
																assign node28007 = (inp[7]) ? 4'b0101 : 4'b0100;
																assign node28010 = (inp[7]) ? 4'b0100 : 4'b0101;
														assign node28013 = (inp[0]) ? node28021 : node28014;
															assign node28014 = (inp[11]) ? node28018 : node28015;
																assign node28015 = (inp[7]) ? 4'b0101 : 4'b0100;
																assign node28018 = (inp[7]) ? 4'b0100 : 4'b0101;
															assign node28021 = (inp[11]) ? node28025 : node28022;
																assign node28022 = (inp[7]) ? 4'b0101 : 4'b0100;
																assign node28025 = (inp[7]) ? 4'b0100 : 4'b0101;
													assign node28028 = (inp[2]) ? node28034 : node28029;
														assign node28029 = (inp[7]) ? 4'b0101 : node28030;
															assign node28030 = (inp[11]) ? 4'b0101 : 4'b0100;
														assign node28034 = (inp[7]) ? node28038 : node28035;
															assign node28035 = (inp[11]) ? 4'b0101 : 4'b0100;
															assign node28038 = (inp[11]) ? 4'b0100 : 4'b0101;
												assign node28041 = (inp[7]) ? node28045 : node28042;
													assign node28042 = (inp[11]) ? 4'b0101 : 4'b0100;
													assign node28045 = (inp[11]) ? 4'b0100 : 4'b0101;
											assign node28048 = (inp[7]) ? node28052 : node28049;
												assign node28049 = (inp[11]) ? 4'b0101 : 4'b0100;
												assign node28052 = (inp[11]) ? 4'b0100 : 4'b0101;
							assign node28055 = (inp[12]) ? node28331 : node28056;
								assign node28056 = (inp[4]) ? node28200 : node28057;
									assign node28057 = (inp[9]) ? node28081 : node28058;
										assign node28058 = (inp[1]) ? node28070 : node28059;
											assign node28059 = (inp[11]) ? node28065 : node28060;
												assign node28060 = (inp[2]) ? 4'b0100 : node28061;
													assign node28061 = (inp[7]) ? 4'b0101 : 4'b0100;
												assign node28065 = (inp[7]) ? node28067 : 4'b0101;
													assign node28067 = (inp[2]) ? 4'b0101 : 4'b0100;
											assign node28070 = (inp[11]) ? node28076 : node28071;
												assign node28071 = (inp[2]) ? 4'b0101 : node28072;
													assign node28072 = (inp[7]) ? 4'b0100 : 4'b0101;
												assign node28076 = (inp[7]) ? node28078 : 4'b0100;
													assign node28078 = (inp[2]) ? 4'b0100 : 4'b0101;
										assign node28081 = (inp[13]) ? node28105 : node28082;
											assign node28082 = (inp[11]) ? node28094 : node28083;
												assign node28083 = (inp[1]) ? node28089 : node28084;
													assign node28084 = (inp[2]) ? 4'b0100 : node28085;
														assign node28085 = (inp[7]) ? 4'b0101 : 4'b0100;
													assign node28089 = (inp[2]) ? 4'b0101 : node28090;
														assign node28090 = (inp[7]) ? 4'b0100 : 4'b0101;
												assign node28094 = (inp[1]) ? node28100 : node28095;
													assign node28095 = (inp[7]) ? node28097 : 4'b0101;
														assign node28097 = (inp[2]) ? 4'b0101 : 4'b0100;
													assign node28100 = (inp[7]) ? node28102 : 4'b0100;
														assign node28102 = (inp[2]) ? 4'b0100 : 4'b0101;
											assign node28105 = (inp[0]) ? node28145 : node28106;
												assign node28106 = (inp[7]) ? node28122 : node28107;
													assign node28107 = (inp[10]) ? node28115 : node28108;
														assign node28108 = (inp[11]) ? node28112 : node28109;
															assign node28109 = (inp[1]) ? 4'b0101 : 4'b0100;
															assign node28112 = (inp[1]) ? 4'b0100 : 4'b0101;
														assign node28115 = (inp[1]) ? node28119 : node28116;
															assign node28116 = (inp[11]) ? 4'b0101 : 4'b0100;
															assign node28119 = (inp[11]) ? 4'b0100 : 4'b0101;
													assign node28122 = (inp[10]) ? node28132 : node28123;
														assign node28123 = (inp[2]) ? 4'b0100 : node28124;
															assign node28124 = (inp[1]) ? node28128 : node28125;
																assign node28125 = (inp[11]) ? 4'b0100 : 4'b0101;
																assign node28128 = (inp[11]) ? 4'b0101 : 4'b0100;
														assign node28132 = (inp[2]) ? node28138 : node28133;
															assign node28133 = (inp[11]) ? 4'b0100 : node28134;
																assign node28134 = (inp[1]) ? 4'b0100 : 4'b0101;
															assign node28138 = (inp[11]) ? node28142 : node28139;
																assign node28139 = (inp[1]) ? 4'b0101 : 4'b0100;
																assign node28142 = (inp[1]) ? 4'b0100 : 4'b0101;
												assign node28145 = (inp[2]) ? node28177 : node28146;
													assign node28146 = (inp[10]) ? node28162 : node28147;
														assign node28147 = (inp[7]) ? node28155 : node28148;
															assign node28148 = (inp[11]) ? node28152 : node28149;
																assign node28149 = (inp[1]) ? 4'b0101 : 4'b0100;
																assign node28152 = (inp[1]) ? 4'b0100 : 4'b0101;
															assign node28155 = (inp[1]) ? node28159 : node28156;
																assign node28156 = (inp[11]) ? 4'b0100 : 4'b0101;
																assign node28159 = (inp[11]) ? 4'b0101 : 4'b0100;
														assign node28162 = (inp[11]) ? node28170 : node28163;
															assign node28163 = (inp[1]) ? node28167 : node28164;
																assign node28164 = (inp[7]) ? 4'b0101 : 4'b0100;
																assign node28167 = (inp[7]) ? 4'b0100 : 4'b0101;
															assign node28170 = (inp[1]) ? node28174 : node28171;
																assign node28171 = (inp[7]) ? 4'b0100 : 4'b0101;
																assign node28174 = (inp[7]) ? 4'b0101 : 4'b0100;
													assign node28177 = (inp[7]) ? node28185 : node28178;
														assign node28178 = (inp[1]) ? node28182 : node28179;
															assign node28179 = (inp[11]) ? 4'b0101 : 4'b0100;
															assign node28182 = (inp[11]) ? 4'b0100 : 4'b0101;
														assign node28185 = (inp[10]) ? node28193 : node28186;
															assign node28186 = (inp[11]) ? node28190 : node28187;
																assign node28187 = (inp[1]) ? 4'b0101 : 4'b0100;
																assign node28190 = (inp[1]) ? 4'b0100 : 4'b0101;
															assign node28193 = (inp[1]) ? node28197 : node28194;
																assign node28194 = (inp[11]) ? 4'b0101 : 4'b0100;
																assign node28197 = (inp[11]) ? 4'b0100 : 4'b0101;
									assign node28200 = (inp[9]) ? node28248 : node28201;
										assign node28201 = (inp[10]) ? node28225 : node28202;
											assign node28202 = (inp[1]) ? node28214 : node28203;
												assign node28203 = (inp[11]) ? node28209 : node28204;
													assign node28204 = (inp[7]) ? 4'b0000 : node28205;
														assign node28205 = (inp[2]) ? 4'b0000 : 4'b0001;
													assign node28209 = (inp[2]) ? 4'b0001 : node28210;
														assign node28210 = (inp[7]) ? 4'b0001 : 4'b0000;
												assign node28214 = (inp[11]) ? node28220 : node28215;
													assign node28215 = (inp[2]) ? 4'b0001 : node28216;
														assign node28216 = (inp[7]) ? 4'b0001 : 4'b0000;
													assign node28220 = (inp[2]) ? 4'b0000 : node28221;
														assign node28221 = (inp[7]) ? 4'b0000 : 4'b0001;
											assign node28225 = (inp[1]) ? node28237 : node28226;
												assign node28226 = (inp[11]) ? node28232 : node28227;
													assign node28227 = (inp[2]) ? 4'b0000 : node28228;
														assign node28228 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node28232 = (inp[2]) ? 4'b0001 : node28233;
														assign node28233 = (inp[7]) ? 4'b0001 : 4'b0000;
												assign node28237 = (inp[11]) ? node28243 : node28238;
													assign node28238 = (inp[2]) ? 4'b0001 : node28239;
														assign node28239 = (inp[7]) ? 4'b0001 : 4'b0000;
													assign node28243 = (inp[2]) ? 4'b0000 : node28244;
														assign node28244 = (inp[7]) ? 4'b0000 : 4'b0001;
										assign node28248 = (inp[0]) ? node28312 : node28249;
											assign node28249 = (inp[2]) ? node28297 : node28250;
												assign node28250 = (inp[13]) ? node28274 : node28251;
													assign node28251 = (inp[10]) ? node28261 : node28252;
														assign node28252 = (inp[1]) ? node28254 : 4'b0001;
															assign node28254 = (inp[7]) ? node28258 : node28255;
																assign node28255 = (inp[11]) ? 4'b0001 : 4'b0000;
																assign node28258 = (inp[11]) ? 4'b0000 : 4'b0001;
														assign node28261 = (inp[7]) ? node28269 : node28262;
															assign node28262 = (inp[11]) ? node28266 : node28263;
																assign node28263 = (inp[1]) ? 4'b0000 : 4'b0001;
																assign node28266 = (inp[1]) ? 4'b0001 : 4'b0000;
															assign node28269 = (inp[1]) ? node28271 : 4'b0000;
																assign node28271 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node28274 = (inp[10]) ? node28282 : node28275;
														assign node28275 = (inp[1]) ? 4'b0000 : node28276;
															assign node28276 = (inp[11]) ? node28278 : 4'b0000;
																assign node28278 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node28282 = (inp[1]) ? node28290 : node28283;
															assign node28283 = (inp[11]) ? node28287 : node28284;
																assign node28284 = (inp[7]) ? 4'b0000 : 4'b0001;
																assign node28287 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node28290 = (inp[7]) ? node28294 : node28291;
																assign node28291 = (inp[11]) ? 4'b0001 : 4'b0000;
																assign node28294 = (inp[11]) ? 4'b0000 : 4'b0001;
												assign node28297 = (inp[7]) ? node28305 : node28298;
													assign node28298 = (inp[11]) ? node28302 : node28299;
														assign node28299 = (inp[1]) ? 4'b0001 : 4'b0000;
														assign node28302 = (inp[1]) ? 4'b0000 : 4'b0001;
													assign node28305 = (inp[1]) ? node28309 : node28306;
														assign node28306 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node28309 = (inp[11]) ? 4'b0000 : 4'b0001;
											assign node28312 = (inp[11]) ? node28320 : node28313;
												assign node28313 = (inp[1]) ? node28315 : 4'b0000;
													assign node28315 = (inp[2]) ? 4'b0001 : node28316;
														assign node28316 = (inp[7]) ? 4'b0001 : 4'b0000;
												assign node28320 = (inp[1]) ? node28326 : node28321;
													assign node28321 = (inp[7]) ? 4'b0001 : node28322;
														assign node28322 = (inp[2]) ? 4'b0001 : 4'b0000;
													assign node28326 = (inp[2]) ? 4'b0000 : node28327;
														assign node28327 = (inp[7]) ? 4'b0000 : 4'b0001;
								assign node28331 = (inp[11]) ? node28337 : node28332;
									assign node28332 = (inp[2]) ? 4'b0001 : node28333;
										assign node28333 = (inp[4]) ? 4'b0001 : 4'b0000;
									assign node28337 = (inp[2]) ? 4'b0000 : node28338;
										assign node28338 = (inp[4]) ? 4'b0000 : 4'b0001;
		assign node28342 = (inp[6]) ? node45374 : node28343;
			assign node28343 = (inp[3]) ? node37603 : node28344;
				assign node28344 = (inp[12]) ? node32842 : node28345;
					assign node28345 = (inp[4]) ? node30479 : node28346;
						assign node28346 = (inp[8]) ? node29776 : node28347;
							assign node28347 = (inp[13]) ? node29059 : node28348;
								assign node28348 = (inp[2]) ? node28716 : node28349;
									assign node28349 = (inp[5]) ? node28535 : node28350;
										assign node28350 = (inp[1]) ? node28442 : node28351;
											assign node28351 = (inp[7]) ? node28395 : node28352;
												assign node28352 = (inp[15]) ? node28372 : node28353;
													assign node28353 = (inp[9]) ? node28365 : node28354;
														assign node28354 = (inp[10]) ? node28360 : node28355;
															assign node28355 = (inp[0]) ? 4'b1000 : node28356;
																assign node28356 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node28360 = (inp[0]) ? 4'b1001 : node28361;
																assign node28361 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node28365 = (inp[10]) ? node28367 : 4'b1001;
															assign node28367 = (inp[11]) ? node28369 : 4'b1000;
																assign node28369 = (inp[0]) ? 4'b1000 : 4'b1001;
													assign node28372 = (inp[9]) ? node28384 : node28373;
														assign node28373 = (inp[10]) ? node28379 : node28374;
															assign node28374 = (inp[0]) ? 4'b1010 : node28375;
																assign node28375 = (inp[11]) ? 4'b1011 : 4'b1010;
															assign node28379 = (inp[11]) ? node28381 : 4'b1011;
																assign node28381 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node28384 = (inp[10]) ? node28390 : node28385;
															assign node28385 = (inp[0]) ? 4'b1011 : node28386;
																assign node28386 = (inp[11]) ? 4'b1010 : 4'b1011;
															assign node28390 = (inp[0]) ? 4'b1010 : node28391;
																assign node28391 = (inp[11]) ? 4'b1011 : 4'b1010;
												assign node28395 = (inp[15]) ? node28425 : node28396;
													assign node28396 = (inp[11]) ? node28410 : node28397;
														assign node28397 = (inp[0]) ? node28405 : node28398;
															assign node28398 = (inp[9]) ? node28402 : node28399;
																assign node28399 = (inp[10]) ? 4'b1011 : 4'b1010;
																assign node28402 = (inp[10]) ? 4'b1010 : 4'b1011;
															assign node28405 = (inp[10]) ? node28407 : 4'b1011;
																assign node28407 = (inp[9]) ? 4'b1010 : 4'b1011;
														assign node28410 = (inp[9]) ? node28418 : node28411;
															assign node28411 = (inp[0]) ? node28415 : node28412;
																assign node28412 = (inp[10]) ? 4'b1010 : 4'b1011;
																assign node28415 = (inp[10]) ? 4'b1011 : 4'b1010;
															assign node28418 = (inp[10]) ? node28422 : node28419;
																assign node28419 = (inp[0]) ? 4'b1011 : 4'b1010;
																assign node28422 = (inp[0]) ? 4'b1010 : 4'b1011;
													assign node28425 = (inp[0]) ? node28435 : node28426;
														assign node28426 = (inp[10]) ? 4'b1101 : node28427;
															assign node28427 = (inp[11]) ? node28431 : node28428;
																assign node28428 = (inp[9]) ? 4'b1101 : 4'b1100;
																assign node28431 = (inp[9]) ? 4'b1100 : 4'b1101;
														assign node28435 = (inp[9]) ? node28439 : node28436;
															assign node28436 = (inp[10]) ? 4'b1101 : 4'b1100;
															assign node28439 = (inp[10]) ? 4'b1100 : 4'b1101;
											assign node28442 = (inp[15]) ? node28488 : node28443;
												assign node28443 = (inp[7]) ? node28467 : node28444;
													assign node28444 = (inp[11]) ? node28452 : node28445;
														assign node28445 = (inp[9]) ? node28449 : node28446;
															assign node28446 = (inp[10]) ? 4'b1001 : 4'b1000;
															assign node28449 = (inp[10]) ? 4'b1000 : 4'b1001;
														assign node28452 = (inp[9]) ? node28460 : node28453;
															assign node28453 = (inp[10]) ? node28457 : node28454;
																assign node28454 = (inp[0]) ? 4'b1000 : 4'b1001;
																assign node28457 = (inp[0]) ? 4'b1001 : 4'b1000;
															assign node28460 = (inp[0]) ? node28464 : node28461;
																assign node28461 = (inp[10]) ? 4'b1001 : 4'b1000;
																assign node28464 = (inp[10]) ? 4'b1000 : 4'b1001;
													assign node28467 = (inp[9]) ? node28477 : node28468;
														assign node28468 = (inp[10]) ? node28474 : node28469;
															assign node28469 = (inp[0]) ? 4'b1010 : node28470;
																assign node28470 = (inp[11]) ? 4'b1011 : 4'b1010;
															assign node28474 = (inp[11]) ? 4'b1010 : 4'b1011;
														assign node28477 = (inp[10]) ? node28483 : node28478;
															assign node28478 = (inp[0]) ? 4'b1011 : node28479;
																assign node28479 = (inp[11]) ? 4'b1010 : 4'b1011;
															assign node28483 = (inp[0]) ? 4'b1010 : node28484;
																assign node28484 = (inp[11]) ? 4'b1011 : 4'b1010;
												assign node28488 = (inp[7]) ? node28512 : node28489;
													assign node28489 = (inp[0]) ? node28503 : node28490;
														assign node28490 = (inp[11]) ? node28496 : node28491;
															assign node28491 = (inp[10]) ? node28493 : 4'b1010;
																assign node28493 = (inp[9]) ? 4'b1010 : 4'b1011;
															assign node28496 = (inp[9]) ? node28500 : node28497;
																assign node28497 = (inp[10]) ? 4'b1011 : 4'b1010;
																assign node28500 = (inp[10]) ? 4'b1010 : 4'b1011;
														assign node28503 = (inp[11]) ? node28505 : 4'b1011;
															assign node28505 = (inp[10]) ? node28509 : node28506;
																assign node28506 = (inp[9]) ? 4'b1011 : 4'b1010;
																assign node28509 = (inp[9]) ? 4'b1010 : 4'b1011;
													assign node28512 = (inp[0]) ? node28528 : node28513;
														assign node28513 = (inp[10]) ? node28521 : node28514;
															assign node28514 = (inp[11]) ? node28518 : node28515;
																assign node28515 = (inp[9]) ? 4'b1000 : 4'b1001;
																assign node28518 = (inp[9]) ? 4'b1001 : 4'b1000;
															assign node28521 = (inp[11]) ? node28525 : node28522;
																assign node28522 = (inp[9]) ? 4'b1001 : 4'b1000;
																assign node28525 = (inp[9]) ? 4'b1000 : 4'b1001;
														assign node28528 = (inp[9]) ? node28532 : node28529;
															assign node28529 = (inp[10]) ? 4'b1000 : 4'b1001;
															assign node28532 = (inp[10]) ? 4'b1001 : 4'b1000;
										assign node28535 = (inp[1]) ? node28625 : node28536;
											assign node28536 = (inp[10]) ? node28580 : node28537;
												assign node28537 = (inp[0]) ? node28561 : node28538;
													assign node28538 = (inp[11]) ? node28552 : node28539;
														assign node28539 = (inp[15]) ? node28545 : node28540;
															assign node28540 = (inp[7]) ? 4'b1110 : node28541;
																assign node28541 = (inp[9]) ? 4'b1101 : 4'b1100;
															assign node28545 = (inp[7]) ? node28549 : node28546;
																assign node28546 = (inp[9]) ? 4'b1111 : 4'b1110;
																assign node28549 = (inp[9]) ? 4'b1100 : 4'b1101;
														assign node28552 = (inp[9]) ? node28556 : node28553;
															assign node28553 = (inp[15]) ? 4'b1101 : 4'b1110;
															assign node28556 = (inp[7]) ? 4'b1100 : node28557;
																assign node28557 = (inp[15]) ? 4'b1110 : 4'b1100;
													assign node28561 = (inp[9]) ? node28571 : node28562;
														assign node28562 = (inp[7]) ? node28566 : node28563;
															assign node28563 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node28566 = (inp[15]) ? node28568 : 4'b1111;
																assign node28568 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node28571 = (inp[7]) ? node28575 : node28572;
															assign node28572 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node28575 = (inp[15]) ? node28577 : 4'b1110;
																assign node28577 = (inp[11]) ? 4'b1100 : 4'b1101;
												assign node28580 = (inp[11]) ? node28598 : node28581;
													assign node28581 = (inp[7]) ? node28587 : node28582;
														assign node28582 = (inp[15]) ? 4'b1111 : node28583;
															assign node28583 = (inp[9]) ? 4'b1100 : 4'b1101;
														assign node28587 = (inp[15]) ? node28591 : node28588;
															assign node28588 = (inp[9]) ? 4'b1111 : 4'b1110;
															assign node28591 = (inp[9]) ? node28595 : node28592;
																assign node28592 = (inp[0]) ? 4'b1101 : 4'b1100;
																assign node28595 = (inp[0]) ? 4'b1100 : 4'b1101;
													assign node28598 = (inp[9]) ? node28612 : node28599;
														assign node28599 = (inp[7]) ? node28607 : node28600;
															assign node28600 = (inp[0]) ? node28604 : node28601;
																assign node28601 = (inp[15]) ? 4'b1110 : 4'b1100;
																assign node28604 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node28607 = (inp[15]) ? 4'b1100 : node28608;
																assign node28608 = (inp[0]) ? 4'b1110 : 4'b1111;
														assign node28612 = (inp[0]) ? node28620 : node28613;
															assign node28613 = (inp[7]) ? node28617 : node28614;
																assign node28614 = (inp[15]) ? 4'b1111 : 4'b1101;
																assign node28617 = (inp[15]) ? 4'b1101 : 4'b1110;
															assign node28620 = (inp[7]) ? 4'b1101 : node28621;
																assign node28621 = (inp[15]) ? 4'b1110 : 4'b1100;
											assign node28625 = (inp[7]) ? node28669 : node28626;
												assign node28626 = (inp[15]) ? node28648 : node28627;
													assign node28627 = (inp[11]) ? node28641 : node28628;
														assign node28628 = (inp[9]) ? node28636 : node28629;
															assign node28629 = (inp[10]) ? node28633 : node28630;
																assign node28630 = (inp[0]) ? 4'b1001 : 4'b1000;
																assign node28633 = (inp[0]) ? 4'b1000 : 4'b1001;
															assign node28636 = (inp[10]) ? node28638 : 4'b1001;
																assign node28638 = (inp[0]) ? 4'b1001 : 4'b1000;
														assign node28641 = (inp[10]) ? node28645 : node28642;
															assign node28642 = (inp[9]) ? 4'b1001 : 4'b1000;
															assign node28645 = (inp[9]) ? 4'b1000 : 4'b1001;
													assign node28648 = (inp[11]) ? node28654 : node28649;
														assign node28649 = (inp[10]) ? 4'b1010 : node28650;
															assign node28650 = (inp[9]) ? 4'b1010 : 4'b1011;
														assign node28654 = (inp[0]) ? node28662 : node28655;
															assign node28655 = (inp[10]) ? node28659 : node28656;
																assign node28656 = (inp[9]) ? 4'b1011 : 4'b1010;
																assign node28659 = (inp[9]) ? 4'b1010 : 4'b1011;
															assign node28662 = (inp[9]) ? node28666 : node28663;
																assign node28663 = (inp[10]) ? 4'b1010 : 4'b1011;
																assign node28666 = (inp[10]) ? 4'b1011 : 4'b1010;
												assign node28669 = (inp[15]) ? node28689 : node28670;
													assign node28670 = (inp[9]) ? node28678 : node28671;
														assign node28671 = (inp[10]) ? 4'b1010 : node28672;
															assign node28672 = (inp[0]) ? node28674 : 4'b1011;
																assign node28674 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node28678 = (inp[10]) ? node28684 : node28679;
															assign node28679 = (inp[11]) ? 4'b1010 : node28680;
																assign node28680 = (inp[0]) ? 4'b1011 : 4'b1010;
															assign node28684 = (inp[11]) ? 4'b1011 : node28685;
																assign node28685 = (inp[0]) ? 4'b1010 : 4'b1011;
													assign node28689 = (inp[11]) ? node28701 : node28690;
														assign node28690 = (inp[0]) ? node28696 : node28691;
															assign node28691 = (inp[9]) ? 4'b1100 : node28692;
																assign node28692 = (inp[10]) ? 4'b1101 : 4'b1100;
															assign node28696 = (inp[10]) ? 4'b1100 : node28697;
																assign node28697 = (inp[9]) ? 4'b1101 : 4'b1100;
														assign node28701 = (inp[0]) ? node28709 : node28702;
															assign node28702 = (inp[9]) ? node28706 : node28703;
																assign node28703 = (inp[10]) ? 4'b1100 : 4'b1101;
																assign node28706 = (inp[10]) ? 4'b1101 : 4'b1100;
															assign node28709 = (inp[10]) ? node28713 : node28710;
																assign node28710 = (inp[9]) ? 4'b1101 : 4'b1100;
																assign node28713 = (inp[9]) ? 4'b1100 : 4'b1101;
									assign node28716 = (inp[5]) ? node28878 : node28717;
										assign node28717 = (inp[15]) ? node28795 : node28718;
											assign node28718 = (inp[7]) ? node28772 : node28719;
												assign node28719 = (inp[0]) ? node28749 : node28720;
													assign node28720 = (inp[11]) ? node28734 : node28721;
														assign node28721 = (inp[1]) ? node28729 : node28722;
															assign node28722 = (inp[10]) ? node28726 : node28723;
																assign node28723 = (inp[9]) ? 4'b1101 : 4'b1100;
																assign node28726 = (inp[9]) ? 4'b1100 : 4'b1101;
															assign node28729 = (inp[9]) ? node28731 : 4'b1101;
																assign node28731 = (inp[10]) ? 4'b1100 : 4'b1101;
														assign node28734 = (inp[1]) ? node28742 : node28735;
															assign node28735 = (inp[10]) ? node28739 : node28736;
																assign node28736 = (inp[9]) ? 4'b1101 : 4'b1100;
																assign node28739 = (inp[9]) ? 4'b1100 : 4'b1101;
															assign node28742 = (inp[9]) ? node28746 : node28743;
																assign node28743 = (inp[10]) ? 4'b1101 : 4'b1100;
																assign node28746 = (inp[10]) ? 4'b1100 : 4'b1101;
													assign node28749 = (inp[9]) ? node28757 : node28750;
														assign node28750 = (inp[11]) ? node28754 : node28751;
															assign node28751 = (inp[10]) ? 4'b1100 : 4'b1101;
															assign node28754 = (inp[10]) ? 4'b1101 : 4'b1100;
														assign node28757 = (inp[1]) ? node28765 : node28758;
															assign node28758 = (inp[10]) ? node28762 : node28759;
																assign node28759 = (inp[11]) ? 4'b1101 : 4'b1100;
																assign node28762 = (inp[11]) ? 4'b1100 : 4'b1101;
															assign node28765 = (inp[10]) ? node28769 : node28766;
																assign node28766 = (inp[11]) ? 4'b1101 : 4'b1100;
																assign node28769 = (inp[11]) ? 4'b1100 : 4'b1101;
												assign node28772 = (inp[10]) ? node28784 : node28773;
													assign node28773 = (inp[9]) ? node28779 : node28774;
														assign node28774 = (inp[0]) ? node28776 : 4'b1110;
															assign node28776 = (inp[11]) ? 4'b1110 : 4'b1111;
														assign node28779 = (inp[11]) ? 4'b1111 : node28780;
															assign node28780 = (inp[0]) ? 4'b1110 : 4'b1111;
													assign node28784 = (inp[9]) ? node28790 : node28785;
														assign node28785 = (inp[0]) ? node28787 : 4'b1111;
															assign node28787 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node28790 = (inp[0]) ? node28792 : 4'b1110;
															assign node28792 = (inp[11]) ? 4'b1110 : 4'b1111;
											assign node28795 = (inp[7]) ? node28829 : node28796;
												assign node28796 = (inp[11]) ? node28816 : node28797;
													assign node28797 = (inp[9]) ? node28807 : node28798;
														assign node28798 = (inp[10]) ? node28804 : node28799;
															assign node28799 = (inp[1]) ? 4'b1111 : node28800;
																assign node28800 = (inp[0]) ? 4'b1111 : 4'b1110;
															assign node28804 = (inp[1]) ? 4'b1110 : 4'b1111;
														assign node28807 = (inp[10]) ? node28813 : node28808;
															assign node28808 = (inp[0]) ? 4'b1110 : node28809;
																assign node28809 = (inp[1]) ? 4'b1110 : 4'b1111;
															assign node28813 = (inp[0]) ? 4'b1111 : 4'b1110;
													assign node28816 = (inp[10]) ? node28824 : node28817;
														assign node28817 = (inp[9]) ? 4'b1111 : node28818;
															assign node28818 = (inp[1]) ? node28820 : 4'b1110;
																assign node28820 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node28824 = (inp[9]) ? 4'b1110 : node28825;
															assign node28825 = (inp[1]) ? 4'b1110 : 4'b1111;
												assign node28829 = (inp[1]) ? node28849 : node28830;
													assign node28830 = (inp[0]) ? node28842 : node28831;
														assign node28831 = (inp[10]) ? node28837 : node28832;
															assign node28832 = (inp[11]) ? node28834 : 4'b1000;
																assign node28834 = (inp[9]) ? 4'b1001 : 4'b1000;
															assign node28837 = (inp[11]) ? node28839 : 4'b1001;
																assign node28839 = (inp[9]) ? 4'b1000 : 4'b1001;
														assign node28842 = (inp[9]) ? node28846 : node28843;
															assign node28843 = (inp[10]) ? 4'b1000 : 4'b1001;
															assign node28846 = (inp[10]) ? 4'b1001 : 4'b1000;
													assign node28849 = (inp[11]) ? node28863 : node28850;
														assign node28850 = (inp[10]) ? node28858 : node28851;
															assign node28851 = (inp[9]) ? node28855 : node28852;
																assign node28852 = (inp[0]) ? 4'b1100 : 4'b1101;
																assign node28855 = (inp[0]) ? 4'b1101 : 4'b1100;
															assign node28858 = (inp[9]) ? node28860 : 4'b1100;
																assign node28860 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node28863 = (inp[0]) ? node28871 : node28864;
															assign node28864 = (inp[9]) ? node28868 : node28865;
																assign node28865 = (inp[10]) ? 4'b1100 : 4'b1101;
																assign node28868 = (inp[10]) ? 4'b1101 : 4'b1100;
															assign node28871 = (inp[9]) ? node28875 : node28872;
																assign node28872 = (inp[10]) ? 4'b1100 : 4'b1101;
																assign node28875 = (inp[10]) ? 4'b1101 : 4'b1100;
										assign node28878 = (inp[1]) ? node28968 : node28879;
											assign node28879 = (inp[0]) ? node28933 : node28880;
												assign node28880 = (inp[9]) ? node28910 : node28881;
													assign node28881 = (inp[10]) ? node28895 : node28882;
														assign node28882 = (inp[15]) ? node28890 : node28883;
															assign node28883 = (inp[7]) ? node28887 : node28884;
																assign node28884 = (inp[11]) ? 4'b1000 : 4'b1001;
																assign node28887 = (inp[11]) ? 4'b1011 : 4'b1010;
															assign node28890 = (inp[7]) ? 4'b1000 : node28891;
																assign node28891 = (inp[11]) ? 4'b1010 : 4'b1011;
														assign node28895 = (inp[11]) ? node28903 : node28896;
															assign node28896 = (inp[7]) ? node28900 : node28897;
																assign node28897 = (inp[15]) ? 4'b1010 : 4'b1000;
																assign node28900 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node28903 = (inp[7]) ? node28907 : node28904;
																assign node28904 = (inp[15]) ? 4'b1011 : 4'b1001;
																assign node28907 = (inp[15]) ? 4'b1001 : 4'b1010;
													assign node28910 = (inp[10]) ? node28922 : node28911;
														assign node28911 = (inp[7]) ? node28919 : node28912;
															assign node28912 = (inp[15]) ? node28916 : node28913;
																assign node28913 = (inp[11]) ? 4'b1001 : 4'b1000;
																assign node28916 = (inp[11]) ? 4'b1011 : 4'b1010;
															assign node28919 = (inp[15]) ? 4'b1001 : 4'b1011;
														assign node28922 = (inp[7]) ? node28928 : node28923;
															assign node28923 = (inp[11]) ? 4'b1000 : node28924;
																assign node28924 = (inp[15]) ? 4'b1011 : 4'b1001;
															assign node28928 = (inp[15]) ? 4'b1000 : node28929;
																assign node28929 = (inp[11]) ? 4'b1011 : 4'b1010;
												assign node28933 = (inp[9]) ? node28953 : node28934;
													assign node28934 = (inp[10]) ? node28944 : node28935;
														assign node28935 = (inp[7]) ? node28939 : node28936;
															assign node28936 = (inp[15]) ? 4'b1011 : 4'b1001;
															assign node28939 = (inp[15]) ? node28941 : 4'b1010;
																assign node28941 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node28944 = (inp[7]) ? node28948 : node28945;
															assign node28945 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node28948 = (inp[15]) ? node28950 : 4'b1011;
																assign node28950 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node28953 = (inp[15]) ? node28961 : node28954;
														assign node28954 = (inp[7]) ? node28958 : node28955;
															assign node28955 = (inp[10]) ? 4'b1001 : 4'b1000;
															assign node28958 = (inp[10]) ? 4'b1010 : 4'b1011;
														assign node28961 = (inp[7]) ? node28963 : 4'b1010;
															assign node28963 = (inp[10]) ? node28965 : 4'b1000;
																assign node28965 = (inp[11]) ? 4'b1000 : 4'b1001;
											assign node28968 = (inp[15]) ? node29014 : node28969;
												assign node28969 = (inp[7]) ? node28991 : node28970;
													assign node28970 = (inp[11]) ? node28978 : node28971;
														assign node28971 = (inp[9]) ? node28975 : node28972;
															assign node28972 = (inp[10]) ? 4'b1100 : 4'b1101;
															assign node28975 = (inp[10]) ? 4'b1101 : 4'b1100;
														assign node28978 = (inp[10]) ? node28986 : node28979;
															assign node28979 = (inp[0]) ? node28983 : node28980;
																assign node28980 = (inp[9]) ? 4'b1101 : 4'b1100;
																assign node28983 = (inp[9]) ? 4'b1100 : 4'b1101;
															assign node28986 = (inp[0]) ? node28988 : 4'b1101;
																assign node28988 = (inp[9]) ? 4'b1101 : 4'b1100;
													assign node28991 = (inp[10]) ? node29003 : node28992;
														assign node28992 = (inp[9]) ? node28998 : node28993;
															assign node28993 = (inp[0]) ? 4'b1110 : node28994;
																assign node28994 = (inp[11]) ? 4'b1111 : 4'b1110;
															assign node28998 = (inp[0]) ? 4'b1111 : node28999;
																assign node28999 = (inp[11]) ? 4'b1110 : 4'b1111;
														assign node29003 = (inp[9]) ? node29009 : node29004;
															assign node29004 = (inp[0]) ? 4'b1111 : node29005;
																assign node29005 = (inp[11]) ? 4'b1110 : 4'b1111;
															assign node29009 = (inp[0]) ? 4'b1110 : node29010;
																assign node29010 = (inp[11]) ? 4'b1111 : 4'b1110;
												assign node29014 = (inp[7]) ? node29036 : node29015;
													assign node29015 = (inp[0]) ? node29023 : node29016;
														assign node29016 = (inp[9]) ? node29020 : node29017;
															assign node29017 = (inp[10]) ? 4'b1110 : 4'b1111;
															assign node29020 = (inp[10]) ? 4'b1111 : 4'b1110;
														assign node29023 = (inp[9]) ? node29031 : node29024;
															assign node29024 = (inp[10]) ? node29028 : node29025;
																assign node29025 = (inp[11]) ? 4'b1111 : 4'b1110;
																assign node29028 = (inp[11]) ? 4'b1110 : 4'b1111;
															assign node29031 = (inp[10]) ? node29033 : 4'b1110;
																assign node29033 = (inp[11]) ? 4'b1111 : 4'b1110;
													assign node29036 = (inp[9]) ? node29048 : node29037;
														assign node29037 = (inp[10]) ? node29043 : node29038;
															assign node29038 = (inp[0]) ? 4'b1001 : node29039;
																assign node29039 = (inp[11]) ? 4'b1000 : 4'b1001;
															assign node29043 = (inp[0]) ? 4'b1000 : node29044;
																assign node29044 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node29048 = (inp[10]) ? node29054 : node29049;
															assign node29049 = (inp[11]) ? node29051 : 4'b1000;
																assign node29051 = (inp[0]) ? 4'b1000 : 4'b1001;
															assign node29054 = (inp[0]) ? 4'b1001 : node29055;
																assign node29055 = (inp[11]) ? 4'b1000 : 4'b1001;
								assign node29059 = (inp[2]) ? node29413 : node29060;
									assign node29060 = (inp[1]) ? node29236 : node29061;
										assign node29061 = (inp[5]) ? node29143 : node29062;
											assign node29062 = (inp[15]) ? node29104 : node29063;
												assign node29063 = (inp[7]) ? node29083 : node29064;
													assign node29064 = (inp[10]) ? node29072 : node29065;
														assign node29065 = (inp[0]) ? 4'b1101 : node29066;
															assign node29066 = (inp[9]) ? node29068 : 4'b1101;
																assign node29068 = (inp[11]) ? 4'b1100 : 4'b1101;
														assign node29072 = (inp[9]) ? node29078 : node29073;
															assign node29073 = (inp[0]) ? 4'b1101 : node29074;
																assign node29074 = (inp[11]) ? 4'b1100 : 4'b1101;
															assign node29078 = (inp[0]) ? 4'b1100 : node29079;
																assign node29079 = (inp[11]) ? 4'b1101 : 4'b1100;
													assign node29083 = (inp[10]) ? node29093 : node29084;
														assign node29084 = (inp[0]) ? 4'b1111 : node29085;
															assign node29085 = (inp[9]) ? node29089 : node29086;
																assign node29086 = (inp[11]) ? 4'b1111 : 4'b1110;
																assign node29089 = (inp[11]) ? 4'b1110 : 4'b1111;
														assign node29093 = (inp[9]) ? node29099 : node29094;
															assign node29094 = (inp[0]) ? 4'b1111 : node29095;
																assign node29095 = (inp[11]) ? 4'b1110 : 4'b1111;
															assign node29099 = (inp[0]) ? 4'b1110 : node29100;
																assign node29100 = (inp[11]) ? 4'b1111 : 4'b1110;
												assign node29104 = (inp[7]) ? node29124 : node29105;
													assign node29105 = (inp[0]) ? node29119 : node29106;
														assign node29106 = (inp[10]) ? node29112 : node29107;
															assign node29107 = (inp[11]) ? node29109 : 4'b1110;
																assign node29109 = (inp[9]) ? 4'b1111 : 4'b1110;
															assign node29112 = (inp[11]) ? node29116 : node29113;
																assign node29113 = (inp[9]) ? 4'b1111 : 4'b1110;
																assign node29116 = (inp[9]) ? 4'b1110 : 4'b1111;
														assign node29119 = (inp[10]) ? node29121 : 4'b1110;
															assign node29121 = (inp[9]) ? 4'b1111 : 4'b1110;
													assign node29124 = (inp[10]) ? node29136 : node29125;
														assign node29125 = (inp[9]) ? node29131 : node29126;
															assign node29126 = (inp[11]) ? 4'b1001 : node29127;
																assign node29127 = (inp[0]) ? 4'b1000 : 4'b1001;
															assign node29131 = (inp[0]) ? node29133 : 4'b1000;
																assign node29133 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node29136 = (inp[9]) ? node29138 : 4'b1000;
															assign node29138 = (inp[11]) ? 4'b1001 : node29139;
																assign node29139 = (inp[0]) ? 4'b1000 : 4'b1001;
											assign node29143 = (inp[11]) ? node29201 : node29144;
												assign node29144 = (inp[15]) ? node29174 : node29145;
													assign node29145 = (inp[7]) ? node29159 : node29146;
														assign node29146 = (inp[10]) ? node29154 : node29147;
															assign node29147 = (inp[9]) ? node29151 : node29148;
																assign node29148 = (inp[0]) ? 4'b1001 : 4'b1000;
																assign node29151 = (inp[0]) ? 4'b1000 : 4'b1001;
															assign node29154 = (inp[0]) ? 4'b1001 : node29155;
																assign node29155 = (inp[9]) ? 4'b1000 : 4'b1001;
														assign node29159 = (inp[0]) ? node29167 : node29160;
															assign node29160 = (inp[9]) ? node29164 : node29161;
																assign node29161 = (inp[10]) ? 4'b1010 : 4'b1011;
																assign node29164 = (inp[10]) ? 4'b1011 : 4'b1010;
															assign node29167 = (inp[10]) ? node29171 : node29168;
																assign node29168 = (inp[9]) ? 4'b1011 : 4'b1010;
																assign node29171 = (inp[9]) ? 4'b1010 : 4'b1011;
													assign node29174 = (inp[7]) ? node29188 : node29175;
														assign node29175 = (inp[9]) ? node29181 : node29176;
															assign node29176 = (inp[10]) ? 4'b1010 : node29177;
																assign node29177 = (inp[0]) ? 4'b1010 : 4'b1011;
															assign node29181 = (inp[0]) ? node29185 : node29182;
																assign node29182 = (inp[10]) ? 4'b1011 : 4'b1010;
																assign node29185 = (inp[10]) ? 4'b1010 : 4'b1011;
														assign node29188 = (inp[0]) ? node29196 : node29189;
															assign node29189 = (inp[10]) ? node29193 : node29190;
																assign node29190 = (inp[9]) ? 4'b1000 : 4'b1001;
																assign node29193 = (inp[9]) ? 4'b1001 : 4'b1000;
															assign node29196 = (inp[9]) ? 4'b1000 : node29197;
																assign node29197 = (inp[10]) ? 4'b1000 : 4'b1001;
												assign node29201 = (inp[9]) ? node29219 : node29202;
													assign node29202 = (inp[7]) ? node29210 : node29203;
														assign node29203 = (inp[15]) ? node29207 : node29204;
															assign node29204 = (inp[10]) ? 4'b1001 : 4'b1000;
															assign node29207 = (inp[10]) ? 4'b1010 : 4'b1011;
														assign node29210 = (inp[15]) ? node29214 : node29211;
															assign node29211 = (inp[10]) ? 4'b1010 : 4'b1011;
															assign node29214 = (inp[10]) ? node29216 : 4'b1001;
																assign node29216 = (inp[0]) ? 4'b1000 : 4'b1001;
													assign node29219 = (inp[10]) ? node29227 : node29220;
														assign node29220 = (inp[7]) ? node29224 : node29221;
															assign node29221 = (inp[15]) ? 4'b1010 : 4'b1001;
															assign node29224 = (inp[15]) ? 4'b1001 : 4'b1010;
														assign node29227 = (inp[15]) ? node29231 : node29228;
															assign node29228 = (inp[7]) ? 4'b1011 : 4'b1000;
															assign node29231 = (inp[7]) ? node29233 : 4'b1011;
																assign node29233 = (inp[0]) ? 4'b1001 : 4'b1000;
										assign node29236 = (inp[7]) ? node29328 : node29237;
											assign node29237 = (inp[15]) ? node29283 : node29238;
												assign node29238 = (inp[5]) ? node29262 : node29239;
													assign node29239 = (inp[11]) ? node29247 : node29240;
														assign node29240 = (inp[10]) ? node29244 : node29241;
															assign node29241 = (inp[9]) ? 4'b1101 : 4'b1100;
															assign node29244 = (inp[9]) ? 4'b1100 : 4'b1101;
														assign node29247 = (inp[0]) ? node29255 : node29248;
															assign node29248 = (inp[10]) ? node29252 : node29249;
																assign node29249 = (inp[9]) ? 4'b1100 : 4'b1101;
																assign node29252 = (inp[9]) ? 4'b1101 : 4'b1100;
															assign node29255 = (inp[9]) ? node29259 : node29256;
																assign node29256 = (inp[10]) ? 4'b1101 : 4'b1100;
																assign node29259 = (inp[10]) ? 4'b1100 : 4'b1101;
													assign node29262 = (inp[0]) ? node29270 : node29263;
														assign node29263 = (inp[9]) ? node29267 : node29264;
															assign node29264 = (inp[10]) ? 4'b1101 : 4'b1100;
															assign node29267 = (inp[10]) ? 4'b1100 : 4'b1101;
														assign node29270 = (inp[9]) ? node29276 : node29271;
															assign node29271 = (inp[11]) ? node29273 : 4'b1100;
																assign node29273 = (inp[10]) ? 4'b1101 : 4'b1100;
															assign node29276 = (inp[11]) ? node29280 : node29277;
																assign node29277 = (inp[10]) ? 4'b1101 : 4'b1100;
																assign node29280 = (inp[10]) ? 4'b1100 : 4'b1101;
												assign node29283 = (inp[0]) ? node29303 : node29284;
													assign node29284 = (inp[10]) ? node29294 : node29285;
														assign node29285 = (inp[9]) ? node29289 : node29286;
															assign node29286 = (inp[11]) ? 4'b1111 : 4'b1110;
															assign node29289 = (inp[11]) ? 4'b1110 : node29290;
																assign node29290 = (inp[5]) ? 4'b1111 : 4'b1110;
														assign node29294 = (inp[9]) ? node29298 : node29295;
															assign node29295 = (inp[11]) ? 4'b1110 : 4'b1111;
															assign node29298 = (inp[5]) ? node29300 : 4'b1111;
																assign node29300 = (inp[11]) ? 4'b1111 : 4'b1110;
													assign node29303 = (inp[5]) ? node29317 : node29304;
														assign node29304 = (inp[10]) ? node29312 : node29305;
															assign node29305 = (inp[11]) ? node29309 : node29306;
																assign node29306 = (inp[9]) ? 4'b1111 : 4'b1110;
																assign node29309 = (inp[9]) ? 4'b1110 : 4'b1111;
															assign node29312 = (inp[11]) ? node29314 : 4'b1111;
																assign node29314 = (inp[9]) ? 4'b1111 : 4'b1110;
														assign node29317 = (inp[11]) ? node29323 : node29318;
															assign node29318 = (inp[9]) ? 4'b1111 : node29319;
																assign node29319 = (inp[10]) ? 4'b1111 : 4'b1110;
															assign node29323 = (inp[9]) ? node29325 : 4'b1111;
																assign node29325 = (inp[10]) ? 4'b1110 : 4'b1111;
											assign node29328 = (inp[15]) ? node29372 : node29329;
												assign node29329 = (inp[9]) ? node29353 : node29330;
													assign node29330 = (inp[0]) ? node29342 : node29331;
														assign node29331 = (inp[10]) ? node29337 : node29332;
															assign node29332 = (inp[11]) ? 4'b1111 : node29333;
																assign node29333 = (inp[5]) ? 4'b1111 : 4'b1110;
															assign node29337 = (inp[11]) ? 4'b1110 : node29338;
																assign node29338 = (inp[5]) ? 4'b1110 : 4'b1111;
														assign node29342 = (inp[10]) ? node29348 : node29343;
															assign node29343 = (inp[5]) ? node29345 : 4'b1110;
																assign node29345 = (inp[11]) ? 4'b1111 : 4'b1110;
															assign node29348 = (inp[11]) ? node29350 : 4'b1111;
																assign node29350 = (inp[5]) ? 4'b1110 : 4'b1111;
													assign node29353 = (inp[5]) ? node29361 : node29354;
														assign node29354 = (inp[10]) ? node29356 : 4'b1111;
															assign node29356 = (inp[11]) ? node29358 : 4'b1110;
																assign node29358 = (inp[0]) ? 4'b1110 : 4'b1111;
														assign node29361 = (inp[10]) ? node29367 : node29362;
															assign node29362 = (inp[11]) ? 4'b1110 : node29363;
																assign node29363 = (inp[0]) ? 4'b1111 : 4'b1110;
															assign node29367 = (inp[11]) ? 4'b1111 : node29368;
																assign node29368 = (inp[0]) ? 4'b1110 : 4'b1111;
												assign node29372 = (inp[5]) ? node29394 : node29373;
													assign node29373 = (inp[11]) ? node29385 : node29374;
														assign node29374 = (inp[0]) ? node29380 : node29375;
															assign node29375 = (inp[10]) ? node29377 : 4'b1100;
																assign node29377 = (inp[9]) ? 4'b1100 : 4'b1101;
															assign node29380 = (inp[10]) ? node29382 : 4'b1101;
																assign node29382 = (inp[9]) ? 4'b1100 : 4'b1101;
														assign node29385 = (inp[10]) ? 4'b1100 : node29386;
															assign node29386 = (inp[0]) ? node29390 : node29387;
																assign node29387 = (inp[9]) ? 4'b1100 : 4'b1101;
																assign node29390 = (inp[9]) ? 4'b1101 : 4'b1100;
													assign node29394 = (inp[10]) ? node29404 : node29395;
														assign node29395 = (inp[9]) ? node29401 : node29396;
															assign node29396 = (inp[11]) ? 4'b1001 : node29397;
																assign node29397 = (inp[0]) ? 4'b1000 : 4'b1001;
															assign node29401 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node29404 = (inp[9]) ? node29410 : node29405;
															assign node29405 = (inp[11]) ? 4'b1000 : node29406;
																assign node29406 = (inp[0]) ? 4'b1001 : 4'b1000;
															assign node29410 = (inp[11]) ? 4'b1001 : 4'b1000;
									assign node29413 = (inp[5]) ? node29621 : node29414;
										assign node29414 = (inp[1]) ? node29508 : node29415;
											assign node29415 = (inp[15]) ? node29471 : node29416;
												assign node29416 = (inp[7]) ? node29442 : node29417;
													assign node29417 = (inp[0]) ? node29427 : node29418;
														assign node29418 = (inp[10]) ? 4'b1000 : node29419;
															assign node29419 = (inp[9]) ? node29423 : node29420;
																assign node29420 = (inp[11]) ? 4'b1000 : 4'b1001;
																assign node29423 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node29427 = (inp[11]) ? node29435 : node29428;
															assign node29428 = (inp[10]) ? node29432 : node29429;
																assign node29429 = (inp[9]) ? 4'b1000 : 4'b1001;
																assign node29432 = (inp[9]) ? 4'b1001 : 4'b1000;
															assign node29435 = (inp[10]) ? node29439 : node29436;
																assign node29436 = (inp[9]) ? 4'b1000 : 4'b1001;
																assign node29439 = (inp[9]) ? 4'b1001 : 4'b1000;
													assign node29442 = (inp[11]) ? node29456 : node29443;
														assign node29443 = (inp[0]) ? node29449 : node29444;
															assign node29444 = (inp[10]) ? 4'b1011 : node29445;
																assign node29445 = (inp[9]) ? 4'b1010 : 4'b1011;
															assign node29449 = (inp[9]) ? node29453 : node29450;
																assign node29450 = (inp[10]) ? 4'b1010 : 4'b1011;
																assign node29453 = (inp[10]) ? 4'b1011 : 4'b1010;
														assign node29456 = (inp[10]) ? node29464 : node29457;
															assign node29457 = (inp[0]) ? node29461 : node29458;
																assign node29458 = (inp[9]) ? 4'b1011 : 4'b1010;
																assign node29461 = (inp[9]) ? 4'b1010 : 4'b1011;
															assign node29464 = (inp[0]) ? node29468 : node29465;
																assign node29465 = (inp[9]) ? 4'b1010 : 4'b1011;
																assign node29468 = (inp[9]) ? 4'b1011 : 4'b1010;
												assign node29471 = (inp[7]) ? node29493 : node29472;
													assign node29472 = (inp[10]) ? node29482 : node29473;
														assign node29473 = (inp[9]) ? node29479 : node29474;
															assign node29474 = (inp[11]) ? node29476 : 4'b1010;
																assign node29476 = (inp[0]) ? 4'b1010 : 4'b1011;
															assign node29479 = (inp[11]) ? 4'b1010 : 4'b1011;
														assign node29482 = (inp[9]) ? node29488 : node29483;
															assign node29483 = (inp[0]) ? 4'b1011 : node29484;
																assign node29484 = (inp[11]) ? 4'b1010 : 4'b1011;
															assign node29488 = (inp[0]) ? 4'b1010 : node29489;
																assign node29489 = (inp[11]) ? 4'b1011 : 4'b1010;
													assign node29493 = (inp[9]) ? node29501 : node29494;
														assign node29494 = (inp[10]) ? node29496 : 4'b1100;
															assign node29496 = (inp[0]) ? 4'b1101 : node29497;
																assign node29497 = (inp[11]) ? 4'b1100 : 4'b1101;
														assign node29501 = (inp[10]) ? 4'b1100 : node29502;
															assign node29502 = (inp[0]) ? 4'b1101 : node29503;
																assign node29503 = (inp[11]) ? 4'b1100 : 4'b1101;
											assign node29508 = (inp[0]) ? node29570 : node29509;
												assign node29509 = (inp[15]) ? node29541 : node29510;
													assign node29510 = (inp[7]) ? node29526 : node29511;
														assign node29511 = (inp[11]) ? node29519 : node29512;
															assign node29512 = (inp[9]) ? node29516 : node29513;
																assign node29513 = (inp[10]) ? 4'b1000 : 4'b1001;
																assign node29516 = (inp[10]) ? 4'b1001 : 4'b1000;
															assign node29519 = (inp[9]) ? node29523 : node29520;
																assign node29520 = (inp[10]) ? 4'b1001 : 4'b1000;
																assign node29523 = (inp[10]) ? 4'b1000 : 4'b1001;
														assign node29526 = (inp[10]) ? node29534 : node29527;
															assign node29527 = (inp[9]) ? node29531 : node29528;
																assign node29528 = (inp[11]) ? 4'b1010 : 4'b1011;
																assign node29531 = (inp[11]) ? 4'b1011 : 4'b1010;
															assign node29534 = (inp[11]) ? node29538 : node29535;
																assign node29535 = (inp[9]) ? 4'b1011 : 4'b1010;
																assign node29538 = (inp[9]) ? 4'b1010 : 4'b1011;
													assign node29541 = (inp[7]) ? node29557 : node29542;
														assign node29542 = (inp[11]) ? node29550 : node29543;
															assign node29543 = (inp[9]) ? node29547 : node29544;
																assign node29544 = (inp[10]) ? 4'b1011 : 4'b1010;
																assign node29547 = (inp[10]) ? 4'b1010 : 4'b1011;
															assign node29550 = (inp[10]) ? node29554 : node29551;
																assign node29551 = (inp[9]) ? 4'b1011 : 4'b1010;
																assign node29554 = (inp[9]) ? 4'b1010 : 4'b1011;
														assign node29557 = (inp[10]) ? node29565 : node29558;
															assign node29558 = (inp[9]) ? node29562 : node29559;
																assign node29559 = (inp[11]) ? 4'b1000 : 4'b1001;
																assign node29562 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node29565 = (inp[11]) ? 4'b1000 : node29566;
																assign node29566 = (inp[9]) ? 4'b1001 : 4'b1000;
												assign node29570 = (inp[11]) ? node29594 : node29571;
													assign node29571 = (inp[7]) ? node29581 : node29572;
														assign node29572 = (inp[15]) ? node29574 : 4'b1001;
															assign node29574 = (inp[9]) ? node29578 : node29575;
																assign node29575 = (inp[10]) ? 4'b1010 : 4'b1011;
																assign node29578 = (inp[10]) ? 4'b1011 : 4'b1010;
														assign node29581 = (inp[15]) ? node29589 : node29582;
															assign node29582 = (inp[10]) ? node29586 : node29583;
																assign node29583 = (inp[9]) ? 4'b1010 : 4'b1011;
																assign node29586 = (inp[9]) ? 4'b1011 : 4'b1010;
															assign node29589 = (inp[10]) ? node29591 : 4'b1001;
																assign node29591 = (inp[9]) ? 4'b1001 : 4'b1000;
													assign node29594 = (inp[7]) ? node29608 : node29595;
														assign node29595 = (inp[15]) ? node29603 : node29596;
															assign node29596 = (inp[9]) ? node29600 : node29597;
																assign node29597 = (inp[10]) ? 4'b1000 : 4'b1001;
																assign node29600 = (inp[10]) ? 4'b1001 : 4'b1000;
															assign node29603 = (inp[9]) ? 4'b1011 : node29604;
																assign node29604 = (inp[10]) ? 4'b1011 : 4'b1010;
														assign node29608 = (inp[15]) ? node29616 : node29609;
															assign node29609 = (inp[10]) ? node29613 : node29610;
																assign node29610 = (inp[9]) ? 4'b1010 : 4'b1011;
																assign node29613 = (inp[9]) ? 4'b1011 : 4'b1010;
															assign node29616 = (inp[9]) ? 4'b1000 : node29617;
																assign node29617 = (inp[10]) ? 4'b1000 : 4'b1001;
										assign node29621 = (inp[1]) ? node29697 : node29622;
											assign node29622 = (inp[7]) ? node29660 : node29623;
												assign node29623 = (inp[15]) ? node29643 : node29624;
													assign node29624 = (inp[0]) ? node29636 : node29625;
														assign node29625 = (inp[11]) ? node29631 : node29626;
															assign node29626 = (inp[10]) ? node29628 : 4'b1101;
																assign node29628 = (inp[9]) ? 4'b1101 : 4'b1100;
															assign node29631 = (inp[9]) ? node29633 : 4'b1100;
																assign node29633 = (inp[10]) ? 4'b1100 : 4'b1101;
														assign node29636 = (inp[9]) ? node29640 : node29637;
															assign node29637 = (inp[10]) ? 4'b1100 : 4'b1101;
															assign node29640 = (inp[10]) ? 4'b1101 : 4'b1100;
													assign node29643 = (inp[10]) ? node29651 : node29644;
														assign node29644 = (inp[9]) ? 4'b1111 : node29645;
															assign node29645 = (inp[11]) ? node29647 : 4'b1110;
																assign node29647 = (inp[0]) ? 4'b1110 : 4'b1111;
														assign node29651 = (inp[9]) ? node29655 : node29652;
															assign node29652 = (inp[11]) ? 4'b1110 : 4'b1111;
															assign node29655 = (inp[11]) ? node29657 : 4'b1110;
																assign node29657 = (inp[0]) ? 4'b1110 : 4'b1111;
												assign node29660 = (inp[15]) ? node29682 : node29661;
													assign node29661 = (inp[11]) ? node29669 : node29662;
														assign node29662 = (inp[9]) ? node29666 : node29663;
															assign node29663 = (inp[10]) ? 4'b1111 : 4'b1110;
															assign node29666 = (inp[10]) ? 4'b1110 : 4'b1111;
														assign node29669 = (inp[0]) ? node29675 : node29670;
															assign node29670 = (inp[9]) ? node29672 : 4'b1111;
																assign node29672 = (inp[10]) ? 4'b1111 : 4'b1110;
															assign node29675 = (inp[9]) ? node29679 : node29676;
																assign node29676 = (inp[10]) ? 4'b1111 : 4'b1110;
																assign node29679 = (inp[10]) ? 4'b1110 : 4'b1111;
													assign node29682 = (inp[9]) ? node29692 : node29683;
														assign node29683 = (inp[10]) ? node29689 : node29684;
															assign node29684 = (inp[11]) ? 4'b1101 : node29685;
																assign node29685 = (inp[0]) ? 4'b1100 : 4'b1101;
															assign node29689 = (inp[11]) ? 4'b1100 : 4'b1101;
														assign node29692 = (inp[10]) ? 4'b1101 : node29693;
															assign node29693 = (inp[11]) ? 4'b1100 : 4'b1101;
											assign node29697 = (inp[15]) ? node29741 : node29698;
												assign node29698 = (inp[7]) ? node29720 : node29699;
													assign node29699 = (inp[0]) ? node29707 : node29700;
														assign node29700 = (inp[10]) ? node29704 : node29701;
															assign node29701 = (inp[9]) ? 4'b1000 : 4'b1001;
															assign node29704 = (inp[9]) ? 4'b1001 : 4'b1000;
														assign node29707 = (inp[9]) ? node29715 : node29708;
															assign node29708 = (inp[10]) ? node29712 : node29709;
																assign node29709 = (inp[11]) ? 4'b1001 : 4'b1000;
																assign node29712 = (inp[11]) ? 4'b1000 : 4'b1001;
															assign node29715 = (inp[11]) ? 4'b1000 : node29716;
																assign node29716 = (inp[10]) ? 4'b1000 : 4'b1001;
													assign node29720 = (inp[11]) ? node29734 : node29721;
														assign node29721 = (inp[9]) ? node29729 : node29722;
															assign node29722 = (inp[0]) ? node29726 : node29723;
																assign node29723 = (inp[10]) ? 4'b1011 : 4'b1010;
																assign node29726 = (inp[10]) ? 4'b1010 : 4'b1011;
															assign node29729 = (inp[10]) ? 4'b1011 : node29730;
																assign node29730 = (inp[0]) ? 4'b1010 : 4'b1011;
														assign node29734 = (inp[9]) ? node29738 : node29735;
															assign node29735 = (inp[10]) ? 4'b1011 : 4'b1010;
															assign node29738 = (inp[10]) ? 4'b1010 : 4'b1011;
												assign node29741 = (inp[7]) ? node29759 : node29742;
													assign node29742 = (inp[9]) ? node29748 : node29743;
														assign node29743 = (inp[10]) ? node29745 : 4'b1011;
															assign node29745 = (inp[0]) ? 4'b1010 : 4'b1011;
														assign node29748 = (inp[10]) ? node29754 : node29749;
															assign node29749 = (inp[0]) ? 4'b1010 : node29750;
																assign node29750 = (inp[11]) ? 4'b1011 : 4'b1010;
															assign node29754 = (inp[0]) ? 4'b1011 : node29755;
																assign node29755 = (inp[11]) ? 4'b1010 : 4'b1011;
													assign node29759 = (inp[10]) ? node29771 : node29760;
														assign node29760 = (inp[9]) ? node29766 : node29761;
															assign node29761 = (inp[0]) ? 4'b1100 : node29762;
																assign node29762 = (inp[11]) ? 4'b1101 : 4'b1100;
															assign node29766 = (inp[11]) ? node29768 : 4'b1101;
																assign node29768 = (inp[0]) ? 4'b1101 : 4'b1100;
														assign node29771 = (inp[9]) ? 4'b1100 : node29772;
															assign node29772 = (inp[11]) ? 4'b1100 : 4'b1101;
							assign node29776 = (inp[10]) ? node30140 : node29777;
								assign node29777 = (inp[0]) ? node29965 : node29778;
									assign node29778 = (inp[2]) ? node29866 : node29779;
										assign node29779 = (inp[1]) ? node29821 : node29780;
											assign node29780 = (inp[5]) ? node29798 : node29781;
												assign node29781 = (inp[11]) ? node29789 : node29782;
													assign node29782 = (inp[13]) ? node29784 : 4'b1000;
														assign node29784 = (inp[7]) ? 4'b1000 : node29785;
															assign node29785 = (inp[15]) ? 4'b1001 : 4'b1000;
													assign node29789 = (inp[7]) ? node29791 : 4'b1001;
														assign node29791 = (inp[15]) ? node29795 : node29792;
															assign node29792 = (inp[13]) ? 4'b1000 : 4'b1001;
															assign node29795 = (inp[13]) ? 4'b1001 : 4'b1000;
												assign node29798 = (inp[7]) ? node29810 : node29799;
													assign node29799 = (inp[15]) ? node29805 : node29800;
														assign node29800 = (inp[13]) ? 4'b1100 : node29801;
															assign node29801 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node29805 = (inp[13]) ? node29807 : 4'b1000;
															assign node29807 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node29810 = (inp[15]) ? node29816 : node29811;
														assign node29811 = (inp[13]) ? node29813 : 4'b1001;
															assign node29813 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node29816 = (inp[13]) ? node29818 : 4'b1101;
															assign node29818 = (inp[11]) ? 4'b1100 : 4'b1101;
											assign node29821 = (inp[5]) ? node29843 : node29822;
												assign node29822 = (inp[13]) ? node29836 : node29823;
													assign node29823 = (inp[7]) ? node29829 : node29824;
														assign node29824 = (inp[15]) ? 4'b1100 : node29825;
															assign node29825 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node29829 = (inp[11]) ? node29833 : node29830;
															assign node29830 = (inp[15]) ? 4'b1101 : 4'b1100;
															assign node29833 = (inp[15]) ? 4'b1100 : 4'b1101;
													assign node29836 = (inp[15]) ? node29838 : 4'b1100;
														assign node29838 = (inp[7]) ? 4'b1100 : node29839;
															assign node29839 = (inp[11]) ? 4'b1101 : 4'b1100;
												assign node29843 = (inp[7]) ? node29855 : node29844;
													assign node29844 = (inp[15]) ? node29850 : node29845;
														assign node29845 = (inp[11]) ? 4'b1000 : node29846;
															assign node29846 = (inp[13]) ? 4'b1001 : 4'b1000;
														assign node29850 = (inp[11]) ? 4'b1100 : node29851;
															assign node29851 = (inp[13]) ? 4'b1100 : 4'b1101;
													assign node29855 = (inp[15]) ? node29861 : node29856;
														assign node29856 = (inp[13]) ? node29858 : 4'b1101;
															assign node29858 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node29861 = (inp[13]) ? node29863 : 4'b1000;
															assign node29863 = (inp[11]) ? 4'b1001 : 4'b1000;
										assign node29866 = (inp[1]) ? node29920 : node29867;
											assign node29867 = (inp[5]) ? node29897 : node29868;
												assign node29868 = (inp[13]) ? node29876 : node29869;
													assign node29869 = (inp[11]) ? 4'b1100 : node29870;
														assign node29870 = (inp[7]) ? node29872 : 4'b1100;
															assign node29872 = (inp[15]) ? 4'b1101 : 4'b1100;
													assign node29876 = (inp[7]) ? node29892 : node29877;
														assign node29877 = (inp[9]) ? node29885 : node29878;
															assign node29878 = (inp[11]) ? node29882 : node29879;
																assign node29879 = (inp[15]) ? 4'b1100 : 4'b1101;
																assign node29882 = (inp[15]) ? 4'b1101 : 4'b1100;
															assign node29885 = (inp[11]) ? node29889 : node29886;
																assign node29886 = (inp[15]) ? 4'b1100 : 4'b1101;
																assign node29889 = (inp[15]) ? 4'b1101 : 4'b1100;
														assign node29892 = (inp[15]) ? 4'b1100 : node29893;
															assign node29893 = (inp[11]) ? 4'b1100 : 4'b1101;
												assign node29897 = (inp[7]) ? node29909 : node29898;
													assign node29898 = (inp[15]) ? node29904 : node29899;
														assign node29899 = (inp[11]) ? node29901 : 4'b1001;
															assign node29901 = (inp[13]) ? 4'b1001 : 4'b1000;
														assign node29904 = (inp[13]) ? 4'b1100 : node29905;
															assign node29905 = (inp[11]) ? 4'b1100 : 4'b1101;
													assign node29909 = (inp[15]) ? node29915 : node29910;
														assign node29910 = (inp[11]) ? node29912 : 4'b1100;
															assign node29912 = (inp[13]) ? 4'b1100 : 4'b1101;
														assign node29915 = (inp[13]) ? node29917 : 4'b1000;
															assign node29917 = (inp[11]) ? 4'b1001 : 4'b1000;
											assign node29920 = (inp[5]) ? node29942 : node29921;
												assign node29921 = (inp[11]) ? node29929 : node29922;
													assign node29922 = (inp[7]) ? node29924 : 4'b1001;
														assign node29924 = (inp[13]) ? 4'b1001 : node29925;
															assign node29925 = (inp[15]) ? 4'b1000 : 4'b1001;
													assign node29929 = (inp[7]) ? node29937 : node29930;
														assign node29930 = (inp[13]) ? node29934 : node29931;
															assign node29931 = (inp[15]) ? 4'b1001 : 4'b1000;
															assign node29934 = (inp[15]) ? 4'b1000 : 4'b1001;
														assign node29937 = (inp[15]) ? 4'b1001 : node29938;
															assign node29938 = (inp[13]) ? 4'b1001 : 4'b1000;
												assign node29942 = (inp[7]) ? node29954 : node29943;
													assign node29943 = (inp[15]) ? node29949 : node29944;
														assign node29944 = (inp[13]) ? 4'b1101 : node29945;
															assign node29945 = (inp[11]) ? 4'b1100 : 4'b1101;
														assign node29949 = (inp[11]) ? 4'b1001 : node29950;
															assign node29950 = (inp[13]) ? 4'b1001 : 4'b1000;
													assign node29954 = (inp[15]) ? node29960 : node29955;
														assign node29955 = (inp[13]) ? node29957 : 4'b1000;
															assign node29957 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node29960 = (inp[11]) ? 4'b1100 : node29961;
															assign node29961 = (inp[13]) ? 4'b1100 : 4'b1101;
									assign node29965 = (inp[1]) ? node30047 : node29966;
										assign node29966 = (inp[2]) ? node30006 : node29967;
											assign node29967 = (inp[5]) ? node29983 : node29968;
												assign node29968 = (inp[11]) ? node29974 : node29969;
													assign node29969 = (inp[15]) ? node29971 : 4'b1001;
														assign node29971 = (inp[7]) ? 4'b1001 : 4'b1000;
													assign node29974 = (inp[13]) ? node29980 : node29975;
														assign node29975 = (inp[15]) ? node29977 : 4'b1000;
															assign node29977 = (inp[7]) ? 4'b1001 : 4'b1000;
														assign node29980 = (inp[15]) ? 4'b1000 : 4'b1001;
												assign node29983 = (inp[7]) ? node29995 : node29984;
													assign node29984 = (inp[15]) ? node29990 : node29985;
														assign node29985 = (inp[13]) ? 4'b1101 : node29986;
															assign node29986 = (inp[11]) ? 4'b1100 : 4'b1101;
														assign node29990 = (inp[11]) ? node29992 : 4'b1001;
															assign node29992 = (inp[13]) ? 4'b1000 : 4'b1001;
													assign node29995 = (inp[15]) ? node30001 : node29996;
														assign node29996 = (inp[11]) ? 4'b1000 : node29997;
															assign node29997 = (inp[13]) ? 4'b1001 : 4'b1000;
														assign node30001 = (inp[11]) ? node30003 : 4'b1100;
															assign node30003 = (inp[13]) ? 4'b1101 : 4'b1100;
											assign node30006 = (inp[5]) ? node30024 : node30007;
												assign node30007 = (inp[13]) ? node30015 : node30008;
													assign node30008 = (inp[15]) ? node30010 : 4'b1101;
														assign node30010 = (inp[7]) ? node30012 : 4'b1101;
															assign node30012 = (inp[11]) ? 4'b1101 : 4'b1100;
													assign node30015 = (inp[15]) ? node30019 : node30016;
														assign node30016 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node30019 = (inp[7]) ? 4'b1101 : node30020;
															assign node30020 = (inp[11]) ? 4'b1100 : 4'b1101;
												assign node30024 = (inp[15]) ? node30036 : node30025;
													assign node30025 = (inp[7]) ? node30031 : node30026;
														assign node30026 = (inp[11]) ? node30028 : 4'b1000;
															assign node30028 = (inp[13]) ? 4'b1000 : 4'b1001;
														assign node30031 = (inp[13]) ? 4'b1101 : node30032;
															assign node30032 = (inp[11]) ? 4'b1100 : 4'b1101;
													assign node30036 = (inp[7]) ? node30042 : node30037;
														assign node30037 = (inp[11]) ? 4'b1101 : node30038;
															assign node30038 = (inp[13]) ? 4'b1101 : 4'b1100;
														assign node30042 = (inp[13]) ? node30044 : 4'b1001;
															assign node30044 = (inp[11]) ? 4'b1000 : 4'b1001;
										assign node30047 = (inp[2]) ? node30095 : node30048;
											assign node30048 = (inp[5]) ? node30076 : node30049;
												assign node30049 = (inp[11]) ? node30057 : node30050;
													assign node30050 = (inp[7]) ? node30052 : 4'b1101;
														assign node30052 = (inp[15]) ? node30054 : 4'b1101;
															assign node30054 = (inp[13]) ? 4'b1101 : 4'b1100;
													assign node30057 = (inp[7]) ? node30071 : node30058;
														assign node30058 = (inp[9]) ? node30066 : node30059;
															assign node30059 = (inp[13]) ? node30063 : node30060;
																assign node30060 = (inp[15]) ? 4'b1101 : 4'b1100;
																assign node30063 = (inp[15]) ? 4'b1100 : 4'b1101;
															assign node30066 = (inp[13]) ? node30068 : 4'b1100;
																assign node30068 = (inp[15]) ? 4'b1100 : 4'b1101;
														assign node30071 = (inp[13]) ? 4'b1101 : node30072;
															assign node30072 = (inp[15]) ? 4'b1101 : 4'b1100;
												assign node30076 = (inp[15]) ? node30084 : node30077;
													assign node30077 = (inp[7]) ? 4'b1100 : node30078;
														assign node30078 = (inp[11]) ? 4'b1001 : node30079;
															assign node30079 = (inp[13]) ? 4'b1000 : 4'b1001;
													assign node30084 = (inp[7]) ? node30090 : node30085;
														assign node30085 = (inp[13]) ? 4'b1101 : node30086;
															assign node30086 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node30090 = (inp[11]) ? node30092 : 4'b1001;
															assign node30092 = (inp[13]) ? 4'b1000 : 4'b1001;
											assign node30095 = (inp[5]) ? node30117 : node30096;
												assign node30096 = (inp[13]) ? node30110 : node30097;
													assign node30097 = (inp[7]) ? node30103 : node30098;
														assign node30098 = (inp[15]) ? 4'b1000 : node30099;
															assign node30099 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node30103 = (inp[15]) ? node30107 : node30104;
															assign node30104 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node30107 = (inp[11]) ? 4'b1000 : 4'b1001;
													assign node30110 = (inp[7]) ? 4'b1000 : node30111;
														assign node30111 = (inp[15]) ? node30113 : 4'b1000;
															assign node30113 = (inp[11]) ? 4'b1001 : 4'b1000;
												assign node30117 = (inp[7]) ? node30129 : node30118;
													assign node30118 = (inp[15]) ? node30124 : node30119;
														assign node30119 = (inp[13]) ? 4'b1100 : node30120;
															assign node30120 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node30124 = (inp[13]) ? 4'b1000 : node30125;
															assign node30125 = (inp[11]) ? 4'b1000 : 4'b1001;
													assign node30129 = (inp[15]) ? node30135 : node30130;
														assign node30130 = (inp[13]) ? node30132 : 4'b1001;
															assign node30132 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node30135 = (inp[13]) ? 4'b1101 : node30136;
															assign node30136 = (inp[11]) ? 4'b1101 : 4'b1100;
								assign node30140 = (inp[0]) ? node30306 : node30141;
									assign node30141 = (inp[2]) ? node30223 : node30142;
										assign node30142 = (inp[1]) ? node30180 : node30143;
											assign node30143 = (inp[5]) ? node30161 : node30144;
												assign node30144 = (inp[11]) ? node30152 : node30145;
													assign node30145 = (inp[7]) ? 4'b1001 : node30146;
														assign node30146 = (inp[15]) ? node30148 : 4'b1001;
															assign node30148 = (inp[13]) ? 4'b1000 : 4'b1001;
													assign node30152 = (inp[13]) ? node30158 : node30153;
														assign node30153 = (inp[15]) ? node30155 : 4'b1000;
															assign node30155 = (inp[7]) ? 4'b1001 : 4'b1000;
														assign node30158 = (inp[15]) ? 4'b1000 : 4'b1001;
												assign node30161 = (inp[7]) ? node30173 : node30162;
													assign node30162 = (inp[15]) ? node30168 : node30163;
														assign node30163 = (inp[11]) ? node30165 : 4'b1101;
															assign node30165 = (inp[13]) ? 4'b1101 : 4'b1100;
														assign node30168 = (inp[13]) ? node30170 : 4'b1001;
															assign node30170 = (inp[11]) ? 4'b1000 : 4'b1001;
													assign node30173 = (inp[15]) ? node30175 : 4'b1000;
														assign node30175 = (inp[13]) ? node30177 : 4'b1100;
															assign node30177 = (inp[11]) ? 4'b1101 : 4'b1100;
											assign node30180 = (inp[5]) ? node30202 : node30181;
												assign node30181 = (inp[13]) ? node30195 : node30182;
													assign node30182 = (inp[7]) ? node30188 : node30183;
														assign node30183 = (inp[15]) ? 4'b1101 : node30184;
															assign node30184 = (inp[9]) ? 4'b1100 : 4'b1101;
														assign node30188 = (inp[15]) ? node30192 : node30189;
															assign node30189 = (inp[11]) ? 4'b1100 : 4'b1101;
															assign node30192 = (inp[11]) ? 4'b1101 : 4'b1100;
													assign node30195 = (inp[15]) ? node30197 : 4'b1101;
														assign node30197 = (inp[7]) ? 4'b1101 : node30198;
															assign node30198 = (inp[11]) ? 4'b1100 : 4'b1101;
												assign node30202 = (inp[15]) ? node30212 : node30203;
													assign node30203 = (inp[7]) ? node30207 : node30204;
														assign node30204 = (inp[13]) ? 4'b1000 : 4'b1001;
														assign node30207 = (inp[11]) ? 4'b1100 : node30208;
															assign node30208 = (inp[13]) ? 4'b1101 : 4'b1100;
													assign node30212 = (inp[7]) ? node30218 : node30213;
														assign node30213 = (inp[11]) ? 4'b1101 : node30214;
															assign node30214 = (inp[13]) ? 4'b1101 : 4'b1100;
														assign node30218 = (inp[13]) ? node30220 : 4'b1001;
															assign node30220 = (inp[11]) ? 4'b1000 : 4'b1001;
										assign node30223 = (inp[1]) ? node30265 : node30224;
											assign node30224 = (inp[5]) ? node30242 : node30225;
												assign node30225 = (inp[13]) ? node30233 : node30226;
													assign node30226 = (inp[15]) ? node30228 : 4'b1101;
														assign node30228 = (inp[11]) ? 4'b1101 : node30229;
															assign node30229 = (inp[7]) ? 4'b1100 : 4'b1101;
													assign node30233 = (inp[15]) ? node30237 : node30234;
														assign node30234 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node30237 = (inp[11]) ? node30239 : 4'b1101;
															assign node30239 = (inp[7]) ? 4'b1101 : 4'b1100;
												assign node30242 = (inp[7]) ? node30254 : node30243;
													assign node30243 = (inp[15]) ? node30249 : node30244;
														assign node30244 = (inp[11]) ? node30246 : 4'b1000;
															assign node30246 = (inp[13]) ? 4'b1000 : 4'b1001;
														assign node30249 = (inp[13]) ? 4'b1101 : node30250;
															assign node30250 = (inp[11]) ? 4'b1101 : 4'b1100;
													assign node30254 = (inp[15]) ? node30260 : node30255;
														assign node30255 = (inp[11]) ? node30257 : 4'b1101;
															assign node30257 = (inp[13]) ? 4'b1101 : 4'b1100;
														assign node30260 = (inp[11]) ? node30262 : 4'b1001;
															assign node30262 = (inp[13]) ? 4'b1000 : 4'b1001;
											assign node30265 = (inp[5]) ? node30283 : node30266;
												assign node30266 = (inp[11]) ? node30274 : node30267;
													assign node30267 = (inp[7]) ? node30269 : 4'b1000;
														assign node30269 = (inp[15]) ? node30271 : 4'b1000;
															assign node30271 = (inp[13]) ? 4'b1000 : 4'b1001;
													assign node30274 = (inp[13]) ? node30278 : node30275;
														assign node30275 = (inp[15]) ? 4'b1000 : 4'b1001;
														assign node30278 = (inp[15]) ? node30280 : 4'b1000;
															assign node30280 = (inp[9]) ? 4'b1000 : 4'b1001;
												assign node30283 = (inp[7]) ? node30295 : node30284;
													assign node30284 = (inp[15]) ? node30290 : node30285;
														assign node30285 = (inp[13]) ? 4'b1100 : node30286;
															assign node30286 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node30290 = (inp[13]) ? 4'b1000 : node30291;
															assign node30291 = (inp[11]) ? 4'b1000 : 4'b1001;
													assign node30295 = (inp[15]) ? node30301 : node30296;
														assign node30296 = (inp[11]) ? 4'b1001 : node30297;
															assign node30297 = (inp[13]) ? 4'b1000 : 4'b1001;
														assign node30301 = (inp[11]) ? 4'b1101 : node30302;
															assign node30302 = (inp[13]) ? 4'b1101 : 4'b1100;
									assign node30306 = (inp[1]) ? node30392 : node30307;
										assign node30307 = (inp[2]) ? node30349 : node30308;
											assign node30308 = (inp[5]) ? node30326 : node30309;
												assign node30309 = (inp[11]) ? node30317 : node30310;
													assign node30310 = (inp[15]) ? node30312 : 4'b1000;
														assign node30312 = (inp[13]) ? node30314 : 4'b1000;
															assign node30314 = (inp[7]) ? 4'b1000 : 4'b1001;
													assign node30317 = (inp[13]) ? node30323 : node30318;
														assign node30318 = (inp[15]) ? node30320 : 4'b1001;
															assign node30320 = (inp[7]) ? 4'b1000 : 4'b1001;
														assign node30323 = (inp[15]) ? 4'b1001 : 4'b1000;
												assign node30326 = (inp[7]) ? node30338 : node30327;
													assign node30327 = (inp[15]) ? node30333 : node30328;
														assign node30328 = (inp[11]) ? node30330 : 4'b1100;
															assign node30330 = (inp[13]) ? 4'b1100 : 4'b1101;
														assign node30333 = (inp[13]) ? node30335 : 4'b1000;
															assign node30335 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node30338 = (inp[15]) ? node30344 : node30339;
														assign node30339 = (inp[11]) ? 4'b1001 : node30340;
															assign node30340 = (inp[13]) ? 4'b1000 : 4'b1001;
														assign node30344 = (inp[11]) ? node30346 : 4'b1101;
															assign node30346 = (inp[13]) ? 4'b1100 : 4'b1101;
											assign node30349 = (inp[5]) ? node30371 : node30350;
												assign node30350 = (inp[11]) ? node30364 : node30351;
													assign node30351 = (inp[7]) ? node30357 : node30352;
														assign node30352 = (inp[15]) ? 4'b1100 : node30353;
															assign node30353 = (inp[13]) ? 4'b1101 : 4'b1100;
														assign node30357 = (inp[15]) ? node30361 : node30358;
															assign node30358 = (inp[13]) ? 4'b1101 : 4'b1100;
															assign node30361 = (inp[13]) ? 4'b1100 : 4'b1101;
													assign node30364 = (inp[15]) ? node30366 : 4'b1100;
														assign node30366 = (inp[7]) ? 4'b1100 : node30367;
															assign node30367 = (inp[13]) ? 4'b1101 : 4'b1100;
												assign node30371 = (inp[15]) ? node30381 : node30372;
													assign node30372 = (inp[7]) ? node30378 : node30373;
														assign node30373 = (inp[11]) ? node30375 : 4'b1001;
															assign node30375 = (inp[13]) ? 4'b1001 : 4'b1000;
														assign node30378 = (inp[13]) ? 4'b1100 : 4'b1101;
													assign node30381 = (inp[7]) ? node30387 : node30382;
														assign node30382 = (inp[11]) ? 4'b1100 : node30383;
															assign node30383 = (inp[13]) ? 4'b1100 : 4'b1101;
														assign node30387 = (inp[13]) ? node30389 : 4'b1000;
															assign node30389 = (inp[11]) ? 4'b1001 : 4'b1000;
										assign node30392 = (inp[2]) ? node30434 : node30393;
											assign node30393 = (inp[5]) ? node30411 : node30394;
												assign node30394 = (inp[13]) ? node30404 : node30395;
													assign node30395 = (inp[15]) ? node30399 : node30396;
														assign node30396 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node30399 = (inp[7]) ? node30401 : 4'b1100;
															assign node30401 = (inp[11]) ? 4'b1100 : 4'b1101;
													assign node30404 = (inp[15]) ? node30406 : 4'b1100;
														assign node30406 = (inp[11]) ? node30408 : 4'b1100;
															assign node30408 = (inp[7]) ? 4'b1100 : 4'b1101;
												assign node30411 = (inp[7]) ? node30423 : node30412;
													assign node30412 = (inp[15]) ? node30418 : node30413;
														assign node30413 = (inp[11]) ? 4'b1000 : node30414;
															assign node30414 = (inp[13]) ? 4'b1001 : 4'b1000;
														assign node30418 = (inp[11]) ? 4'b1100 : node30419;
															assign node30419 = (inp[13]) ? 4'b1100 : 4'b1101;
													assign node30423 = (inp[15]) ? node30429 : node30424;
														assign node30424 = (inp[13]) ? node30426 : 4'b1101;
															assign node30426 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node30429 = (inp[11]) ? node30431 : 4'b1000;
															assign node30431 = (inp[13]) ? 4'b1001 : 4'b1000;
											assign node30434 = (inp[5]) ? node30456 : node30435;
												assign node30435 = (inp[11]) ? node30443 : node30436;
													assign node30436 = (inp[13]) ? 4'b1001 : node30437;
														assign node30437 = (inp[7]) ? node30439 : 4'b1001;
															assign node30439 = (inp[15]) ? 4'b1000 : 4'b1001;
													assign node30443 = (inp[7]) ? node30451 : node30444;
														assign node30444 = (inp[15]) ? node30448 : node30445;
															assign node30445 = (inp[13]) ? 4'b1001 : 4'b1000;
															assign node30448 = (inp[13]) ? 4'b1000 : 4'b1001;
														assign node30451 = (inp[15]) ? 4'b1001 : node30452;
															assign node30452 = (inp[13]) ? 4'b1001 : 4'b1000;
												assign node30456 = (inp[7]) ? node30468 : node30457;
													assign node30457 = (inp[15]) ? node30463 : node30458;
														assign node30458 = (inp[11]) ? node30460 : 4'b1101;
															assign node30460 = (inp[13]) ? 4'b1101 : 4'b1100;
														assign node30463 = (inp[13]) ? 4'b1001 : node30464;
															assign node30464 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node30468 = (inp[15]) ? node30474 : node30469;
														assign node30469 = (inp[13]) ? node30471 : 4'b1000;
															assign node30471 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node30474 = (inp[13]) ? 4'b1100 : node30475;
															assign node30475 = (inp[11]) ? 4'b1100 : 4'b1101;
						assign node30479 = (inp[7]) ? node31771 : node30480;
							assign node30480 = (inp[8]) ? node31228 : node30481;
								assign node30481 = (inp[1]) ? node30849 : node30482;
									assign node30482 = (inp[9]) ? node30660 : node30483;
										assign node30483 = (inp[10]) ? node30581 : node30484;
											assign node30484 = (inp[0]) ? node30534 : node30485;
												assign node30485 = (inp[5]) ? node30511 : node30486;
													assign node30486 = (inp[11]) ? node30496 : node30487;
														assign node30487 = (inp[2]) ? 4'b1101 : node30488;
															assign node30488 = (inp[15]) ? node30492 : node30489;
																assign node30489 = (inp[13]) ? 4'b1100 : 4'b1000;
																assign node30492 = (inp[13]) ? 4'b1001 : 4'b1100;
														assign node30496 = (inp[13]) ? node30504 : node30497;
															assign node30497 = (inp[2]) ? node30501 : node30498;
																assign node30498 = (inp[15]) ? 4'b1101 : 4'b1001;
																assign node30501 = (inp[15]) ? 4'b1001 : 4'b1101;
															assign node30504 = (inp[2]) ? node30508 : node30505;
																assign node30505 = (inp[15]) ? 4'b1001 : 4'b1101;
																assign node30508 = (inp[15]) ? 4'b1100 : 4'b1001;
													assign node30511 = (inp[15]) ? node30521 : node30512;
														assign node30512 = (inp[2]) ? node30518 : node30513;
															assign node30513 = (inp[13]) ? node30515 : 4'b1100;
																assign node30515 = (inp[11]) ? 4'b1000 : 4'b1001;
															assign node30518 = (inp[13]) ? 4'b1100 : 4'b1000;
														assign node30521 = (inp[11]) ? node30529 : node30522;
															assign node30522 = (inp[13]) ? node30526 : node30523;
																assign node30523 = (inp[2]) ? 4'b1100 : 4'b1001;
																assign node30526 = (inp[2]) ? 4'b1000 : 4'b1100;
															assign node30529 = (inp[13]) ? node30531 : 4'b1100;
																assign node30531 = (inp[2]) ? 4'b1001 : 4'b1101;
												assign node30534 = (inp[5]) ? node30556 : node30535;
													assign node30535 = (inp[15]) ? node30547 : node30536;
														assign node30536 = (inp[11]) ? node30542 : node30537;
															assign node30537 = (inp[2]) ? node30539 : 4'b1100;
																assign node30539 = (inp[13]) ? 4'b1000 : 4'b1100;
															assign node30542 = (inp[2]) ? 4'b1000 : node30543;
																assign node30543 = (inp[13]) ? 4'b1100 : 4'b1000;
														assign node30547 = (inp[13]) ? node30551 : node30548;
															assign node30548 = (inp[2]) ? 4'b1000 : 4'b1100;
															assign node30551 = (inp[2]) ? 4'b1101 : node30552;
																assign node30552 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node30556 = (inp[11]) ? node30572 : node30557;
														assign node30557 = (inp[15]) ? node30565 : node30558;
															assign node30558 = (inp[13]) ? node30562 : node30559;
																assign node30559 = (inp[2]) ? 4'b1001 : 4'b1101;
																assign node30562 = (inp[2]) ? 4'b1101 : 4'b1001;
															assign node30565 = (inp[13]) ? node30569 : node30566;
																assign node30566 = (inp[2]) ? 4'b1101 : 4'b1001;
																assign node30569 = (inp[2]) ? 4'b1000 : 4'b1100;
														assign node30572 = (inp[15]) ? node30574 : 4'b1100;
															assign node30574 = (inp[13]) ? node30578 : node30575;
																assign node30575 = (inp[2]) ? 4'b1100 : 4'b1001;
																assign node30578 = (inp[2]) ? 4'b1000 : 4'b1100;
											assign node30581 = (inp[15]) ? node30621 : node30582;
												assign node30582 = (inp[13]) ? node30602 : node30583;
													assign node30583 = (inp[2]) ? node30591 : node30584;
														assign node30584 = (inp[5]) ? node30586 : 4'b1001;
															assign node30586 = (inp[11]) ? 4'b1101 : node30587;
																assign node30587 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node30591 = (inp[5]) ? node30597 : node30592;
															assign node30592 = (inp[11]) ? 4'b1100 : node30593;
																assign node30593 = (inp[0]) ? 4'b1101 : 4'b1100;
															assign node30597 = (inp[11]) ? 4'b1001 : node30598;
																assign node30598 = (inp[0]) ? 4'b1000 : 4'b1001;
													assign node30602 = (inp[5]) ? node30614 : node30603;
														assign node30603 = (inp[2]) ? node30609 : node30604;
															assign node30604 = (inp[0]) ? 4'b1101 : node30605;
																assign node30605 = (inp[11]) ? 4'b1100 : 4'b1101;
															assign node30609 = (inp[11]) ? node30611 : 4'b1001;
																assign node30611 = (inp[0]) ? 4'b1001 : 4'b1000;
														assign node30614 = (inp[2]) ? node30616 : 4'b1000;
															assign node30616 = (inp[11]) ? 4'b1101 : node30617;
																assign node30617 = (inp[0]) ? 4'b1100 : 4'b1101;
												assign node30621 = (inp[13]) ? node30641 : node30622;
													assign node30622 = (inp[5]) ? node30634 : node30623;
														assign node30623 = (inp[2]) ? node30629 : node30624;
															assign node30624 = (inp[11]) ? node30626 : 4'b1101;
																assign node30626 = (inp[0]) ? 4'b1101 : 4'b1100;
															assign node30629 = (inp[11]) ? node30631 : 4'b1001;
																assign node30631 = (inp[0]) ? 4'b1001 : 4'b1000;
														assign node30634 = (inp[2]) ? node30638 : node30635;
															assign node30635 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node30638 = (inp[0]) ? 4'b1100 : 4'b1101;
													assign node30641 = (inp[5]) ? node30649 : node30642;
														assign node30642 = (inp[2]) ? 4'b1100 : node30643;
															assign node30643 = (inp[11]) ? 4'b1000 : node30644;
																assign node30644 = (inp[0]) ? 4'b1001 : 4'b1000;
														assign node30649 = (inp[2]) ? node30655 : node30650;
															assign node30650 = (inp[0]) ? 4'b1101 : node30651;
																assign node30651 = (inp[11]) ? 4'b1100 : 4'b1101;
															assign node30655 = (inp[0]) ? 4'b1001 : node30656;
																assign node30656 = (inp[11]) ? 4'b1000 : 4'b1001;
										assign node30660 = (inp[10]) ? node30750 : node30661;
											assign node30661 = (inp[2]) ? node30697 : node30662;
												assign node30662 = (inp[15]) ? node30684 : node30663;
													assign node30663 = (inp[5]) ? node30675 : node30664;
														assign node30664 = (inp[13]) ? node30670 : node30665;
															assign node30665 = (inp[11]) ? node30667 : 4'b1001;
																assign node30667 = (inp[0]) ? 4'b1001 : 4'b1000;
															assign node30670 = (inp[0]) ? 4'b1101 : node30671;
																assign node30671 = (inp[11]) ? 4'b1100 : 4'b1101;
														assign node30675 = (inp[13]) ? node30679 : node30676;
															assign node30676 = (inp[11]) ? 4'b1101 : 4'b1100;
															assign node30679 = (inp[0]) ? 4'b1000 : node30680;
																assign node30680 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node30684 = (inp[0]) ? node30688 : node30685;
														assign node30685 = (inp[11]) ? 4'b1100 : 4'b1000;
														assign node30688 = (inp[13]) ? node30692 : node30689;
															assign node30689 = (inp[5]) ? 4'b1000 : 4'b1101;
															assign node30692 = (inp[5]) ? 4'b1101 : node30693;
																assign node30693 = (inp[11]) ? 4'b1000 : 4'b1001;
												assign node30697 = (inp[5]) ? node30721 : node30698;
													assign node30698 = (inp[11]) ? node30708 : node30699;
														assign node30699 = (inp[13]) ? node30705 : node30700;
															assign node30700 = (inp[15]) ? 4'b1001 : node30701;
																assign node30701 = (inp[0]) ? 4'b1101 : 4'b1100;
															assign node30705 = (inp[15]) ? 4'b1100 : 4'b1001;
														assign node30708 = (inp[15]) ? node30714 : node30709;
															assign node30709 = (inp[13]) ? node30711 : 4'b1100;
																assign node30711 = (inp[0]) ? 4'b1001 : 4'b1000;
															assign node30714 = (inp[13]) ? node30718 : node30715;
																assign node30715 = (inp[0]) ? 4'b1001 : 4'b1000;
																assign node30718 = (inp[0]) ? 4'b1100 : 4'b1101;
													assign node30721 = (inp[0]) ? node30737 : node30722;
														assign node30722 = (inp[11]) ? node30730 : node30723;
															assign node30723 = (inp[13]) ? node30727 : node30724;
																assign node30724 = (inp[15]) ? 4'b1101 : 4'b1001;
																assign node30727 = (inp[15]) ? 4'b1001 : 4'b1101;
															assign node30730 = (inp[15]) ? node30734 : node30731;
																assign node30731 = (inp[13]) ? 4'b1101 : 4'b1001;
																assign node30734 = (inp[13]) ? 4'b1000 : 4'b1101;
														assign node30737 = (inp[11]) ? node30745 : node30738;
															assign node30738 = (inp[13]) ? node30742 : node30739;
																assign node30739 = (inp[15]) ? 4'b1100 : 4'b1000;
																assign node30742 = (inp[15]) ? 4'b1001 : 4'b1100;
															assign node30745 = (inp[13]) ? node30747 : 4'b1101;
																assign node30747 = (inp[15]) ? 4'b1001 : 4'b1101;
											assign node30750 = (inp[11]) ? node30802 : node30751;
												assign node30751 = (inp[5]) ? node30779 : node30752;
													assign node30752 = (inp[2]) ? node30766 : node30753;
														assign node30753 = (inp[0]) ? node30759 : node30754;
															assign node30754 = (inp[13]) ? 4'b1100 : node30755;
																assign node30755 = (inp[15]) ? 4'b1100 : 4'b1000;
															assign node30759 = (inp[15]) ? node30763 : node30760;
																assign node30760 = (inp[13]) ? 4'b1100 : 4'b1000;
																assign node30763 = (inp[13]) ? 4'b1000 : 4'b1100;
														assign node30766 = (inp[0]) ? node30772 : node30767;
															assign node30767 = (inp[13]) ? node30769 : 4'b1101;
																assign node30769 = (inp[15]) ? 4'b1101 : 4'b1000;
															assign node30772 = (inp[13]) ? node30776 : node30773;
																assign node30773 = (inp[15]) ? 4'b1000 : 4'b1100;
																assign node30776 = (inp[15]) ? 4'b1101 : 4'b1000;
													assign node30779 = (inp[13]) ? node30793 : node30780;
														assign node30780 = (inp[0]) ? node30786 : node30781;
															assign node30781 = (inp[2]) ? 4'b1100 : node30782;
																assign node30782 = (inp[15]) ? 4'b1001 : 4'b1100;
															assign node30786 = (inp[15]) ? node30790 : node30787;
																assign node30787 = (inp[2]) ? 4'b1001 : 4'b1101;
																assign node30790 = (inp[2]) ? 4'b1101 : 4'b1001;
														assign node30793 = (inp[15]) ? node30799 : node30794;
															assign node30794 = (inp[2]) ? node30796 : 4'b1001;
																assign node30796 = (inp[0]) ? 4'b1101 : 4'b1100;
															assign node30799 = (inp[2]) ? 4'b1000 : 4'b1100;
												assign node30802 = (inp[5]) ? node30832 : node30803;
													assign node30803 = (inp[0]) ? node30817 : node30804;
														assign node30804 = (inp[15]) ? node30812 : node30805;
															assign node30805 = (inp[2]) ? node30809 : node30806;
																assign node30806 = (inp[13]) ? 4'b1101 : 4'b1001;
																assign node30809 = (inp[13]) ? 4'b1001 : 4'b1101;
															assign node30812 = (inp[2]) ? node30814 : 4'b1001;
																assign node30814 = (inp[13]) ? 4'b1100 : 4'b1001;
														assign node30817 = (inp[2]) ? node30825 : node30818;
															assign node30818 = (inp[15]) ? node30822 : node30819;
																assign node30819 = (inp[13]) ? 4'b1100 : 4'b1000;
																assign node30822 = (inp[13]) ? 4'b1001 : 4'b1100;
															assign node30825 = (inp[13]) ? node30829 : node30826;
																assign node30826 = (inp[15]) ? 4'b1000 : 4'b1101;
																assign node30829 = (inp[15]) ? 4'b1101 : 4'b1000;
													assign node30832 = (inp[15]) ? node30842 : node30833;
														assign node30833 = (inp[2]) ? node30839 : node30834;
															assign node30834 = (inp[13]) ? node30836 : 4'b1100;
																assign node30836 = (inp[0]) ? 4'b1001 : 4'b1000;
															assign node30839 = (inp[13]) ? 4'b1100 : 4'b1000;
														assign node30842 = (inp[13]) ? node30846 : node30843;
															assign node30843 = (inp[2]) ? 4'b1100 : 4'b1001;
															assign node30846 = (inp[0]) ? 4'b1100 : 4'b1001;
									assign node30849 = (inp[15]) ? node31035 : node30850;
										assign node30850 = (inp[2]) ? node30942 : node30851;
											assign node30851 = (inp[13]) ? node30899 : node30852;
												assign node30852 = (inp[5]) ? node30876 : node30853;
													assign node30853 = (inp[10]) ? node30865 : node30854;
														assign node30854 = (inp[9]) ? node30860 : node30855;
															assign node30855 = (inp[11]) ? node30857 : 4'b1000;
																assign node30857 = (inp[0]) ? 4'b1000 : 4'b1001;
															assign node30860 = (inp[0]) ? 4'b1001 : node30861;
																assign node30861 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node30865 = (inp[9]) ? node30871 : node30866;
															assign node30866 = (inp[11]) ? node30868 : 4'b1001;
																assign node30868 = (inp[0]) ? 4'b1001 : 4'b1000;
															assign node30871 = (inp[0]) ? 4'b1000 : node30872;
																assign node30872 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node30876 = (inp[9]) ? node30888 : node30877;
														assign node30877 = (inp[10]) ? node30883 : node30878;
															assign node30878 = (inp[0]) ? 4'b1001 : node30879;
																assign node30879 = (inp[11]) ? 4'b1000 : 4'b1001;
															assign node30883 = (inp[0]) ? 4'b1000 : node30884;
																assign node30884 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node30888 = (inp[10]) ? node30894 : node30889;
															assign node30889 = (inp[11]) ? node30891 : 4'b1000;
																assign node30891 = (inp[0]) ? 4'b1000 : 4'b1001;
															assign node30894 = (inp[11]) ? node30896 : 4'b1001;
																assign node30896 = (inp[0]) ? 4'b1001 : 4'b1000;
												assign node30899 = (inp[5]) ? node30921 : node30900;
													assign node30900 = (inp[11]) ? node30908 : node30901;
														assign node30901 = (inp[10]) ? node30905 : node30902;
															assign node30902 = (inp[9]) ? 4'b1101 : 4'b1100;
															assign node30905 = (inp[9]) ? 4'b1100 : 4'b1101;
														assign node30908 = (inp[10]) ? node30916 : node30909;
															assign node30909 = (inp[0]) ? node30913 : node30910;
																assign node30910 = (inp[9]) ? 4'b1100 : 4'b1101;
																assign node30913 = (inp[9]) ? 4'b1101 : 4'b1100;
															assign node30916 = (inp[9]) ? 4'b1101 : node30917;
																assign node30917 = (inp[0]) ? 4'b1101 : 4'b1100;
													assign node30921 = (inp[9]) ? node30933 : node30922;
														assign node30922 = (inp[10]) ? node30928 : node30923;
															assign node30923 = (inp[0]) ? 4'b1101 : node30924;
																assign node30924 = (inp[11]) ? 4'b1100 : 4'b1101;
															assign node30928 = (inp[0]) ? 4'b1100 : node30929;
																assign node30929 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node30933 = (inp[0]) ? 4'b1100 : node30934;
															assign node30934 = (inp[11]) ? node30938 : node30935;
																assign node30935 = (inp[10]) ? 4'b1101 : 4'b1100;
																assign node30938 = (inp[10]) ? 4'b1100 : 4'b1101;
											assign node30942 = (inp[13]) ? node30980 : node30943;
												assign node30943 = (inp[11]) ? node30965 : node30944;
													assign node30944 = (inp[0]) ? node30950 : node30945;
														assign node30945 = (inp[10]) ? 4'b1100 : node30946;
															assign node30946 = (inp[9]) ? 4'b1100 : 4'b1101;
														assign node30950 = (inp[9]) ? node30958 : node30951;
															assign node30951 = (inp[5]) ? node30955 : node30952;
																assign node30952 = (inp[10]) ? 4'b1101 : 4'b1100;
																assign node30955 = (inp[10]) ? 4'b1100 : 4'b1101;
															assign node30958 = (inp[5]) ? node30962 : node30959;
																assign node30959 = (inp[10]) ? 4'b1100 : 4'b1101;
																assign node30962 = (inp[10]) ? 4'b1101 : 4'b1100;
													assign node30965 = (inp[9]) ? node30973 : node30966;
														assign node30966 = (inp[10]) ? node30970 : node30967;
															assign node30967 = (inp[5]) ? 4'b1100 : 4'b1101;
															assign node30970 = (inp[5]) ? 4'b1101 : 4'b1100;
														assign node30973 = (inp[10]) ? node30977 : node30974;
															assign node30974 = (inp[5]) ? 4'b1101 : 4'b1100;
															assign node30977 = (inp[5]) ? 4'b1100 : 4'b1101;
												assign node30980 = (inp[10]) ? node31012 : node30981;
													assign node30981 = (inp[0]) ? node30997 : node30982;
														assign node30982 = (inp[11]) ? node30990 : node30983;
															assign node30983 = (inp[9]) ? node30987 : node30984;
																assign node30984 = (inp[5]) ? 4'b1001 : 4'b1000;
																assign node30987 = (inp[5]) ? 4'b1000 : 4'b1001;
															assign node30990 = (inp[5]) ? node30994 : node30991;
																assign node30991 = (inp[9]) ? 4'b1000 : 4'b1001;
																assign node30994 = (inp[9]) ? 4'b1001 : 4'b1000;
														assign node30997 = (inp[11]) ? node31005 : node30998;
															assign node30998 = (inp[5]) ? node31002 : node30999;
																assign node30999 = (inp[9]) ? 4'b1001 : 4'b1000;
																assign node31002 = (inp[9]) ? 4'b1000 : 4'b1001;
															assign node31005 = (inp[9]) ? node31009 : node31006;
																assign node31006 = (inp[5]) ? 4'b1001 : 4'b1000;
																assign node31009 = (inp[5]) ? 4'b1000 : 4'b1001;
													assign node31012 = (inp[5]) ? node31024 : node31013;
														assign node31013 = (inp[9]) ? node31019 : node31014;
															assign node31014 = (inp[11]) ? node31016 : 4'b1001;
																assign node31016 = (inp[0]) ? 4'b1001 : 4'b1000;
															assign node31019 = (inp[0]) ? 4'b1000 : node31020;
																assign node31020 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node31024 = (inp[9]) ? node31030 : node31025;
															assign node31025 = (inp[0]) ? 4'b1000 : node31026;
																assign node31026 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node31030 = (inp[11]) ? node31032 : 4'b1001;
																assign node31032 = (inp[0]) ? 4'b1001 : 4'b1000;
										assign node31035 = (inp[13]) ? node31133 : node31036;
											assign node31036 = (inp[2]) ? node31078 : node31037;
												assign node31037 = (inp[5]) ? node31059 : node31038;
													assign node31038 = (inp[9]) ? node31050 : node31039;
														assign node31039 = (inp[10]) ? node31045 : node31040;
															assign node31040 = (inp[0]) ? node31042 : 4'b1100;
																assign node31042 = (inp[11]) ? 4'b1100 : 4'b1101;
															assign node31045 = (inp[11]) ? 4'b1101 : node31046;
																assign node31046 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node31050 = (inp[10]) ? node31054 : node31051;
															assign node31051 = (inp[11]) ? 4'b1101 : 4'b1100;
															assign node31054 = (inp[0]) ? node31056 : 4'b1100;
																assign node31056 = (inp[11]) ? 4'b1100 : 4'b1101;
													assign node31059 = (inp[10]) ? node31067 : node31060;
														assign node31060 = (inp[9]) ? node31062 : 4'b1101;
															assign node31062 = (inp[11]) ? 4'b1100 : node31063;
																assign node31063 = (inp[0]) ? 4'b1101 : 4'b1100;
														assign node31067 = (inp[9]) ? node31073 : node31068;
															assign node31068 = (inp[0]) ? node31070 : 4'b1100;
																assign node31070 = (inp[11]) ? 4'b1100 : 4'b1101;
															assign node31073 = (inp[0]) ? node31075 : 4'b1101;
																assign node31075 = (inp[11]) ? 4'b1101 : 4'b1100;
												assign node31078 = (inp[0]) ? node31102 : node31079;
													assign node31079 = (inp[10]) ? node31087 : node31080;
														assign node31080 = (inp[9]) ? node31084 : node31081;
															assign node31081 = (inp[5]) ? 4'b1001 : 4'b1000;
															assign node31084 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node31087 = (inp[11]) ? node31095 : node31088;
															assign node31088 = (inp[9]) ? node31092 : node31089;
																assign node31089 = (inp[5]) ? 4'b1000 : 4'b1001;
																assign node31092 = (inp[5]) ? 4'b1001 : 4'b1000;
															assign node31095 = (inp[5]) ? node31099 : node31096;
																assign node31096 = (inp[9]) ? 4'b1000 : 4'b1001;
																assign node31099 = (inp[9]) ? 4'b1001 : 4'b1000;
													assign node31102 = (inp[9]) ? node31118 : node31103;
														assign node31103 = (inp[10]) ? node31111 : node31104;
															assign node31104 = (inp[11]) ? node31108 : node31105;
																assign node31105 = (inp[5]) ? 4'b1000 : 4'b1001;
																assign node31108 = (inp[5]) ? 4'b1001 : 4'b1000;
															assign node31111 = (inp[11]) ? node31115 : node31112;
																assign node31112 = (inp[5]) ? 4'b1001 : 4'b1000;
																assign node31115 = (inp[5]) ? 4'b1000 : 4'b1001;
														assign node31118 = (inp[5]) ? node31126 : node31119;
															assign node31119 = (inp[11]) ? node31123 : node31120;
																assign node31120 = (inp[10]) ? 4'b1001 : 4'b1000;
																assign node31123 = (inp[10]) ? 4'b1000 : 4'b1001;
															assign node31126 = (inp[10]) ? node31130 : node31127;
																assign node31127 = (inp[11]) ? 4'b1000 : 4'b1001;
																assign node31130 = (inp[11]) ? 4'b1001 : 4'b1000;
											assign node31133 = (inp[2]) ? node31183 : node31134;
												assign node31134 = (inp[11]) ? node31162 : node31135;
													assign node31135 = (inp[0]) ? node31149 : node31136;
														assign node31136 = (inp[5]) ? node31144 : node31137;
															assign node31137 = (inp[9]) ? node31141 : node31138;
																assign node31138 = (inp[10]) ? 4'b1001 : 4'b1000;
																assign node31141 = (inp[10]) ? 4'b1000 : 4'b1001;
															assign node31144 = (inp[10]) ? 4'b1001 : node31145;
																assign node31145 = (inp[9]) ? 4'b1000 : 4'b1001;
														assign node31149 = (inp[9]) ? node31155 : node31150;
															assign node31150 = (inp[5]) ? 4'b1000 : node31151;
																assign node31151 = (inp[10]) ? 4'b1001 : 4'b1000;
															assign node31155 = (inp[5]) ? node31159 : node31156;
																assign node31156 = (inp[10]) ? 4'b1000 : 4'b1001;
																assign node31159 = (inp[10]) ? 4'b1001 : 4'b1000;
													assign node31162 = (inp[9]) ? node31174 : node31163;
														assign node31163 = (inp[0]) ? node31169 : node31164;
															assign node31164 = (inp[5]) ? 4'b1001 : node31165;
																assign node31165 = (inp[10]) ? 4'b1000 : 4'b1001;
															assign node31169 = (inp[5]) ? 4'b1000 : node31170;
																assign node31170 = (inp[10]) ? 4'b1001 : 4'b1000;
														assign node31174 = (inp[0]) ? node31176 : 4'b1000;
															assign node31176 = (inp[10]) ? node31180 : node31177;
																assign node31177 = (inp[5]) ? 4'b1000 : 4'b1001;
																assign node31180 = (inp[5]) ? 4'b1001 : 4'b1000;
												assign node31183 = (inp[11]) ? node31213 : node31184;
													assign node31184 = (inp[0]) ? node31200 : node31185;
														assign node31185 = (inp[10]) ? node31193 : node31186;
															assign node31186 = (inp[5]) ? node31190 : node31187;
																assign node31187 = (inp[9]) ? 4'b1100 : 4'b1101;
																assign node31190 = (inp[9]) ? 4'b1101 : 4'b1100;
															assign node31193 = (inp[9]) ? node31197 : node31194;
																assign node31194 = (inp[5]) ? 4'b1101 : 4'b1100;
																assign node31197 = (inp[5]) ? 4'b1100 : 4'b1101;
														assign node31200 = (inp[5]) ? node31208 : node31201;
															assign node31201 = (inp[9]) ? node31205 : node31202;
																assign node31202 = (inp[10]) ? 4'b1101 : 4'b1100;
																assign node31205 = (inp[10]) ? 4'b1100 : 4'b1101;
															assign node31208 = (inp[10]) ? node31210 : 4'b1100;
																assign node31210 = (inp[9]) ? 4'b1101 : 4'b1100;
													assign node31213 = (inp[10]) ? node31221 : node31214;
														assign node31214 = (inp[5]) ? node31218 : node31215;
															assign node31215 = (inp[9]) ? 4'b1100 : 4'b1101;
															assign node31218 = (inp[9]) ? 4'b1101 : 4'b1100;
														assign node31221 = (inp[9]) ? node31225 : node31222;
															assign node31222 = (inp[5]) ? 4'b1101 : 4'b1100;
															assign node31225 = (inp[5]) ? 4'b1100 : 4'b1101;
								assign node31228 = (inp[11]) ? node31524 : node31229;
									assign node31229 = (inp[2]) ? node31397 : node31230;
										assign node31230 = (inp[13]) ? node31308 : node31231;
											assign node31231 = (inp[15]) ? node31279 : node31232;
												assign node31232 = (inp[5]) ? node31248 : node31233;
													assign node31233 = (inp[1]) ? node31241 : node31234;
														assign node31234 = (inp[0]) ? node31238 : node31235;
															assign node31235 = (inp[10]) ? 4'b1011 : 4'b1010;
															assign node31238 = (inp[10]) ? 4'b1010 : 4'b1011;
														assign node31241 = (inp[0]) ? node31245 : node31242;
															assign node31242 = (inp[10]) ? 4'b1111 : 4'b1110;
															assign node31245 = (inp[10]) ? 4'b1110 : 4'b1111;
													assign node31248 = (inp[1]) ? node31264 : node31249;
														assign node31249 = (inp[9]) ? node31257 : node31250;
															assign node31250 = (inp[0]) ? node31254 : node31251;
																assign node31251 = (inp[10]) ? 4'b1111 : 4'b1110;
																assign node31254 = (inp[10]) ? 4'b1110 : 4'b1111;
															assign node31257 = (inp[0]) ? node31261 : node31258;
																assign node31258 = (inp[10]) ? 4'b1111 : 4'b1110;
																assign node31261 = (inp[10]) ? 4'b1110 : 4'b1111;
														assign node31264 = (inp[9]) ? node31272 : node31265;
															assign node31265 = (inp[0]) ? node31269 : node31266;
																assign node31266 = (inp[10]) ? 4'b1010 : 4'b1011;
																assign node31269 = (inp[10]) ? 4'b1011 : 4'b1010;
															assign node31272 = (inp[0]) ? node31276 : node31273;
																assign node31273 = (inp[10]) ? 4'b1010 : 4'b1011;
																assign node31276 = (inp[10]) ? 4'b1011 : 4'b1010;
												assign node31279 = (inp[10]) ? node31293 : node31280;
													assign node31280 = (inp[0]) ? node31288 : node31281;
														assign node31281 = (inp[5]) ? node31285 : node31282;
															assign node31282 = (inp[1]) ? 4'b1011 : 4'b1110;
															assign node31285 = (inp[1]) ? 4'b1111 : 4'b1011;
														assign node31288 = (inp[5]) ? node31290 : 4'b1111;
															assign node31290 = (inp[1]) ? 4'b1110 : 4'b1010;
													assign node31293 = (inp[0]) ? node31301 : node31294;
														assign node31294 = (inp[1]) ? node31298 : node31295;
															assign node31295 = (inp[5]) ? 4'b1010 : 4'b1111;
															assign node31298 = (inp[5]) ? 4'b1110 : 4'b1010;
														assign node31301 = (inp[5]) ? node31305 : node31302;
															assign node31302 = (inp[1]) ? 4'b1011 : 4'b1110;
															assign node31305 = (inp[1]) ? 4'b1111 : 4'b1011;
											assign node31308 = (inp[15]) ? node31354 : node31309;
												assign node31309 = (inp[1]) ? node31331 : node31310;
													assign node31310 = (inp[5]) ? node31318 : node31311;
														assign node31311 = (inp[0]) ? node31315 : node31312;
															assign node31312 = (inp[10]) ? 4'b1011 : 4'b1010;
															assign node31315 = (inp[10]) ? 4'b1010 : 4'b1011;
														assign node31318 = (inp[9]) ? node31324 : node31319;
															assign node31319 = (inp[0]) ? 4'b1111 : node31320;
																assign node31320 = (inp[10]) ? 4'b1110 : 4'b1111;
															assign node31324 = (inp[0]) ? node31328 : node31325;
																assign node31325 = (inp[10]) ? 4'b1110 : 4'b1111;
																assign node31328 = (inp[10]) ? 4'b1111 : 4'b1110;
													assign node31331 = (inp[5]) ? node31347 : node31332;
														assign node31332 = (inp[9]) ? node31340 : node31333;
															assign node31333 = (inp[10]) ? node31337 : node31334;
																assign node31334 = (inp[0]) ? 4'b1111 : 4'b1110;
																assign node31337 = (inp[0]) ? 4'b1110 : 4'b1111;
															assign node31340 = (inp[0]) ? node31344 : node31341;
																assign node31341 = (inp[10]) ? 4'b1111 : 4'b1110;
																assign node31344 = (inp[10]) ? 4'b1110 : 4'b1111;
														assign node31347 = (inp[10]) ? node31351 : node31348;
															assign node31348 = (inp[0]) ? 4'b1010 : 4'b1011;
															assign node31351 = (inp[0]) ? 4'b1011 : 4'b1010;
												assign node31354 = (inp[5]) ? node31376 : node31355;
													assign node31355 = (inp[1]) ? node31369 : node31356;
														assign node31356 = (inp[9]) ? node31364 : node31357;
															assign node31357 = (inp[10]) ? node31361 : node31358;
																assign node31358 = (inp[0]) ? 4'b1110 : 4'b1111;
																assign node31361 = (inp[0]) ? 4'b1111 : 4'b1110;
															assign node31364 = (inp[10]) ? 4'b1111 : node31365;
																assign node31365 = (inp[0]) ? 4'b1110 : 4'b1111;
														assign node31369 = (inp[0]) ? node31373 : node31370;
															assign node31370 = (inp[10]) ? 4'b1011 : 4'b1010;
															assign node31373 = (inp[10]) ? 4'b1010 : 4'b1011;
													assign node31376 = (inp[1]) ? node31390 : node31377;
														assign node31377 = (inp[9]) ? node31383 : node31378;
															assign node31378 = (inp[10]) ? node31380 : 4'b1010;
																assign node31380 = (inp[0]) ? 4'b1010 : 4'b1011;
															assign node31383 = (inp[0]) ? node31387 : node31384;
																assign node31384 = (inp[10]) ? 4'b1011 : 4'b1010;
																assign node31387 = (inp[10]) ? 4'b1010 : 4'b1011;
														assign node31390 = (inp[10]) ? node31394 : node31391;
															assign node31391 = (inp[0]) ? 4'b1110 : 4'b1111;
															assign node31394 = (inp[0]) ? 4'b1111 : 4'b1110;
										assign node31397 = (inp[5]) ? node31469 : node31398;
											assign node31398 = (inp[1]) ? node31446 : node31399;
												assign node31399 = (inp[15]) ? node31415 : node31400;
													assign node31400 = (inp[0]) ? node31408 : node31401;
														assign node31401 = (inp[9]) ? node31403 : 4'b1110;
															assign node31403 = (inp[13]) ? node31405 : 4'b1110;
																assign node31405 = (inp[10]) ? 4'b1111 : 4'b1110;
														assign node31408 = (inp[10]) ? node31412 : node31409;
															assign node31409 = (inp[13]) ? 4'b1111 : 4'b1110;
															assign node31412 = (inp[13]) ? 4'b1110 : 4'b1111;
													assign node31415 = (inp[9]) ? node31431 : node31416;
														assign node31416 = (inp[10]) ? node31424 : node31417;
															assign node31417 = (inp[0]) ? node31421 : node31418;
																assign node31418 = (inp[13]) ? 4'b1011 : 4'b1010;
																assign node31421 = (inp[13]) ? 4'b1010 : 4'b1011;
															assign node31424 = (inp[0]) ? node31428 : node31425;
																assign node31425 = (inp[13]) ? 4'b1010 : 4'b1011;
																assign node31428 = (inp[13]) ? 4'b1011 : 4'b1010;
														assign node31431 = (inp[10]) ? node31439 : node31432;
															assign node31432 = (inp[0]) ? node31436 : node31433;
																assign node31433 = (inp[13]) ? 4'b1011 : 4'b1010;
																assign node31436 = (inp[13]) ? 4'b1010 : 4'b1011;
															assign node31439 = (inp[0]) ? node31443 : node31440;
																assign node31440 = (inp[13]) ? 4'b1010 : 4'b1011;
																assign node31443 = (inp[13]) ? 4'b1011 : 4'b1010;
												assign node31446 = (inp[15]) ? node31462 : node31447;
													assign node31447 = (inp[9]) ? node31455 : node31448;
														assign node31448 = (inp[0]) ? node31452 : node31449;
															assign node31449 = (inp[10]) ? 4'b1011 : 4'b1010;
															assign node31452 = (inp[10]) ? 4'b1010 : 4'b1011;
														assign node31455 = (inp[10]) ? node31459 : node31456;
															assign node31456 = (inp[0]) ? 4'b1011 : 4'b1010;
															assign node31459 = (inp[0]) ? 4'b1010 : 4'b1011;
													assign node31462 = (inp[10]) ? node31466 : node31463;
														assign node31463 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node31466 = (inp[0]) ? 4'b1110 : 4'b1111;
											assign node31469 = (inp[0]) ? node31495 : node31470;
												assign node31470 = (inp[15]) ? node31488 : node31471;
													assign node31471 = (inp[1]) ? node31479 : node31472;
														assign node31472 = (inp[9]) ? node31474 : 4'b1011;
															assign node31474 = (inp[13]) ? 4'b1010 : node31475;
																assign node31475 = (inp[10]) ? 4'b1011 : 4'b1010;
														assign node31479 = (inp[9]) ? 4'b1111 : node31480;
															assign node31480 = (inp[13]) ? node31484 : node31481;
																assign node31481 = (inp[10]) ? 4'b1111 : 4'b1110;
																assign node31484 = (inp[10]) ? 4'b1110 : 4'b1111;
													assign node31488 = (inp[1]) ? node31492 : node31489;
														assign node31489 = (inp[10]) ? 4'b1111 : 4'b1110;
														assign node31492 = (inp[10]) ? 4'b1010 : 4'b1011;
												assign node31495 = (inp[15]) ? node31517 : node31496;
													assign node31496 = (inp[1]) ? node31512 : node31497;
														assign node31497 = (inp[9]) ? node31505 : node31498;
															assign node31498 = (inp[10]) ? node31502 : node31499;
																assign node31499 = (inp[13]) ? 4'b1010 : 4'b1011;
																assign node31502 = (inp[13]) ? 4'b1011 : 4'b1010;
															assign node31505 = (inp[10]) ? node31509 : node31506;
																assign node31506 = (inp[13]) ? 4'b1010 : 4'b1011;
																assign node31509 = (inp[13]) ? 4'b1011 : 4'b1010;
														assign node31512 = (inp[13]) ? node31514 : 4'b1111;
															assign node31514 = (inp[10]) ? 4'b1111 : 4'b1110;
													assign node31517 = (inp[1]) ? node31521 : node31518;
														assign node31518 = (inp[10]) ? 4'b1110 : 4'b1111;
														assign node31521 = (inp[10]) ? 4'b1011 : 4'b1010;
									assign node31524 = (inp[15]) ? node31664 : node31525;
										assign node31525 = (inp[13]) ? node31597 : node31526;
											assign node31526 = (inp[10]) ? node31558 : node31527;
												assign node31527 = (inp[2]) ? node31543 : node31528;
													assign node31528 = (inp[0]) ? node31536 : node31529;
														assign node31529 = (inp[5]) ? node31533 : node31530;
															assign node31530 = (inp[1]) ? 4'b1111 : 4'b1011;
															assign node31533 = (inp[1]) ? 4'b1010 : 4'b1110;
														assign node31536 = (inp[5]) ? node31540 : node31537;
															assign node31537 = (inp[1]) ? 4'b1110 : 4'b1010;
															assign node31540 = (inp[1]) ? 4'b1011 : 4'b1111;
													assign node31543 = (inp[1]) ? node31551 : node31544;
														assign node31544 = (inp[5]) ? node31548 : node31545;
															assign node31545 = (inp[0]) ? 4'b1110 : 4'b1111;
															assign node31548 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node31551 = (inp[5]) ? node31555 : node31552;
															assign node31552 = (inp[0]) ? 4'b1010 : 4'b1011;
															assign node31555 = (inp[0]) ? 4'b1111 : 4'b1110;
												assign node31558 = (inp[5]) ? node31582 : node31559;
													assign node31559 = (inp[0]) ? node31575 : node31560;
														assign node31560 = (inp[9]) ? node31568 : node31561;
															assign node31561 = (inp[2]) ? node31565 : node31562;
																assign node31562 = (inp[1]) ? 4'b1110 : 4'b1010;
																assign node31565 = (inp[1]) ? 4'b1010 : 4'b1110;
															assign node31568 = (inp[2]) ? node31572 : node31569;
																assign node31569 = (inp[1]) ? 4'b1110 : 4'b1010;
																assign node31572 = (inp[1]) ? 4'b1010 : 4'b1110;
														assign node31575 = (inp[2]) ? node31579 : node31576;
															assign node31576 = (inp[1]) ? 4'b1111 : 4'b1011;
															assign node31579 = (inp[1]) ? 4'b1011 : 4'b1111;
													assign node31582 = (inp[0]) ? node31590 : node31583;
														assign node31583 = (inp[2]) ? node31587 : node31584;
															assign node31584 = (inp[1]) ? 4'b1011 : 4'b1111;
															assign node31587 = (inp[1]) ? 4'b1111 : 4'b1011;
														assign node31590 = (inp[2]) ? node31594 : node31591;
															assign node31591 = (inp[1]) ? 4'b1010 : 4'b1110;
															assign node31594 = (inp[1]) ? 4'b1110 : 4'b1010;
											assign node31597 = (inp[1]) ? node31627 : node31598;
												assign node31598 = (inp[0]) ? node31612 : node31599;
													assign node31599 = (inp[10]) ? node31605 : node31600;
														assign node31600 = (inp[2]) ? 4'b1010 : node31601;
															assign node31601 = (inp[5]) ? 4'b1110 : 4'b1010;
														assign node31605 = (inp[5]) ? node31609 : node31606;
															assign node31606 = (inp[2]) ? 4'b1110 : 4'b1011;
															assign node31609 = (inp[2]) ? 4'b1011 : 4'b1111;
													assign node31612 = (inp[10]) ? node31620 : node31613;
														assign node31613 = (inp[5]) ? node31617 : node31614;
															assign node31614 = (inp[2]) ? 4'b1110 : 4'b1011;
															assign node31617 = (inp[2]) ? 4'b1011 : 4'b1111;
														assign node31620 = (inp[5]) ? node31624 : node31621;
															assign node31621 = (inp[2]) ? 4'b1111 : 4'b1010;
															assign node31624 = (inp[2]) ? 4'b1010 : 4'b1110;
												assign node31627 = (inp[2]) ? node31649 : node31628;
													assign node31628 = (inp[5]) ? node31634 : node31629;
														assign node31629 = (inp[0]) ? node31631 : 4'b1111;
															assign node31631 = (inp[10]) ? 4'b1110 : 4'b1111;
														assign node31634 = (inp[9]) ? node31642 : node31635;
															assign node31635 = (inp[10]) ? node31639 : node31636;
																assign node31636 = (inp[0]) ? 4'b1010 : 4'b1011;
																assign node31639 = (inp[0]) ? 4'b1011 : 4'b1010;
															assign node31642 = (inp[0]) ? node31646 : node31643;
																assign node31643 = (inp[10]) ? 4'b1010 : 4'b1011;
																assign node31646 = (inp[10]) ? 4'b1011 : 4'b1010;
													assign node31649 = (inp[5]) ? node31657 : node31650;
														assign node31650 = (inp[10]) ? node31654 : node31651;
															assign node31651 = (inp[0]) ? 4'b1011 : 4'b1010;
															assign node31654 = (inp[0]) ? 4'b1010 : 4'b1011;
														assign node31657 = (inp[10]) ? node31661 : node31658;
															assign node31658 = (inp[0]) ? 4'b1111 : 4'b1110;
															assign node31661 = (inp[0]) ? 4'b1110 : 4'b1111;
										assign node31664 = (inp[1]) ? node31704 : node31665;
											assign node31665 = (inp[0]) ? node31685 : node31666;
												assign node31666 = (inp[10]) ? node31676 : node31667;
													assign node31667 = (inp[5]) ? node31671 : node31668;
														assign node31668 = (inp[2]) ? 4'b1011 : 4'b1111;
														assign node31671 = (inp[2]) ? node31673 : 4'b1010;
															assign node31673 = (inp[13]) ? 4'b1111 : 4'b1110;
													assign node31676 = (inp[5]) ? node31680 : node31677;
														assign node31677 = (inp[2]) ? 4'b1010 : 4'b1110;
														assign node31680 = (inp[2]) ? node31682 : 4'b1011;
															assign node31682 = (inp[13]) ? 4'b1110 : 4'b1111;
												assign node31685 = (inp[10]) ? node31695 : node31686;
													assign node31686 = (inp[5]) ? node31690 : node31687;
														assign node31687 = (inp[2]) ? 4'b1010 : 4'b1110;
														assign node31690 = (inp[2]) ? node31692 : 4'b1011;
															assign node31692 = (inp[13]) ? 4'b1110 : 4'b1111;
													assign node31695 = (inp[5]) ? node31699 : node31696;
														assign node31696 = (inp[2]) ? 4'b1011 : 4'b1111;
														assign node31699 = (inp[2]) ? node31701 : 4'b1010;
															assign node31701 = (inp[13]) ? 4'b1111 : 4'b1110;
											assign node31704 = (inp[2]) ? node31734 : node31705;
												assign node31705 = (inp[5]) ? node31711 : node31706;
													assign node31706 = (inp[0]) ? 4'b1010 : node31707;
														assign node31707 = (inp[10]) ? 4'b1011 : 4'b1010;
													assign node31711 = (inp[0]) ? node31727 : node31712;
														assign node31712 = (inp[9]) ? node31720 : node31713;
															assign node31713 = (inp[10]) ? node31717 : node31714;
																assign node31714 = (inp[13]) ? 4'b1110 : 4'b1111;
																assign node31717 = (inp[13]) ? 4'b1111 : 4'b1110;
															assign node31720 = (inp[13]) ? node31724 : node31721;
																assign node31721 = (inp[10]) ? 4'b1110 : 4'b1111;
																assign node31724 = (inp[10]) ? 4'b1111 : 4'b1110;
														assign node31727 = (inp[13]) ? node31731 : node31728;
															assign node31728 = (inp[10]) ? 4'b1111 : 4'b1110;
															assign node31731 = (inp[10]) ? 4'b1110 : 4'b1111;
												assign node31734 = (inp[5]) ? node31756 : node31735;
													assign node31735 = (inp[0]) ? node31749 : node31736;
														assign node31736 = (inp[9]) ? node31744 : node31737;
															assign node31737 = (inp[13]) ? node31741 : node31738;
																assign node31738 = (inp[10]) ? 4'b1111 : 4'b1110;
																assign node31741 = (inp[10]) ? 4'b1110 : 4'b1111;
															assign node31744 = (inp[10]) ? 4'b1111 : node31745;
																assign node31745 = (inp[13]) ? 4'b1111 : 4'b1110;
														assign node31749 = (inp[13]) ? node31753 : node31750;
															assign node31750 = (inp[10]) ? 4'b1110 : 4'b1111;
															assign node31753 = (inp[10]) ? 4'b1111 : 4'b1110;
													assign node31756 = (inp[13]) ? node31764 : node31757;
														assign node31757 = (inp[10]) ? node31761 : node31758;
															assign node31758 = (inp[0]) ? 4'b1010 : 4'b1011;
															assign node31761 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node31764 = (inp[0]) ? node31768 : node31765;
															assign node31765 = (inp[10]) ? 4'b1011 : 4'b1010;
															assign node31768 = (inp[10]) ? 4'b1010 : 4'b1011;
							assign node31771 = (inp[11]) ? node32313 : node31772;
								assign node31772 = (inp[9]) ? node32046 : node31773;
									assign node31773 = (inp[10]) ? node31925 : node31774;
										assign node31774 = (inp[8]) ? node31856 : node31775;
											assign node31775 = (inp[0]) ? node31815 : node31776;
												assign node31776 = (inp[1]) ? node31804 : node31777;
													assign node31777 = (inp[5]) ? node31791 : node31778;
														assign node31778 = (inp[15]) ? node31786 : node31779;
															assign node31779 = (inp[2]) ? node31783 : node31780;
																assign node31780 = (inp[13]) ? 4'b1110 : 4'b1010;
																assign node31783 = (inp[13]) ? 4'b1010 : 4'b1111;
															assign node31786 = (inp[13]) ? node31788 : 4'b1110;
																assign node31788 = (inp[2]) ? 4'b1011 : 4'b1111;
														assign node31791 = (inp[2]) ? node31799 : node31792;
															assign node31792 = (inp[13]) ? node31796 : node31793;
																assign node31793 = (inp[15]) ? 4'b1110 : 4'b1111;
																assign node31796 = (inp[15]) ? 4'b1011 : 4'b1010;
															assign node31799 = (inp[13]) ? 4'b1111 : node31800;
																assign node31800 = (inp[15]) ? 4'b1010 : 4'b1011;
													assign node31804 = (inp[13]) ? node31812 : node31805;
														assign node31805 = (inp[2]) ? node31809 : node31806;
															assign node31806 = (inp[15]) ? 4'b1011 : 4'b1010;
															assign node31809 = (inp[15]) ? 4'b1110 : 4'b1111;
														assign node31812 = (inp[2]) ? 4'b1010 : 4'b1110;
												assign node31815 = (inp[15]) ? node31835 : node31816;
													assign node31816 = (inp[2]) ? node31824 : node31817;
														assign node31817 = (inp[13]) ? 4'b1110 : node31818;
															assign node31818 = (inp[1]) ? 4'b1010 : node31819;
																assign node31819 = (inp[5]) ? 4'b1110 : 4'b1010;
														assign node31824 = (inp[13]) ? node31830 : node31825;
															assign node31825 = (inp[5]) ? node31827 : 4'b1110;
																assign node31827 = (inp[1]) ? 4'b1110 : 4'b1010;
															assign node31830 = (inp[1]) ? 4'b1010 : node31831;
																assign node31831 = (inp[5]) ? 4'b1110 : 4'b1010;
													assign node31835 = (inp[13]) ? node31845 : node31836;
														assign node31836 = (inp[1]) ? 4'b1111 : node31837;
															assign node31837 = (inp[5]) ? node31841 : node31838;
																assign node31838 = (inp[2]) ? 4'b1110 : 4'b1011;
																assign node31841 = (inp[2]) ? 4'b1010 : 4'b1110;
														assign node31845 = (inp[2]) ? node31851 : node31846;
															assign node31846 = (inp[5]) ? node31848 : 4'b1110;
																assign node31848 = (inp[1]) ? 4'b1110 : 4'b1010;
															assign node31851 = (inp[1]) ? 4'b1010 : node31852;
																assign node31852 = (inp[5]) ? 4'b1111 : 4'b1010;
											assign node31856 = (inp[0]) ? node31894 : node31857;
												assign node31857 = (inp[15]) ? node31879 : node31858;
													assign node31858 = (inp[13]) ? node31866 : node31859;
														assign node31859 = (inp[1]) ? node31863 : node31860;
															assign node31860 = (inp[2]) ? 4'b1111 : 4'b1010;
															assign node31863 = (inp[2]) ? 4'b1010 : 4'b1110;
														assign node31866 = (inp[5]) ? node31872 : node31867;
															assign node31867 = (inp[1]) ? 4'b1010 : node31868;
																assign node31868 = (inp[2]) ? 4'b1110 : 4'b1010;
															assign node31872 = (inp[1]) ? node31876 : node31873;
																assign node31873 = (inp[2]) ? 4'b1110 : 4'b1010;
																assign node31876 = (inp[2]) ? 4'b1010 : 4'b1110;
													assign node31879 = (inp[13]) ? node31887 : node31880;
														assign node31880 = (inp[1]) ? node31884 : node31881;
															assign node31881 = (inp[2]) ? 4'b1110 : 4'b1010;
															assign node31884 = (inp[2]) ? 4'b1011 : 4'b1111;
														assign node31887 = (inp[1]) ? node31891 : node31888;
															assign node31888 = (inp[2]) ? 4'b1111 : 4'b1010;
															assign node31891 = (inp[2]) ? 4'b1010 : 4'b1110;
												assign node31894 = (inp[13]) ? node31908 : node31895;
													assign node31895 = (inp[1]) ? node31901 : node31896;
														assign node31896 = (inp[2]) ? node31898 : 4'b1011;
															assign node31898 = (inp[15]) ? 4'b1111 : 4'b1110;
														assign node31901 = (inp[2]) ? node31905 : node31902;
															assign node31902 = (inp[15]) ? 4'b1110 : 4'b1111;
															assign node31905 = (inp[15]) ? 4'b1010 : 4'b1011;
													assign node31908 = (inp[5]) ? node31916 : node31909;
														assign node31909 = (inp[2]) ? node31913 : node31910;
															assign node31910 = (inp[1]) ? 4'b1111 : 4'b1011;
															assign node31913 = (inp[1]) ? 4'b1011 : 4'b1111;
														assign node31916 = (inp[15]) ? node31922 : node31917;
															assign node31917 = (inp[1]) ? 4'b1111 : node31918;
																assign node31918 = (inp[2]) ? 4'b1111 : 4'b1011;
															assign node31922 = (inp[1]) ? 4'b1011 : 4'b1110;
										assign node31925 = (inp[8]) ? node31987 : node31926;
											assign node31926 = (inp[13]) ? node31960 : node31927;
												assign node31927 = (inp[2]) ? node31941 : node31928;
													assign node31928 = (inp[1]) ? node31938 : node31929;
														assign node31929 = (inp[5]) ? node31933 : node31930;
															assign node31930 = (inp[0]) ? 4'b1010 : 4'b1011;
															assign node31933 = (inp[0]) ? 4'b1111 : node31934;
																assign node31934 = (inp[15]) ? 4'b1111 : 4'b1110;
														assign node31938 = (inp[15]) ? 4'b1010 : 4'b1011;
													assign node31941 = (inp[1]) ? node31953 : node31942;
														assign node31942 = (inp[5]) ? node31948 : node31943;
															assign node31943 = (inp[15]) ? 4'b1111 : node31944;
																assign node31944 = (inp[0]) ? 4'b1111 : 4'b1110;
															assign node31948 = (inp[15]) ? 4'b1011 : node31949;
																assign node31949 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node31953 = (inp[0]) ? node31957 : node31954;
															assign node31954 = (inp[15]) ? 4'b1111 : 4'b1110;
															assign node31957 = (inp[15]) ? 4'b1110 : 4'b1111;
												assign node31960 = (inp[2]) ? node31974 : node31961;
													assign node31961 = (inp[1]) ? 4'b1111 : node31962;
														assign node31962 = (inp[5]) ? node31968 : node31963;
															assign node31963 = (inp[15]) ? node31965 : 4'b1111;
																assign node31965 = (inp[0]) ? 4'b1111 : 4'b1110;
															assign node31968 = (inp[15]) ? node31970 : 4'b1011;
																assign node31970 = (inp[0]) ? 4'b1011 : 4'b1010;
													assign node31974 = (inp[1]) ? 4'b1011 : node31975;
														assign node31975 = (inp[5]) ? node31981 : node31976;
															assign node31976 = (inp[0]) ? 4'b1011 : node31977;
																assign node31977 = (inp[15]) ? 4'b1010 : 4'b1011;
															assign node31981 = (inp[0]) ? node31983 : 4'b1110;
																assign node31983 = (inp[15]) ? 4'b1110 : 4'b1111;
											assign node31987 = (inp[0]) ? node32009 : node31988;
												assign node31988 = (inp[13]) ? node32000 : node31989;
													assign node31989 = (inp[2]) ? node31995 : node31990;
														assign node31990 = (inp[1]) ? node31992 : 4'b1011;
															assign node31992 = (inp[15]) ? 4'b1110 : 4'b1111;
														assign node31995 = (inp[1]) ? node31997 : 4'b1110;
															assign node31997 = (inp[15]) ? 4'b1010 : 4'b1011;
													assign node32000 = (inp[2]) ? node32004 : node32001;
														assign node32001 = (inp[1]) ? 4'b1111 : 4'b1011;
														assign node32004 = (inp[1]) ? 4'b1011 : node32005;
															assign node32005 = (inp[15]) ? 4'b1110 : 4'b1111;
												assign node32009 = (inp[15]) ? node32033 : node32010;
													assign node32010 = (inp[13]) ? node32018 : node32011;
														assign node32011 = (inp[1]) ? node32015 : node32012;
															assign node32012 = (inp[2]) ? 4'b1111 : 4'b1010;
															assign node32015 = (inp[2]) ? 4'b1010 : 4'b1110;
														assign node32018 = (inp[5]) ? node32026 : node32019;
															assign node32019 = (inp[1]) ? node32023 : node32020;
																assign node32020 = (inp[2]) ? 4'b1110 : 4'b1010;
																assign node32023 = (inp[2]) ? 4'b1010 : 4'b1110;
															assign node32026 = (inp[2]) ? node32030 : node32027;
																assign node32027 = (inp[1]) ? 4'b1110 : 4'b1010;
																assign node32030 = (inp[1]) ? 4'b1010 : 4'b1110;
													assign node32033 = (inp[1]) ? node32039 : node32034;
														assign node32034 = (inp[2]) ? node32036 : 4'b1010;
															assign node32036 = (inp[13]) ? 4'b1111 : 4'b1110;
														assign node32039 = (inp[13]) ? node32043 : node32040;
															assign node32040 = (inp[2]) ? 4'b1011 : 4'b1111;
															assign node32043 = (inp[2]) ? 4'b1010 : 4'b1110;
									assign node32046 = (inp[10]) ? node32180 : node32047;
										assign node32047 = (inp[0]) ? node32111 : node32048;
											assign node32048 = (inp[8]) ? node32088 : node32049;
												assign node32049 = (inp[13]) ? node32071 : node32050;
													assign node32050 = (inp[15]) ? node32060 : node32051;
														assign node32051 = (inp[2]) ? node32055 : node32052;
															assign node32052 = (inp[1]) ? 4'b1011 : 4'b1110;
															assign node32055 = (inp[1]) ? 4'b1110 : node32056;
																assign node32056 = (inp[5]) ? 4'b1010 : 4'b1110;
														assign node32060 = (inp[2]) ? node32066 : node32061;
															assign node32061 = (inp[1]) ? 4'b1010 : node32062;
																assign node32062 = (inp[5]) ? 4'b1111 : 4'b1011;
															assign node32066 = (inp[1]) ? 4'b1111 : node32067;
																assign node32067 = (inp[5]) ? 4'b1011 : 4'b1111;
													assign node32071 = (inp[1]) ? node32085 : node32072;
														assign node32072 = (inp[15]) ? node32080 : node32073;
															assign node32073 = (inp[2]) ? node32077 : node32074;
																assign node32074 = (inp[5]) ? 4'b1011 : 4'b1111;
																assign node32077 = (inp[5]) ? 4'b1110 : 4'b1011;
															assign node32080 = (inp[2]) ? 4'b1010 : node32081;
																assign node32081 = (inp[5]) ? 4'b1010 : 4'b1110;
														assign node32085 = (inp[2]) ? 4'b1011 : 4'b1111;
												assign node32088 = (inp[13]) ? node32102 : node32089;
													assign node32089 = (inp[1]) ? node32095 : node32090;
														assign node32090 = (inp[2]) ? node32092 : 4'b1010;
															assign node32092 = (inp[15]) ? 4'b1110 : 4'b1111;
														assign node32095 = (inp[15]) ? node32099 : node32096;
															assign node32096 = (inp[2]) ? 4'b1010 : 4'b1110;
															assign node32099 = (inp[2]) ? 4'b1011 : 4'b1111;
													assign node32102 = (inp[1]) ? node32108 : node32103;
														assign node32103 = (inp[2]) ? node32105 : 4'b1010;
															assign node32105 = (inp[15]) ? 4'b1111 : 4'b1110;
														assign node32108 = (inp[2]) ? 4'b1010 : 4'b1110;
											assign node32111 = (inp[15]) ? node32145 : node32112;
												assign node32112 = (inp[2]) ? node32128 : node32113;
													assign node32113 = (inp[1]) ? node32123 : node32114;
														assign node32114 = (inp[8]) ? 4'b1011 : node32115;
															assign node32115 = (inp[5]) ? node32119 : node32116;
																assign node32116 = (inp[13]) ? 4'b1111 : 4'b1011;
																assign node32119 = (inp[13]) ? 4'b1011 : 4'b1111;
														assign node32123 = (inp[13]) ? 4'b1111 : node32124;
															assign node32124 = (inp[8]) ? 4'b1111 : 4'b1011;
													assign node32128 = (inp[1]) ? node32140 : node32129;
														assign node32129 = (inp[8]) ? node32137 : node32130;
															assign node32130 = (inp[13]) ? node32134 : node32131;
																assign node32131 = (inp[5]) ? 4'b1011 : 4'b1111;
																assign node32134 = (inp[5]) ? 4'b1111 : 4'b1011;
															assign node32137 = (inp[13]) ? 4'b1111 : 4'b1110;
														assign node32140 = (inp[8]) ? 4'b1011 : node32141;
															assign node32141 = (inp[13]) ? 4'b1011 : 4'b1111;
												assign node32145 = (inp[13]) ? node32165 : node32146;
													assign node32146 = (inp[1]) ? node32160 : node32147;
														assign node32147 = (inp[2]) ? node32155 : node32148;
															assign node32148 = (inp[5]) ? node32152 : node32149;
																assign node32149 = (inp[8]) ? 4'b1011 : 4'b1010;
																assign node32152 = (inp[8]) ? 4'b1011 : 4'b1111;
															assign node32155 = (inp[8]) ? 4'b1111 : node32156;
																assign node32156 = (inp[5]) ? 4'b1011 : 4'b1111;
														assign node32160 = (inp[8]) ? node32162 : 4'b1010;
															assign node32162 = (inp[2]) ? 4'b1010 : 4'b1110;
													assign node32165 = (inp[2]) ? node32173 : node32166;
														assign node32166 = (inp[1]) ? 4'b1111 : node32167;
															assign node32167 = (inp[8]) ? 4'b1011 : node32168;
																assign node32168 = (inp[5]) ? 4'b1011 : 4'b1111;
														assign node32173 = (inp[1]) ? 4'b1011 : node32174;
															assign node32174 = (inp[5]) ? 4'b1110 : node32175;
																assign node32175 = (inp[8]) ? 4'b1110 : 4'b1011;
										assign node32180 = (inp[0]) ? node32242 : node32181;
											assign node32181 = (inp[8]) ? node32219 : node32182;
												assign node32182 = (inp[1]) ? node32208 : node32183;
													assign node32183 = (inp[2]) ? node32193 : node32184;
														assign node32184 = (inp[15]) ? node32190 : node32185;
															assign node32185 = (inp[5]) ? 4'b1111 : node32186;
																assign node32186 = (inp[13]) ? 4'b1110 : 4'b1010;
															assign node32190 = (inp[5]) ? 4'b1110 : 4'b1111;
														assign node32193 = (inp[15]) ? node32201 : node32194;
															assign node32194 = (inp[13]) ? node32198 : node32195;
																assign node32195 = (inp[5]) ? 4'b1011 : 4'b1111;
																assign node32198 = (inp[5]) ? 4'b1111 : 4'b1010;
															assign node32201 = (inp[13]) ? node32205 : node32202;
																assign node32202 = (inp[5]) ? 4'b1010 : 4'b1110;
																assign node32205 = (inp[5]) ? 4'b1111 : 4'b1011;
													assign node32208 = (inp[13]) ? node32216 : node32209;
														assign node32209 = (inp[2]) ? node32213 : node32210;
															assign node32210 = (inp[15]) ? 4'b1011 : 4'b1010;
															assign node32213 = (inp[15]) ? 4'b1110 : 4'b1111;
														assign node32216 = (inp[2]) ? 4'b1010 : 4'b1110;
												assign node32219 = (inp[15]) ? node32229 : node32220;
													assign node32220 = (inp[1]) ? node32226 : node32221;
														assign node32221 = (inp[2]) ? node32223 : 4'b1011;
															assign node32223 = (inp[13]) ? 4'b1111 : 4'b1110;
														assign node32226 = (inp[2]) ? 4'b1011 : 4'b1111;
													assign node32229 = (inp[2]) ? node32235 : node32230;
														assign node32230 = (inp[1]) ? node32232 : 4'b1011;
															assign node32232 = (inp[13]) ? 4'b1111 : 4'b1110;
														assign node32235 = (inp[1]) ? node32239 : node32236;
															assign node32236 = (inp[13]) ? 4'b1110 : 4'b1111;
															assign node32239 = (inp[5]) ? 4'b1011 : 4'b1010;
											assign node32242 = (inp[15]) ? node32276 : node32243;
												assign node32243 = (inp[8]) ? node32261 : node32244;
													assign node32244 = (inp[13]) ? node32256 : node32245;
														assign node32245 = (inp[2]) ? node32251 : node32246;
															assign node32246 = (inp[1]) ? 4'b1010 : node32247;
																assign node32247 = (inp[5]) ? 4'b1110 : 4'b1010;
															assign node32251 = (inp[1]) ? 4'b1110 : node32252;
																assign node32252 = (inp[5]) ? 4'b1010 : 4'b1110;
														assign node32256 = (inp[2]) ? 4'b1010 : node32257;
															assign node32257 = (inp[1]) ? 4'b1110 : 4'b1010;
													assign node32261 = (inp[13]) ? node32269 : node32262;
														assign node32262 = (inp[2]) ? node32266 : node32263;
															assign node32263 = (inp[1]) ? 4'b1110 : 4'b1010;
															assign node32266 = (inp[1]) ? 4'b1010 : 4'b1111;
														assign node32269 = (inp[2]) ? node32273 : node32270;
															assign node32270 = (inp[1]) ? 4'b1110 : 4'b1010;
															assign node32273 = (inp[1]) ? 4'b1010 : 4'b1110;
												assign node32276 = (inp[13]) ? node32302 : node32277;
													assign node32277 = (inp[1]) ? node32287 : node32278;
														assign node32278 = (inp[2]) ? node32282 : node32279;
															assign node32279 = (inp[8]) ? 4'b1010 : 4'b1011;
															assign node32282 = (inp[8]) ? 4'b1110 : node32283;
																assign node32283 = (inp[5]) ? 4'b1010 : 4'b1110;
														assign node32287 = (inp[5]) ? node32295 : node32288;
															assign node32288 = (inp[8]) ? node32292 : node32289;
																assign node32289 = (inp[2]) ? 4'b1111 : 4'b1011;
																assign node32292 = (inp[2]) ? 4'b1011 : 4'b1111;
															assign node32295 = (inp[2]) ? node32299 : node32296;
																assign node32296 = (inp[8]) ? 4'b1111 : 4'b1011;
																assign node32299 = (inp[8]) ? 4'b1011 : 4'b1111;
													assign node32302 = (inp[1]) ? node32310 : node32303;
														assign node32303 = (inp[2]) ? node32305 : 4'b1010;
															assign node32305 = (inp[8]) ? 4'b1111 : node32306;
																assign node32306 = (inp[5]) ? 4'b1111 : 4'b1010;
														assign node32310 = (inp[2]) ? 4'b1010 : 4'b1110;
								assign node32313 = (inp[9]) ? node32603 : node32314;
									assign node32314 = (inp[10]) ? node32452 : node32315;
										assign node32315 = (inp[0]) ? node32395 : node32316;
											assign node32316 = (inp[15]) ? node32354 : node32317;
												assign node32317 = (inp[8]) ? node32335 : node32318;
													assign node32318 = (inp[13]) ? node32328 : node32319;
														assign node32319 = (inp[2]) ? node32325 : node32320;
															assign node32320 = (inp[1]) ? 4'b1011 : node32321;
																assign node32321 = (inp[5]) ? 4'b1111 : 4'b1011;
															assign node32325 = (inp[5]) ? 4'b1011 : 4'b1111;
														assign node32328 = (inp[2]) ? node32330 : 4'b1111;
															assign node32330 = (inp[5]) ? node32332 : 4'b1011;
																assign node32332 = (inp[1]) ? 4'b1011 : 4'b1111;
													assign node32335 = (inp[13]) ? node32347 : node32336;
														assign node32336 = (inp[5]) ? node32342 : node32337;
															assign node32337 = (inp[2]) ? 4'b1111 : node32338;
																assign node32338 = (inp[1]) ? 4'b1111 : 4'b1011;
															assign node32342 = (inp[1]) ? 4'b1011 : node32343;
																assign node32343 = (inp[2]) ? 4'b1111 : 4'b1011;
														assign node32347 = (inp[5]) ? 4'b1010 : node32348;
															assign node32348 = (inp[1]) ? node32350 : 4'b1111;
																assign node32350 = (inp[2]) ? 4'b1010 : 4'b1110;
												assign node32354 = (inp[1]) ? node32372 : node32355;
													assign node32355 = (inp[2]) ? node32363 : node32356;
														assign node32356 = (inp[13]) ? 4'b1011 : node32357;
															assign node32357 = (inp[8]) ? 4'b1010 : node32358;
																assign node32358 = (inp[5]) ? 4'b1111 : 4'b1010;
														assign node32363 = (inp[8]) ? 4'b1111 : node32364;
															assign node32364 = (inp[5]) ? node32368 : node32365;
																assign node32365 = (inp[13]) ? 4'b1011 : 4'b1111;
																assign node32368 = (inp[13]) ? 4'b1110 : 4'b1011;
													assign node32372 = (inp[13]) ? node32388 : node32373;
														assign node32373 = (inp[5]) ? node32381 : node32374;
															assign node32374 = (inp[8]) ? node32378 : node32375;
																assign node32375 = (inp[2]) ? 4'b1110 : 4'b1010;
																assign node32378 = (inp[2]) ? 4'b1010 : 4'b1110;
															assign node32381 = (inp[2]) ? node32385 : node32382;
																assign node32382 = (inp[8]) ? 4'b1110 : 4'b1010;
																assign node32385 = (inp[8]) ? 4'b1010 : 4'b1110;
														assign node32388 = (inp[8]) ? node32392 : node32389;
															assign node32389 = (inp[2]) ? 4'b1011 : 4'b1111;
															assign node32392 = (inp[2]) ? 4'b1010 : 4'b1110;
											assign node32395 = (inp[1]) ? node32429 : node32396;
												assign node32396 = (inp[2]) ? node32418 : node32397;
													assign node32397 = (inp[8]) ? node32411 : node32398;
														assign node32398 = (inp[5]) ? node32404 : node32399;
															assign node32399 = (inp[13]) ? node32401 : 4'b1010;
																assign node32401 = (inp[15]) ? 4'b1111 : 4'b1110;
															assign node32404 = (inp[13]) ? node32408 : node32405;
																assign node32405 = (inp[15]) ? 4'b1110 : 4'b1111;
																assign node32408 = (inp[15]) ? 4'b1011 : 4'b1010;
														assign node32411 = (inp[15]) ? node32415 : node32412;
															assign node32412 = (inp[13]) ? 4'b1011 : 4'b1010;
															assign node32415 = (inp[13]) ? 4'b1010 : 4'b1011;
													assign node32418 = (inp[8]) ? 4'b1110 : node32419;
														assign node32419 = (inp[13]) ? 4'b1111 : node32420;
															assign node32420 = (inp[5]) ? node32424 : node32421;
																assign node32421 = (inp[15]) ? 4'b1110 : 4'b1111;
																assign node32424 = (inp[15]) ? 4'b1010 : 4'b1011;
												assign node32429 = (inp[2]) ? node32441 : node32430;
													assign node32430 = (inp[8]) ? node32436 : node32431;
														assign node32431 = (inp[13]) ? 4'b1110 : node32432;
															assign node32432 = (inp[15]) ? 4'b1011 : 4'b1010;
														assign node32436 = (inp[13]) ? 4'b1111 : node32437;
															assign node32437 = (inp[15]) ? 4'b1111 : 4'b1110;
													assign node32441 = (inp[8]) ? node32447 : node32442;
														assign node32442 = (inp[13]) ? 4'b1010 : node32443;
															assign node32443 = (inp[15]) ? 4'b1110 : 4'b1111;
														assign node32447 = (inp[15]) ? 4'b1011 : node32448;
															assign node32448 = (inp[13]) ? 4'b1011 : 4'b1010;
										assign node32452 = (inp[0]) ? node32528 : node32453;
											assign node32453 = (inp[15]) ? node32499 : node32454;
												assign node32454 = (inp[13]) ? node32478 : node32455;
													assign node32455 = (inp[8]) ? node32463 : node32456;
														assign node32456 = (inp[1]) ? node32460 : node32457;
															assign node32457 = (inp[2]) ? 4'b1010 : 4'b1110;
															assign node32460 = (inp[2]) ? 4'b1110 : 4'b1010;
														assign node32463 = (inp[5]) ? node32471 : node32464;
															assign node32464 = (inp[1]) ? node32468 : node32465;
																assign node32465 = (inp[2]) ? 4'b1110 : 4'b1010;
																assign node32468 = (inp[2]) ? 4'b1010 : 4'b1110;
															assign node32471 = (inp[1]) ? node32475 : node32472;
																assign node32472 = (inp[2]) ? 4'b1110 : 4'b1010;
																assign node32475 = (inp[2]) ? 4'b1010 : 4'b1110;
													assign node32478 = (inp[8]) ? node32490 : node32479;
														assign node32479 = (inp[2]) ? node32485 : node32480;
															assign node32480 = (inp[5]) ? node32482 : 4'b1110;
																assign node32482 = (inp[1]) ? 4'b1110 : 4'b1010;
															assign node32485 = (inp[1]) ? 4'b1010 : node32486;
																assign node32486 = (inp[5]) ? 4'b1110 : 4'b1010;
														assign node32490 = (inp[5]) ? node32492 : 4'b1011;
															assign node32492 = (inp[1]) ? node32496 : node32493;
																assign node32493 = (inp[2]) ? 4'b1110 : 4'b1011;
																assign node32496 = (inp[2]) ? 4'b1011 : 4'b1111;
												assign node32499 = (inp[1]) ? node32517 : node32500;
													assign node32500 = (inp[2]) ? node32508 : node32501;
														assign node32501 = (inp[13]) ? node32503 : 4'b1011;
															assign node32503 = (inp[5]) ? 4'b1010 : node32504;
																assign node32504 = (inp[8]) ? 4'b1010 : 4'b1110;
														assign node32508 = (inp[8]) ? 4'b1110 : node32509;
															assign node32509 = (inp[13]) ? node32513 : node32510;
																assign node32510 = (inp[5]) ? 4'b1010 : 4'b1110;
																assign node32513 = (inp[5]) ? 4'b1111 : 4'b1010;
													assign node32517 = (inp[2]) ? node32523 : node32518;
														assign node32518 = (inp[8]) ? 4'b1111 : node32519;
															assign node32519 = (inp[13]) ? 4'b1110 : 4'b1011;
														assign node32523 = (inp[8]) ? 4'b1011 : node32524;
															assign node32524 = (inp[13]) ? 4'b1010 : 4'b1111;
											assign node32528 = (inp[15]) ? node32570 : node32529;
												assign node32529 = (inp[13]) ? node32551 : node32530;
													assign node32530 = (inp[8]) ? node32536 : node32531;
														assign node32531 = (inp[2]) ? node32533 : 4'b1011;
															assign node32533 = (inp[5]) ? 4'b1010 : 4'b1110;
														assign node32536 = (inp[5]) ? node32544 : node32537;
															assign node32537 = (inp[2]) ? node32541 : node32538;
																assign node32538 = (inp[1]) ? 4'b1111 : 4'b1011;
																assign node32541 = (inp[1]) ? 4'b1011 : 4'b1111;
															assign node32544 = (inp[1]) ? node32548 : node32545;
																assign node32545 = (inp[2]) ? 4'b1111 : 4'b1011;
																assign node32548 = (inp[2]) ? 4'b1011 : 4'b1111;
													assign node32551 = (inp[8]) ? node32563 : node32552;
														assign node32552 = (inp[2]) ? node32558 : node32553;
															assign node32553 = (inp[5]) ? node32555 : 4'b1111;
																assign node32555 = (inp[1]) ? 4'b1111 : 4'b1011;
															assign node32558 = (inp[1]) ? 4'b1011 : node32559;
																assign node32559 = (inp[5]) ? 4'b1110 : 4'b1011;
														assign node32563 = (inp[1]) ? node32567 : node32564;
															assign node32564 = (inp[2]) ? 4'b1111 : 4'b1010;
															assign node32567 = (inp[2]) ? 4'b1010 : 4'b1110;
												assign node32570 = (inp[8]) ? node32594 : node32571;
													assign node32571 = (inp[13]) ? node32583 : node32572;
														assign node32572 = (inp[2]) ? node32578 : node32573;
															assign node32573 = (inp[1]) ? 4'b1010 : node32574;
																assign node32574 = (inp[5]) ? 4'b1111 : 4'b1011;
															assign node32578 = (inp[1]) ? 4'b1111 : node32579;
																assign node32579 = (inp[5]) ? 4'b1011 : 4'b1111;
														assign node32583 = (inp[1]) ? node32591 : node32584;
															assign node32584 = (inp[2]) ? node32588 : node32585;
																assign node32585 = (inp[5]) ? 4'b1010 : 4'b1110;
																assign node32588 = (inp[5]) ? 4'b1110 : 4'b1010;
															assign node32591 = (inp[2]) ? 4'b1011 : 4'b1111;
													assign node32594 = (inp[1]) ? node32600 : node32595;
														assign node32595 = (inp[2]) ? 4'b1111 : node32596;
															assign node32596 = (inp[13]) ? 4'b1011 : 4'b1010;
														assign node32600 = (inp[2]) ? 4'b1010 : 4'b1110;
									assign node32603 = (inp[10]) ? node32725 : node32604;
										assign node32604 = (inp[0]) ? node32672 : node32605;
											assign node32605 = (inp[8]) ? node32651 : node32606;
												assign node32606 = (inp[15]) ? node32630 : node32607;
													assign node32607 = (inp[1]) ? node32623 : node32608;
														assign node32608 = (inp[2]) ? node32616 : node32609;
															assign node32609 = (inp[13]) ? node32613 : node32610;
																assign node32610 = (inp[5]) ? 4'b1110 : 4'b1010;
																assign node32613 = (inp[5]) ? 4'b1010 : 4'b1110;
															assign node32616 = (inp[5]) ? node32620 : node32617;
																assign node32617 = (inp[13]) ? 4'b1010 : 4'b1110;
																assign node32620 = (inp[13]) ? 4'b1110 : 4'b1010;
														assign node32623 = (inp[2]) ? node32627 : node32624;
															assign node32624 = (inp[13]) ? 4'b1110 : 4'b1010;
															assign node32627 = (inp[13]) ? 4'b1010 : 4'b1110;
													assign node32630 = (inp[13]) ? node32640 : node32631;
														assign node32631 = (inp[5]) ? node32637 : node32632;
															assign node32632 = (inp[2]) ? node32634 : 4'b1011;
																assign node32634 = (inp[1]) ? 4'b1111 : 4'b1110;
															assign node32637 = (inp[2]) ? 4'b1010 : 4'b1110;
														assign node32640 = (inp[2]) ? node32646 : node32641;
															assign node32641 = (inp[5]) ? node32643 : 4'b1110;
																assign node32643 = (inp[1]) ? 4'b1110 : 4'b1010;
															assign node32646 = (inp[1]) ? 4'b1010 : node32647;
																assign node32647 = (inp[5]) ? 4'b1111 : 4'b1010;
												assign node32651 = (inp[1]) ? node32661 : node32652;
													assign node32652 = (inp[2]) ? 4'b1111 : node32653;
														assign node32653 = (inp[13]) ? node32657 : node32654;
															assign node32654 = (inp[15]) ? 4'b1010 : 4'b1011;
															assign node32657 = (inp[15]) ? 4'b1011 : 4'b1010;
													assign node32661 = (inp[2]) ? node32667 : node32662;
														assign node32662 = (inp[13]) ? 4'b1110 : node32663;
															assign node32663 = (inp[15]) ? 4'b1110 : 4'b1111;
														assign node32667 = (inp[13]) ? 4'b1010 : node32668;
															assign node32668 = (inp[15]) ? 4'b1010 : 4'b1011;
											assign node32672 = (inp[1]) ? node32706 : node32673;
												assign node32673 = (inp[2]) ? node32693 : node32674;
													assign node32674 = (inp[8]) ? node32688 : node32675;
														assign node32675 = (inp[13]) ? node32681 : node32676;
															assign node32676 = (inp[5]) ? node32678 : 4'b1011;
																assign node32678 = (inp[15]) ? 4'b1111 : 4'b1110;
															assign node32681 = (inp[15]) ? node32685 : node32682;
																assign node32682 = (inp[5]) ? 4'b1011 : 4'b1111;
																assign node32685 = (inp[5]) ? 4'b1010 : 4'b1110;
														assign node32688 = (inp[13]) ? 4'b1010 : node32689;
															assign node32689 = (inp[15]) ? 4'b1011 : 4'b1010;
													assign node32693 = (inp[8]) ? 4'b1110 : node32694;
														assign node32694 = (inp[5]) ? node32700 : node32695;
															assign node32695 = (inp[13]) ? node32697 : 4'b1110;
																assign node32697 = (inp[15]) ? 4'b1010 : 4'b1011;
															assign node32700 = (inp[13]) ? 4'b1110 : node32701;
																assign node32701 = (inp[15]) ? 4'b1011 : 4'b1010;
												assign node32706 = (inp[13]) ? node32722 : node32707;
													assign node32707 = (inp[15]) ? node32715 : node32708;
														assign node32708 = (inp[2]) ? node32712 : node32709;
															assign node32709 = (inp[8]) ? 4'b1110 : 4'b1011;
															assign node32712 = (inp[8]) ? 4'b1010 : 4'b1110;
														assign node32715 = (inp[2]) ? node32719 : node32716;
															assign node32716 = (inp[8]) ? 4'b1111 : 4'b1010;
															assign node32719 = (inp[8]) ? 4'b1011 : 4'b1111;
													assign node32722 = (inp[2]) ? 4'b1011 : 4'b1111;
										assign node32725 = (inp[0]) ? node32789 : node32726;
											assign node32726 = (inp[8]) ? node32768 : node32727;
												assign node32727 = (inp[15]) ? node32749 : node32728;
													assign node32728 = (inp[1]) ? node32742 : node32729;
														assign node32729 = (inp[2]) ? node32735 : node32730;
															assign node32730 = (inp[5]) ? node32732 : 4'b1011;
																assign node32732 = (inp[13]) ? 4'b1011 : 4'b1111;
															assign node32735 = (inp[13]) ? node32739 : node32736;
																assign node32736 = (inp[5]) ? 4'b1011 : 4'b1111;
																assign node32739 = (inp[5]) ? 4'b1111 : 4'b1011;
														assign node32742 = (inp[2]) ? node32746 : node32743;
															assign node32743 = (inp[13]) ? 4'b1111 : 4'b1011;
															assign node32746 = (inp[13]) ? 4'b1011 : 4'b1111;
													assign node32749 = (inp[13]) ? node32759 : node32750;
														assign node32750 = (inp[2]) ? node32756 : node32751;
															assign node32751 = (inp[1]) ? 4'b1010 : node32752;
																assign node32752 = (inp[5]) ? 4'b1111 : 4'b1010;
															assign node32756 = (inp[1]) ? 4'b1110 : 4'b1111;
														assign node32759 = (inp[5]) ? node32763 : node32760;
															assign node32760 = (inp[2]) ? 4'b1011 : 4'b1111;
															assign node32763 = (inp[2]) ? node32765 : 4'b1011;
																assign node32765 = (inp[1]) ? 4'b1011 : 4'b1110;
												assign node32768 = (inp[1]) ? node32778 : node32769;
													assign node32769 = (inp[2]) ? 4'b1110 : node32770;
														assign node32770 = (inp[15]) ? node32774 : node32771;
															assign node32771 = (inp[13]) ? 4'b1011 : 4'b1010;
															assign node32774 = (inp[13]) ? 4'b1010 : 4'b1011;
													assign node32778 = (inp[2]) ? node32784 : node32779;
														assign node32779 = (inp[15]) ? 4'b1111 : node32780;
															assign node32780 = (inp[13]) ? 4'b1111 : 4'b1110;
														assign node32784 = (inp[13]) ? 4'b1011 : node32785;
															assign node32785 = (inp[15]) ? 4'b1011 : 4'b1010;
											assign node32789 = (inp[1]) ? node32823 : node32790;
												assign node32790 = (inp[2]) ? node32810 : node32791;
													assign node32791 = (inp[8]) ? node32803 : node32792;
														assign node32792 = (inp[13]) ? node32798 : node32793;
															assign node32793 = (inp[5]) ? node32795 : 4'b1010;
																assign node32795 = (inp[15]) ? 4'b1110 : 4'b1111;
															assign node32798 = (inp[15]) ? 4'b1111 : node32799;
																assign node32799 = (inp[5]) ? 4'b1010 : 4'b1110;
														assign node32803 = (inp[13]) ? node32807 : node32804;
															assign node32804 = (inp[15]) ? 4'b1010 : 4'b1011;
															assign node32807 = (inp[15]) ? 4'b1011 : 4'b1010;
													assign node32810 = (inp[8]) ? 4'b1111 : node32811;
														assign node32811 = (inp[13]) ? node32817 : node32812;
															assign node32812 = (inp[5]) ? 4'b1010 : node32813;
																assign node32813 = (inp[15]) ? 4'b1110 : 4'b1111;
															assign node32817 = (inp[15]) ? node32819 : 4'b1010;
																assign node32819 = (inp[5]) ? 4'b1111 : 4'b1011;
												assign node32823 = (inp[2]) ? node32833 : node32824;
													assign node32824 = (inp[13]) ? 4'b1110 : node32825;
														assign node32825 = (inp[8]) ? node32829 : node32826;
															assign node32826 = (inp[15]) ? 4'b1011 : 4'b1010;
															assign node32829 = (inp[15]) ? 4'b1110 : 4'b1111;
													assign node32833 = (inp[13]) ? 4'b1010 : node32834;
														assign node32834 = (inp[15]) ? node32838 : node32835;
															assign node32835 = (inp[8]) ? 4'b1011 : 4'b1111;
															assign node32838 = (inp[8]) ? 4'b1010 : 4'b1110;
					assign node32842 = (inp[4]) ? node35142 : node32843;
						assign node32843 = (inp[8]) ? node34269 : node32844;
							assign node32844 = (inp[9]) ? node33490 : node32845;
								assign node32845 = (inp[13]) ? node33173 : node32846;
									assign node32846 = (inp[10]) ? node33010 : node32847;
										assign node32847 = (inp[5]) ? node32925 : node32848;
											assign node32848 = (inp[2]) ? node32890 : node32849;
												assign node32849 = (inp[1]) ? node32871 : node32850;
													assign node32850 = (inp[7]) ? node32862 : node32851;
														assign node32851 = (inp[15]) ? node32857 : node32852;
															assign node32852 = (inp[11]) ? node32854 : 4'b1010;
																assign node32854 = (inp[0]) ? 4'b1010 : 4'b1011;
															assign node32857 = (inp[11]) ? node32859 : 4'b1100;
																assign node32859 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node32862 = (inp[15]) ? node32866 : node32863;
															assign node32863 = (inp[11]) ? 4'b1100 : 4'b1101;
															assign node32866 = (inp[0]) ? 4'b1011 : node32867;
																assign node32867 = (inp[11]) ? 4'b1010 : 4'b1011;
													assign node32871 = (inp[7]) ? node32879 : node32872;
														assign node32872 = (inp[15]) ? 4'b1101 : node32873;
															assign node32873 = (inp[0]) ? 4'b1111 : node32874;
																assign node32874 = (inp[11]) ? 4'b1110 : 4'b1111;
														assign node32879 = (inp[15]) ? node32885 : node32880;
															assign node32880 = (inp[0]) ? node32882 : 4'b1101;
																assign node32882 = (inp[11]) ? 4'b1101 : 4'b1100;
															assign node32885 = (inp[0]) ? node32887 : 4'b1010;
																assign node32887 = (inp[11]) ? 4'b1010 : 4'b1011;
												assign node32890 = (inp[15]) ? node32906 : node32891;
													assign node32891 = (inp[7]) ? node32899 : node32892;
														assign node32892 = (inp[1]) ? node32896 : node32893;
															assign node32893 = (inp[11]) ? 4'b1110 : 4'b1111;
															assign node32896 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node32899 = (inp[1]) ? node32903 : node32900;
															assign node32900 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node32903 = (inp[0]) ? 4'b1001 : 4'b1000;
													assign node32906 = (inp[7]) ? node32914 : node32907;
														assign node32907 = (inp[0]) ? node32909 : 4'b1000;
															assign node32909 = (inp[11]) ? node32911 : 4'b1001;
																assign node32911 = (inp[1]) ? 4'b1000 : 4'b1001;
														assign node32914 = (inp[1]) ? node32920 : node32915;
															assign node32915 = (inp[11]) ? 4'b1111 : node32916;
																assign node32916 = (inp[0]) ? 4'b1110 : 4'b1111;
															assign node32920 = (inp[0]) ? 4'b1111 : node32921;
																assign node32921 = (inp[11]) ? 4'b1110 : 4'b1111;
											assign node32925 = (inp[2]) ? node32969 : node32926;
												assign node32926 = (inp[15]) ? node32946 : node32927;
													assign node32927 = (inp[7]) ? node32935 : node32928;
														assign node32928 = (inp[1]) ? node32932 : node32929;
															assign node32929 = (inp[11]) ? 4'b1010 : 4'b1011;
															assign node32932 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node32935 = (inp[1]) ? node32941 : node32936;
															assign node32936 = (inp[11]) ? node32938 : 4'b1000;
																assign node32938 = (inp[0]) ? 4'b1000 : 4'b1001;
															assign node32941 = (inp[0]) ? 4'b1101 : node32942;
																assign node32942 = (inp[11]) ? 4'b1100 : 4'b1101;
													assign node32946 = (inp[7]) ? node32958 : node32947;
														assign node32947 = (inp[1]) ? node32953 : node32948;
															assign node32948 = (inp[11]) ? 4'b1000 : node32949;
																assign node32949 = (inp[0]) ? 4'b1001 : 4'b1000;
															assign node32953 = (inp[11]) ? node32955 : 4'b1100;
																assign node32955 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node32958 = (inp[1]) ? node32964 : node32959;
															assign node32959 = (inp[11]) ? node32961 : 4'b1110;
																assign node32961 = (inp[0]) ? 4'b1110 : 4'b1111;
															assign node32964 = (inp[0]) ? 4'b1010 : node32965;
																assign node32965 = (inp[11]) ? 4'b1011 : 4'b1010;
												assign node32969 = (inp[15]) ? node32989 : node32970;
													assign node32970 = (inp[7]) ? node32980 : node32971;
														assign node32971 = (inp[1]) ? node32977 : node32972;
															assign node32972 = (inp[11]) ? node32974 : 4'b1111;
																assign node32974 = (inp[0]) ? 4'b1111 : 4'b1110;
															assign node32977 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node32980 = (inp[1]) ? node32986 : node32981;
															assign node32981 = (inp[0]) ? node32983 : 4'b1100;
																assign node32983 = (inp[11]) ? 4'b1100 : 4'b1101;
															assign node32986 = (inp[0]) ? 4'b1000 : 4'b1001;
													assign node32989 = (inp[7]) ? node32999 : node32990;
														assign node32990 = (inp[1]) ? node32994 : node32991;
															assign node32991 = (inp[11]) ? 4'b1100 : 4'b1101;
															assign node32994 = (inp[11]) ? node32996 : 4'b1001;
																assign node32996 = (inp[0]) ? 4'b1001 : 4'b1000;
														assign node32999 = (inp[1]) ? node33005 : node33000;
															assign node33000 = (inp[0]) ? 4'b1011 : node33001;
																assign node33001 = (inp[11]) ? 4'b1010 : 4'b1011;
															assign node33005 = (inp[11]) ? 4'b1110 : node33006;
																assign node33006 = (inp[0]) ? 4'b1111 : 4'b1110;
										assign node33010 = (inp[11]) ? node33078 : node33011;
											assign node33011 = (inp[15]) ? node33043 : node33012;
												assign node33012 = (inp[7]) ? node33028 : node33013;
													assign node33013 = (inp[2]) ? node33021 : node33014;
														assign node33014 = (inp[0]) ? 4'b1011 : node33015;
															assign node33015 = (inp[1]) ? node33017 : 4'b1011;
																assign node33017 = (inp[5]) ? 4'b1010 : 4'b1110;
														assign node33021 = (inp[1]) ? node33025 : node33022;
															assign node33022 = (inp[5]) ? 4'b1110 : 4'b1111;
															assign node33025 = (inp[5]) ? 4'b1111 : 4'b1011;
													assign node33028 = (inp[2]) ? node33036 : node33029;
														assign node33029 = (inp[1]) ? 4'b1100 : node33030;
															assign node33030 = (inp[5]) ? 4'b1001 : node33031;
																assign node33031 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node33036 = (inp[1]) ? 4'b1001 : node33037;
															assign node33037 = (inp[5]) ? 4'b1100 : node33038;
																assign node33038 = (inp[0]) ? 4'b1001 : 4'b1000;
												assign node33043 = (inp[7]) ? node33063 : node33044;
													assign node33044 = (inp[2]) ? node33054 : node33045;
														assign node33045 = (inp[5]) ? node33049 : node33046;
															assign node33046 = (inp[1]) ? 4'b1100 : 4'b1101;
															assign node33049 = (inp[1]) ? 4'b1101 : node33050;
																assign node33050 = (inp[0]) ? 4'b1000 : 4'b1001;
														assign node33054 = (inp[1]) ? node33058 : node33055;
															assign node33055 = (inp[5]) ? 4'b1100 : 4'b1000;
															assign node33058 = (inp[0]) ? 4'b1000 : node33059;
																assign node33059 = (inp[5]) ? 4'b1000 : 4'b1001;
													assign node33063 = (inp[2]) ? node33069 : node33064;
														assign node33064 = (inp[5]) ? node33066 : 4'b1010;
															assign node33066 = (inp[1]) ? 4'b1011 : 4'b1111;
														assign node33069 = (inp[1]) ? node33073 : node33070;
															assign node33070 = (inp[5]) ? 4'b1010 : 4'b1111;
															assign node33073 = (inp[0]) ? 4'b1110 : node33074;
																assign node33074 = (inp[5]) ? 4'b1111 : 4'b1110;
											assign node33078 = (inp[1]) ? node33126 : node33079;
												assign node33079 = (inp[2]) ? node33099 : node33080;
													assign node33080 = (inp[15]) ? node33086 : node33081;
														assign node33081 = (inp[7]) ? node33083 : 4'b1011;
															assign node33083 = (inp[5]) ? 4'b1001 : 4'b1101;
														assign node33086 = (inp[7]) ? node33092 : node33087;
															assign node33087 = (inp[5]) ? 4'b1001 : node33088;
																assign node33088 = (inp[0]) ? 4'b1101 : 4'b1100;
															assign node33092 = (inp[5]) ? node33096 : node33093;
																assign node33093 = (inp[0]) ? 4'b1010 : 4'b1011;
																assign node33096 = (inp[0]) ? 4'b1111 : 4'b1110;
													assign node33099 = (inp[0]) ? node33115 : node33100;
														assign node33100 = (inp[5]) ? node33108 : node33101;
															assign node33101 = (inp[7]) ? node33105 : node33102;
																assign node33102 = (inp[15]) ? 4'b1001 : 4'b1111;
																assign node33105 = (inp[15]) ? 4'b1110 : 4'b1000;
															assign node33108 = (inp[7]) ? node33112 : node33109;
																assign node33109 = (inp[15]) ? 4'b1101 : 4'b1111;
																assign node33112 = (inp[15]) ? 4'b1011 : 4'b1101;
														assign node33115 = (inp[7]) ? node33119 : node33116;
															assign node33116 = (inp[15]) ? 4'b1100 : 4'b1110;
															assign node33119 = (inp[15]) ? node33123 : node33120;
																assign node33120 = (inp[5]) ? 4'b1101 : 4'b1000;
																assign node33123 = (inp[5]) ? 4'b1010 : 4'b1110;
												assign node33126 = (inp[2]) ? node33150 : node33127;
													assign node33127 = (inp[15]) ? node33139 : node33128;
														assign node33128 = (inp[7]) ? node33134 : node33129;
															assign node33129 = (inp[5]) ? 4'b1010 : node33130;
																assign node33130 = (inp[0]) ? 4'b1110 : 4'b1111;
															assign node33134 = (inp[5]) ? node33136 : 4'b1100;
																assign node33136 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node33139 = (inp[7]) ? node33145 : node33140;
															assign node33140 = (inp[0]) ? node33142 : 4'b1100;
																assign node33142 = (inp[5]) ? 4'b1101 : 4'b1100;
															assign node33145 = (inp[0]) ? 4'b1011 : node33146;
																assign node33146 = (inp[5]) ? 4'b1010 : 4'b1011;
													assign node33150 = (inp[5]) ? node33160 : node33151;
														assign node33151 = (inp[7]) ? node33157 : node33152;
															assign node33152 = (inp[15]) ? 4'b1001 : node33153;
																assign node33153 = (inp[0]) ? 4'b1011 : 4'b1010;
															assign node33157 = (inp[15]) ? 4'b1111 : 4'b1001;
														assign node33160 = (inp[7]) ? node33168 : node33161;
															assign node33161 = (inp[15]) ? node33165 : node33162;
																assign node33162 = (inp[0]) ? 4'b1111 : 4'b1110;
																assign node33165 = (inp[0]) ? 4'b1000 : 4'b1001;
															assign node33168 = (inp[15]) ? 4'b1111 : node33169;
																assign node33169 = (inp[0]) ? 4'b1001 : 4'b1000;
									assign node33173 = (inp[7]) ? node33331 : node33174;
										assign node33174 = (inp[15]) ? node33258 : node33175;
											assign node33175 = (inp[2]) ? node33219 : node33176;
												assign node33176 = (inp[5]) ? node33198 : node33177;
													assign node33177 = (inp[1]) ? node33187 : node33178;
														assign node33178 = (inp[10]) ? node33184 : node33179;
															assign node33179 = (inp[0]) ? 4'b1110 : node33180;
																assign node33180 = (inp[11]) ? 4'b1111 : 4'b1110;
															assign node33184 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node33187 = (inp[10]) ? node33193 : node33188;
															assign node33188 = (inp[11]) ? 4'b1011 : node33189;
																assign node33189 = (inp[0]) ? 4'b1010 : 4'b1011;
															assign node33193 = (inp[11]) ? 4'b1010 : node33194;
																assign node33194 = (inp[0]) ? 4'b1011 : 4'b1010;
													assign node33198 = (inp[1]) ? node33210 : node33199;
														assign node33199 = (inp[10]) ? node33205 : node33200;
															assign node33200 = (inp[11]) ? 4'b1110 : node33201;
																assign node33201 = (inp[0]) ? 4'b1111 : 4'b1110;
															assign node33205 = (inp[11]) ? 4'b1111 : node33206;
																assign node33206 = (inp[0]) ? 4'b1110 : 4'b1111;
														assign node33210 = (inp[10]) ? node33216 : node33211;
															assign node33211 = (inp[11]) ? 4'b1111 : node33212;
																assign node33212 = (inp[0]) ? 4'b1110 : 4'b1111;
															assign node33216 = (inp[0]) ? 4'b1111 : 4'b1110;
												assign node33219 = (inp[1]) ? node33241 : node33220;
													assign node33220 = (inp[10]) ? node33230 : node33221;
														assign node33221 = (inp[11]) ? node33225 : node33222;
															assign node33222 = (inp[5]) ? 4'b1010 : 4'b1011;
															assign node33225 = (inp[5]) ? 4'b1011 : node33226;
																assign node33226 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node33230 = (inp[5]) ? node33236 : node33231;
															assign node33231 = (inp[11]) ? node33233 : 4'b1010;
																assign node33233 = (inp[0]) ? 4'b1010 : 4'b1011;
															assign node33236 = (inp[0]) ? node33238 : 4'b1010;
																assign node33238 = (inp[11]) ? 4'b1010 : 4'b1011;
													assign node33241 = (inp[5]) ? node33251 : node33242;
														assign node33242 = (inp[11]) ? node33244 : 4'b1110;
															assign node33244 = (inp[10]) ? node33248 : node33245;
																assign node33245 = (inp[0]) ? 4'b1110 : 4'b1111;
																assign node33248 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node33251 = (inp[10]) ? node33253 : 4'b1010;
															assign node33253 = (inp[0]) ? node33255 : 4'b1011;
																assign node33255 = (inp[11]) ? 4'b1011 : 4'b1010;
											assign node33258 = (inp[2]) ? node33288 : node33259;
												assign node33259 = (inp[10]) ? node33279 : node33260;
													assign node33260 = (inp[5]) ? node33270 : node33261;
														assign node33261 = (inp[11]) ? node33265 : node33262;
															assign node33262 = (inp[0]) ? 4'b1000 : 4'b1001;
															assign node33265 = (inp[1]) ? node33267 : 4'b1001;
																assign node33267 = (inp[0]) ? 4'b1001 : 4'b1000;
														assign node33270 = (inp[1]) ? node33276 : node33271;
															assign node33271 = (inp[11]) ? 4'b1101 : node33272;
																assign node33272 = (inp[0]) ? 4'b1100 : 4'b1101;
															assign node33276 = (inp[0]) ? 4'b1000 : 4'b1001;
													assign node33279 = (inp[1]) ? 4'b1000 : node33280;
														assign node33280 = (inp[5]) ? node33282 : 4'b1000;
															assign node33282 = (inp[11]) ? 4'b1100 : node33283;
																assign node33283 = (inp[0]) ? 4'b1101 : 4'b1100;
												assign node33288 = (inp[5]) ? node33310 : node33289;
													assign node33289 = (inp[11]) ? node33301 : node33290;
														assign node33290 = (inp[10]) ? node33296 : node33291;
															assign node33291 = (inp[0]) ? 4'b1100 : node33292;
																assign node33292 = (inp[1]) ? 4'b1101 : 4'b1100;
															assign node33296 = (inp[1]) ? node33298 : 4'b1101;
																assign node33298 = (inp[0]) ? 4'b1101 : 4'b1100;
														assign node33301 = (inp[10]) ? node33307 : node33302;
															assign node33302 = (inp[1]) ? 4'b1101 : node33303;
																assign node33303 = (inp[0]) ? 4'b1100 : 4'b1101;
															assign node33307 = (inp[1]) ? 4'b1100 : 4'b1101;
													assign node33310 = (inp[1]) ? node33322 : node33311;
														assign node33311 = (inp[10]) ? node33317 : node33312;
															assign node33312 = (inp[11]) ? 4'b1000 : node33313;
																assign node33313 = (inp[0]) ? 4'b1001 : 4'b1000;
															assign node33317 = (inp[0]) ? node33319 : 4'b1001;
																assign node33319 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node33322 = (inp[0]) ? 4'b1100 : node33323;
															assign node33323 = (inp[11]) ? node33327 : node33324;
																assign node33324 = (inp[10]) ? 4'b1101 : 4'b1100;
																assign node33327 = (inp[10]) ? 4'b1100 : 4'b1101;
										assign node33331 = (inp[15]) ? node33421 : node33332;
											assign node33332 = (inp[2]) ? node33372 : node33333;
												assign node33333 = (inp[1]) ? node33353 : node33334;
													assign node33334 = (inp[5]) ? node33342 : node33335;
														assign node33335 = (inp[10]) ? node33337 : 4'b1001;
															assign node33337 = (inp[11]) ? node33339 : 4'b1000;
																assign node33339 = (inp[0]) ? 4'b1000 : 4'b1001;
														assign node33342 = (inp[10]) ? node33348 : node33343;
															assign node33343 = (inp[0]) ? 4'b1100 : node33344;
																assign node33344 = (inp[11]) ? 4'b1101 : 4'b1100;
															assign node33348 = (inp[0]) ? 4'b1101 : node33349;
																assign node33349 = (inp[11]) ? 4'b1100 : 4'b1101;
													assign node33353 = (inp[10]) ? node33365 : node33354;
														assign node33354 = (inp[0]) ? node33360 : node33355;
															assign node33355 = (inp[5]) ? 4'b1001 : node33356;
																assign node33356 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node33360 = (inp[5]) ? node33362 : 4'b1000;
																assign node33362 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node33365 = (inp[11]) ? node33367 : 4'b1001;
															assign node33367 = (inp[5]) ? 4'b1000 : node33368;
																assign node33368 = (inp[0]) ? 4'b1001 : 4'b1000;
												assign node33372 = (inp[5]) ? node33402 : node33373;
													assign node33373 = (inp[11]) ? node33387 : node33374;
														assign node33374 = (inp[0]) ? node33380 : node33375;
															assign node33375 = (inp[1]) ? 4'b1100 : node33376;
																assign node33376 = (inp[10]) ? 4'b1100 : 4'b1101;
															assign node33380 = (inp[10]) ? node33384 : node33381;
																assign node33381 = (inp[1]) ? 4'b1101 : 4'b1100;
																assign node33384 = (inp[1]) ? 4'b1100 : 4'b1101;
														assign node33387 = (inp[0]) ? node33395 : node33388;
															assign node33388 = (inp[10]) ? node33392 : node33389;
																assign node33389 = (inp[1]) ? 4'b1100 : 4'b1101;
																assign node33392 = (inp[1]) ? 4'b1101 : 4'b1100;
															assign node33395 = (inp[1]) ? node33399 : node33396;
																assign node33396 = (inp[10]) ? 4'b1100 : 4'b1101;
																assign node33399 = (inp[10]) ? 4'b1101 : 4'b1100;
													assign node33402 = (inp[1]) ? node33412 : node33403;
														assign node33403 = (inp[11]) ? node33407 : node33404;
															assign node33404 = (inp[10]) ? 4'b1000 : 4'b1001;
															assign node33407 = (inp[10]) ? node33409 : 4'b1000;
																assign node33409 = (inp[0]) ? 4'b1000 : 4'b1001;
														assign node33412 = (inp[10]) ? node33418 : node33413;
															assign node33413 = (inp[0]) ? 4'b1100 : node33414;
																assign node33414 = (inp[11]) ? 4'b1101 : 4'b1100;
															assign node33418 = (inp[11]) ? 4'b1100 : 4'b1101;
											assign node33421 = (inp[2]) ? node33463 : node33422;
												assign node33422 = (inp[1]) ? node33442 : node33423;
													assign node33423 = (inp[5]) ? node33431 : node33424;
														assign node33424 = (inp[10]) ? node33426 : 4'b1110;
															assign node33426 = (inp[11]) ? node33428 : 4'b1111;
																assign node33428 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node33431 = (inp[10]) ? node33437 : node33432;
															assign node33432 = (inp[0]) ? node33434 : 4'b1011;
																assign node33434 = (inp[11]) ? 4'b1011 : 4'b1010;
															assign node33437 = (inp[11]) ? 4'b1010 : node33438;
																assign node33438 = (inp[0]) ? 4'b1011 : 4'b1010;
													assign node33442 = (inp[10]) ? node33452 : node33443;
														assign node33443 = (inp[5]) ? node33447 : node33444;
															assign node33444 = (inp[11]) ? 4'b1111 : 4'b1110;
															assign node33447 = (inp[0]) ? 4'b1111 : node33448;
																assign node33448 = (inp[11]) ? 4'b1110 : 4'b1111;
														assign node33452 = (inp[11]) ? node33458 : node33453;
															assign node33453 = (inp[0]) ? node33455 : 4'b1110;
																assign node33455 = (inp[5]) ? 4'b1110 : 4'b1111;
															assign node33458 = (inp[5]) ? node33460 : 4'b1110;
																assign node33460 = (inp[0]) ? 4'b1110 : 4'b1111;
												assign node33463 = (inp[1]) ? node33477 : node33464;
													assign node33464 = (inp[5]) ? node33470 : node33465;
														assign node33465 = (inp[10]) ? node33467 : 4'b1011;
															assign node33467 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node33470 = (inp[10]) ? node33474 : node33471;
															assign node33471 = (inp[11]) ? 4'b1111 : 4'b1110;
															assign node33474 = (inp[0]) ? 4'b1111 : 4'b1110;
													assign node33477 = (inp[10]) ? node33483 : node33478;
														assign node33478 = (inp[0]) ? 4'b1010 : node33479;
															assign node33479 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node33483 = (inp[0]) ? node33485 : 4'b1011;
															assign node33485 = (inp[11]) ? 4'b1011 : node33486;
																assign node33486 = (inp[5]) ? 4'b1011 : 4'b1010;
								assign node33490 = (inp[10]) ? node33874 : node33491;
									assign node33491 = (inp[13]) ? node33675 : node33492;
										assign node33492 = (inp[11]) ? node33578 : node33493;
											assign node33493 = (inp[2]) ? node33535 : node33494;
												assign node33494 = (inp[1]) ? node33514 : node33495;
													assign node33495 = (inp[15]) ? node33505 : node33496;
														assign node33496 = (inp[7]) ? node33502 : node33497;
															assign node33497 = (inp[0]) ? node33499 : 4'b1011;
																assign node33499 = (inp[5]) ? 4'b1010 : 4'b1011;
															assign node33502 = (inp[5]) ? 4'b1001 : 4'b1101;
														assign node33505 = (inp[7]) ? node33511 : node33506;
															assign node33506 = (inp[5]) ? node33508 : 4'b1101;
																assign node33508 = (inp[0]) ? 4'b1000 : 4'b1001;
															assign node33511 = (inp[5]) ? 4'b1111 : 4'b1010;
													assign node33514 = (inp[15]) ? node33526 : node33515;
														assign node33515 = (inp[7]) ? node33521 : node33516;
															assign node33516 = (inp[5]) ? node33518 : 4'b1110;
																assign node33518 = (inp[0]) ? 4'b1011 : 4'b1010;
															assign node33521 = (inp[0]) ? node33523 : 4'b1100;
																assign node33523 = (inp[5]) ? 4'b1100 : 4'b1101;
														assign node33526 = (inp[7]) ? node33530 : node33527;
															assign node33527 = (inp[5]) ? 4'b1101 : 4'b1100;
															assign node33530 = (inp[0]) ? node33532 : 4'b1011;
																assign node33532 = (inp[5]) ? 4'b1011 : 4'b1010;
												assign node33535 = (inp[1]) ? node33559 : node33536;
													assign node33536 = (inp[7]) ? node33546 : node33537;
														assign node33537 = (inp[15]) ? node33543 : node33538;
															assign node33538 = (inp[0]) ? 4'b1110 : node33539;
																assign node33539 = (inp[5]) ? 4'b1110 : 4'b1111;
															assign node33543 = (inp[5]) ? 4'b1100 : 4'b1000;
														assign node33546 = (inp[15]) ? node33554 : node33547;
															assign node33547 = (inp[5]) ? node33551 : node33548;
																assign node33548 = (inp[0]) ? 4'b1001 : 4'b1000;
																assign node33551 = (inp[0]) ? 4'b1100 : 4'b1101;
															assign node33554 = (inp[5]) ? 4'b1010 : node33555;
																assign node33555 = (inp[0]) ? 4'b1111 : 4'b1110;
													assign node33559 = (inp[0]) ? node33569 : node33560;
														assign node33560 = (inp[5]) ? node33566 : node33561;
															assign node33561 = (inp[15]) ? 4'b1001 : node33562;
																assign node33562 = (inp[7]) ? 4'b1001 : 4'b1011;
															assign node33566 = (inp[7]) ? 4'b1001 : 4'b1000;
														assign node33569 = (inp[15]) ? node33575 : node33570;
															assign node33570 = (inp[7]) ? node33572 : 4'b1111;
																assign node33572 = (inp[5]) ? 4'b1001 : 4'b1000;
															assign node33575 = (inp[7]) ? 4'b1110 : 4'b1000;
											assign node33578 = (inp[5]) ? node33628 : node33579;
												assign node33579 = (inp[0]) ? node33601 : node33580;
													assign node33580 = (inp[2]) ? node33592 : node33581;
														assign node33581 = (inp[7]) ? node33587 : node33582;
															assign node33582 = (inp[15]) ? 4'b1100 : node33583;
																assign node33583 = (inp[1]) ? 4'b1111 : 4'b1010;
															assign node33587 = (inp[15]) ? 4'b1011 : node33588;
																assign node33588 = (inp[1]) ? 4'b1100 : 4'b1101;
														assign node33592 = (inp[1]) ? node33596 : node33593;
															assign node33593 = (inp[15]) ? 4'b1110 : 4'b1111;
															assign node33596 = (inp[7]) ? 4'b1111 : node33597;
																assign node33597 = (inp[15]) ? 4'b1001 : 4'b1010;
													assign node33601 = (inp[2]) ? node33615 : node33602;
														assign node33602 = (inp[1]) ? node33608 : node33603;
															assign node33603 = (inp[7]) ? 4'b1010 : node33604;
																assign node33604 = (inp[15]) ? 4'b1101 : 4'b1011;
															assign node33608 = (inp[15]) ? node33612 : node33609;
																assign node33609 = (inp[7]) ? 4'b1100 : 4'b1110;
																assign node33612 = (inp[7]) ? 4'b1011 : 4'b1100;
														assign node33615 = (inp[1]) ? node33621 : node33616;
															assign node33616 = (inp[7]) ? 4'b1000 : node33617;
																assign node33617 = (inp[15]) ? 4'b1000 : 4'b1111;
															assign node33621 = (inp[15]) ? node33625 : node33622;
																assign node33622 = (inp[7]) ? 4'b1001 : 4'b1011;
																assign node33625 = (inp[7]) ? 4'b1110 : 4'b1001;
												assign node33628 = (inp[2]) ? node33650 : node33629;
													assign node33629 = (inp[7]) ? node33637 : node33630;
														assign node33630 = (inp[15]) ? node33634 : node33631;
															assign node33631 = (inp[1]) ? 4'b1010 : 4'b1011;
															assign node33634 = (inp[1]) ? 4'b1101 : 4'b1001;
														assign node33637 = (inp[15]) ? node33645 : node33638;
															assign node33638 = (inp[1]) ? node33642 : node33639;
																assign node33639 = (inp[0]) ? 4'b1001 : 4'b1000;
																assign node33642 = (inp[0]) ? 4'b1100 : 4'b1101;
															assign node33645 = (inp[1]) ? 4'b1011 : node33646;
																assign node33646 = (inp[0]) ? 4'b1111 : 4'b1110;
													assign node33650 = (inp[15]) ? node33664 : node33651;
														assign node33651 = (inp[7]) ? node33659 : node33652;
															assign node33652 = (inp[0]) ? node33656 : node33653;
																assign node33653 = (inp[1]) ? 4'b1110 : 4'b1111;
																assign node33656 = (inp[1]) ? 4'b1111 : 4'b1110;
															assign node33659 = (inp[1]) ? node33661 : 4'b1101;
																assign node33661 = (inp[0]) ? 4'b1001 : 4'b1000;
														assign node33664 = (inp[7]) ? node33670 : node33665;
															assign node33665 = (inp[1]) ? node33667 : 4'b1101;
																assign node33667 = (inp[0]) ? 4'b1000 : 4'b1001;
															assign node33670 = (inp[1]) ? 4'b1111 : node33671;
																assign node33671 = (inp[0]) ? 4'b1010 : 4'b1011;
										assign node33675 = (inp[11]) ? node33785 : node33676;
											assign node33676 = (inp[0]) ? node33728 : node33677;
												assign node33677 = (inp[2]) ? node33703 : node33678;
													assign node33678 = (inp[1]) ? node33692 : node33679;
														assign node33679 = (inp[5]) ? node33687 : node33680;
															assign node33680 = (inp[15]) ? node33684 : node33681;
																assign node33681 = (inp[7]) ? 4'b1000 : 4'b1111;
																assign node33684 = (inp[7]) ? 4'b1111 : 4'b1000;
															assign node33687 = (inp[15]) ? 4'b1100 : node33688;
																assign node33688 = (inp[7]) ? 4'b1101 : 4'b1111;
														assign node33692 = (inp[7]) ? node33698 : node33693;
															assign node33693 = (inp[15]) ? 4'b1000 : node33694;
																assign node33694 = (inp[5]) ? 4'b1110 : 4'b1010;
															assign node33698 = (inp[15]) ? 4'b1110 : node33699;
																assign node33699 = (inp[5]) ? 4'b1000 : 4'b1001;
													assign node33703 = (inp[1]) ? node33717 : node33704;
														assign node33704 = (inp[15]) ? node33710 : node33705;
															assign node33705 = (inp[7]) ? node33707 : 4'b1010;
																assign node33707 = (inp[5]) ? 4'b1000 : 4'b1100;
															assign node33710 = (inp[7]) ? node33714 : node33711;
																assign node33711 = (inp[5]) ? 4'b1001 : 4'b1101;
																assign node33714 = (inp[5]) ? 4'b1111 : 4'b1010;
														assign node33717 = (inp[5]) ? node33721 : node33718;
															assign node33718 = (inp[7]) ? 4'b1101 : 4'b1111;
															assign node33721 = (inp[7]) ? node33725 : node33722;
																assign node33722 = (inp[15]) ? 4'b1101 : 4'b1011;
																assign node33725 = (inp[15]) ? 4'b1011 : 4'b1101;
												assign node33728 = (inp[2]) ? node33758 : node33729;
													assign node33729 = (inp[1]) ? node33745 : node33730;
														assign node33730 = (inp[15]) ? node33738 : node33731;
															assign node33731 = (inp[7]) ? node33735 : node33732;
																assign node33732 = (inp[5]) ? 4'b1110 : 4'b1111;
																assign node33735 = (inp[5]) ? 4'b1101 : 4'b1000;
															assign node33738 = (inp[7]) ? node33742 : node33739;
																assign node33739 = (inp[5]) ? 4'b1101 : 4'b1001;
																assign node33742 = (inp[5]) ? 4'b1011 : 4'b1111;
														assign node33745 = (inp[15]) ? node33751 : node33746;
															assign node33746 = (inp[7]) ? 4'b1001 : node33747;
																assign node33747 = (inp[5]) ? 4'b1111 : 4'b1011;
															assign node33751 = (inp[7]) ? node33755 : node33752;
																assign node33752 = (inp[5]) ? 4'b1001 : 4'b1000;
																assign node33755 = (inp[5]) ? 4'b1110 : 4'b1111;
													assign node33758 = (inp[5]) ? node33770 : node33759;
														assign node33759 = (inp[15]) ? node33767 : node33760;
															assign node33760 = (inp[7]) ? node33764 : node33761;
																assign node33761 = (inp[1]) ? 4'b1111 : 4'b1010;
																assign node33764 = (inp[1]) ? 4'b1100 : 4'b1101;
															assign node33767 = (inp[7]) ? 4'b1010 : 4'b1101;
														assign node33770 = (inp[1]) ? node33778 : node33771;
															assign node33771 = (inp[15]) ? node33775 : node33772;
																assign node33772 = (inp[7]) ? 4'b1000 : 4'b1011;
																assign node33775 = (inp[7]) ? 4'b1111 : 4'b1000;
															assign node33778 = (inp[7]) ? node33782 : node33779;
																assign node33779 = (inp[15]) ? 4'b1101 : 4'b1010;
																assign node33782 = (inp[15]) ? 4'b1011 : 4'b1101;
											assign node33785 = (inp[2]) ? node33829 : node33786;
												assign node33786 = (inp[1]) ? node33810 : node33787;
													assign node33787 = (inp[15]) ? node33801 : node33788;
														assign node33788 = (inp[7]) ? node33794 : node33789;
															assign node33789 = (inp[5]) ? 4'b1111 : node33790;
																assign node33790 = (inp[0]) ? 4'b1111 : 4'b1110;
															assign node33794 = (inp[5]) ? node33798 : node33795;
																assign node33795 = (inp[0]) ? 4'b1000 : 4'b1001;
																assign node33798 = (inp[0]) ? 4'b1101 : 4'b1100;
														assign node33801 = (inp[7]) ? node33805 : node33802;
															assign node33802 = (inp[5]) ? 4'b1100 : 4'b1000;
															assign node33805 = (inp[5]) ? 4'b1010 : node33806;
																assign node33806 = (inp[0]) ? 4'b1111 : 4'b1110;
													assign node33810 = (inp[15]) ? node33820 : node33811;
														assign node33811 = (inp[7]) ? node33815 : node33812;
															assign node33812 = (inp[5]) ? 4'b1110 : 4'b1010;
															assign node33815 = (inp[5]) ? 4'b1000 : node33816;
																assign node33816 = (inp[0]) ? 4'b1001 : 4'b1000;
														assign node33820 = (inp[7]) ? node33826 : node33821;
															assign node33821 = (inp[5]) ? 4'b1000 : node33822;
																assign node33822 = (inp[0]) ? 4'b1000 : 4'b1001;
															assign node33826 = (inp[5]) ? 4'b1111 : 4'b1110;
												assign node33829 = (inp[1]) ? node33855 : node33830;
													assign node33830 = (inp[15]) ? node33842 : node33831;
														assign node33831 = (inp[7]) ? node33837 : node33832;
															assign node33832 = (inp[5]) ? 4'b1010 : node33833;
																assign node33833 = (inp[0]) ? 4'b1010 : 4'b1011;
															assign node33837 = (inp[0]) ? node33839 : 4'b1001;
																assign node33839 = (inp[5]) ? 4'b1000 : 4'b1100;
														assign node33842 = (inp[7]) ? node33848 : node33843;
															assign node33843 = (inp[5]) ? 4'b1001 : node33844;
																assign node33844 = (inp[0]) ? 4'b1101 : 4'b1100;
															assign node33848 = (inp[5]) ? node33852 : node33849;
																assign node33849 = (inp[0]) ? 4'b1010 : 4'b1011;
																assign node33852 = (inp[0]) ? 4'b1111 : 4'b1110;
													assign node33855 = (inp[7]) ? node33867 : node33856;
														assign node33856 = (inp[15]) ? node33862 : node33857;
															assign node33857 = (inp[0]) ? node33859 : 4'b1110;
																assign node33859 = (inp[5]) ? 4'b1011 : 4'b1111;
															assign node33862 = (inp[0]) ? node33864 : 4'b1100;
																assign node33864 = (inp[5]) ? 4'b1101 : 4'b1100;
														assign node33867 = (inp[15]) ? node33869 : 4'b1101;
															assign node33869 = (inp[5]) ? node33871 : 4'b1011;
																assign node33871 = (inp[0]) ? 4'b1011 : 4'b1010;
									assign node33874 = (inp[13]) ? node34084 : node33875;
										assign node33875 = (inp[11]) ? node33983 : node33876;
											assign node33876 = (inp[0]) ? node33936 : node33877;
												assign node33877 = (inp[5]) ? node33905 : node33878;
													assign node33878 = (inp[2]) ? node33894 : node33879;
														assign node33879 = (inp[1]) ? node33887 : node33880;
															assign node33880 = (inp[7]) ? node33884 : node33881;
																assign node33881 = (inp[15]) ? 4'b1100 : 4'b1010;
																assign node33884 = (inp[15]) ? 4'b1011 : 4'b1100;
															assign node33887 = (inp[7]) ? node33891 : node33888;
																assign node33888 = (inp[15]) ? 4'b1101 : 4'b1111;
																assign node33891 = (inp[15]) ? 4'b1010 : 4'b1101;
														assign node33894 = (inp[1]) ? node33900 : node33895;
															assign node33895 = (inp[7]) ? node33897 : 4'b1001;
																assign node33897 = (inp[15]) ? 4'b1111 : 4'b1001;
															assign node33900 = (inp[7]) ? 4'b1000 : node33901;
																assign node33901 = (inp[15]) ? 4'b1000 : 4'b1010;
													assign node33905 = (inp[2]) ? node33921 : node33906;
														assign node33906 = (inp[15]) ? node33914 : node33907;
															assign node33907 = (inp[1]) ? node33911 : node33908;
																assign node33908 = (inp[7]) ? 4'b1000 : 4'b1010;
																assign node33911 = (inp[7]) ? 4'b1101 : 4'b1011;
															assign node33914 = (inp[7]) ? node33918 : node33915;
																assign node33915 = (inp[1]) ? 4'b1100 : 4'b1000;
																assign node33918 = (inp[1]) ? 4'b1010 : 4'b1110;
														assign node33921 = (inp[1]) ? node33929 : node33922;
															assign node33922 = (inp[7]) ? node33926 : node33923;
																assign node33923 = (inp[15]) ? 4'b1101 : 4'b1111;
																assign node33926 = (inp[15]) ? 4'b1011 : 4'b1100;
															assign node33929 = (inp[7]) ? node33933 : node33930;
																assign node33930 = (inp[15]) ? 4'b1001 : 4'b1110;
																assign node33933 = (inp[15]) ? 4'b1110 : 4'b1000;
												assign node33936 = (inp[5]) ? node33958 : node33937;
													assign node33937 = (inp[2]) ? node33945 : node33938;
														assign node33938 = (inp[15]) ? 4'b1011 : node33939;
															assign node33939 = (inp[7]) ? 4'b1101 : node33940;
																assign node33940 = (inp[1]) ? 4'b1111 : 4'b1010;
														assign node33945 = (inp[15]) ? node33953 : node33946;
															assign node33946 = (inp[7]) ? node33950 : node33947;
																assign node33947 = (inp[1]) ? 4'b1010 : 4'b1111;
																assign node33950 = (inp[1]) ? 4'b1001 : 4'b1000;
															assign node33953 = (inp[7]) ? node33955 : 4'b1001;
																assign node33955 = (inp[1]) ? 4'b1111 : 4'b1110;
													assign node33958 = (inp[2]) ? node33970 : node33959;
														assign node33959 = (inp[7]) ? node33965 : node33960;
															assign node33960 = (inp[1]) ? 4'b1100 : node33961;
																assign node33961 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node33965 = (inp[15]) ? node33967 : 4'b1000;
																assign node33967 = (inp[1]) ? 4'b1010 : 4'b1110;
														assign node33970 = (inp[1]) ? node33976 : node33971;
															assign node33971 = (inp[15]) ? 4'b1101 : node33972;
																assign node33972 = (inp[7]) ? 4'b1101 : 4'b1111;
															assign node33976 = (inp[15]) ? node33980 : node33977;
																assign node33977 = (inp[7]) ? 4'b1000 : 4'b1110;
																assign node33980 = (inp[7]) ? 4'b1111 : 4'b1001;
											assign node33983 = (inp[1]) ? node34037 : node33984;
												assign node33984 = (inp[2]) ? node34014 : node33985;
													assign node33985 = (inp[0]) ? node34001 : node33986;
														assign node33986 = (inp[7]) ? node33994 : node33987;
															assign node33987 = (inp[15]) ? node33991 : node33988;
																assign node33988 = (inp[5]) ? 4'b1010 : 4'b1011;
																assign node33991 = (inp[5]) ? 4'b1000 : 4'b1101;
															assign node33994 = (inp[5]) ? node33998 : node33995;
																assign node33995 = (inp[15]) ? 4'b1010 : 4'b1100;
																assign node33998 = (inp[15]) ? 4'b1111 : 4'b1001;
														assign node34001 = (inp[7]) ? node34007 : node34002;
															assign node34002 = (inp[15]) ? node34004 : 4'b1010;
																assign node34004 = (inp[5]) ? 4'b1000 : 4'b1100;
															assign node34007 = (inp[15]) ? node34011 : node34008;
																assign node34008 = (inp[5]) ? 4'b1000 : 4'b1100;
																assign node34011 = (inp[5]) ? 4'b1110 : 4'b1011;
													assign node34014 = (inp[0]) ? node34024 : node34015;
														assign node34015 = (inp[15]) ? node34019 : node34016;
															assign node34016 = (inp[7]) ? 4'b1100 : 4'b1110;
															assign node34019 = (inp[7]) ? 4'b1010 : node34020;
																assign node34020 = (inp[5]) ? 4'b1100 : 4'b1000;
														assign node34024 = (inp[15]) ? node34032 : node34025;
															assign node34025 = (inp[7]) ? node34029 : node34026;
																assign node34026 = (inp[5]) ? 4'b1111 : 4'b1110;
																assign node34029 = (inp[5]) ? 4'b1100 : 4'b1001;
															assign node34032 = (inp[7]) ? node34034 : 4'b1101;
																assign node34034 = (inp[5]) ? 4'b1011 : 4'b1111;
												assign node34037 = (inp[2]) ? node34059 : node34038;
													assign node34038 = (inp[15]) ? node34050 : node34039;
														assign node34039 = (inp[7]) ? node34045 : node34040;
															assign node34040 = (inp[5]) ? 4'b1011 : node34041;
																assign node34041 = (inp[0]) ? 4'b1111 : 4'b1110;
															assign node34045 = (inp[0]) ? 4'b1101 : node34046;
																assign node34046 = (inp[5]) ? 4'b1100 : 4'b1101;
														assign node34050 = (inp[7]) ? node34054 : node34051;
															assign node34051 = (inp[5]) ? 4'b1100 : 4'b1101;
															assign node34054 = (inp[5]) ? node34056 : 4'b1010;
																assign node34056 = (inp[0]) ? 4'b1010 : 4'b1011;
													assign node34059 = (inp[5]) ? node34071 : node34060;
														assign node34060 = (inp[7]) ? node34066 : node34061;
															assign node34061 = (inp[15]) ? 4'b1000 : node34062;
																assign node34062 = (inp[0]) ? 4'b1010 : 4'b1011;
															assign node34066 = (inp[15]) ? node34068 : 4'b1000;
																assign node34068 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node34071 = (inp[15]) ? node34079 : node34072;
															assign node34072 = (inp[7]) ? node34076 : node34073;
																assign node34073 = (inp[0]) ? 4'b1110 : 4'b1111;
																assign node34076 = (inp[0]) ? 4'b1000 : 4'b1001;
															assign node34079 = (inp[7]) ? 4'b1110 : node34080;
																assign node34080 = (inp[0]) ? 4'b1001 : 4'b1000;
										assign node34084 = (inp[11]) ? node34184 : node34085;
											assign node34085 = (inp[0]) ? node34133 : node34086;
												assign node34086 = (inp[2]) ? node34106 : node34087;
													assign node34087 = (inp[15]) ? node34097 : node34088;
														assign node34088 = (inp[1]) ? node34092 : node34089;
															assign node34089 = (inp[7]) ? 4'b1100 : 4'b1110;
															assign node34092 = (inp[7]) ? node34094 : 4'b1011;
																assign node34094 = (inp[5]) ? 4'b1001 : 4'b1000;
														assign node34097 = (inp[7]) ? node34103 : node34098;
															assign node34098 = (inp[1]) ? 4'b1001 : node34099;
																assign node34099 = (inp[5]) ? 4'b1101 : 4'b1001;
															assign node34103 = (inp[1]) ? 4'b1111 : 4'b1011;
													assign node34106 = (inp[1]) ? node34120 : node34107;
														assign node34107 = (inp[15]) ? node34113 : node34108;
															assign node34108 = (inp[7]) ? node34110 : 4'b1011;
																assign node34110 = (inp[5]) ? 4'b1001 : 4'b1101;
															assign node34113 = (inp[7]) ? node34117 : node34114;
																assign node34114 = (inp[5]) ? 4'b1000 : 4'b1100;
																assign node34117 = (inp[5]) ? 4'b1110 : 4'b1011;
														assign node34120 = (inp[5]) ? node34128 : node34121;
															assign node34121 = (inp[15]) ? node34125 : node34122;
																assign node34122 = (inp[7]) ? 4'b1100 : 4'b1110;
																assign node34125 = (inp[7]) ? 4'b1010 : 4'b1101;
															assign node34128 = (inp[15]) ? node34130 : 4'b1010;
																assign node34130 = (inp[7]) ? 4'b1010 : 4'b1100;
												assign node34133 = (inp[2]) ? node34159 : node34134;
													assign node34134 = (inp[5]) ? node34148 : node34135;
														assign node34135 = (inp[1]) ? node34141 : node34136;
															assign node34136 = (inp[7]) ? 4'b1110 : node34137;
																assign node34137 = (inp[15]) ? 4'b1000 : 4'b1110;
															assign node34141 = (inp[15]) ? node34145 : node34142;
																assign node34142 = (inp[7]) ? 4'b1000 : 4'b1010;
																assign node34145 = (inp[7]) ? 4'b1110 : 4'b1001;
														assign node34148 = (inp[7]) ? node34152 : node34149;
															assign node34149 = (inp[1]) ? 4'b1110 : 4'b1111;
															assign node34152 = (inp[15]) ? node34156 : node34153;
																assign node34153 = (inp[1]) ? 4'b1000 : 4'b1100;
																assign node34156 = (inp[1]) ? 4'b1111 : 4'b1010;
													assign node34159 = (inp[5]) ? node34169 : node34160;
														assign node34160 = (inp[7]) ? node34166 : node34161;
															assign node34161 = (inp[15]) ? 4'b1100 : node34162;
																assign node34162 = (inp[1]) ? 4'b1110 : 4'b1011;
															assign node34166 = (inp[15]) ? 4'b1011 : 4'b1101;
														assign node34169 = (inp[7]) ? node34177 : node34170;
															assign node34170 = (inp[15]) ? node34174 : node34171;
																assign node34171 = (inp[1]) ? 4'b1011 : 4'b1010;
																assign node34174 = (inp[1]) ? 4'b1100 : 4'b1001;
															assign node34177 = (inp[15]) ? node34181 : node34178;
																assign node34178 = (inp[1]) ? 4'b1100 : 4'b1001;
																assign node34181 = (inp[1]) ? 4'b1010 : 4'b1110;
											assign node34184 = (inp[2]) ? node34226 : node34185;
												assign node34185 = (inp[1]) ? node34205 : node34186;
													assign node34186 = (inp[15]) ? node34196 : node34187;
														assign node34187 = (inp[7]) ? node34193 : node34188;
															assign node34188 = (inp[5]) ? 4'b1110 : node34189;
																assign node34189 = (inp[0]) ? 4'b1110 : 4'b1111;
															assign node34193 = (inp[0]) ? 4'b1001 : 4'b1000;
														assign node34196 = (inp[7]) ? node34200 : node34197;
															assign node34197 = (inp[5]) ? 4'b1101 : 4'b1001;
															assign node34200 = (inp[5]) ? 4'b1011 : node34201;
																assign node34201 = (inp[0]) ? 4'b1110 : 4'b1111;
													assign node34205 = (inp[7]) ? node34215 : node34206;
														assign node34206 = (inp[15]) ? node34210 : node34207;
															assign node34207 = (inp[5]) ? 4'b1111 : 4'b1011;
															assign node34210 = (inp[0]) ? 4'b1001 : node34211;
																assign node34211 = (inp[5]) ? 4'b1001 : 4'b1000;
														assign node34215 = (inp[15]) ? node34221 : node34216;
															assign node34216 = (inp[5]) ? 4'b1001 : node34217;
																assign node34217 = (inp[0]) ? 4'b1000 : 4'b1001;
															assign node34221 = (inp[0]) ? 4'b1111 : node34222;
																assign node34222 = (inp[5]) ? 4'b1110 : 4'b1111;
												assign node34226 = (inp[5]) ? node34246 : node34227;
													assign node34227 = (inp[15]) ? node34237 : node34228;
														assign node34228 = (inp[7]) ? node34234 : node34229;
															assign node34229 = (inp[1]) ? node34231 : 4'b1011;
																assign node34231 = (inp[0]) ? 4'b1110 : 4'b1111;
															assign node34234 = (inp[1]) ? 4'b1100 : 4'b1101;
														assign node34237 = (inp[7]) ? node34241 : node34238;
															assign node34238 = (inp[1]) ? 4'b1101 : 4'b1100;
															assign node34241 = (inp[0]) ? node34243 : 4'b1010;
																assign node34243 = (inp[1]) ? 4'b1010 : 4'b1011;
													assign node34246 = (inp[0]) ? node34258 : node34247;
														assign node34247 = (inp[7]) ? node34253 : node34248;
															assign node34248 = (inp[15]) ? node34250 : 4'b1010;
																assign node34250 = (inp[1]) ? 4'b1101 : 4'b1000;
															assign node34253 = (inp[15]) ? node34255 : 4'b1101;
																assign node34255 = (inp[1]) ? 4'b1011 : 4'b1111;
														assign node34258 = (inp[15]) ? node34264 : node34259;
															assign node34259 = (inp[1]) ? 4'b1010 : node34260;
																assign node34260 = (inp[7]) ? 4'b1001 : 4'b1011;
															assign node34264 = (inp[7]) ? node34266 : 4'b1000;
																assign node34266 = (inp[1]) ? 4'b1010 : 4'b1110;
							assign node34269 = (inp[11]) ? node34799 : node34270;
								assign node34270 = (inp[5]) ? node34522 : node34271;
									assign node34271 = (inp[10]) ? node34403 : node34272;
										assign node34272 = (inp[0]) ? node34324 : node34273;
											assign node34273 = (inp[7]) ? node34301 : node34274;
												assign node34274 = (inp[2]) ? node34290 : node34275;
													assign node34275 = (inp[13]) ? node34283 : node34276;
														assign node34276 = (inp[15]) ? node34280 : node34277;
															assign node34277 = (inp[1]) ? 4'b1111 : 4'b1010;
															assign node34280 = (inp[1]) ? 4'b1010 : 4'b1110;
														assign node34283 = (inp[1]) ? node34287 : node34284;
															assign node34284 = (inp[15]) ? 4'b1111 : 4'b1010;
															assign node34287 = (inp[15]) ? 4'b1011 : 4'b1111;
													assign node34290 = (inp[1]) ? node34298 : node34291;
														assign node34291 = (inp[15]) ? node34295 : node34292;
															assign node34292 = (inp[13]) ? 4'b1111 : 4'b1110;
															assign node34295 = (inp[13]) ? 4'b1010 : 4'b1011;
														assign node34298 = (inp[15]) ? 4'b1110 : 4'b1010;
												assign node34301 = (inp[2]) ? node34313 : node34302;
													assign node34302 = (inp[1]) ? node34310 : node34303;
														assign node34303 = (inp[15]) ? node34307 : node34304;
															assign node34304 = (inp[13]) ? 4'b1111 : 4'b1110;
															assign node34307 = (inp[13]) ? 4'b1010 : 4'b1011;
														assign node34310 = (inp[15]) ? 4'b1110 : 4'b1010;
													assign node34313 = (inp[15]) ? node34321 : node34314;
														assign node34314 = (inp[1]) ? node34318 : node34315;
															assign node34315 = (inp[13]) ? 4'b1010 : 4'b1011;
															assign node34318 = (inp[13]) ? 4'b1111 : 4'b1110;
														assign node34321 = (inp[1]) ? 4'b1011 : 4'b1111;
											assign node34324 = (inp[13]) ? node34364 : node34325;
												assign node34325 = (inp[2]) ? node34349 : node34326;
													assign node34326 = (inp[9]) ? node34336 : node34327;
														assign node34327 = (inp[1]) ? node34329 : 4'b1111;
															assign node34329 = (inp[15]) ? node34333 : node34330;
																assign node34330 = (inp[7]) ? 4'b1011 : 4'b1110;
																assign node34333 = (inp[7]) ? 4'b1111 : 4'b1011;
														assign node34336 = (inp[1]) ? node34342 : node34337;
															assign node34337 = (inp[15]) ? 4'b1010 : node34338;
																assign node34338 = (inp[7]) ? 4'b1111 : 4'b1011;
															assign node34342 = (inp[15]) ? node34346 : node34343;
																assign node34343 = (inp[7]) ? 4'b1011 : 4'b1110;
																assign node34346 = (inp[7]) ? 4'b1111 : 4'b1011;
													assign node34349 = (inp[7]) ? node34357 : node34350;
														assign node34350 = (inp[1]) ? node34354 : node34351;
															assign node34351 = (inp[15]) ? 4'b1010 : 4'b1111;
															assign node34354 = (inp[15]) ? 4'b1111 : 4'b1011;
														assign node34357 = (inp[15]) ? node34361 : node34358;
															assign node34358 = (inp[1]) ? 4'b1111 : 4'b1010;
															assign node34361 = (inp[1]) ? 4'b1010 : 4'b1110;
												assign node34364 = (inp[15]) ? node34382 : node34365;
													assign node34365 = (inp[7]) ? node34373 : node34366;
														assign node34366 = (inp[2]) ? node34370 : node34367;
															assign node34367 = (inp[1]) ? 4'b1110 : 4'b1011;
															assign node34370 = (inp[1]) ? 4'b1011 : 4'b1110;
														assign node34373 = (inp[9]) ? node34375 : 4'b1110;
															assign node34375 = (inp[2]) ? node34379 : node34376;
																assign node34376 = (inp[1]) ? 4'b1011 : 4'b1110;
																assign node34379 = (inp[1]) ? 4'b1110 : 4'b1011;
													assign node34382 = (inp[1]) ? node34390 : node34383;
														assign node34383 = (inp[2]) ? node34387 : node34384;
															assign node34384 = (inp[7]) ? 4'b1011 : 4'b1110;
															assign node34387 = (inp[7]) ? 4'b1110 : 4'b1011;
														assign node34390 = (inp[9]) ? node34396 : node34391;
															assign node34391 = (inp[7]) ? 4'b1010 : node34392;
																assign node34392 = (inp[2]) ? 4'b1111 : 4'b1010;
															assign node34396 = (inp[2]) ? node34400 : node34397;
																assign node34397 = (inp[7]) ? 4'b1111 : 4'b1010;
																assign node34400 = (inp[7]) ? 4'b1010 : 4'b1111;
										assign node34403 = (inp[0]) ? node34475 : node34404;
											assign node34404 = (inp[15]) ? node34450 : node34405;
												assign node34405 = (inp[13]) ? node34421 : node34406;
													assign node34406 = (inp[1]) ? node34414 : node34407;
														assign node34407 = (inp[7]) ? node34411 : node34408;
															assign node34408 = (inp[2]) ? 4'b1111 : 4'b1011;
															assign node34411 = (inp[2]) ? 4'b1010 : 4'b1111;
														assign node34414 = (inp[2]) ? node34418 : node34415;
															assign node34415 = (inp[7]) ? 4'b1011 : 4'b1110;
															assign node34418 = (inp[7]) ? 4'b1111 : 4'b1011;
													assign node34421 = (inp[7]) ? node34437 : node34422;
														assign node34422 = (inp[9]) ? node34430 : node34423;
															assign node34423 = (inp[1]) ? node34427 : node34424;
																assign node34424 = (inp[2]) ? 4'b1110 : 4'b1011;
																assign node34427 = (inp[2]) ? 4'b1011 : 4'b1110;
															assign node34430 = (inp[1]) ? node34434 : node34431;
																assign node34431 = (inp[2]) ? 4'b1110 : 4'b1011;
																assign node34434 = (inp[2]) ? 4'b1011 : 4'b1110;
														assign node34437 = (inp[9]) ? node34445 : node34438;
															assign node34438 = (inp[2]) ? node34442 : node34439;
																assign node34439 = (inp[1]) ? 4'b1011 : 4'b1110;
																assign node34442 = (inp[1]) ? 4'b1110 : 4'b1011;
															assign node34445 = (inp[1]) ? node34447 : 4'b1011;
																assign node34447 = (inp[2]) ? 4'b1110 : 4'b1011;
												assign node34450 = (inp[1]) ? node34466 : node34451;
													assign node34451 = (inp[13]) ? node34459 : node34452;
														assign node34452 = (inp[2]) ? node34456 : node34453;
															assign node34453 = (inp[7]) ? 4'b1010 : 4'b1111;
															assign node34456 = (inp[7]) ? 4'b1110 : 4'b1010;
														assign node34459 = (inp[7]) ? node34463 : node34460;
															assign node34460 = (inp[2]) ? 4'b1011 : 4'b1110;
															assign node34463 = (inp[2]) ? 4'b1110 : 4'b1011;
													assign node34466 = (inp[2]) ? node34472 : node34467;
														assign node34467 = (inp[7]) ? 4'b1111 : node34468;
															assign node34468 = (inp[13]) ? 4'b1010 : 4'b1011;
														assign node34472 = (inp[7]) ? 4'b1010 : 4'b1111;
											assign node34475 = (inp[7]) ? node34499 : node34476;
												assign node34476 = (inp[2]) ? node34488 : node34477;
													assign node34477 = (inp[1]) ? node34483 : node34478;
														assign node34478 = (inp[15]) ? node34480 : 4'b1010;
															assign node34480 = (inp[13]) ? 4'b1111 : 4'b1110;
														assign node34483 = (inp[15]) ? node34485 : 4'b1111;
															assign node34485 = (inp[13]) ? 4'b1011 : 4'b1010;
													assign node34488 = (inp[1]) ? node34496 : node34489;
														assign node34489 = (inp[15]) ? node34493 : node34490;
															assign node34490 = (inp[13]) ? 4'b1111 : 4'b1110;
															assign node34493 = (inp[13]) ? 4'b1010 : 4'b1011;
														assign node34496 = (inp[15]) ? 4'b1110 : 4'b1010;
												assign node34499 = (inp[2]) ? node34511 : node34500;
													assign node34500 = (inp[1]) ? node34508 : node34501;
														assign node34501 = (inp[15]) ? node34505 : node34502;
															assign node34502 = (inp[13]) ? 4'b1111 : 4'b1110;
															assign node34505 = (inp[13]) ? 4'b1010 : 4'b1011;
														assign node34508 = (inp[15]) ? 4'b1110 : 4'b1010;
													assign node34511 = (inp[15]) ? node34519 : node34512;
														assign node34512 = (inp[1]) ? node34516 : node34513;
															assign node34513 = (inp[13]) ? 4'b1010 : 4'b1011;
															assign node34516 = (inp[13]) ? 4'b1111 : 4'b1110;
														assign node34519 = (inp[1]) ? 4'b1011 : 4'b1111;
									assign node34522 = (inp[1]) ? node34608 : node34523;
										assign node34523 = (inp[2]) ? node34555 : node34524;
											assign node34524 = (inp[0]) ? node34540 : node34525;
												assign node34525 = (inp[10]) ? node34533 : node34526;
													assign node34526 = (inp[7]) ? 4'b1010 : node34527;
														assign node34527 = (inp[15]) ? 4'b1010 : node34528;
															assign node34528 = (inp[13]) ? 4'b1011 : 4'b1010;
													assign node34533 = (inp[15]) ? 4'b1011 : node34534;
														assign node34534 = (inp[13]) ? node34536 : 4'b1011;
															assign node34536 = (inp[7]) ? 4'b1011 : 4'b1010;
												assign node34540 = (inp[10]) ? node34548 : node34541;
													assign node34541 = (inp[15]) ? 4'b1011 : node34542;
														assign node34542 = (inp[13]) ? node34544 : 4'b1011;
															assign node34544 = (inp[7]) ? 4'b1011 : 4'b1010;
													assign node34548 = (inp[15]) ? 4'b1010 : node34549;
														assign node34549 = (inp[7]) ? 4'b1010 : node34550;
															assign node34550 = (inp[13]) ? 4'b1011 : 4'b1010;
											assign node34555 = (inp[13]) ? node34579 : node34556;
												assign node34556 = (inp[0]) ? node34568 : node34557;
													assign node34557 = (inp[10]) ? node34563 : node34558;
														assign node34558 = (inp[7]) ? node34560 : 4'b1111;
															assign node34560 = (inp[15]) ? 4'b1111 : 4'b1110;
														assign node34563 = (inp[7]) ? node34565 : 4'b1110;
															assign node34565 = (inp[15]) ? 4'b1110 : 4'b1111;
													assign node34568 = (inp[10]) ? node34574 : node34569;
														assign node34569 = (inp[15]) ? 4'b1110 : node34570;
															assign node34570 = (inp[7]) ? 4'b1111 : 4'b1110;
														assign node34574 = (inp[7]) ? node34576 : 4'b1111;
															assign node34576 = (inp[15]) ? 4'b1111 : 4'b1110;
												assign node34579 = (inp[0]) ? node34593 : node34580;
													assign node34580 = (inp[7]) ? node34588 : node34581;
														assign node34581 = (inp[15]) ? node34585 : node34582;
															assign node34582 = (inp[10]) ? 4'b1110 : 4'b1111;
															assign node34585 = (inp[10]) ? 4'b1111 : 4'b1110;
														assign node34588 = (inp[10]) ? 4'b1110 : node34589;
															assign node34589 = (inp[15]) ? 4'b1110 : 4'b1111;
													assign node34593 = (inp[9]) ? node34601 : node34594;
														assign node34594 = (inp[10]) ? node34598 : node34595;
															assign node34595 = (inp[15]) ? 4'b1111 : 4'b1110;
															assign node34598 = (inp[15]) ? 4'b1110 : 4'b1111;
														assign node34601 = (inp[15]) ? node34605 : node34602;
															assign node34602 = (inp[10]) ? 4'b1111 : 4'b1110;
															assign node34605 = (inp[10]) ? 4'b1110 : 4'b1111;
										assign node34608 = (inp[2]) ? node34714 : node34609;
											assign node34609 = (inp[7]) ? node34665 : node34610;
												assign node34610 = (inp[0]) ? node34634 : node34611;
													assign node34611 = (inp[10]) ? node34619 : node34612;
														assign node34612 = (inp[15]) ? node34616 : node34613;
															assign node34613 = (inp[13]) ? 4'b1110 : 4'b1111;
															assign node34616 = (inp[13]) ? 4'b1111 : 4'b1110;
														assign node34619 = (inp[9]) ? node34627 : node34620;
															assign node34620 = (inp[13]) ? node34624 : node34621;
																assign node34621 = (inp[15]) ? 4'b1111 : 4'b1110;
																assign node34624 = (inp[15]) ? 4'b1110 : 4'b1111;
															assign node34627 = (inp[13]) ? node34631 : node34628;
																assign node34628 = (inp[15]) ? 4'b1111 : 4'b1110;
																assign node34631 = (inp[15]) ? 4'b1110 : 4'b1111;
													assign node34634 = (inp[10]) ? node34650 : node34635;
														assign node34635 = (inp[9]) ? node34643 : node34636;
															assign node34636 = (inp[13]) ? node34640 : node34637;
																assign node34637 = (inp[15]) ? 4'b1111 : 4'b1110;
																assign node34640 = (inp[15]) ? 4'b1110 : 4'b1111;
															assign node34643 = (inp[13]) ? node34647 : node34644;
																assign node34644 = (inp[15]) ? 4'b1111 : 4'b1110;
																assign node34647 = (inp[15]) ? 4'b1110 : 4'b1111;
														assign node34650 = (inp[9]) ? node34658 : node34651;
															assign node34651 = (inp[13]) ? node34655 : node34652;
																assign node34652 = (inp[15]) ? 4'b1110 : 4'b1111;
																assign node34655 = (inp[15]) ? 4'b1111 : 4'b1110;
															assign node34658 = (inp[15]) ? node34662 : node34659;
																assign node34659 = (inp[13]) ? 4'b1110 : 4'b1111;
																assign node34662 = (inp[13]) ? 4'b1111 : 4'b1110;
												assign node34665 = (inp[9]) ? node34685 : node34666;
													assign node34666 = (inp[10]) ? node34678 : node34667;
														assign node34667 = (inp[0]) ? node34673 : node34668;
															assign node34668 = (inp[13]) ? 4'b1111 : node34669;
																assign node34669 = (inp[15]) ? 4'b1110 : 4'b1111;
															assign node34673 = (inp[13]) ? 4'b1110 : node34674;
																assign node34674 = (inp[15]) ? 4'b1111 : 4'b1110;
														assign node34678 = (inp[0]) ? node34680 : 4'b1110;
															assign node34680 = (inp[13]) ? 4'b1111 : node34681;
																assign node34681 = (inp[15]) ? 4'b1110 : 4'b1111;
													assign node34685 = (inp[13]) ? node34699 : node34686;
														assign node34686 = (inp[0]) ? node34692 : node34687;
															assign node34687 = (inp[15]) ? node34689 : 4'b1110;
																assign node34689 = (inp[10]) ? 4'b1111 : 4'b1110;
															assign node34692 = (inp[10]) ? node34696 : node34693;
																assign node34693 = (inp[15]) ? 4'b1111 : 4'b1110;
																assign node34696 = (inp[15]) ? 4'b1110 : 4'b1111;
														assign node34699 = (inp[15]) ? node34707 : node34700;
															assign node34700 = (inp[10]) ? node34704 : node34701;
																assign node34701 = (inp[0]) ? 4'b1110 : 4'b1111;
																assign node34704 = (inp[0]) ? 4'b1111 : 4'b1110;
															assign node34707 = (inp[10]) ? node34711 : node34708;
																assign node34708 = (inp[0]) ? 4'b1110 : 4'b1111;
																assign node34711 = (inp[0]) ? 4'b1111 : 4'b1110;
											assign node34714 = (inp[7]) ? node34754 : node34715;
												assign node34715 = (inp[0]) ? node34731 : node34716;
													assign node34716 = (inp[13]) ? node34724 : node34717;
														assign node34717 = (inp[10]) ? node34721 : node34718;
															assign node34718 = (inp[15]) ? 4'b1011 : 4'b1010;
															assign node34721 = (inp[15]) ? 4'b1010 : 4'b1011;
														assign node34724 = (inp[10]) ? node34728 : node34725;
															assign node34725 = (inp[15]) ? 4'b1010 : 4'b1011;
															assign node34728 = (inp[15]) ? 4'b1011 : 4'b1010;
													assign node34731 = (inp[9]) ? node34741 : node34732;
														assign node34732 = (inp[10]) ? node34734 : 4'b1010;
															assign node34734 = (inp[13]) ? node34738 : node34735;
																assign node34735 = (inp[15]) ? 4'b1011 : 4'b1010;
																assign node34738 = (inp[15]) ? 4'b1010 : 4'b1011;
														assign node34741 = (inp[10]) ? node34749 : node34742;
															assign node34742 = (inp[13]) ? node34746 : node34743;
																assign node34743 = (inp[15]) ? 4'b1010 : 4'b1011;
																assign node34746 = (inp[15]) ? 4'b1011 : 4'b1010;
															assign node34749 = (inp[15]) ? node34751 : 4'b1011;
																assign node34751 = (inp[13]) ? 4'b1010 : 4'b1011;
												assign node34754 = (inp[15]) ? node34770 : node34755;
													assign node34755 = (inp[9]) ? node34763 : node34756;
														assign node34756 = (inp[10]) ? node34760 : node34757;
															assign node34757 = (inp[0]) ? 4'b1011 : 4'b1010;
															assign node34760 = (inp[0]) ? 4'b1010 : 4'b1011;
														assign node34763 = (inp[10]) ? node34767 : node34764;
															assign node34764 = (inp[0]) ? 4'b1011 : 4'b1010;
															assign node34767 = (inp[0]) ? 4'b1010 : 4'b1011;
													assign node34770 = (inp[9]) ? node34786 : node34771;
														assign node34771 = (inp[13]) ? node34779 : node34772;
															assign node34772 = (inp[10]) ? node34776 : node34773;
																assign node34773 = (inp[0]) ? 4'b1010 : 4'b1011;
																assign node34776 = (inp[0]) ? 4'b1011 : 4'b1010;
															assign node34779 = (inp[0]) ? node34783 : node34780;
																assign node34780 = (inp[10]) ? 4'b1011 : 4'b1010;
																assign node34783 = (inp[10]) ? 4'b1010 : 4'b1011;
														assign node34786 = (inp[13]) ? node34794 : node34787;
															assign node34787 = (inp[10]) ? node34791 : node34788;
																assign node34788 = (inp[0]) ? 4'b1010 : 4'b1011;
																assign node34791 = (inp[0]) ? 4'b1011 : 4'b1010;
															assign node34794 = (inp[0]) ? 4'b1010 : node34795;
																assign node34795 = (inp[10]) ? 4'b1011 : 4'b1010;
								assign node34799 = (inp[10]) ? node34977 : node34800;
									assign node34800 = (inp[0]) ? node34886 : node34801;
										assign node34801 = (inp[2]) ? node34843 : node34802;
											assign node34802 = (inp[1]) ? node34822 : node34803;
												assign node34803 = (inp[5]) ? node34813 : node34804;
													assign node34804 = (inp[7]) ? node34810 : node34805;
														assign node34805 = (inp[15]) ? 4'b1111 : node34806;
															assign node34806 = (inp[13]) ? 4'b1010 : 4'b1011;
														assign node34810 = (inp[15]) ? 4'b1010 : 4'b1110;
													assign node34813 = (inp[13]) ? node34819 : node34814;
														assign node34814 = (inp[15]) ? 4'b1010 : node34815;
															assign node34815 = (inp[7]) ? 4'b1011 : 4'b1010;
														assign node34819 = (inp[15]) ? 4'b1011 : 4'b1010;
												assign node34822 = (inp[5]) ? node34836 : node34823;
													assign node34823 = (inp[15]) ? node34831 : node34824;
														assign node34824 = (inp[7]) ? node34828 : node34825;
															assign node34825 = (inp[13]) ? 4'b1111 : 4'b1110;
															assign node34828 = (inp[13]) ? 4'b1010 : 4'b1011;
														assign node34831 = (inp[7]) ? node34833 : 4'b1011;
															assign node34833 = (inp[9]) ? 4'b1111 : 4'b1110;
													assign node34836 = (inp[15]) ? 4'b1111 : node34837;
														assign node34837 = (inp[13]) ? 4'b1111 : node34838;
															assign node34838 = (inp[7]) ? 4'b1110 : 4'b1111;
											assign node34843 = (inp[1]) ? node34861 : node34844;
												assign node34844 = (inp[5]) ? node34854 : node34845;
													assign node34845 = (inp[7]) ? node34849 : node34846;
														assign node34846 = (inp[15]) ? 4'b1010 : 4'b1110;
														assign node34849 = (inp[15]) ? node34851 : 4'b1011;
															assign node34851 = (inp[13]) ? 4'b1110 : 4'b1111;
													assign node34854 = (inp[7]) ? 4'b1110 : node34855;
														assign node34855 = (inp[15]) ? 4'b1110 : node34856;
															assign node34856 = (inp[13]) ? 4'b1111 : 4'b1110;
												assign node34861 = (inp[5]) ? node34879 : node34862;
													assign node34862 = (inp[13]) ? node34870 : node34863;
														assign node34863 = (inp[7]) ? node34867 : node34864;
															assign node34864 = (inp[15]) ? 4'b1110 : 4'b1011;
															assign node34867 = (inp[15]) ? 4'b1011 : 4'b1110;
														assign node34870 = (inp[9]) ? 4'b1010 : node34871;
															assign node34871 = (inp[7]) ? node34875 : node34872;
																assign node34872 = (inp[15]) ? 4'b1111 : 4'b1010;
																assign node34875 = (inp[15]) ? 4'b1010 : 4'b1110;
													assign node34879 = (inp[7]) ? node34881 : 4'b1010;
														assign node34881 = (inp[13]) ? 4'b1010 : node34882;
															assign node34882 = (inp[15]) ? 4'b1010 : 4'b1011;
										assign node34886 = (inp[2]) ? node34936 : node34887;
											assign node34887 = (inp[1]) ? node34907 : node34888;
												assign node34888 = (inp[5]) ? node34898 : node34889;
													assign node34889 = (inp[7]) ? node34895 : node34890;
														assign node34890 = (inp[15]) ? 4'b1110 : node34891;
															assign node34891 = (inp[13]) ? 4'b1011 : 4'b1010;
														assign node34895 = (inp[15]) ? 4'b1011 : 4'b1111;
													assign node34898 = (inp[13]) ? node34904 : node34899;
														assign node34899 = (inp[15]) ? 4'b1011 : node34900;
															assign node34900 = (inp[7]) ? 4'b1010 : 4'b1011;
														assign node34904 = (inp[15]) ? 4'b1010 : 4'b1011;
												assign node34907 = (inp[5]) ? node34929 : node34908;
													assign node34908 = (inp[13]) ? node34922 : node34909;
														assign node34909 = (inp[9]) ? node34917 : node34910;
															assign node34910 = (inp[7]) ? node34914 : node34911;
																assign node34911 = (inp[15]) ? 4'b1010 : 4'b1111;
																assign node34914 = (inp[15]) ? 4'b1111 : 4'b1010;
															assign node34917 = (inp[15]) ? 4'b1111 : node34918;
																assign node34918 = (inp[7]) ? 4'b1010 : 4'b1111;
														assign node34922 = (inp[15]) ? node34926 : node34923;
															assign node34923 = (inp[7]) ? 4'b1011 : 4'b1110;
															assign node34926 = (inp[7]) ? 4'b1110 : 4'b1010;
													assign node34929 = (inp[15]) ? 4'b1110 : node34930;
														assign node34930 = (inp[13]) ? 4'b1110 : node34931;
															assign node34931 = (inp[7]) ? 4'b1111 : 4'b1110;
											assign node34936 = (inp[1]) ? node34954 : node34937;
												assign node34937 = (inp[5]) ? node34947 : node34938;
													assign node34938 = (inp[7]) ? node34942 : node34939;
														assign node34939 = (inp[15]) ? 4'b1011 : 4'b1111;
														assign node34942 = (inp[15]) ? node34944 : 4'b1010;
															assign node34944 = (inp[13]) ? 4'b1111 : 4'b1110;
													assign node34947 = (inp[15]) ? 4'b1111 : node34948;
														assign node34948 = (inp[13]) ? node34950 : 4'b1111;
															assign node34950 = (inp[7]) ? 4'b1111 : 4'b1110;
												assign node34954 = (inp[5]) ? node34970 : node34955;
													assign node34955 = (inp[13]) ? node34963 : node34956;
														assign node34956 = (inp[7]) ? node34960 : node34957;
															assign node34957 = (inp[15]) ? 4'b1111 : 4'b1010;
															assign node34960 = (inp[15]) ? 4'b1010 : 4'b1111;
														assign node34963 = (inp[7]) ? node34967 : node34964;
															assign node34964 = (inp[15]) ? 4'b1110 : 4'b1011;
															assign node34967 = (inp[15]) ? 4'b1011 : 4'b1111;
													assign node34970 = (inp[13]) ? 4'b1011 : node34971;
														assign node34971 = (inp[7]) ? node34973 : 4'b1011;
															assign node34973 = (inp[15]) ? 4'b1011 : 4'b1010;
									assign node34977 = (inp[0]) ? node35061 : node34978;
										assign node34978 = (inp[2]) ? node35020 : node34979;
											assign node34979 = (inp[1]) ? node34999 : node34980;
												assign node34980 = (inp[5]) ? node34990 : node34981;
													assign node34981 = (inp[7]) ? node34987 : node34982;
														assign node34982 = (inp[15]) ? 4'b1110 : node34983;
															assign node34983 = (inp[13]) ? 4'b1011 : 4'b1010;
														assign node34987 = (inp[15]) ? 4'b1011 : 4'b1111;
													assign node34990 = (inp[13]) ? node34996 : node34991;
														assign node34991 = (inp[15]) ? 4'b1011 : node34992;
															assign node34992 = (inp[7]) ? 4'b1010 : 4'b1011;
														assign node34996 = (inp[15]) ? 4'b1010 : 4'b1011;
												assign node34999 = (inp[5]) ? node35013 : node35000;
													assign node35000 = (inp[7]) ? node35006 : node35001;
														assign node35001 = (inp[15]) ? 4'b1010 : node35002;
															assign node35002 = (inp[13]) ? 4'b1110 : 4'b1111;
														assign node35006 = (inp[15]) ? node35010 : node35007;
															assign node35007 = (inp[13]) ? 4'b1011 : 4'b1010;
															assign node35010 = (inp[13]) ? 4'b1110 : 4'b1111;
													assign node35013 = (inp[13]) ? 4'b1110 : node35014;
														assign node35014 = (inp[15]) ? 4'b1110 : node35015;
															assign node35015 = (inp[7]) ? 4'b1111 : 4'b1110;
											assign node35020 = (inp[1]) ? node35038 : node35021;
												assign node35021 = (inp[5]) ? node35031 : node35022;
													assign node35022 = (inp[7]) ? node35026 : node35023;
														assign node35023 = (inp[15]) ? 4'b1011 : 4'b1111;
														assign node35026 = (inp[15]) ? node35028 : 4'b1010;
															assign node35028 = (inp[13]) ? 4'b1111 : 4'b1110;
													assign node35031 = (inp[15]) ? 4'b1111 : node35032;
														assign node35032 = (inp[13]) ? node35034 : 4'b1111;
															assign node35034 = (inp[7]) ? 4'b1111 : 4'b1110;
												assign node35038 = (inp[5]) ? node35054 : node35039;
													assign node35039 = (inp[13]) ? node35047 : node35040;
														assign node35040 = (inp[15]) ? node35044 : node35041;
															assign node35041 = (inp[7]) ? 4'b1111 : 4'b1010;
															assign node35044 = (inp[7]) ? 4'b1010 : 4'b1111;
														assign node35047 = (inp[7]) ? node35051 : node35048;
															assign node35048 = (inp[15]) ? 4'b1110 : 4'b1011;
															assign node35051 = (inp[15]) ? 4'b1011 : 4'b1111;
													assign node35054 = (inp[13]) ? 4'b1011 : node35055;
														assign node35055 = (inp[7]) ? node35057 : 4'b1011;
															assign node35057 = (inp[15]) ? 4'b1011 : 4'b1010;
										assign node35061 = (inp[2]) ? node35101 : node35062;
											assign node35062 = (inp[1]) ? node35082 : node35063;
												assign node35063 = (inp[5]) ? node35073 : node35064;
													assign node35064 = (inp[7]) ? node35070 : node35065;
														assign node35065 = (inp[15]) ? 4'b1111 : node35066;
															assign node35066 = (inp[13]) ? 4'b1010 : 4'b1011;
														assign node35070 = (inp[15]) ? 4'b1010 : 4'b1110;
													assign node35073 = (inp[13]) ? node35079 : node35074;
														assign node35074 = (inp[7]) ? node35076 : 4'b1010;
															assign node35076 = (inp[15]) ? 4'b1010 : 4'b1011;
														assign node35079 = (inp[15]) ? 4'b1011 : 4'b1010;
												assign node35082 = (inp[5]) ? node35094 : node35083;
													assign node35083 = (inp[7]) ? node35089 : node35084;
														assign node35084 = (inp[15]) ? 4'b1011 : node35085;
															assign node35085 = (inp[13]) ? 4'b1111 : 4'b1110;
														assign node35089 = (inp[15]) ? 4'b1110 : node35090;
															assign node35090 = (inp[13]) ? 4'b1010 : 4'b1011;
													assign node35094 = (inp[13]) ? 4'b1111 : node35095;
														assign node35095 = (inp[7]) ? node35097 : 4'b1111;
															assign node35097 = (inp[15]) ? 4'b1111 : 4'b1110;
											assign node35101 = (inp[1]) ? node35119 : node35102;
												assign node35102 = (inp[5]) ? node35112 : node35103;
													assign node35103 = (inp[7]) ? node35107 : node35104;
														assign node35104 = (inp[15]) ? 4'b1010 : 4'b1110;
														assign node35107 = (inp[15]) ? node35109 : 4'b1011;
															assign node35109 = (inp[13]) ? 4'b1110 : 4'b1111;
													assign node35112 = (inp[13]) ? node35114 : 4'b1110;
														assign node35114 = (inp[7]) ? 4'b1110 : node35115;
															assign node35115 = (inp[15]) ? 4'b1110 : 4'b1111;
												assign node35119 = (inp[5]) ? node35133 : node35120;
													assign node35120 = (inp[7]) ? node35128 : node35121;
														assign node35121 = (inp[15]) ? node35125 : node35122;
															assign node35122 = (inp[13]) ? 4'b1010 : 4'b1011;
															assign node35125 = (inp[13]) ? 4'b1111 : 4'b1110;
														assign node35128 = (inp[15]) ? node35130 : 4'b1110;
															assign node35130 = (inp[13]) ? 4'b1010 : 4'b1011;
													assign node35133 = (inp[13]) ? 4'b1010 : node35134;
														assign node35134 = (inp[9]) ? node35136 : 4'b1010;
															assign node35136 = (inp[15]) ? 4'b1010 : node35137;
																assign node35137 = (inp[7]) ? 4'b1011 : 4'b1010;
						assign node35142 = (inp[7]) ? node36636 : node35143;
							assign node35143 = (inp[8]) ? node35923 : node35144;
								assign node35144 = (inp[15]) ? node35480 : node35145;
									assign node35145 = (inp[2]) ? node35307 : node35146;
										assign node35146 = (inp[13]) ? node35218 : node35147;
											assign node35147 = (inp[5]) ? node35181 : node35148;
												assign node35148 = (inp[1]) ? node35162 : node35149;
													assign node35149 = (inp[10]) ? node35153 : node35150;
														assign node35150 = (inp[9]) ? 4'b1111 : 4'b1110;
														assign node35153 = (inp[9]) ? node35159 : node35154;
															assign node35154 = (inp[11]) ? node35156 : 4'b1111;
																assign node35156 = (inp[0]) ? 4'b1111 : 4'b1110;
															assign node35159 = (inp[0]) ? 4'b1110 : 4'b1111;
													assign node35162 = (inp[10]) ? node35174 : node35163;
														assign node35163 = (inp[9]) ? node35169 : node35164;
															assign node35164 = (inp[11]) ? 4'b1011 : node35165;
																assign node35165 = (inp[0]) ? 4'b1010 : 4'b1011;
															assign node35169 = (inp[0]) ? node35171 : 4'b1010;
																assign node35171 = (inp[11]) ? 4'b1010 : 4'b1011;
														assign node35174 = (inp[9]) ? 4'b1011 : node35175;
															assign node35175 = (inp[0]) ? node35177 : 4'b1010;
																assign node35177 = (inp[11]) ? 4'b1010 : 4'b1011;
												assign node35181 = (inp[1]) ? node35201 : node35182;
													assign node35182 = (inp[11]) ? node35192 : node35183;
														assign node35183 = (inp[0]) ? node35185 : 4'b1111;
															assign node35185 = (inp[9]) ? node35189 : node35186;
																assign node35186 = (inp[10]) ? 4'b1110 : 4'b1111;
																assign node35189 = (inp[10]) ? 4'b1111 : 4'b1110;
														assign node35192 = (inp[0]) ? 4'b1111 : node35193;
															assign node35193 = (inp[9]) ? node35197 : node35194;
																assign node35194 = (inp[10]) ? 4'b1111 : 4'b1110;
																assign node35197 = (inp[10]) ? 4'b1110 : 4'b1111;
													assign node35201 = (inp[10]) ? node35213 : node35202;
														assign node35202 = (inp[9]) ? node35208 : node35203;
															assign node35203 = (inp[0]) ? 4'b1110 : node35204;
																assign node35204 = (inp[11]) ? 4'b1111 : 4'b1110;
															assign node35208 = (inp[0]) ? 4'b1111 : node35209;
																assign node35209 = (inp[11]) ? 4'b1110 : 4'b1111;
														assign node35213 = (inp[9]) ? 4'b1110 : node35214;
															assign node35214 = (inp[0]) ? 4'b1111 : 4'b1110;
											assign node35218 = (inp[5]) ? node35258 : node35219;
												assign node35219 = (inp[1]) ? node35237 : node35220;
													assign node35220 = (inp[10]) ? node35228 : node35221;
														assign node35221 = (inp[9]) ? 4'b1011 : node35222;
															assign node35222 = (inp[11]) ? 4'b1010 : node35223;
																assign node35223 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node35228 = (inp[9]) ? node35232 : node35229;
															assign node35229 = (inp[11]) ? 4'b1011 : 4'b1010;
															assign node35232 = (inp[0]) ? node35234 : 4'b1010;
																assign node35234 = (inp[11]) ? 4'b1010 : 4'b1011;
													assign node35237 = (inp[9]) ? node35247 : node35238;
														assign node35238 = (inp[10]) ? node35244 : node35239;
															assign node35239 = (inp[0]) ? node35241 : 4'b1111;
																assign node35241 = (inp[11]) ? 4'b1111 : 4'b1110;
															assign node35244 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node35247 = (inp[10]) ? node35253 : node35248;
															assign node35248 = (inp[0]) ? node35250 : 4'b1110;
																assign node35250 = (inp[11]) ? 4'b1110 : 4'b1111;
															assign node35253 = (inp[11]) ? 4'b1111 : node35254;
																assign node35254 = (inp[0]) ? 4'b1110 : 4'b1111;
												assign node35258 = (inp[9]) ? node35282 : node35259;
													assign node35259 = (inp[0]) ? node35267 : node35260;
														assign node35260 = (inp[10]) ? node35264 : node35261;
															assign node35261 = (inp[1]) ? 4'b1010 : 4'b1011;
															assign node35264 = (inp[1]) ? 4'b1011 : 4'b1010;
														assign node35267 = (inp[11]) ? node35275 : node35268;
															assign node35268 = (inp[10]) ? node35272 : node35269;
																assign node35269 = (inp[1]) ? 4'b1011 : 4'b1010;
																assign node35272 = (inp[1]) ? 4'b1010 : 4'b1011;
															assign node35275 = (inp[1]) ? node35279 : node35276;
																assign node35276 = (inp[10]) ? 4'b1010 : 4'b1011;
																assign node35279 = (inp[10]) ? 4'b1011 : 4'b1010;
													assign node35282 = (inp[11]) ? node35292 : node35283;
														assign node35283 = (inp[0]) ? node35285 : 4'b1010;
															assign node35285 = (inp[1]) ? node35289 : node35286;
																assign node35286 = (inp[10]) ? 4'b1010 : 4'b1011;
																assign node35289 = (inp[10]) ? 4'b1011 : 4'b1010;
														assign node35292 = (inp[0]) ? node35300 : node35293;
															assign node35293 = (inp[1]) ? node35297 : node35294;
																assign node35294 = (inp[10]) ? 4'b1011 : 4'b1010;
																assign node35297 = (inp[10]) ? 4'b1010 : 4'b1011;
															assign node35300 = (inp[10]) ? node35304 : node35301;
																assign node35301 = (inp[1]) ? 4'b1011 : 4'b1010;
																assign node35304 = (inp[1]) ? 4'b1010 : 4'b1011;
										assign node35307 = (inp[13]) ? node35395 : node35308;
											assign node35308 = (inp[5]) ? node35342 : node35309;
												assign node35309 = (inp[1]) ? node35321 : node35310;
													assign node35310 = (inp[9]) ? node35316 : node35311;
														assign node35311 = (inp[10]) ? node35313 : 4'b1010;
															assign node35313 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node35316 = (inp[10]) ? node35318 : 4'b1011;
															assign node35318 = (inp[0]) ? 4'b1010 : 4'b1011;
													assign node35321 = (inp[9]) ? node35331 : node35322;
														assign node35322 = (inp[10]) ? node35328 : node35323;
															assign node35323 = (inp[0]) ? 4'b1111 : node35324;
																assign node35324 = (inp[11]) ? 4'b1110 : 4'b1111;
															assign node35328 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node35331 = (inp[10]) ? node35337 : node35332;
															assign node35332 = (inp[0]) ? 4'b1110 : node35333;
																assign node35333 = (inp[11]) ? 4'b1111 : 4'b1110;
															assign node35337 = (inp[11]) ? node35339 : 4'b1111;
																assign node35339 = (inp[0]) ? 4'b1111 : 4'b1110;
												assign node35342 = (inp[10]) ? node35372 : node35343;
													assign node35343 = (inp[11]) ? node35359 : node35344;
														assign node35344 = (inp[0]) ? node35352 : node35345;
															assign node35345 = (inp[1]) ? node35349 : node35346;
																assign node35346 = (inp[9]) ? 4'b1010 : 4'b1011;
																assign node35349 = (inp[9]) ? 4'b1011 : 4'b1010;
															assign node35352 = (inp[1]) ? node35356 : node35353;
																assign node35353 = (inp[9]) ? 4'b1010 : 4'b1011;
																assign node35356 = (inp[9]) ? 4'b1011 : 4'b1010;
														assign node35359 = (inp[9]) ? node35365 : node35360;
															assign node35360 = (inp[1]) ? node35362 : 4'b1010;
																assign node35362 = (inp[0]) ? 4'b1010 : 4'b1011;
															assign node35365 = (inp[0]) ? node35369 : node35366;
																assign node35366 = (inp[1]) ? 4'b1010 : 4'b1011;
																assign node35369 = (inp[1]) ? 4'b1011 : 4'b1010;
													assign node35372 = (inp[0]) ? node35388 : node35373;
														assign node35373 = (inp[1]) ? node35381 : node35374;
															assign node35374 = (inp[11]) ? node35378 : node35375;
																assign node35375 = (inp[9]) ? 4'b1011 : 4'b1010;
																assign node35378 = (inp[9]) ? 4'b1010 : 4'b1011;
															assign node35381 = (inp[11]) ? node35385 : node35382;
																assign node35382 = (inp[9]) ? 4'b1010 : 4'b1011;
																assign node35385 = (inp[9]) ? 4'b1011 : 4'b1010;
														assign node35388 = (inp[1]) ? node35392 : node35389;
															assign node35389 = (inp[9]) ? 4'b1011 : 4'b1010;
															assign node35392 = (inp[9]) ? 4'b1010 : 4'b1011;
											assign node35395 = (inp[1]) ? node35441 : node35396;
												assign node35396 = (inp[5]) ? node35420 : node35397;
													assign node35397 = (inp[11]) ? node35405 : node35398;
														assign node35398 = (inp[9]) ? node35402 : node35399;
															assign node35399 = (inp[10]) ? 4'b1111 : 4'b1110;
															assign node35402 = (inp[10]) ? 4'b1110 : 4'b1111;
														assign node35405 = (inp[0]) ? node35413 : node35406;
															assign node35406 = (inp[10]) ? node35410 : node35407;
																assign node35407 = (inp[9]) ? 4'b1110 : 4'b1111;
																assign node35410 = (inp[9]) ? 4'b1111 : 4'b1110;
															assign node35413 = (inp[10]) ? node35417 : node35414;
																assign node35414 = (inp[9]) ? 4'b1111 : 4'b1110;
																assign node35417 = (inp[9]) ? 4'b1110 : 4'b1111;
													assign node35420 = (inp[10]) ? node35432 : node35421;
														assign node35421 = (inp[9]) ? node35427 : node35422;
															assign node35422 = (inp[0]) ? 4'b1111 : node35423;
																assign node35423 = (inp[11]) ? 4'b1110 : 4'b1111;
															assign node35427 = (inp[0]) ? 4'b1110 : node35428;
																assign node35428 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node35432 = (inp[9]) ? node35438 : node35433;
															assign node35433 = (inp[11]) ? node35435 : 4'b1110;
																assign node35435 = (inp[0]) ? 4'b1110 : 4'b1111;
															assign node35438 = (inp[0]) ? 4'b1111 : 4'b1110;
												assign node35441 = (inp[5]) ? node35463 : node35442;
													assign node35442 = (inp[10]) ? node35454 : node35443;
														assign node35443 = (inp[9]) ? node35449 : node35444;
															assign node35444 = (inp[11]) ? 4'b1011 : node35445;
																assign node35445 = (inp[0]) ? 4'b1010 : 4'b1011;
															assign node35449 = (inp[11]) ? 4'b1010 : node35450;
																assign node35450 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node35454 = (inp[9]) ? node35458 : node35455;
															assign node35455 = (inp[11]) ? 4'b1010 : 4'b1011;
															assign node35458 = (inp[11]) ? 4'b1011 : node35459;
																assign node35459 = (inp[0]) ? 4'b1010 : 4'b1011;
													assign node35463 = (inp[9]) ? node35469 : node35464;
														assign node35464 = (inp[0]) ? node35466 : 4'b1111;
															assign node35466 = (inp[10]) ? 4'b1111 : 4'b1110;
														assign node35469 = (inp[10]) ? node35475 : node35470;
															assign node35470 = (inp[11]) ? node35472 : 4'b1111;
																assign node35472 = (inp[0]) ? 4'b1111 : 4'b1110;
															assign node35475 = (inp[0]) ? 4'b1110 : node35476;
																assign node35476 = (inp[11]) ? 4'b1111 : 4'b1110;
									assign node35480 = (inp[0]) ? node35702 : node35481;
										assign node35481 = (inp[11]) ? node35597 : node35482;
											assign node35482 = (inp[1]) ? node35540 : node35483;
												assign node35483 = (inp[10]) ? node35511 : node35484;
													assign node35484 = (inp[13]) ? node35496 : node35485;
														assign node35485 = (inp[2]) ? node35489 : node35486;
															assign node35486 = (inp[5]) ? 4'b1011 : 4'b1010;
															assign node35489 = (inp[5]) ? node35493 : node35490;
																assign node35490 = (inp[9]) ? 4'b1111 : 4'b1110;
																assign node35493 = (inp[9]) ? 4'b1110 : 4'b1111;
														assign node35496 = (inp[2]) ? node35504 : node35497;
															assign node35497 = (inp[5]) ? node35501 : node35498;
																assign node35498 = (inp[9]) ? 4'b1110 : 4'b1111;
																assign node35501 = (inp[9]) ? 4'b1111 : 4'b1110;
															assign node35504 = (inp[9]) ? node35508 : node35505;
																assign node35505 = (inp[5]) ? 4'b1010 : 4'b1011;
																assign node35508 = (inp[5]) ? 4'b1011 : 4'b1010;
													assign node35511 = (inp[9]) ? node35527 : node35512;
														assign node35512 = (inp[13]) ? node35520 : node35513;
															assign node35513 = (inp[2]) ? node35517 : node35514;
																assign node35514 = (inp[5]) ? 4'b1010 : 4'b1011;
																assign node35517 = (inp[5]) ? 4'b1110 : 4'b1111;
															assign node35520 = (inp[2]) ? node35524 : node35521;
																assign node35521 = (inp[5]) ? 4'b1111 : 4'b1110;
																assign node35524 = (inp[5]) ? 4'b1011 : 4'b1010;
														assign node35527 = (inp[5]) ? node35535 : node35528;
															assign node35528 = (inp[13]) ? node35532 : node35529;
																assign node35529 = (inp[2]) ? 4'b1110 : 4'b1010;
																assign node35532 = (inp[2]) ? 4'b1011 : 4'b1111;
															assign node35535 = (inp[13]) ? node35537 : 4'b1011;
																assign node35537 = (inp[2]) ? 4'b1010 : 4'b1110;
												assign node35540 = (inp[13]) ? node35568 : node35541;
													assign node35541 = (inp[9]) ? node35555 : node35542;
														assign node35542 = (inp[10]) ? node35548 : node35543;
															assign node35543 = (inp[2]) ? node35545 : 4'b1011;
																assign node35545 = (inp[5]) ? 4'b1110 : 4'b1010;
															assign node35548 = (inp[5]) ? node35552 : node35549;
																assign node35549 = (inp[2]) ? 4'b1011 : 4'b1111;
																assign node35552 = (inp[2]) ? 4'b1111 : 4'b1010;
														assign node35555 = (inp[10]) ? node35563 : node35556;
															assign node35556 = (inp[5]) ? node35560 : node35557;
																assign node35557 = (inp[2]) ? 4'b1011 : 4'b1111;
																assign node35560 = (inp[2]) ? 4'b1111 : 4'b1010;
															assign node35563 = (inp[5]) ? 4'b1011 : node35564;
																assign node35564 = (inp[2]) ? 4'b1010 : 4'b1110;
													assign node35568 = (inp[2]) ? node35584 : node35569;
														assign node35569 = (inp[5]) ? node35577 : node35570;
															assign node35570 = (inp[10]) ? node35574 : node35571;
																assign node35571 = (inp[9]) ? 4'b1010 : 4'b1011;
																assign node35574 = (inp[9]) ? 4'b1011 : 4'b1010;
															assign node35577 = (inp[9]) ? node35581 : node35578;
																assign node35578 = (inp[10]) ? 4'b1111 : 4'b1110;
																assign node35581 = (inp[10]) ? 4'b1110 : 4'b1111;
														assign node35584 = (inp[5]) ? node35592 : node35585;
															assign node35585 = (inp[9]) ? node35589 : node35586;
																assign node35586 = (inp[10]) ? 4'b1110 : 4'b1111;
																assign node35589 = (inp[10]) ? 4'b1111 : 4'b1110;
															assign node35592 = (inp[10]) ? 4'b1011 : node35593;
																assign node35593 = (inp[9]) ? 4'b1011 : 4'b1010;
											assign node35597 = (inp[1]) ? node35645 : node35598;
												assign node35598 = (inp[9]) ? node35626 : node35599;
													assign node35599 = (inp[10]) ? node35611 : node35600;
														assign node35600 = (inp[5]) ? node35606 : node35601;
															assign node35601 = (inp[13]) ? node35603 : 4'b1111;
																assign node35603 = (inp[2]) ? 4'b1011 : 4'b1111;
															assign node35606 = (inp[2]) ? 4'b1110 : node35607;
																assign node35607 = (inp[13]) ? 4'b1110 : 4'b1011;
														assign node35611 = (inp[5]) ? node35619 : node35612;
															assign node35612 = (inp[2]) ? node35616 : node35613;
																assign node35613 = (inp[13]) ? 4'b1110 : 4'b1011;
																assign node35616 = (inp[13]) ? 4'b1010 : 4'b1110;
															assign node35619 = (inp[2]) ? node35623 : node35620;
																assign node35620 = (inp[13]) ? 4'b1111 : 4'b1010;
																assign node35623 = (inp[13]) ? 4'b1011 : 4'b1111;
													assign node35626 = (inp[2]) ? node35636 : node35627;
														assign node35627 = (inp[13]) ? node35629 : 4'b1010;
															assign node35629 = (inp[5]) ? node35633 : node35630;
																assign node35630 = (inp[10]) ? 4'b1111 : 4'b1110;
																assign node35633 = (inp[10]) ? 4'b1110 : 4'b1111;
														assign node35636 = (inp[13]) ? 4'b1011 : node35637;
															assign node35637 = (inp[5]) ? node35641 : node35638;
																assign node35638 = (inp[10]) ? 4'b1111 : 4'b1110;
																assign node35641 = (inp[10]) ? 4'b1110 : 4'b1111;
												assign node35645 = (inp[5]) ? node35671 : node35646;
													assign node35646 = (inp[10]) ? node35660 : node35647;
														assign node35647 = (inp[9]) ? node35655 : node35648;
															assign node35648 = (inp[2]) ? node35652 : node35649;
																assign node35649 = (inp[13]) ? 4'b1011 : 4'b1111;
																assign node35652 = (inp[13]) ? 4'b1110 : 4'b1011;
															assign node35655 = (inp[2]) ? 4'b1111 : node35656;
																assign node35656 = (inp[13]) ? 4'b1010 : 4'b1110;
														assign node35660 = (inp[2]) ? node35664 : node35661;
															assign node35661 = (inp[13]) ? 4'b1011 : 4'b1111;
															assign node35664 = (inp[13]) ? node35668 : node35665;
																assign node35665 = (inp[9]) ? 4'b1011 : 4'b1010;
																assign node35668 = (inp[9]) ? 4'b1110 : 4'b1111;
													assign node35671 = (inp[13]) ? node35687 : node35672;
														assign node35672 = (inp[2]) ? node35680 : node35673;
															assign node35673 = (inp[9]) ? node35677 : node35674;
																assign node35674 = (inp[10]) ? 4'b1011 : 4'b1010;
																assign node35677 = (inp[10]) ? 4'b1010 : 4'b1011;
															assign node35680 = (inp[10]) ? node35684 : node35681;
																assign node35681 = (inp[9]) ? 4'b1111 : 4'b1110;
																assign node35684 = (inp[9]) ? 4'b1110 : 4'b1111;
														assign node35687 = (inp[2]) ? node35695 : node35688;
															assign node35688 = (inp[9]) ? node35692 : node35689;
																assign node35689 = (inp[10]) ? 4'b1110 : 4'b1111;
																assign node35692 = (inp[10]) ? 4'b1111 : 4'b1110;
															assign node35695 = (inp[9]) ? node35699 : node35696;
																assign node35696 = (inp[10]) ? 4'b1010 : 4'b1011;
																assign node35699 = (inp[10]) ? 4'b1011 : 4'b1010;
										assign node35702 = (inp[11]) ? node35822 : node35703;
											assign node35703 = (inp[1]) ? node35765 : node35704;
												assign node35704 = (inp[5]) ? node35734 : node35705;
													assign node35705 = (inp[2]) ? node35721 : node35706;
														assign node35706 = (inp[13]) ? node35714 : node35707;
															assign node35707 = (inp[9]) ? node35711 : node35708;
																assign node35708 = (inp[10]) ? 4'b1010 : 4'b1011;
																assign node35711 = (inp[10]) ? 4'b1011 : 4'b1010;
															assign node35714 = (inp[10]) ? node35718 : node35715;
																assign node35715 = (inp[9]) ? 4'b1111 : 4'b1110;
																assign node35718 = (inp[9]) ? 4'b1110 : 4'b1111;
														assign node35721 = (inp[13]) ? node35727 : node35722;
															assign node35722 = (inp[10]) ? 4'b1111 : node35723;
																assign node35723 = (inp[9]) ? 4'b1111 : 4'b1110;
															assign node35727 = (inp[9]) ? node35731 : node35728;
																assign node35728 = (inp[10]) ? 4'b1011 : 4'b1010;
																assign node35731 = (inp[10]) ? 4'b1010 : 4'b1011;
													assign node35734 = (inp[2]) ? node35750 : node35735;
														assign node35735 = (inp[13]) ? node35743 : node35736;
															assign node35736 = (inp[10]) ? node35740 : node35737;
																assign node35737 = (inp[9]) ? 4'b1011 : 4'b1010;
																assign node35740 = (inp[9]) ? 4'b1010 : 4'b1011;
															assign node35743 = (inp[10]) ? node35747 : node35744;
																assign node35744 = (inp[9]) ? 4'b1110 : 4'b1111;
																assign node35747 = (inp[9]) ? 4'b1111 : 4'b1110;
														assign node35750 = (inp[13]) ? node35758 : node35751;
															assign node35751 = (inp[9]) ? node35755 : node35752;
																assign node35752 = (inp[10]) ? 4'b1110 : 4'b1111;
																assign node35755 = (inp[10]) ? 4'b1111 : 4'b1110;
															assign node35758 = (inp[9]) ? node35762 : node35759;
																assign node35759 = (inp[10]) ? 4'b1010 : 4'b1011;
																assign node35762 = (inp[10]) ? 4'b1011 : 4'b1010;
												assign node35765 = (inp[2]) ? node35797 : node35766;
													assign node35766 = (inp[10]) ? node35782 : node35767;
														assign node35767 = (inp[9]) ? node35775 : node35768;
															assign node35768 = (inp[13]) ? node35772 : node35769;
																assign node35769 = (inp[5]) ? 4'b1011 : 4'b1110;
																assign node35772 = (inp[5]) ? 4'b1110 : 4'b1010;
															assign node35775 = (inp[5]) ? node35779 : node35776;
																assign node35776 = (inp[13]) ? 4'b1011 : 4'b1111;
																assign node35779 = (inp[13]) ? 4'b1111 : 4'b1010;
														assign node35782 = (inp[9]) ? node35790 : node35783;
															assign node35783 = (inp[5]) ? node35787 : node35784;
																assign node35784 = (inp[13]) ? 4'b1011 : 4'b1111;
																assign node35787 = (inp[13]) ? 4'b1111 : 4'b1010;
															assign node35790 = (inp[5]) ? node35794 : node35791;
																assign node35791 = (inp[13]) ? 4'b1010 : 4'b1110;
																assign node35794 = (inp[13]) ? 4'b1110 : 4'b1011;
													assign node35797 = (inp[13]) ? node35809 : node35798;
														assign node35798 = (inp[5]) ? node35802 : node35799;
															assign node35799 = (inp[10]) ? 4'b1011 : 4'b1010;
															assign node35802 = (inp[9]) ? node35806 : node35803;
																assign node35803 = (inp[10]) ? 4'b1110 : 4'b1111;
																assign node35806 = (inp[10]) ? 4'b1111 : 4'b1110;
														assign node35809 = (inp[5]) ? node35817 : node35810;
															assign node35810 = (inp[10]) ? node35814 : node35811;
																assign node35811 = (inp[9]) ? 4'b1110 : 4'b1111;
																assign node35814 = (inp[9]) ? 4'b1111 : 4'b1110;
															assign node35817 = (inp[9]) ? node35819 : 4'b1011;
																assign node35819 = (inp[10]) ? 4'b1010 : 4'b1011;
											assign node35822 = (inp[9]) ? node35872 : node35823;
												assign node35823 = (inp[10]) ? node35849 : node35824;
													assign node35824 = (inp[5]) ? node35840 : node35825;
														assign node35825 = (inp[13]) ? node35833 : node35826;
															assign node35826 = (inp[2]) ? node35830 : node35827;
																assign node35827 = (inp[1]) ? 4'b1110 : 4'b1010;
																assign node35830 = (inp[1]) ? 4'b1010 : 4'b1110;
															assign node35833 = (inp[1]) ? node35837 : node35834;
																assign node35834 = (inp[2]) ? 4'b1011 : 4'b1111;
																assign node35837 = (inp[2]) ? 4'b1111 : 4'b1011;
														assign node35840 = (inp[13]) ? node35846 : node35841;
															assign node35841 = (inp[2]) ? node35843 : 4'b1011;
																assign node35843 = (inp[1]) ? 4'b1110 : 4'b1111;
															assign node35846 = (inp[2]) ? 4'b1010 : 4'b1110;
													assign node35849 = (inp[13]) ? node35861 : node35850;
														assign node35850 = (inp[5]) ? node35858 : node35851;
															assign node35851 = (inp[1]) ? node35855 : node35852;
																assign node35852 = (inp[2]) ? 4'b1111 : 4'b1011;
																assign node35855 = (inp[2]) ? 4'b1011 : 4'b1111;
															assign node35858 = (inp[2]) ? 4'b1111 : 4'b1010;
														assign node35861 = (inp[5]) ? node35869 : node35862;
															assign node35862 = (inp[2]) ? node35866 : node35863;
																assign node35863 = (inp[1]) ? 4'b1010 : 4'b1110;
																assign node35866 = (inp[1]) ? 4'b1110 : 4'b1010;
															assign node35869 = (inp[2]) ? 4'b1011 : 4'b1111;
												assign node35872 = (inp[10]) ? node35900 : node35873;
													assign node35873 = (inp[1]) ? node35885 : node35874;
														assign node35874 = (inp[5]) ? node35880 : node35875;
															assign node35875 = (inp[13]) ? node35877 : 4'b1111;
																assign node35877 = (inp[2]) ? 4'b1010 : 4'b1110;
															assign node35880 = (inp[13]) ? 4'b1111 : node35881;
																assign node35881 = (inp[2]) ? 4'b1110 : 4'b1010;
														assign node35885 = (inp[5]) ? node35893 : node35886;
															assign node35886 = (inp[13]) ? node35890 : node35887;
																assign node35887 = (inp[2]) ? 4'b1011 : 4'b1111;
																assign node35890 = (inp[2]) ? 4'b1110 : 4'b1010;
															assign node35893 = (inp[2]) ? node35897 : node35894;
																assign node35894 = (inp[13]) ? 4'b1111 : 4'b1010;
																assign node35897 = (inp[13]) ? 4'b1011 : 4'b1111;
													assign node35900 = (inp[5]) ? node35914 : node35901;
														assign node35901 = (inp[13]) ? node35909 : node35902;
															assign node35902 = (inp[2]) ? node35906 : node35903;
																assign node35903 = (inp[1]) ? 4'b1110 : 4'b1010;
																assign node35906 = (inp[1]) ? 4'b1010 : 4'b1110;
															assign node35909 = (inp[1]) ? node35911 : 4'b1011;
																assign node35911 = (inp[2]) ? 4'b1111 : 4'b1011;
														assign node35914 = (inp[13]) ? node35920 : node35915;
															assign node35915 = (inp[2]) ? node35917 : 4'b1011;
																assign node35917 = (inp[1]) ? 4'b1110 : 4'b1111;
															assign node35920 = (inp[2]) ? 4'b1010 : 4'b1110;
								assign node35923 = (inp[9]) ? node36273 : node35924;
									assign node35924 = (inp[2]) ? node36088 : node35925;
										assign node35925 = (inp[5]) ? node36015 : node35926;
											assign node35926 = (inp[11]) ? node35966 : node35927;
												assign node35927 = (inp[1]) ? node35951 : node35928;
													assign node35928 = (inp[15]) ? node35944 : node35929;
														assign node35929 = (inp[10]) ? node35937 : node35930;
															assign node35930 = (inp[0]) ? node35934 : node35931;
																assign node35931 = (inp[13]) ? 4'b1001 : 4'b1000;
																assign node35934 = (inp[13]) ? 4'b1000 : 4'b1001;
															assign node35937 = (inp[13]) ? node35941 : node35938;
																assign node35938 = (inp[0]) ? 4'b1000 : 4'b1001;
																assign node35941 = (inp[0]) ? 4'b1001 : 4'b1000;
														assign node35944 = (inp[10]) ? node35948 : node35945;
															assign node35945 = (inp[0]) ? 4'b1101 : 4'b1100;
															assign node35948 = (inp[0]) ? 4'b1100 : 4'b1101;
													assign node35951 = (inp[15]) ? node35959 : node35952;
														assign node35952 = (inp[13]) ? 4'b1100 : node35953;
															assign node35953 = (inp[0]) ? node35955 : 4'b1101;
																assign node35955 = (inp[10]) ? 4'b1101 : 4'b1100;
														assign node35959 = (inp[10]) ? node35963 : node35960;
															assign node35960 = (inp[0]) ? 4'b1001 : 4'b1000;
															assign node35963 = (inp[0]) ? 4'b1000 : 4'b1001;
												assign node35966 = (inp[0]) ? node35984 : node35967;
													assign node35967 = (inp[15]) ? node35975 : node35968;
														assign node35968 = (inp[1]) ? node35972 : node35969;
															assign node35969 = (inp[10]) ? 4'b1001 : 4'b1000;
															assign node35972 = (inp[10]) ? 4'b1100 : 4'b1101;
														assign node35975 = (inp[1]) ? 4'b1000 : node35976;
															assign node35976 = (inp[13]) ? node35980 : node35977;
																assign node35977 = (inp[10]) ? 4'b1101 : 4'b1100;
																assign node35980 = (inp[10]) ? 4'b1100 : 4'b1101;
													assign node35984 = (inp[13]) ? node36000 : node35985;
														assign node35985 = (inp[10]) ? node35993 : node35986;
															assign node35986 = (inp[15]) ? node35990 : node35987;
																assign node35987 = (inp[1]) ? 4'b1100 : 4'b1001;
																assign node35990 = (inp[1]) ? 4'b1001 : 4'b1101;
															assign node35993 = (inp[15]) ? node35997 : node35994;
																assign node35994 = (inp[1]) ? 4'b1101 : 4'b1000;
																assign node35997 = (inp[1]) ? 4'b1000 : 4'b1100;
														assign node36000 = (inp[10]) ? node36008 : node36001;
															assign node36001 = (inp[15]) ? node36005 : node36002;
																assign node36002 = (inp[1]) ? 4'b1100 : 4'b1001;
																assign node36005 = (inp[1]) ? 4'b1000 : 4'b1100;
															assign node36008 = (inp[15]) ? node36012 : node36009;
																assign node36009 = (inp[1]) ? 4'b1101 : 4'b1000;
																assign node36012 = (inp[1]) ? 4'b1001 : 4'b1101;
											assign node36015 = (inp[10]) ? node36055 : node36016;
												assign node36016 = (inp[13]) ? node36032 : node36017;
													assign node36017 = (inp[15]) ? node36027 : node36018;
														assign node36018 = (inp[1]) ? node36024 : node36019;
															assign node36019 = (inp[0]) ? 4'b1100 : node36020;
																assign node36020 = (inp[11]) ? 4'b1100 : 4'b1101;
															assign node36024 = (inp[0]) ? 4'b1001 : 4'b1000;
														assign node36027 = (inp[1]) ? 4'b1101 : node36028;
															assign node36028 = (inp[0]) ? 4'b1000 : 4'b1001;
													assign node36032 = (inp[0]) ? node36046 : node36033;
														assign node36033 = (inp[11]) ? node36041 : node36034;
															assign node36034 = (inp[1]) ? node36038 : node36035;
																assign node36035 = (inp[15]) ? 4'b1001 : 4'b1101;
																assign node36038 = (inp[15]) ? 4'b1100 : 4'b1001;
															assign node36041 = (inp[1]) ? node36043 : 4'b1000;
																assign node36043 = (inp[15]) ? 4'b1100 : 4'b1000;
														assign node36046 = (inp[15]) ? node36052 : node36047;
															assign node36047 = (inp[11]) ? 4'b1001 : node36048;
																assign node36048 = (inp[1]) ? 4'b1000 : 4'b1100;
															assign node36052 = (inp[1]) ? 4'b1101 : 4'b1001;
												assign node36055 = (inp[1]) ? node36073 : node36056;
													assign node36056 = (inp[15]) ? node36066 : node36057;
														assign node36057 = (inp[11]) ? node36061 : node36058;
															assign node36058 = (inp[0]) ? 4'b1101 : 4'b1100;
															assign node36061 = (inp[13]) ? 4'b1100 : node36062;
																assign node36062 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node36066 = (inp[0]) ? 4'b1001 : node36067;
															assign node36067 = (inp[13]) ? node36069 : 4'b1000;
																assign node36069 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node36073 = (inp[15]) ? node36077 : node36074;
														assign node36074 = (inp[0]) ? 4'b1000 : 4'b1001;
														assign node36077 = (inp[0]) ? node36083 : node36078;
															assign node36078 = (inp[11]) ? 4'b1101 : node36079;
																assign node36079 = (inp[13]) ? 4'b1101 : 4'b1100;
															assign node36083 = (inp[13]) ? 4'b1100 : node36084;
																assign node36084 = (inp[11]) ? 4'b1100 : 4'b1101;
										assign node36088 = (inp[0]) ? node36190 : node36089;
											assign node36089 = (inp[11]) ? node36141 : node36090;
												assign node36090 = (inp[13]) ? node36118 : node36091;
													assign node36091 = (inp[1]) ? node36107 : node36092;
														assign node36092 = (inp[10]) ? node36100 : node36093;
															assign node36093 = (inp[5]) ? node36097 : node36094;
																assign node36094 = (inp[15]) ? 4'b1000 : 4'b1100;
																assign node36097 = (inp[15]) ? 4'b1101 : 4'b1001;
															assign node36100 = (inp[5]) ? node36104 : node36101;
																assign node36101 = (inp[15]) ? 4'b1001 : 4'b1101;
																assign node36104 = (inp[15]) ? 4'b1100 : 4'b1000;
														assign node36107 = (inp[5]) ? node36111 : node36108;
															assign node36108 = (inp[15]) ? 4'b1100 : 4'b1000;
															assign node36111 = (inp[15]) ? node36115 : node36112;
																assign node36112 = (inp[10]) ? 4'b1101 : 4'b1100;
																assign node36115 = (inp[10]) ? 4'b1000 : 4'b1001;
													assign node36118 = (inp[10]) ? node36130 : node36119;
														assign node36119 = (inp[15]) ? node36123 : node36120;
															assign node36120 = (inp[1]) ? 4'b1000 : 4'b1001;
															assign node36123 = (inp[1]) ? node36127 : node36124;
																assign node36124 = (inp[5]) ? 4'b1100 : 4'b1000;
																assign node36127 = (inp[5]) ? 4'b1000 : 4'b1101;
														assign node36130 = (inp[1]) ? node36134 : node36131;
															assign node36131 = (inp[15]) ? 4'b1001 : 4'b1000;
															assign node36134 = (inp[5]) ? node36138 : node36135;
																assign node36135 = (inp[15]) ? 4'b1100 : 4'b1001;
																assign node36138 = (inp[15]) ? 4'b1001 : 4'b1101;
												assign node36141 = (inp[15]) ? node36171 : node36142;
													assign node36142 = (inp[10]) ? node36158 : node36143;
														assign node36143 = (inp[13]) ? node36151 : node36144;
															assign node36144 = (inp[5]) ? node36148 : node36145;
																assign node36145 = (inp[1]) ? 4'b1001 : 4'b1101;
																assign node36148 = (inp[1]) ? 4'b1101 : 4'b1000;
															assign node36151 = (inp[1]) ? node36155 : node36152;
																assign node36152 = (inp[5]) ? 4'b1001 : 4'b1100;
																assign node36155 = (inp[5]) ? 4'b1100 : 4'b1001;
														assign node36158 = (inp[13]) ? node36164 : node36159;
															assign node36159 = (inp[5]) ? 4'b1100 : node36160;
																assign node36160 = (inp[1]) ? 4'b1000 : 4'b1100;
															assign node36164 = (inp[1]) ? node36168 : node36165;
																assign node36165 = (inp[5]) ? 4'b1000 : 4'b1101;
																assign node36168 = (inp[5]) ? 4'b1101 : 4'b1000;
													assign node36171 = (inp[10]) ? node36181 : node36172;
														assign node36172 = (inp[5]) ? node36178 : node36173;
															assign node36173 = (inp[1]) ? 4'b1101 : node36174;
																assign node36174 = (inp[13]) ? 4'b1001 : 4'b1000;
															assign node36178 = (inp[1]) ? 4'b1000 : 4'b1100;
														assign node36181 = (inp[5]) ? node36187 : node36182;
															assign node36182 = (inp[1]) ? 4'b1100 : node36183;
																assign node36183 = (inp[13]) ? 4'b1000 : 4'b1001;
															assign node36187 = (inp[1]) ? 4'b1001 : 4'b1101;
											assign node36190 = (inp[10]) ? node36234 : node36191;
												assign node36191 = (inp[11]) ? node36217 : node36192;
													assign node36192 = (inp[13]) ? node36208 : node36193;
														assign node36193 = (inp[5]) ? node36201 : node36194;
															assign node36194 = (inp[15]) ? node36198 : node36195;
																assign node36195 = (inp[1]) ? 4'b1000 : 4'b1101;
																assign node36198 = (inp[1]) ? 4'b1101 : 4'b1001;
															assign node36201 = (inp[15]) ? node36205 : node36202;
																assign node36202 = (inp[1]) ? 4'b1101 : 4'b1000;
																assign node36205 = (inp[1]) ? 4'b1000 : 4'b1100;
														assign node36208 = (inp[5]) ? 4'b1101 : node36209;
															assign node36209 = (inp[15]) ? node36213 : node36210;
																assign node36210 = (inp[1]) ? 4'b1001 : 4'b1101;
																assign node36213 = (inp[1]) ? 4'b1100 : 4'b1001;
													assign node36217 = (inp[5]) ? node36227 : node36218;
														assign node36218 = (inp[1]) ? node36224 : node36219;
															assign node36219 = (inp[15]) ? 4'b1000 : node36220;
																assign node36220 = (inp[13]) ? 4'b1101 : 4'b1100;
															assign node36224 = (inp[15]) ? 4'b1100 : 4'b1000;
														assign node36227 = (inp[15]) ? node36231 : node36228;
															assign node36228 = (inp[1]) ? 4'b1100 : 4'b1000;
															assign node36231 = (inp[1]) ? 4'b1001 : 4'b1101;
												assign node36234 = (inp[15]) ? node36256 : node36235;
													assign node36235 = (inp[11]) ? node36243 : node36236;
														assign node36236 = (inp[5]) ? node36240 : node36237;
															assign node36237 = (inp[1]) ? 4'b1000 : 4'b1100;
															assign node36240 = (inp[1]) ? 4'b1100 : 4'b1001;
														assign node36243 = (inp[1]) ? node36251 : node36244;
															assign node36244 = (inp[5]) ? node36248 : node36245;
																assign node36245 = (inp[13]) ? 4'b1100 : 4'b1101;
																assign node36248 = (inp[13]) ? 4'b1001 : 4'b1000;
															assign node36251 = (inp[5]) ? node36253 : 4'b1001;
																assign node36253 = (inp[13]) ? 4'b1100 : 4'b1101;
													assign node36256 = (inp[5]) ? node36266 : node36257;
														assign node36257 = (inp[1]) ? node36263 : node36258;
															assign node36258 = (inp[13]) ? node36260 : 4'b1000;
																assign node36260 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node36263 = (inp[13]) ? 4'b1101 : 4'b1100;
														assign node36266 = (inp[1]) ? 4'b1000 : node36267;
															assign node36267 = (inp[13]) ? 4'b1100 : node36268;
																assign node36268 = (inp[11]) ? 4'b1100 : 4'b1101;
									assign node36273 = (inp[11]) ? node36447 : node36274;
										assign node36274 = (inp[0]) ? node36362 : node36275;
											assign node36275 = (inp[10]) ? node36321 : node36276;
												assign node36276 = (inp[5]) ? node36302 : node36277;
													assign node36277 = (inp[15]) ? node36291 : node36278;
														assign node36278 = (inp[13]) ? node36284 : node36279;
															assign node36279 = (inp[1]) ? node36281 : 4'b1000;
																assign node36281 = (inp[2]) ? 4'b1001 : 4'b1101;
															assign node36284 = (inp[2]) ? node36288 : node36285;
																assign node36285 = (inp[1]) ? 4'b1100 : 4'b1001;
																assign node36288 = (inp[1]) ? 4'b1000 : 4'b1100;
														assign node36291 = (inp[13]) ? node36297 : node36292;
															assign node36292 = (inp[1]) ? 4'b1100 : node36293;
																assign node36293 = (inp[2]) ? 4'b1000 : 4'b1100;
															assign node36297 = (inp[2]) ? 4'b1101 : node36298;
																assign node36298 = (inp[1]) ? 4'b1000 : 4'b1100;
													assign node36302 = (inp[2]) ? node36312 : node36303;
														assign node36303 = (inp[1]) ? node36307 : node36304;
															assign node36304 = (inp[15]) ? 4'b1001 : 4'b1101;
															assign node36307 = (inp[15]) ? 4'b1101 : node36308;
																assign node36308 = (inp[13]) ? 4'b1001 : 4'b1000;
														assign node36312 = (inp[1]) ? node36316 : node36313;
															assign node36313 = (inp[15]) ? 4'b1100 : 4'b1001;
															assign node36316 = (inp[15]) ? node36318 : 4'b1100;
																assign node36318 = (inp[13]) ? 4'b1000 : 4'b1001;
												assign node36321 = (inp[5]) ? node36341 : node36322;
													assign node36322 = (inp[1]) ? node36330 : node36323;
														assign node36323 = (inp[15]) ? node36327 : node36324;
															assign node36324 = (inp[2]) ? 4'b1101 : 4'b1001;
															assign node36327 = (inp[2]) ? 4'b1001 : 4'b1101;
														assign node36330 = (inp[15]) ? node36336 : node36331;
															assign node36331 = (inp[13]) ? 4'b1001 : node36332;
																assign node36332 = (inp[2]) ? 4'b1000 : 4'b1100;
															assign node36336 = (inp[2]) ? node36338 : 4'b1001;
																assign node36338 = (inp[13]) ? 4'b1100 : 4'b1101;
													assign node36341 = (inp[1]) ? node36351 : node36342;
														assign node36342 = (inp[2]) ? node36346 : node36343;
															assign node36343 = (inp[15]) ? 4'b1000 : 4'b1100;
															assign node36346 = (inp[15]) ? node36348 : 4'b1000;
																assign node36348 = (inp[13]) ? 4'b1101 : 4'b1100;
														assign node36351 = (inp[15]) ? node36357 : node36352;
															assign node36352 = (inp[2]) ? 4'b1101 : node36353;
																assign node36353 = (inp[13]) ? 4'b1000 : 4'b1001;
															assign node36357 = (inp[13]) ? node36359 : 4'b1000;
																assign node36359 = (inp[2]) ? 4'b1001 : 4'b1101;
											assign node36362 = (inp[10]) ? node36404 : node36363;
												assign node36363 = (inp[5]) ? node36383 : node36364;
													assign node36364 = (inp[1]) ? node36372 : node36365;
														assign node36365 = (inp[2]) ? node36369 : node36366;
															assign node36366 = (inp[15]) ? 4'b1101 : 4'b1001;
															assign node36369 = (inp[15]) ? 4'b1001 : 4'b1101;
														assign node36372 = (inp[15]) ? node36380 : node36373;
															assign node36373 = (inp[13]) ? node36377 : node36374;
																assign node36374 = (inp[2]) ? 4'b1000 : 4'b1100;
																assign node36377 = (inp[2]) ? 4'b1001 : 4'b1101;
															assign node36380 = (inp[13]) ? 4'b1100 : 4'b1101;
													assign node36383 = (inp[1]) ? node36395 : node36384;
														assign node36384 = (inp[13]) ? node36390 : node36385;
															assign node36385 = (inp[15]) ? node36387 : 4'b1100;
																assign node36387 = (inp[2]) ? 4'b1100 : 4'b1000;
															assign node36390 = (inp[15]) ? 4'b1101 : node36391;
																assign node36391 = (inp[2]) ? 4'b1000 : 4'b1100;
														assign node36395 = (inp[15]) ? node36399 : node36396;
															assign node36396 = (inp[2]) ? 4'b1101 : 4'b1001;
															assign node36399 = (inp[2]) ? 4'b1001 : node36400;
																assign node36400 = (inp[13]) ? 4'b1101 : 4'b1100;
												assign node36404 = (inp[5]) ? node36428 : node36405;
													assign node36405 = (inp[15]) ? node36419 : node36406;
														assign node36406 = (inp[13]) ? node36414 : node36407;
															assign node36407 = (inp[1]) ? node36411 : node36408;
																assign node36408 = (inp[2]) ? 4'b1100 : 4'b1000;
																assign node36411 = (inp[2]) ? 4'b1001 : 4'b1101;
															assign node36414 = (inp[1]) ? node36416 : 4'b1001;
																assign node36416 = (inp[2]) ? 4'b1000 : 4'b1100;
														assign node36419 = (inp[1]) ? node36423 : node36420;
															assign node36420 = (inp[2]) ? 4'b1000 : 4'b1100;
															assign node36423 = (inp[2]) ? node36425 : 4'b1000;
																assign node36425 = (inp[13]) ? 4'b1101 : 4'b1100;
													assign node36428 = (inp[1]) ? node36436 : node36429;
														assign node36429 = (inp[2]) ? node36433 : node36430;
															assign node36430 = (inp[15]) ? 4'b1001 : 4'b1101;
															assign node36433 = (inp[15]) ? 4'b1100 : 4'b1001;
														assign node36436 = (inp[2]) ? node36442 : node36437;
															assign node36437 = (inp[15]) ? node36439 : 4'b1001;
																assign node36439 = (inp[13]) ? 4'b1100 : 4'b1101;
															assign node36442 = (inp[15]) ? node36444 : 4'b1100;
																assign node36444 = (inp[13]) ? 4'b1000 : 4'b1001;
										assign node36447 = (inp[15]) ? node36535 : node36448;
											assign node36448 = (inp[1]) ? node36488 : node36449;
												assign node36449 = (inp[2]) ? node36467 : node36450;
													assign node36450 = (inp[5]) ? node36458 : node36451;
														assign node36451 = (inp[0]) ? node36455 : node36452;
															assign node36452 = (inp[10]) ? 4'b1001 : 4'b1000;
															assign node36455 = (inp[10]) ? 4'b1000 : 4'b1001;
														assign node36458 = (inp[0]) ? node36460 : 4'b1100;
															assign node36460 = (inp[10]) ? node36464 : node36461;
																assign node36461 = (inp[13]) ? 4'b1100 : 4'b1101;
																assign node36464 = (inp[13]) ? 4'b1101 : 4'b1100;
													assign node36467 = (inp[5]) ? node36475 : node36468;
														assign node36468 = (inp[0]) ? 4'b1100 : node36469;
															assign node36469 = (inp[13]) ? node36471 : 4'b1101;
																assign node36471 = (inp[10]) ? 4'b1101 : 4'b1100;
														assign node36475 = (inp[0]) ? node36481 : node36476;
															assign node36476 = (inp[10]) ? 4'b1001 : node36477;
																assign node36477 = (inp[13]) ? 4'b1001 : 4'b1000;
															assign node36481 = (inp[13]) ? node36485 : node36482;
																assign node36482 = (inp[10]) ? 4'b1000 : 4'b1001;
																assign node36485 = (inp[10]) ? 4'b1001 : 4'b1000;
												assign node36488 = (inp[5]) ? node36506 : node36489;
													assign node36489 = (inp[2]) ? node36497 : node36490;
														assign node36490 = (inp[0]) ? node36494 : node36491;
															assign node36491 = (inp[10]) ? 4'b1100 : 4'b1101;
															assign node36494 = (inp[10]) ? 4'b1101 : 4'b1100;
														assign node36497 = (inp[13]) ? node36499 : 4'b1000;
															assign node36499 = (inp[10]) ? node36503 : node36500;
																assign node36500 = (inp[0]) ? 4'b1000 : 4'b1001;
																assign node36503 = (inp[0]) ? 4'b1001 : 4'b1000;
													assign node36506 = (inp[2]) ? node36520 : node36507;
														assign node36507 = (inp[13]) ? node36515 : node36508;
															assign node36508 = (inp[10]) ? node36512 : node36509;
																assign node36509 = (inp[0]) ? 4'b1001 : 4'b1000;
																assign node36512 = (inp[0]) ? 4'b1000 : 4'b1001;
															assign node36515 = (inp[0]) ? node36517 : 4'b1000;
																assign node36517 = (inp[10]) ? 4'b1000 : 4'b1001;
														assign node36520 = (inp[0]) ? node36528 : node36521;
															assign node36521 = (inp[13]) ? node36525 : node36522;
																assign node36522 = (inp[10]) ? 4'b1100 : 4'b1101;
																assign node36525 = (inp[10]) ? 4'b1101 : 4'b1100;
															assign node36528 = (inp[13]) ? node36532 : node36529;
																assign node36529 = (inp[10]) ? 4'b1101 : 4'b1100;
																assign node36532 = (inp[10]) ? 4'b1100 : 4'b1101;
											assign node36535 = (inp[1]) ? node36577 : node36536;
												assign node36536 = (inp[0]) ? node36560 : node36537;
													assign node36537 = (inp[5]) ? node36551 : node36538;
														assign node36538 = (inp[2]) ? node36546 : node36539;
															assign node36539 = (inp[13]) ? node36543 : node36540;
																assign node36540 = (inp[10]) ? 4'b1101 : 4'b1100;
																assign node36543 = (inp[10]) ? 4'b1100 : 4'b1101;
															assign node36546 = (inp[10]) ? 4'b1001 : node36547;
																assign node36547 = (inp[13]) ? 4'b1001 : 4'b1000;
														assign node36551 = (inp[2]) ? node36557 : node36552;
															assign node36552 = (inp[13]) ? 4'b1000 : node36553;
																assign node36553 = (inp[10]) ? 4'b1000 : 4'b1001;
															assign node36557 = (inp[10]) ? 4'b1101 : 4'b1100;
													assign node36560 = (inp[10]) ? node36568 : node36561;
														assign node36561 = (inp[5]) ? node36565 : node36562;
															assign node36562 = (inp[13]) ? 4'b1100 : 4'b1101;
															assign node36565 = (inp[2]) ? 4'b1101 : 4'b1001;
														assign node36568 = (inp[5]) ? node36574 : node36569;
															assign node36569 = (inp[2]) ? node36571 : 4'b1100;
																assign node36571 = (inp[13]) ? 4'b1001 : 4'b1000;
															assign node36574 = (inp[2]) ? 4'b1100 : 4'b1001;
												assign node36577 = (inp[13]) ? node36605 : node36578;
													assign node36578 = (inp[2]) ? node36590 : node36579;
														assign node36579 = (inp[5]) ? node36585 : node36580;
															assign node36580 = (inp[10]) ? 4'b1001 : node36581;
																assign node36581 = (inp[0]) ? 4'b1001 : 4'b1000;
															assign node36585 = (inp[0]) ? 4'b1101 : node36586;
																assign node36586 = (inp[10]) ? 4'b1101 : 4'b1100;
														assign node36590 = (inp[5]) ? node36598 : node36591;
															assign node36591 = (inp[10]) ? node36595 : node36592;
																assign node36592 = (inp[0]) ? 4'b1100 : 4'b1101;
																assign node36595 = (inp[0]) ? 4'b1101 : 4'b1100;
															assign node36598 = (inp[0]) ? node36602 : node36599;
																assign node36599 = (inp[10]) ? 4'b1001 : 4'b1000;
																assign node36602 = (inp[10]) ? 4'b1000 : 4'b1001;
													assign node36605 = (inp[5]) ? node36621 : node36606;
														assign node36606 = (inp[2]) ? node36614 : node36607;
															assign node36607 = (inp[10]) ? node36611 : node36608;
																assign node36608 = (inp[0]) ? 4'b1000 : 4'b1001;
																assign node36611 = (inp[0]) ? 4'b1001 : 4'b1000;
															assign node36614 = (inp[10]) ? node36618 : node36615;
																assign node36615 = (inp[0]) ? 4'b1100 : 4'b1101;
																assign node36618 = (inp[0]) ? 4'b1101 : 4'b1100;
														assign node36621 = (inp[2]) ? node36629 : node36622;
															assign node36622 = (inp[0]) ? node36626 : node36623;
																assign node36623 = (inp[10]) ? 4'b1101 : 4'b1100;
																assign node36626 = (inp[10]) ? 4'b1100 : 4'b1101;
															assign node36629 = (inp[10]) ? node36633 : node36630;
																assign node36630 = (inp[0]) ? 4'b1001 : 4'b1000;
																assign node36633 = (inp[0]) ? 4'b1000 : 4'b1001;
							assign node36636 = (inp[15]) ? node37106 : node36637;
								assign node36637 = (inp[13]) ? node36889 : node36638;
									assign node36638 = (inp[2]) ? node36778 : node36639;
										assign node36639 = (inp[8]) ? node36715 : node36640;
											assign node36640 = (inp[1]) ? node36692 : node36641;
												assign node36641 = (inp[5]) ? node36671 : node36642;
													assign node36642 = (inp[11]) ? node36658 : node36643;
														assign node36643 = (inp[0]) ? node36651 : node36644;
															assign node36644 = (inp[10]) ? node36648 : node36645;
																assign node36645 = (inp[9]) ? 4'b1000 : 4'b1001;
																assign node36648 = (inp[9]) ? 4'b1001 : 4'b1000;
															assign node36651 = (inp[9]) ? node36655 : node36652;
																assign node36652 = (inp[10]) ? 4'b1000 : 4'b1001;
																assign node36655 = (inp[10]) ? 4'b1001 : 4'b1000;
														assign node36658 = (inp[9]) ? node36664 : node36659;
															assign node36659 = (inp[10]) ? 4'b1000 : node36660;
																assign node36660 = (inp[0]) ? 4'b1001 : 4'b1000;
															assign node36664 = (inp[10]) ? node36668 : node36665;
																assign node36665 = (inp[0]) ? 4'b1000 : 4'b1001;
																assign node36668 = (inp[0]) ? 4'b1001 : 4'b1000;
													assign node36671 = (inp[0]) ? node36679 : node36672;
														assign node36672 = (inp[9]) ? node36676 : node36673;
															assign node36673 = (inp[10]) ? 4'b1101 : 4'b1100;
															assign node36676 = (inp[10]) ? 4'b1100 : 4'b1101;
														assign node36679 = (inp[11]) ? node36685 : node36680;
															assign node36680 = (inp[10]) ? 4'b1101 : node36681;
																assign node36681 = (inp[9]) ? 4'b1100 : 4'b1101;
															assign node36685 = (inp[9]) ? node36689 : node36686;
																assign node36686 = (inp[10]) ? 4'b1101 : 4'b1100;
																assign node36689 = (inp[10]) ? 4'b1100 : 4'b1101;
												assign node36692 = (inp[10]) ? node36704 : node36693;
													assign node36693 = (inp[9]) ? node36699 : node36694;
														assign node36694 = (inp[0]) ? 4'b1000 : node36695;
															assign node36695 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node36699 = (inp[11]) ? node36701 : 4'b1001;
															assign node36701 = (inp[0]) ? 4'b1001 : 4'b1000;
													assign node36704 = (inp[9]) ? node36710 : node36705;
														assign node36705 = (inp[0]) ? 4'b1001 : node36706;
															assign node36706 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node36710 = (inp[0]) ? 4'b1000 : node36711;
															assign node36711 = (inp[11]) ? 4'b1001 : 4'b1000;
											assign node36715 = (inp[1]) ? node36747 : node36716;
												assign node36716 = (inp[11]) ? node36724 : node36717;
													assign node36717 = (inp[0]) ? node36721 : node36718;
														assign node36718 = (inp[10]) ? 4'b1000 : 4'b1001;
														assign node36721 = (inp[10]) ? 4'b1001 : 4'b1000;
													assign node36724 = (inp[9]) ? node36740 : node36725;
														assign node36725 = (inp[5]) ? node36733 : node36726;
															assign node36726 = (inp[0]) ? node36730 : node36727;
																assign node36727 = (inp[10]) ? 4'b1001 : 4'b1000;
																assign node36730 = (inp[10]) ? 4'b1000 : 4'b1001;
															assign node36733 = (inp[0]) ? node36737 : node36734;
																assign node36734 = (inp[10]) ? 4'b1001 : 4'b1000;
																assign node36737 = (inp[10]) ? 4'b1000 : 4'b1001;
														assign node36740 = (inp[0]) ? node36744 : node36741;
															assign node36741 = (inp[10]) ? 4'b1001 : 4'b1000;
															assign node36744 = (inp[10]) ? 4'b1000 : 4'b1001;
												assign node36747 = (inp[9]) ? node36763 : node36748;
													assign node36748 = (inp[11]) ? node36756 : node36749;
														assign node36749 = (inp[10]) ? node36753 : node36750;
															assign node36750 = (inp[0]) ? 4'b1101 : 4'b1100;
															assign node36753 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node36756 = (inp[10]) ? node36760 : node36757;
															assign node36757 = (inp[0]) ? 4'b1100 : 4'b1101;
															assign node36760 = (inp[0]) ? 4'b1101 : 4'b1100;
													assign node36763 = (inp[10]) ? node36771 : node36764;
														assign node36764 = (inp[0]) ? node36768 : node36765;
															assign node36765 = (inp[11]) ? 4'b1101 : 4'b1100;
															assign node36768 = (inp[11]) ? 4'b1100 : 4'b1101;
														assign node36771 = (inp[0]) ? node36775 : node36772;
															assign node36772 = (inp[11]) ? 4'b1100 : 4'b1101;
															assign node36775 = (inp[11]) ? 4'b1101 : 4'b1100;
										assign node36778 = (inp[8]) ? node36842 : node36779;
											assign node36779 = (inp[1]) ? node36821 : node36780;
												assign node36780 = (inp[5]) ? node36800 : node36781;
													assign node36781 = (inp[10]) ? node36791 : node36782;
														assign node36782 = (inp[9]) ? node36788 : node36783;
															assign node36783 = (inp[11]) ? 4'b1100 : node36784;
																assign node36784 = (inp[0]) ? 4'b1101 : 4'b1100;
															assign node36788 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node36791 = (inp[9]) ? node36797 : node36792;
															assign node36792 = (inp[0]) ? node36794 : 4'b1101;
																assign node36794 = (inp[11]) ? 4'b1101 : 4'b1100;
															assign node36797 = (inp[0]) ? 4'b1101 : 4'b1100;
													assign node36800 = (inp[10]) ? node36812 : node36801;
														assign node36801 = (inp[9]) ? node36807 : node36802;
															assign node36802 = (inp[11]) ? 4'b1000 : node36803;
																assign node36803 = (inp[0]) ? 4'b1001 : 4'b1000;
															assign node36807 = (inp[0]) ? node36809 : 4'b1001;
																assign node36809 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node36812 = (inp[0]) ? node36814 : 4'b1001;
															assign node36814 = (inp[11]) ? node36818 : node36815;
																assign node36815 = (inp[9]) ? 4'b1001 : 4'b1000;
																assign node36818 = (inp[9]) ? 4'b1000 : 4'b1001;
												assign node36821 = (inp[10]) ? node36833 : node36822;
													assign node36822 = (inp[9]) ? node36828 : node36823;
														assign node36823 = (inp[11]) ? 4'b1101 : node36824;
															assign node36824 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node36828 = (inp[11]) ? 4'b1100 : node36829;
															assign node36829 = (inp[0]) ? 4'b1101 : 4'b1100;
													assign node36833 = (inp[9]) ? node36839 : node36834;
														assign node36834 = (inp[0]) ? node36836 : 4'b1100;
															assign node36836 = (inp[11]) ? 4'b1100 : 4'b1101;
														assign node36839 = (inp[0]) ? 4'b1100 : 4'b1101;
											assign node36842 = (inp[1]) ? node36866 : node36843;
												assign node36843 = (inp[11]) ? node36859 : node36844;
													assign node36844 = (inp[9]) ? node36852 : node36845;
														assign node36845 = (inp[10]) ? node36849 : node36846;
															assign node36846 = (inp[0]) ? 4'b1101 : 4'b1100;
															assign node36849 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node36852 = (inp[0]) ? node36856 : node36853;
															assign node36853 = (inp[10]) ? 4'b1101 : 4'b1100;
															assign node36856 = (inp[10]) ? 4'b1100 : 4'b1101;
													assign node36859 = (inp[10]) ? node36863 : node36860;
														assign node36860 = (inp[0]) ? 4'b1101 : 4'b1100;
														assign node36863 = (inp[0]) ? 4'b1100 : 4'b1101;
												assign node36866 = (inp[0]) ? node36874 : node36867;
													assign node36867 = (inp[11]) ? node36871 : node36868;
														assign node36868 = (inp[10]) ? 4'b1001 : 4'b1000;
														assign node36871 = (inp[10]) ? 4'b1000 : 4'b1001;
													assign node36874 = (inp[5]) ? node36882 : node36875;
														assign node36875 = (inp[11]) ? node36879 : node36876;
															assign node36876 = (inp[10]) ? 4'b1000 : 4'b1001;
															assign node36879 = (inp[10]) ? 4'b1001 : 4'b1000;
														assign node36882 = (inp[10]) ? node36886 : node36883;
															assign node36883 = (inp[11]) ? 4'b1000 : 4'b1001;
															assign node36886 = (inp[11]) ? 4'b1001 : 4'b1000;
									assign node36889 = (inp[2]) ? node36999 : node36890;
										assign node36890 = (inp[1]) ? node36962 : node36891;
											assign node36891 = (inp[8]) ? node36929 : node36892;
												assign node36892 = (inp[5]) ? node36906 : node36893;
													assign node36893 = (inp[10]) ? node36899 : node36894;
														assign node36894 = (inp[9]) ? node36896 : 4'b1101;
															assign node36896 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node36899 = (inp[9]) ? node36901 : 4'b1100;
															assign node36901 = (inp[0]) ? 4'b1101 : node36902;
																assign node36902 = (inp[11]) ? 4'b1100 : 4'b1101;
													assign node36906 = (inp[0]) ? node36922 : node36907;
														assign node36907 = (inp[10]) ? node36915 : node36908;
															assign node36908 = (inp[9]) ? node36912 : node36909;
																assign node36909 = (inp[11]) ? 4'b1000 : 4'b1001;
																assign node36912 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node36915 = (inp[9]) ? node36919 : node36916;
																assign node36916 = (inp[11]) ? 4'b1001 : 4'b1000;
																assign node36919 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node36922 = (inp[9]) ? node36926 : node36923;
															assign node36923 = (inp[10]) ? 4'b1000 : 4'b1001;
															assign node36926 = (inp[10]) ? 4'b1001 : 4'b1000;
												assign node36929 = (inp[5]) ? node36937 : node36930;
													assign node36930 = (inp[0]) ? node36934 : node36931;
														assign node36931 = (inp[10]) ? 4'b1000 : 4'b1001;
														assign node36934 = (inp[10]) ? 4'b1001 : 4'b1000;
													assign node36937 = (inp[9]) ? node36947 : node36938;
														assign node36938 = (inp[11]) ? node36940 : 4'b1000;
															assign node36940 = (inp[0]) ? node36944 : node36941;
																assign node36941 = (inp[10]) ? 4'b1000 : 4'b1001;
																assign node36944 = (inp[10]) ? 4'b1001 : 4'b1000;
														assign node36947 = (inp[11]) ? node36955 : node36948;
															assign node36948 = (inp[0]) ? node36952 : node36949;
																assign node36949 = (inp[10]) ? 4'b1000 : 4'b1001;
																assign node36952 = (inp[10]) ? 4'b1001 : 4'b1000;
															assign node36955 = (inp[0]) ? node36959 : node36956;
																assign node36956 = (inp[10]) ? 4'b1000 : 4'b1001;
																assign node36959 = (inp[10]) ? 4'b1001 : 4'b1000;
											assign node36962 = (inp[9]) ? node36986 : node36963;
												assign node36963 = (inp[10]) ? node36973 : node36964;
													assign node36964 = (inp[0]) ? node36970 : node36965;
														assign node36965 = (inp[8]) ? 4'b1100 : node36966;
															assign node36966 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node36970 = (inp[8]) ? 4'b1101 : 4'b1100;
													assign node36973 = (inp[11]) ? node36979 : node36974;
														assign node36974 = (inp[0]) ? node36976 : 4'b1101;
															assign node36976 = (inp[8]) ? 4'b1100 : 4'b1101;
														assign node36979 = (inp[8]) ? node36983 : node36980;
															assign node36980 = (inp[0]) ? 4'b1101 : 4'b1100;
															assign node36983 = (inp[0]) ? 4'b1100 : 4'b1101;
												assign node36986 = (inp[10]) ? node36994 : node36987;
													assign node36987 = (inp[0]) ? 4'b1101 : node36988;
														assign node36988 = (inp[8]) ? 4'b1100 : node36989;
															assign node36989 = (inp[11]) ? 4'b1100 : 4'b1101;
													assign node36994 = (inp[0]) ? 4'b1100 : node36995;
														assign node36995 = (inp[11]) ? 4'b1101 : 4'b1100;
										assign node36999 = (inp[1]) ? node37067 : node37000;
											assign node37000 = (inp[5]) ? node37032 : node37001;
												assign node37001 = (inp[8]) ? node37017 : node37002;
													assign node37002 = (inp[11]) ? node37010 : node37003;
														assign node37003 = (inp[10]) ? node37007 : node37004;
															assign node37004 = (inp[9]) ? 4'b1000 : 4'b1001;
															assign node37007 = (inp[9]) ? 4'b1001 : 4'b1000;
														assign node37010 = (inp[10]) ? 4'b1001 : node37011;
															assign node37011 = (inp[0]) ? 4'b1000 : node37012;
																assign node37012 = (inp[9]) ? 4'b1001 : 4'b1000;
													assign node37017 = (inp[0]) ? node37025 : node37018;
														assign node37018 = (inp[10]) ? node37022 : node37019;
															assign node37019 = (inp[11]) ? 4'b1100 : 4'b1101;
															assign node37022 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node37025 = (inp[11]) ? node37029 : node37026;
															assign node37026 = (inp[10]) ? 4'b1101 : 4'b1100;
															assign node37029 = (inp[10]) ? 4'b1100 : 4'b1101;
												assign node37032 = (inp[0]) ? node37044 : node37033;
													assign node37033 = (inp[10]) ? node37035 : 4'b1100;
														assign node37035 = (inp[11]) ? node37039 : node37036;
															assign node37036 = (inp[8]) ? 4'b1100 : 4'b1101;
															assign node37039 = (inp[9]) ? node37041 : 4'b1101;
																assign node37041 = (inp[8]) ? 4'b1101 : 4'b1100;
													assign node37044 = (inp[8]) ? node37060 : node37045;
														assign node37045 = (inp[9]) ? node37053 : node37046;
															assign node37046 = (inp[10]) ? node37050 : node37047;
																assign node37047 = (inp[11]) ? 4'b1100 : 4'b1101;
																assign node37050 = (inp[11]) ? 4'b1101 : 4'b1100;
															assign node37053 = (inp[11]) ? node37057 : node37054;
																assign node37054 = (inp[10]) ? 4'b1101 : 4'b1100;
																assign node37057 = (inp[10]) ? 4'b1100 : 4'b1101;
														assign node37060 = (inp[10]) ? node37064 : node37061;
															assign node37061 = (inp[11]) ? 4'b1101 : 4'b1100;
															assign node37064 = (inp[11]) ? 4'b1100 : 4'b1101;
											assign node37067 = (inp[9]) ? node37091 : node37068;
												assign node37068 = (inp[10]) ? node37082 : node37069;
													assign node37069 = (inp[11]) ? node37075 : node37070;
														assign node37070 = (inp[0]) ? node37072 : 4'b1000;
															assign node37072 = (inp[8]) ? 4'b1001 : 4'b1000;
														assign node37075 = (inp[0]) ? node37079 : node37076;
															assign node37076 = (inp[8]) ? 4'b1000 : 4'b1001;
															assign node37079 = (inp[8]) ? 4'b1001 : 4'b1000;
													assign node37082 = (inp[8]) ? node37088 : node37083;
														assign node37083 = (inp[0]) ? 4'b1001 : node37084;
															assign node37084 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node37088 = (inp[0]) ? 4'b1000 : 4'b1001;
												assign node37091 = (inp[10]) ? node37099 : node37092;
													assign node37092 = (inp[0]) ? 4'b1001 : node37093;
														assign node37093 = (inp[8]) ? 4'b1000 : node37094;
															assign node37094 = (inp[11]) ? 4'b1000 : 4'b1001;
													assign node37099 = (inp[0]) ? 4'b1000 : node37100;
														assign node37100 = (inp[8]) ? 4'b1001 : node37101;
															assign node37101 = (inp[11]) ? 4'b1001 : 4'b1000;
								assign node37106 = (inp[2]) ? node37332 : node37107;
									assign node37107 = (inp[1]) ? node37251 : node37108;
										assign node37108 = (inp[8]) ? node37210 : node37109;
											assign node37109 = (inp[5]) ? node37161 : node37110;
												assign node37110 = (inp[13]) ? node37138 : node37111;
													assign node37111 = (inp[0]) ? node37125 : node37112;
														assign node37112 = (inp[11]) ? node37118 : node37113;
															assign node37113 = (inp[9]) ? node37115 : 4'b1000;
																assign node37115 = (inp[10]) ? 4'b1001 : 4'b1000;
															assign node37118 = (inp[10]) ? node37122 : node37119;
																assign node37119 = (inp[9]) ? 4'b1000 : 4'b1001;
																assign node37122 = (inp[9]) ? 4'b1001 : 4'b1000;
														assign node37125 = (inp[9]) ? node37131 : node37126;
															assign node37126 = (inp[10]) ? 4'b1001 : node37127;
																assign node37127 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node37131 = (inp[10]) ? node37135 : node37132;
																assign node37132 = (inp[11]) ? 4'b1000 : 4'b1001;
																assign node37135 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node37138 = (inp[10]) ? node37150 : node37139;
														assign node37139 = (inp[9]) ? node37145 : node37140;
															assign node37140 = (inp[0]) ? node37142 : 4'b1100;
																assign node37142 = (inp[11]) ? 4'b1100 : 4'b1101;
															assign node37145 = (inp[11]) ? 4'b1101 : node37146;
																assign node37146 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node37150 = (inp[9]) ? node37156 : node37151;
															assign node37151 = (inp[11]) ? 4'b1101 : node37152;
																assign node37152 = (inp[0]) ? 4'b1100 : 4'b1101;
															assign node37156 = (inp[11]) ? 4'b1100 : node37157;
																assign node37157 = (inp[0]) ? 4'b1101 : 4'b1100;
												assign node37161 = (inp[13]) ? node37179 : node37162;
													assign node37162 = (inp[10]) ? node37174 : node37163;
														assign node37163 = (inp[9]) ? node37169 : node37164;
															assign node37164 = (inp[11]) ? node37166 : 4'b1101;
																assign node37166 = (inp[0]) ? 4'b1101 : 4'b1100;
															assign node37169 = (inp[0]) ? 4'b1100 : node37170;
																assign node37170 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node37174 = (inp[9]) ? node37176 : 4'b1100;
															assign node37176 = (inp[11]) ? 4'b1100 : 4'b1101;
													assign node37179 = (inp[11]) ? node37195 : node37180;
														assign node37180 = (inp[10]) ? node37188 : node37181;
															assign node37181 = (inp[0]) ? node37185 : node37182;
																assign node37182 = (inp[9]) ? 4'b1001 : 4'b1000;
																assign node37185 = (inp[9]) ? 4'b1000 : 4'b1001;
															assign node37188 = (inp[9]) ? node37192 : node37189;
																assign node37189 = (inp[0]) ? 4'b1000 : 4'b1001;
																assign node37192 = (inp[0]) ? 4'b1001 : 4'b1000;
														assign node37195 = (inp[0]) ? node37203 : node37196;
															assign node37196 = (inp[10]) ? node37200 : node37197;
																assign node37197 = (inp[9]) ? 4'b1001 : 4'b1000;
																assign node37200 = (inp[9]) ? 4'b1000 : 4'b1001;
															assign node37203 = (inp[10]) ? node37207 : node37204;
																assign node37204 = (inp[9]) ? 4'b1001 : 4'b1000;
																assign node37207 = (inp[9]) ? 4'b1000 : 4'b1001;
											assign node37210 = (inp[13]) ? node37218 : node37211;
												assign node37211 = (inp[0]) ? node37215 : node37212;
													assign node37212 = (inp[10]) ? 4'b1000 : 4'b1001;
													assign node37215 = (inp[10]) ? 4'b1001 : 4'b1000;
												assign node37218 = (inp[0]) ? node37242 : node37219;
													assign node37219 = (inp[5]) ? node37227 : node37220;
														assign node37220 = (inp[11]) ? node37224 : node37221;
															assign node37221 = (inp[10]) ? 4'b1000 : 4'b1001;
															assign node37224 = (inp[10]) ? 4'b1001 : 4'b1000;
														assign node37227 = (inp[9]) ? node37235 : node37228;
															assign node37228 = (inp[10]) ? node37232 : node37229;
																assign node37229 = (inp[11]) ? 4'b1000 : 4'b1001;
																assign node37232 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node37235 = (inp[10]) ? node37239 : node37236;
																assign node37236 = (inp[11]) ? 4'b1000 : 4'b1001;
																assign node37239 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node37242 = (inp[9]) ? 4'b1000 : node37243;
														assign node37243 = (inp[11]) ? node37247 : node37244;
															assign node37244 = (inp[10]) ? 4'b1001 : 4'b1000;
															assign node37247 = (inp[10]) ? 4'b1000 : 4'b1001;
										assign node37251 = (inp[8]) ? node37309 : node37252;
											assign node37252 = (inp[13]) ? node37276 : node37253;
												assign node37253 = (inp[9]) ? node37265 : node37254;
													assign node37254 = (inp[10]) ? node37260 : node37255;
														assign node37255 = (inp[0]) ? 4'b1001 : node37256;
															assign node37256 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node37260 = (inp[0]) ? 4'b1000 : node37261;
															assign node37261 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node37265 = (inp[10]) ? node37271 : node37266;
														assign node37266 = (inp[0]) ? 4'b1000 : node37267;
															assign node37267 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node37271 = (inp[11]) ? node37273 : 4'b1001;
															assign node37273 = (inp[0]) ? 4'b1001 : 4'b1000;
												assign node37276 = (inp[0]) ? node37294 : node37277;
													assign node37277 = (inp[10]) ? node37285 : node37278;
														assign node37278 = (inp[5]) ? 4'b1101 : node37279;
															assign node37279 = (inp[9]) ? 4'b1101 : node37280;
																assign node37280 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node37285 = (inp[5]) ? node37289 : node37286;
															assign node37286 = (inp[9]) ? 4'b1101 : 4'b1100;
															assign node37289 = (inp[9]) ? node37291 : 4'b1101;
																assign node37291 = (inp[11]) ? 4'b1101 : 4'b1100;
													assign node37294 = (inp[11]) ? node37302 : node37295;
														assign node37295 = (inp[9]) ? node37299 : node37296;
															assign node37296 = (inp[10]) ? 4'b1101 : 4'b1100;
															assign node37299 = (inp[10]) ? 4'b1100 : 4'b1101;
														assign node37302 = (inp[9]) ? node37306 : node37303;
															assign node37303 = (inp[10]) ? 4'b1101 : 4'b1100;
															assign node37306 = (inp[10]) ? 4'b1100 : 4'b1101;
											assign node37309 = (inp[0]) ? node37321 : node37310;
												assign node37310 = (inp[10]) ? node37316 : node37311;
													assign node37311 = (inp[13]) ? 4'b1100 : node37312;
														assign node37312 = (inp[11]) ? 4'b1100 : 4'b1101;
													assign node37316 = (inp[13]) ? 4'b1101 : node37317;
														assign node37317 = (inp[11]) ? 4'b1101 : 4'b1100;
												assign node37321 = (inp[10]) ? node37327 : node37322;
													assign node37322 = (inp[11]) ? 4'b1101 : node37323;
														assign node37323 = (inp[13]) ? 4'b1101 : 4'b1100;
													assign node37327 = (inp[11]) ? 4'b1100 : node37328;
														assign node37328 = (inp[13]) ? 4'b1100 : 4'b1101;
									assign node37332 = (inp[1]) ? node37498 : node37333;
										assign node37333 = (inp[8]) ? node37431 : node37334;
											assign node37334 = (inp[11]) ? node37384 : node37335;
												assign node37335 = (inp[0]) ? node37361 : node37336;
													assign node37336 = (inp[5]) ? node37352 : node37337;
														assign node37337 = (inp[13]) ? node37345 : node37338;
															assign node37338 = (inp[10]) ? node37342 : node37339;
																assign node37339 = (inp[9]) ? 4'b1100 : 4'b1101;
																assign node37342 = (inp[9]) ? 4'b1101 : 4'b1100;
															assign node37345 = (inp[9]) ? node37349 : node37346;
																assign node37346 = (inp[10]) ? 4'b1001 : 4'b1000;
																assign node37349 = (inp[10]) ? 4'b1000 : 4'b1001;
														assign node37352 = (inp[13]) ? 4'b1101 : node37353;
															assign node37353 = (inp[9]) ? node37357 : node37354;
																assign node37354 = (inp[10]) ? 4'b1000 : 4'b1001;
																assign node37357 = (inp[10]) ? 4'b1001 : 4'b1000;
													assign node37361 = (inp[9]) ? node37371 : node37362;
														assign node37362 = (inp[10]) ? 4'b1101 : node37363;
															assign node37363 = (inp[5]) ? node37367 : node37364;
																assign node37364 = (inp[13]) ? 4'b1001 : 4'b1101;
																assign node37367 = (inp[13]) ? 4'b1100 : 4'b1001;
														assign node37371 = (inp[10]) ? node37377 : node37372;
															assign node37372 = (inp[13]) ? 4'b1101 : node37373;
																assign node37373 = (inp[5]) ? 4'b1000 : 4'b1100;
															assign node37377 = (inp[13]) ? node37381 : node37378;
																assign node37378 = (inp[5]) ? 4'b1001 : 4'b1101;
																assign node37381 = (inp[5]) ? 4'b1100 : 4'b1001;
												assign node37384 = (inp[9]) ? node37414 : node37385;
													assign node37385 = (inp[10]) ? node37401 : node37386;
														assign node37386 = (inp[0]) ? node37394 : node37387;
															assign node37387 = (inp[5]) ? node37391 : node37388;
																assign node37388 = (inp[13]) ? 4'b1000 : 4'b1100;
																assign node37391 = (inp[13]) ? 4'b1101 : 4'b1000;
															assign node37394 = (inp[13]) ? node37398 : node37395;
																assign node37395 = (inp[5]) ? 4'b1001 : 4'b1101;
																assign node37398 = (inp[5]) ? 4'b1100 : 4'b1000;
														assign node37401 = (inp[0]) ? node37407 : node37402;
															assign node37402 = (inp[5]) ? 4'b1001 : node37403;
																assign node37403 = (inp[13]) ? 4'b1001 : 4'b1101;
															assign node37407 = (inp[13]) ? node37411 : node37408;
																assign node37408 = (inp[5]) ? 4'b1000 : 4'b1100;
																assign node37411 = (inp[5]) ? 4'b1101 : 4'b1001;
													assign node37414 = (inp[10]) ? node37422 : node37415;
														assign node37415 = (inp[5]) ? node37419 : node37416;
															assign node37416 = (inp[13]) ? 4'b1001 : 4'b1100;
															assign node37419 = (inp[13]) ? 4'b1100 : 4'b1001;
														assign node37422 = (inp[5]) ? node37426 : node37423;
															assign node37423 = (inp[13]) ? 4'b1000 : 4'b1100;
															assign node37426 = (inp[13]) ? node37428 : 4'b1000;
																assign node37428 = (inp[0]) ? 4'b1100 : 4'b1101;
											assign node37431 = (inp[5]) ? node37455 : node37432;
												assign node37432 = (inp[10]) ? node37444 : node37433;
													assign node37433 = (inp[0]) ? node37439 : node37434;
														assign node37434 = (inp[11]) ? 4'b1100 : node37435;
															assign node37435 = (inp[13]) ? 4'b1100 : 4'b1101;
														assign node37439 = (inp[13]) ? 4'b1101 : node37440;
															assign node37440 = (inp[11]) ? 4'b1101 : 4'b1100;
													assign node37444 = (inp[0]) ? node37450 : node37445;
														assign node37445 = (inp[11]) ? 4'b1101 : node37446;
															assign node37446 = (inp[13]) ? 4'b1101 : 4'b1100;
														assign node37450 = (inp[13]) ? 4'b1100 : node37451;
															assign node37451 = (inp[11]) ? 4'b1100 : 4'b1101;
												assign node37455 = (inp[13]) ? node37477 : node37456;
													assign node37456 = (inp[11]) ? node37464 : node37457;
														assign node37457 = (inp[10]) ? node37461 : node37458;
															assign node37458 = (inp[9]) ? 4'b1100 : 4'b1101;
															assign node37461 = (inp[0]) ? 4'b1101 : 4'b1100;
														assign node37464 = (inp[9]) ? node37472 : node37465;
															assign node37465 = (inp[10]) ? node37469 : node37466;
																assign node37466 = (inp[0]) ? 4'b1101 : 4'b1100;
																assign node37469 = (inp[0]) ? 4'b1100 : 4'b1101;
															assign node37472 = (inp[10]) ? node37474 : 4'b1101;
																assign node37474 = (inp[0]) ? 4'b1100 : 4'b1101;
													assign node37477 = (inp[11]) ? node37493 : node37478;
														assign node37478 = (inp[9]) ? node37486 : node37479;
															assign node37479 = (inp[0]) ? node37483 : node37480;
																assign node37480 = (inp[10]) ? 4'b1101 : 4'b1100;
																assign node37483 = (inp[10]) ? 4'b1100 : 4'b1101;
															assign node37486 = (inp[10]) ? node37490 : node37487;
																assign node37487 = (inp[0]) ? 4'b1101 : 4'b1100;
																assign node37490 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node37493 = (inp[9]) ? 4'b1100 : node37494;
															assign node37494 = (inp[0]) ? 4'b1101 : 4'b1100;
										assign node37498 = (inp[13]) ? node37564 : node37499;
											assign node37499 = (inp[8]) ? node37521 : node37500;
												assign node37500 = (inp[9]) ? node37510 : node37501;
													assign node37501 = (inp[10]) ? node37507 : node37502;
														assign node37502 = (inp[11]) ? 4'b1100 : node37503;
															assign node37503 = (inp[0]) ? 4'b1101 : 4'b1100;
														assign node37507 = (inp[5]) ? 4'b1101 : 4'b1100;
													assign node37510 = (inp[10]) ? node37516 : node37511;
														assign node37511 = (inp[11]) ? 4'b1101 : node37512;
															assign node37512 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node37516 = (inp[0]) ? node37518 : 4'b1100;
															assign node37518 = (inp[11]) ? 4'b1100 : 4'b1101;
												assign node37521 = (inp[5]) ? node37543 : node37522;
													assign node37522 = (inp[0]) ? node37530 : node37523;
														assign node37523 = (inp[10]) ? node37527 : node37524;
															assign node37524 = (inp[11]) ? 4'b1000 : 4'b1001;
															assign node37527 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node37530 = (inp[9]) ? node37536 : node37531;
															assign node37531 = (inp[11]) ? 4'b1000 : node37532;
																assign node37532 = (inp[10]) ? 4'b1001 : 4'b1000;
															assign node37536 = (inp[10]) ? node37540 : node37537;
																assign node37537 = (inp[11]) ? 4'b1001 : 4'b1000;
																assign node37540 = (inp[11]) ? 4'b1000 : 4'b1001;
													assign node37543 = (inp[0]) ? node37557 : node37544;
														assign node37544 = (inp[9]) ? node37550 : node37545;
															assign node37545 = (inp[11]) ? node37547 : 4'b1001;
																assign node37547 = (inp[10]) ? 4'b1001 : 4'b1000;
															assign node37550 = (inp[11]) ? node37554 : node37551;
																assign node37551 = (inp[10]) ? 4'b1000 : 4'b1001;
																assign node37554 = (inp[10]) ? 4'b1001 : 4'b1000;
														assign node37557 = (inp[10]) ? node37561 : node37558;
															assign node37558 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node37561 = (inp[11]) ? 4'b1000 : 4'b1001;
											assign node37564 = (inp[8]) ? node37596 : node37565;
												assign node37565 = (inp[0]) ? node37589 : node37566;
													assign node37566 = (inp[11]) ? node37574 : node37567;
														assign node37567 = (inp[9]) ? node37571 : node37568;
															assign node37568 = (inp[10]) ? 4'b1001 : 4'b1000;
															assign node37571 = (inp[10]) ? 4'b1000 : 4'b1001;
														assign node37574 = (inp[5]) ? node37582 : node37575;
															assign node37575 = (inp[10]) ? node37579 : node37576;
																assign node37576 = (inp[9]) ? 4'b1000 : 4'b1001;
																assign node37579 = (inp[9]) ? 4'b1001 : 4'b1000;
															assign node37582 = (inp[9]) ? node37586 : node37583;
																assign node37583 = (inp[10]) ? 4'b1000 : 4'b1001;
																assign node37586 = (inp[10]) ? 4'b1001 : 4'b1000;
													assign node37589 = (inp[9]) ? node37593 : node37590;
														assign node37590 = (inp[10]) ? 4'b1001 : 4'b1000;
														assign node37593 = (inp[10]) ? 4'b1000 : 4'b1001;
												assign node37596 = (inp[0]) ? node37600 : node37597;
													assign node37597 = (inp[10]) ? 4'b1001 : 4'b1000;
													assign node37600 = (inp[10]) ? 4'b1000 : 4'b1001;
				assign node37603 = (inp[12]) ? node41821 : node37604;
					assign node37604 = (inp[8]) ? node40414 : node37605;
						assign node37605 = (inp[7]) ? node39085 : node37606;
							assign node37606 = (inp[15]) ? node38284 : node37607;
								assign node37607 = (inp[4]) ? node37943 : node37608;
									assign node37608 = (inp[0]) ? node37778 : node37609;
										assign node37609 = (inp[1]) ? node37699 : node37610;
											assign node37610 = (inp[10]) ? node37654 : node37611;
												assign node37611 = (inp[13]) ? node37635 : node37612;
													assign node37612 = (inp[2]) ? node37624 : node37613;
														assign node37613 = (inp[5]) ? node37619 : node37614;
															assign node37614 = (inp[9]) ? 4'b0010 : node37615;
																assign node37615 = (inp[11]) ? 4'b0011 : 4'b0010;
															assign node37619 = (inp[11]) ? node37621 : 4'b0110;
																assign node37621 = (inp[9]) ? 4'b0110 : 4'b0111;
														assign node37624 = (inp[5]) ? node37628 : node37625;
															assign node37625 = (inp[9]) ? 4'b0111 : 4'b0110;
															assign node37628 = (inp[11]) ? node37632 : node37629;
																assign node37629 = (inp[9]) ? 4'b0010 : 4'b0011;
																assign node37632 = (inp[9]) ? 4'b0011 : 4'b0010;
													assign node37635 = (inp[9]) ? node37645 : node37636;
														assign node37636 = (inp[2]) ? node37642 : node37637;
															assign node37637 = (inp[5]) ? node37639 : 4'b0110;
																assign node37639 = (inp[11]) ? 4'b0010 : 4'b0011;
															assign node37642 = (inp[5]) ? 4'b0111 : 4'b0011;
														assign node37645 = (inp[2]) ? node37651 : node37646;
															assign node37646 = (inp[5]) ? node37648 : 4'b0111;
																assign node37648 = (inp[11]) ? 4'b0011 : 4'b0010;
															assign node37651 = (inp[5]) ? 4'b0110 : 4'b0010;
												assign node37654 = (inp[9]) ? node37678 : node37655;
													assign node37655 = (inp[5]) ? node37665 : node37656;
														assign node37656 = (inp[13]) ? node37662 : node37657;
															assign node37657 = (inp[2]) ? 4'b0111 : node37658;
																assign node37658 = (inp[11]) ? 4'b0010 : 4'b0011;
															assign node37662 = (inp[2]) ? 4'b0010 : 4'b0111;
														assign node37665 = (inp[2]) ? node37673 : node37666;
															assign node37666 = (inp[13]) ? node37670 : node37667;
																assign node37667 = (inp[11]) ? 4'b0110 : 4'b0111;
																assign node37670 = (inp[11]) ? 4'b0011 : 4'b0010;
															assign node37673 = (inp[13]) ? 4'b0110 : node37674;
																assign node37674 = (inp[11]) ? 4'b0011 : 4'b0010;
													assign node37678 = (inp[13]) ? node37692 : node37679;
														assign node37679 = (inp[5]) ? node37685 : node37680;
															assign node37680 = (inp[2]) ? 4'b0110 : node37681;
																assign node37681 = (inp[11]) ? 4'b0011 : 4'b0010;
															assign node37685 = (inp[2]) ? node37689 : node37686;
																assign node37686 = (inp[11]) ? 4'b0111 : 4'b0110;
																assign node37689 = (inp[11]) ? 4'b0010 : 4'b0011;
														assign node37692 = (inp[5]) ? node37696 : node37693;
															assign node37693 = (inp[2]) ? 4'b0011 : 4'b0110;
															assign node37696 = (inp[2]) ? 4'b0111 : 4'b0011;
											assign node37699 = (inp[2]) ? node37739 : node37700;
												assign node37700 = (inp[13]) ? node37724 : node37701;
													assign node37701 = (inp[9]) ? node37713 : node37702;
														assign node37702 = (inp[10]) ? node37708 : node37703;
															assign node37703 = (inp[11]) ? node37705 : 4'b0110;
																assign node37705 = (inp[5]) ? 4'b0110 : 4'b0111;
															assign node37708 = (inp[5]) ? 4'b0111 : node37709;
																assign node37709 = (inp[11]) ? 4'b0110 : 4'b0111;
														assign node37713 = (inp[10]) ? node37719 : node37714;
															assign node37714 = (inp[5]) ? 4'b0111 : node37715;
																assign node37715 = (inp[11]) ? 4'b0110 : 4'b0111;
															assign node37719 = (inp[5]) ? 4'b0110 : node37720;
																assign node37720 = (inp[11]) ? 4'b0111 : 4'b0110;
													assign node37724 = (inp[10]) ? node37734 : node37725;
														assign node37725 = (inp[9]) ? node37729 : node37726;
															assign node37726 = (inp[11]) ? 4'b0010 : 4'b0011;
															assign node37729 = (inp[11]) ? node37731 : 4'b0010;
																assign node37731 = (inp[5]) ? 4'b0010 : 4'b0011;
														assign node37734 = (inp[9]) ? node37736 : 4'b0010;
															assign node37736 = (inp[11]) ? 4'b0010 : 4'b0011;
												assign node37739 = (inp[13]) ? node37759 : node37740;
													assign node37740 = (inp[9]) ? node37748 : node37741;
														assign node37741 = (inp[10]) ? 4'b0010 : node37742;
															assign node37742 = (inp[5]) ? 4'b0011 : node37743;
																assign node37743 = (inp[11]) ? 4'b0010 : 4'b0011;
														assign node37748 = (inp[10]) ? node37754 : node37749;
															assign node37749 = (inp[5]) ? 4'b0010 : node37750;
																assign node37750 = (inp[11]) ? 4'b0011 : 4'b0010;
															assign node37754 = (inp[5]) ? 4'b0011 : node37755;
																assign node37755 = (inp[11]) ? 4'b0010 : 4'b0011;
													assign node37759 = (inp[10]) ? node37767 : node37760;
														assign node37760 = (inp[5]) ? node37762 : 4'b0110;
															assign node37762 = (inp[9]) ? node37764 : 4'b0110;
																assign node37764 = (inp[11]) ? 4'b0110 : 4'b0111;
														assign node37767 = (inp[9]) ? node37773 : node37768;
															assign node37768 = (inp[5]) ? node37770 : 4'b0110;
																assign node37770 = (inp[11]) ? 4'b0110 : 4'b0111;
															assign node37773 = (inp[5]) ? node37775 : 4'b0111;
																assign node37775 = (inp[11]) ? 4'b0111 : 4'b0110;
										assign node37778 = (inp[10]) ? node37870 : node37779;
											assign node37779 = (inp[9]) ? node37817 : node37780;
												assign node37780 = (inp[2]) ? node37792 : node37781;
													assign node37781 = (inp[13]) ? node37787 : node37782;
														assign node37782 = (inp[5]) ? 4'b0111 : node37783;
															assign node37783 = (inp[1]) ? 4'b0111 : 4'b0011;
														assign node37787 = (inp[5]) ? 4'b0010 : node37788;
															assign node37788 = (inp[1]) ? 4'b0010 : 4'b0111;
													assign node37792 = (inp[13]) ? node37804 : node37793;
														assign node37793 = (inp[1]) ? node37799 : node37794;
															assign node37794 = (inp[5]) ? 4'b0010 : node37795;
																assign node37795 = (inp[11]) ? 4'b0111 : 4'b0110;
															assign node37799 = (inp[11]) ? 4'b0010 : node37800;
																assign node37800 = (inp[5]) ? 4'b0011 : 4'b0010;
														assign node37804 = (inp[11]) ? node37810 : node37805;
															assign node37805 = (inp[1]) ? 4'b0111 : node37806;
																assign node37806 = (inp[5]) ? 4'b0111 : 4'b0011;
															assign node37810 = (inp[1]) ? node37814 : node37811;
																assign node37811 = (inp[5]) ? 4'b0110 : 4'b0010;
																assign node37814 = (inp[5]) ? 4'b0111 : 4'b0110;
												assign node37817 = (inp[11]) ? node37845 : node37818;
													assign node37818 = (inp[5]) ? node37834 : node37819;
														assign node37819 = (inp[1]) ? node37827 : node37820;
															assign node37820 = (inp[13]) ? node37824 : node37821;
																assign node37821 = (inp[2]) ? 4'b0111 : 4'b0010;
																assign node37824 = (inp[2]) ? 4'b0010 : 4'b0111;
															assign node37827 = (inp[2]) ? node37831 : node37828;
																assign node37828 = (inp[13]) ? 4'b0011 : 4'b0110;
																assign node37831 = (inp[13]) ? 4'b0110 : 4'b0011;
														assign node37834 = (inp[2]) ? node37842 : node37835;
															assign node37835 = (inp[13]) ? node37839 : node37836;
																assign node37836 = (inp[1]) ? 4'b0111 : 4'b0110;
																assign node37839 = (inp[1]) ? 4'b0010 : 4'b0011;
															assign node37842 = (inp[13]) ? 4'b0110 : 4'b0010;
													assign node37845 = (inp[2]) ? node37857 : node37846;
														assign node37846 = (inp[13]) ? node37852 : node37847;
															assign node37847 = (inp[1]) ? 4'b0110 : node37848;
																assign node37848 = (inp[5]) ? 4'b0110 : 4'b0010;
															assign node37852 = (inp[1]) ? 4'b0011 : node37853;
																assign node37853 = (inp[5]) ? 4'b0011 : 4'b0110;
														assign node37857 = (inp[13]) ? node37863 : node37858;
															assign node37858 = (inp[5]) ? 4'b0011 : node37859;
																assign node37859 = (inp[1]) ? 4'b0011 : 4'b0110;
															assign node37863 = (inp[5]) ? node37867 : node37864;
																assign node37864 = (inp[1]) ? 4'b0111 : 4'b0011;
																assign node37867 = (inp[1]) ? 4'b0110 : 4'b0111;
											assign node37870 = (inp[5]) ? node37904 : node37871;
												assign node37871 = (inp[1]) ? node37887 : node37872;
													assign node37872 = (inp[13]) ? node37878 : node37873;
														assign node37873 = (inp[2]) ? 4'b0110 : node37874;
															assign node37874 = (inp[9]) ? 4'b0011 : 4'b0010;
														assign node37878 = (inp[2]) ? 4'b0010 : node37879;
															assign node37879 = (inp[9]) ? node37883 : node37880;
																assign node37880 = (inp[11]) ? 4'b0110 : 4'b0111;
																assign node37883 = (inp[11]) ? 4'b0111 : 4'b0110;
													assign node37887 = (inp[9]) ? node37897 : node37888;
														assign node37888 = (inp[13]) ? node37892 : node37889;
															assign node37889 = (inp[2]) ? 4'b0011 : 4'b0110;
															assign node37892 = (inp[2]) ? node37894 : 4'b0011;
																assign node37894 = (inp[11]) ? 4'b0111 : 4'b0110;
														assign node37897 = (inp[2]) ? node37901 : node37898;
															assign node37898 = (inp[13]) ? 4'b0010 : 4'b0111;
															assign node37901 = (inp[13]) ? 4'b0110 : 4'b0010;
												assign node37904 = (inp[9]) ? node37928 : node37905;
													assign node37905 = (inp[11]) ? node37919 : node37906;
														assign node37906 = (inp[2]) ? node37914 : node37907;
															assign node37907 = (inp[13]) ? node37911 : node37908;
																assign node37908 = (inp[1]) ? 4'b0111 : 4'b0110;
																assign node37911 = (inp[1]) ? 4'b0010 : 4'b0011;
															assign node37914 = (inp[13]) ? 4'b0110 : node37915;
																assign node37915 = (inp[1]) ? 4'b0010 : 4'b0011;
														assign node37919 = (inp[2]) ? node37923 : node37920;
															assign node37920 = (inp[13]) ? 4'b0011 : 4'b0110;
															assign node37923 = (inp[13]) ? node37925 : 4'b0011;
																assign node37925 = (inp[1]) ? 4'b0110 : 4'b0111;
													assign node37928 = (inp[2]) ? node37936 : node37929;
														assign node37929 = (inp[13]) ? node37933 : node37930;
															assign node37930 = (inp[1]) ? 4'b0110 : 4'b0111;
															assign node37933 = (inp[1]) ? 4'b0011 : 4'b0010;
														assign node37936 = (inp[13]) ? node37938 : 4'b0010;
															assign node37938 = (inp[1]) ? 4'b0111 : node37939;
																assign node37939 = (inp[11]) ? 4'b0110 : 4'b0111;
									assign node37943 = (inp[13]) ? node38119 : node37944;
										assign node37944 = (inp[2]) ? node38032 : node37945;
											assign node37945 = (inp[5]) ? node37985 : node37946;
												assign node37946 = (inp[9]) ? node37966 : node37947;
													assign node37947 = (inp[10]) ? node37959 : node37948;
														assign node37948 = (inp[0]) ? node37954 : node37949;
															assign node37949 = (inp[1]) ? 4'b0000 : node37950;
																assign node37950 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node37954 = (inp[1]) ? node37956 : 4'b0001;
																assign node37956 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node37959 = (inp[0]) ? 4'b0000 : node37960;
															assign node37960 = (inp[11]) ? node37962 : 4'b0001;
																assign node37962 = (inp[1]) ? 4'b0001 : 4'b0000;
													assign node37966 = (inp[10]) ? node37978 : node37967;
														assign node37967 = (inp[0]) ? node37973 : node37968;
															assign node37968 = (inp[11]) ? node37970 : 4'b0001;
																assign node37970 = (inp[1]) ? 4'b0001 : 4'b0000;
															assign node37973 = (inp[11]) ? 4'b0000 : node37974;
																assign node37974 = (inp[1]) ? 4'b0001 : 4'b0000;
														assign node37978 = (inp[1]) ? node37980 : 4'b0001;
															assign node37980 = (inp[11]) ? node37982 : 4'b0000;
																assign node37982 = (inp[0]) ? 4'b0001 : 4'b0000;
												assign node37985 = (inp[1]) ? node38009 : node37986;
													assign node37986 = (inp[11]) ? node37996 : node37987;
														assign node37987 = (inp[0]) ? node37989 : 4'b0000;
															assign node37989 = (inp[10]) ? node37993 : node37990;
																assign node37990 = (inp[9]) ? 4'b0001 : 4'b0000;
																assign node37993 = (inp[9]) ? 4'b0000 : 4'b0001;
														assign node37996 = (inp[0]) ? node38002 : node37997;
															assign node37997 = (inp[10]) ? 4'b0001 : node37998;
																assign node37998 = (inp[9]) ? 4'b0001 : 4'b0000;
															assign node38002 = (inp[9]) ? node38006 : node38003;
																assign node38003 = (inp[10]) ? 4'b0001 : 4'b0000;
																assign node38006 = (inp[10]) ? 4'b0000 : 4'b0001;
													assign node38009 = (inp[9]) ? node38021 : node38010;
														assign node38010 = (inp[10]) ? node38016 : node38011;
															assign node38011 = (inp[11]) ? 4'b0100 : node38012;
																assign node38012 = (inp[0]) ? 4'b0100 : 4'b0101;
															assign node38016 = (inp[11]) ? 4'b0101 : node38017;
																assign node38017 = (inp[0]) ? 4'b0101 : 4'b0100;
														assign node38021 = (inp[10]) ? node38027 : node38022;
															assign node38022 = (inp[11]) ? 4'b0101 : node38023;
																assign node38023 = (inp[0]) ? 4'b0101 : 4'b0100;
															assign node38027 = (inp[11]) ? 4'b0100 : node38028;
																assign node38028 = (inp[0]) ? 4'b0100 : 4'b0101;
											assign node38032 = (inp[1]) ? node38076 : node38033;
												assign node38033 = (inp[5]) ? node38053 : node38034;
													assign node38034 = (inp[11]) ? node38042 : node38035;
														assign node38035 = (inp[10]) ? node38039 : node38036;
															assign node38036 = (inp[9]) ? 4'b0100 : 4'b0101;
															assign node38039 = (inp[9]) ? 4'b0101 : 4'b0100;
														assign node38042 = (inp[9]) ? node38048 : node38043;
															assign node38043 = (inp[10]) ? node38045 : 4'b0100;
																assign node38045 = (inp[0]) ? 4'b0101 : 4'b0100;
															assign node38048 = (inp[10]) ? node38050 : 4'b0101;
																assign node38050 = (inp[0]) ? 4'b0100 : 4'b0101;
													assign node38053 = (inp[11]) ? node38061 : node38054;
														assign node38054 = (inp[10]) ? node38058 : node38055;
															assign node38055 = (inp[9]) ? 4'b0101 : 4'b0100;
															assign node38058 = (inp[9]) ? 4'b0100 : 4'b0101;
														assign node38061 = (inp[0]) ? node38069 : node38062;
															assign node38062 = (inp[10]) ? node38066 : node38063;
																assign node38063 = (inp[9]) ? 4'b0101 : 4'b0100;
																assign node38066 = (inp[9]) ? 4'b0100 : 4'b0101;
															assign node38069 = (inp[10]) ? node38073 : node38070;
																assign node38070 = (inp[9]) ? 4'b0100 : 4'b0101;
																assign node38073 = (inp[9]) ? 4'b0101 : 4'b0100;
												assign node38076 = (inp[5]) ? node38098 : node38077;
													assign node38077 = (inp[0]) ? node38091 : node38078;
														assign node38078 = (inp[11]) ? node38084 : node38079;
															assign node38079 = (inp[10]) ? node38081 : 4'b0101;
																assign node38081 = (inp[9]) ? 4'b0100 : 4'b0101;
															assign node38084 = (inp[9]) ? node38088 : node38085;
																assign node38085 = (inp[10]) ? 4'b0100 : 4'b0101;
																assign node38088 = (inp[10]) ? 4'b0101 : 4'b0100;
														assign node38091 = (inp[9]) ? node38095 : node38092;
															assign node38092 = (inp[10]) ? 4'b0100 : 4'b0101;
															assign node38095 = (inp[10]) ? 4'b0101 : 4'b0100;
													assign node38098 = (inp[9]) ? node38108 : node38099;
														assign node38099 = (inp[11]) ? 4'b0001 : node38100;
															assign node38100 = (inp[0]) ? node38104 : node38101;
																assign node38101 = (inp[10]) ? 4'b0000 : 4'b0001;
																assign node38104 = (inp[10]) ? 4'b0001 : 4'b0000;
														assign node38108 = (inp[10]) ? node38114 : node38109;
															assign node38109 = (inp[11]) ? 4'b0001 : node38110;
																assign node38110 = (inp[0]) ? 4'b0001 : 4'b0000;
															assign node38114 = (inp[0]) ? 4'b0000 : node38115;
																assign node38115 = (inp[11]) ? 4'b0000 : 4'b0001;
										assign node38119 = (inp[2]) ? node38199 : node38120;
											assign node38120 = (inp[1]) ? node38166 : node38121;
												assign node38121 = (inp[10]) ? node38145 : node38122;
													assign node38122 = (inp[11]) ? node38130 : node38123;
														assign node38123 = (inp[9]) ? node38127 : node38124;
															assign node38124 = (inp[5]) ? 4'b0101 : 4'b0100;
															assign node38127 = (inp[5]) ? 4'b0100 : 4'b0101;
														assign node38130 = (inp[0]) ? node38138 : node38131;
															assign node38131 = (inp[5]) ? node38135 : node38132;
																assign node38132 = (inp[9]) ? 4'b0101 : 4'b0100;
																assign node38135 = (inp[9]) ? 4'b0100 : 4'b0101;
															assign node38138 = (inp[5]) ? node38142 : node38139;
																assign node38139 = (inp[9]) ? 4'b0100 : 4'b0101;
																assign node38142 = (inp[9]) ? 4'b0101 : 4'b0100;
													assign node38145 = (inp[9]) ? node38157 : node38146;
														assign node38146 = (inp[5]) ? node38152 : node38147;
															assign node38147 = (inp[0]) ? node38149 : 4'b0101;
																assign node38149 = (inp[11]) ? 4'b0100 : 4'b0101;
															assign node38152 = (inp[0]) ? node38154 : 4'b0100;
																assign node38154 = (inp[11]) ? 4'b0101 : 4'b0100;
														assign node38157 = (inp[5]) ? node38161 : node38158;
															assign node38158 = (inp[0]) ? 4'b0101 : 4'b0100;
															assign node38161 = (inp[0]) ? node38163 : 4'b0101;
																assign node38163 = (inp[11]) ? 4'b0100 : 4'b0101;
												assign node38166 = (inp[5]) ? node38182 : node38167;
													assign node38167 = (inp[10]) ? node38173 : node38168;
														assign node38168 = (inp[9]) ? node38170 : 4'b0100;
															assign node38170 = (inp[0]) ? 4'b0101 : 4'b0100;
														assign node38173 = (inp[9]) ? node38179 : node38174;
															assign node38174 = (inp[11]) ? 4'b0101 : node38175;
																assign node38175 = (inp[0]) ? 4'b0101 : 4'b0100;
															assign node38179 = (inp[0]) ? 4'b0100 : 4'b0101;
													assign node38182 = (inp[9]) ? node38188 : node38183;
														assign node38183 = (inp[10]) ? 4'b0000 : node38184;
															assign node38184 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node38188 = (inp[10]) ? node38194 : node38189;
															assign node38189 = (inp[11]) ? 4'b0000 : node38190;
																assign node38190 = (inp[0]) ? 4'b0000 : 4'b0001;
															assign node38194 = (inp[11]) ? 4'b0001 : node38195;
																assign node38195 = (inp[0]) ? 4'b0001 : 4'b0000;
											assign node38199 = (inp[1]) ? node38251 : node38200;
												assign node38200 = (inp[11]) ? node38230 : node38201;
													assign node38201 = (inp[5]) ? node38217 : node38202;
														assign node38202 = (inp[0]) ? node38210 : node38203;
															assign node38203 = (inp[10]) ? node38207 : node38204;
																assign node38204 = (inp[9]) ? 4'b0001 : 4'b0000;
																assign node38207 = (inp[9]) ? 4'b0000 : 4'b0001;
															assign node38210 = (inp[10]) ? node38214 : node38211;
																assign node38211 = (inp[9]) ? 4'b0001 : 4'b0000;
																assign node38214 = (inp[9]) ? 4'b0000 : 4'b0001;
														assign node38217 = (inp[0]) ? node38225 : node38218;
															assign node38218 = (inp[9]) ? node38222 : node38219;
																assign node38219 = (inp[10]) ? 4'b0000 : 4'b0001;
																assign node38222 = (inp[10]) ? 4'b0001 : 4'b0000;
															assign node38225 = (inp[9]) ? 4'b0000 : node38226;
																assign node38226 = (inp[10]) ? 4'b0000 : 4'b0001;
													assign node38230 = (inp[10]) ? node38240 : node38231;
														assign node38231 = (inp[5]) ? node38233 : 4'b0000;
															assign node38233 = (inp[0]) ? node38237 : node38234;
																assign node38234 = (inp[9]) ? 4'b0000 : 4'b0001;
																assign node38237 = (inp[9]) ? 4'b0001 : 4'b0000;
														assign node38240 = (inp[0]) ? node38246 : node38241;
															assign node38241 = (inp[9]) ? 4'b0000 : node38242;
																assign node38242 = (inp[5]) ? 4'b0000 : 4'b0001;
															assign node38246 = (inp[5]) ? 4'b0001 : node38247;
																assign node38247 = (inp[9]) ? 4'b0001 : 4'b0000;
												assign node38251 = (inp[5]) ? node38263 : node38252;
													assign node38252 = (inp[10]) ? node38258 : node38253;
														assign node38253 = (inp[11]) ? node38255 : 4'b0001;
															assign node38255 = (inp[9]) ? 4'b0001 : 4'b0000;
														assign node38258 = (inp[9]) ? 4'b0000 : node38259;
															assign node38259 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node38263 = (inp[11]) ? node38271 : node38264;
														assign node38264 = (inp[10]) ? node38268 : node38265;
															assign node38265 = (inp[9]) ? 4'b0100 : 4'b0101;
															assign node38268 = (inp[9]) ? 4'b0101 : 4'b0100;
														assign node38271 = (inp[10]) ? node38277 : node38272;
															assign node38272 = (inp[9]) ? 4'b0100 : node38273;
																assign node38273 = (inp[0]) ? 4'b0100 : 4'b0101;
															assign node38277 = (inp[0]) ? node38281 : node38278;
																assign node38278 = (inp[9]) ? 4'b0101 : 4'b0100;
																assign node38281 = (inp[9]) ? 4'b0100 : 4'b0101;
								assign node38284 = (inp[11]) ? node38686 : node38285;
									assign node38285 = (inp[2]) ? node38487 : node38286;
										assign node38286 = (inp[4]) ? node38384 : node38287;
											assign node38287 = (inp[13]) ? node38337 : node38288;
												assign node38288 = (inp[5]) ? node38314 : node38289;
													assign node38289 = (inp[1]) ? node38299 : node38290;
														assign node38290 = (inp[9]) ? 4'b0000 : node38291;
															assign node38291 = (inp[10]) ? node38295 : node38292;
																assign node38292 = (inp[0]) ? 4'b0001 : 4'b0000;
																assign node38295 = (inp[0]) ? 4'b0000 : 4'b0001;
														assign node38299 = (inp[9]) ? node38307 : node38300;
															assign node38300 = (inp[10]) ? node38304 : node38301;
																assign node38301 = (inp[0]) ? 4'b0000 : 4'b0001;
																assign node38304 = (inp[0]) ? 4'b0001 : 4'b0000;
															assign node38307 = (inp[10]) ? node38311 : node38308;
																assign node38308 = (inp[0]) ? 4'b0001 : 4'b0000;
																assign node38311 = (inp[0]) ? 4'b0000 : 4'b0001;
													assign node38314 = (inp[1]) ? node38322 : node38315;
														assign node38315 = (inp[9]) ? node38319 : node38316;
															assign node38316 = (inp[10]) ? 4'b0001 : 4'b0000;
															assign node38319 = (inp[10]) ? 4'b0000 : 4'b0001;
														assign node38322 = (inp[0]) ? node38330 : node38323;
															assign node38323 = (inp[10]) ? node38327 : node38324;
																assign node38324 = (inp[9]) ? 4'b0100 : 4'b0101;
																assign node38327 = (inp[9]) ? 4'b0101 : 4'b0100;
															assign node38330 = (inp[10]) ? node38334 : node38331;
																assign node38331 = (inp[9]) ? 4'b0101 : 4'b0100;
																assign node38334 = (inp[9]) ? 4'b0100 : 4'b0101;
												assign node38337 = (inp[5]) ? node38359 : node38338;
													assign node38338 = (inp[10]) ? node38352 : node38339;
														assign node38339 = (inp[0]) ? node38347 : node38340;
															assign node38340 = (inp[1]) ? node38344 : node38341;
																assign node38341 = (inp[9]) ? 4'b0100 : 4'b0101;
																assign node38344 = (inp[9]) ? 4'b0101 : 4'b0100;
															assign node38347 = (inp[1]) ? node38349 : 4'b0100;
																assign node38349 = (inp[9]) ? 4'b0101 : 4'b0100;
														assign node38352 = (inp[9]) ? node38356 : node38353;
															assign node38353 = (inp[1]) ? 4'b0101 : 4'b0100;
															assign node38356 = (inp[1]) ? 4'b0100 : 4'b0101;
													assign node38359 = (inp[1]) ? node38369 : node38360;
														assign node38360 = (inp[10]) ? 4'b0100 : node38361;
															assign node38361 = (inp[0]) ? node38365 : node38362;
																assign node38362 = (inp[9]) ? 4'b0101 : 4'b0100;
																assign node38365 = (inp[9]) ? 4'b0100 : 4'b0101;
														assign node38369 = (inp[9]) ? node38377 : node38370;
															assign node38370 = (inp[0]) ? node38374 : node38371;
																assign node38371 = (inp[10]) ? 4'b0000 : 4'b0001;
																assign node38374 = (inp[10]) ? 4'b0001 : 4'b0000;
															assign node38377 = (inp[10]) ? node38381 : node38378;
																assign node38378 = (inp[0]) ? 4'b0001 : 4'b0000;
																assign node38381 = (inp[0]) ? 4'b0000 : 4'b0001;
											assign node38384 = (inp[13]) ? node38436 : node38385;
												assign node38385 = (inp[5]) ? node38415 : node38386;
													assign node38386 = (inp[0]) ? node38402 : node38387;
														assign node38387 = (inp[9]) ? node38395 : node38388;
															assign node38388 = (inp[10]) ? node38392 : node38389;
																assign node38389 = (inp[1]) ? 4'b0101 : 4'b0100;
																assign node38392 = (inp[1]) ? 4'b0100 : 4'b0101;
															assign node38395 = (inp[1]) ? node38399 : node38396;
																assign node38396 = (inp[10]) ? 4'b0100 : 4'b0101;
																assign node38399 = (inp[10]) ? 4'b0101 : 4'b0100;
														assign node38402 = (inp[1]) ? node38410 : node38403;
															assign node38403 = (inp[10]) ? node38407 : node38404;
																assign node38404 = (inp[9]) ? 4'b0100 : 4'b0101;
																assign node38407 = (inp[9]) ? 4'b0101 : 4'b0100;
															assign node38410 = (inp[10]) ? 4'b0101 : node38411;
																assign node38411 = (inp[9]) ? 4'b0101 : 4'b0100;
													assign node38415 = (inp[1]) ? node38423 : node38416;
														assign node38416 = (inp[9]) ? node38418 : 4'b0101;
															assign node38418 = (inp[0]) ? 4'b0100 : node38419;
																assign node38419 = (inp[10]) ? 4'b0101 : 4'b0100;
														assign node38423 = (inp[10]) ? node38429 : node38424;
															assign node38424 = (inp[0]) ? 4'b0001 : node38425;
																assign node38425 = (inp[9]) ? 4'b0001 : 4'b0000;
															assign node38429 = (inp[0]) ? node38433 : node38430;
																assign node38430 = (inp[9]) ? 4'b0000 : 4'b0001;
																assign node38433 = (inp[9]) ? 4'b0001 : 4'b0000;
												assign node38436 = (inp[5]) ? node38464 : node38437;
													assign node38437 = (inp[0]) ? node38451 : node38438;
														assign node38438 = (inp[10]) ? node38444 : node38439;
															assign node38439 = (inp[9]) ? node38441 : 4'b0001;
																assign node38441 = (inp[1]) ? 4'b0000 : 4'b0001;
															assign node38444 = (inp[1]) ? node38448 : node38445;
																assign node38445 = (inp[9]) ? 4'b0000 : 4'b0001;
																assign node38448 = (inp[9]) ? 4'b0001 : 4'b0000;
														assign node38451 = (inp[9]) ? node38459 : node38452;
															assign node38452 = (inp[1]) ? node38456 : node38453;
																assign node38453 = (inp[10]) ? 4'b0000 : 4'b0001;
																assign node38456 = (inp[10]) ? 4'b0001 : 4'b0000;
															assign node38459 = (inp[10]) ? 4'b0000 : node38460;
																assign node38460 = (inp[1]) ? 4'b0001 : 4'b0000;
													assign node38464 = (inp[1]) ? node38480 : node38465;
														assign node38465 = (inp[10]) ? node38473 : node38466;
															assign node38466 = (inp[9]) ? node38470 : node38467;
																assign node38467 = (inp[0]) ? 4'b0000 : 4'b0001;
																assign node38470 = (inp[0]) ? 4'b0001 : 4'b0000;
															assign node38473 = (inp[9]) ? node38477 : node38474;
																assign node38474 = (inp[0]) ? 4'b0001 : 4'b0000;
																assign node38477 = (inp[0]) ? 4'b0000 : 4'b0001;
														assign node38480 = (inp[9]) ? node38484 : node38481;
															assign node38481 = (inp[10]) ? 4'b0100 : 4'b0101;
															assign node38484 = (inp[10]) ? 4'b0101 : 4'b0100;
										assign node38487 = (inp[1]) ? node38585 : node38488;
											assign node38488 = (inp[5]) ? node38526 : node38489;
												assign node38489 = (inp[9]) ? node38507 : node38490;
													assign node38490 = (inp[4]) ? node38498 : node38491;
														assign node38491 = (inp[13]) ? node38495 : node38492;
															assign node38492 = (inp[10]) ? 4'b0101 : 4'b0100;
															assign node38495 = (inp[10]) ? 4'b0001 : 4'b0000;
														assign node38498 = (inp[13]) ? node38504 : node38499;
															assign node38499 = (inp[10]) ? 4'b0000 : node38500;
																assign node38500 = (inp[0]) ? 4'b0001 : 4'b0000;
															assign node38504 = (inp[10]) ? 4'b0100 : 4'b0101;
													assign node38507 = (inp[10]) ? node38517 : node38508;
														assign node38508 = (inp[4]) ? node38512 : node38509;
															assign node38509 = (inp[13]) ? 4'b0001 : 4'b0101;
															assign node38512 = (inp[13]) ? 4'b0100 : node38513;
																assign node38513 = (inp[0]) ? 4'b0000 : 4'b0001;
														assign node38517 = (inp[4]) ? node38521 : node38518;
															assign node38518 = (inp[13]) ? 4'b0000 : 4'b0100;
															assign node38521 = (inp[13]) ? 4'b0101 : node38522;
																assign node38522 = (inp[0]) ? 4'b0001 : 4'b0000;
												assign node38526 = (inp[9]) ? node38554 : node38527;
													assign node38527 = (inp[10]) ? node38541 : node38528;
														assign node38528 = (inp[0]) ? node38534 : node38529;
															assign node38529 = (inp[13]) ? node38531 : 4'b0001;
																assign node38531 = (inp[4]) ? 4'b0100 : 4'b0001;
															assign node38534 = (inp[13]) ? node38538 : node38535;
																assign node38535 = (inp[4]) ? 4'b0000 : 4'b0100;
																assign node38538 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node38541 = (inp[0]) ? node38549 : node38542;
															assign node38542 = (inp[13]) ? node38546 : node38543;
																assign node38543 = (inp[4]) ? 4'b0000 : 4'b0100;
																assign node38546 = (inp[4]) ? 4'b0101 : 4'b0000;
															assign node38549 = (inp[4]) ? 4'b0001 : node38550;
																assign node38550 = (inp[13]) ? 4'b0001 : 4'b0101;
													assign node38554 = (inp[10]) ? node38570 : node38555;
														assign node38555 = (inp[0]) ? node38563 : node38556;
															assign node38556 = (inp[4]) ? node38560 : node38557;
																assign node38557 = (inp[13]) ? 4'b0000 : 4'b0100;
																assign node38560 = (inp[13]) ? 4'b0101 : 4'b0000;
															assign node38563 = (inp[13]) ? node38567 : node38564;
																assign node38564 = (inp[4]) ? 4'b0001 : 4'b0101;
																assign node38567 = (inp[4]) ? 4'b0101 : 4'b0001;
														assign node38570 = (inp[0]) ? node38578 : node38571;
															assign node38571 = (inp[13]) ? node38575 : node38572;
																assign node38572 = (inp[4]) ? 4'b0001 : 4'b0101;
																assign node38575 = (inp[4]) ? 4'b0100 : 4'b0001;
															assign node38578 = (inp[4]) ? node38582 : node38579;
																assign node38579 = (inp[13]) ? 4'b0000 : 4'b0100;
																assign node38582 = (inp[13]) ? 4'b0100 : 4'b0000;
											assign node38585 = (inp[5]) ? node38645 : node38586;
												assign node38586 = (inp[0]) ? node38618 : node38587;
													assign node38587 = (inp[10]) ? node38603 : node38588;
														assign node38588 = (inp[9]) ? node38596 : node38589;
															assign node38589 = (inp[13]) ? node38593 : node38590;
																assign node38590 = (inp[4]) ? 4'b0001 : 4'b0101;
																assign node38593 = (inp[4]) ? 4'b0100 : 4'b0001;
															assign node38596 = (inp[13]) ? node38600 : node38597;
																assign node38597 = (inp[4]) ? 4'b0000 : 4'b0100;
																assign node38600 = (inp[4]) ? 4'b0101 : 4'b0000;
														assign node38603 = (inp[9]) ? node38611 : node38604;
															assign node38604 = (inp[4]) ? node38608 : node38605;
																assign node38605 = (inp[13]) ? 4'b0000 : 4'b0100;
																assign node38608 = (inp[13]) ? 4'b0101 : 4'b0000;
															assign node38611 = (inp[4]) ? node38615 : node38612;
																assign node38612 = (inp[13]) ? 4'b0001 : 4'b0101;
																assign node38615 = (inp[13]) ? 4'b0100 : 4'b0001;
													assign node38618 = (inp[9]) ? node38630 : node38619;
														assign node38619 = (inp[10]) ? node38625 : node38620;
															assign node38620 = (inp[4]) ? node38622 : 4'b0101;
																assign node38622 = (inp[13]) ? 4'b0100 : 4'b0000;
															assign node38625 = (inp[4]) ? 4'b0101 : node38626;
																assign node38626 = (inp[13]) ? 4'b0000 : 4'b0100;
														assign node38630 = (inp[10]) ? node38638 : node38631;
															assign node38631 = (inp[4]) ? node38635 : node38632;
																assign node38632 = (inp[13]) ? 4'b0000 : 4'b0100;
																assign node38635 = (inp[13]) ? 4'b0101 : 4'b0001;
															assign node38638 = (inp[4]) ? node38642 : node38639;
																assign node38639 = (inp[13]) ? 4'b0001 : 4'b0101;
																assign node38642 = (inp[13]) ? 4'b0100 : 4'b0000;
												assign node38645 = (inp[0]) ? node38663 : node38646;
													assign node38646 = (inp[4]) ? node38654 : node38647;
														assign node38647 = (inp[13]) ? node38649 : 4'b0000;
															assign node38649 = (inp[9]) ? node38651 : 4'b0100;
																assign node38651 = (inp[10]) ? 4'b0101 : 4'b0100;
														assign node38654 = (inp[13]) ? 4'b0000 : node38655;
															assign node38655 = (inp[9]) ? node38659 : node38656;
																assign node38656 = (inp[10]) ? 4'b0100 : 4'b0101;
																assign node38659 = (inp[10]) ? 4'b0101 : 4'b0100;
													assign node38663 = (inp[10]) ? node38673 : node38664;
														assign node38664 = (inp[9]) ? node38666 : 4'b0001;
															assign node38666 = (inp[4]) ? node38670 : node38667;
																assign node38667 = (inp[13]) ? 4'b0100 : 4'b0000;
																assign node38670 = (inp[13]) ? 4'b0000 : 4'b0100;
														assign node38673 = (inp[9]) ? node38681 : node38674;
															assign node38674 = (inp[4]) ? node38678 : node38675;
																assign node38675 = (inp[13]) ? 4'b0100 : 4'b0000;
																assign node38678 = (inp[13]) ? 4'b0000 : 4'b0100;
															assign node38681 = (inp[4]) ? 4'b0101 : node38682;
																assign node38682 = (inp[13]) ? 4'b0101 : 4'b0001;
									assign node38686 = (inp[2]) ? node38872 : node38687;
										assign node38687 = (inp[5]) ? node38791 : node38688;
											assign node38688 = (inp[4]) ? node38746 : node38689;
												assign node38689 = (inp[13]) ? node38717 : node38690;
													assign node38690 = (inp[1]) ? node38704 : node38691;
														assign node38691 = (inp[0]) ? node38699 : node38692;
															assign node38692 = (inp[9]) ? node38696 : node38693;
																assign node38693 = (inp[10]) ? 4'b0000 : 4'b0001;
																assign node38696 = (inp[10]) ? 4'b0001 : 4'b0000;
															assign node38699 = (inp[9]) ? 4'b0001 : node38700;
																assign node38700 = (inp[10]) ? 4'b0000 : 4'b0001;
														assign node38704 = (inp[0]) ? node38712 : node38705;
															assign node38705 = (inp[10]) ? node38709 : node38706;
																assign node38706 = (inp[9]) ? 4'b0001 : 4'b0000;
																assign node38709 = (inp[9]) ? 4'b0000 : 4'b0001;
															assign node38712 = (inp[10]) ? 4'b0000 : node38713;
																assign node38713 = (inp[9]) ? 4'b0001 : 4'b0000;
													assign node38717 = (inp[1]) ? node38731 : node38718;
														assign node38718 = (inp[0]) ? node38726 : node38719;
															assign node38719 = (inp[9]) ? node38723 : node38720;
																assign node38720 = (inp[10]) ? 4'b0100 : 4'b0101;
																assign node38723 = (inp[10]) ? 4'b0101 : 4'b0100;
															assign node38726 = (inp[9]) ? 4'b0100 : node38727;
																assign node38727 = (inp[10]) ? 4'b0101 : 4'b0100;
														assign node38731 = (inp[10]) ? node38739 : node38732;
															assign node38732 = (inp[9]) ? node38736 : node38733;
																assign node38733 = (inp[0]) ? 4'b0101 : 4'b0100;
																assign node38736 = (inp[0]) ? 4'b0100 : 4'b0101;
															assign node38739 = (inp[9]) ? node38743 : node38740;
																assign node38740 = (inp[0]) ? 4'b0100 : 4'b0101;
																assign node38743 = (inp[0]) ? 4'b0101 : 4'b0100;
												assign node38746 = (inp[13]) ? node38762 : node38747;
													assign node38747 = (inp[9]) ? node38755 : node38748;
														assign node38748 = (inp[10]) ? node38752 : node38749;
															assign node38749 = (inp[1]) ? 4'b0100 : 4'b0101;
															assign node38752 = (inp[1]) ? 4'b0101 : 4'b0100;
														assign node38755 = (inp[1]) ? node38759 : node38756;
															assign node38756 = (inp[10]) ? 4'b0101 : 4'b0100;
															assign node38759 = (inp[10]) ? 4'b0100 : 4'b0101;
													assign node38762 = (inp[0]) ? node38776 : node38763;
														assign node38763 = (inp[9]) ? node38769 : node38764;
															assign node38764 = (inp[10]) ? node38766 : 4'b0001;
																assign node38766 = (inp[1]) ? 4'b0001 : 4'b0000;
															assign node38769 = (inp[10]) ? node38773 : node38770;
																assign node38770 = (inp[1]) ? 4'b0001 : 4'b0000;
																assign node38773 = (inp[1]) ? 4'b0000 : 4'b0001;
														assign node38776 = (inp[9]) ? node38784 : node38777;
															assign node38777 = (inp[1]) ? node38781 : node38778;
																assign node38778 = (inp[10]) ? 4'b0000 : 4'b0001;
																assign node38781 = (inp[10]) ? 4'b0001 : 4'b0000;
															assign node38784 = (inp[1]) ? node38788 : node38785;
																assign node38785 = (inp[10]) ? 4'b0001 : 4'b0000;
																assign node38788 = (inp[10]) ? 4'b0000 : 4'b0001;
											assign node38791 = (inp[10]) ? node38835 : node38792;
												assign node38792 = (inp[9]) ? node38816 : node38793;
													assign node38793 = (inp[13]) ? node38801 : node38794;
														assign node38794 = (inp[1]) ? node38798 : node38795;
															assign node38795 = (inp[4]) ? 4'b0100 : 4'b0000;
															assign node38798 = (inp[4]) ? 4'b0001 : 4'b0100;
														assign node38801 = (inp[0]) ? node38809 : node38802;
															assign node38802 = (inp[1]) ? node38806 : node38803;
																assign node38803 = (inp[4]) ? 4'b0000 : 4'b0101;
																assign node38806 = (inp[4]) ? 4'b0101 : 4'b0000;
															assign node38809 = (inp[1]) ? node38813 : node38810;
																assign node38810 = (inp[4]) ? 4'b0000 : 4'b0101;
																assign node38813 = (inp[4]) ? 4'b0100 : 4'b0000;
													assign node38816 = (inp[1]) ? node38826 : node38817;
														assign node38817 = (inp[4]) ? node38823 : node38818;
															assign node38818 = (inp[13]) ? 4'b0100 : node38819;
																assign node38819 = (inp[0]) ? 4'b0000 : 4'b0001;
															assign node38823 = (inp[13]) ? 4'b0001 : 4'b0101;
														assign node38826 = (inp[4]) ? node38830 : node38827;
															assign node38827 = (inp[13]) ? 4'b0001 : 4'b0101;
															assign node38830 = (inp[13]) ? node38832 : 4'b0000;
																assign node38832 = (inp[0]) ? 4'b0101 : 4'b0100;
												assign node38835 = (inp[9]) ? node38853 : node38836;
													assign node38836 = (inp[4]) ? node38844 : node38837;
														assign node38837 = (inp[13]) ? node38841 : node38838;
															assign node38838 = (inp[1]) ? 4'b0101 : 4'b0001;
															assign node38841 = (inp[1]) ? 4'b0001 : 4'b0100;
														assign node38844 = (inp[1]) ? node38848 : node38845;
															assign node38845 = (inp[13]) ? 4'b0001 : 4'b0101;
															assign node38848 = (inp[13]) ? node38850 : 4'b0000;
																assign node38850 = (inp[0]) ? 4'b0101 : 4'b0100;
													assign node38853 = (inp[13]) ? node38863 : node38854;
														assign node38854 = (inp[1]) ? node38860 : node38855;
															assign node38855 = (inp[4]) ? 4'b0100 : node38856;
																assign node38856 = (inp[0]) ? 4'b0001 : 4'b0000;
															assign node38860 = (inp[4]) ? 4'b0001 : 4'b0100;
														assign node38863 = (inp[1]) ? node38867 : node38864;
															assign node38864 = (inp[4]) ? 4'b0000 : 4'b0101;
															assign node38867 = (inp[4]) ? node38869 : 4'b0000;
																assign node38869 = (inp[0]) ? 4'b0100 : 4'b0101;
										assign node38872 = (inp[0]) ? node38972 : node38873;
											assign node38873 = (inp[13]) ? node38927 : node38874;
												assign node38874 = (inp[4]) ? node38900 : node38875;
													assign node38875 = (inp[5]) ? node38889 : node38876;
														assign node38876 = (inp[9]) ? node38884 : node38877;
															assign node38877 = (inp[1]) ? node38881 : node38878;
																assign node38878 = (inp[10]) ? 4'b0101 : 4'b0100;
																assign node38881 = (inp[10]) ? 4'b0100 : 4'b0101;
															assign node38884 = (inp[10]) ? node38886 : 4'b0101;
																assign node38886 = (inp[1]) ? 4'b0101 : 4'b0100;
														assign node38889 = (inp[1]) ? node38893 : node38890;
															assign node38890 = (inp[10]) ? 4'b0100 : 4'b0101;
															assign node38893 = (inp[10]) ? node38897 : node38894;
																assign node38894 = (inp[9]) ? 4'b0000 : 4'b0001;
																assign node38897 = (inp[9]) ? 4'b0001 : 4'b0000;
													assign node38900 = (inp[5]) ? node38916 : node38901;
														assign node38901 = (inp[9]) ? node38909 : node38902;
															assign node38902 = (inp[10]) ? node38906 : node38903;
																assign node38903 = (inp[1]) ? 4'b0000 : 4'b0001;
																assign node38906 = (inp[1]) ? 4'b0001 : 4'b0000;
															assign node38909 = (inp[1]) ? node38913 : node38910;
																assign node38910 = (inp[10]) ? 4'b0001 : 4'b0000;
																assign node38913 = (inp[10]) ? 4'b0000 : 4'b0001;
														assign node38916 = (inp[1]) ? node38922 : node38917;
															assign node38917 = (inp[10]) ? 4'b0001 : node38918;
																assign node38918 = (inp[9]) ? 4'b0001 : 4'b0000;
															assign node38922 = (inp[10]) ? 4'b0101 : node38923;
																assign node38923 = (inp[9]) ? 4'b0100 : 4'b0101;
												assign node38927 = (inp[4]) ? node38947 : node38928;
													assign node38928 = (inp[1]) ? node38936 : node38929;
														assign node38929 = (inp[9]) ? node38933 : node38930;
															assign node38930 = (inp[10]) ? 4'b0001 : 4'b0000;
															assign node38933 = (inp[10]) ? 4'b0000 : 4'b0001;
														assign node38936 = (inp[5]) ? node38942 : node38937;
															assign node38937 = (inp[10]) ? node38939 : 4'b0000;
																assign node38939 = (inp[9]) ? 4'b0001 : 4'b0000;
															assign node38942 = (inp[9]) ? node38944 : 4'b0101;
																assign node38944 = (inp[10]) ? 4'b0101 : 4'b0100;
													assign node38947 = (inp[1]) ? node38961 : node38948;
														assign node38948 = (inp[9]) ? node38956 : node38949;
															assign node38949 = (inp[10]) ? node38953 : node38950;
																assign node38950 = (inp[5]) ? 4'b0100 : 4'b0101;
																assign node38953 = (inp[5]) ? 4'b0101 : 4'b0100;
															assign node38956 = (inp[5]) ? node38958 : 4'b0101;
																assign node38958 = (inp[10]) ? 4'b0100 : 4'b0101;
														assign node38961 = (inp[5]) ? node38967 : node38962;
															assign node38962 = (inp[9]) ? 4'b0100 : node38963;
																assign node38963 = (inp[10]) ? 4'b0101 : 4'b0100;
															assign node38967 = (inp[10]) ? node38969 : 4'b0000;
																assign node38969 = (inp[9]) ? 4'b0001 : 4'b0000;
											assign node38972 = (inp[4]) ? node39028 : node38973;
												assign node38973 = (inp[13]) ? node39005 : node38974;
													assign node38974 = (inp[5]) ? node38990 : node38975;
														assign node38975 = (inp[9]) ? node38983 : node38976;
															assign node38976 = (inp[10]) ? node38980 : node38977;
																assign node38977 = (inp[1]) ? 4'b0100 : 4'b0101;
																assign node38980 = (inp[1]) ? 4'b0101 : 4'b0100;
															assign node38983 = (inp[10]) ? node38987 : node38984;
																assign node38984 = (inp[1]) ? 4'b0101 : 4'b0100;
																assign node38987 = (inp[1]) ? 4'b0100 : 4'b0101;
														assign node38990 = (inp[1]) ? node38998 : node38991;
															assign node38991 = (inp[9]) ? node38995 : node38992;
																assign node38992 = (inp[10]) ? 4'b0101 : 4'b0100;
																assign node38995 = (inp[10]) ? 4'b0100 : 4'b0101;
															assign node38998 = (inp[10]) ? node39002 : node38999;
																assign node38999 = (inp[9]) ? 4'b0000 : 4'b0001;
																assign node39002 = (inp[9]) ? 4'b0001 : 4'b0000;
													assign node39005 = (inp[1]) ? node39015 : node39006;
														assign node39006 = (inp[9]) ? 4'b0000 : node39007;
															assign node39007 = (inp[5]) ? node39011 : node39008;
																assign node39008 = (inp[10]) ? 4'b0000 : 4'b0001;
																assign node39011 = (inp[10]) ? 4'b0001 : 4'b0000;
														assign node39015 = (inp[5]) ? node39021 : node39016;
															assign node39016 = (inp[10]) ? node39018 : 4'b0001;
																assign node39018 = (inp[9]) ? 4'b0000 : 4'b0001;
															assign node39021 = (inp[10]) ? node39025 : node39022;
																assign node39022 = (inp[9]) ? 4'b0101 : 4'b0100;
																assign node39025 = (inp[9]) ? 4'b0100 : 4'b0101;
												assign node39028 = (inp[13]) ? node39060 : node39029;
													assign node39029 = (inp[5]) ? node39045 : node39030;
														assign node39030 = (inp[1]) ? node39038 : node39031;
															assign node39031 = (inp[10]) ? node39035 : node39032;
																assign node39032 = (inp[9]) ? 4'b0000 : 4'b0001;
																assign node39035 = (inp[9]) ? 4'b0001 : 4'b0000;
															assign node39038 = (inp[9]) ? node39042 : node39039;
																assign node39039 = (inp[10]) ? 4'b0001 : 4'b0000;
																assign node39042 = (inp[10]) ? 4'b0000 : 4'b0001;
														assign node39045 = (inp[1]) ? node39053 : node39046;
															assign node39046 = (inp[10]) ? node39050 : node39047;
																assign node39047 = (inp[9]) ? 4'b0001 : 4'b0000;
																assign node39050 = (inp[9]) ? 4'b0000 : 4'b0001;
															assign node39053 = (inp[9]) ? node39057 : node39054;
																assign node39054 = (inp[10]) ? 4'b0101 : 4'b0100;
																assign node39057 = (inp[10]) ? 4'b0100 : 4'b0101;
													assign node39060 = (inp[1]) ? node39074 : node39061;
														assign node39061 = (inp[5]) ? node39067 : node39062;
															assign node39062 = (inp[9]) ? 4'b0101 : node39063;
																assign node39063 = (inp[10]) ? 4'b0101 : 4'b0100;
															assign node39067 = (inp[9]) ? node39071 : node39068;
																assign node39068 = (inp[10]) ? 4'b0100 : 4'b0101;
																assign node39071 = (inp[10]) ? 4'b0101 : 4'b0100;
														assign node39074 = (inp[5]) ? node39078 : node39075;
															assign node39075 = (inp[9]) ? 4'b0100 : 4'b0101;
															assign node39078 = (inp[9]) ? node39082 : node39079;
																assign node39079 = (inp[10]) ? 4'b0001 : 4'b0000;
																assign node39082 = (inp[10]) ? 4'b0000 : 4'b0001;
							assign node39085 = (inp[4]) ? node39783 : node39086;
								assign node39086 = (inp[15]) ? node39444 : node39087;
									assign node39087 = (inp[10]) ? node39249 : node39088;
										assign node39088 = (inp[2]) ? node39166 : node39089;
											assign node39089 = (inp[13]) ? node39131 : node39090;
												assign node39090 = (inp[5]) ? node39108 : node39091;
													assign node39091 = (inp[1]) ? node39101 : node39092;
														assign node39092 = (inp[9]) ? node39096 : node39093;
															assign node39093 = (inp[0]) ? 4'b0101 : 4'b0100;
															assign node39096 = (inp[11]) ? 4'b0100 : node39097;
																assign node39097 = (inp[0]) ? 4'b0100 : 4'b0101;
														assign node39101 = (inp[9]) ? node39103 : 4'b0000;
															assign node39103 = (inp[0]) ? node39105 : 4'b0001;
																assign node39105 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node39108 = (inp[9]) ? node39120 : node39109;
														assign node39109 = (inp[0]) ? node39115 : node39110;
															assign node39110 = (inp[11]) ? 4'b0001 : node39111;
																assign node39111 = (inp[1]) ? 4'b0000 : 4'b0001;
															assign node39115 = (inp[1]) ? 4'b0001 : node39116;
																assign node39116 = (inp[11]) ? 4'b0000 : 4'b0001;
														assign node39120 = (inp[0]) ? node39126 : node39121;
															assign node39121 = (inp[1]) ? node39123 : 4'b0000;
																assign node39123 = (inp[11]) ? 4'b0000 : 4'b0001;
															assign node39126 = (inp[11]) ? node39128 : 4'b0000;
																assign node39128 = (inp[1]) ? 4'b0000 : 4'b0001;
												assign node39131 = (inp[1]) ? node39149 : node39132;
													assign node39132 = (inp[5]) ? node39140 : node39133;
														assign node39133 = (inp[9]) ? node39135 : 4'b0000;
															assign node39135 = (inp[11]) ? 4'b0001 : node39136;
																assign node39136 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node39140 = (inp[9]) ? node39144 : node39141;
															assign node39141 = (inp[0]) ? 4'b0101 : 4'b0100;
															assign node39144 = (inp[11]) ? 4'b0100 : node39145;
																assign node39145 = (inp[0]) ? 4'b0100 : 4'b0101;
													assign node39149 = (inp[9]) ? node39157 : node39150;
														assign node39150 = (inp[11]) ? 4'b0100 : node39151;
															assign node39151 = (inp[0]) ? 4'b0100 : node39152;
																assign node39152 = (inp[5]) ? 4'b0100 : 4'b0101;
														assign node39157 = (inp[11]) ? node39163 : node39158;
															assign node39158 = (inp[0]) ? 4'b0101 : node39159;
																assign node39159 = (inp[5]) ? 4'b0101 : 4'b0100;
															assign node39163 = (inp[0]) ? 4'b0100 : 4'b0101;
											assign node39166 = (inp[13]) ? node39208 : node39167;
												assign node39167 = (inp[1]) ? node39189 : node39168;
													assign node39168 = (inp[5]) ? node39178 : node39169;
														assign node39169 = (inp[9]) ? node39173 : node39170;
															assign node39170 = (inp[0]) ? 4'b0000 : 4'b0001;
															assign node39173 = (inp[0]) ? 4'b0001 : node39174;
																assign node39174 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node39178 = (inp[9]) ? node39184 : node39179;
															assign node39179 = (inp[11]) ? 4'b0101 : node39180;
																assign node39180 = (inp[0]) ? 4'b0101 : 4'b0100;
															assign node39184 = (inp[0]) ? 4'b0100 : node39185;
																assign node39185 = (inp[11]) ? 4'b0100 : 4'b0101;
													assign node39189 = (inp[9]) ? node39199 : node39190;
														assign node39190 = (inp[5]) ? node39196 : node39191;
															assign node39191 = (inp[11]) ? 4'b0100 : node39192;
																assign node39192 = (inp[0]) ? 4'b0100 : 4'b0101;
															assign node39196 = (inp[0]) ? 4'b0101 : 4'b0100;
														assign node39199 = (inp[0]) ? node39203 : node39200;
															assign node39200 = (inp[11]) ? 4'b0101 : 4'b0100;
															assign node39203 = (inp[11]) ? node39205 : 4'b0101;
																assign node39205 = (inp[5]) ? 4'b0100 : 4'b0101;
												assign node39208 = (inp[1]) ? node39228 : node39209;
													assign node39209 = (inp[5]) ? node39219 : node39210;
														assign node39210 = (inp[9]) ? node39216 : node39211;
															assign node39211 = (inp[0]) ? node39213 : 4'b0101;
																assign node39213 = (inp[11]) ? 4'b0100 : 4'b0101;
															assign node39216 = (inp[0]) ? 4'b0101 : 4'b0100;
														assign node39219 = (inp[9]) ? node39223 : node39220;
															assign node39220 = (inp[0]) ? 4'b0000 : 4'b0001;
															assign node39223 = (inp[0]) ? 4'b0001 : node39224;
																assign node39224 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node39228 = (inp[9]) ? node39238 : node39229;
														assign node39229 = (inp[0]) ? node39235 : node39230;
															assign node39230 = (inp[5]) ? 4'b0001 : node39231;
																assign node39231 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node39235 = (inp[5]) ? 4'b0000 : 4'b0001;
														assign node39238 = (inp[5]) ? node39244 : node39239;
															assign node39239 = (inp[0]) ? 4'b0000 : node39240;
																assign node39240 = (inp[11]) ? 4'b0000 : 4'b0001;
															assign node39244 = (inp[11]) ? node39246 : 4'b0000;
																assign node39246 = (inp[0]) ? 4'b0001 : 4'b0000;
										assign node39249 = (inp[11]) ? node39345 : node39250;
											assign node39250 = (inp[13]) ? node39296 : node39251;
												assign node39251 = (inp[2]) ? node39271 : node39252;
													assign node39252 = (inp[5]) ? node39262 : node39253;
														assign node39253 = (inp[1]) ? node39259 : node39254;
															assign node39254 = (inp[0]) ? node39256 : 4'b0100;
																assign node39256 = (inp[9]) ? 4'b0101 : 4'b0100;
															assign node39259 = (inp[9]) ? 4'b0000 : 4'b0001;
														assign node39262 = (inp[9]) ? node39268 : node39263;
															assign node39263 = (inp[0]) ? 4'b0000 : node39264;
																assign node39264 = (inp[1]) ? 4'b0001 : 4'b0000;
															assign node39268 = (inp[1]) ? 4'b0000 : 4'b0001;
													assign node39271 = (inp[5]) ? node39285 : node39272;
														assign node39272 = (inp[1]) ? node39280 : node39273;
															assign node39273 = (inp[0]) ? node39277 : node39274;
																assign node39274 = (inp[9]) ? 4'b0001 : 4'b0000;
																assign node39277 = (inp[9]) ? 4'b0000 : 4'b0001;
															assign node39280 = (inp[9]) ? 4'b0100 : node39281;
																assign node39281 = (inp[0]) ? 4'b0101 : 4'b0100;
														assign node39285 = (inp[9]) ? node39291 : node39286;
															assign node39286 = (inp[1]) ? 4'b0101 : node39287;
																assign node39287 = (inp[0]) ? 4'b0100 : 4'b0101;
															assign node39291 = (inp[1]) ? 4'b0100 : node39292;
																assign node39292 = (inp[0]) ? 4'b0101 : 4'b0100;
												assign node39296 = (inp[2]) ? node39322 : node39297;
													assign node39297 = (inp[5]) ? node39311 : node39298;
														assign node39298 = (inp[1]) ? node39304 : node39299;
															assign node39299 = (inp[0]) ? 4'b0001 : node39300;
																assign node39300 = (inp[9]) ? 4'b0001 : 4'b0000;
															assign node39304 = (inp[9]) ? node39308 : node39305;
																assign node39305 = (inp[0]) ? 4'b0101 : 4'b0100;
																assign node39308 = (inp[0]) ? 4'b0100 : 4'b0101;
														assign node39311 = (inp[9]) ? node39317 : node39312;
															assign node39312 = (inp[1]) ? 4'b0101 : node39313;
																assign node39313 = (inp[0]) ? 4'b0100 : 4'b0101;
															assign node39317 = (inp[1]) ? 4'b0100 : node39318;
																assign node39318 = (inp[0]) ? 4'b0101 : 4'b0100;
													assign node39322 = (inp[1]) ? node39334 : node39323;
														assign node39323 = (inp[5]) ? node39327 : node39324;
															assign node39324 = (inp[9]) ? 4'b0101 : 4'b0100;
															assign node39327 = (inp[9]) ? node39331 : node39328;
																assign node39328 = (inp[0]) ? 4'b0001 : 4'b0000;
																assign node39331 = (inp[0]) ? 4'b0000 : 4'b0001;
														assign node39334 = (inp[9]) ? node39340 : node39335;
															assign node39335 = (inp[5]) ? 4'b0000 : node39336;
																assign node39336 = (inp[0]) ? 4'b0000 : 4'b0001;
															assign node39340 = (inp[0]) ? 4'b0001 : node39341;
																assign node39341 = (inp[5]) ? 4'b0001 : 4'b0000;
											assign node39345 = (inp[0]) ? node39397 : node39346;
												assign node39346 = (inp[1]) ? node39376 : node39347;
													assign node39347 = (inp[9]) ? node39361 : node39348;
														assign node39348 = (inp[13]) ? node39356 : node39349;
															assign node39349 = (inp[2]) ? node39353 : node39350;
																assign node39350 = (inp[5]) ? 4'b0000 : 4'b0100;
																assign node39353 = (inp[5]) ? 4'b0100 : 4'b0001;
															assign node39356 = (inp[5]) ? 4'b0001 : node39357;
																assign node39357 = (inp[2]) ? 4'b0100 : 4'b0001;
														assign node39361 = (inp[2]) ? node39369 : node39362;
															assign node39362 = (inp[5]) ? node39366 : node39363;
																assign node39363 = (inp[13]) ? 4'b0000 : 4'b0101;
																assign node39366 = (inp[13]) ? 4'b0101 : 4'b0001;
															assign node39369 = (inp[5]) ? node39373 : node39370;
																assign node39370 = (inp[13]) ? 4'b0101 : 4'b0000;
																assign node39373 = (inp[13]) ? 4'b0000 : 4'b0101;
													assign node39376 = (inp[9]) ? node39388 : node39377;
														assign node39377 = (inp[5]) ? node39383 : node39378;
															assign node39378 = (inp[2]) ? 4'b0101 : node39379;
																assign node39379 = (inp[13]) ? 4'b0101 : 4'b0001;
															assign node39383 = (inp[2]) ? node39385 : 4'b0101;
																assign node39385 = (inp[13]) ? 4'b0000 : 4'b0101;
														assign node39388 = (inp[13]) ? node39394 : node39389;
															assign node39389 = (inp[2]) ? 4'b0100 : node39390;
																assign node39390 = (inp[5]) ? 4'b0001 : 4'b0000;
															assign node39394 = (inp[2]) ? 4'b0001 : 4'b0100;
												assign node39397 = (inp[5]) ? node39425 : node39398;
													assign node39398 = (inp[1]) ? node39410 : node39399;
														assign node39399 = (inp[9]) ? node39403 : node39400;
															assign node39400 = (inp[13]) ? 4'b0101 : 4'b0100;
															assign node39403 = (inp[2]) ? node39407 : node39404;
																assign node39404 = (inp[13]) ? 4'b0000 : 4'b0101;
																assign node39407 = (inp[13]) ? 4'b0100 : 4'b0000;
														assign node39410 = (inp[9]) ? node39418 : node39411;
															assign node39411 = (inp[2]) ? node39415 : node39412;
																assign node39412 = (inp[13]) ? 4'b0101 : 4'b0000;
																assign node39415 = (inp[13]) ? 4'b0000 : 4'b0101;
															assign node39418 = (inp[13]) ? node39422 : node39419;
																assign node39419 = (inp[2]) ? 4'b0100 : 4'b0001;
																assign node39422 = (inp[2]) ? 4'b0001 : 4'b0100;
													assign node39425 = (inp[9]) ? node39435 : node39426;
														assign node39426 = (inp[2]) ? node39432 : node39427;
															assign node39427 = (inp[13]) ? 4'b0100 : node39428;
																assign node39428 = (inp[1]) ? 4'b0000 : 4'b0001;
															assign node39432 = (inp[13]) ? 4'b0001 : 4'b0100;
														assign node39435 = (inp[13]) ? node39441 : node39436;
															assign node39436 = (inp[2]) ? 4'b0101 : node39437;
																assign node39437 = (inp[1]) ? 4'b0001 : 4'b0000;
															assign node39441 = (inp[2]) ? 4'b0000 : 4'b0101;
									assign node39444 = (inp[10]) ? node39598 : node39445;
										assign node39445 = (inp[1]) ? node39523 : node39446;
											assign node39446 = (inp[5]) ? node39488 : node39447;
												assign node39447 = (inp[9]) ? node39469 : node39448;
													assign node39448 = (inp[0]) ? node39462 : node39449;
														assign node39449 = (inp[13]) ? node39455 : node39450;
															assign node39450 = (inp[2]) ? node39452 : 4'b0010;
																assign node39452 = (inp[11]) ? 4'b0110 : 4'b0111;
															assign node39455 = (inp[2]) ? node39459 : node39456;
																assign node39456 = (inp[11]) ? 4'b0111 : 4'b0110;
																assign node39459 = (inp[11]) ? 4'b0010 : 4'b0011;
														assign node39462 = (inp[2]) ? node39466 : node39463;
															assign node39463 = (inp[11]) ? 4'b0011 : 4'b0010;
															assign node39466 = (inp[13]) ? 4'b0010 : 4'b0110;
													assign node39469 = (inp[2]) ? node39481 : node39470;
														assign node39470 = (inp[13]) ? node39476 : node39471;
															assign node39471 = (inp[11]) ? node39473 : 4'b0011;
																assign node39473 = (inp[0]) ? 4'b0010 : 4'b0011;
															assign node39476 = (inp[0]) ? 4'b0110 : node39477;
																assign node39477 = (inp[11]) ? 4'b0110 : 4'b0111;
														assign node39481 = (inp[13]) ? node39483 : 4'b0110;
															assign node39483 = (inp[11]) ? 4'b0011 : node39484;
																assign node39484 = (inp[0]) ? 4'b0011 : 4'b0010;
												assign node39488 = (inp[9]) ? node39510 : node39489;
													assign node39489 = (inp[0]) ? node39497 : node39490;
														assign node39490 = (inp[2]) ? node39494 : node39491;
															assign node39491 = (inp[13]) ? 4'b0011 : 4'b0111;
															assign node39494 = (inp[11]) ? 4'b0111 : 4'b0110;
														assign node39497 = (inp[11]) ? node39503 : node39498;
															assign node39498 = (inp[2]) ? 4'b0010 : node39499;
																assign node39499 = (inp[13]) ? 4'b0011 : 4'b0111;
															assign node39503 = (inp[2]) ? node39507 : node39504;
																assign node39504 = (inp[13]) ? 4'b0010 : 4'b0110;
																assign node39507 = (inp[13]) ? 4'b0111 : 4'b0011;
													assign node39510 = (inp[13]) ? node39518 : node39511;
														assign node39511 = (inp[2]) ? 4'b0011 : node39512;
															assign node39512 = (inp[0]) ? node39514 : 4'b0110;
																assign node39514 = (inp[11]) ? 4'b0111 : 4'b0110;
														assign node39518 = (inp[2]) ? 4'b0110 : node39519;
															assign node39519 = (inp[0]) ? 4'b0011 : 4'b0010;
											assign node39523 = (inp[9]) ? node39565 : node39524;
												assign node39524 = (inp[2]) ? node39546 : node39525;
													assign node39525 = (inp[13]) ? node39535 : node39526;
														assign node39526 = (inp[5]) ? node39530 : node39527;
															assign node39527 = (inp[11]) ? 4'b0110 : 4'b0111;
															assign node39530 = (inp[0]) ? node39532 : 4'b0110;
																assign node39532 = (inp[11]) ? 4'b0111 : 4'b0110;
														assign node39535 = (inp[5]) ? node39541 : node39536;
															assign node39536 = (inp[11]) ? 4'b0010 : node39537;
																assign node39537 = (inp[0]) ? 4'b0010 : 4'b0011;
															assign node39541 = (inp[11]) ? node39543 : 4'b0010;
																assign node39543 = (inp[0]) ? 4'b0011 : 4'b0010;
													assign node39546 = (inp[13]) ? node39554 : node39547;
														assign node39547 = (inp[11]) ? node39549 : 4'b0011;
															assign node39549 = (inp[0]) ? node39551 : 4'b0011;
																assign node39551 = (inp[5]) ? 4'b0010 : 4'b0011;
														assign node39554 = (inp[5]) ? node39560 : node39555;
															assign node39555 = (inp[0]) ? node39557 : 4'b0111;
																assign node39557 = (inp[11]) ? 4'b0110 : 4'b0111;
															assign node39560 = (inp[0]) ? 4'b0110 : node39561;
																assign node39561 = (inp[11]) ? 4'b0110 : 4'b0111;
												assign node39565 = (inp[2]) ? node39585 : node39566;
													assign node39566 = (inp[13]) ? node39574 : node39567;
														assign node39567 = (inp[11]) ? 4'b0111 : node39568;
															assign node39568 = (inp[5]) ? 4'b0111 : node39569;
																assign node39569 = (inp[0]) ? 4'b0111 : 4'b0110;
														assign node39574 = (inp[0]) ? node39580 : node39575;
															assign node39575 = (inp[5]) ? 4'b0011 : node39576;
																assign node39576 = (inp[11]) ? 4'b0011 : 4'b0010;
															assign node39580 = (inp[11]) ? node39582 : 4'b0011;
																assign node39582 = (inp[5]) ? 4'b0010 : 4'b0011;
													assign node39585 = (inp[13]) ? node39593 : node39586;
														assign node39586 = (inp[5]) ? node39588 : 4'b0010;
															assign node39588 = (inp[11]) ? node39590 : 4'b0010;
																assign node39590 = (inp[0]) ? 4'b0011 : 4'b0010;
														assign node39593 = (inp[11]) ? 4'b0111 : node39594;
															assign node39594 = (inp[0]) ? 4'b0111 : 4'b0110;
										assign node39598 = (inp[11]) ? node39684 : node39599;
											assign node39599 = (inp[5]) ? node39653 : node39600;
												assign node39600 = (inp[2]) ? node39626 : node39601;
													assign node39601 = (inp[9]) ? node39613 : node39602;
														assign node39602 = (inp[13]) ? node39608 : node39603;
															assign node39603 = (inp[0]) ? node39605 : 4'b0110;
																assign node39605 = (inp[1]) ? 4'b0111 : 4'b0011;
															assign node39608 = (inp[1]) ? 4'b0010 : node39609;
																assign node39609 = (inp[0]) ? 4'b0110 : 4'b0111;
														assign node39613 = (inp[0]) ? node39621 : node39614;
															assign node39614 = (inp[1]) ? node39618 : node39615;
																assign node39615 = (inp[13]) ? 4'b0110 : 4'b0010;
																assign node39618 = (inp[13]) ? 4'b0011 : 4'b0111;
															assign node39621 = (inp[1]) ? node39623 : 4'b0111;
																assign node39623 = (inp[13]) ? 4'b0010 : 4'b0110;
													assign node39626 = (inp[9]) ? node39642 : node39627;
														assign node39627 = (inp[0]) ? node39635 : node39628;
															assign node39628 = (inp[1]) ? node39632 : node39629;
																assign node39629 = (inp[13]) ? 4'b0010 : 4'b0110;
																assign node39632 = (inp[13]) ? 4'b0110 : 4'b0011;
															assign node39635 = (inp[1]) ? node39639 : node39636;
																assign node39636 = (inp[13]) ? 4'b0011 : 4'b0111;
																assign node39639 = (inp[13]) ? 4'b0110 : 4'b0010;
														assign node39642 = (inp[0]) ? node39648 : node39643;
															assign node39643 = (inp[1]) ? node39645 : 4'b0111;
																assign node39645 = (inp[13]) ? 4'b0111 : 4'b0010;
															assign node39648 = (inp[1]) ? 4'b0111 : node39649;
																assign node39649 = (inp[13]) ? 4'b0010 : 4'b0110;
												assign node39653 = (inp[2]) ? node39669 : node39654;
													assign node39654 = (inp[13]) ? node39662 : node39655;
														assign node39655 = (inp[1]) ? node39659 : node39656;
															assign node39656 = (inp[9]) ? 4'b0111 : 4'b0110;
															assign node39659 = (inp[9]) ? 4'b0110 : 4'b0111;
														assign node39662 = (inp[1]) ? node39666 : node39663;
															assign node39663 = (inp[9]) ? 4'b0011 : 4'b0010;
															assign node39666 = (inp[9]) ? 4'b0010 : 4'b0011;
													assign node39669 = (inp[13]) ? node39677 : node39670;
														assign node39670 = (inp[9]) ? node39674 : node39671;
															assign node39671 = (inp[1]) ? 4'b0010 : 4'b0011;
															assign node39674 = (inp[1]) ? 4'b0011 : 4'b0010;
														assign node39677 = (inp[9]) ? 4'b0111 : node39678;
															assign node39678 = (inp[0]) ? 4'b0110 : node39679;
																assign node39679 = (inp[1]) ? 4'b0110 : 4'b0111;
											assign node39684 = (inp[9]) ? node39734 : node39685;
												assign node39685 = (inp[5]) ? node39705 : node39686;
													assign node39686 = (inp[1]) ? node39696 : node39687;
														assign node39687 = (inp[2]) ? node39693 : node39688;
															assign node39688 = (inp[13]) ? 4'b0110 : node39689;
																assign node39689 = (inp[0]) ? 4'b0010 : 4'b0011;
															assign node39693 = (inp[13]) ? 4'b0011 : 4'b0111;
														assign node39696 = (inp[2]) ? node39700 : node39697;
															assign node39697 = (inp[13]) ? 4'b0011 : 4'b0111;
															assign node39700 = (inp[13]) ? node39702 : 4'b0010;
																assign node39702 = (inp[0]) ? 4'b0111 : 4'b0110;
													assign node39705 = (inp[1]) ? node39719 : node39706;
														assign node39706 = (inp[0]) ? node39714 : node39707;
															assign node39707 = (inp[13]) ? node39711 : node39708;
																assign node39708 = (inp[2]) ? 4'b0011 : 4'b0110;
																assign node39711 = (inp[2]) ? 4'b0110 : 4'b0010;
															assign node39714 = (inp[2]) ? 4'b0110 : node39715;
																assign node39715 = (inp[13]) ? 4'b0011 : 4'b0111;
														assign node39719 = (inp[0]) ? node39727 : node39720;
															assign node39720 = (inp[2]) ? node39724 : node39721;
																assign node39721 = (inp[13]) ? 4'b0011 : 4'b0111;
																assign node39724 = (inp[13]) ? 4'b0111 : 4'b0010;
															assign node39727 = (inp[2]) ? node39731 : node39728;
																assign node39728 = (inp[13]) ? 4'b0010 : 4'b0110;
																assign node39731 = (inp[13]) ? 4'b0111 : 4'b0011;
												assign node39734 = (inp[1]) ? node39762 : node39735;
													assign node39735 = (inp[13]) ? node39749 : node39736;
														assign node39736 = (inp[5]) ? node39742 : node39737;
															assign node39737 = (inp[2]) ? 4'b0110 : node39738;
																assign node39738 = (inp[0]) ? 4'b0011 : 4'b0010;
															assign node39742 = (inp[2]) ? node39746 : node39743;
																assign node39743 = (inp[0]) ? 4'b0110 : 4'b0111;
																assign node39746 = (inp[0]) ? 4'b0011 : 4'b0010;
														assign node39749 = (inp[0]) ? node39755 : node39750;
															assign node39750 = (inp[5]) ? node39752 : 4'b0111;
																assign node39752 = (inp[2]) ? 4'b0111 : 4'b0011;
															assign node39755 = (inp[2]) ? node39759 : node39756;
																assign node39756 = (inp[5]) ? 4'b0010 : 4'b0111;
																assign node39759 = (inp[5]) ? 4'b0111 : 4'b0010;
													assign node39762 = (inp[0]) ? node39770 : node39763;
														assign node39763 = (inp[2]) ? node39767 : node39764;
															assign node39764 = (inp[13]) ? 4'b0010 : 4'b0110;
															assign node39767 = (inp[5]) ? 4'b0110 : 4'b0111;
														assign node39770 = (inp[2]) ? node39778 : node39771;
															assign node39771 = (inp[13]) ? node39775 : node39772;
																assign node39772 = (inp[5]) ? 4'b0111 : 4'b0110;
																assign node39775 = (inp[5]) ? 4'b0011 : 4'b0010;
															assign node39778 = (inp[5]) ? node39780 : 4'b0011;
																assign node39780 = (inp[13]) ? 4'b0110 : 4'b0010;
								assign node39783 = (inp[11]) ? node40103 : node39784;
									assign node39784 = (inp[10]) ? node39956 : node39785;
										assign node39785 = (inp[9]) ? node39875 : node39786;
											assign node39786 = (inp[1]) ? node39840 : node39787;
												assign node39787 = (inp[0]) ? node39809 : node39788;
													assign node39788 = (inp[15]) ? node39802 : node39789;
														assign node39789 = (inp[13]) ? node39795 : node39790;
															assign node39790 = (inp[2]) ? node39792 : 4'b0010;
																assign node39792 = (inp[5]) ? 4'b0111 : 4'b0010;
															assign node39795 = (inp[2]) ? node39799 : node39796;
																assign node39796 = (inp[5]) ? 4'b0110 : 4'b0011;
																assign node39799 = (inp[5]) ? 4'b0010 : 4'b0110;
														assign node39802 = (inp[5]) ? 4'b0010 : node39803;
															assign node39803 = (inp[2]) ? 4'b0110 : node39804;
																assign node39804 = (inp[13]) ? 4'b0010 : 4'b0110;
													assign node39809 = (inp[13]) ? node39825 : node39810;
														assign node39810 = (inp[15]) ? node39818 : node39811;
															assign node39811 = (inp[5]) ? node39815 : node39812;
																assign node39812 = (inp[2]) ? 4'b0011 : 4'b0111;
																assign node39815 = (inp[2]) ? 4'b0111 : 4'b0011;
															assign node39818 = (inp[2]) ? node39822 : node39819;
																assign node39819 = (inp[5]) ? 4'b0010 : 4'b0110;
																assign node39822 = (inp[5]) ? 4'b0111 : 4'b0010;
														assign node39825 = (inp[15]) ? node39833 : node39826;
															assign node39826 = (inp[5]) ? node39830 : node39827;
																assign node39827 = (inp[2]) ? 4'b0110 : 4'b0010;
																assign node39830 = (inp[2]) ? 4'b0010 : 4'b0110;
															assign node39833 = (inp[5]) ? node39837 : node39834;
																assign node39834 = (inp[2]) ? 4'b0111 : 4'b0010;
																assign node39837 = (inp[2]) ? 4'b0011 : 4'b0111;
												assign node39840 = (inp[0]) ? node39864 : node39841;
													assign node39841 = (inp[15]) ? node39849 : node39842;
														assign node39842 = (inp[13]) ? node39846 : node39843;
															assign node39843 = (inp[2]) ? 4'b0110 : 4'b0010;
															assign node39846 = (inp[2]) ? 4'b0011 : 4'b0111;
														assign node39849 = (inp[5]) ? node39857 : node39850;
															assign node39850 = (inp[13]) ? node39854 : node39851;
																assign node39851 = (inp[2]) ? 4'b0111 : 4'b0011;
																assign node39854 = (inp[2]) ? 4'b0011 : 4'b0111;
															assign node39857 = (inp[2]) ? node39861 : node39858;
																assign node39858 = (inp[13]) ? 4'b0111 : 4'b0011;
																assign node39861 = (inp[13]) ? 4'b0011 : 4'b0111;
													assign node39864 = (inp[13]) ? node39872 : node39865;
														assign node39865 = (inp[2]) ? node39869 : node39866;
															assign node39866 = (inp[15]) ? 4'b0011 : 4'b0010;
															assign node39869 = (inp[15]) ? 4'b0110 : 4'b0111;
														assign node39872 = (inp[2]) ? 4'b0010 : 4'b0110;
											assign node39875 = (inp[1]) ? node39933 : node39876;
												assign node39876 = (inp[0]) ? node39906 : node39877;
													assign node39877 = (inp[15]) ? node39891 : node39878;
														assign node39878 = (inp[13]) ? node39886 : node39879;
															assign node39879 = (inp[5]) ? node39883 : node39880;
																assign node39880 = (inp[2]) ? 4'b0011 : 4'b0111;
																assign node39883 = (inp[2]) ? 4'b0110 : 4'b0011;
															assign node39886 = (inp[5]) ? node39888 : 4'b0111;
																assign node39888 = (inp[2]) ? 4'b0011 : 4'b0111;
														assign node39891 = (inp[5]) ? node39899 : node39892;
															assign node39892 = (inp[13]) ? node39896 : node39893;
																assign node39893 = (inp[2]) ? 4'b0011 : 4'b0111;
																assign node39896 = (inp[2]) ? 4'b0111 : 4'b0011;
															assign node39899 = (inp[13]) ? node39903 : node39900;
																assign node39900 = (inp[2]) ? 4'b0111 : 4'b0011;
																assign node39903 = (inp[2]) ? 4'b0011 : 4'b0111;
													assign node39906 = (inp[5]) ? node39920 : node39907;
														assign node39907 = (inp[2]) ? node39913 : node39908;
															assign node39908 = (inp[13]) ? 4'b0011 : node39909;
																assign node39909 = (inp[15]) ? 4'b0111 : 4'b0110;
															assign node39913 = (inp[13]) ? node39917 : node39914;
																assign node39914 = (inp[15]) ? 4'b0011 : 4'b0010;
																assign node39917 = (inp[15]) ? 4'b0110 : 4'b0111;
														assign node39920 = (inp[13]) ? node39926 : node39921;
															assign node39921 = (inp[2]) ? 4'b0110 : node39922;
																assign node39922 = (inp[15]) ? 4'b0011 : 4'b0010;
															assign node39926 = (inp[2]) ? node39930 : node39927;
																assign node39927 = (inp[15]) ? 4'b0110 : 4'b0111;
																assign node39930 = (inp[15]) ? 4'b0010 : 4'b0011;
												assign node39933 = (inp[0]) ? node39945 : node39934;
													assign node39934 = (inp[13]) ? node39942 : node39935;
														assign node39935 = (inp[2]) ? node39939 : node39936;
															assign node39936 = (inp[15]) ? 4'b0010 : 4'b0011;
															assign node39939 = (inp[15]) ? 4'b0110 : 4'b0111;
														assign node39942 = (inp[2]) ? 4'b0010 : 4'b0110;
													assign node39945 = (inp[13]) ? node39953 : node39946;
														assign node39946 = (inp[2]) ? node39950 : node39947;
															assign node39947 = (inp[15]) ? 4'b0010 : 4'b0011;
															assign node39950 = (inp[15]) ? 4'b0111 : 4'b0110;
														assign node39953 = (inp[2]) ? 4'b0011 : 4'b0111;
										assign node39956 = (inp[9]) ? node40026 : node39957;
											assign node39957 = (inp[1]) ? node40003 : node39958;
												assign node39958 = (inp[0]) ? node39978 : node39959;
													assign node39959 = (inp[15]) ? node39969 : node39960;
														assign node39960 = (inp[2]) ? 4'b0011 : node39961;
															assign node39961 = (inp[13]) ? node39965 : node39962;
																assign node39962 = (inp[5]) ? 4'b0011 : 4'b0111;
																assign node39965 = (inp[5]) ? 4'b0111 : 4'b0010;
														assign node39969 = (inp[13]) ? node39971 : 4'b0111;
															assign node39971 = (inp[5]) ? node39975 : node39972;
																assign node39972 = (inp[2]) ? 4'b0111 : 4'b0011;
																assign node39975 = (inp[2]) ? 4'b0011 : 4'b0111;
													assign node39978 = (inp[13]) ? node39994 : node39979;
														assign node39979 = (inp[15]) ? node39987 : node39980;
															assign node39980 = (inp[5]) ? node39984 : node39981;
																assign node39981 = (inp[2]) ? 4'b0010 : 4'b0110;
																assign node39984 = (inp[2]) ? 4'b0110 : 4'b0010;
															assign node39987 = (inp[5]) ? node39991 : node39988;
																assign node39988 = (inp[2]) ? 4'b0011 : 4'b0111;
																assign node39991 = (inp[2]) ? 4'b0110 : 4'b0011;
														assign node39994 = (inp[2]) ? node39996 : 4'b0011;
															assign node39996 = (inp[15]) ? node40000 : node39997;
																assign node39997 = (inp[5]) ? 4'b0011 : 4'b0111;
																assign node40000 = (inp[5]) ? 4'b0010 : 4'b0110;
												assign node40003 = (inp[0]) ? node40015 : node40004;
													assign node40004 = (inp[13]) ? node40012 : node40005;
														assign node40005 = (inp[15]) ? node40009 : node40006;
															assign node40006 = (inp[2]) ? 4'b0111 : 4'b0011;
															assign node40009 = (inp[2]) ? 4'b0110 : 4'b0010;
														assign node40012 = (inp[2]) ? 4'b0010 : 4'b0110;
													assign node40015 = (inp[13]) ? node40023 : node40016;
														assign node40016 = (inp[2]) ? node40020 : node40017;
															assign node40017 = (inp[15]) ? 4'b0010 : 4'b0011;
															assign node40020 = (inp[15]) ? 4'b0111 : 4'b0110;
														assign node40023 = (inp[2]) ? 4'b0011 : 4'b0111;
											assign node40026 = (inp[1]) ? node40080 : node40027;
												assign node40027 = (inp[0]) ? node40059 : node40028;
													assign node40028 = (inp[15]) ? node40044 : node40029;
														assign node40029 = (inp[13]) ? node40037 : node40030;
															assign node40030 = (inp[5]) ? node40034 : node40031;
																assign node40031 = (inp[2]) ? 4'b0010 : 4'b0110;
																assign node40034 = (inp[2]) ? 4'b0111 : 4'b0010;
															assign node40037 = (inp[2]) ? node40041 : node40038;
																assign node40038 = (inp[5]) ? 4'b0110 : 4'b0011;
																assign node40041 = (inp[5]) ? 4'b0010 : 4'b0110;
														assign node40044 = (inp[5]) ? node40052 : node40045;
															assign node40045 = (inp[2]) ? node40049 : node40046;
																assign node40046 = (inp[13]) ? 4'b0010 : 4'b0110;
																assign node40049 = (inp[13]) ? 4'b0110 : 4'b0010;
															assign node40052 = (inp[13]) ? node40056 : node40053;
																assign node40053 = (inp[2]) ? 4'b0110 : 4'b0010;
																assign node40056 = (inp[2]) ? 4'b0010 : 4'b0110;
													assign node40059 = (inp[2]) ? node40069 : node40060;
														assign node40060 = (inp[5]) ? node40062 : 4'b0010;
															assign node40062 = (inp[13]) ? node40066 : node40063;
																assign node40063 = (inp[15]) ? 4'b0010 : 4'b0011;
																assign node40066 = (inp[15]) ? 4'b0111 : 4'b0110;
														assign node40069 = (inp[13]) ? node40073 : node40070;
															assign node40070 = (inp[5]) ? 4'b0111 : 4'b0011;
															assign node40073 = (inp[15]) ? node40077 : node40074;
																assign node40074 = (inp[5]) ? 4'b0010 : 4'b0110;
																assign node40077 = (inp[5]) ? 4'b0011 : 4'b0111;
												assign node40080 = (inp[0]) ? node40092 : node40081;
													assign node40081 = (inp[13]) ? node40089 : node40082;
														assign node40082 = (inp[2]) ? node40086 : node40083;
															assign node40083 = (inp[15]) ? 4'b0011 : 4'b0010;
															assign node40086 = (inp[15]) ? 4'b0111 : 4'b0110;
														assign node40089 = (inp[2]) ? 4'b0011 : 4'b0111;
													assign node40092 = (inp[13]) ? node40100 : node40093;
														assign node40093 = (inp[2]) ? node40097 : node40094;
															assign node40094 = (inp[15]) ? 4'b0011 : 4'b0010;
															assign node40097 = (inp[15]) ? 4'b0110 : 4'b0111;
														assign node40100 = (inp[2]) ? 4'b0010 : 4'b0110;
									assign node40103 = (inp[13]) ? node40287 : node40104;
										assign node40104 = (inp[2]) ? node40196 : node40105;
											assign node40105 = (inp[1]) ? node40149 : node40106;
												assign node40106 = (inp[5]) ? node40128 : node40107;
													assign node40107 = (inp[15]) ? node40115 : node40108;
														assign node40108 = (inp[9]) ? node40112 : node40109;
															assign node40109 = (inp[10]) ? 4'b0110 : 4'b0111;
															assign node40112 = (inp[10]) ? 4'b0111 : 4'b0110;
														assign node40115 = (inp[0]) ? node40123 : node40116;
															assign node40116 = (inp[10]) ? node40120 : node40117;
																assign node40117 = (inp[9]) ? 4'b0111 : 4'b0110;
																assign node40120 = (inp[9]) ? 4'b0110 : 4'b0111;
															assign node40123 = (inp[10]) ? node40125 : 4'b0111;
																assign node40125 = (inp[9]) ? 4'b0111 : 4'b0110;
													assign node40128 = (inp[0]) ? node40142 : node40129;
														assign node40129 = (inp[10]) ? node40135 : node40130;
															assign node40130 = (inp[15]) ? 4'b0011 : node40131;
																assign node40131 = (inp[9]) ? 4'b0010 : 4'b0011;
															assign node40135 = (inp[9]) ? node40139 : node40136;
																assign node40136 = (inp[15]) ? 4'b0011 : 4'b0010;
																assign node40139 = (inp[15]) ? 4'b0010 : 4'b0011;
														assign node40142 = (inp[10]) ? node40146 : node40143;
															assign node40143 = (inp[9]) ? 4'b0010 : 4'b0011;
															assign node40146 = (inp[9]) ? 4'b0011 : 4'b0010;
												assign node40149 = (inp[15]) ? node40165 : node40150;
													assign node40150 = (inp[9]) ? node40158 : node40151;
														assign node40151 = (inp[0]) ? node40155 : node40152;
															assign node40152 = (inp[10]) ? 4'b0011 : 4'b0010;
															assign node40155 = (inp[10]) ? 4'b0010 : 4'b0011;
														assign node40158 = (inp[10]) ? node40162 : node40159;
															assign node40159 = (inp[0]) ? 4'b0010 : 4'b0011;
															assign node40162 = (inp[0]) ? 4'b0011 : 4'b0010;
													assign node40165 = (inp[10]) ? node40181 : node40166;
														assign node40166 = (inp[5]) ? node40174 : node40167;
															assign node40167 = (inp[0]) ? node40171 : node40168;
																assign node40168 = (inp[9]) ? 4'b0010 : 4'b0011;
																assign node40171 = (inp[9]) ? 4'b0011 : 4'b0010;
															assign node40174 = (inp[0]) ? node40178 : node40175;
																assign node40175 = (inp[9]) ? 4'b0010 : 4'b0011;
																assign node40178 = (inp[9]) ? 4'b0011 : 4'b0010;
														assign node40181 = (inp[5]) ? node40189 : node40182;
															assign node40182 = (inp[9]) ? node40186 : node40183;
																assign node40183 = (inp[0]) ? 4'b0011 : 4'b0010;
																assign node40186 = (inp[0]) ? 4'b0010 : 4'b0011;
															assign node40189 = (inp[0]) ? node40193 : node40190;
																assign node40190 = (inp[9]) ? 4'b0011 : 4'b0010;
																assign node40193 = (inp[9]) ? 4'b0010 : 4'b0011;
											assign node40196 = (inp[1]) ? node40242 : node40197;
												assign node40197 = (inp[5]) ? node40221 : node40198;
													assign node40198 = (inp[9]) ? node40210 : node40199;
														assign node40199 = (inp[10]) ? node40205 : node40200;
															assign node40200 = (inp[15]) ? node40202 : 4'b0011;
																assign node40202 = (inp[0]) ? 4'b0011 : 4'b0010;
															assign node40205 = (inp[0]) ? 4'b0010 : node40206;
																assign node40206 = (inp[15]) ? 4'b0011 : 4'b0010;
														assign node40210 = (inp[10]) ? node40216 : node40211;
															assign node40211 = (inp[0]) ? 4'b0010 : node40212;
																assign node40212 = (inp[15]) ? 4'b0011 : 4'b0010;
															assign node40216 = (inp[0]) ? 4'b0011 : node40217;
																assign node40217 = (inp[15]) ? 4'b0010 : 4'b0011;
													assign node40221 = (inp[9]) ? node40233 : node40222;
														assign node40222 = (inp[10]) ? node40228 : node40223;
															assign node40223 = (inp[15]) ? 4'b0111 : node40224;
																assign node40224 = (inp[0]) ? 4'b0110 : 4'b0111;
															assign node40228 = (inp[15]) ? 4'b0110 : node40229;
																assign node40229 = (inp[0]) ? 4'b0111 : 4'b0110;
														assign node40233 = (inp[0]) ? node40235 : 4'b0111;
															assign node40235 = (inp[10]) ? node40239 : node40236;
																assign node40236 = (inp[15]) ? 4'b0110 : 4'b0111;
																assign node40239 = (inp[15]) ? 4'b0111 : 4'b0110;
												assign node40242 = (inp[0]) ? node40272 : node40243;
													assign node40243 = (inp[5]) ? node40259 : node40244;
														assign node40244 = (inp[9]) ? node40252 : node40245;
															assign node40245 = (inp[15]) ? node40249 : node40246;
																assign node40246 = (inp[10]) ? 4'b0110 : 4'b0111;
																assign node40249 = (inp[10]) ? 4'b0111 : 4'b0110;
															assign node40252 = (inp[15]) ? node40256 : node40253;
																assign node40253 = (inp[10]) ? 4'b0111 : 4'b0110;
																assign node40256 = (inp[10]) ? 4'b0110 : 4'b0111;
														assign node40259 = (inp[9]) ? node40265 : node40260;
															assign node40260 = (inp[10]) ? 4'b0111 : node40261;
																assign node40261 = (inp[15]) ? 4'b0110 : 4'b0111;
															assign node40265 = (inp[10]) ? node40269 : node40266;
																assign node40266 = (inp[15]) ? 4'b0111 : 4'b0110;
																assign node40269 = (inp[15]) ? 4'b0110 : 4'b0111;
													assign node40272 = (inp[9]) ? node40280 : node40273;
														assign node40273 = (inp[15]) ? node40277 : node40274;
															assign node40274 = (inp[10]) ? 4'b0110 : 4'b0111;
															assign node40277 = (inp[10]) ? 4'b0111 : 4'b0110;
														assign node40280 = (inp[15]) ? node40284 : node40281;
															assign node40281 = (inp[10]) ? 4'b0111 : 4'b0110;
															assign node40284 = (inp[10]) ? 4'b0110 : 4'b0111;
										assign node40287 = (inp[2]) ? node40353 : node40288;
											assign node40288 = (inp[1]) ? node40322 : node40289;
												assign node40289 = (inp[5]) ? node40307 : node40290;
													assign node40290 = (inp[10]) ? node40298 : node40291;
														assign node40291 = (inp[9]) ? 4'b0011 : node40292;
															assign node40292 = (inp[15]) ? node40294 : 4'b0010;
																assign node40294 = (inp[0]) ? 4'b0011 : 4'b0010;
														assign node40298 = (inp[9]) ? node40302 : node40299;
															assign node40299 = (inp[0]) ? 4'b0010 : 4'b0011;
															assign node40302 = (inp[15]) ? node40304 : 4'b0010;
																assign node40304 = (inp[0]) ? 4'b0011 : 4'b0010;
													assign node40307 = (inp[10]) ? node40313 : node40308;
														assign node40308 = (inp[9]) ? 4'b0110 : node40309;
															assign node40309 = (inp[15]) ? 4'b0111 : 4'b0110;
														assign node40313 = (inp[15]) ? node40319 : node40314;
															assign node40314 = (inp[9]) ? 4'b0110 : node40315;
																assign node40315 = (inp[0]) ? 4'b0110 : 4'b0111;
															assign node40319 = (inp[9]) ? 4'b0111 : 4'b0110;
												assign node40322 = (inp[0]) ? node40346 : node40323;
													assign node40323 = (inp[15]) ? node40339 : node40324;
														assign node40324 = (inp[5]) ? node40332 : node40325;
															assign node40325 = (inp[10]) ? node40329 : node40326;
																assign node40326 = (inp[9]) ? 4'b0111 : 4'b0110;
																assign node40329 = (inp[9]) ? 4'b0110 : 4'b0111;
															assign node40332 = (inp[10]) ? node40336 : node40333;
																assign node40333 = (inp[9]) ? 4'b0111 : 4'b0110;
																assign node40336 = (inp[9]) ? 4'b0110 : 4'b0111;
														assign node40339 = (inp[5]) ? 4'b0110 : node40340;
															assign node40340 = (inp[9]) ? node40342 : 4'b0110;
																assign node40342 = (inp[10]) ? 4'b0110 : 4'b0111;
													assign node40346 = (inp[9]) ? node40350 : node40347;
														assign node40347 = (inp[10]) ? 4'b0111 : 4'b0110;
														assign node40350 = (inp[10]) ? 4'b0110 : 4'b0111;
											assign node40353 = (inp[5]) ? node40383 : node40354;
												assign node40354 = (inp[1]) ? node40370 : node40355;
													assign node40355 = (inp[10]) ? node40365 : node40356;
														assign node40356 = (inp[9]) ? node40362 : node40357;
															assign node40357 = (inp[15]) ? 4'b0111 : node40358;
																assign node40358 = (inp[0]) ? 4'b0111 : 4'b0110;
															assign node40362 = (inp[0]) ? 4'b0110 : 4'b0111;
														assign node40365 = (inp[9]) ? node40367 : 4'b0110;
															assign node40367 = (inp[0]) ? 4'b0111 : 4'b0110;
													assign node40370 = (inp[15]) ? node40376 : node40371;
														assign node40371 = (inp[10]) ? 4'b0010 : node40372;
															assign node40372 = (inp[9]) ? 4'b0011 : 4'b0010;
														assign node40376 = (inp[10]) ? node40380 : node40377;
															assign node40377 = (inp[9]) ? 4'b0011 : 4'b0010;
															assign node40380 = (inp[9]) ? 4'b0010 : 4'b0011;
												assign node40383 = (inp[9]) ? node40399 : node40384;
													assign node40384 = (inp[10]) ? node40392 : node40385;
														assign node40385 = (inp[1]) ? 4'b0010 : node40386;
															assign node40386 = (inp[0]) ? 4'b0011 : node40387;
																assign node40387 = (inp[15]) ? 4'b0011 : 4'b0010;
														assign node40392 = (inp[1]) ? 4'b0011 : node40393;
															assign node40393 = (inp[15]) ? 4'b0010 : node40394;
																assign node40394 = (inp[0]) ? 4'b0010 : 4'b0011;
													assign node40399 = (inp[10]) ? node40407 : node40400;
														assign node40400 = (inp[1]) ? 4'b0011 : node40401;
															assign node40401 = (inp[15]) ? 4'b0010 : node40402;
																assign node40402 = (inp[0]) ? 4'b0010 : 4'b0011;
														assign node40407 = (inp[1]) ? 4'b0010 : node40408;
															assign node40408 = (inp[15]) ? 4'b0011 : node40409;
																assign node40409 = (inp[0]) ? 4'b0011 : 4'b0010;
						assign node40414 = (inp[4]) ? node41216 : node40415;
							assign node40415 = (inp[2]) ? node40791 : node40416;
								assign node40416 = (inp[15]) ? node40562 : node40417;
									assign node40417 = (inp[10]) ? node40495 : node40418;
										assign node40418 = (inp[13]) ? node40470 : node40419;
											assign node40419 = (inp[11]) ? node40441 : node40420;
												assign node40420 = (inp[1]) ? node40428 : node40421;
													assign node40421 = (inp[7]) ? node40425 : node40422;
														assign node40422 = (inp[5]) ? 4'b0110 : 4'b0010;
														assign node40425 = (inp[5]) ? 4'b0011 : 4'b0110;
													assign node40428 = (inp[0]) ? node40434 : node40429;
														assign node40429 = (inp[5]) ? node40431 : 4'b0110;
															assign node40431 = (inp[7]) ? 4'b0010 : 4'b0110;
														assign node40434 = (inp[5]) ? node40438 : node40435;
															assign node40435 = (inp[7]) ? 4'b0110 : 4'b0010;
															assign node40438 = (inp[7]) ? 4'b0010 : 4'b0110;
												assign node40441 = (inp[1]) ? node40463 : node40442;
													assign node40442 = (inp[9]) ? node40450 : node40443;
														assign node40443 = (inp[7]) ? node40447 : node40444;
															assign node40444 = (inp[5]) ? 4'b0111 : 4'b0011;
															assign node40447 = (inp[5]) ? 4'b0011 : 4'b0111;
														assign node40450 = (inp[0]) ? node40456 : node40451;
															assign node40451 = (inp[5]) ? 4'b0111 : node40452;
																assign node40452 = (inp[7]) ? 4'b0111 : 4'b0011;
															assign node40456 = (inp[7]) ? node40460 : node40457;
																assign node40457 = (inp[5]) ? 4'b0111 : 4'b0011;
																assign node40460 = (inp[5]) ? 4'b0011 : 4'b0111;
													assign node40463 = (inp[5]) ? node40467 : node40464;
														assign node40464 = (inp[7]) ? 4'b0110 : 4'b0010;
														assign node40467 = (inp[7]) ? 4'b0011 : 4'b0110;
											assign node40470 = (inp[11]) ? node40480 : node40471;
												assign node40471 = (inp[5]) ? node40475 : node40472;
													assign node40472 = (inp[7]) ? 4'b0111 : 4'b0011;
													assign node40475 = (inp[7]) ? node40477 : 4'b0111;
														assign node40477 = (inp[1]) ? 4'b0011 : 4'b0010;
												assign node40480 = (inp[1]) ? node40488 : node40481;
													assign node40481 = (inp[5]) ? node40485 : node40482;
														assign node40482 = (inp[7]) ? 4'b0110 : 4'b0010;
														assign node40485 = (inp[7]) ? 4'b0010 : 4'b0110;
													assign node40488 = (inp[5]) ? node40492 : node40489;
														assign node40489 = (inp[7]) ? 4'b0111 : 4'b0011;
														assign node40492 = (inp[7]) ? 4'b0010 : 4'b0111;
										assign node40495 = (inp[13]) ? node40537 : node40496;
											assign node40496 = (inp[1]) ? node40528 : node40497;
												assign node40497 = (inp[11]) ? node40505 : node40498;
													assign node40498 = (inp[7]) ? node40502 : node40499;
														assign node40499 = (inp[5]) ? 4'b0111 : 4'b0011;
														assign node40502 = (inp[5]) ? 4'b0010 : 4'b0111;
													assign node40505 = (inp[9]) ? node40515 : node40506;
														assign node40506 = (inp[0]) ? node40508 : 4'b0010;
															assign node40508 = (inp[7]) ? node40512 : node40509;
																assign node40509 = (inp[5]) ? 4'b0110 : 4'b0010;
																assign node40512 = (inp[5]) ? 4'b0010 : 4'b0110;
														assign node40515 = (inp[0]) ? node40523 : node40516;
															assign node40516 = (inp[7]) ? node40520 : node40517;
																assign node40517 = (inp[5]) ? 4'b0110 : 4'b0010;
																assign node40520 = (inp[5]) ? 4'b0010 : 4'b0110;
															assign node40523 = (inp[5]) ? node40525 : 4'b0110;
																assign node40525 = (inp[7]) ? 4'b0010 : 4'b0110;
												assign node40528 = (inp[7]) ? node40532 : node40529;
													assign node40529 = (inp[5]) ? 4'b0111 : 4'b0011;
													assign node40532 = (inp[5]) ? node40534 : 4'b0111;
														assign node40534 = (inp[11]) ? 4'b0010 : 4'b0011;
											assign node40537 = (inp[11]) ? node40547 : node40538;
												assign node40538 = (inp[5]) ? node40542 : node40539;
													assign node40539 = (inp[7]) ? 4'b0110 : 4'b0010;
													assign node40542 = (inp[7]) ? node40544 : 4'b0110;
														assign node40544 = (inp[1]) ? 4'b0010 : 4'b0011;
												assign node40547 = (inp[1]) ? node40555 : node40548;
													assign node40548 = (inp[7]) ? node40552 : node40549;
														assign node40549 = (inp[5]) ? 4'b0111 : 4'b0011;
														assign node40552 = (inp[5]) ? 4'b0011 : 4'b0111;
													assign node40555 = (inp[5]) ? node40559 : node40556;
														assign node40556 = (inp[7]) ? 4'b0110 : 4'b0010;
														assign node40559 = (inp[7]) ? 4'b0011 : 4'b0110;
									assign node40562 = (inp[11]) ? node40648 : node40563;
										assign node40563 = (inp[0]) ? node40571 : node40564;
											assign node40564 = (inp[10]) ? node40568 : node40565;
												assign node40565 = (inp[1]) ? 4'b0011 : 4'b0010;
												assign node40568 = (inp[1]) ? 4'b0010 : 4'b0011;
											assign node40571 = (inp[13]) ? node40611 : node40572;
												assign node40572 = (inp[9]) ? node40594 : node40573;
													assign node40573 = (inp[5]) ? node40587 : node40574;
														assign node40574 = (inp[7]) ? node40582 : node40575;
															assign node40575 = (inp[10]) ? node40579 : node40576;
																assign node40576 = (inp[1]) ? 4'b0011 : 4'b0010;
																assign node40579 = (inp[1]) ? 4'b0010 : 4'b0011;
															assign node40582 = (inp[1]) ? 4'b0011 : node40583;
																assign node40583 = (inp[10]) ? 4'b0011 : 4'b0010;
														assign node40587 = (inp[1]) ? node40591 : node40588;
															assign node40588 = (inp[10]) ? 4'b0011 : 4'b0010;
															assign node40591 = (inp[10]) ? 4'b0010 : 4'b0011;
													assign node40594 = (inp[5]) ? node40604 : node40595;
														assign node40595 = (inp[7]) ? node40597 : 4'b0010;
															assign node40597 = (inp[10]) ? node40601 : node40598;
																assign node40598 = (inp[1]) ? 4'b0011 : 4'b0010;
																assign node40601 = (inp[1]) ? 4'b0010 : 4'b0011;
														assign node40604 = (inp[1]) ? node40608 : node40605;
															assign node40605 = (inp[10]) ? 4'b0011 : 4'b0010;
															assign node40608 = (inp[10]) ? 4'b0010 : 4'b0011;
												assign node40611 = (inp[5]) ? node40635 : node40612;
													assign node40612 = (inp[9]) ? node40628 : node40613;
														assign node40613 = (inp[7]) ? node40621 : node40614;
															assign node40614 = (inp[10]) ? node40618 : node40615;
																assign node40615 = (inp[1]) ? 4'b0011 : 4'b0010;
																assign node40618 = (inp[1]) ? 4'b0010 : 4'b0011;
															assign node40621 = (inp[10]) ? node40625 : node40622;
																assign node40622 = (inp[1]) ? 4'b0011 : 4'b0010;
																assign node40625 = (inp[1]) ? 4'b0010 : 4'b0011;
														assign node40628 = (inp[1]) ? node40632 : node40629;
															assign node40629 = (inp[10]) ? 4'b0011 : 4'b0010;
															assign node40632 = (inp[10]) ? 4'b0010 : 4'b0011;
													assign node40635 = (inp[7]) ? node40643 : node40636;
														assign node40636 = (inp[1]) ? node40640 : node40637;
															assign node40637 = (inp[10]) ? 4'b0011 : 4'b0010;
															assign node40640 = (inp[10]) ? 4'b0010 : 4'b0011;
														assign node40643 = (inp[10]) ? node40645 : 4'b0010;
															assign node40645 = (inp[1]) ? 4'b0010 : 4'b0011;
										assign node40648 = (inp[13]) ? node40718 : node40649;
											assign node40649 = (inp[5]) ? node40695 : node40650;
												assign node40650 = (inp[9]) ? node40664 : node40651;
													assign node40651 = (inp[1]) ? node40657 : node40652;
														assign node40652 = (inp[7]) ? node40654 : 4'b0010;
															assign node40654 = (inp[10]) ? 4'b0011 : 4'b0010;
														assign node40657 = (inp[10]) ? node40661 : node40658;
															assign node40658 = (inp[7]) ? 4'b0011 : 4'b0010;
															assign node40661 = (inp[7]) ? 4'b0010 : 4'b0011;
													assign node40664 = (inp[0]) ? node40680 : node40665;
														assign node40665 = (inp[7]) ? node40673 : node40666;
															assign node40666 = (inp[1]) ? node40670 : node40667;
																assign node40667 = (inp[10]) ? 4'b0010 : 4'b0011;
																assign node40670 = (inp[10]) ? 4'b0011 : 4'b0010;
															assign node40673 = (inp[1]) ? node40677 : node40674;
																assign node40674 = (inp[10]) ? 4'b0011 : 4'b0010;
																assign node40677 = (inp[10]) ? 4'b0010 : 4'b0011;
														assign node40680 = (inp[10]) ? node40688 : node40681;
															assign node40681 = (inp[7]) ? node40685 : node40682;
																assign node40682 = (inp[1]) ? 4'b0010 : 4'b0011;
																assign node40685 = (inp[1]) ? 4'b0011 : 4'b0010;
															assign node40688 = (inp[1]) ? node40692 : node40689;
																assign node40689 = (inp[7]) ? 4'b0011 : 4'b0010;
																assign node40692 = (inp[7]) ? 4'b0010 : 4'b0011;
												assign node40695 = (inp[7]) ? node40711 : node40696;
													assign node40696 = (inp[0]) ? node40704 : node40697;
														assign node40697 = (inp[1]) ? node40701 : node40698;
															assign node40698 = (inp[10]) ? 4'b0011 : 4'b0010;
															assign node40701 = (inp[10]) ? 4'b0010 : 4'b0011;
														assign node40704 = (inp[9]) ? 4'b0011 : node40705;
															assign node40705 = (inp[1]) ? 4'b0011 : node40706;
																assign node40706 = (inp[10]) ? 4'b0011 : 4'b0010;
													assign node40711 = (inp[1]) ? node40715 : node40712;
														assign node40712 = (inp[10]) ? 4'b0010 : 4'b0011;
														assign node40715 = (inp[10]) ? 4'b0011 : 4'b0010;
											assign node40718 = (inp[5]) ? node40760 : node40719;
												assign node40719 = (inp[9]) ? node40735 : node40720;
													assign node40720 = (inp[10]) ? node40728 : node40721;
														assign node40721 = (inp[0]) ? 4'b0011 : node40722;
															assign node40722 = (inp[1]) ? 4'b0011 : node40723;
																assign node40723 = (inp[7]) ? 4'b0010 : 4'b0011;
														assign node40728 = (inp[7]) ? node40732 : node40729;
															assign node40729 = (inp[1]) ? 4'b0011 : 4'b0010;
															assign node40732 = (inp[1]) ? 4'b0010 : 4'b0011;
													assign node40735 = (inp[7]) ? node40749 : node40736;
														assign node40736 = (inp[0]) ? node40742 : node40737;
															assign node40737 = (inp[10]) ? node40739 : 4'b0010;
																assign node40739 = (inp[1]) ? 4'b0011 : 4'b0010;
															assign node40742 = (inp[1]) ? node40746 : node40743;
																assign node40743 = (inp[10]) ? 4'b0010 : 4'b0011;
																assign node40746 = (inp[10]) ? 4'b0011 : 4'b0010;
														assign node40749 = (inp[0]) ? node40755 : node40750;
															assign node40750 = (inp[1]) ? node40752 : 4'b0011;
																assign node40752 = (inp[10]) ? 4'b0010 : 4'b0011;
															assign node40755 = (inp[10]) ? 4'b0011 : node40756;
																assign node40756 = (inp[1]) ? 4'b0011 : 4'b0010;
												assign node40760 = (inp[9]) ? node40776 : node40761;
													assign node40761 = (inp[10]) ? node40769 : node40762;
														assign node40762 = (inp[7]) ? node40766 : node40763;
															assign node40763 = (inp[1]) ? 4'b0011 : 4'b0010;
															assign node40766 = (inp[1]) ? 4'b0010 : 4'b0011;
														assign node40769 = (inp[7]) ? node40773 : node40770;
															assign node40770 = (inp[1]) ? 4'b0010 : 4'b0011;
															assign node40773 = (inp[1]) ? 4'b0011 : 4'b0010;
													assign node40776 = (inp[10]) ? node40784 : node40777;
														assign node40777 = (inp[7]) ? node40781 : node40778;
															assign node40778 = (inp[1]) ? 4'b0011 : 4'b0010;
															assign node40781 = (inp[1]) ? 4'b0010 : 4'b0011;
														assign node40784 = (inp[7]) ? node40788 : node40785;
															assign node40785 = (inp[1]) ? 4'b0010 : 4'b0011;
															assign node40788 = (inp[1]) ? 4'b0011 : 4'b0010;
								assign node40791 = (inp[15]) ? node41075 : node40792;
									assign node40792 = (inp[9]) ? node40970 : node40793;
										assign node40793 = (inp[1]) ? node40877 : node40794;
											assign node40794 = (inp[5]) ? node40830 : node40795;
												assign node40795 = (inp[7]) ? node40815 : node40796;
													assign node40796 = (inp[11]) ? node40802 : node40797;
														assign node40797 = (inp[10]) ? node40799 : 4'b0110;
															assign node40799 = (inp[13]) ? 4'b0110 : 4'b0111;
														assign node40802 = (inp[0]) ? node40808 : node40803;
															assign node40803 = (inp[10]) ? 4'b0110 : node40804;
																assign node40804 = (inp[13]) ? 4'b0111 : 4'b0110;
															assign node40808 = (inp[10]) ? node40812 : node40809;
																assign node40809 = (inp[13]) ? 4'b0111 : 4'b0110;
																assign node40812 = (inp[13]) ? 4'b0110 : 4'b0111;
													assign node40815 = (inp[13]) ? node40823 : node40816;
														assign node40816 = (inp[11]) ? node40820 : node40817;
															assign node40817 = (inp[10]) ? 4'b0010 : 4'b0011;
															assign node40820 = (inp[10]) ? 4'b0011 : 4'b0010;
														assign node40823 = (inp[11]) ? node40827 : node40824;
															assign node40824 = (inp[10]) ? 4'b0011 : 4'b0010;
															assign node40827 = (inp[10]) ? 4'b0010 : 4'b0011;
												assign node40830 = (inp[7]) ? node40854 : node40831;
													assign node40831 = (inp[11]) ? node40839 : node40832;
														assign node40832 = (inp[13]) ? node40836 : node40833;
															assign node40833 = (inp[10]) ? 4'b0010 : 4'b0011;
															assign node40836 = (inp[10]) ? 4'b0011 : 4'b0010;
														assign node40839 = (inp[0]) ? node40847 : node40840;
															assign node40840 = (inp[10]) ? node40844 : node40841;
																assign node40841 = (inp[13]) ? 4'b0011 : 4'b0010;
																assign node40844 = (inp[13]) ? 4'b0010 : 4'b0011;
															assign node40847 = (inp[10]) ? node40851 : node40848;
																assign node40848 = (inp[13]) ? 4'b0011 : 4'b0010;
																assign node40851 = (inp[13]) ? 4'b0010 : 4'b0011;
													assign node40854 = (inp[10]) ? node40862 : node40855;
														assign node40855 = (inp[13]) ? node40859 : node40856;
															assign node40856 = (inp[11]) ? 4'b0111 : 4'b0110;
															assign node40859 = (inp[11]) ? 4'b0110 : 4'b0111;
														assign node40862 = (inp[0]) ? node40870 : node40863;
															assign node40863 = (inp[11]) ? node40867 : node40864;
																assign node40864 = (inp[13]) ? 4'b0110 : 4'b0111;
																assign node40867 = (inp[13]) ? 4'b0111 : 4'b0110;
															assign node40870 = (inp[11]) ? node40874 : node40871;
																assign node40871 = (inp[13]) ? 4'b0110 : 4'b0111;
																assign node40874 = (inp[13]) ? 4'b0111 : 4'b0110;
											assign node40877 = (inp[11]) ? node40909 : node40878;
												assign node40878 = (inp[13]) ? node40894 : node40879;
													assign node40879 = (inp[10]) ? node40887 : node40880;
														assign node40880 = (inp[7]) ? node40884 : node40881;
															assign node40881 = (inp[5]) ? 4'b0011 : 4'b0111;
															assign node40884 = (inp[5]) ? 4'b0110 : 4'b0011;
														assign node40887 = (inp[5]) ? node40891 : node40888;
															assign node40888 = (inp[7]) ? 4'b0010 : 4'b0110;
															assign node40891 = (inp[7]) ? 4'b0111 : 4'b0010;
													assign node40894 = (inp[10]) ? node40902 : node40895;
														assign node40895 = (inp[5]) ? node40899 : node40896;
															assign node40896 = (inp[7]) ? 4'b0010 : 4'b0110;
															assign node40899 = (inp[7]) ? 4'b0111 : 4'b0010;
														assign node40902 = (inp[5]) ? node40906 : node40903;
															assign node40903 = (inp[7]) ? 4'b0011 : 4'b0111;
															assign node40906 = (inp[7]) ? 4'b0110 : 4'b0011;
												assign node40909 = (inp[13]) ? node40941 : node40910;
													assign node40910 = (inp[0]) ? node40926 : node40911;
														assign node40911 = (inp[10]) ? node40919 : node40912;
															assign node40912 = (inp[5]) ? node40916 : node40913;
																assign node40913 = (inp[7]) ? 4'b0011 : 4'b0110;
																assign node40916 = (inp[7]) ? 4'b0110 : 4'b0011;
															assign node40919 = (inp[7]) ? node40923 : node40920;
																assign node40920 = (inp[5]) ? 4'b0010 : 4'b0111;
																assign node40923 = (inp[5]) ? 4'b0111 : 4'b0010;
														assign node40926 = (inp[5]) ? node40934 : node40927;
															assign node40927 = (inp[7]) ? node40931 : node40928;
																assign node40928 = (inp[10]) ? 4'b0111 : 4'b0110;
																assign node40931 = (inp[10]) ? 4'b0010 : 4'b0011;
															assign node40934 = (inp[7]) ? node40938 : node40935;
																assign node40935 = (inp[10]) ? 4'b0010 : 4'b0011;
																assign node40938 = (inp[10]) ? 4'b0111 : 4'b0110;
													assign node40941 = (inp[0]) ? node40957 : node40942;
														assign node40942 = (inp[5]) ? node40950 : node40943;
															assign node40943 = (inp[7]) ? node40947 : node40944;
																assign node40944 = (inp[10]) ? 4'b0110 : 4'b0111;
																assign node40947 = (inp[10]) ? 4'b0011 : 4'b0010;
															assign node40950 = (inp[7]) ? node40954 : node40951;
																assign node40951 = (inp[10]) ? 4'b0011 : 4'b0010;
																assign node40954 = (inp[10]) ? 4'b0110 : 4'b0111;
														assign node40957 = (inp[10]) ? node40965 : node40958;
															assign node40958 = (inp[5]) ? node40962 : node40959;
																assign node40959 = (inp[7]) ? 4'b0010 : 4'b0111;
																assign node40962 = (inp[7]) ? 4'b0111 : 4'b0010;
															assign node40965 = (inp[7]) ? node40967 : 4'b0011;
																assign node40967 = (inp[5]) ? 4'b0110 : 4'b0011;
										assign node40970 = (inp[5]) ? node41028 : node40971;
											assign node40971 = (inp[7]) ? node41001 : node40972;
												assign node40972 = (inp[1]) ? node40980 : node40973;
													assign node40973 = (inp[13]) ? node40977 : node40974;
														assign node40974 = (inp[10]) ? 4'b0111 : 4'b0110;
														assign node40977 = (inp[10]) ? 4'b0110 : 4'b0111;
													assign node40980 = (inp[0]) ? node40990 : node40981;
														assign node40981 = (inp[11]) ? node40983 : 4'b0110;
															assign node40983 = (inp[13]) ? node40987 : node40984;
																assign node40984 = (inp[10]) ? 4'b0111 : 4'b0110;
																assign node40987 = (inp[10]) ? 4'b0110 : 4'b0111;
														assign node40990 = (inp[11]) ? node40996 : node40991;
															assign node40991 = (inp[10]) ? 4'b0111 : node40992;
																assign node40992 = (inp[13]) ? 4'b0110 : 4'b0111;
															assign node40996 = (inp[10]) ? 4'b0110 : node40997;
																assign node40997 = (inp[13]) ? 4'b0111 : 4'b0110;
												assign node41001 = (inp[1]) ? node41021 : node41002;
													assign node41002 = (inp[0]) ? node41016 : node41003;
														assign node41003 = (inp[10]) ? node41011 : node41004;
															assign node41004 = (inp[13]) ? node41008 : node41005;
																assign node41005 = (inp[11]) ? 4'b0010 : 4'b0011;
																assign node41008 = (inp[11]) ? 4'b0011 : 4'b0010;
															assign node41011 = (inp[13]) ? 4'b0011 : node41012;
																assign node41012 = (inp[11]) ? 4'b0011 : 4'b0010;
														assign node41016 = (inp[11]) ? node41018 : 4'b0011;
															assign node41018 = (inp[13]) ? 4'b0010 : 4'b0011;
													assign node41021 = (inp[10]) ? node41025 : node41022;
														assign node41022 = (inp[13]) ? 4'b0010 : 4'b0011;
														assign node41025 = (inp[13]) ? 4'b0011 : 4'b0010;
											assign node41028 = (inp[7]) ? node41050 : node41029;
												assign node41029 = (inp[11]) ? node41037 : node41030;
													assign node41030 = (inp[13]) ? node41034 : node41031;
														assign node41031 = (inp[10]) ? 4'b0010 : 4'b0011;
														assign node41034 = (inp[10]) ? 4'b0011 : 4'b0010;
													assign node41037 = (inp[1]) ? node41045 : node41038;
														assign node41038 = (inp[13]) ? node41042 : node41039;
															assign node41039 = (inp[10]) ? 4'b0011 : 4'b0010;
															assign node41042 = (inp[10]) ? 4'b0010 : 4'b0011;
														assign node41045 = (inp[10]) ? 4'b0011 : node41046;
															assign node41046 = (inp[13]) ? 4'b0010 : 4'b0011;
												assign node41050 = (inp[11]) ? node41058 : node41051;
													assign node41051 = (inp[13]) ? node41055 : node41052;
														assign node41052 = (inp[10]) ? 4'b0111 : 4'b0110;
														assign node41055 = (inp[10]) ? 4'b0110 : 4'b0111;
													assign node41058 = (inp[0]) ? node41066 : node41059;
														assign node41059 = (inp[10]) ? node41061 : 4'b0111;
															assign node41061 = (inp[13]) ? 4'b0111 : node41062;
																assign node41062 = (inp[1]) ? 4'b0111 : 4'b0110;
														assign node41066 = (inp[13]) ? node41068 : 4'b0111;
															assign node41068 = (inp[1]) ? node41072 : node41069;
																assign node41069 = (inp[10]) ? 4'b0111 : 4'b0110;
																assign node41072 = (inp[10]) ? 4'b0110 : 4'b0111;
									assign node41075 = (inp[9]) ? node41115 : node41076;
										assign node41076 = (inp[10]) ? node41096 : node41077;
											assign node41077 = (inp[1]) ? node41087 : node41078;
												assign node41078 = (inp[11]) ? 4'b0110 : node41079;
													assign node41079 = (inp[5]) ? node41083 : node41080;
														assign node41080 = (inp[7]) ? 4'b0111 : 4'b0110;
														assign node41083 = (inp[7]) ? 4'b0110 : 4'b0111;
												assign node41087 = (inp[11]) ? 4'b0111 : node41088;
													assign node41088 = (inp[5]) ? node41092 : node41089;
														assign node41089 = (inp[7]) ? 4'b0110 : 4'b0111;
														assign node41092 = (inp[7]) ? 4'b0111 : 4'b0110;
											assign node41096 = (inp[1]) ? node41106 : node41097;
												assign node41097 = (inp[11]) ? 4'b0111 : node41098;
													assign node41098 = (inp[7]) ? node41102 : node41099;
														assign node41099 = (inp[5]) ? 4'b0110 : 4'b0111;
														assign node41102 = (inp[5]) ? 4'b0111 : 4'b0110;
												assign node41106 = (inp[11]) ? 4'b0110 : node41107;
													assign node41107 = (inp[7]) ? node41111 : node41108;
														assign node41108 = (inp[5]) ? 4'b0111 : 4'b0110;
														assign node41111 = (inp[5]) ? 4'b0110 : 4'b0111;
										assign node41115 = (inp[13]) ? node41155 : node41116;
											assign node41116 = (inp[10]) ? node41136 : node41117;
												assign node41117 = (inp[1]) ? node41127 : node41118;
													assign node41118 = (inp[11]) ? 4'b0110 : node41119;
														assign node41119 = (inp[7]) ? node41123 : node41120;
															assign node41120 = (inp[5]) ? 4'b0111 : 4'b0110;
															assign node41123 = (inp[5]) ? 4'b0110 : 4'b0111;
													assign node41127 = (inp[11]) ? 4'b0111 : node41128;
														assign node41128 = (inp[5]) ? node41132 : node41129;
															assign node41129 = (inp[7]) ? 4'b0110 : 4'b0111;
															assign node41132 = (inp[7]) ? 4'b0111 : 4'b0110;
												assign node41136 = (inp[1]) ? node41146 : node41137;
													assign node41137 = (inp[11]) ? 4'b0111 : node41138;
														assign node41138 = (inp[7]) ? node41142 : node41139;
															assign node41139 = (inp[5]) ? 4'b0110 : 4'b0111;
															assign node41142 = (inp[5]) ? 4'b0111 : 4'b0110;
													assign node41146 = (inp[11]) ? 4'b0110 : node41147;
														assign node41147 = (inp[7]) ? node41151 : node41148;
															assign node41148 = (inp[5]) ? 4'b0111 : 4'b0110;
															assign node41151 = (inp[5]) ? 4'b0110 : 4'b0111;
											assign node41155 = (inp[1]) ? node41191 : node41156;
												assign node41156 = (inp[10]) ? node41174 : node41157;
													assign node41157 = (inp[11]) ? 4'b0110 : node41158;
														assign node41158 = (inp[0]) ? node41166 : node41159;
															assign node41159 = (inp[5]) ? node41163 : node41160;
																assign node41160 = (inp[7]) ? 4'b0111 : 4'b0110;
																assign node41163 = (inp[7]) ? 4'b0110 : 4'b0111;
															assign node41166 = (inp[5]) ? node41170 : node41167;
																assign node41167 = (inp[7]) ? 4'b0111 : 4'b0110;
																assign node41170 = (inp[7]) ? 4'b0110 : 4'b0111;
													assign node41174 = (inp[11]) ? 4'b0111 : node41175;
														assign node41175 = (inp[0]) ? node41183 : node41176;
															assign node41176 = (inp[5]) ? node41180 : node41177;
																assign node41177 = (inp[7]) ? 4'b0110 : 4'b0111;
																assign node41180 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node41183 = (inp[5]) ? node41187 : node41184;
																assign node41184 = (inp[7]) ? 4'b0110 : 4'b0111;
																assign node41187 = (inp[7]) ? 4'b0111 : 4'b0110;
												assign node41191 = (inp[10]) ? node41201 : node41192;
													assign node41192 = (inp[11]) ? 4'b0111 : node41193;
														assign node41193 = (inp[7]) ? node41197 : node41194;
															assign node41194 = (inp[5]) ? 4'b0110 : 4'b0111;
															assign node41197 = (inp[5]) ? 4'b0111 : 4'b0110;
													assign node41201 = (inp[11]) ? 4'b0110 : node41202;
														assign node41202 = (inp[0]) ? node41208 : node41203;
															assign node41203 = (inp[5]) ? node41205 : 4'b0111;
																assign node41205 = (inp[7]) ? 4'b0110 : 4'b0111;
															assign node41208 = (inp[7]) ? node41212 : node41209;
																assign node41209 = (inp[5]) ? 4'b0111 : 4'b0110;
																assign node41212 = (inp[5]) ? 4'b0110 : 4'b0111;
							assign node41216 = (inp[2]) ? node41516 : node41217;
								assign node41217 = (inp[15]) ? node41429 : node41218;
									assign node41218 = (inp[7]) ? node41386 : node41219;
										assign node41219 = (inp[9]) ? node41307 : node41220;
											assign node41220 = (inp[11]) ? node41258 : node41221;
												assign node41221 = (inp[5]) ? node41233 : node41222;
													assign node41222 = (inp[1]) ? node41228 : node41223;
														assign node41223 = (inp[13]) ? node41225 : 4'b0010;
															assign node41225 = (inp[10]) ? 4'b0010 : 4'b0011;
														assign node41228 = (inp[10]) ? node41230 : 4'b0010;
															assign node41230 = (inp[13]) ? 4'b0010 : 4'b0011;
													assign node41233 = (inp[1]) ? node41249 : node41234;
														assign node41234 = (inp[0]) ? node41242 : node41235;
															assign node41235 = (inp[13]) ? node41239 : node41236;
																assign node41236 = (inp[10]) ? 4'b0010 : 4'b0011;
																assign node41239 = (inp[10]) ? 4'b0011 : 4'b0010;
															assign node41242 = (inp[13]) ? node41246 : node41243;
																assign node41243 = (inp[10]) ? 4'b0010 : 4'b0011;
																assign node41246 = (inp[10]) ? 4'b0011 : 4'b0010;
														assign node41249 = (inp[0]) ? node41253 : node41250;
															assign node41250 = (inp[10]) ? 4'b0010 : 4'b0011;
															assign node41253 = (inp[13]) ? node41255 : 4'b0010;
																assign node41255 = (inp[10]) ? 4'b0011 : 4'b0010;
												assign node41258 = (inp[13]) ? node41288 : node41259;
													assign node41259 = (inp[5]) ? node41273 : node41260;
														assign node41260 = (inp[0]) ? node41266 : node41261;
															assign node41261 = (inp[10]) ? node41263 : 4'b0011;
																assign node41263 = (inp[1]) ? 4'b0011 : 4'b0010;
															assign node41266 = (inp[1]) ? node41270 : node41267;
																assign node41267 = (inp[10]) ? 4'b0010 : 4'b0011;
																assign node41270 = (inp[10]) ? 4'b0011 : 4'b0010;
														assign node41273 = (inp[0]) ? node41281 : node41274;
															assign node41274 = (inp[10]) ? node41278 : node41275;
																assign node41275 = (inp[1]) ? 4'b0011 : 4'b0010;
																assign node41278 = (inp[1]) ? 4'b0010 : 4'b0011;
															assign node41281 = (inp[1]) ? node41285 : node41282;
																assign node41282 = (inp[10]) ? 4'b0011 : 4'b0010;
																assign node41285 = (inp[10]) ? 4'b0010 : 4'b0011;
													assign node41288 = (inp[1]) ? node41302 : node41289;
														assign node41289 = (inp[0]) ? node41295 : node41290;
															assign node41290 = (inp[5]) ? node41292 : 4'b0011;
																assign node41292 = (inp[10]) ? 4'b0010 : 4'b0011;
															assign node41295 = (inp[5]) ? node41299 : node41296;
																assign node41296 = (inp[10]) ? 4'b0011 : 4'b0010;
																assign node41299 = (inp[10]) ? 4'b0010 : 4'b0011;
														assign node41302 = (inp[10]) ? node41304 : 4'b0010;
															assign node41304 = (inp[5]) ? 4'b0011 : 4'b0010;
											assign node41307 = (inp[11]) ? node41357 : node41308;
												assign node41308 = (inp[1]) ? node41332 : node41309;
													assign node41309 = (inp[10]) ? node41325 : node41310;
														assign node41310 = (inp[0]) ? node41318 : node41311;
															assign node41311 = (inp[5]) ? node41315 : node41312;
																assign node41312 = (inp[13]) ? 4'b0011 : 4'b0010;
																assign node41315 = (inp[13]) ? 4'b0010 : 4'b0011;
															assign node41318 = (inp[5]) ? node41322 : node41319;
																assign node41319 = (inp[13]) ? 4'b0011 : 4'b0010;
																assign node41322 = (inp[13]) ? 4'b0010 : 4'b0011;
														assign node41325 = (inp[13]) ? node41329 : node41326;
															assign node41326 = (inp[5]) ? 4'b0010 : 4'b0011;
															assign node41329 = (inp[5]) ? 4'b0011 : 4'b0010;
													assign node41332 = (inp[5]) ? node41342 : node41333;
														assign node41333 = (inp[0]) ? 4'b0011 : node41334;
															assign node41334 = (inp[10]) ? node41338 : node41335;
																assign node41335 = (inp[13]) ? 4'b0011 : 4'b0010;
																assign node41338 = (inp[13]) ? 4'b0010 : 4'b0011;
														assign node41342 = (inp[0]) ? node41350 : node41343;
															assign node41343 = (inp[10]) ? node41347 : node41344;
																assign node41344 = (inp[13]) ? 4'b0010 : 4'b0011;
																assign node41347 = (inp[13]) ? 4'b0011 : 4'b0010;
															assign node41350 = (inp[10]) ? node41354 : node41351;
																assign node41351 = (inp[13]) ? 4'b0010 : 4'b0011;
																assign node41354 = (inp[13]) ? 4'b0011 : 4'b0010;
												assign node41357 = (inp[10]) ? node41371 : node41358;
													assign node41358 = (inp[13]) ? node41364 : node41359;
														assign node41359 = (inp[1]) ? node41361 : 4'b0010;
															assign node41361 = (inp[5]) ? 4'b0011 : 4'b0010;
														assign node41364 = (inp[1]) ? node41368 : node41365;
															assign node41365 = (inp[5]) ? 4'b0011 : 4'b0010;
															assign node41368 = (inp[5]) ? 4'b0010 : 4'b0011;
													assign node41371 = (inp[13]) ? node41379 : node41372;
														assign node41372 = (inp[1]) ? node41376 : node41373;
															assign node41373 = (inp[5]) ? 4'b0011 : 4'b0010;
															assign node41376 = (inp[5]) ? 4'b0010 : 4'b0011;
														assign node41379 = (inp[5]) ? node41383 : node41380;
															assign node41380 = (inp[1]) ? 4'b0010 : 4'b0011;
															assign node41383 = (inp[1]) ? 4'b0011 : 4'b0010;
										assign node41386 = (inp[11]) ? node41394 : node41387;
											assign node41387 = (inp[10]) ? node41391 : node41388;
												assign node41388 = (inp[13]) ? 4'b0111 : 4'b0110;
												assign node41391 = (inp[13]) ? 4'b0110 : 4'b0111;
											assign node41394 = (inp[1]) ? node41422 : node41395;
												assign node41395 = (inp[0]) ? node41403 : node41396;
													assign node41396 = (inp[13]) ? node41400 : node41397;
														assign node41397 = (inp[10]) ? 4'b0110 : 4'b0111;
														assign node41400 = (inp[10]) ? 4'b0111 : 4'b0110;
													assign node41403 = (inp[9]) ? node41409 : node41404;
														assign node41404 = (inp[10]) ? 4'b0110 : node41405;
															assign node41405 = (inp[13]) ? 4'b0110 : 4'b0111;
														assign node41409 = (inp[5]) ? node41417 : node41410;
															assign node41410 = (inp[10]) ? node41414 : node41411;
																assign node41411 = (inp[13]) ? 4'b0110 : 4'b0111;
																assign node41414 = (inp[13]) ? 4'b0111 : 4'b0110;
															assign node41417 = (inp[13]) ? 4'b0111 : node41418;
																assign node41418 = (inp[10]) ? 4'b0110 : 4'b0111;
												assign node41422 = (inp[13]) ? node41426 : node41423;
													assign node41423 = (inp[10]) ? 4'b0111 : 4'b0110;
													assign node41426 = (inp[10]) ? 4'b0110 : 4'b0111;
									assign node41429 = (inp[10]) ? node41473 : node41430;
										assign node41430 = (inp[1]) ? node41440 : node41431;
											assign node41431 = (inp[7]) ? 4'b0110 : node41432;
												assign node41432 = (inp[11]) ? node41436 : node41433;
													assign node41433 = (inp[5]) ? 4'b0111 : 4'b0110;
													assign node41436 = (inp[5]) ? 4'b0110 : 4'b0111;
											assign node41440 = (inp[7]) ? 4'b0111 : node41441;
												assign node41441 = (inp[0]) ? node41465 : node41442;
													assign node41442 = (inp[13]) ? node41458 : node41443;
														assign node41443 = (inp[9]) ? node41451 : node41444;
															assign node41444 = (inp[5]) ? node41448 : node41445;
																assign node41445 = (inp[11]) ? 4'b0110 : 4'b0111;
																assign node41448 = (inp[11]) ? 4'b0111 : 4'b0110;
															assign node41451 = (inp[11]) ? node41455 : node41452;
																assign node41452 = (inp[5]) ? 4'b0110 : 4'b0111;
																assign node41455 = (inp[5]) ? 4'b0111 : 4'b0110;
														assign node41458 = (inp[5]) ? node41462 : node41459;
															assign node41459 = (inp[11]) ? 4'b0110 : 4'b0111;
															assign node41462 = (inp[11]) ? 4'b0111 : 4'b0110;
													assign node41465 = (inp[11]) ? node41469 : node41466;
														assign node41466 = (inp[5]) ? 4'b0110 : 4'b0111;
														assign node41469 = (inp[5]) ? 4'b0111 : 4'b0110;
										assign node41473 = (inp[1]) ? node41507 : node41474;
											assign node41474 = (inp[7]) ? 4'b0111 : node41475;
												assign node41475 = (inp[0]) ? node41491 : node41476;
													assign node41476 = (inp[13]) ? node41484 : node41477;
														assign node41477 = (inp[5]) ? node41481 : node41478;
															assign node41478 = (inp[11]) ? 4'b0110 : 4'b0111;
															assign node41481 = (inp[11]) ? 4'b0111 : 4'b0110;
														assign node41484 = (inp[11]) ? node41488 : node41485;
															assign node41485 = (inp[5]) ? 4'b0110 : 4'b0111;
															assign node41488 = (inp[5]) ? 4'b0111 : 4'b0110;
													assign node41491 = (inp[13]) ? node41499 : node41492;
														assign node41492 = (inp[11]) ? node41496 : node41493;
															assign node41493 = (inp[5]) ? 4'b0110 : 4'b0111;
															assign node41496 = (inp[5]) ? 4'b0111 : 4'b0110;
														assign node41499 = (inp[5]) ? node41503 : node41500;
															assign node41500 = (inp[11]) ? 4'b0110 : 4'b0111;
															assign node41503 = (inp[11]) ? 4'b0111 : 4'b0110;
											assign node41507 = (inp[7]) ? 4'b0110 : node41508;
												assign node41508 = (inp[5]) ? node41512 : node41509;
													assign node41509 = (inp[11]) ? 4'b0111 : 4'b0110;
													assign node41512 = (inp[11]) ? 4'b0110 : 4'b0111;
								assign node41516 = (inp[7]) ? node41710 : node41517;
									assign node41517 = (inp[15]) ? node41589 : node41518;
										assign node41518 = (inp[5]) ? node41566 : node41519;
											assign node41519 = (inp[0]) ? node41543 : node41520;
												assign node41520 = (inp[11]) ? node41536 : node41521;
													assign node41521 = (inp[13]) ? node41529 : node41522;
														assign node41522 = (inp[10]) ? node41526 : node41523;
															assign node41523 = (inp[1]) ? 4'b0110 : 4'b0111;
															assign node41526 = (inp[1]) ? 4'b0111 : 4'b0110;
														assign node41529 = (inp[1]) ? node41533 : node41530;
															assign node41530 = (inp[10]) ? 4'b0111 : 4'b0110;
															assign node41533 = (inp[10]) ? 4'b0110 : 4'b0111;
													assign node41536 = (inp[10]) ? node41540 : node41537;
														assign node41537 = (inp[13]) ? 4'b0110 : 4'b0111;
														assign node41540 = (inp[13]) ? 4'b0111 : 4'b0110;
												assign node41543 = (inp[13]) ? node41555 : node41544;
													assign node41544 = (inp[10]) ? node41550 : node41545;
														assign node41545 = (inp[1]) ? node41547 : 4'b0111;
															assign node41547 = (inp[11]) ? 4'b0111 : 4'b0110;
														assign node41550 = (inp[11]) ? 4'b0110 : node41551;
															assign node41551 = (inp[1]) ? 4'b0111 : 4'b0110;
													assign node41555 = (inp[10]) ? node41561 : node41556;
														assign node41556 = (inp[11]) ? 4'b0110 : node41557;
															assign node41557 = (inp[1]) ? 4'b0111 : 4'b0110;
														assign node41561 = (inp[11]) ? 4'b0111 : node41562;
															assign node41562 = (inp[1]) ? 4'b0110 : 4'b0111;
											assign node41566 = (inp[10]) ? node41578 : node41567;
												assign node41567 = (inp[13]) ? node41573 : node41568;
													assign node41568 = (inp[11]) ? 4'b0110 : node41569;
														assign node41569 = (inp[1]) ? 4'b0111 : 4'b0110;
													assign node41573 = (inp[11]) ? 4'b0111 : node41574;
														assign node41574 = (inp[1]) ? 4'b0110 : 4'b0111;
												assign node41578 = (inp[13]) ? node41584 : node41579;
													assign node41579 = (inp[1]) ? node41581 : 4'b0111;
														assign node41581 = (inp[11]) ? 4'b0111 : 4'b0110;
													assign node41584 = (inp[1]) ? node41586 : 4'b0110;
														assign node41586 = (inp[11]) ? 4'b0110 : 4'b0111;
										assign node41589 = (inp[10]) ? node41635 : node41590;
											assign node41590 = (inp[1]) ? node41628 : node41591;
												assign node41591 = (inp[13]) ? node41615 : node41592;
													assign node41592 = (inp[9]) ? node41608 : node41593;
														assign node41593 = (inp[0]) ? node41601 : node41594;
															assign node41594 = (inp[11]) ? node41598 : node41595;
																assign node41595 = (inp[5]) ? 4'b0011 : 4'b0010;
																assign node41598 = (inp[5]) ? 4'b0010 : 4'b0011;
															assign node41601 = (inp[5]) ? node41605 : node41602;
																assign node41602 = (inp[11]) ? 4'b0011 : 4'b0010;
																assign node41605 = (inp[11]) ? 4'b0010 : 4'b0011;
														assign node41608 = (inp[11]) ? node41612 : node41609;
															assign node41609 = (inp[5]) ? 4'b0011 : 4'b0010;
															assign node41612 = (inp[5]) ? 4'b0010 : 4'b0011;
													assign node41615 = (inp[9]) ? node41621 : node41616;
														assign node41616 = (inp[11]) ? 4'b0010 : node41617;
															assign node41617 = (inp[5]) ? 4'b0011 : 4'b0010;
														assign node41621 = (inp[11]) ? node41625 : node41622;
															assign node41622 = (inp[5]) ? 4'b0011 : 4'b0010;
															assign node41625 = (inp[5]) ? 4'b0010 : 4'b0011;
												assign node41628 = (inp[5]) ? node41632 : node41629;
													assign node41629 = (inp[11]) ? 4'b0010 : 4'b0011;
													assign node41632 = (inp[11]) ? 4'b0011 : 4'b0010;
											assign node41635 = (inp[0]) ? node41667 : node41636;
												assign node41636 = (inp[5]) ? node41652 : node41637;
													assign node41637 = (inp[13]) ? node41645 : node41638;
														assign node41638 = (inp[1]) ? node41642 : node41639;
															assign node41639 = (inp[11]) ? 4'b0010 : 4'b0011;
															assign node41642 = (inp[11]) ? 4'b0011 : 4'b0010;
														assign node41645 = (inp[11]) ? node41649 : node41646;
															assign node41646 = (inp[1]) ? 4'b0010 : 4'b0011;
															assign node41649 = (inp[1]) ? 4'b0011 : 4'b0010;
													assign node41652 = (inp[9]) ? node41660 : node41653;
														assign node41653 = (inp[1]) ? node41657 : node41654;
															assign node41654 = (inp[11]) ? 4'b0011 : 4'b0010;
															assign node41657 = (inp[11]) ? 4'b0010 : 4'b0011;
														assign node41660 = (inp[1]) ? node41664 : node41661;
															assign node41661 = (inp[11]) ? 4'b0011 : 4'b0010;
															assign node41664 = (inp[11]) ? 4'b0010 : 4'b0011;
												assign node41667 = (inp[9]) ? node41689 : node41668;
													assign node41668 = (inp[13]) ? node41684 : node41669;
														assign node41669 = (inp[11]) ? node41677 : node41670;
															assign node41670 = (inp[5]) ? node41674 : node41671;
																assign node41671 = (inp[1]) ? 4'b0010 : 4'b0011;
																assign node41674 = (inp[1]) ? 4'b0011 : 4'b0010;
															assign node41677 = (inp[1]) ? node41681 : node41678;
																assign node41678 = (inp[5]) ? 4'b0011 : 4'b0010;
																assign node41681 = (inp[5]) ? 4'b0010 : 4'b0011;
														assign node41684 = (inp[1]) ? 4'b0010 : node41685;
															assign node41685 = (inp[11]) ? 4'b0011 : 4'b0010;
													assign node41689 = (inp[11]) ? node41697 : node41690;
														assign node41690 = (inp[5]) ? node41694 : node41691;
															assign node41691 = (inp[1]) ? 4'b0010 : 4'b0011;
															assign node41694 = (inp[1]) ? 4'b0011 : 4'b0010;
														assign node41697 = (inp[13]) ? node41703 : node41698;
															assign node41698 = (inp[5]) ? 4'b0010 : node41699;
																assign node41699 = (inp[1]) ? 4'b0011 : 4'b0010;
															assign node41703 = (inp[5]) ? node41707 : node41704;
																assign node41704 = (inp[1]) ? 4'b0011 : 4'b0010;
																assign node41707 = (inp[1]) ? 4'b0010 : 4'b0011;
									assign node41710 = (inp[15]) ? node41768 : node41711;
										assign node41711 = (inp[1]) ? node41761 : node41712;
											assign node41712 = (inp[5]) ? node41746 : node41713;
												assign node41713 = (inp[10]) ? node41721 : node41714;
													assign node41714 = (inp[11]) ? node41718 : node41715;
														assign node41715 = (inp[13]) ? 4'b0011 : 4'b0010;
														assign node41718 = (inp[13]) ? 4'b0010 : 4'b0011;
													assign node41721 = (inp[9]) ? node41731 : node41722;
														assign node41722 = (inp[0]) ? node41724 : 4'b0010;
															assign node41724 = (inp[11]) ? node41728 : node41725;
																assign node41725 = (inp[13]) ? 4'b0010 : 4'b0011;
																assign node41728 = (inp[13]) ? 4'b0011 : 4'b0010;
														assign node41731 = (inp[0]) ? node41739 : node41732;
															assign node41732 = (inp[11]) ? node41736 : node41733;
																assign node41733 = (inp[13]) ? 4'b0010 : 4'b0011;
																assign node41736 = (inp[13]) ? 4'b0011 : 4'b0010;
															assign node41739 = (inp[13]) ? node41743 : node41740;
																assign node41740 = (inp[11]) ? 4'b0010 : 4'b0011;
																assign node41743 = (inp[11]) ? 4'b0011 : 4'b0010;
												assign node41746 = (inp[13]) ? node41754 : node41747;
													assign node41747 = (inp[11]) ? node41751 : node41748;
														assign node41748 = (inp[10]) ? 4'b0011 : 4'b0010;
														assign node41751 = (inp[10]) ? 4'b0010 : 4'b0011;
													assign node41754 = (inp[10]) ? node41758 : node41755;
														assign node41755 = (inp[11]) ? 4'b0010 : 4'b0011;
														assign node41758 = (inp[11]) ? 4'b0011 : 4'b0010;
											assign node41761 = (inp[10]) ? node41765 : node41762;
												assign node41762 = (inp[13]) ? 4'b0011 : 4'b0010;
												assign node41765 = (inp[13]) ? 4'b0010 : 4'b0011;
										assign node41768 = (inp[9]) ? node41814 : node41769;
											assign node41769 = (inp[5]) ? node41793 : node41770;
												assign node41770 = (inp[11]) ? node41778 : node41771;
													assign node41771 = (inp[1]) ? node41775 : node41772;
														assign node41772 = (inp[10]) ? 4'b0011 : 4'b0010;
														assign node41775 = (inp[10]) ? 4'b0010 : 4'b0011;
													assign node41778 = (inp[13]) ? node41786 : node41779;
														assign node41779 = (inp[10]) ? node41783 : node41780;
															assign node41780 = (inp[1]) ? 4'b0011 : 4'b0010;
															assign node41783 = (inp[1]) ? 4'b0010 : 4'b0011;
														assign node41786 = (inp[10]) ? node41790 : node41787;
															assign node41787 = (inp[1]) ? 4'b0011 : 4'b0010;
															assign node41790 = (inp[1]) ? 4'b0010 : 4'b0011;
												assign node41793 = (inp[11]) ? node41807 : node41794;
													assign node41794 = (inp[13]) ? node41802 : node41795;
														assign node41795 = (inp[1]) ? node41799 : node41796;
															assign node41796 = (inp[10]) ? 4'b0011 : 4'b0010;
															assign node41799 = (inp[10]) ? 4'b0010 : 4'b0011;
														assign node41802 = (inp[10]) ? 4'b0011 : node41803;
															assign node41803 = (inp[1]) ? 4'b0011 : 4'b0010;
													assign node41807 = (inp[1]) ? node41811 : node41808;
														assign node41808 = (inp[10]) ? 4'b0011 : 4'b0010;
														assign node41811 = (inp[10]) ? 4'b0010 : 4'b0011;
											assign node41814 = (inp[10]) ? node41818 : node41815;
												assign node41815 = (inp[1]) ? 4'b0011 : 4'b0010;
												assign node41818 = (inp[1]) ? 4'b0010 : 4'b0011;
					assign node41821 = (inp[8]) ? node44523 : node41822;
						assign node41822 = (inp[7]) ? node43208 : node41823;
							assign node41823 = (inp[4]) ? node42481 : node41824;
								assign node41824 = (inp[15]) ? node42176 : node41825;
									assign node41825 = (inp[5]) ? node42009 : node41826;
										assign node41826 = (inp[1]) ? node41928 : node41827;
											assign node41827 = (inp[2]) ? node41881 : node41828;
												assign node41828 = (inp[13]) ? node41850 : node41829;
													assign node41829 = (inp[11]) ? node41843 : node41830;
														assign node41830 = (inp[10]) ? node41836 : node41831;
															assign node41831 = (inp[9]) ? 4'b0101 : node41832;
																assign node41832 = (inp[0]) ? 4'b0101 : 4'b0100;
															assign node41836 = (inp[0]) ? node41840 : node41837;
																assign node41837 = (inp[9]) ? 4'b0100 : 4'b0101;
																assign node41840 = (inp[9]) ? 4'b0101 : 4'b0100;
														assign node41843 = (inp[10]) ? node41847 : node41844;
															assign node41844 = (inp[9]) ? 4'b0100 : 4'b0101;
															assign node41847 = (inp[9]) ? 4'b0101 : 4'b0100;
													assign node41850 = (inp[0]) ? node41866 : node41851;
														assign node41851 = (inp[9]) ? node41859 : node41852;
															assign node41852 = (inp[10]) ? node41856 : node41853;
																assign node41853 = (inp[11]) ? 4'b0000 : 4'b0001;
																assign node41856 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node41859 = (inp[11]) ? node41863 : node41860;
																assign node41860 = (inp[10]) ? 4'b0001 : 4'b0000;
																assign node41863 = (inp[10]) ? 4'b0000 : 4'b0001;
														assign node41866 = (inp[11]) ? node41874 : node41867;
															assign node41867 = (inp[9]) ? node41871 : node41868;
																assign node41868 = (inp[10]) ? 4'b0001 : 4'b0000;
																assign node41871 = (inp[10]) ? 4'b0000 : 4'b0001;
															assign node41874 = (inp[9]) ? node41878 : node41875;
																assign node41875 = (inp[10]) ? 4'b0001 : 4'b0000;
																assign node41878 = (inp[10]) ? 4'b0000 : 4'b0001;
												assign node41881 = (inp[13]) ? node41907 : node41882;
													assign node41882 = (inp[11]) ? node41892 : node41883;
														assign node41883 = (inp[0]) ? node41885 : 4'b0001;
															assign node41885 = (inp[9]) ? node41889 : node41886;
																assign node41886 = (inp[10]) ? 4'b0001 : 4'b0000;
																assign node41889 = (inp[10]) ? 4'b0000 : 4'b0001;
														assign node41892 = (inp[0]) ? node41900 : node41893;
															assign node41893 = (inp[9]) ? node41897 : node41894;
																assign node41894 = (inp[10]) ? 4'b0001 : 4'b0000;
																assign node41897 = (inp[10]) ? 4'b0000 : 4'b0001;
															assign node41900 = (inp[10]) ? node41904 : node41901;
																assign node41901 = (inp[9]) ? 4'b0001 : 4'b0000;
																assign node41904 = (inp[9]) ? 4'b0000 : 4'b0001;
													assign node41907 = (inp[9]) ? node41919 : node41908;
														assign node41908 = (inp[10]) ? node41914 : node41909;
															assign node41909 = (inp[11]) ? node41911 : 4'b0101;
																assign node41911 = (inp[0]) ? 4'b0100 : 4'b0101;
															assign node41914 = (inp[0]) ? node41916 : 4'b0100;
																assign node41916 = (inp[11]) ? 4'b0101 : 4'b0100;
														assign node41919 = (inp[10]) ? node41923 : node41920;
															assign node41920 = (inp[11]) ? 4'b0101 : 4'b0100;
															assign node41923 = (inp[11]) ? node41925 : 4'b0101;
																assign node41925 = (inp[0]) ? 4'b0100 : 4'b0101;
											assign node41928 = (inp[13]) ? node41968 : node41929;
												assign node41929 = (inp[2]) ? node41947 : node41930;
													assign node41930 = (inp[10]) ? node41940 : node41931;
														assign node41931 = (inp[9]) ? node41935 : node41932;
															assign node41932 = (inp[0]) ? 4'b0000 : 4'b0001;
															assign node41935 = (inp[11]) ? node41937 : 4'b0000;
																assign node41937 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node41940 = (inp[9]) ? 4'b0001 : node41941;
															assign node41941 = (inp[11]) ? node41943 : 4'b0000;
																assign node41943 = (inp[0]) ? 4'b0001 : 4'b0000;
													assign node41947 = (inp[0]) ? node41961 : node41948;
														assign node41948 = (inp[9]) ? node41956 : node41949;
															assign node41949 = (inp[10]) ? node41953 : node41950;
																assign node41950 = (inp[11]) ? 4'b0101 : 4'b0100;
																assign node41953 = (inp[11]) ? 4'b0100 : 4'b0101;
															assign node41956 = (inp[10]) ? 4'b0100 : node41957;
																assign node41957 = (inp[11]) ? 4'b0100 : 4'b0101;
														assign node41961 = (inp[10]) ? node41965 : node41962;
															assign node41962 = (inp[9]) ? 4'b0100 : 4'b0101;
															assign node41965 = (inp[9]) ? 4'b0101 : 4'b0100;
												assign node41968 = (inp[2]) ? node41992 : node41969;
													assign node41969 = (inp[9]) ? node41981 : node41970;
														assign node41970 = (inp[10]) ? node41976 : node41971;
															assign node41971 = (inp[0]) ? 4'b0101 : node41972;
																assign node41972 = (inp[11]) ? 4'b0101 : 4'b0100;
															assign node41976 = (inp[11]) ? 4'b0100 : node41977;
																assign node41977 = (inp[0]) ? 4'b0100 : 4'b0101;
														assign node41981 = (inp[10]) ? node41987 : node41982;
															assign node41982 = (inp[0]) ? 4'b0100 : node41983;
																assign node41983 = (inp[11]) ? 4'b0100 : 4'b0101;
															assign node41987 = (inp[0]) ? 4'b0101 : node41988;
																assign node41988 = (inp[11]) ? 4'b0101 : 4'b0100;
													assign node41992 = (inp[11]) ? node42004 : node41993;
														assign node41993 = (inp[9]) ? node41999 : node41994;
															assign node41994 = (inp[10]) ? node41996 : 4'b0000;
																assign node41996 = (inp[0]) ? 4'b0001 : 4'b0000;
															assign node41999 = (inp[10]) ? 4'b0001 : node42000;
																assign node42000 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node42004 = (inp[10]) ? 4'b0001 : node42005;
															assign node42005 = (inp[9]) ? 4'b0001 : 4'b0000;
										assign node42009 = (inp[0]) ? node42085 : node42010;
											assign node42010 = (inp[13]) ? node42048 : node42011;
												assign node42011 = (inp[2]) ? node42027 : node42012;
													assign node42012 = (inp[9]) ? node42022 : node42013;
														assign node42013 = (inp[10]) ? node42019 : node42014;
															assign node42014 = (inp[11]) ? node42016 : 4'b0000;
																assign node42016 = (inp[1]) ? 4'b0001 : 4'b0000;
															assign node42019 = (inp[1]) ? 4'b0000 : 4'b0001;
														assign node42022 = (inp[10]) ? 4'b0000 : node42023;
															assign node42023 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node42027 = (inp[10]) ? node42039 : node42028;
														assign node42028 = (inp[9]) ? node42034 : node42029;
															assign node42029 = (inp[1]) ? 4'b0100 : node42030;
																assign node42030 = (inp[11]) ? 4'b0100 : 4'b0101;
															assign node42034 = (inp[11]) ? 4'b0101 : node42035;
																assign node42035 = (inp[1]) ? 4'b0101 : 4'b0100;
														assign node42039 = (inp[9]) ? node42043 : node42040;
															assign node42040 = (inp[1]) ? 4'b0101 : 4'b0100;
															assign node42043 = (inp[1]) ? 4'b0100 : node42044;
																assign node42044 = (inp[11]) ? 4'b0100 : 4'b0101;
												assign node42048 = (inp[2]) ? node42062 : node42049;
													assign node42049 = (inp[10]) ? node42057 : node42050;
														assign node42050 = (inp[9]) ? node42054 : node42051;
															assign node42051 = (inp[11]) ? 4'b0100 : 4'b0101;
															assign node42054 = (inp[11]) ? 4'b0101 : 4'b0100;
														assign node42057 = (inp[9]) ? 4'b0100 : node42058;
															assign node42058 = (inp[1]) ? 4'b0101 : 4'b0100;
													assign node42062 = (inp[10]) ? node42074 : node42063;
														assign node42063 = (inp[9]) ? node42069 : node42064;
															assign node42064 = (inp[11]) ? 4'b0001 : node42065;
																assign node42065 = (inp[1]) ? 4'b0001 : 4'b0000;
															assign node42069 = (inp[1]) ? 4'b0000 : node42070;
																assign node42070 = (inp[11]) ? 4'b0000 : 4'b0001;
														assign node42074 = (inp[9]) ? node42080 : node42075;
															assign node42075 = (inp[11]) ? 4'b0000 : node42076;
																assign node42076 = (inp[1]) ? 4'b0000 : 4'b0001;
															assign node42080 = (inp[11]) ? 4'b0001 : node42081;
																assign node42081 = (inp[1]) ? 4'b0001 : 4'b0000;
											assign node42085 = (inp[1]) ? node42125 : node42086;
												assign node42086 = (inp[9]) ? node42106 : node42087;
													assign node42087 = (inp[10]) ? node42097 : node42088;
														assign node42088 = (inp[13]) ? node42094 : node42089;
															assign node42089 = (inp[2]) ? 4'b0100 : node42090;
																assign node42090 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node42094 = (inp[2]) ? 4'b0001 : 4'b0100;
														assign node42097 = (inp[2]) ? node42103 : node42098;
															assign node42098 = (inp[13]) ? 4'b0101 : node42099;
																assign node42099 = (inp[11]) ? 4'b0000 : 4'b0001;
															assign node42103 = (inp[13]) ? 4'b0000 : 4'b0101;
													assign node42106 = (inp[10]) ? node42116 : node42107;
														assign node42107 = (inp[2]) ? node42113 : node42108;
															assign node42108 = (inp[13]) ? 4'b0101 : node42109;
																assign node42109 = (inp[11]) ? 4'b0000 : 4'b0001;
															assign node42113 = (inp[13]) ? 4'b0000 : 4'b0101;
														assign node42116 = (inp[2]) ? node42122 : node42117;
															assign node42117 = (inp[13]) ? 4'b0100 : node42118;
																assign node42118 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node42122 = (inp[13]) ? 4'b0001 : 4'b0100;
												assign node42125 = (inp[2]) ? node42149 : node42126;
													assign node42126 = (inp[13]) ? node42134 : node42127;
														assign node42127 = (inp[10]) ? node42131 : node42128;
															assign node42128 = (inp[9]) ? 4'b0000 : 4'b0001;
															assign node42131 = (inp[9]) ? 4'b0001 : 4'b0000;
														assign node42134 = (inp[11]) ? node42142 : node42135;
															assign node42135 = (inp[10]) ? node42139 : node42136;
																assign node42136 = (inp[9]) ? 4'b0101 : 4'b0100;
																assign node42139 = (inp[9]) ? 4'b0100 : 4'b0101;
															assign node42142 = (inp[9]) ? node42146 : node42143;
																assign node42143 = (inp[10]) ? 4'b0100 : 4'b0101;
																assign node42146 = (inp[10]) ? 4'b0101 : 4'b0100;
													assign node42149 = (inp[13]) ? node42163 : node42150;
														assign node42150 = (inp[9]) ? node42158 : node42151;
															assign node42151 = (inp[10]) ? node42155 : node42152;
																assign node42152 = (inp[11]) ? 4'b0101 : 4'b0100;
																assign node42155 = (inp[11]) ? 4'b0100 : 4'b0101;
															assign node42158 = (inp[10]) ? 4'b0100 : node42159;
																assign node42159 = (inp[11]) ? 4'b0100 : 4'b0101;
														assign node42163 = (inp[11]) ? node42171 : node42164;
															assign node42164 = (inp[10]) ? node42168 : node42165;
																assign node42165 = (inp[9]) ? 4'b0000 : 4'b0001;
																assign node42168 = (inp[9]) ? 4'b0001 : 4'b0000;
															assign node42171 = (inp[9]) ? 4'b0000 : node42172;
																assign node42172 = (inp[10]) ? 4'b0001 : 4'b0000;
									assign node42176 = (inp[2]) ? node42318 : node42177;
										assign node42177 = (inp[13]) ? node42257 : node42178;
											assign node42178 = (inp[1]) ? node42214 : node42179;
												assign node42179 = (inp[5]) ? node42201 : node42180;
													assign node42180 = (inp[9]) ? node42192 : node42181;
														assign node42181 = (inp[10]) ? node42187 : node42182;
															assign node42182 = (inp[0]) ? 4'b0111 : node42183;
																assign node42183 = (inp[11]) ? 4'b0111 : 4'b0110;
															assign node42187 = (inp[0]) ? 4'b0110 : node42188;
																assign node42188 = (inp[11]) ? 4'b0110 : 4'b0111;
														assign node42192 = (inp[10]) ? node42196 : node42193;
															assign node42193 = (inp[0]) ? 4'b0110 : 4'b0111;
															assign node42196 = (inp[11]) ? 4'b0111 : node42197;
																assign node42197 = (inp[0]) ? 4'b0111 : 4'b0110;
													assign node42201 = (inp[9]) ? node42207 : node42202;
														assign node42202 = (inp[10]) ? 4'b0011 : node42203;
															assign node42203 = (inp[0]) ? 4'b0011 : 4'b0010;
														assign node42207 = (inp[10]) ? node42211 : node42208;
															assign node42208 = (inp[11]) ? 4'b0010 : 4'b0011;
															assign node42211 = (inp[11]) ? 4'b0011 : 4'b0010;
												assign node42214 = (inp[0]) ? node42234 : node42215;
													assign node42215 = (inp[5]) ? node42227 : node42216;
														assign node42216 = (inp[9]) ? node42222 : node42217;
															assign node42217 = (inp[11]) ? node42219 : 4'b0011;
																assign node42219 = (inp[10]) ? 4'b0010 : 4'b0011;
															assign node42222 = (inp[10]) ? node42224 : 4'b0010;
																assign node42224 = (inp[11]) ? 4'b0011 : 4'b0010;
														assign node42227 = (inp[9]) ? node42231 : node42228;
															assign node42228 = (inp[10]) ? 4'b0011 : 4'b0010;
															assign node42231 = (inp[10]) ? 4'b0010 : 4'b0011;
													assign node42234 = (inp[11]) ? node42250 : node42235;
														assign node42235 = (inp[5]) ? node42243 : node42236;
															assign node42236 = (inp[9]) ? node42240 : node42237;
																assign node42237 = (inp[10]) ? 4'b0010 : 4'b0011;
																assign node42240 = (inp[10]) ? 4'b0011 : 4'b0010;
															assign node42243 = (inp[10]) ? node42247 : node42244;
																assign node42244 = (inp[9]) ? 4'b0011 : 4'b0010;
																assign node42247 = (inp[9]) ? 4'b0010 : 4'b0011;
														assign node42250 = (inp[9]) ? node42254 : node42251;
															assign node42251 = (inp[10]) ? 4'b0010 : 4'b0011;
															assign node42254 = (inp[10]) ? 4'b0011 : 4'b0010;
											assign node42257 = (inp[5]) ? node42295 : node42258;
												assign node42258 = (inp[1]) ? node42276 : node42259;
													assign node42259 = (inp[9]) ? node42271 : node42260;
														assign node42260 = (inp[10]) ? node42266 : node42261;
															assign node42261 = (inp[11]) ? 4'b0011 : node42262;
																assign node42262 = (inp[0]) ? 4'b0011 : 4'b0010;
															assign node42266 = (inp[11]) ? 4'b0010 : node42267;
																assign node42267 = (inp[0]) ? 4'b0010 : 4'b0011;
														assign node42271 = (inp[10]) ? node42273 : 4'b0010;
															assign node42273 = (inp[11]) ? 4'b0011 : 4'b0010;
													assign node42276 = (inp[9]) ? node42288 : node42277;
														assign node42277 = (inp[10]) ? node42283 : node42278;
															assign node42278 = (inp[11]) ? node42280 : 4'b0111;
																assign node42280 = (inp[0]) ? 4'b0110 : 4'b0111;
															assign node42283 = (inp[0]) ? node42285 : 4'b0110;
																assign node42285 = (inp[11]) ? 4'b0111 : 4'b0110;
														assign node42288 = (inp[10]) ? 4'b0111 : node42289;
															assign node42289 = (inp[11]) ? node42291 : 4'b0110;
																assign node42291 = (inp[0]) ? 4'b0111 : 4'b0110;
												assign node42295 = (inp[9]) ? node42307 : node42296;
													assign node42296 = (inp[10]) ? node42302 : node42297;
														assign node42297 = (inp[0]) ? 4'b0111 : node42298;
															assign node42298 = (inp[11]) ? 4'b0111 : 4'b0110;
														assign node42302 = (inp[11]) ? 4'b0110 : node42303;
															assign node42303 = (inp[0]) ? 4'b0110 : 4'b0111;
													assign node42307 = (inp[10]) ? node42313 : node42308;
														assign node42308 = (inp[0]) ? 4'b0110 : node42309;
															assign node42309 = (inp[11]) ? 4'b0110 : 4'b0111;
														assign node42313 = (inp[11]) ? 4'b0111 : node42314;
															assign node42314 = (inp[0]) ? 4'b0111 : 4'b0110;
										assign node42318 = (inp[13]) ? node42408 : node42319;
											assign node42319 = (inp[1]) ? node42361 : node42320;
												assign node42320 = (inp[5]) ? node42342 : node42321;
													assign node42321 = (inp[0]) ? node42335 : node42322;
														assign node42322 = (inp[9]) ? node42328 : node42323;
															assign node42323 = (inp[10]) ? 4'b0010 : node42324;
																assign node42324 = (inp[11]) ? 4'b0010 : 4'b0011;
															assign node42328 = (inp[11]) ? node42332 : node42329;
																assign node42329 = (inp[10]) ? 4'b0011 : 4'b0010;
																assign node42332 = (inp[10]) ? 4'b0010 : 4'b0011;
														assign node42335 = (inp[10]) ? node42339 : node42336;
															assign node42336 = (inp[9]) ? 4'b0011 : 4'b0010;
															assign node42339 = (inp[9]) ? 4'b0010 : 4'b0011;
													assign node42342 = (inp[9]) ? node42352 : node42343;
														assign node42343 = (inp[10]) ? node42347 : node42344;
															assign node42344 = (inp[11]) ? 4'b0110 : 4'b0111;
															assign node42347 = (inp[11]) ? 4'b0111 : node42348;
																assign node42348 = (inp[0]) ? 4'b0111 : 4'b0110;
														assign node42352 = (inp[10]) ? node42356 : node42353;
															assign node42353 = (inp[11]) ? 4'b0111 : 4'b0110;
															assign node42356 = (inp[0]) ? 4'b0110 : node42357;
																assign node42357 = (inp[11]) ? 4'b0110 : 4'b0111;
												assign node42361 = (inp[10]) ? node42385 : node42362;
													assign node42362 = (inp[9]) ? node42374 : node42363;
														assign node42363 = (inp[5]) ? node42369 : node42364;
															assign node42364 = (inp[0]) ? node42366 : 4'b0110;
																assign node42366 = (inp[11]) ? 4'b0111 : 4'b0110;
															assign node42369 = (inp[0]) ? 4'b0110 : node42370;
																assign node42370 = (inp[11]) ? 4'b0110 : 4'b0111;
														assign node42374 = (inp[0]) ? node42380 : node42375;
															assign node42375 = (inp[11]) ? 4'b0111 : node42376;
																assign node42376 = (inp[5]) ? 4'b0110 : 4'b0111;
															assign node42380 = (inp[11]) ? node42382 : 4'b0111;
																assign node42382 = (inp[5]) ? 4'b0111 : 4'b0110;
													assign node42385 = (inp[9]) ? node42397 : node42386;
														assign node42386 = (inp[0]) ? node42392 : node42387;
															assign node42387 = (inp[5]) ? node42389 : 4'b0111;
																assign node42389 = (inp[11]) ? 4'b0111 : 4'b0110;
															assign node42392 = (inp[5]) ? 4'b0111 : node42393;
																assign node42393 = (inp[11]) ? 4'b0110 : 4'b0111;
														assign node42397 = (inp[5]) ? node42403 : node42398;
															assign node42398 = (inp[11]) ? node42400 : 4'b0110;
																assign node42400 = (inp[0]) ? 4'b0111 : 4'b0110;
															assign node42403 = (inp[11]) ? 4'b0110 : node42404;
																assign node42404 = (inp[0]) ? 4'b0110 : 4'b0111;
											assign node42408 = (inp[5]) ? node42458 : node42409;
												assign node42409 = (inp[1]) ? node42431 : node42410;
													assign node42410 = (inp[0]) ? node42416 : node42411;
														assign node42411 = (inp[9]) ? 4'b0111 : node42412;
															assign node42412 = (inp[10]) ? 4'b0111 : 4'b0110;
														assign node42416 = (inp[11]) ? node42424 : node42417;
															assign node42417 = (inp[9]) ? node42421 : node42418;
																assign node42418 = (inp[10]) ? 4'b0111 : 4'b0110;
																assign node42421 = (inp[10]) ? 4'b0110 : 4'b0111;
															assign node42424 = (inp[9]) ? node42428 : node42425;
																assign node42425 = (inp[10]) ? 4'b0110 : 4'b0111;
																assign node42428 = (inp[10]) ? 4'b0111 : 4'b0110;
													assign node42431 = (inp[11]) ? node42445 : node42432;
														assign node42432 = (inp[0]) ? node42440 : node42433;
															assign node42433 = (inp[10]) ? node42437 : node42434;
																assign node42434 = (inp[9]) ? 4'b0011 : 4'b0010;
																assign node42437 = (inp[9]) ? 4'b0010 : 4'b0011;
															assign node42440 = (inp[10]) ? node42442 : 4'b0010;
																assign node42442 = (inp[9]) ? 4'b0010 : 4'b0011;
														assign node42445 = (inp[10]) ? node42451 : node42446;
															assign node42446 = (inp[0]) ? node42448 : 4'b0011;
																assign node42448 = (inp[9]) ? 4'b0010 : 4'b0011;
															assign node42451 = (inp[0]) ? node42455 : node42452;
																assign node42452 = (inp[9]) ? 4'b0010 : 4'b0011;
																assign node42455 = (inp[9]) ? 4'b0011 : 4'b0010;
												assign node42458 = (inp[9]) ? node42470 : node42459;
													assign node42459 = (inp[10]) ? node42465 : node42460;
														assign node42460 = (inp[11]) ? 4'b0010 : node42461;
															assign node42461 = (inp[0]) ? 4'b0010 : 4'b0011;
														assign node42465 = (inp[0]) ? 4'b0011 : node42466;
															assign node42466 = (inp[11]) ? 4'b0011 : 4'b0010;
													assign node42470 = (inp[10]) ? node42476 : node42471;
														assign node42471 = (inp[11]) ? 4'b0011 : node42472;
															assign node42472 = (inp[0]) ? 4'b0011 : 4'b0010;
														assign node42476 = (inp[11]) ? 4'b0010 : node42477;
															assign node42477 = (inp[0]) ? 4'b0010 : 4'b0011;
								assign node42481 = (inp[5]) ? node42875 : node42482;
									assign node42482 = (inp[9]) ? node42666 : node42483;
										assign node42483 = (inp[15]) ? node42585 : node42484;
											assign node42484 = (inp[0]) ? node42532 : node42485;
												assign node42485 = (inp[13]) ? node42505 : node42486;
													assign node42486 = (inp[10]) ? node42496 : node42487;
														assign node42487 = (inp[1]) ? node42493 : node42488;
															assign node42488 = (inp[2]) ? node42490 : 4'b0010;
																assign node42490 = (inp[11]) ? 4'b0111 : 4'b0110;
															assign node42493 = (inp[2]) ? 4'b0011 : 4'b0111;
														assign node42496 = (inp[1]) ? node42502 : node42497;
															assign node42497 = (inp[2]) ? node42499 : 4'b0011;
																assign node42499 = (inp[11]) ? 4'b0110 : 4'b0111;
															assign node42502 = (inp[2]) ? 4'b0010 : 4'b0110;
													assign node42505 = (inp[10]) ? node42519 : node42506;
														assign node42506 = (inp[2]) ? node42512 : node42507;
															assign node42507 = (inp[1]) ? 4'b0010 : node42508;
																assign node42508 = (inp[11]) ? 4'b0110 : 4'b0111;
															assign node42512 = (inp[1]) ? node42516 : node42513;
																assign node42513 = (inp[11]) ? 4'b0010 : 4'b0011;
																assign node42516 = (inp[11]) ? 4'b0111 : 4'b0110;
														assign node42519 = (inp[2]) ? node42525 : node42520;
															assign node42520 = (inp[1]) ? 4'b0011 : node42521;
																assign node42521 = (inp[11]) ? 4'b0111 : 4'b0110;
															assign node42525 = (inp[1]) ? node42529 : node42526;
																assign node42526 = (inp[11]) ? 4'b0011 : 4'b0010;
																assign node42529 = (inp[11]) ? 4'b0110 : 4'b0111;
												assign node42532 = (inp[11]) ? node42558 : node42533;
													assign node42533 = (inp[13]) ? node42549 : node42534;
														assign node42534 = (inp[10]) ? node42542 : node42535;
															assign node42535 = (inp[1]) ? node42539 : node42536;
																assign node42536 = (inp[2]) ? 4'b0111 : 4'b0010;
																assign node42539 = (inp[2]) ? 4'b0011 : 4'b0111;
															assign node42542 = (inp[1]) ? node42546 : node42543;
																assign node42543 = (inp[2]) ? 4'b0110 : 4'b0011;
																assign node42546 = (inp[2]) ? 4'b0010 : 4'b0110;
														assign node42549 = (inp[10]) ? node42553 : node42550;
															assign node42550 = (inp[1]) ? 4'b0111 : 4'b0110;
															assign node42553 = (inp[1]) ? 4'b0011 : node42554;
																assign node42554 = (inp[2]) ? 4'b0011 : 4'b0111;
													assign node42558 = (inp[2]) ? node42572 : node42559;
														assign node42559 = (inp[13]) ? node42565 : node42560;
															assign node42560 = (inp[1]) ? node42562 : 4'b0011;
																assign node42562 = (inp[10]) ? 4'b0111 : 4'b0110;
															assign node42565 = (inp[1]) ? node42569 : node42566;
																assign node42566 = (inp[10]) ? 4'b0111 : 4'b0110;
																assign node42569 = (inp[10]) ? 4'b0010 : 4'b0011;
														assign node42572 = (inp[1]) ? node42578 : node42573;
															assign node42573 = (inp[13]) ? node42575 : 4'b0110;
																assign node42575 = (inp[10]) ? 4'b0011 : 4'b0010;
															assign node42578 = (inp[13]) ? node42582 : node42579;
																assign node42579 = (inp[10]) ? 4'b0011 : 4'b0010;
																assign node42582 = (inp[10]) ? 4'b0110 : 4'b0111;
											assign node42585 = (inp[2]) ? node42629 : node42586;
												assign node42586 = (inp[10]) ? node42610 : node42587;
													assign node42587 = (inp[0]) ? node42597 : node42588;
														assign node42588 = (inp[1]) ? node42592 : node42589;
															assign node42589 = (inp[13]) ? 4'b0010 : 4'b0110;
															assign node42592 = (inp[13]) ? node42594 : 4'b0010;
																assign node42594 = (inp[11]) ? 4'b0111 : 4'b0110;
														assign node42597 = (inp[11]) ? node42603 : node42598;
															assign node42598 = (inp[13]) ? 4'b0111 : node42599;
																assign node42599 = (inp[1]) ? 4'b0010 : 4'b0110;
															assign node42603 = (inp[13]) ? node42607 : node42604;
																assign node42604 = (inp[1]) ? 4'b0011 : 4'b0111;
																assign node42607 = (inp[1]) ? 4'b0111 : 4'b0011;
													assign node42610 = (inp[0]) ? node42620 : node42611;
														assign node42611 = (inp[13]) ? node42615 : node42612;
															assign node42612 = (inp[1]) ? 4'b0011 : 4'b0111;
															assign node42615 = (inp[1]) ? node42617 : 4'b0011;
																assign node42617 = (inp[11]) ? 4'b0110 : 4'b0111;
														assign node42620 = (inp[1]) ? 4'b0110 : node42621;
															assign node42621 = (inp[11]) ? node42625 : node42622;
																assign node42622 = (inp[13]) ? 4'b0011 : 4'b0111;
																assign node42625 = (inp[13]) ? 4'b0010 : 4'b0110;
												assign node42629 = (inp[10]) ? node42645 : node42630;
													assign node42630 = (inp[0]) ? node42638 : node42631;
														assign node42631 = (inp[11]) ? node42633 : 4'b0110;
															assign node42633 = (inp[1]) ? 4'b0111 : node42634;
																assign node42634 = (inp[13]) ? 4'b0111 : 4'b0010;
														assign node42638 = (inp[1]) ? node42642 : node42639;
															assign node42639 = (inp[13]) ? 4'b0111 : 4'b0011;
															assign node42642 = (inp[13]) ? 4'b0011 : 4'b0111;
													assign node42645 = (inp[0]) ? node42659 : node42646;
														assign node42646 = (inp[11]) ? node42654 : node42647;
															assign node42647 = (inp[13]) ? node42651 : node42648;
																assign node42648 = (inp[1]) ? 4'b0111 : 4'b0011;
																assign node42651 = (inp[1]) ? 4'b0011 : 4'b0111;
															assign node42654 = (inp[13]) ? node42656 : 4'b0011;
																assign node42656 = (inp[1]) ? 4'b0010 : 4'b0110;
														assign node42659 = (inp[1]) ? node42663 : node42660;
															assign node42660 = (inp[13]) ? 4'b0110 : 4'b0010;
															assign node42663 = (inp[13]) ? 4'b0010 : 4'b0110;
										assign node42666 = (inp[11]) ? node42762 : node42667;
											assign node42667 = (inp[10]) ? node42717 : node42668;
												assign node42668 = (inp[15]) ? node42694 : node42669;
													assign node42669 = (inp[1]) ? node42685 : node42670;
														assign node42670 = (inp[0]) ? node42678 : node42671;
															assign node42671 = (inp[13]) ? node42675 : node42672;
																assign node42672 = (inp[2]) ? 4'b0111 : 4'b0011;
																assign node42675 = (inp[2]) ? 4'b0010 : 4'b0110;
															assign node42678 = (inp[2]) ? node42682 : node42679;
																assign node42679 = (inp[13]) ? 4'b0111 : 4'b0011;
																assign node42682 = (inp[13]) ? 4'b0011 : 4'b0110;
														assign node42685 = (inp[13]) ? node42689 : node42686;
															assign node42686 = (inp[2]) ? 4'b0010 : 4'b0110;
															assign node42689 = (inp[2]) ? node42691 : 4'b0011;
																assign node42691 = (inp[0]) ? 4'b0110 : 4'b0111;
													assign node42694 = (inp[13]) ? node42708 : node42695;
														assign node42695 = (inp[0]) ? node42703 : node42696;
															assign node42696 = (inp[2]) ? node42700 : node42697;
																assign node42697 = (inp[1]) ? 4'b0011 : 4'b0111;
																assign node42700 = (inp[1]) ? 4'b0111 : 4'b0011;
															assign node42703 = (inp[2]) ? 4'b0011 : node42704;
																assign node42704 = (inp[1]) ? 4'b0011 : 4'b0111;
														assign node42708 = (inp[2]) ? node42710 : 4'b0011;
															assign node42710 = (inp[1]) ? node42714 : node42711;
																assign node42711 = (inp[0]) ? 4'b0110 : 4'b0111;
																assign node42714 = (inp[0]) ? 4'b0010 : 4'b0011;
												assign node42717 = (inp[15]) ? node42739 : node42718;
													assign node42718 = (inp[1]) ? node42730 : node42719;
														assign node42719 = (inp[13]) ? node42725 : node42720;
															assign node42720 = (inp[2]) ? node42722 : 4'b0010;
																assign node42722 = (inp[0]) ? 4'b0111 : 4'b0110;
															assign node42725 = (inp[2]) ? node42727 : 4'b0111;
																assign node42727 = (inp[0]) ? 4'b0010 : 4'b0011;
														assign node42730 = (inp[13]) ? node42734 : node42731;
															assign node42731 = (inp[2]) ? 4'b0011 : 4'b0111;
															assign node42734 = (inp[2]) ? node42736 : 4'b0010;
																assign node42736 = (inp[0]) ? 4'b0111 : 4'b0110;
													assign node42739 = (inp[0]) ? node42749 : node42740;
														assign node42740 = (inp[1]) ? node42742 : 4'b0110;
															assign node42742 = (inp[2]) ? node42746 : node42743;
																assign node42743 = (inp[13]) ? 4'b0110 : 4'b0010;
																assign node42746 = (inp[13]) ? 4'b0010 : 4'b0110;
														assign node42749 = (inp[13]) ? node42757 : node42750;
															assign node42750 = (inp[2]) ? node42754 : node42751;
																assign node42751 = (inp[1]) ? 4'b0010 : 4'b0110;
																assign node42754 = (inp[1]) ? 4'b0111 : 4'b0010;
															assign node42757 = (inp[2]) ? 4'b0111 : node42758;
																assign node42758 = (inp[1]) ? 4'b0111 : 4'b0010;
											assign node42762 = (inp[10]) ? node42820 : node42763;
												assign node42763 = (inp[0]) ? node42791 : node42764;
													assign node42764 = (inp[1]) ? node42778 : node42765;
														assign node42765 = (inp[2]) ? node42771 : node42766;
															assign node42766 = (inp[13]) ? node42768 : 4'b0111;
																assign node42768 = (inp[15]) ? 4'b0011 : 4'b0111;
															assign node42771 = (inp[15]) ? node42775 : node42772;
																assign node42772 = (inp[13]) ? 4'b0011 : 4'b0110;
																assign node42775 = (inp[13]) ? 4'b0110 : 4'b0011;
														assign node42778 = (inp[2]) ? node42786 : node42779;
															assign node42779 = (inp[15]) ? node42783 : node42780;
																assign node42780 = (inp[13]) ? 4'b0011 : 4'b0110;
																assign node42783 = (inp[13]) ? 4'b0110 : 4'b0011;
															assign node42786 = (inp[13]) ? 4'b0010 : node42787;
																assign node42787 = (inp[15]) ? 4'b0110 : 4'b0010;
													assign node42791 = (inp[15]) ? node42807 : node42792;
														assign node42792 = (inp[13]) ? node42800 : node42793;
															assign node42793 = (inp[1]) ? node42797 : node42794;
																assign node42794 = (inp[2]) ? 4'b0110 : 4'b0010;
																assign node42797 = (inp[2]) ? 4'b0011 : 4'b0111;
															assign node42800 = (inp[1]) ? node42804 : node42801;
																assign node42801 = (inp[2]) ? 4'b0011 : 4'b0111;
																assign node42804 = (inp[2]) ? 4'b0110 : 4'b0010;
														assign node42807 = (inp[13]) ? node42815 : node42808;
															assign node42808 = (inp[1]) ? node42812 : node42809;
																assign node42809 = (inp[2]) ? 4'b0010 : 4'b0110;
																assign node42812 = (inp[2]) ? 4'b0110 : 4'b0010;
															assign node42815 = (inp[1]) ? 4'b0110 : node42816;
																assign node42816 = (inp[2]) ? 4'b0110 : 4'b0010;
												assign node42820 = (inp[0]) ? node42848 : node42821;
													assign node42821 = (inp[1]) ? node42835 : node42822;
														assign node42822 = (inp[2]) ? node42830 : node42823;
															assign node42823 = (inp[13]) ? node42827 : node42824;
																assign node42824 = (inp[15]) ? 4'b0110 : 4'b0010;
																assign node42827 = (inp[15]) ? 4'b0010 : 4'b0110;
															assign node42830 = (inp[15]) ? node42832 : 4'b0010;
																assign node42832 = (inp[13]) ? 4'b0111 : 4'b0010;
														assign node42835 = (inp[2]) ? node42843 : node42836;
															assign node42836 = (inp[13]) ? node42840 : node42837;
																assign node42837 = (inp[15]) ? 4'b0010 : 4'b0111;
																assign node42840 = (inp[15]) ? 4'b0111 : 4'b0010;
															assign node42843 = (inp[15]) ? node42845 : 4'b0011;
																assign node42845 = (inp[13]) ? 4'b0011 : 4'b0111;
													assign node42848 = (inp[15]) ? node42862 : node42849;
														assign node42849 = (inp[13]) ? node42855 : node42850;
															assign node42850 = (inp[1]) ? 4'b0010 : node42851;
																assign node42851 = (inp[2]) ? 4'b0111 : 4'b0011;
															assign node42855 = (inp[1]) ? node42859 : node42856;
																assign node42856 = (inp[2]) ? 4'b0010 : 4'b0110;
																assign node42859 = (inp[2]) ? 4'b0111 : 4'b0011;
														assign node42862 = (inp[1]) ? node42870 : node42863;
															assign node42863 = (inp[2]) ? node42867 : node42864;
																assign node42864 = (inp[13]) ? 4'b0011 : 4'b0111;
																assign node42867 = (inp[13]) ? 4'b0111 : 4'b0011;
															assign node42870 = (inp[2]) ? 4'b0011 : node42871;
																assign node42871 = (inp[13]) ? 4'b0111 : 4'b0011;
									assign node42875 = (inp[10]) ? node43029 : node42876;
										assign node42876 = (inp[9]) ? node42958 : node42877;
											assign node42877 = (inp[0]) ? node42919 : node42878;
												assign node42878 = (inp[11]) ? node42900 : node42879;
													assign node42879 = (inp[15]) ? node42895 : node42880;
														assign node42880 = (inp[1]) ? node42888 : node42881;
															assign node42881 = (inp[2]) ? node42885 : node42882;
																assign node42882 = (inp[13]) ? 4'b0010 : 4'b0111;
																assign node42885 = (inp[13]) ? 4'b0111 : 4'b0011;
															assign node42888 = (inp[13]) ? node42892 : node42889;
																assign node42889 = (inp[2]) ? 4'b0010 : 4'b0110;
																assign node42892 = (inp[2]) ? 4'b0111 : 4'b0011;
														assign node42895 = (inp[13]) ? 4'b0011 : node42896;
															assign node42896 = (inp[2]) ? 4'b0111 : 4'b0011;
													assign node42900 = (inp[2]) ? node42908 : node42901;
														assign node42901 = (inp[15]) ? node42905 : node42902;
															assign node42902 = (inp[13]) ? 4'b0011 : 4'b0110;
															assign node42905 = (inp[13]) ? 4'b0110 : 4'b0011;
														assign node42908 = (inp[1]) ? node42912 : node42909;
															assign node42909 = (inp[15]) ? 4'b0010 : 4'b0111;
															assign node42912 = (inp[13]) ? node42916 : node42913;
																assign node42913 = (inp[15]) ? 4'b0110 : 4'b0010;
																assign node42916 = (inp[15]) ? 4'b0010 : 4'b0110;
												assign node42919 = (inp[15]) ? node42943 : node42920;
													assign node42920 = (inp[1]) ? node42930 : node42921;
														assign node42921 = (inp[13]) ? node42925 : node42922;
															assign node42922 = (inp[2]) ? 4'b0010 : 4'b0110;
															assign node42925 = (inp[2]) ? node42927 : 4'b0011;
																assign node42927 = (inp[11]) ? 4'b0110 : 4'b0111;
														assign node42930 = (inp[2]) ? node42938 : node42931;
															assign node42931 = (inp[13]) ? node42935 : node42932;
																assign node42932 = (inp[11]) ? 4'b0111 : 4'b0110;
																assign node42935 = (inp[11]) ? 4'b0010 : 4'b0011;
															assign node42938 = (inp[13]) ? 4'b0110 : node42939;
																assign node42939 = (inp[11]) ? 4'b0011 : 4'b0010;
													assign node42943 = (inp[11]) ? node42951 : node42944;
														assign node42944 = (inp[13]) ? node42948 : node42945;
															assign node42945 = (inp[2]) ? 4'b0110 : 4'b0011;
															assign node42948 = (inp[2]) ? 4'b0010 : 4'b0110;
														assign node42951 = (inp[13]) ? node42955 : node42952;
															assign node42952 = (inp[2]) ? 4'b0110 : 4'b0010;
															assign node42955 = (inp[2]) ? 4'b0010 : 4'b0110;
											assign node42958 = (inp[0]) ? node43000 : node42959;
												assign node42959 = (inp[11]) ? node42985 : node42960;
													assign node42960 = (inp[15]) ? node42972 : node42961;
														assign node42961 = (inp[13]) ? node42967 : node42962;
															assign node42962 = (inp[2]) ? 4'b0011 : node42963;
																assign node42963 = (inp[1]) ? 4'b0111 : 4'b0110;
															assign node42967 = (inp[2]) ? 4'b0110 : node42968;
																assign node42968 = (inp[1]) ? 4'b0010 : 4'b0011;
														assign node42972 = (inp[1]) ? node42978 : node42973;
															assign node42973 = (inp[2]) ? 4'b0010 : node42974;
																assign node42974 = (inp[13]) ? 4'b0110 : 4'b0010;
															assign node42978 = (inp[13]) ? node42982 : node42979;
																assign node42979 = (inp[2]) ? 4'b0110 : 4'b0010;
																assign node42982 = (inp[2]) ? 4'b0010 : 4'b0110;
													assign node42985 = (inp[2]) ? node42993 : node42986;
														assign node42986 = (inp[15]) ? node42990 : node42987;
															assign node42987 = (inp[13]) ? 4'b0010 : 4'b0111;
															assign node42990 = (inp[13]) ? 4'b0111 : 4'b0010;
														assign node42993 = (inp[13]) ? node42997 : node42994;
															assign node42994 = (inp[15]) ? 4'b0111 : 4'b0011;
															assign node42997 = (inp[15]) ? 4'b0011 : 4'b0110;
												assign node43000 = (inp[15]) ? node43020 : node43001;
													assign node43001 = (inp[2]) ? node43011 : node43002;
														assign node43002 = (inp[13]) ? node43006 : node43003;
															assign node43003 = (inp[1]) ? 4'b0110 : 4'b0111;
															assign node43006 = (inp[11]) ? node43008 : 4'b0010;
																assign node43008 = (inp[1]) ? 4'b0011 : 4'b0010;
														assign node43011 = (inp[13]) ? node43017 : node43012;
															assign node43012 = (inp[11]) ? node43014 : 4'b0011;
																assign node43014 = (inp[1]) ? 4'b0010 : 4'b0011;
															assign node43017 = (inp[11]) ? 4'b0111 : 4'b0110;
													assign node43020 = (inp[13]) ? node43026 : node43021;
														assign node43021 = (inp[2]) ? 4'b0111 : node43022;
															assign node43022 = (inp[11]) ? 4'b0011 : 4'b0010;
														assign node43026 = (inp[2]) ? 4'b0011 : 4'b0111;
										assign node43029 = (inp[9]) ? node43105 : node43030;
											assign node43030 = (inp[11]) ? node43076 : node43031;
												assign node43031 = (inp[0]) ? node43053 : node43032;
													assign node43032 = (inp[15]) ? node43046 : node43033;
														assign node43033 = (inp[1]) ? node43041 : node43034;
															assign node43034 = (inp[13]) ? node43038 : node43035;
																assign node43035 = (inp[2]) ? 4'b0010 : 4'b0110;
																assign node43038 = (inp[2]) ? 4'b0110 : 4'b0011;
															assign node43041 = (inp[13]) ? 4'b0110 : node43042;
																assign node43042 = (inp[2]) ? 4'b0011 : 4'b0111;
														assign node43046 = (inp[2]) ? node43050 : node43047;
															assign node43047 = (inp[13]) ? 4'b0110 : 4'b0010;
															assign node43050 = (inp[13]) ? 4'b0010 : 4'b0110;
													assign node43053 = (inp[2]) ? node43069 : node43054;
														assign node43054 = (inp[1]) ? node43062 : node43055;
															assign node43055 = (inp[13]) ? node43059 : node43056;
																assign node43056 = (inp[15]) ? 4'b0010 : 4'b0111;
																assign node43059 = (inp[15]) ? 4'b0111 : 4'b0010;
															assign node43062 = (inp[15]) ? node43066 : node43063;
																assign node43063 = (inp[13]) ? 4'b0010 : 4'b0111;
																assign node43066 = (inp[13]) ? 4'b0111 : 4'b0010;
														assign node43069 = (inp[13]) ? node43073 : node43070;
															assign node43070 = (inp[15]) ? 4'b0111 : 4'b0011;
															assign node43073 = (inp[15]) ? 4'b0011 : 4'b0110;
												assign node43076 = (inp[2]) ? node43090 : node43077;
													assign node43077 = (inp[15]) ? node43085 : node43078;
														assign node43078 = (inp[13]) ? 4'b0010 : node43079;
															assign node43079 = (inp[1]) ? node43081 : 4'b0111;
																assign node43081 = (inp[0]) ? 4'b0110 : 4'b0111;
														assign node43085 = (inp[13]) ? 4'b0111 : node43086;
															assign node43086 = (inp[0]) ? 4'b0011 : 4'b0010;
													assign node43090 = (inp[15]) ? node43102 : node43091;
														assign node43091 = (inp[13]) ? node43097 : node43092;
															assign node43092 = (inp[1]) ? node43094 : 4'b0011;
																assign node43094 = (inp[0]) ? 4'b0010 : 4'b0011;
															assign node43097 = (inp[1]) ? 4'b0111 : node43098;
																assign node43098 = (inp[0]) ? 4'b0111 : 4'b0110;
														assign node43102 = (inp[13]) ? 4'b0011 : 4'b0111;
											assign node43105 = (inp[0]) ? node43163 : node43106;
												assign node43106 = (inp[11]) ? node43136 : node43107;
													assign node43107 = (inp[15]) ? node43121 : node43108;
														assign node43108 = (inp[1]) ? node43116 : node43109;
															assign node43109 = (inp[13]) ? node43113 : node43110;
																assign node43110 = (inp[2]) ? 4'b0011 : 4'b0111;
																assign node43113 = (inp[2]) ? 4'b0111 : 4'b0010;
															assign node43116 = (inp[13]) ? 4'b0111 : node43117;
																assign node43117 = (inp[2]) ? 4'b0010 : 4'b0110;
														assign node43121 = (inp[1]) ? node43129 : node43122;
															assign node43122 = (inp[2]) ? node43126 : node43123;
																assign node43123 = (inp[13]) ? 4'b0111 : 4'b0011;
																assign node43126 = (inp[13]) ? 4'b0011 : 4'b0111;
															assign node43129 = (inp[2]) ? node43133 : node43130;
																assign node43130 = (inp[13]) ? 4'b0111 : 4'b0011;
																assign node43133 = (inp[13]) ? 4'b0011 : 4'b0111;
													assign node43136 = (inp[2]) ? node43152 : node43137;
														assign node43137 = (inp[1]) ? node43145 : node43138;
															assign node43138 = (inp[15]) ? node43142 : node43139;
																assign node43139 = (inp[13]) ? 4'b0011 : 4'b0110;
																assign node43142 = (inp[13]) ? 4'b0110 : 4'b0011;
															assign node43145 = (inp[13]) ? node43149 : node43146;
																assign node43146 = (inp[15]) ? 4'b0011 : 4'b0110;
																assign node43149 = (inp[15]) ? 4'b0110 : 4'b0011;
														assign node43152 = (inp[1]) ? node43158 : node43153;
															assign node43153 = (inp[13]) ? 4'b0111 : node43154;
																assign node43154 = (inp[15]) ? 4'b0110 : 4'b0010;
															assign node43158 = (inp[15]) ? 4'b0010 : node43159;
																assign node43159 = (inp[13]) ? 4'b0110 : 4'b0010;
												assign node43163 = (inp[15]) ? node43187 : node43164;
													assign node43164 = (inp[1]) ? node43172 : node43165;
														assign node43165 = (inp[11]) ? 4'b0110 : node43166;
															assign node43166 = (inp[13]) ? node43168 : 4'b0110;
																assign node43168 = (inp[2]) ? 4'b0111 : 4'b0011;
														assign node43172 = (inp[11]) ? node43180 : node43173;
															assign node43173 = (inp[2]) ? node43177 : node43174;
																assign node43174 = (inp[13]) ? 4'b0011 : 4'b0110;
																assign node43177 = (inp[13]) ? 4'b0110 : 4'b0010;
															assign node43180 = (inp[13]) ? node43184 : node43181;
																assign node43181 = (inp[2]) ? 4'b0011 : 4'b0111;
																assign node43184 = (inp[2]) ? 4'b0110 : 4'b0010;
													assign node43187 = (inp[11]) ? node43193 : node43188;
														assign node43188 = (inp[2]) ? node43190 : 4'b0110;
															assign node43190 = (inp[13]) ? 4'b0010 : 4'b0110;
														assign node43193 = (inp[1]) ? node43201 : node43194;
															assign node43194 = (inp[13]) ? node43198 : node43195;
																assign node43195 = (inp[2]) ? 4'b0110 : 4'b0010;
																assign node43198 = (inp[2]) ? 4'b0010 : 4'b0110;
															assign node43201 = (inp[2]) ? node43205 : node43202;
																assign node43202 = (inp[13]) ? 4'b0110 : 4'b0010;
																assign node43205 = (inp[13]) ? 4'b0010 : 4'b0110;
							assign node43208 = (inp[15]) ? node43874 : node43209;
								assign node43209 = (inp[4]) ? node43597 : node43210;
									assign node43210 = (inp[5]) ? node43412 : node43211;
										assign node43211 = (inp[1]) ? node43323 : node43212;
											assign node43212 = (inp[0]) ? node43274 : node43213;
												assign node43213 = (inp[13]) ? node43243 : node43214;
													assign node43214 = (inp[2]) ? node43228 : node43215;
														assign node43215 = (inp[11]) ? node43221 : node43216;
															assign node43216 = (inp[10]) ? 4'b0110 : node43217;
																assign node43217 = (inp[9]) ? 4'b0111 : 4'b0110;
															assign node43221 = (inp[10]) ? node43225 : node43222;
																assign node43222 = (inp[9]) ? 4'b0111 : 4'b0110;
																assign node43225 = (inp[9]) ? 4'b0110 : 4'b0111;
														assign node43228 = (inp[11]) ? node43236 : node43229;
															assign node43229 = (inp[10]) ? node43233 : node43230;
																assign node43230 = (inp[9]) ? 4'b0010 : 4'b0011;
																assign node43233 = (inp[9]) ? 4'b0011 : 4'b0010;
															assign node43236 = (inp[9]) ? node43240 : node43237;
																assign node43237 = (inp[10]) ? 4'b0010 : 4'b0011;
																assign node43240 = (inp[10]) ? 4'b0011 : 4'b0010;
													assign node43243 = (inp[2]) ? node43259 : node43244;
														assign node43244 = (inp[11]) ? node43252 : node43245;
															assign node43245 = (inp[10]) ? node43249 : node43246;
																assign node43246 = (inp[9]) ? 4'b0010 : 4'b0011;
																assign node43249 = (inp[9]) ? 4'b0011 : 4'b0010;
															assign node43252 = (inp[9]) ? node43256 : node43253;
																assign node43253 = (inp[10]) ? 4'b0010 : 4'b0011;
																assign node43256 = (inp[10]) ? 4'b0011 : 4'b0010;
														assign node43259 = (inp[9]) ? node43267 : node43260;
															assign node43260 = (inp[11]) ? node43264 : node43261;
																assign node43261 = (inp[10]) ? 4'b0111 : 4'b0110;
																assign node43264 = (inp[10]) ? 4'b0110 : 4'b0111;
															assign node43267 = (inp[10]) ? node43271 : node43268;
																assign node43268 = (inp[11]) ? 4'b0110 : 4'b0111;
																assign node43271 = (inp[11]) ? 4'b0111 : 4'b0110;
												assign node43274 = (inp[10]) ? node43296 : node43275;
													assign node43275 = (inp[9]) ? node43289 : node43276;
														assign node43276 = (inp[11]) ? node43282 : node43277;
															assign node43277 = (inp[13]) ? node43279 : 4'b0011;
																assign node43279 = (inp[2]) ? 4'b0111 : 4'b0011;
															assign node43282 = (inp[2]) ? node43286 : node43283;
																assign node43283 = (inp[13]) ? 4'b0010 : 4'b0111;
																assign node43286 = (inp[13]) ? 4'b0111 : 4'b0010;
														assign node43289 = (inp[11]) ? 4'b0011 : node43290;
															assign node43290 = (inp[13]) ? 4'b0010 : node43291;
																assign node43291 = (inp[2]) ? 4'b0010 : 4'b0111;
													assign node43296 = (inp[13]) ? node43312 : node43297;
														assign node43297 = (inp[2]) ? node43305 : node43298;
															assign node43298 = (inp[11]) ? node43302 : node43299;
																assign node43299 = (inp[9]) ? 4'b0110 : 4'b0111;
																assign node43302 = (inp[9]) ? 4'b0111 : 4'b0110;
															assign node43305 = (inp[9]) ? node43309 : node43306;
																assign node43306 = (inp[11]) ? 4'b0011 : 4'b0010;
																assign node43309 = (inp[11]) ? 4'b0010 : 4'b0011;
														assign node43312 = (inp[2]) ? node43320 : node43313;
															assign node43313 = (inp[9]) ? node43317 : node43314;
																assign node43314 = (inp[11]) ? 4'b0011 : 4'b0010;
																assign node43317 = (inp[11]) ? 4'b0010 : 4'b0011;
															assign node43320 = (inp[9]) ? 4'b0111 : 4'b0110;
											assign node43323 = (inp[9]) ? node43365 : node43324;
												assign node43324 = (inp[2]) ? node43344 : node43325;
													assign node43325 = (inp[13]) ? node43337 : node43326;
														assign node43326 = (inp[10]) ? node43332 : node43327;
															assign node43327 = (inp[0]) ? 4'b0111 : node43328;
																assign node43328 = (inp[11]) ? 4'b0111 : 4'b0110;
															assign node43332 = (inp[0]) ? 4'b0110 : node43333;
																assign node43333 = (inp[11]) ? 4'b0110 : 4'b0111;
														assign node43337 = (inp[10]) ? 4'b0011 : node43338;
															assign node43338 = (inp[11]) ? 4'b0010 : node43339;
																assign node43339 = (inp[0]) ? 4'b0010 : 4'b0011;
													assign node43344 = (inp[13]) ? node43354 : node43345;
														assign node43345 = (inp[10]) ? node43351 : node43346;
															assign node43346 = (inp[0]) ? 4'b0010 : node43347;
																assign node43347 = (inp[11]) ? 4'b0010 : 4'b0011;
															assign node43351 = (inp[0]) ? 4'b0011 : 4'b0010;
														assign node43354 = (inp[10]) ? node43360 : node43355;
															assign node43355 = (inp[0]) ? node43357 : 4'b0111;
																assign node43357 = (inp[11]) ? 4'b0110 : 4'b0111;
															assign node43360 = (inp[0]) ? node43362 : 4'b0110;
																assign node43362 = (inp[11]) ? 4'b0111 : 4'b0110;
												assign node43365 = (inp[0]) ? node43393 : node43366;
													assign node43366 = (inp[10]) ? node43382 : node43367;
														assign node43367 = (inp[11]) ? node43375 : node43368;
															assign node43368 = (inp[13]) ? node43372 : node43369;
																assign node43369 = (inp[2]) ? 4'b0010 : 4'b0111;
																assign node43372 = (inp[2]) ? 4'b0110 : 4'b0010;
															assign node43375 = (inp[2]) ? node43379 : node43376;
																assign node43376 = (inp[13]) ? 4'b0011 : 4'b0110;
																assign node43379 = (inp[13]) ? 4'b0110 : 4'b0011;
														assign node43382 = (inp[13]) ? node43388 : node43383;
															assign node43383 = (inp[2]) ? node43385 : 4'b0110;
																assign node43385 = (inp[11]) ? 4'b0010 : 4'b0011;
															assign node43388 = (inp[2]) ? 4'b0111 : node43389;
																assign node43389 = (inp[11]) ? 4'b0010 : 4'b0011;
													assign node43393 = (inp[10]) ? node43403 : node43394;
														assign node43394 = (inp[2]) ? node43398 : node43395;
															assign node43395 = (inp[13]) ? 4'b0011 : 4'b0110;
															assign node43398 = (inp[13]) ? node43400 : 4'b0011;
																assign node43400 = (inp[11]) ? 4'b0111 : 4'b0110;
														assign node43403 = (inp[13]) ? node43407 : node43404;
															assign node43404 = (inp[2]) ? 4'b0010 : 4'b0111;
															assign node43407 = (inp[2]) ? node43409 : 4'b0010;
																assign node43409 = (inp[11]) ? 4'b0110 : 4'b0111;
										assign node43412 = (inp[9]) ? node43508 : node43413;
											assign node43413 = (inp[10]) ? node43461 : node43414;
												assign node43414 = (inp[11]) ? node43438 : node43415;
													assign node43415 = (inp[0]) ? node43431 : node43416;
														assign node43416 = (inp[1]) ? node43424 : node43417;
															assign node43417 = (inp[2]) ? node43421 : node43418;
																assign node43418 = (inp[13]) ? 4'b0011 : 4'b0110;
																assign node43421 = (inp[13]) ? 4'b0111 : 4'b0011;
															assign node43424 = (inp[13]) ? node43428 : node43425;
																assign node43425 = (inp[2]) ? 4'b0110 : 4'b0011;
																assign node43428 = (inp[2]) ? 4'b0011 : 4'b0110;
														assign node43431 = (inp[1]) ? node43433 : 4'b0111;
															assign node43433 = (inp[13]) ? node43435 : 4'b0111;
																assign node43435 = (inp[2]) ? 4'b0010 : 4'b0111;
													assign node43438 = (inp[13]) ? node43452 : node43439;
														assign node43439 = (inp[0]) ? node43445 : node43440;
															assign node43440 = (inp[2]) ? node43442 : 4'b0111;
																assign node43442 = (inp[1]) ? 4'b0111 : 4'b0010;
															assign node43445 = (inp[2]) ? node43449 : node43446;
																assign node43446 = (inp[1]) ? 4'b0010 : 4'b0111;
																assign node43449 = (inp[1]) ? 4'b0111 : 4'b0010;
														assign node43452 = (inp[2]) ? node43456 : node43453;
															assign node43453 = (inp[1]) ? 4'b0111 : 4'b0010;
															assign node43456 = (inp[1]) ? 4'b0010 : node43457;
																assign node43457 = (inp[0]) ? 4'b0110 : 4'b0111;
												assign node43461 = (inp[1]) ? node43489 : node43462;
													assign node43462 = (inp[11]) ? node43474 : node43463;
														assign node43463 = (inp[2]) ? node43469 : node43464;
															assign node43464 = (inp[13]) ? 4'b0011 : node43465;
																assign node43465 = (inp[0]) ? 4'b0110 : 4'b0111;
															assign node43469 = (inp[13]) ? 4'b0110 : node43470;
																assign node43470 = (inp[0]) ? 4'b0011 : 4'b0010;
														assign node43474 = (inp[0]) ? node43482 : node43475;
															assign node43475 = (inp[13]) ? node43479 : node43476;
																assign node43476 = (inp[2]) ? 4'b0011 : 4'b0110;
																assign node43479 = (inp[2]) ? 4'b0110 : 4'b0011;
															assign node43482 = (inp[13]) ? node43486 : node43483;
																assign node43483 = (inp[2]) ? 4'b0011 : 4'b0110;
																assign node43486 = (inp[2]) ? 4'b0111 : 4'b0011;
													assign node43489 = (inp[11]) ? node43503 : node43490;
														assign node43490 = (inp[2]) ? node43496 : node43491;
															assign node43491 = (inp[13]) ? node43493 : 4'b0010;
																assign node43493 = (inp[0]) ? 4'b0110 : 4'b0111;
															assign node43496 = (inp[13]) ? node43500 : node43497;
																assign node43497 = (inp[0]) ? 4'b0110 : 4'b0111;
																assign node43500 = (inp[0]) ? 4'b0011 : 4'b0010;
														assign node43503 = (inp[2]) ? 4'b0110 : node43504;
															assign node43504 = (inp[13]) ? 4'b0110 : 4'b0011;
											assign node43508 = (inp[10]) ? node43552 : node43509;
												assign node43509 = (inp[11]) ? node43535 : node43510;
													assign node43510 = (inp[13]) ? node43522 : node43511;
														assign node43511 = (inp[0]) ? node43517 : node43512;
															assign node43512 = (inp[2]) ? node43514 : 4'b0010;
																assign node43514 = (inp[1]) ? 4'b0111 : 4'b0010;
															assign node43517 = (inp[1]) ? node43519 : 4'b0110;
																assign node43519 = (inp[2]) ? 4'b0110 : 4'b0010;
														assign node43522 = (inp[1]) ? node43528 : node43523;
															assign node43523 = (inp[2]) ? 4'b0110 : node43524;
																assign node43524 = (inp[0]) ? 4'b0011 : 4'b0010;
															assign node43528 = (inp[2]) ? node43532 : node43529;
																assign node43529 = (inp[0]) ? 4'b0110 : 4'b0111;
																assign node43532 = (inp[0]) ? 4'b0011 : 4'b0010;
													assign node43535 = (inp[2]) ? node43545 : node43536;
														assign node43536 = (inp[13]) ? node43542 : node43537;
															assign node43537 = (inp[1]) ? node43539 : 4'b0110;
																assign node43539 = (inp[0]) ? 4'b0011 : 4'b0010;
															assign node43542 = (inp[1]) ? 4'b0110 : 4'b0011;
														assign node43545 = (inp[1]) ? 4'b0011 : node43546;
															assign node43546 = (inp[0]) ? node43548 : 4'b0110;
																assign node43548 = (inp[13]) ? 4'b0111 : 4'b0011;
												assign node43552 = (inp[0]) ? node43574 : node43553;
													assign node43553 = (inp[13]) ? node43563 : node43554;
														assign node43554 = (inp[11]) ? node43556 : 4'b0110;
															assign node43556 = (inp[2]) ? node43560 : node43557;
																assign node43557 = (inp[1]) ? 4'b0011 : 4'b0111;
																assign node43560 = (inp[1]) ? 4'b0111 : 4'b0010;
														assign node43563 = (inp[2]) ? node43571 : node43564;
															assign node43564 = (inp[1]) ? node43568 : node43565;
																assign node43565 = (inp[11]) ? 4'b0010 : 4'b0011;
																assign node43568 = (inp[11]) ? 4'b0111 : 4'b0110;
															assign node43571 = (inp[1]) ? 4'b0011 : 4'b0111;
													assign node43574 = (inp[2]) ? node43590 : node43575;
														assign node43575 = (inp[11]) ? node43583 : node43576;
															assign node43576 = (inp[1]) ? node43580 : node43577;
																assign node43577 = (inp[13]) ? 4'b0010 : 4'b0111;
																assign node43580 = (inp[13]) ? 4'b0111 : 4'b0011;
															assign node43583 = (inp[13]) ? node43587 : node43584;
																assign node43584 = (inp[1]) ? 4'b0010 : 4'b0111;
																assign node43587 = (inp[1]) ? 4'b0111 : 4'b0010;
														assign node43590 = (inp[1]) ? 4'b0010 : node43591;
															assign node43591 = (inp[13]) ? node43593 : 4'b0010;
																assign node43593 = (inp[11]) ? 4'b0110 : 4'b0111;
									assign node43597 = (inp[10]) ? node43749 : node43598;
										assign node43598 = (inp[9]) ? node43678 : node43599;
											assign node43599 = (inp[11]) ? node43639 : node43600;
												assign node43600 = (inp[13]) ? node43624 : node43601;
													assign node43601 = (inp[2]) ? node43611 : node43602;
														assign node43602 = (inp[1]) ? 4'b0000 : node43603;
															assign node43603 = (inp[0]) ? node43607 : node43604;
																assign node43604 = (inp[5]) ? 4'b0001 : 4'b0101;
																assign node43607 = (inp[5]) ? 4'b0000 : 4'b0100;
														assign node43611 = (inp[5]) ? node43619 : node43612;
															assign node43612 = (inp[1]) ? node43616 : node43613;
																assign node43613 = (inp[0]) ? 4'b0000 : 4'b0001;
																assign node43616 = (inp[0]) ? 4'b0101 : 4'b0100;
															assign node43619 = (inp[0]) ? node43621 : 4'b0100;
																assign node43621 = (inp[1]) ? 4'b0101 : 4'b0100;
													assign node43624 = (inp[2]) ? node43632 : node43625;
														assign node43625 = (inp[1]) ? node43629 : node43626;
															assign node43626 = (inp[5]) ? 4'b0101 : 4'b0001;
															assign node43629 = (inp[0]) ? 4'b0100 : 4'b0101;
														assign node43632 = (inp[1]) ? node43636 : node43633;
															assign node43633 = (inp[5]) ? 4'b0001 : 4'b0101;
															assign node43636 = (inp[0]) ? 4'b0000 : 4'b0001;
												assign node43639 = (inp[13]) ? node43661 : node43640;
													assign node43640 = (inp[1]) ? node43656 : node43641;
														assign node43641 = (inp[0]) ? node43649 : node43642;
															assign node43642 = (inp[2]) ? node43646 : node43643;
																assign node43643 = (inp[5]) ? 4'b0000 : 4'b0100;
																assign node43646 = (inp[5]) ? 4'b0100 : 4'b0000;
															assign node43649 = (inp[2]) ? node43653 : node43650;
																assign node43650 = (inp[5]) ? 4'b0000 : 4'b0100;
																assign node43653 = (inp[5]) ? 4'b0101 : 4'b0000;
														assign node43656 = (inp[2]) ? 4'b0101 : node43657;
															assign node43657 = (inp[0]) ? 4'b0001 : 4'b0000;
													assign node43661 = (inp[1]) ? node43675 : node43662;
														assign node43662 = (inp[0]) ? node43668 : node43663;
															assign node43663 = (inp[5]) ? 4'b0001 : node43664;
																assign node43664 = (inp[2]) ? 4'b0101 : 4'b0001;
															assign node43668 = (inp[5]) ? node43672 : node43669;
																assign node43669 = (inp[2]) ? 4'b0100 : 4'b0001;
																assign node43672 = (inp[2]) ? 4'b0000 : 4'b0100;
														assign node43675 = (inp[2]) ? 4'b0000 : 4'b0100;
											assign node43678 = (inp[1]) ? node43726 : node43679;
												assign node43679 = (inp[13]) ? node43705 : node43680;
													assign node43680 = (inp[11]) ? node43696 : node43681;
														assign node43681 = (inp[0]) ? node43689 : node43682;
															assign node43682 = (inp[2]) ? node43686 : node43683;
																assign node43683 = (inp[5]) ? 4'b0000 : 4'b0100;
																assign node43686 = (inp[5]) ? 4'b0101 : 4'b0000;
															assign node43689 = (inp[2]) ? node43693 : node43690;
																assign node43690 = (inp[5]) ? 4'b0001 : 4'b0101;
																assign node43693 = (inp[5]) ? 4'b0101 : 4'b0001;
														assign node43696 = (inp[2]) ? node43700 : node43697;
															assign node43697 = (inp[5]) ? 4'b0001 : 4'b0101;
															assign node43700 = (inp[5]) ? node43702 : 4'b0001;
																assign node43702 = (inp[0]) ? 4'b0100 : 4'b0101;
													assign node43705 = (inp[11]) ? node43711 : node43706;
														assign node43706 = (inp[5]) ? 4'b0100 : node43707;
															assign node43707 = (inp[2]) ? 4'b0100 : 4'b0000;
														assign node43711 = (inp[0]) ? node43719 : node43712;
															assign node43712 = (inp[5]) ? node43716 : node43713;
																assign node43713 = (inp[2]) ? 4'b0100 : 4'b0000;
																assign node43716 = (inp[2]) ? 4'b0000 : 4'b0100;
															assign node43719 = (inp[2]) ? node43723 : node43720;
																assign node43720 = (inp[5]) ? 4'b0101 : 4'b0000;
																assign node43723 = (inp[5]) ? 4'b0001 : 4'b0101;
												assign node43726 = (inp[13]) ? node43738 : node43727;
													assign node43727 = (inp[2]) ? node43733 : node43728;
														assign node43728 = (inp[11]) ? node43730 : 4'b0001;
															assign node43730 = (inp[0]) ? 4'b0000 : 4'b0001;
														assign node43733 = (inp[11]) ? 4'b0100 : node43734;
															assign node43734 = (inp[0]) ? 4'b0100 : 4'b0101;
													assign node43738 = (inp[2]) ? node43744 : node43739;
														assign node43739 = (inp[11]) ? 4'b0101 : node43740;
															assign node43740 = (inp[0]) ? 4'b0101 : 4'b0100;
														assign node43744 = (inp[11]) ? 4'b0001 : node43745;
															assign node43745 = (inp[0]) ? 4'b0001 : 4'b0000;
										assign node43749 = (inp[9]) ? node43817 : node43750;
											assign node43750 = (inp[0]) ? node43786 : node43751;
												assign node43751 = (inp[1]) ? node43771 : node43752;
													assign node43752 = (inp[13]) ? node43762 : node43753;
														assign node43753 = (inp[11]) ? 4'b0101 : node43754;
															assign node43754 = (inp[5]) ? node43758 : node43755;
																assign node43755 = (inp[2]) ? 4'b0000 : 4'b0100;
																assign node43758 = (inp[2]) ? 4'b0101 : 4'b0000;
														assign node43762 = (inp[2]) ? node43768 : node43763;
															assign node43763 = (inp[5]) ? 4'b0100 : node43764;
																assign node43764 = (inp[11]) ? 4'b0000 : 4'b0001;
															assign node43768 = (inp[5]) ? 4'b0000 : 4'b0100;
													assign node43771 = (inp[11]) ? node43779 : node43772;
														assign node43772 = (inp[13]) ? node43776 : node43773;
															assign node43773 = (inp[5]) ? 4'b0101 : 4'b0001;
															assign node43776 = (inp[2]) ? 4'b0000 : 4'b0100;
														assign node43779 = (inp[13]) ? node43783 : node43780;
															assign node43780 = (inp[2]) ? 4'b0100 : 4'b0001;
															assign node43783 = (inp[2]) ? 4'b0001 : 4'b0101;
												assign node43786 = (inp[13]) ? node43802 : node43787;
													assign node43787 = (inp[1]) ? node43797 : node43788;
														assign node43788 = (inp[5]) ? node43792 : node43789;
															assign node43789 = (inp[2]) ? 4'b0001 : 4'b0101;
															assign node43792 = (inp[2]) ? node43794 : 4'b0001;
																assign node43794 = (inp[11]) ? 4'b0100 : 4'b0101;
														assign node43797 = (inp[2]) ? 4'b0100 : node43798;
															assign node43798 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node43802 = (inp[1]) ? node43814 : node43803;
														assign node43803 = (inp[11]) ? node43809 : node43804;
															assign node43804 = (inp[2]) ? 4'b0000 : node43805;
																assign node43805 = (inp[5]) ? 4'b0100 : 4'b0000;
															assign node43809 = (inp[2]) ? 4'b0101 : node43810;
																assign node43810 = (inp[5]) ? 4'b0101 : 4'b0000;
														assign node43814 = (inp[2]) ? 4'b0001 : 4'b0101;
											assign node43817 = (inp[2]) ? node43845 : node43818;
												assign node43818 = (inp[13]) ? node43832 : node43819;
													assign node43819 = (inp[1]) ? node43827 : node43820;
														assign node43820 = (inp[5]) ? node43822 : 4'b0100;
															assign node43822 = (inp[11]) ? 4'b0000 : node43823;
																assign node43823 = (inp[0]) ? 4'b0000 : 4'b0001;
														assign node43827 = (inp[0]) ? node43829 : 4'b0000;
															assign node43829 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node43832 = (inp[1]) ? node43842 : node43833;
														assign node43833 = (inp[5]) ? node43837 : node43834;
															assign node43834 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node43837 = (inp[0]) ? node43839 : 4'b0101;
																assign node43839 = (inp[11]) ? 4'b0100 : 4'b0101;
														assign node43842 = (inp[0]) ? 4'b0100 : 4'b0101;
												assign node43845 = (inp[13]) ? node43859 : node43846;
													assign node43846 = (inp[1]) ? node43854 : node43847;
														assign node43847 = (inp[5]) ? 4'b0100 : node43848;
															assign node43848 = (inp[11]) ? 4'b0000 : node43849;
																assign node43849 = (inp[0]) ? 4'b0000 : 4'b0001;
														assign node43854 = (inp[0]) ? 4'b0101 : node43855;
															assign node43855 = (inp[11]) ? 4'b0101 : 4'b0100;
													assign node43859 = (inp[1]) ? node43869 : node43860;
														assign node43860 = (inp[5]) ? node43866 : node43861;
															assign node43861 = (inp[11]) ? node43863 : 4'b0101;
																assign node43863 = (inp[0]) ? 4'b0100 : 4'b0101;
															assign node43866 = (inp[11]) ? 4'b0000 : 4'b0001;
														assign node43869 = (inp[0]) ? 4'b0000 : node43870;
															assign node43870 = (inp[11]) ? 4'b0000 : 4'b0001;
								assign node43874 = (inp[10]) ? node44206 : node43875;
									assign node43875 = (inp[9]) ? node44037 : node43876;
										assign node43876 = (inp[0]) ? node43956 : node43877;
											assign node43877 = (inp[11]) ? node43917 : node43878;
												assign node43878 = (inp[4]) ? node43896 : node43879;
													assign node43879 = (inp[2]) ? node43887 : node43880;
														assign node43880 = (inp[13]) ? 4'b0100 : node43881;
															assign node43881 = (inp[1]) ? node43883 : 4'b0101;
																assign node43883 = (inp[5]) ? 4'b0000 : 4'b0001;
														assign node43887 = (inp[13]) ? node43891 : node43888;
															assign node43888 = (inp[1]) ? 4'b0101 : 4'b0000;
															assign node43891 = (inp[5]) ? 4'b0001 : node43892;
																assign node43892 = (inp[1]) ? 4'b0001 : 4'b0101;
													assign node43896 = (inp[13]) ? node43908 : node43897;
														assign node43897 = (inp[2]) ? node43903 : node43898;
															assign node43898 = (inp[5]) ? 4'b0001 : node43899;
																assign node43899 = (inp[1]) ? 4'b0001 : 4'b0101;
															assign node43903 = (inp[5]) ? 4'b0101 : node43904;
																assign node43904 = (inp[1]) ? 4'b0101 : 4'b0001;
														assign node43908 = (inp[2]) ? node43912 : node43909;
															assign node43909 = (inp[5]) ? 4'b0101 : 4'b0001;
															assign node43912 = (inp[5]) ? 4'b0001 : node43913;
																assign node43913 = (inp[1]) ? 4'b0001 : 4'b0101;
												assign node43917 = (inp[5]) ? node43945 : node43918;
													assign node43918 = (inp[1]) ? node43932 : node43919;
														assign node43919 = (inp[13]) ? node43925 : node43920;
															assign node43920 = (inp[2]) ? 4'b0001 : node43921;
																assign node43921 = (inp[4]) ? 4'b0101 : 4'b0100;
															assign node43925 = (inp[2]) ? node43929 : node43926;
																assign node43926 = (inp[4]) ? 4'b0001 : 4'b0000;
																assign node43929 = (inp[4]) ? 4'b0100 : 4'b0101;
														assign node43932 = (inp[4]) ? node43938 : node43933;
															assign node43933 = (inp[2]) ? node43935 : 4'b0000;
																assign node43935 = (inp[13]) ? 4'b0001 : 4'b0101;
															assign node43938 = (inp[13]) ? node43942 : node43939;
																assign node43939 = (inp[2]) ? 4'b0100 : 4'b0001;
																assign node43942 = (inp[2]) ? 4'b0000 : 4'b0100;
													assign node43945 = (inp[2]) ? node43953 : node43946;
														assign node43946 = (inp[13]) ? node43950 : node43947;
															assign node43947 = (inp[4]) ? 4'b0001 : 4'b0000;
															assign node43950 = (inp[4]) ? 4'b0100 : 4'b0101;
														assign node43953 = (inp[13]) ? 4'b0000 : 4'b0100;
											assign node43956 = (inp[11]) ? node43994 : node43957;
												assign node43957 = (inp[5]) ? node43983 : node43958;
													assign node43958 = (inp[13]) ? node43970 : node43959;
														assign node43959 = (inp[1]) ? node43965 : node43960;
															assign node43960 = (inp[2]) ? 4'b0001 : node43961;
																assign node43961 = (inp[4]) ? 4'b0101 : 4'b0100;
															assign node43965 = (inp[2]) ? node43967 : 4'b0001;
																assign node43967 = (inp[4]) ? 4'b0100 : 4'b0101;
														assign node43970 = (inp[1]) ? node43978 : node43971;
															assign node43971 = (inp[2]) ? node43975 : node43972;
																assign node43972 = (inp[4]) ? 4'b0001 : 4'b0000;
																assign node43975 = (inp[4]) ? 4'b0100 : 4'b0101;
															assign node43978 = (inp[2]) ? node43980 : 4'b0100;
																assign node43980 = (inp[4]) ? 4'b0000 : 4'b0001;
													assign node43983 = (inp[2]) ? node43991 : node43984;
														assign node43984 = (inp[13]) ? node43988 : node43985;
															assign node43985 = (inp[4]) ? 4'b0001 : 4'b0000;
															assign node43988 = (inp[4]) ? 4'b0100 : 4'b0101;
														assign node43991 = (inp[13]) ? 4'b0000 : 4'b0100;
												assign node43994 = (inp[4]) ? node44018 : node43995;
													assign node43995 = (inp[2]) ? node44007 : node43996;
														assign node43996 = (inp[5]) ? node44004 : node43997;
															assign node43997 = (inp[13]) ? node44001 : node43998;
																assign node43998 = (inp[1]) ? 4'b0000 : 4'b0100;
																assign node44001 = (inp[1]) ? 4'b0101 : 4'b0000;
															assign node44004 = (inp[13]) ? 4'b0101 : 4'b0001;
														assign node44007 = (inp[13]) ? node44013 : node44008;
															assign node44008 = (inp[5]) ? 4'b0100 : node44009;
																assign node44009 = (inp[1]) ? 4'b0100 : 4'b0001;
															assign node44013 = (inp[1]) ? 4'b0000 : node44014;
																assign node44014 = (inp[5]) ? 4'b0000 : 4'b0100;
													assign node44018 = (inp[13]) ? node44028 : node44019;
														assign node44019 = (inp[2]) ? node44023 : node44020;
															assign node44020 = (inp[1]) ? 4'b0000 : 4'b0100;
															assign node44023 = (inp[5]) ? 4'b0100 : node44024;
																assign node44024 = (inp[1]) ? 4'b0100 : 4'b0000;
														assign node44028 = (inp[2]) ? node44032 : node44029;
															assign node44029 = (inp[1]) ? 4'b0100 : 4'b0000;
															assign node44032 = (inp[1]) ? 4'b0000 : node44033;
																assign node44033 = (inp[5]) ? 4'b0000 : 4'b0100;
										assign node44037 = (inp[0]) ? node44117 : node44038;
											assign node44038 = (inp[11]) ? node44080 : node44039;
												assign node44039 = (inp[4]) ? node44059 : node44040;
													assign node44040 = (inp[2]) ? node44052 : node44041;
														assign node44041 = (inp[5]) ? node44049 : node44042;
															assign node44042 = (inp[1]) ? node44046 : node44043;
																assign node44043 = (inp[13]) ? 4'b0000 : 4'b0100;
																assign node44046 = (inp[13]) ? 4'b0101 : 4'b0000;
															assign node44049 = (inp[13]) ? 4'b0101 : 4'b0001;
														assign node44052 = (inp[13]) ? 4'b0000 : node44053;
															assign node44053 = (inp[1]) ? 4'b0100 : node44054;
																assign node44054 = (inp[5]) ? 4'b0100 : 4'b0001;
													assign node44059 = (inp[1]) ? node44067 : node44060;
														assign node44060 = (inp[2]) ? 4'b0000 : node44061;
															assign node44061 = (inp[13]) ? 4'b0000 : node44062;
																assign node44062 = (inp[5]) ? 4'b0000 : 4'b0100;
														assign node44067 = (inp[5]) ? node44073 : node44068;
															assign node44068 = (inp[13]) ? node44070 : 4'b0100;
																assign node44070 = (inp[2]) ? 4'b0000 : 4'b0100;
															assign node44073 = (inp[13]) ? node44077 : node44074;
																assign node44074 = (inp[2]) ? 4'b0100 : 4'b0000;
																assign node44077 = (inp[2]) ? 4'b0000 : 4'b0100;
												assign node44080 = (inp[5]) ? node44106 : node44081;
													assign node44081 = (inp[1]) ? node44093 : node44082;
														assign node44082 = (inp[13]) ? node44088 : node44083;
															assign node44083 = (inp[2]) ? 4'b0000 : node44084;
																assign node44084 = (inp[4]) ? 4'b0100 : 4'b0101;
															assign node44088 = (inp[2]) ? node44090 : 4'b0000;
																assign node44090 = (inp[4]) ? 4'b0101 : 4'b0100;
														assign node44093 = (inp[13]) ? node44101 : node44094;
															assign node44094 = (inp[2]) ? node44098 : node44095;
																assign node44095 = (inp[4]) ? 4'b0000 : 4'b0001;
																assign node44098 = (inp[4]) ? 4'b0101 : 4'b0100;
															assign node44101 = (inp[2]) ? node44103 : 4'b0101;
																assign node44103 = (inp[4]) ? 4'b0001 : 4'b0000;
													assign node44106 = (inp[2]) ? node44114 : node44107;
														assign node44107 = (inp[13]) ? node44111 : node44108;
															assign node44108 = (inp[4]) ? 4'b0000 : 4'b0001;
															assign node44111 = (inp[4]) ? 4'b0101 : 4'b0100;
														assign node44114 = (inp[13]) ? 4'b0001 : 4'b0101;
											assign node44117 = (inp[11]) ? node44153 : node44118;
												assign node44118 = (inp[5]) ? node44142 : node44119;
													assign node44119 = (inp[1]) ? node44131 : node44120;
														assign node44120 = (inp[4]) ? node44124 : node44121;
															assign node44121 = (inp[13]) ? 4'b0100 : 4'b0101;
															assign node44124 = (inp[13]) ? node44128 : node44125;
																assign node44125 = (inp[2]) ? 4'b0000 : 4'b0100;
																assign node44128 = (inp[2]) ? 4'b0101 : 4'b0000;
														assign node44131 = (inp[13]) ? node44137 : node44132;
															assign node44132 = (inp[2]) ? 4'b0100 : node44133;
																assign node44133 = (inp[4]) ? 4'b0000 : 4'b0001;
															assign node44137 = (inp[2]) ? node44139 : 4'b0101;
																assign node44139 = (inp[4]) ? 4'b0001 : 4'b0000;
													assign node44142 = (inp[2]) ? node44150 : node44143;
														assign node44143 = (inp[13]) ? node44147 : node44144;
															assign node44144 = (inp[4]) ? 4'b0000 : 4'b0001;
															assign node44147 = (inp[4]) ? 4'b0101 : 4'b0100;
														assign node44150 = (inp[13]) ? 4'b0001 : 4'b0101;
												assign node44153 = (inp[4]) ? node44177 : node44154;
													assign node44154 = (inp[2]) ? node44166 : node44155;
														assign node44155 = (inp[5]) ? node44163 : node44156;
															assign node44156 = (inp[13]) ? node44160 : node44157;
																assign node44157 = (inp[1]) ? 4'b0001 : 4'b0101;
																assign node44160 = (inp[1]) ? 4'b0100 : 4'b0001;
															assign node44163 = (inp[13]) ? 4'b0100 : 4'b0000;
														assign node44166 = (inp[13]) ? node44172 : node44167;
															assign node44167 = (inp[5]) ? 4'b0101 : node44168;
																assign node44168 = (inp[1]) ? 4'b0101 : 4'b0000;
															assign node44172 = (inp[5]) ? 4'b0001 : node44173;
																assign node44173 = (inp[1]) ? 4'b0001 : 4'b0101;
													assign node44177 = (inp[1]) ? node44191 : node44178;
														assign node44178 = (inp[13]) ? node44186 : node44179;
															assign node44179 = (inp[2]) ? node44183 : node44180;
																assign node44180 = (inp[5]) ? 4'b0001 : 4'b0101;
																assign node44183 = (inp[5]) ? 4'b0101 : 4'b0001;
															assign node44186 = (inp[5]) ? 4'b0101 : node44187;
																assign node44187 = (inp[2]) ? 4'b0101 : 4'b0001;
														assign node44191 = (inp[5]) ? node44199 : node44192;
															assign node44192 = (inp[2]) ? node44196 : node44193;
																assign node44193 = (inp[13]) ? 4'b0101 : 4'b0001;
																assign node44196 = (inp[13]) ? 4'b0001 : 4'b0101;
															assign node44199 = (inp[13]) ? node44203 : node44200;
																assign node44200 = (inp[2]) ? 4'b0101 : 4'b0001;
																assign node44203 = (inp[2]) ? 4'b0001 : 4'b0101;
									assign node44206 = (inp[9]) ? node44354 : node44207;
										assign node44207 = (inp[0]) ? node44293 : node44208;
											assign node44208 = (inp[11]) ? node44252 : node44209;
												assign node44209 = (inp[4]) ? node44231 : node44210;
													assign node44210 = (inp[2]) ? node44222 : node44211;
														assign node44211 = (inp[5]) ? node44219 : node44212;
															assign node44212 = (inp[13]) ? node44216 : node44213;
																assign node44213 = (inp[1]) ? 4'b0000 : 4'b0100;
																assign node44216 = (inp[1]) ? 4'b0101 : 4'b0000;
															assign node44219 = (inp[13]) ? 4'b0101 : 4'b0001;
														assign node44222 = (inp[13]) ? node44228 : node44223;
															assign node44223 = (inp[1]) ? 4'b0100 : node44224;
																assign node44224 = (inp[5]) ? 4'b0100 : 4'b0001;
															assign node44228 = (inp[1]) ? 4'b0000 : 4'b0100;
													assign node44231 = (inp[2]) ? node44243 : node44232;
														assign node44232 = (inp[13]) ? node44238 : node44233;
															assign node44233 = (inp[1]) ? 4'b0000 : node44234;
																assign node44234 = (inp[5]) ? 4'b0000 : 4'b0100;
															assign node44238 = (inp[5]) ? 4'b0100 : node44239;
																assign node44239 = (inp[1]) ? 4'b0100 : 4'b0000;
														assign node44243 = (inp[13]) ? node44249 : node44244;
															assign node44244 = (inp[5]) ? 4'b0100 : node44245;
																assign node44245 = (inp[1]) ? 4'b0100 : 4'b0000;
															assign node44249 = (inp[1]) ? 4'b0000 : 4'b0100;
												assign node44252 = (inp[5]) ? node44282 : node44253;
													assign node44253 = (inp[2]) ? node44267 : node44254;
														assign node44254 = (inp[4]) ? node44260 : node44255;
															assign node44255 = (inp[13]) ? 4'b0001 : node44256;
																assign node44256 = (inp[1]) ? 4'b0001 : 4'b0101;
															assign node44260 = (inp[13]) ? node44264 : node44261;
																assign node44261 = (inp[1]) ? 4'b0000 : 4'b0100;
																assign node44264 = (inp[1]) ? 4'b0101 : 4'b0000;
														assign node44267 = (inp[4]) ? node44275 : node44268;
															assign node44268 = (inp[13]) ? node44272 : node44269;
																assign node44269 = (inp[1]) ? 4'b0100 : 4'b0000;
																assign node44272 = (inp[1]) ? 4'b0000 : 4'b0100;
															assign node44275 = (inp[13]) ? node44279 : node44276;
																assign node44276 = (inp[1]) ? 4'b0101 : 4'b0000;
																assign node44279 = (inp[1]) ? 4'b0001 : 4'b0101;
													assign node44282 = (inp[2]) ? node44290 : node44283;
														assign node44283 = (inp[13]) ? node44287 : node44284;
															assign node44284 = (inp[4]) ? 4'b0000 : 4'b0001;
															assign node44287 = (inp[4]) ? 4'b0101 : 4'b0100;
														assign node44290 = (inp[13]) ? 4'b0001 : 4'b0101;
											assign node44293 = (inp[2]) ? node44333 : node44294;
												assign node44294 = (inp[13]) ? node44322 : node44295;
													assign node44295 = (inp[5]) ? node44307 : node44296;
														assign node44296 = (inp[1]) ? node44302 : node44297;
															assign node44297 = (inp[11]) ? 4'b0101 : node44298;
																assign node44298 = (inp[4]) ? 4'b0100 : 4'b0101;
															assign node44302 = (inp[4]) ? node44304 : 4'b0001;
																assign node44304 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node44307 = (inp[1]) ? node44315 : node44308;
															assign node44308 = (inp[4]) ? node44312 : node44309;
																assign node44309 = (inp[11]) ? 4'b0000 : 4'b0001;
																assign node44312 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node44315 = (inp[4]) ? node44319 : node44316;
																assign node44316 = (inp[11]) ? 4'b0000 : 4'b0001;
																assign node44319 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node44322 = (inp[5]) ? node44330 : node44323;
														assign node44323 = (inp[1]) ? node44327 : node44324;
															assign node44324 = (inp[4]) ? 4'b0000 : 4'b0001;
															assign node44327 = (inp[11]) ? 4'b0100 : 4'b0101;
														assign node44330 = (inp[4]) ? 4'b0101 : 4'b0100;
												assign node44333 = (inp[13]) ? node44345 : node44334;
													assign node44334 = (inp[5]) ? 4'b0101 : node44335;
														assign node44335 = (inp[1]) ? node44339 : node44336;
															assign node44336 = (inp[4]) ? 4'b0001 : 4'b0000;
															assign node44339 = (inp[11]) ? 4'b0101 : node44340;
																assign node44340 = (inp[4]) ? 4'b0101 : 4'b0100;
													assign node44345 = (inp[1]) ? node44349 : node44346;
														assign node44346 = (inp[5]) ? 4'b0001 : 4'b0101;
														assign node44349 = (inp[4]) ? 4'b0001 : node44350;
															assign node44350 = (inp[11]) ? 4'b0001 : 4'b0000;
										assign node44354 = (inp[11]) ? node44438 : node44355;
											assign node44355 = (inp[0]) ? node44397 : node44356;
												assign node44356 = (inp[4]) ? node44378 : node44357;
													assign node44357 = (inp[2]) ? node44369 : node44358;
														assign node44358 = (inp[5]) ? node44366 : node44359;
															assign node44359 = (inp[1]) ? node44363 : node44360;
																assign node44360 = (inp[13]) ? 4'b0001 : 4'b0101;
																assign node44363 = (inp[13]) ? 4'b0100 : 4'b0001;
															assign node44366 = (inp[13]) ? 4'b0100 : 4'b0000;
														assign node44369 = (inp[13]) ? node44373 : node44370;
															assign node44370 = (inp[1]) ? 4'b0101 : 4'b0000;
															assign node44373 = (inp[1]) ? 4'b0001 : node44374;
																assign node44374 = (inp[5]) ? 4'b0001 : 4'b0101;
													assign node44378 = (inp[5]) ? node44388 : node44379;
														assign node44379 = (inp[1]) ? node44381 : 4'b0001;
															assign node44381 = (inp[2]) ? node44385 : node44382;
																assign node44382 = (inp[13]) ? 4'b0101 : 4'b0001;
																assign node44385 = (inp[13]) ? 4'b0001 : 4'b0101;
														assign node44388 = (inp[1]) ? 4'b0101 : node44389;
															assign node44389 = (inp[13]) ? node44393 : node44390;
																assign node44390 = (inp[2]) ? 4'b0101 : 4'b0001;
																assign node44393 = (inp[2]) ? 4'b0001 : 4'b0101;
												assign node44397 = (inp[5]) ? node44427 : node44398;
													assign node44398 = (inp[1]) ? node44414 : node44399;
														assign node44399 = (inp[4]) ? node44407 : node44400;
															assign node44400 = (inp[2]) ? node44404 : node44401;
																assign node44401 = (inp[13]) ? 4'b0000 : 4'b0100;
																assign node44404 = (inp[13]) ? 4'b0101 : 4'b0001;
															assign node44407 = (inp[13]) ? node44411 : node44408;
																assign node44408 = (inp[2]) ? 4'b0001 : 4'b0101;
																assign node44411 = (inp[2]) ? 4'b0100 : 4'b0001;
														assign node44414 = (inp[13]) ? node44422 : node44415;
															assign node44415 = (inp[2]) ? node44419 : node44416;
																assign node44416 = (inp[4]) ? 4'b0001 : 4'b0000;
																assign node44419 = (inp[4]) ? 4'b0100 : 4'b0101;
															assign node44422 = (inp[2]) ? node44424 : 4'b0100;
																assign node44424 = (inp[4]) ? 4'b0000 : 4'b0001;
													assign node44427 = (inp[2]) ? node44435 : node44428;
														assign node44428 = (inp[13]) ? node44432 : node44429;
															assign node44429 = (inp[4]) ? 4'b0001 : 4'b0000;
															assign node44432 = (inp[4]) ? 4'b0100 : 4'b0101;
														assign node44435 = (inp[13]) ? 4'b0000 : 4'b0100;
											assign node44438 = (inp[0]) ? node44476 : node44439;
												assign node44439 = (inp[5]) ? node44465 : node44440;
													assign node44440 = (inp[1]) ? node44454 : node44441;
														assign node44441 = (inp[2]) ? node44449 : node44442;
															assign node44442 = (inp[4]) ? node44446 : node44443;
																assign node44443 = (inp[13]) ? 4'b0000 : 4'b0100;
																assign node44446 = (inp[13]) ? 4'b0001 : 4'b0101;
															assign node44449 = (inp[13]) ? node44451 : 4'b0001;
																assign node44451 = (inp[4]) ? 4'b0100 : 4'b0101;
														assign node44454 = (inp[2]) ? node44458 : node44455;
															assign node44455 = (inp[13]) ? 4'b0100 : 4'b0000;
															assign node44458 = (inp[4]) ? node44462 : node44459;
																assign node44459 = (inp[13]) ? 4'b0001 : 4'b0101;
																assign node44462 = (inp[13]) ? 4'b0000 : 4'b0100;
													assign node44465 = (inp[2]) ? node44473 : node44466;
														assign node44466 = (inp[13]) ? node44470 : node44467;
															assign node44467 = (inp[4]) ? 4'b0001 : 4'b0000;
															assign node44470 = (inp[4]) ? 4'b0100 : 4'b0101;
														assign node44473 = (inp[13]) ? 4'b0000 : 4'b0100;
												assign node44476 = (inp[4]) ? node44494 : node44477;
													assign node44477 = (inp[2]) ? node44487 : node44478;
														assign node44478 = (inp[5]) ? node44484 : node44479;
															assign node44479 = (inp[1]) ? 4'b0101 : node44480;
																assign node44480 = (inp[13]) ? 4'b0000 : 4'b0100;
															assign node44484 = (inp[13]) ? 4'b0101 : 4'b0001;
														assign node44487 = (inp[13]) ? node44489 : 4'b0100;
															assign node44489 = (inp[1]) ? 4'b0000 : node44490;
																assign node44490 = (inp[5]) ? 4'b0000 : 4'b0100;
													assign node44494 = (inp[5]) ? node44510 : node44495;
														assign node44495 = (inp[13]) ? node44503 : node44496;
															assign node44496 = (inp[2]) ? node44500 : node44497;
																assign node44497 = (inp[1]) ? 4'b0000 : 4'b0100;
																assign node44500 = (inp[1]) ? 4'b0100 : 4'b0000;
															assign node44503 = (inp[1]) ? node44507 : node44504;
																assign node44504 = (inp[2]) ? 4'b0100 : 4'b0000;
																assign node44507 = (inp[2]) ? 4'b0000 : 4'b0100;
														assign node44510 = (inp[1]) ? node44518 : node44511;
															assign node44511 = (inp[13]) ? node44515 : node44512;
																assign node44512 = (inp[2]) ? 4'b0100 : 4'b0000;
																assign node44515 = (inp[2]) ? 4'b0000 : 4'b0100;
															assign node44518 = (inp[13]) ? node44520 : 4'b0000;
																assign node44520 = (inp[2]) ? 4'b0000 : 4'b0100;
						assign node44523 = (inp[2]) ? node45059 : node44524;
							assign node44524 = (inp[15]) ? node45020 : node44525;
								assign node44525 = (inp[7]) ? node44757 : node44526;
									assign node44526 = (inp[5]) ? node44660 : node44527;
										assign node44527 = (inp[4]) ? node44591 : node44528;
											assign node44528 = (inp[11]) ? node44584 : node44529;
												assign node44529 = (inp[0]) ? node44559 : node44530;
													assign node44530 = (inp[10]) ? node44546 : node44531;
														assign node44531 = (inp[9]) ? node44539 : node44532;
															assign node44532 = (inp[1]) ? node44536 : node44533;
																assign node44533 = (inp[13]) ? 4'b0101 : 4'b0100;
																assign node44536 = (inp[13]) ? 4'b0100 : 4'b0101;
															assign node44539 = (inp[1]) ? node44543 : node44540;
																assign node44540 = (inp[13]) ? 4'b0101 : 4'b0100;
																assign node44543 = (inp[13]) ? 4'b0100 : 4'b0101;
														assign node44546 = (inp[9]) ? node44554 : node44547;
															assign node44547 = (inp[13]) ? node44551 : node44548;
																assign node44548 = (inp[1]) ? 4'b0100 : 4'b0101;
																assign node44551 = (inp[1]) ? 4'b0101 : 4'b0100;
															assign node44554 = (inp[1]) ? 4'b0100 : node44555;
																assign node44555 = (inp[13]) ? 4'b0100 : 4'b0101;
													assign node44559 = (inp[9]) ? node44575 : node44560;
														assign node44560 = (inp[13]) ? node44568 : node44561;
															assign node44561 = (inp[1]) ? node44565 : node44562;
																assign node44562 = (inp[10]) ? 4'b0101 : 4'b0100;
																assign node44565 = (inp[10]) ? 4'b0100 : 4'b0101;
															assign node44568 = (inp[1]) ? node44572 : node44569;
																assign node44569 = (inp[10]) ? 4'b0100 : 4'b0101;
																assign node44572 = (inp[10]) ? 4'b0101 : 4'b0100;
														assign node44575 = (inp[13]) ? 4'b0101 : node44576;
															assign node44576 = (inp[10]) ? node44580 : node44577;
																assign node44577 = (inp[1]) ? 4'b0101 : 4'b0100;
																assign node44580 = (inp[1]) ? 4'b0100 : 4'b0101;
												assign node44584 = (inp[13]) ? node44588 : node44585;
													assign node44585 = (inp[10]) ? 4'b0100 : 4'b0101;
													assign node44588 = (inp[10]) ? 4'b0101 : 4'b0100;
											assign node44591 = (inp[9]) ? node44635 : node44592;
												assign node44592 = (inp[0]) ? node44612 : node44593;
													assign node44593 = (inp[11]) ? node44605 : node44594;
														assign node44594 = (inp[1]) ? node44600 : node44595;
															assign node44595 = (inp[13]) ? node44597 : 4'b0000;
																assign node44597 = (inp[10]) ? 4'b0000 : 4'b0001;
															assign node44600 = (inp[13]) ? 4'b0001 : node44601;
																assign node44601 = (inp[10]) ? 4'b0001 : 4'b0000;
														assign node44605 = (inp[13]) ? 4'b0000 : node44606;
															assign node44606 = (inp[10]) ? node44608 : 4'b0000;
																assign node44608 = (inp[1]) ? 4'b0000 : 4'b0001;
													assign node44612 = (inp[10]) ? node44624 : node44613;
														assign node44613 = (inp[13]) ? node44619 : node44614;
															assign node44614 = (inp[11]) ? node44616 : 4'b0000;
																assign node44616 = (inp[1]) ? 4'b0001 : 4'b0000;
															assign node44619 = (inp[1]) ? node44621 : 4'b0001;
																assign node44621 = (inp[11]) ? 4'b0000 : 4'b0001;
														assign node44624 = (inp[13]) ? node44630 : node44625;
															assign node44625 = (inp[1]) ? node44627 : 4'b0001;
																assign node44627 = (inp[11]) ? 4'b0000 : 4'b0001;
															assign node44630 = (inp[11]) ? node44632 : 4'b0000;
																assign node44632 = (inp[1]) ? 4'b0001 : 4'b0000;
												assign node44635 = (inp[11]) ? node44643 : node44636;
													assign node44636 = (inp[10]) ? node44640 : node44637;
														assign node44637 = (inp[13]) ? 4'b0001 : 4'b0000;
														assign node44640 = (inp[13]) ? 4'b0000 : 4'b0001;
													assign node44643 = (inp[1]) ? node44651 : node44644;
														assign node44644 = (inp[13]) ? node44648 : node44645;
															assign node44645 = (inp[10]) ? 4'b0001 : 4'b0000;
															assign node44648 = (inp[10]) ? 4'b0000 : 4'b0001;
														assign node44651 = (inp[0]) ? node44653 : 4'b0001;
															assign node44653 = (inp[13]) ? node44657 : node44654;
																assign node44654 = (inp[10]) ? 4'b0000 : 4'b0001;
																assign node44657 = (inp[10]) ? 4'b0001 : 4'b0000;
										assign node44660 = (inp[10]) ? node44734 : node44661;
											assign node44661 = (inp[1]) ? node44689 : node44662;
												assign node44662 = (inp[11]) ? node44682 : node44663;
													assign node44663 = (inp[9]) ? node44669 : node44664;
														assign node44664 = (inp[4]) ? node44666 : 4'b0000;
															assign node44666 = (inp[13]) ? 4'b0000 : 4'b0001;
														assign node44669 = (inp[0]) ? node44677 : node44670;
															assign node44670 = (inp[4]) ? node44674 : node44671;
																assign node44671 = (inp[13]) ? 4'b0001 : 4'b0000;
																assign node44674 = (inp[13]) ? 4'b0000 : 4'b0001;
															assign node44677 = (inp[13]) ? node44679 : 4'b0000;
																assign node44679 = (inp[4]) ? 4'b0000 : 4'b0001;
													assign node44682 = (inp[4]) ? node44686 : node44683;
														assign node44683 = (inp[13]) ? 4'b0001 : 4'b0000;
														assign node44686 = (inp[13]) ? 4'b0000 : 4'b0001;
												assign node44689 = (inp[0]) ? node44705 : node44690;
													assign node44690 = (inp[9]) ? node44696 : node44691;
														assign node44691 = (inp[4]) ? node44693 : 4'b0000;
															assign node44693 = (inp[11]) ? 4'b0000 : 4'b0001;
														assign node44696 = (inp[4]) ? node44698 : 4'b0001;
															assign node44698 = (inp[13]) ? node44702 : node44699;
																assign node44699 = (inp[11]) ? 4'b0000 : 4'b0001;
																assign node44702 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node44705 = (inp[9]) ? node44721 : node44706;
														assign node44706 = (inp[11]) ? node44714 : node44707;
															assign node44707 = (inp[13]) ? node44711 : node44708;
																assign node44708 = (inp[4]) ? 4'b0001 : 4'b0000;
																assign node44711 = (inp[4]) ? 4'b0000 : 4'b0001;
															assign node44714 = (inp[13]) ? node44718 : node44715;
																assign node44715 = (inp[4]) ? 4'b0000 : 4'b0001;
																assign node44718 = (inp[4]) ? 4'b0001 : 4'b0000;
														assign node44721 = (inp[4]) ? node44727 : node44722;
															assign node44722 = (inp[11]) ? 4'b0000 : node44723;
																assign node44723 = (inp[13]) ? 4'b0001 : 4'b0000;
															assign node44727 = (inp[13]) ? node44731 : node44728;
																assign node44728 = (inp[11]) ? 4'b0000 : 4'b0001;
																assign node44731 = (inp[11]) ? 4'b0001 : 4'b0000;
											assign node44734 = (inp[4]) ? node44746 : node44735;
												assign node44735 = (inp[13]) ? node44741 : node44736;
													assign node44736 = (inp[1]) ? node44738 : 4'b0001;
														assign node44738 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node44741 = (inp[1]) ? node44743 : 4'b0000;
														assign node44743 = (inp[11]) ? 4'b0001 : 4'b0000;
												assign node44746 = (inp[13]) ? node44752 : node44747;
													assign node44747 = (inp[11]) ? node44749 : 4'b0000;
														assign node44749 = (inp[1]) ? 4'b0001 : 4'b0000;
													assign node44752 = (inp[11]) ? node44754 : 4'b0001;
														assign node44754 = (inp[1]) ? 4'b0000 : 4'b0001;
									assign node44757 = (inp[5]) ? node44863 : node44758;
										assign node44758 = (inp[4]) ? node44782 : node44759;
											assign node44759 = (inp[13]) ? node44771 : node44760;
												assign node44760 = (inp[10]) ? node44766 : node44761;
													assign node44761 = (inp[11]) ? 4'b0000 : node44762;
														assign node44762 = (inp[1]) ? 4'b0000 : 4'b0001;
													assign node44766 = (inp[11]) ? 4'b0001 : node44767;
														assign node44767 = (inp[1]) ? 4'b0001 : 4'b0000;
												assign node44771 = (inp[10]) ? node44777 : node44772;
													assign node44772 = (inp[1]) ? 4'b0001 : node44773;
														assign node44773 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node44777 = (inp[1]) ? 4'b0000 : node44778;
														assign node44778 = (inp[11]) ? 4'b0000 : 4'b0001;
											assign node44782 = (inp[1]) ? node44834 : node44783;
												assign node44783 = (inp[9]) ? node44811 : node44784;
													assign node44784 = (inp[13]) ? node44798 : node44785;
														assign node44785 = (inp[0]) ? node44793 : node44786;
															assign node44786 = (inp[11]) ? node44790 : node44787;
																assign node44787 = (inp[10]) ? 4'b0100 : 4'b0101;
																assign node44790 = (inp[10]) ? 4'b0101 : 4'b0100;
															assign node44793 = (inp[11]) ? node44795 : 4'b0100;
																assign node44795 = (inp[10]) ? 4'b0101 : 4'b0100;
														assign node44798 = (inp[0]) ? node44806 : node44799;
															assign node44799 = (inp[10]) ? node44803 : node44800;
																assign node44800 = (inp[11]) ? 4'b0101 : 4'b0100;
																assign node44803 = (inp[11]) ? 4'b0100 : 4'b0101;
															assign node44806 = (inp[10]) ? node44808 : 4'b0101;
																assign node44808 = (inp[11]) ? 4'b0100 : 4'b0101;
													assign node44811 = (inp[0]) ? node44821 : node44812;
														assign node44812 = (inp[11]) ? 4'b0100 : node44813;
															assign node44813 = (inp[10]) ? node44817 : node44814;
																assign node44814 = (inp[13]) ? 4'b0100 : 4'b0101;
																assign node44817 = (inp[13]) ? 4'b0101 : 4'b0100;
														assign node44821 = (inp[10]) ? node44829 : node44822;
															assign node44822 = (inp[13]) ? node44826 : node44823;
																assign node44823 = (inp[11]) ? 4'b0100 : 4'b0101;
																assign node44826 = (inp[11]) ? 4'b0101 : 4'b0100;
															assign node44829 = (inp[13]) ? 4'b0100 : node44830;
																assign node44830 = (inp[11]) ? 4'b0101 : 4'b0100;
												assign node44834 = (inp[11]) ? node44842 : node44835;
													assign node44835 = (inp[13]) ? node44839 : node44836;
														assign node44836 = (inp[10]) ? 4'b0101 : 4'b0100;
														assign node44839 = (inp[10]) ? 4'b0100 : 4'b0101;
													assign node44842 = (inp[9]) ? node44856 : node44843;
														assign node44843 = (inp[0]) ? node44851 : node44844;
															assign node44844 = (inp[13]) ? node44848 : node44845;
																assign node44845 = (inp[10]) ? 4'b0101 : 4'b0100;
																assign node44848 = (inp[10]) ? 4'b0100 : 4'b0101;
															assign node44851 = (inp[10]) ? node44853 : 4'b0101;
																assign node44853 = (inp[13]) ? 4'b0100 : 4'b0101;
														assign node44856 = (inp[13]) ? node44860 : node44857;
															assign node44857 = (inp[10]) ? 4'b0101 : 4'b0100;
															assign node44860 = (inp[10]) ? 4'b0100 : 4'b0101;
										assign node44863 = (inp[11]) ? node44943 : node44864;
											assign node44864 = (inp[0]) ? node44912 : node44865;
												assign node44865 = (inp[1]) ? node44897 : node44866;
													assign node44866 = (inp[9]) ? node44882 : node44867;
														assign node44867 = (inp[13]) ? node44875 : node44868;
															assign node44868 = (inp[10]) ? node44872 : node44869;
																assign node44869 = (inp[4]) ? 4'b0101 : 4'b0100;
																assign node44872 = (inp[4]) ? 4'b0100 : 4'b0101;
															assign node44875 = (inp[4]) ? node44879 : node44876;
																assign node44876 = (inp[10]) ? 4'b0100 : 4'b0101;
																assign node44879 = (inp[10]) ? 4'b0101 : 4'b0100;
														assign node44882 = (inp[10]) ? node44890 : node44883;
															assign node44883 = (inp[13]) ? node44887 : node44884;
																assign node44884 = (inp[4]) ? 4'b0101 : 4'b0100;
																assign node44887 = (inp[4]) ? 4'b0100 : 4'b0101;
															assign node44890 = (inp[13]) ? node44894 : node44891;
																assign node44891 = (inp[4]) ? 4'b0100 : 4'b0101;
																assign node44894 = (inp[4]) ? 4'b0101 : 4'b0100;
													assign node44897 = (inp[13]) ? node44905 : node44898;
														assign node44898 = (inp[4]) ? node44902 : node44899;
															assign node44899 = (inp[10]) ? 4'b0100 : 4'b0101;
															assign node44902 = (inp[10]) ? 4'b0101 : 4'b0100;
														assign node44905 = (inp[4]) ? node44909 : node44906;
															assign node44906 = (inp[10]) ? 4'b0101 : 4'b0100;
															assign node44909 = (inp[10]) ? 4'b0100 : 4'b0101;
												assign node44912 = (inp[10]) ? node44928 : node44913;
													assign node44913 = (inp[13]) ? node44921 : node44914;
														assign node44914 = (inp[1]) ? node44918 : node44915;
															assign node44915 = (inp[4]) ? 4'b0101 : 4'b0100;
															assign node44918 = (inp[4]) ? 4'b0100 : 4'b0101;
														assign node44921 = (inp[1]) ? node44925 : node44922;
															assign node44922 = (inp[4]) ? 4'b0100 : 4'b0101;
															assign node44925 = (inp[4]) ? 4'b0101 : 4'b0100;
													assign node44928 = (inp[4]) ? node44936 : node44929;
														assign node44929 = (inp[13]) ? node44933 : node44930;
															assign node44930 = (inp[1]) ? 4'b0100 : 4'b0101;
															assign node44933 = (inp[1]) ? 4'b0101 : 4'b0100;
														assign node44936 = (inp[9]) ? 4'b0100 : node44937;
															assign node44937 = (inp[13]) ? node44939 : 4'b0100;
																assign node44939 = (inp[1]) ? 4'b0100 : 4'b0101;
											assign node44943 = (inp[9]) ? node44971 : node44944;
												assign node44944 = (inp[10]) ? node44964 : node44945;
													assign node44945 = (inp[1]) ? node44957 : node44946;
														assign node44946 = (inp[0]) ? node44952 : node44947;
															assign node44947 = (inp[4]) ? 4'b0100 : node44948;
																assign node44948 = (inp[13]) ? 4'b0100 : 4'b0101;
															assign node44952 = (inp[13]) ? node44954 : 4'b0101;
																assign node44954 = (inp[4]) ? 4'b0101 : 4'b0100;
														assign node44957 = (inp[13]) ? node44961 : node44958;
															assign node44958 = (inp[4]) ? 4'b0100 : 4'b0101;
															assign node44961 = (inp[4]) ? 4'b0101 : 4'b0100;
													assign node44964 = (inp[13]) ? node44968 : node44965;
														assign node44965 = (inp[4]) ? 4'b0101 : 4'b0100;
														assign node44968 = (inp[4]) ? 4'b0100 : 4'b0101;
												assign node44971 = (inp[4]) ? node44995 : node44972;
													assign node44972 = (inp[0]) ? node44986 : node44973;
														assign node44973 = (inp[1]) ? node44979 : node44974;
															assign node44974 = (inp[13]) ? 4'b0100 : node44975;
																assign node44975 = (inp[10]) ? 4'b0100 : 4'b0101;
															assign node44979 = (inp[10]) ? node44983 : node44980;
																assign node44980 = (inp[13]) ? 4'b0100 : 4'b0101;
																assign node44983 = (inp[13]) ? 4'b0101 : 4'b0100;
														assign node44986 = (inp[1]) ? node44988 : 4'b0101;
															assign node44988 = (inp[13]) ? node44992 : node44989;
																assign node44989 = (inp[10]) ? 4'b0100 : 4'b0101;
																assign node44992 = (inp[10]) ? 4'b0101 : 4'b0100;
													assign node44995 = (inp[1]) ? node45011 : node44996;
														assign node44996 = (inp[0]) ? node45004 : node44997;
															assign node44997 = (inp[13]) ? node45001 : node44998;
																assign node44998 = (inp[10]) ? 4'b0101 : 4'b0100;
																assign node45001 = (inp[10]) ? 4'b0100 : 4'b0101;
															assign node45004 = (inp[13]) ? node45008 : node45005;
																assign node45005 = (inp[10]) ? 4'b0101 : 4'b0100;
																assign node45008 = (inp[10]) ? 4'b0100 : 4'b0101;
														assign node45011 = (inp[0]) ? 4'b0100 : node45012;
															assign node45012 = (inp[10]) ? node45016 : node45013;
																assign node45013 = (inp[13]) ? 4'b0101 : 4'b0100;
																assign node45016 = (inp[13]) ? 4'b0100 : 4'b0101;
								assign node45020 = (inp[7]) ? node45044 : node45021;
									assign node45021 = (inp[10]) ? node45031 : node45022;
										assign node45022 = (inp[5]) ? node45028 : node45023;
											assign node45023 = (inp[4]) ? 4'b0100 : node45024;
												assign node45024 = (inp[11]) ? 4'b0101 : 4'b0100;
											assign node45028 = (inp[4]) ? 4'b0101 : 4'b0100;
										assign node45031 = (inp[11]) ? node45037 : node45032;
											assign node45032 = (inp[5]) ? node45034 : 4'b0101;
												assign node45034 = (inp[4]) ? 4'b0100 : 4'b0101;
											assign node45037 = (inp[4]) ? node45041 : node45038;
												assign node45038 = (inp[5]) ? 4'b0101 : 4'b0100;
												assign node45041 = (inp[5]) ? 4'b0100 : 4'b0101;
									assign node45044 = (inp[10]) ? node45052 : node45045;
										assign node45045 = (inp[4]) ? 4'b0101 : node45046;
											assign node45046 = (inp[11]) ? 4'b0100 : node45047;
												assign node45047 = (inp[5]) ? 4'b0100 : 4'b0101;
										assign node45052 = (inp[4]) ? 4'b0100 : node45053;
											assign node45053 = (inp[5]) ? 4'b0101 : node45054;
												assign node45054 = (inp[11]) ? 4'b0101 : 4'b0100;
							assign node45059 = (inp[15]) ? node45347 : node45060;
								assign node45060 = (inp[7]) ? node45246 : node45061;
									assign node45061 = (inp[4]) ? node45109 : node45062;
										assign node45062 = (inp[5]) ? node45086 : node45063;
											assign node45063 = (inp[13]) ? node45075 : node45064;
												assign node45064 = (inp[10]) ? node45070 : node45065;
													assign node45065 = (inp[1]) ? 4'b0000 : node45066;
														assign node45066 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node45070 = (inp[11]) ? 4'b0001 : node45071;
														assign node45071 = (inp[1]) ? 4'b0001 : 4'b0000;
												assign node45075 = (inp[10]) ? node45081 : node45076;
													assign node45076 = (inp[11]) ? 4'b0001 : node45077;
														assign node45077 = (inp[1]) ? 4'b0001 : 4'b0000;
													assign node45081 = (inp[11]) ? 4'b0000 : node45082;
														assign node45082 = (inp[1]) ? 4'b0000 : 4'b0001;
											assign node45086 = (inp[13]) ? node45098 : node45087;
												assign node45087 = (inp[10]) ? node45093 : node45088;
													assign node45088 = (inp[11]) ? 4'b0100 : node45089;
														assign node45089 = (inp[1]) ? 4'b0100 : 4'b0101;
													assign node45093 = (inp[1]) ? 4'b0101 : node45094;
														assign node45094 = (inp[11]) ? 4'b0101 : 4'b0100;
												assign node45098 = (inp[10]) ? node45104 : node45099;
													assign node45099 = (inp[11]) ? 4'b0101 : node45100;
														assign node45100 = (inp[1]) ? 4'b0101 : 4'b0100;
													assign node45104 = (inp[11]) ? 4'b0100 : node45105;
														assign node45105 = (inp[1]) ? 4'b0100 : 4'b0101;
										assign node45109 = (inp[0]) ? node45191 : node45110;
											assign node45110 = (inp[1]) ? node45158 : node45111;
												assign node45111 = (inp[5]) ? node45135 : node45112;
													assign node45112 = (inp[11]) ? node45120 : node45113;
														assign node45113 = (inp[13]) ? node45117 : node45114;
															assign node45114 = (inp[10]) ? 4'b0101 : 4'b0100;
															assign node45117 = (inp[10]) ? 4'b0100 : 4'b0101;
														assign node45120 = (inp[9]) ? node45128 : node45121;
															assign node45121 = (inp[10]) ? node45125 : node45122;
																assign node45122 = (inp[13]) ? 4'b0100 : 4'b0101;
																assign node45125 = (inp[13]) ? 4'b0101 : 4'b0100;
															assign node45128 = (inp[10]) ? node45132 : node45129;
																assign node45129 = (inp[13]) ? 4'b0100 : 4'b0101;
																assign node45132 = (inp[13]) ? 4'b0101 : 4'b0100;
													assign node45135 = (inp[13]) ? node45151 : node45136;
														assign node45136 = (inp[9]) ? node45144 : node45137;
															assign node45137 = (inp[10]) ? node45141 : node45138;
																assign node45138 = (inp[11]) ? 4'b0100 : 4'b0101;
																assign node45141 = (inp[11]) ? 4'b0101 : 4'b0100;
															assign node45144 = (inp[11]) ? node45148 : node45145;
																assign node45145 = (inp[10]) ? 4'b0100 : 4'b0101;
																assign node45148 = (inp[10]) ? 4'b0101 : 4'b0100;
														assign node45151 = (inp[10]) ? node45155 : node45152;
															assign node45152 = (inp[11]) ? 4'b0101 : 4'b0100;
															assign node45155 = (inp[11]) ? 4'b0100 : 4'b0101;
												assign node45158 = (inp[11]) ? node45174 : node45159;
													assign node45159 = (inp[5]) ? node45167 : node45160;
														assign node45160 = (inp[10]) ? node45164 : node45161;
															assign node45161 = (inp[13]) ? 4'b0100 : 4'b0101;
															assign node45164 = (inp[13]) ? 4'b0101 : 4'b0100;
														assign node45167 = (inp[10]) ? node45171 : node45168;
															assign node45168 = (inp[13]) ? 4'b0101 : 4'b0100;
															assign node45171 = (inp[13]) ? 4'b0100 : 4'b0101;
													assign node45174 = (inp[10]) ? node45182 : node45175;
														assign node45175 = (inp[13]) ? node45179 : node45176;
															assign node45176 = (inp[5]) ? 4'b0100 : 4'b0101;
															assign node45179 = (inp[5]) ? 4'b0101 : 4'b0100;
														assign node45182 = (inp[9]) ? node45184 : 4'b0100;
															assign node45184 = (inp[13]) ? node45188 : node45185;
																assign node45185 = (inp[5]) ? 4'b0101 : 4'b0100;
																assign node45188 = (inp[5]) ? 4'b0100 : 4'b0101;
											assign node45191 = (inp[1]) ? node45231 : node45192;
												assign node45192 = (inp[11]) ? node45208 : node45193;
													assign node45193 = (inp[5]) ? node45201 : node45194;
														assign node45194 = (inp[13]) ? node45198 : node45195;
															assign node45195 = (inp[10]) ? 4'b0101 : 4'b0100;
															assign node45198 = (inp[10]) ? 4'b0100 : 4'b0101;
														assign node45201 = (inp[13]) ? node45205 : node45202;
															assign node45202 = (inp[10]) ? 4'b0100 : 4'b0101;
															assign node45205 = (inp[10]) ? 4'b0101 : 4'b0100;
													assign node45208 = (inp[10]) ? node45224 : node45209;
														assign node45209 = (inp[9]) ? node45217 : node45210;
															assign node45210 = (inp[5]) ? node45214 : node45211;
																assign node45211 = (inp[13]) ? 4'b0100 : 4'b0101;
																assign node45214 = (inp[13]) ? 4'b0101 : 4'b0100;
															assign node45217 = (inp[5]) ? node45221 : node45218;
																assign node45218 = (inp[13]) ? 4'b0100 : 4'b0101;
																assign node45221 = (inp[13]) ? 4'b0101 : 4'b0100;
														assign node45224 = (inp[13]) ? node45228 : node45225;
															assign node45225 = (inp[5]) ? 4'b0101 : 4'b0100;
															assign node45228 = (inp[5]) ? 4'b0100 : 4'b0101;
												assign node45231 = (inp[13]) ? node45239 : node45232;
													assign node45232 = (inp[10]) ? node45236 : node45233;
														assign node45233 = (inp[5]) ? 4'b0100 : 4'b0101;
														assign node45236 = (inp[5]) ? 4'b0101 : 4'b0100;
													assign node45239 = (inp[5]) ? node45243 : node45240;
														assign node45240 = (inp[10]) ? 4'b0101 : 4'b0100;
														assign node45243 = (inp[10]) ? 4'b0100 : 4'b0101;
									assign node45246 = (inp[5]) ? node45324 : node45247;
										assign node45247 = (inp[4]) ? node45271 : node45248;
											assign node45248 = (inp[10]) ? node45260 : node45249;
												assign node45249 = (inp[13]) ? node45255 : node45250;
													assign node45250 = (inp[1]) ? node45252 : 4'b0101;
														assign node45252 = (inp[11]) ? 4'b0100 : 4'b0101;
													assign node45255 = (inp[1]) ? node45257 : 4'b0100;
														assign node45257 = (inp[11]) ? 4'b0101 : 4'b0100;
												assign node45260 = (inp[13]) ? node45266 : node45261;
													assign node45261 = (inp[11]) ? node45263 : 4'b0100;
														assign node45263 = (inp[1]) ? 4'b0101 : 4'b0100;
													assign node45266 = (inp[1]) ? node45268 : 4'b0101;
														assign node45268 = (inp[11]) ? 4'b0100 : 4'b0101;
											assign node45271 = (inp[1]) ? node45309 : node45272;
												assign node45272 = (inp[9]) ? node45294 : node45273;
													assign node45273 = (inp[0]) ? node45281 : node45274;
														assign node45274 = (inp[10]) ? 4'b0001 : node45275;
															assign node45275 = (inp[11]) ? node45277 : 4'b0001;
																assign node45277 = (inp[13]) ? 4'b0001 : 4'b0000;
														assign node45281 = (inp[10]) ? node45287 : node45282;
															assign node45282 = (inp[11]) ? 4'b0001 : node45283;
																assign node45283 = (inp[13]) ? 4'b0000 : 4'b0001;
															assign node45287 = (inp[13]) ? node45291 : node45288;
																assign node45288 = (inp[11]) ? 4'b0001 : 4'b0000;
																assign node45291 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node45294 = (inp[13]) ? node45302 : node45295;
														assign node45295 = (inp[10]) ? node45299 : node45296;
															assign node45296 = (inp[11]) ? 4'b0000 : 4'b0001;
															assign node45299 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node45302 = (inp[10]) ? node45306 : node45303;
															assign node45303 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node45306 = (inp[11]) ? 4'b0000 : 4'b0001;
												assign node45309 = (inp[9]) ? node45317 : node45310;
													assign node45310 = (inp[13]) ? node45314 : node45311;
														assign node45311 = (inp[10]) ? 4'b0001 : 4'b0000;
														assign node45314 = (inp[10]) ? 4'b0000 : 4'b0001;
													assign node45317 = (inp[10]) ? node45321 : node45318;
														assign node45318 = (inp[13]) ? 4'b0001 : 4'b0000;
														assign node45321 = (inp[13]) ? 4'b0000 : 4'b0001;
										assign node45324 = (inp[13]) ? node45336 : node45325;
											assign node45325 = (inp[10]) ? node45331 : node45326;
												assign node45326 = (inp[11]) ? 4'b0000 : node45327;
													assign node45327 = (inp[1]) ? 4'b0000 : 4'b0001;
												assign node45331 = (inp[1]) ? 4'b0001 : node45332;
													assign node45332 = (inp[11]) ? 4'b0001 : 4'b0000;
											assign node45336 = (inp[10]) ? node45342 : node45337;
												assign node45337 = (inp[1]) ? 4'b0001 : node45338;
													assign node45338 = (inp[11]) ? 4'b0001 : 4'b0000;
												assign node45342 = (inp[1]) ? 4'b0000 : node45343;
													assign node45343 = (inp[11]) ? 4'b0000 : 4'b0001;
								assign node45347 = (inp[10]) ? node45361 : node45348;
									assign node45348 = (inp[5]) ? 4'b0001 : node45349;
										assign node45349 = (inp[7]) ? node45355 : node45350;
											assign node45350 = (inp[4]) ? 4'b0000 : node45351;
												assign node45351 = (inp[11]) ? 4'b0000 : 4'b0001;
											assign node45355 = (inp[4]) ? 4'b0001 : node45356;
												assign node45356 = (inp[11]) ? 4'b0001 : 4'b0000;
									assign node45361 = (inp[5]) ? 4'b0000 : node45362;
										assign node45362 = (inp[7]) ? node45368 : node45363;
											assign node45363 = (inp[4]) ? 4'b0001 : node45364;
												assign node45364 = (inp[11]) ? 4'b0001 : 4'b0000;
											assign node45368 = (inp[4]) ? 4'b0000 : node45369;
												assign node45369 = (inp[11]) ? 4'b0000 : 4'b0001;
			assign node45374 = (inp[4]) ? node51076 : node45375;
				assign node45375 = (inp[3]) ? node48909 : node45376;
					assign node45376 = (inp[7]) ? node47518 : node45377;
						assign node45377 = (inp[8]) ? node46337 : node45378;
							assign node45378 = (inp[5]) ? node45774 : node45379;
								assign node45379 = (inp[15]) ? node45565 : node45380;
									assign node45380 = (inp[12]) ? node45440 : node45381;
										assign node45381 = (inp[13]) ? node45425 : node45382;
											assign node45382 = (inp[1]) ? node45418 : node45383;
												assign node45383 = (inp[10]) ? node45403 : node45384;
													assign node45384 = (inp[11]) ? node45398 : node45385;
														assign node45385 = (inp[0]) ? node45393 : node45386;
															assign node45386 = (inp[2]) ? node45390 : node45387;
																assign node45387 = (inp[9]) ? 4'b0001 : 4'b0000;
																assign node45390 = (inp[9]) ? 4'b0000 : 4'b0001;
															assign node45393 = (inp[9]) ? node45395 : 4'b0000;
																assign node45395 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node45398 = (inp[9]) ? 4'b0000 : node45399;
															assign node45399 = (inp[2]) ? 4'b0001 : 4'b0000;
													assign node45403 = (inp[0]) ? node45411 : node45404;
														assign node45404 = (inp[9]) ? node45408 : node45405;
															assign node45405 = (inp[2]) ? 4'b0001 : 4'b0000;
															assign node45408 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node45411 = (inp[9]) ? node45415 : node45412;
															assign node45412 = (inp[2]) ? 4'b0001 : 4'b0000;
															assign node45415 = (inp[2]) ? 4'b0000 : 4'b0001;
												assign node45418 = (inp[9]) ? node45422 : node45419;
													assign node45419 = (inp[2]) ? 4'b0001 : 4'b0000;
													assign node45422 = (inp[2]) ? 4'b0000 : 4'b0001;
											assign node45425 = (inp[1]) ? node45433 : node45426;
												assign node45426 = (inp[2]) ? node45430 : node45427;
													assign node45427 = (inp[9]) ? 4'b0101 : 4'b0100;
													assign node45430 = (inp[9]) ? 4'b0100 : 4'b0101;
												assign node45433 = (inp[9]) ? node45437 : node45434;
													assign node45434 = (inp[2]) ? 4'b0101 : 4'b0100;
													assign node45437 = (inp[2]) ? 4'b0100 : 4'b0101;
										assign node45440 = (inp[13]) ? node45478 : node45441;
											assign node45441 = (inp[1]) ? node45471 : node45442;
												assign node45442 = (inp[10]) ? node45464 : node45443;
													assign node45443 = (inp[0]) ? node45457 : node45444;
														assign node45444 = (inp[11]) ? node45450 : node45445;
															assign node45445 = (inp[9]) ? node45447 : 4'b0101;
																assign node45447 = (inp[2]) ? 4'b0100 : 4'b0101;
															assign node45450 = (inp[2]) ? node45454 : node45451;
																assign node45451 = (inp[9]) ? 4'b0101 : 4'b0100;
																assign node45454 = (inp[9]) ? 4'b0100 : 4'b0101;
														assign node45457 = (inp[9]) ? node45461 : node45458;
															assign node45458 = (inp[2]) ? 4'b0101 : 4'b0100;
															assign node45461 = (inp[2]) ? 4'b0100 : 4'b0101;
													assign node45464 = (inp[2]) ? node45468 : node45465;
														assign node45465 = (inp[9]) ? 4'b0101 : 4'b0100;
														assign node45468 = (inp[9]) ? 4'b0100 : 4'b0101;
												assign node45471 = (inp[9]) ? node45475 : node45472;
													assign node45472 = (inp[2]) ? 4'b0100 : 4'b0101;
													assign node45475 = (inp[2]) ? 4'b0101 : 4'b0100;
											assign node45478 = (inp[0]) ? node45518 : node45479;
												assign node45479 = (inp[1]) ? node45495 : node45480;
													assign node45480 = (inp[10]) ? node45488 : node45481;
														assign node45481 = (inp[2]) ? node45485 : node45482;
															assign node45482 = (inp[9]) ? 4'b0001 : 4'b0000;
															assign node45485 = (inp[9]) ? 4'b0000 : 4'b0001;
														assign node45488 = (inp[9]) ? node45492 : node45489;
															assign node45489 = (inp[2]) ? 4'b0001 : 4'b0000;
															assign node45492 = (inp[2]) ? 4'b0000 : 4'b0001;
													assign node45495 = (inp[10]) ? node45503 : node45496;
														assign node45496 = (inp[9]) ? node45500 : node45497;
															assign node45497 = (inp[2]) ? 4'b0000 : 4'b0001;
															assign node45500 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node45503 = (inp[11]) ? node45511 : node45504;
															assign node45504 = (inp[9]) ? node45508 : node45505;
																assign node45505 = (inp[2]) ? 4'b0000 : 4'b0001;
																assign node45508 = (inp[2]) ? 4'b0001 : 4'b0000;
															assign node45511 = (inp[9]) ? node45515 : node45512;
																assign node45512 = (inp[2]) ? 4'b0000 : 4'b0001;
																assign node45515 = (inp[2]) ? 4'b0001 : 4'b0000;
												assign node45518 = (inp[10]) ? node45534 : node45519;
													assign node45519 = (inp[1]) ? node45527 : node45520;
														assign node45520 = (inp[2]) ? node45524 : node45521;
															assign node45521 = (inp[9]) ? 4'b0000 : 4'b0001;
															assign node45524 = (inp[9]) ? 4'b0001 : 4'b0000;
														assign node45527 = (inp[9]) ? node45531 : node45528;
															assign node45528 = (inp[2]) ? 4'b0001 : 4'b0000;
															assign node45531 = (inp[2]) ? 4'b0000 : 4'b0001;
													assign node45534 = (inp[1]) ? node45550 : node45535;
														assign node45535 = (inp[11]) ? node45543 : node45536;
															assign node45536 = (inp[2]) ? node45540 : node45537;
																assign node45537 = (inp[9]) ? 4'b0000 : 4'b0001;
																assign node45540 = (inp[9]) ? 4'b0001 : 4'b0000;
															assign node45543 = (inp[2]) ? node45547 : node45544;
																assign node45544 = (inp[9]) ? 4'b0000 : 4'b0001;
																assign node45547 = (inp[9]) ? 4'b0001 : 4'b0000;
														assign node45550 = (inp[11]) ? node45558 : node45551;
															assign node45551 = (inp[2]) ? node45555 : node45552;
																assign node45552 = (inp[9]) ? 4'b0001 : 4'b0000;
																assign node45555 = (inp[9]) ? 4'b0000 : 4'b0001;
															assign node45558 = (inp[2]) ? node45562 : node45559;
																assign node45559 = (inp[9]) ? 4'b0001 : 4'b0000;
																assign node45562 = (inp[9]) ? 4'b0000 : 4'b0001;
									assign node45565 = (inp[10]) ? node45657 : node45566;
										assign node45566 = (inp[13]) ? node45618 : node45567;
											assign node45567 = (inp[9]) ? node45599 : node45568;
												assign node45568 = (inp[2]) ? node45590 : node45569;
													assign node45569 = (inp[0]) ? node45583 : node45570;
														assign node45570 = (inp[11]) ? node45578 : node45571;
															assign node45571 = (inp[12]) ? node45575 : node45572;
																assign node45572 = (inp[1]) ? 4'b0100 : 4'b0000;
																assign node45575 = (inp[1]) ? 4'b0000 : 4'b0100;
															assign node45578 = (inp[12]) ? 4'b0100 : node45579;
																assign node45579 = (inp[1]) ? 4'b0100 : 4'b0000;
														assign node45583 = (inp[1]) ? node45587 : node45584;
															assign node45584 = (inp[12]) ? 4'b0100 : 4'b0000;
															assign node45587 = (inp[12]) ? 4'b0000 : 4'b0101;
													assign node45590 = (inp[1]) ? node45594 : node45591;
														assign node45591 = (inp[12]) ? 4'b0101 : 4'b0001;
														assign node45594 = (inp[12]) ? 4'b0001 : node45595;
															assign node45595 = (inp[0]) ? 4'b0100 : 4'b0101;
												assign node45599 = (inp[2]) ? node45609 : node45600;
													assign node45600 = (inp[1]) ? node45604 : node45601;
														assign node45601 = (inp[12]) ? 4'b0101 : 4'b0001;
														assign node45604 = (inp[12]) ? 4'b0001 : node45605;
															assign node45605 = (inp[0]) ? 4'b0100 : 4'b0101;
													assign node45609 = (inp[12]) ? node45615 : node45610;
														assign node45610 = (inp[1]) ? node45612 : 4'b0000;
															assign node45612 = (inp[0]) ? 4'b0101 : 4'b0100;
														assign node45615 = (inp[1]) ? 4'b0000 : 4'b0100;
											assign node45618 = (inp[2]) ? node45638 : node45619;
												assign node45619 = (inp[9]) ? node45629 : node45620;
													assign node45620 = (inp[12]) ? node45624 : node45621;
														assign node45621 = (inp[1]) ? 4'b0000 : 4'b0101;
														assign node45624 = (inp[1]) ? 4'b0101 : node45625;
															assign node45625 = (inp[0]) ? 4'b0000 : 4'b0001;
													assign node45629 = (inp[12]) ? node45633 : node45630;
														assign node45630 = (inp[1]) ? 4'b0001 : 4'b0100;
														assign node45633 = (inp[1]) ? 4'b0100 : node45634;
															assign node45634 = (inp[0]) ? 4'b0001 : 4'b0000;
												assign node45638 = (inp[9]) ? node45648 : node45639;
													assign node45639 = (inp[12]) ? node45643 : node45640;
														assign node45640 = (inp[1]) ? 4'b0001 : 4'b0100;
														assign node45643 = (inp[1]) ? 4'b0100 : node45644;
															assign node45644 = (inp[0]) ? 4'b0001 : 4'b0000;
													assign node45648 = (inp[1]) ? node45654 : node45649;
														assign node45649 = (inp[12]) ? node45651 : 4'b0101;
															assign node45651 = (inp[0]) ? 4'b0000 : 4'b0001;
														assign node45654 = (inp[12]) ? 4'b0101 : 4'b0000;
										assign node45657 = (inp[12]) ? node45711 : node45658;
											assign node45658 = (inp[2]) ? node45692 : node45659;
												assign node45659 = (inp[0]) ? node45675 : node45660;
													assign node45660 = (inp[9]) ? node45668 : node45661;
														assign node45661 = (inp[13]) ? node45665 : node45662;
															assign node45662 = (inp[1]) ? 4'b0100 : 4'b0000;
															assign node45665 = (inp[1]) ? 4'b0000 : 4'b0101;
														assign node45668 = (inp[13]) ? node45672 : node45669;
															assign node45669 = (inp[1]) ? 4'b0101 : 4'b0001;
															assign node45672 = (inp[1]) ? 4'b0001 : 4'b0100;
													assign node45675 = (inp[9]) ? node45683 : node45676;
														assign node45676 = (inp[13]) ? node45680 : node45677;
															assign node45677 = (inp[1]) ? 4'b0101 : 4'b0000;
															assign node45680 = (inp[1]) ? 4'b0000 : 4'b0101;
														assign node45683 = (inp[11]) ? 4'b0100 : node45684;
															assign node45684 = (inp[1]) ? node45688 : node45685;
																assign node45685 = (inp[13]) ? 4'b0100 : 4'b0001;
																assign node45688 = (inp[13]) ? 4'b0001 : 4'b0100;
												assign node45692 = (inp[9]) ? node45702 : node45693;
													assign node45693 = (inp[13]) ? node45699 : node45694;
														assign node45694 = (inp[1]) ? node45696 : 4'b0001;
															assign node45696 = (inp[0]) ? 4'b0100 : 4'b0101;
														assign node45699 = (inp[1]) ? 4'b0001 : 4'b0100;
													assign node45702 = (inp[1]) ? node45706 : node45703;
														assign node45703 = (inp[13]) ? 4'b0101 : 4'b0000;
														assign node45706 = (inp[13]) ? 4'b0000 : node45707;
															assign node45707 = (inp[0]) ? 4'b0101 : 4'b0100;
											assign node45711 = (inp[1]) ? node45757 : node45712;
												assign node45712 = (inp[13]) ? node45736 : node45713;
													assign node45713 = (inp[11]) ? node45729 : node45714;
														assign node45714 = (inp[0]) ? node45722 : node45715;
															assign node45715 = (inp[9]) ? node45719 : node45716;
																assign node45716 = (inp[2]) ? 4'b0101 : 4'b0100;
																assign node45719 = (inp[2]) ? 4'b0100 : 4'b0101;
															assign node45722 = (inp[9]) ? node45726 : node45723;
																assign node45723 = (inp[2]) ? 4'b0101 : 4'b0100;
																assign node45726 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node45729 = (inp[9]) ? node45733 : node45730;
															assign node45730 = (inp[2]) ? 4'b0101 : 4'b0100;
															assign node45733 = (inp[2]) ? 4'b0100 : 4'b0101;
													assign node45736 = (inp[9]) ? node45752 : node45737;
														assign node45737 = (inp[11]) ? node45745 : node45738;
															assign node45738 = (inp[0]) ? node45742 : node45739;
																assign node45739 = (inp[2]) ? 4'b0000 : 4'b0001;
																assign node45742 = (inp[2]) ? 4'b0001 : 4'b0000;
															assign node45745 = (inp[2]) ? node45749 : node45746;
																assign node45746 = (inp[0]) ? 4'b0000 : 4'b0001;
																assign node45749 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node45752 = (inp[2]) ? node45754 : 4'b0000;
															assign node45754 = (inp[0]) ? 4'b0000 : 4'b0001;
												assign node45757 = (inp[13]) ? node45767 : node45758;
													assign node45758 = (inp[0]) ? node45760 : 4'b0001;
														assign node45760 = (inp[11]) ? 4'b0000 : node45761;
															assign node45761 = (inp[9]) ? 4'b0001 : node45762;
																assign node45762 = (inp[2]) ? 4'b0001 : 4'b0000;
													assign node45767 = (inp[9]) ? node45771 : node45768;
														assign node45768 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node45771 = (inp[2]) ? 4'b0101 : 4'b0100;
								assign node45774 = (inp[0]) ? node46052 : node45775;
									assign node45775 = (inp[10]) ? node45887 : node45776;
										assign node45776 = (inp[9]) ? node45834 : node45777;
											assign node45777 = (inp[2]) ? node45807 : node45778;
												assign node45778 = (inp[13]) ? node45792 : node45779;
													assign node45779 = (inp[12]) ? node45785 : node45780;
														assign node45780 = (inp[15]) ? node45782 : 4'b0000;
															assign node45782 = (inp[1]) ? 4'b0101 : 4'b0000;
														assign node45785 = (inp[15]) ? node45789 : node45786;
															assign node45786 = (inp[11]) ? 4'b0101 : 4'b0100;
															assign node45789 = (inp[1]) ? 4'b0000 : 4'b0100;
													assign node45792 = (inp[12]) ? node45800 : node45793;
														assign node45793 = (inp[1]) ? node45797 : node45794;
															assign node45794 = (inp[15]) ? 4'b0101 : 4'b0100;
															assign node45797 = (inp[15]) ? 4'b0000 : 4'b0100;
														assign node45800 = (inp[1]) ? node45804 : node45801;
															assign node45801 = (inp[15]) ? 4'b0000 : 4'b0001;
															assign node45804 = (inp[15]) ? 4'b0101 : 4'b0000;
												assign node45807 = (inp[13]) ? node45821 : node45808;
													assign node45808 = (inp[12]) ? node45814 : node45809;
														assign node45809 = (inp[1]) ? node45811 : 4'b0001;
															assign node45811 = (inp[15]) ? 4'b0100 : 4'b0001;
														assign node45814 = (inp[15]) ? node45818 : node45815;
															assign node45815 = (inp[1]) ? 4'b0100 : 4'b0101;
															assign node45818 = (inp[1]) ? 4'b0001 : 4'b0101;
													assign node45821 = (inp[12]) ? node45827 : node45822;
														assign node45822 = (inp[15]) ? node45824 : 4'b0101;
															assign node45824 = (inp[1]) ? 4'b0001 : 4'b0100;
														assign node45827 = (inp[15]) ? node45831 : node45828;
															assign node45828 = (inp[1]) ? 4'b0001 : 4'b0000;
															assign node45831 = (inp[1]) ? 4'b0100 : 4'b0001;
											assign node45834 = (inp[2]) ? node45860 : node45835;
												assign node45835 = (inp[13]) ? node45847 : node45836;
													assign node45836 = (inp[12]) ? node45842 : node45837;
														assign node45837 = (inp[1]) ? node45839 : 4'b0001;
															assign node45839 = (inp[15]) ? 4'b0100 : 4'b0001;
														assign node45842 = (inp[1]) ? node45844 : 4'b0101;
															assign node45844 = (inp[11]) ? 4'b0100 : 4'b0001;
													assign node45847 = (inp[12]) ? node45853 : node45848;
														assign node45848 = (inp[15]) ? node45850 : 4'b0101;
															assign node45850 = (inp[1]) ? 4'b0001 : 4'b0100;
														assign node45853 = (inp[1]) ? node45857 : node45854;
															assign node45854 = (inp[15]) ? 4'b0001 : 4'b0000;
															assign node45857 = (inp[15]) ? 4'b0100 : 4'b0001;
												assign node45860 = (inp[15]) ? node45872 : node45861;
													assign node45861 = (inp[12]) ? node45865 : node45862;
														assign node45862 = (inp[13]) ? 4'b0100 : 4'b0000;
														assign node45865 = (inp[13]) ? node45869 : node45866;
															assign node45866 = (inp[1]) ? 4'b0101 : 4'b0100;
															assign node45869 = (inp[1]) ? 4'b0000 : 4'b0001;
													assign node45872 = (inp[12]) ? node45880 : node45873;
														assign node45873 = (inp[1]) ? node45877 : node45874;
															assign node45874 = (inp[13]) ? 4'b0101 : 4'b0000;
															assign node45877 = (inp[13]) ? 4'b0000 : 4'b0101;
														assign node45880 = (inp[1]) ? node45884 : node45881;
															assign node45881 = (inp[13]) ? 4'b0000 : 4'b0100;
															assign node45884 = (inp[13]) ? 4'b0101 : 4'b0000;
										assign node45887 = (inp[1]) ? node45989 : node45888;
											assign node45888 = (inp[11]) ? node45946 : node45889;
												assign node45889 = (inp[15]) ? node45919 : node45890;
													assign node45890 = (inp[12]) ? node45904 : node45891;
														assign node45891 = (inp[13]) ? node45897 : node45892;
															assign node45892 = (inp[9]) ? node45894 : 4'b0000;
																assign node45894 = (inp[2]) ? 4'b0000 : 4'b0001;
															assign node45897 = (inp[2]) ? node45901 : node45898;
																assign node45898 = (inp[9]) ? 4'b0101 : 4'b0100;
																assign node45901 = (inp[9]) ? 4'b0100 : 4'b0101;
														assign node45904 = (inp[13]) ? node45912 : node45905;
															assign node45905 = (inp[2]) ? node45909 : node45906;
																assign node45906 = (inp[9]) ? 4'b0101 : 4'b0100;
																assign node45909 = (inp[9]) ? 4'b0100 : 4'b0101;
															assign node45912 = (inp[9]) ? node45916 : node45913;
																assign node45913 = (inp[2]) ? 4'b0000 : 4'b0001;
																assign node45916 = (inp[2]) ? 4'b0001 : 4'b0000;
													assign node45919 = (inp[13]) ? node45933 : node45920;
														assign node45920 = (inp[12]) ? node45926 : node45921;
															assign node45921 = (inp[9]) ? 4'b0000 : node45922;
																assign node45922 = (inp[2]) ? 4'b0001 : 4'b0000;
															assign node45926 = (inp[9]) ? node45930 : node45927;
																assign node45927 = (inp[2]) ? 4'b0101 : 4'b0100;
																assign node45930 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node45933 = (inp[12]) ? node45941 : node45934;
															assign node45934 = (inp[2]) ? node45938 : node45935;
																assign node45935 = (inp[9]) ? 4'b0100 : 4'b0101;
																assign node45938 = (inp[9]) ? 4'b0101 : 4'b0100;
															assign node45941 = (inp[2]) ? 4'b0000 : node45942;
																assign node45942 = (inp[9]) ? 4'b0001 : 4'b0000;
												assign node45946 = (inp[12]) ? node45964 : node45947;
													assign node45947 = (inp[13]) ? node45955 : node45948;
														assign node45948 = (inp[2]) ? node45952 : node45949;
															assign node45949 = (inp[9]) ? 4'b0001 : 4'b0000;
															assign node45952 = (inp[9]) ? 4'b0000 : 4'b0001;
														assign node45955 = (inp[15]) ? 4'b0100 : node45956;
															assign node45956 = (inp[2]) ? node45960 : node45957;
																assign node45957 = (inp[9]) ? 4'b0101 : 4'b0100;
																assign node45960 = (inp[9]) ? 4'b0100 : 4'b0101;
													assign node45964 = (inp[13]) ? node45974 : node45965;
														assign node45965 = (inp[15]) ? node45967 : 4'b0100;
															assign node45967 = (inp[2]) ? node45971 : node45968;
																assign node45968 = (inp[9]) ? 4'b0101 : 4'b0100;
																assign node45971 = (inp[9]) ? 4'b0100 : 4'b0101;
														assign node45974 = (inp[15]) ? node45982 : node45975;
															assign node45975 = (inp[2]) ? node45979 : node45976;
																assign node45976 = (inp[9]) ? 4'b0000 : 4'b0001;
																assign node45979 = (inp[9]) ? 4'b0001 : 4'b0000;
															assign node45982 = (inp[2]) ? node45986 : node45983;
																assign node45983 = (inp[9]) ? 4'b0001 : 4'b0000;
																assign node45986 = (inp[9]) ? 4'b0000 : 4'b0001;
											assign node45989 = (inp[9]) ? node46021 : node45990;
												assign node45990 = (inp[2]) ? node46006 : node45991;
													assign node45991 = (inp[13]) ? node45999 : node45992;
														assign node45992 = (inp[15]) ? node45996 : node45993;
															assign node45993 = (inp[12]) ? 4'b0101 : 4'b0000;
															assign node45996 = (inp[12]) ? 4'b0000 : 4'b0101;
														assign node45999 = (inp[12]) ? node46003 : node46000;
															assign node46000 = (inp[15]) ? 4'b0000 : 4'b0100;
															assign node46003 = (inp[15]) ? 4'b0101 : 4'b0000;
													assign node46006 = (inp[12]) ? node46014 : node46007;
														assign node46007 = (inp[15]) ? node46011 : node46008;
															assign node46008 = (inp[13]) ? 4'b0101 : 4'b0001;
															assign node46011 = (inp[13]) ? 4'b0001 : 4'b0100;
														assign node46014 = (inp[13]) ? node46018 : node46015;
															assign node46015 = (inp[15]) ? 4'b0001 : 4'b0100;
															assign node46018 = (inp[15]) ? 4'b0100 : 4'b0001;
												assign node46021 = (inp[2]) ? node46037 : node46022;
													assign node46022 = (inp[15]) ? node46030 : node46023;
														assign node46023 = (inp[13]) ? node46027 : node46024;
															assign node46024 = (inp[12]) ? 4'b0100 : 4'b0001;
															assign node46027 = (inp[12]) ? 4'b0001 : 4'b0101;
														assign node46030 = (inp[12]) ? node46034 : node46031;
															assign node46031 = (inp[13]) ? 4'b0001 : 4'b0100;
															assign node46034 = (inp[13]) ? 4'b0100 : 4'b0001;
													assign node46037 = (inp[12]) ? node46045 : node46038;
														assign node46038 = (inp[15]) ? node46042 : node46039;
															assign node46039 = (inp[13]) ? 4'b0100 : 4'b0000;
															assign node46042 = (inp[13]) ? 4'b0000 : 4'b0101;
														assign node46045 = (inp[15]) ? node46049 : node46046;
															assign node46046 = (inp[13]) ? 4'b0000 : 4'b0101;
															assign node46049 = (inp[13]) ? 4'b0101 : 4'b0000;
									assign node46052 = (inp[10]) ? node46212 : node46053;
										assign node46053 = (inp[12]) ? node46123 : node46054;
											assign node46054 = (inp[13]) ? node46084 : node46055;
												assign node46055 = (inp[1]) ? node46071 : node46056;
													assign node46056 = (inp[11]) ? node46064 : node46057;
														assign node46057 = (inp[9]) ? node46061 : node46058;
															assign node46058 = (inp[2]) ? 4'b0000 : 4'b0001;
															assign node46061 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node46064 = (inp[2]) ? node46068 : node46065;
															assign node46065 = (inp[9]) ? 4'b0000 : 4'b0001;
															assign node46068 = (inp[9]) ? 4'b0001 : 4'b0000;
													assign node46071 = (inp[15]) ? node46079 : node46072;
														assign node46072 = (inp[2]) ? node46076 : node46073;
															assign node46073 = (inp[9]) ? 4'b0000 : 4'b0001;
															assign node46076 = (inp[9]) ? 4'b0001 : 4'b0000;
														assign node46079 = (inp[2]) ? 4'b0101 : node46080;
															assign node46080 = (inp[9]) ? 4'b0100 : 4'b0101;
												assign node46084 = (inp[15]) ? node46100 : node46085;
													assign node46085 = (inp[11]) ? node46093 : node46086;
														assign node46086 = (inp[9]) ? node46090 : node46087;
															assign node46087 = (inp[2]) ? 4'b0100 : 4'b0101;
															assign node46090 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node46093 = (inp[9]) ? node46097 : node46094;
															assign node46094 = (inp[2]) ? 4'b0100 : 4'b0101;
															assign node46097 = (inp[2]) ? 4'b0101 : 4'b0100;
													assign node46100 = (inp[1]) ? node46116 : node46101;
														assign node46101 = (inp[11]) ? node46109 : node46102;
															assign node46102 = (inp[2]) ? node46106 : node46103;
																assign node46103 = (inp[9]) ? 4'b0101 : 4'b0100;
																assign node46106 = (inp[9]) ? 4'b0100 : 4'b0101;
															assign node46109 = (inp[2]) ? node46113 : node46110;
																assign node46110 = (inp[9]) ? 4'b0101 : 4'b0100;
																assign node46113 = (inp[9]) ? 4'b0100 : 4'b0101;
														assign node46116 = (inp[2]) ? node46120 : node46117;
															assign node46117 = (inp[9]) ? 4'b0000 : 4'b0001;
															assign node46120 = (inp[9]) ? 4'b0001 : 4'b0000;
											assign node46123 = (inp[13]) ? node46163 : node46124;
												assign node46124 = (inp[15]) ? node46140 : node46125;
													assign node46125 = (inp[9]) ? node46133 : node46126;
														assign node46126 = (inp[1]) ? node46130 : node46127;
															assign node46127 = (inp[2]) ? 4'b0100 : 4'b0101;
															assign node46130 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node46133 = (inp[2]) ? node46137 : node46134;
															assign node46134 = (inp[1]) ? 4'b0101 : 4'b0100;
															assign node46137 = (inp[1]) ? 4'b0100 : 4'b0101;
													assign node46140 = (inp[1]) ? node46156 : node46141;
														assign node46141 = (inp[11]) ? node46149 : node46142;
															assign node46142 = (inp[2]) ? node46146 : node46143;
																assign node46143 = (inp[9]) ? 4'b0100 : 4'b0101;
																assign node46146 = (inp[9]) ? 4'b0101 : 4'b0100;
															assign node46149 = (inp[9]) ? node46153 : node46150;
																assign node46150 = (inp[2]) ? 4'b0100 : 4'b0101;
																assign node46153 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node46156 = (inp[2]) ? node46160 : node46157;
															assign node46157 = (inp[9]) ? 4'b0000 : 4'b0001;
															assign node46160 = (inp[9]) ? 4'b0001 : 4'b0000;
												assign node46163 = (inp[1]) ? node46195 : node46164;
													assign node46164 = (inp[11]) ? node46180 : node46165;
														assign node46165 = (inp[2]) ? node46173 : node46166;
															assign node46166 = (inp[9]) ? node46170 : node46167;
																assign node46167 = (inp[15]) ? 4'b0000 : 4'b0001;
																assign node46170 = (inp[15]) ? 4'b0001 : 4'b0000;
															assign node46173 = (inp[9]) ? node46177 : node46174;
																assign node46174 = (inp[15]) ? 4'b0001 : 4'b0000;
																assign node46177 = (inp[15]) ? 4'b0000 : 4'b0001;
														assign node46180 = (inp[2]) ? node46188 : node46181;
															assign node46181 = (inp[15]) ? node46185 : node46182;
																assign node46182 = (inp[9]) ? 4'b0000 : 4'b0001;
																assign node46185 = (inp[9]) ? 4'b0001 : 4'b0000;
															assign node46188 = (inp[9]) ? node46192 : node46189;
																assign node46189 = (inp[15]) ? 4'b0001 : 4'b0000;
																assign node46192 = (inp[15]) ? 4'b0000 : 4'b0001;
													assign node46195 = (inp[15]) ? node46201 : node46196;
														assign node46196 = (inp[9]) ? node46198 : 4'b0000;
															assign node46198 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node46201 = (inp[11]) ? node46207 : node46202;
															assign node46202 = (inp[9]) ? 4'b0100 : node46203;
																assign node46203 = (inp[2]) ? 4'b0101 : 4'b0100;
															assign node46207 = (inp[2]) ? node46209 : 4'b0101;
																assign node46209 = (inp[9]) ? 4'b0100 : 4'b0101;
										assign node46212 = (inp[12]) ? node46268 : node46213;
											assign node46213 = (inp[13]) ? node46245 : node46214;
												assign node46214 = (inp[1]) ? node46222 : node46215;
													assign node46215 = (inp[2]) ? node46219 : node46216;
														assign node46216 = (inp[9]) ? 4'b0000 : 4'b0001;
														assign node46219 = (inp[9]) ? 4'b0001 : 4'b0000;
													assign node46222 = (inp[15]) ? node46230 : node46223;
														assign node46223 = (inp[2]) ? node46227 : node46224;
															assign node46224 = (inp[9]) ? 4'b0000 : 4'b0001;
															assign node46227 = (inp[9]) ? 4'b0001 : 4'b0000;
														assign node46230 = (inp[11]) ? node46238 : node46231;
															assign node46231 = (inp[9]) ? node46235 : node46232;
																assign node46232 = (inp[2]) ? 4'b0100 : 4'b0101;
																assign node46235 = (inp[2]) ? 4'b0101 : 4'b0100;
															assign node46238 = (inp[2]) ? node46242 : node46239;
																assign node46239 = (inp[9]) ? 4'b0100 : 4'b0101;
																assign node46242 = (inp[9]) ? 4'b0101 : 4'b0100;
												assign node46245 = (inp[15]) ? node46253 : node46246;
													assign node46246 = (inp[9]) ? node46250 : node46247;
														assign node46247 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node46250 = (inp[2]) ? 4'b0101 : 4'b0100;
													assign node46253 = (inp[1]) ? node46261 : node46254;
														assign node46254 = (inp[2]) ? node46258 : node46255;
															assign node46255 = (inp[9]) ? 4'b0101 : 4'b0100;
															assign node46258 = (inp[9]) ? 4'b0100 : 4'b0101;
														assign node46261 = (inp[2]) ? node46265 : node46262;
															assign node46262 = (inp[9]) ? 4'b0000 : 4'b0001;
															assign node46265 = (inp[9]) ? 4'b0001 : 4'b0000;
											assign node46268 = (inp[13]) ? node46298 : node46269;
												assign node46269 = (inp[15]) ? node46285 : node46270;
													assign node46270 = (inp[9]) ? node46278 : node46271;
														assign node46271 = (inp[2]) ? node46275 : node46272;
															assign node46272 = (inp[1]) ? 4'b0100 : 4'b0101;
															assign node46275 = (inp[1]) ? 4'b0101 : 4'b0100;
														assign node46278 = (inp[1]) ? node46282 : node46279;
															assign node46279 = (inp[2]) ? 4'b0101 : 4'b0100;
															assign node46282 = (inp[2]) ? 4'b0100 : 4'b0101;
													assign node46285 = (inp[1]) ? node46291 : node46286;
														assign node46286 = (inp[9]) ? 4'b0101 : node46287;
															assign node46287 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node46291 = (inp[9]) ? node46295 : node46292;
															assign node46292 = (inp[2]) ? 4'b0000 : 4'b0001;
															assign node46295 = (inp[2]) ? 4'b0001 : 4'b0000;
												assign node46298 = (inp[1]) ? node46322 : node46299;
													assign node46299 = (inp[2]) ? node46307 : node46300;
														assign node46300 = (inp[15]) ? node46304 : node46301;
															assign node46301 = (inp[9]) ? 4'b0000 : 4'b0001;
															assign node46304 = (inp[9]) ? 4'b0001 : 4'b0000;
														assign node46307 = (inp[11]) ? node46315 : node46308;
															assign node46308 = (inp[15]) ? node46312 : node46309;
																assign node46309 = (inp[9]) ? 4'b0001 : 4'b0000;
																assign node46312 = (inp[9]) ? 4'b0000 : 4'b0001;
															assign node46315 = (inp[9]) ? node46319 : node46316;
																assign node46316 = (inp[15]) ? 4'b0001 : 4'b0000;
																assign node46319 = (inp[15]) ? 4'b0000 : 4'b0001;
													assign node46322 = (inp[15]) ? node46330 : node46323;
														assign node46323 = (inp[2]) ? node46327 : node46324;
															assign node46324 = (inp[9]) ? 4'b0001 : 4'b0000;
															assign node46327 = (inp[9]) ? 4'b0000 : 4'b0001;
														assign node46330 = (inp[11]) ? node46332 : 4'b0101;
															assign node46332 = (inp[9]) ? node46334 : 4'b0100;
																assign node46334 = (inp[2]) ? 4'b0100 : 4'b0101;
							assign node46337 = (inp[11]) ? node46925 : node46338;
								assign node46338 = (inp[9]) ? node46658 : node46339;
									assign node46339 = (inp[12]) ? node46493 : node46340;
										assign node46340 = (inp[1]) ? node46412 : node46341;
											assign node46341 = (inp[10]) ? node46379 : node46342;
												assign node46342 = (inp[0]) ? node46362 : node46343;
													assign node46343 = (inp[2]) ? node46353 : node46344;
														assign node46344 = (inp[13]) ? node46346 : 4'b0010;
															assign node46346 = (inp[5]) ? node46350 : node46347;
																assign node46347 = (inp[15]) ? 4'b0011 : 4'b0010;
																assign node46350 = (inp[15]) ? 4'b0010 : 4'b0011;
														assign node46353 = (inp[13]) ? node46355 : 4'b0011;
															assign node46355 = (inp[15]) ? node46359 : node46356;
																assign node46356 = (inp[5]) ? 4'b0010 : 4'b0011;
																assign node46359 = (inp[5]) ? 4'b0011 : 4'b0010;
													assign node46362 = (inp[2]) ? node46370 : node46363;
														assign node46363 = (inp[13]) ? node46365 : 4'b0011;
															assign node46365 = (inp[5]) ? node46367 : 4'b0011;
																assign node46367 = (inp[15]) ? 4'b0011 : 4'b0010;
														assign node46370 = (inp[13]) ? node46372 : 4'b0010;
															assign node46372 = (inp[5]) ? node46376 : node46373;
																assign node46373 = (inp[15]) ? 4'b0011 : 4'b0010;
																assign node46376 = (inp[15]) ? 4'b0010 : 4'b0011;
												assign node46379 = (inp[5]) ? node46395 : node46380;
													assign node46380 = (inp[15]) ? node46388 : node46381;
														assign node46381 = (inp[2]) ? node46385 : node46382;
															assign node46382 = (inp[0]) ? 4'b0011 : 4'b0010;
															assign node46385 = (inp[0]) ? 4'b0010 : 4'b0011;
														assign node46388 = (inp[2]) ? node46390 : 4'b0010;
															assign node46390 = (inp[0]) ? node46392 : 4'b0010;
																assign node46392 = (inp[13]) ? 4'b0011 : 4'b0010;
													assign node46395 = (inp[0]) ? node46407 : node46396;
														assign node46396 = (inp[2]) ? node46402 : node46397;
															assign node46397 = (inp[15]) ? 4'b0010 : node46398;
																assign node46398 = (inp[13]) ? 4'b0011 : 4'b0010;
															assign node46402 = (inp[13]) ? node46404 : 4'b0011;
																assign node46404 = (inp[15]) ? 4'b0011 : 4'b0010;
														assign node46407 = (inp[2]) ? 4'b0010 : node46408;
															assign node46408 = (inp[15]) ? 4'b0011 : 4'b0010;
											assign node46412 = (inp[13]) ? node46456 : node46413;
												assign node46413 = (inp[10]) ? node46437 : node46414;
													assign node46414 = (inp[0]) ? node46426 : node46415;
														assign node46415 = (inp[2]) ? node46421 : node46416;
															assign node46416 = (inp[5]) ? node46418 : 4'b0110;
																assign node46418 = (inp[15]) ? 4'b0111 : 4'b0110;
															assign node46421 = (inp[5]) ? node46423 : 4'b0111;
																assign node46423 = (inp[15]) ? 4'b0110 : 4'b0111;
														assign node46426 = (inp[2]) ? node46432 : node46427;
															assign node46427 = (inp[5]) ? node46429 : 4'b0111;
																assign node46429 = (inp[15]) ? 4'b0110 : 4'b0111;
															assign node46432 = (inp[15]) ? node46434 : 4'b0110;
																assign node46434 = (inp[5]) ? 4'b0111 : 4'b0110;
													assign node46437 = (inp[0]) ? node46449 : node46438;
														assign node46438 = (inp[2]) ? node46444 : node46439;
															assign node46439 = (inp[15]) ? node46441 : 4'b0110;
																assign node46441 = (inp[5]) ? 4'b0111 : 4'b0110;
															assign node46444 = (inp[5]) ? node46446 : 4'b0111;
																assign node46446 = (inp[15]) ? 4'b0110 : 4'b0111;
														assign node46449 = (inp[2]) ? 4'b0110 : node46450;
															assign node46450 = (inp[15]) ? node46452 : 4'b0111;
																assign node46452 = (inp[5]) ? 4'b0110 : 4'b0111;
												assign node46456 = (inp[15]) ? node46486 : node46457;
													assign node46457 = (inp[10]) ? node46471 : node46458;
														assign node46458 = (inp[2]) ? node46464 : node46459;
															assign node46459 = (inp[5]) ? 4'b0110 : node46460;
																assign node46460 = (inp[0]) ? 4'b0111 : 4'b0110;
															assign node46464 = (inp[5]) ? node46468 : node46465;
																assign node46465 = (inp[0]) ? 4'b0110 : 4'b0111;
																assign node46468 = (inp[0]) ? 4'b0111 : 4'b0110;
														assign node46471 = (inp[2]) ? node46479 : node46472;
															assign node46472 = (inp[5]) ? node46476 : node46473;
																assign node46473 = (inp[0]) ? 4'b0111 : 4'b0110;
																assign node46476 = (inp[0]) ? 4'b0110 : 4'b0111;
															assign node46479 = (inp[0]) ? node46483 : node46480;
																assign node46480 = (inp[5]) ? 4'b0110 : 4'b0111;
																assign node46483 = (inp[5]) ? 4'b0111 : 4'b0110;
													assign node46486 = (inp[0]) ? node46490 : node46487;
														assign node46487 = (inp[2]) ? 4'b0111 : 4'b0110;
														assign node46490 = (inp[2]) ? 4'b0110 : 4'b0111;
										assign node46493 = (inp[1]) ? node46577 : node46494;
											assign node46494 = (inp[13]) ? node46516 : node46495;
												assign node46495 = (inp[5]) ? node46509 : node46496;
													assign node46496 = (inp[10]) ? node46502 : node46497;
														assign node46497 = (inp[0]) ? node46499 : 4'b0110;
															assign node46499 = (inp[2]) ? 4'b0110 : 4'b0111;
														assign node46502 = (inp[2]) ? node46506 : node46503;
															assign node46503 = (inp[0]) ? 4'b0111 : 4'b0110;
															assign node46506 = (inp[0]) ? 4'b0110 : 4'b0111;
													assign node46509 = (inp[2]) ? node46513 : node46510;
														assign node46510 = (inp[0]) ? 4'b0111 : 4'b0110;
														assign node46513 = (inp[0]) ? 4'b0110 : 4'b0111;
												assign node46516 = (inp[5]) ? node46546 : node46517;
													assign node46517 = (inp[10]) ? node46533 : node46518;
														assign node46518 = (inp[15]) ? node46526 : node46519;
															assign node46519 = (inp[0]) ? node46523 : node46520;
																assign node46520 = (inp[2]) ? 4'b0111 : 4'b0110;
																assign node46523 = (inp[2]) ? 4'b0110 : 4'b0111;
															assign node46526 = (inp[0]) ? node46530 : node46527;
																assign node46527 = (inp[2]) ? 4'b0110 : 4'b0111;
																assign node46530 = (inp[2]) ? 4'b0111 : 4'b0110;
														assign node46533 = (inp[0]) ? node46539 : node46534;
															assign node46534 = (inp[15]) ? node46536 : 4'b0111;
																assign node46536 = (inp[2]) ? 4'b0110 : 4'b0111;
															assign node46539 = (inp[2]) ? node46543 : node46540;
																assign node46540 = (inp[15]) ? 4'b0110 : 4'b0111;
																assign node46543 = (inp[15]) ? 4'b0111 : 4'b0110;
													assign node46546 = (inp[0]) ? node46562 : node46547;
														assign node46547 = (inp[10]) ? node46555 : node46548;
															assign node46548 = (inp[15]) ? node46552 : node46549;
																assign node46549 = (inp[2]) ? 4'b0110 : 4'b0111;
																assign node46552 = (inp[2]) ? 4'b0111 : 4'b0110;
															assign node46555 = (inp[15]) ? node46559 : node46556;
																assign node46556 = (inp[2]) ? 4'b0110 : 4'b0111;
																assign node46559 = (inp[2]) ? 4'b0111 : 4'b0110;
														assign node46562 = (inp[10]) ? node46570 : node46563;
															assign node46563 = (inp[15]) ? node46567 : node46564;
																assign node46564 = (inp[2]) ? 4'b0111 : 4'b0110;
																assign node46567 = (inp[2]) ? 4'b0110 : 4'b0111;
															assign node46570 = (inp[15]) ? node46574 : node46571;
																assign node46571 = (inp[2]) ? 4'b0111 : 4'b0110;
																assign node46574 = (inp[2]) ? 4'b0110 : 4'b0111;
											assign node46577 = (inp[10]) ? node46615 : node46578;
												assign node46578 = (inp[5]) ? node46608 : node46579;
													assign node46579 = (inp[2]) ? node46595 : node46580;
														assign node46580 = (inp[15]) ? node46588 : node46581;
															assign node46581 = (inp[0]) ? node46585 : node46582;
																assign node46582 = (inp[13]) ? 4'b0010 : 4'b0011;
																assign node46585 = (inp[13]) ? 4'b0011 : 4'b0010;
															assign node46588 = (inp[0]) ? node46592 : node46589;
																assign node46589 = (inp[13]) ? 4'b0011 : 4'b0010;
																assign node46592 = (inp[13]) ? 4'b0010 : 4'b0011;
														assign node46595 = (inp[13]) ? node46603 : node46596;
															assign node46596 = (inp[15]) ? node46600 : node46597;
																assign node46597 = (inp[0]) ? 4'b0011 : 4'b0010;
																assign node46600 = (inp[0]) ? 4'b0010 : 4'b0011;
															assign node46603 = (inp[15]) ? node46605 : 4'b0011;
																assign node46605 = (inp[0]) ? 4'b0011 : 4'b0010;
													assign node46608 = (inp[0]) ? node46612 : node46609;
														assign node46609 = (inp[2]) ? 4'b0011 : 4'b0010;
														assign node46612 = (inp[2]) ? 4'b0010 : 4'b0011;
												assign node46615 = (inp[13]) ? node46639 : node46616;
													assign node46616 = (inp[5]) ? node46632 : node46617;
														assign node46617 = (inp[2]) ? node46625 : node46618;
															assign node46618 = (inp[15]) ? node46622 : node46619;
																assign node46619 = (inp[0]) ? 4'b0010 : 4'b0011;
																assign node46622 = (inp[0]) ? 4'b0011 : 4'b0010;
															assign node46625 = (inp[0]) ? node46629 : node46626;
																assign node46626 = (inp[15]) ? 4'b0011 : 4'b0010;
																assign node46629 = (inp[15]) ? 4'b0010 : 4'b0011;
														assign node46632 = (inp[2]) ? node46636 : node46633;
															assign node46633 = (inp[0]) ? 4'b0011 : 4'b0010;
															assign node46636 = (inp[0]) ? 4'b0010 : 4'b0011;
													assign node46639 = (inp[15]) ? node46645 : node46640;
														assign node46640 = (inp[2]) ? node46642 : 4'b0011;
															assign node46642 = (inp[0]) ? 4'b0010 : 4'b0011;
														assign node46645 = (inp[2]) ? node46653 : node46646;
															assign node46646 = (inp[5]) ? node46650 : node46647;
																assign node46647 = (inp[0]) ? 4'b0010 : 4'b0011;
																assign node46650 = (inp[0]) ? 4'b0011 : 4'b0010;
															assign node46653 = (inp[0]) ? 4'b0011 : node46654;
																assign node46654 = (inp[5]) ? 4'b0011 : 4'b0010;
									assign node46658 = (inp[12]) ? node46772 : node46659;
										assign node46659 = (inp[1]) ? node46723 : node46660;
											assign node46660 = (inp[15]) ? node46684 : node46661;
												assign node46661 = (inp[0]) ? node46673 : node46662;
													assign node46662 = (inp[2]) ? node46668 : node46663;
														assign node46663 = (inp[5]) ? node46665 : 4'b0010;
															assign node46665 = (inp[13]) ? 4'b0011 : 4'b0010;
														assign node46668 = (inp[5]) ? node46670 : 4'b0011;
															assign node46670 = (inp[13]) ? 4'b0010 : 4'b0011;
													assign node46673 = (inp[2]) ? node46679 : node46674;
														assign node46674 = (inp[5]) ? node46676 : 4'b0011;
															assign node46676 = (inp[13]) ? 4'b0010 : 4'b0011;
														assign node46679 = (inp[13]) ? node46681 : 4'b0010;
															assign node46681 = (inp[5]) ? 4'b0011 : 4'b0010;
												assign node46684 = (inp[10]) ? node46700 : node46685;
													assign node46685 = (inp[0]) ? node46693 : node46686;
														assign node46686 = (inp[2]) ? 4'b0011 : node46687;
															assign node46687 = (inp[13]) ? node46689 : 4'b0010;
																assign node46689 = (inp[5]) ? 4'b0010 : 4'b0011;
														assign node46693 = (inp[2]) ? node46695 : 4'b0011;
															assign node46695 = (inp[13]) ? node46697 : 4'b0010;
																assign node46697 = (inp[5]) ? 4'b0010 : 4'b0011;
													assign node46700 = (inp[13]) ? node46708 : node46701;
														assign node46701 = (inp[2]) ? node46705 : node46702;
															assign node46702 = (inp[0]) ? 4'b0011 : 4'b0010;
															assign node46705 = (inp[0]) ? 4'b0010 : 4'b0011;
														assign node46708 = (inp[2]) ? node46716 : node46709;
															assign node46709 = (inp[0]) ? node46713 : node46710;
																assign node46710 = (inp[5]) ? 4'b0010 : 4'b0011;
																assign node46713 = (inp[5]) ? 4'b0011 : 4'b0010;
															assign node46716 = (inp[5]) ? node46720 : node46717;
																assign node46717 = (inp[0]) ? 4'b0011 : 4'b0010;
																assign node46720 = (inp[0]) ? 4'b0010 : 4'b0011;
											assign node46723 = (inp[2]) ? node46745 : node46724;
												assign node46724 = (inp[0]) ? node46734 : node46725;
													assign node46725 = (inp[5]) ? node46727 : 4'b0110;
														assign node46727 = (inp[13]) ? node46731 : node46728;
															assign node46728 = (inp[15]) ? 4'b0111 : 4'b0110;
															assign node46731 = (inp[15]) ? 4'b0110 : 4'b0111;
													assign node46734 = (inp[5]) ? node46736 : 4'b0111;
														assign node46736 = (inp[10]) ? 4'b0111 : node46737;
															assign node46737 = (inp[15]) ? node46741 : node46738;
																assign node46738 = (inp[13]) ? 4'b0110 : 4'b0111;
																assign node46741 = (inp[13]) ? 4'b0111 : 4'b0110;
												assign node46745 = (inp[0]) ? node46755 : node46746;
													assign node46746 = (inp[5]) ? node46748 : 4'b0111;
														assign node46748 = (inp[13]) ? node46752 : node46749;
															assign node46749 = (inp[15]) ? 4'b0110 : 4'b0111;
															assign node46752 = (inp[15]) ? 4'b0111 : 4'b0110;
													assign node46755 = (inp[5]) ? node46757 : 4'b0110;
														assign node46757 = (inp[10]) ? node46765 : node46758;
															assign node46758 = (inp[13]) ? node46762 : node46759;
																assign node46759 = (inp[15]) ? 4'b0111 : 4'b0110;
																assign node46762 = (inp[15]) ? 4'b0110 : 4'b0111;
															assign node46765 = (inp[15]) ? node46769 : node46766;
																assign node46766 = (inp[13]) ? 4'b0111 : 4'b0110;
																assign node46769 = (inp[13]) ? 4'b0110 : 4'b0111;
										assign node46772 = (inp[1]) ? node46844 : node46773;
											assign node46773 = (inp[15]) ? node46805 : node46774;
												assign node46774 = (inp[5]) ? node46782 : node46775;
													assign node46775 = (inp[2]) ? node46779 : node46776;
														assign node46776 = (inp[0]) ? 4'b0111 : 4'b0110;
														assign node46779 = (inp[0]) ? 4'b0110 : 4'b0111;
													assign node46782 = (inp[0]) ? node46790 : node46783;
														assign node46783 = (inp[13]) ? node46787 : node46784;
															assign node46784 = (inp[2]) ? 4'b0111 : 4'b0110;
															assign node46787 = (inp[2]) ? 4'b0110 : 4'b0111;
														assign node46790 = (inp[10]) ? node46798 : node46791;
															assign node46791 = (inp[2]) ? node46795 : node46792;
																assign node46792 = (inp[13]) ? 4'b0110 : 4'b0111;
																assign node46795 = (inp[13]) ? 4'b0111 : 4'b0110;
															assign node46798 = (inp[2]) ? node46802 : node46799;
																assign node46799 = (inp[13]) ? 4'b0110 : 4'b0111;
																assign node46802 = (inp[13]) ? 4'b0111 : 4'b0110;
												assign node46805 = (inp[10]) ? node46829 : node46806;
													assign node46806 = (inp[0]) ? node46818 : node46807;
														assign node46807 = (inp[2]) ? node46813 : node46808;
															assign node46808 = (inp[5]) ? 4'b0110 : node46809;
																assign node46809 = (inp[13]) ? 4'b0111 : 4'b0110;
															assign node46813 = (inp[13]) ? node46815 : 4'b0111;
																assign node46815 = (inp[5]) ? 4'b0111 : 4'b0110;
														assign node46818 = (inp[2]) ? node46824 : node46819;
															assign node46819 = (inp[5]) ? 4'b0111 : node46820;
																assign node46820 = (inp[13]) ? 4'b0110 : 4'b0111;
															assign node46824 = (inp[5]) ? 4'b0110 : node46825;
																assign node46825 = (inp[13]) ? 4'b0111 : 4'b0110;
													assign node46829 = (inp[2]) ? node46837 : node46830;
														assign node46830 = (inp[0]) ? node46832 : 4'b0110;
															assign node46832 = (inp[5]) ? 4'b0111 : node46833;
																assign node46833 = (inp[13]) ? 4'b0110 : 4'b0111;
														assign node46837 = (inp[0]) ? 4'b0110 : node46838;
															assign node46838 = (inp[13]) ? node46840 : 4'b0111;
																assign node46840 = (inp[5]) ? 4'b0111 : 4'b0110;
											assign node46844 = (inp[10]) ? node46888 : node46845;
												assign node46845 = (inp[13]) ? node46869 : node46846;
													assign node46846 = (inp[5]) ? node46862 : node46847;
														assign node46847 = (inp[15]) ? node46855 : node46848;
															assign node46848 = (inp[2]) ? node46852 : node46849;
																assign node46849 = (inp[0]) ? 4'b0010 : 4'b0011;
																assign node46852 = (inp[0]) ? 4'b0011 : 4'b0010;
															assign node46855 = (inp[0]) ? node46859 : node46856;
																assign node46856 = (inp[2]) ? 4'b0011 : 4'b0010;
																assign node46859 = (inp[2]) ? 4'b0010 : 4'b0011;
														assign node46862 = (inp[0]) ? node46866 : node46863;
															assign node46863 = (inp[2]) ? 4'b0011 : 4'b0010;
															assign node46866 = (inp[2]) ? 4'b0010 : 4'b0011;
													assign node46869 = (inp[2]) ? node46877 : node46870;
														assign node46870 = (inp[0]) ? node46872 : 4'b0010;
															assign node46872 = (inp[15]) ? node46874 : 4'b0011;
																assign node46874 = (inp[5]) ? 4'b0011 : 4'b0010;
														assign node46877 = (inp[0]) ? node46883 : node46878;
															assign node46878 = (inp[15]) ? node46880 : 4'b0011;
																assign node46880 = (inp[5]) ? 4'b0011 : 4'b0010;
															assign node46883 = (inp[5]) ? 4'b0010 : node46884;
																assign node46884 = (inp[15]) ? 4'b0011 : 4'b0010;
												assign node46888 = (inp[2]) ? node46906 : node46889;
													assign node46889 = (inp[0]) ? node46897 : node46890;
														assign node46890 = (inp[5]) ? 4'b0010 : node46891;
															assign node46891 = (inp[15]) ? node46893 : 4'b0011;
																assign node46893 = (inp[13]) ? 4'b0011 : 4'b0010;
														assign node46897 = (inp[5]) ? 4'b0011 : node46898;
															assign node46898 = (inp[15]) ? node46902 : node46899;
																assign node46899 = (inp[13]) ? 4'b0011 : 4'b0010;
																assign node46902 = (inp[13]) ? 4'b0010 : 4'b0011;
													assign node46906 = (inp[0]) ? node46916 : node46907;
														assign node46907 = (inp[5]) ? 4'b0011 : node46908;
															assign node46908 = (inp[13]) ? node46912 : node46909;
																assign node46909 = (inp[15]) ? 4'b0011 : 4'b0010;
																assign node46912 = (inp[15]) ? 4'b0010 : 4'b0011;
														assign node46916 = (inp[5]) ? 4'b0010 : node46917;
															assign node46917 = (inp[13]) ? node46921 : node46918;
																assign node46918 = (inp[15]) ? 4'b0010 : 4'b0011;
																assign node46921 = (inp[15]) ? 4'b0011 : 4'b0010;
								assign node46925 = (inp[9]) ? node47195 : node46926;
									assign node46926 = (inp[15]) ? node47038 : node46927;
										assign node46927 = (inp[12]) ? node46975 : node46928;
											assign node46928 = (inp[1]) ? node46952 : node46929;
												assign node46929 = (inp[2]) ? node46941 : node46930;
													assign node46930 = (inp[0]) ? node46936 : node46931;
														assign node46931 = (inp[5]) ? node46933 : 4'b0010;
															assign node46933 = (inp[13]) ? 4'b0011 : 4'b0010;
														assign node46936 = (inp[5]) ? node46938 : 4'b0011;
															assign node46938 = (inp[13]) ? 4'b0010 : 4'b0011;
													assign node46941 = (inp[0]) ? node46947 : node46942;
														assign node46942 = (inp[13]) ? node46944 : 4'b0011;
															assign node46944 = (inp[5]) ? 4'b0010 : 4'b0011;
														assign node46947 = (inp[13]) ? node46949 : 4'b0010;
															assign node46949 = (inp[5]) ? 4'b0011 : 4'b0010;
												assign node46952 = (inp[13]) ? node46960 : node46953;
													assign node46953 = (inp[2]) ? node46957 : node46954;
														assign node46954 = (inp[0]) ? 4'b0111 : 4'b0110;
														assign node46957 = (inp[0]) ? 4'b0110 : 4'b0111;
													assign node46960 = (inp[0]) ? node46968 : node46961;
														assign node46961 = (inp[5]) ? node46965 : node46962;
															assign node46962 = (inp[2]) ? 4'b0111 : 4'b0110;
															assign node46965 = (inp[2]) ? 4'b0110 : 4'b0111;
														assign node46968 = (inp[2]) ? node46972 : node46969;
															assign node46969 = (inp[5]) ? 4'b0110 : 4'b0111;
															assign node46972 = (inp[5]) ? 4'b0111 : 4'b0110;
											assign node46975 = (inp[1]) ? node47015 : node46976;
												assign node46976 = (inp[10]) ? node46994 : node46977;
													assign node46977 = (inp[2]) ? node46983 : node46978;
														assign node46978 = (inp[0]) ? node46980 : 4'b0110;
															assign node46980 = (inp[5]) ? 4'b0110 : 4'b0111;
														assign node46983 = (inp[0]) ? node46989 : node46984;
															assign node46984 = (inp[5]) ? node46986 : 4'b0111;
																assign node46986 = (inp[13]) ? 4'b0110 : 4'b0111;
															assign node46989 = (inp[13]) ? node46991 : 4'b0110;
																assign node46991 = (inp[5]) ? 4'b0111 : 4'b0110;
													assign node46994 = (inp[13]) ? node47002 : node46995;
														assign node46995 = (inp[2]) ? node46999 : node46996;
															assign node46996 = (inp[0]) ? 4'b0111 : 4'b0110;
															assign node46999 = (inp[0]) ? 4'b0110 : 4'b0111;
														assign node47002 = (inp[5]) ? node47010 : node47003;
															assign node47003 = (inp[2]) ? node47007 : node47004;
																assign node47004 = (inp[0]) ? 4'b0111 : 4'b0110;
																assign node47007 = (inp[0]) ? 4'b0110 : 4'b0111;
															assign node47010 = (inp[0]) ? 4'b0111 : node47011;
																assign node47011 = (inp[2]) ? 4'b0110 : 4'b0111;
												assign node47015 = (inp[0]) ? node47027 : node47016;
													assign node47016 = (inp[2]) ? node47022 : node47017;
														assign node47017 = (inp[13]) ? 4'b0010 : node47018;
															assign node47018 = (inp[5]) ? 4'b0010 : 4'b0011;
														assign node47022 = (inp[5]) ? 4'b0011 : node47023;
															assign node47023 = (inp[13]) ? 4'b0011 : 4'b0010;
													assign node47027 = (inp[2]) ? node47033 : node47028;
														assign node47028 = (inp[13]) ? 4'b0011 : node47029;
															assign node47029 = (inp[5]) ? 4'b0011 : 4'b0010;
														assign node47033 = (inp[5]) ? 4'b0010 : node47034;
															assign node47034 = (inp[13]) ? 4'b0010 : 4'b0011;
										assign node47038 = (inp[5]) ? node47100 : node47039;
											assign node47039 = (inp[0]) ? node47069 : node47040;
												assign node47040 = (inp[2]) ? node47054 : node47041;
													assign node47041 = (inp[13]) ? node47049 : node47042;
														assign node47042 = (inp[1]) ? node47046 : node47043;
															assign node47043 = (inp[12]) ? 4'b0110 : 4'b0010;
															assign node47046 = (inp[10]) ? 4'b0010 : 4'b0110;
														assign node47049 = (inp[1]) ? 4'b0011 : node47050;
															assign node47050 = (inp[12]) ? 4'b0111 : 4'b0011;
													assign node47054 = (inp[13]) ? node47062 : node47055;
														assign node47055 = (inp[12]) ? node47059 : node47056;
															assign node47056 = (inp[1]) ? 4'b0111 : 4'b0011;
															assign node47059 = (inp[1]) ? 4'b0011 : 4'b0111;
														assign node47062 = (inp[12]) ? node47066 : node47063;
															assign node47063 = (inp[1]) ? 4'b0111 : 4'b0010;
															assign node47066 = (inp[1]) ? 4'b0010 : 4'b0110;
												assign node47069 = (inp[2]) ? node47085 : node47070;
													assign node47070 = (inp[13]) ? node47078 : node47071;
														assign node47071 = (inp[1]) ? node47075 : node47072;
															assign node47072 = (inp[12]) ? 4'b0111 : 4'b0011;
															assign node47075 = (inp[12]) ? 4'b0011 : 4'b0111;
														assign node47078 = (inp[12]) ? node47082 : node47079;
															assign node47079 = (inp[1]) ? 4'b0111 : 4'b0010;
															assign node47082 = (inp[1]) ? 4'b0010 : 4'b0110;
													assign node47085 = (inp[13]) ? node47091 : node47086;
														assign node47086 = (inp[12]) ? 4'b0010 : node47087;
															assign node47087 = (inp[1]) ? 4'b0110 : 4'b0010;
														assign node47091 = (inp[10]) ? 4'b0011 : node47092;
															assign node47092 = (inp[1]) ? node47096 : node47093;
																assign node47093 = (inp[12]) ? 4'b0111 : 4'b0011;
																assign node47096 = (inp[12]) ? 4'b0011 : 4'b0110;
											assign node47100 = (inp[10]) ? node47148 : node47101;
												assign node47101 = (inp[0]) ? node47119 : node47102;
													assign node47102 = (inp[2]) ? node47110 : node47103;
														assign node47103 = (inp[1]) ? node47107 : node47104;
															assign node47104 = (inp[12]) ? 4'b0110 : 4'b0010;
															assign node47107 = (inp[12]) ? 4'b0010 : 4'b0110;
														assign node47110 = (inp[13]) ? 4'b0011 : node47111;
															assign node47111 = (inp[12]) ? node47115 : node47112;
																assign node47112 = (inp[1]) ? 4'b0110 : 4'b0011;
																assign node47115 = (inp[1]) ? 4'b0011 : 4'b0111;
													assign node47119 = (inp[2]) ? node47133 : node47120;
														assign node47120 = (inp[13]) ? node47126 : node47121;
															assign node47121 = (inp[12]) ? 4'b0011 : node47122;
																assign node47122 = (inp[1]) ? 4'b0110 : 4'b0011;
															assign node47126 = (inp[1]) ? node47130 : node47127;
																assign node47127 = (inp[12]) ? 4'b0111 : 4'b0011;
																assign node47130 = (inp[12]) ? 4'b0011 : 4'b0111;
														assign node47133 = (inp[13]) ? node47141 : node47134;
															assign node47134 = (inp[1]) ? node47138 : node47135;
																assign node47135 = (inp[12]) ? 4'b0110 : 4'b0010;
																assign node47138 = (inp[12]) ? 4'b0010 : 4'b0111;
															assign node47141 = (inp[12]) ? node47145 : node47142;
																assign node47142 = (inp[1]) ? 4'b0110 : 4'b0010;
																assign node47145 = (inp[1]) ? 4'b0010 : 4'b0110;
												assign node47148 = (inp[2]) ? node47176 : node47149;
													assign node47149 = (inp[0]) ? node47163 : node47150;
														assign node47150 = (inp[13]) ? node47156 : node47151;
															assign node47151 = (inp[1]) ? 4'b0010 : node47152;
																assign node47152 = (inp[12]) ? 4'b0110 : 4'b0010;
															assign node47156 = (inp[1]) ? node47160 : node47157;
																assign node47157 = (inp[12]) ? 4'b0110 : 4'b0010;
																assign node47160 = (inp[12]) ? 4'b0010 : 4'b0110;
														assign node47163 = (inp[13]) ? node47169 : node47164;
															assign node47164 = (inp[1]) ? 4'b0011 : node47165;
																assign node47165 = (inp[12]) ? 4'b0111 : 4'b0011;
															assign node47169 = (inp[1]) ? node47173 : node47170;
																assign node47170 = (inp[12]) ? 4'b0111 : 4'b0011;
																assign node47173 = (inp[12]) ? 4'b0011 : 4'b0111;
													assign node47176 = (inp[0]) ? node47186 : node47177;
														assign node47177 = (inp[12]) ? node47183 : node47178;
															assign node47178 = (inp[1]) ? node47180 : 4'b0011;
																assign node47180 = (inp[13]) ? 4'b0111 : 4'b0110;
															assign node47183 = (inp[1]) ? 4'b0011 : 4'b0111;
														assign node47186 = (inp[12]) ? node47192 : node47187;
															assign node47187 = (inp[1]) ? node47189 : 4'b0010;
																assign node47189 = (inp[13]) ? 4'b0110 : 4'b0111;
															assign node47192 = (inp[1]) ? 4'b0010 : 4'b0110;
									assign node47195 = (inp[13]) ? node47397 : node47196;
										assign node47196 = (inp[10]) ? node47302 : node47197;
											assign node47197 = (inp[15]) ? node47249 : node47198;
												assign node47198 = (inp[5]) ? node47222 : node47199;
													assign node47199 = (inp[1]) ? node47215 : node47200;
														assign node47200 = (inp[12]) ? node47208 : node47201;
															assign node47201 = (inp[2]) ? node47205 : node47202;
																assign node47202 = (inp[0]) ? 4'b0011 : 4'b0010;
																assign node47205 = (inp[0]) ? 4'b0010 : 4'b0011;
															assign node47208 = (inp[0]) ? node47212 : node47209;
																assign node47209 = (inp[2]) ? 4'b0111 : 4'b0110;
																assign node47212 = (inp[2]) ? 4'b0110 : 4'b0111;
														assign node47215 = (inp[12]) ? node47217 : 4'b0111;
															assign node47217 = (inp[0]) ? node47219 : 4'b0011;
																assign node47219 = (inp[2]) ? 4'b0011 : 4'b0010;
													assign node47222 = (inp[0]) ? node47234 : node47223;
														assign node47223 = (inp[2]) ? node47229 : node47224;
															assign node47224 = (inp[1]) ? node47226 : 4'b0010;
																assign node47226 = (inp[12]) ? 4'b0010 : 4'b0110;
															assign node47229 = (inp[12]) ? node47231 : 4'b0011;
																assign node47231 = (inp[1]) ? 4'b0011 : 4'b0111;
														assign node47234 = (inp[2]) ? node47242 : node47235;
															assign node47235 = (inp[12]) ? node47239 : node47236;
																assign node47236 = (inp[1]) ? 4'b0111 : 4'b0011;
																assign node47239 = (inp[1]) ? 4'b0011 : 4'b0111;
															assign node47242 = (inp[12]) ? node47246 : node47243;
																assign node47243 = (inp[1]) ? 4'b0110 : 4'b0010;
																assign node47246 = (inp[1]) ? 4'b0010 : 4'b0110;
												assign node47249 = (inp[12]) ? node47273 : node47250;
													assign node47250 = (inp[1]) ? node47258 : node47251;
														assign node47251 = (inp[5]) ? node47253 : 4'b0011;
															assign node47253 = (inp[0]) ? 4'b0010 : node47254;
																assign node47254 = (inp[2]) ? 4'b0011 : 4'b0010;
														assign node47258 = (inp[0]) ? node47266 : node47259;
															assign node47259 = (inp[5]) ? node47263 : node47260;
																assign node47260 = (inp[2]) ? 4'b0111 : 4'b0110;
																assign node47263 = (inp[2]) ? 4'b0110 : 4'b0111;
															assign node47266 = (inp[2]) ? node47270 : node47267;
																assign node47267 = (inp[5]) ? 4'b0110 : 4'b0111;
																assign node47270 = (inp[5]) ? 4'b0111 : 4'b0110;
													assign node47273 = (inp[1]) ? node47287 : node47274;
														assign node47274 = (inp[5]) ? node47280 : node47275;
															assign node47275 = (inp[2]) ? 4'b0110 : node47276;
																assign node47276 = (inp[0]) ? 4'b0111 : 4'b0110;
															assign node47280 = (inp[2]) ? node47284 : node47281;
																assign node47281 = (inp[0]) ? 4'b0111 : 4'b0110;
																assign node47284 = (inp[0]) ? 4'b0110 : 4'b0111;
														assign node47287 = (inp[5]) ? node47295 : node47288;
															assign node47288 = (inp[2]) ? node47292 : node47289;
																assign node47289 = (inp[0]) ? 4'b0011 : 4'b0010;
																assign node47292 = (inp[0]) ? 4'b0010 : 4'b0011;
															assign node47295 = (inp[0]) ? node47299 : node47296;
																assign node47296 = (inp[2]) ? 4'b0011 : 4'b0010;
																assign node47299 = (inp[2]) ? 4'b0010 : 4'b0011;
											assign node47302 = (inp[12]) ? node47362 : node47303;
												assign node47303 = (inp[1]) ? node47331 : node47304;
													assign node47304 = (inp[15]) ? node47320 : node47305;
														assign node47305 = (inp[5]) ? node47313 : node47306;
															assign node47306 = (inp[2]) ? node47310 : node47307;
																assign node47307 = (inp[0]) ? 4'b0011 : 4'b0010;
																assign node47310 = (inp[0]) ? 4'b0010 : 4'b0011;
															assign node47313 = (inp[2]) ? node47317 : node47314;
																assign node47314 = (inp[0]) ? 4'b0011 : 4'b0010;
																assign node47317 = (inp[0]) ? 4'b0010 : 4'b0011;
														assign node47320 = (inp[5]) ? node47326 : node47321;
															assign node47321 = (inp[0]) ? 4'b0010 : node47322;
																assign node47322 = (inp[2]) ? 4'b0011 : 4'b0010;
															assign node47326 = (inp[0]) ? node47328 : 4'b0010;
																assign node47328 = (inp[2]) ? 4'b0010 : 4'b0011;
													assign node47331 = (inp[15]) ? node47347 : node47332;
														assign node47332 = (inp[5]) ? node47340 : node47333;
															assign node47333 = (inp[0]) ? node47337 : node47334;
																assign node47334 = (inp[2]) ? 4'b0111 : 4'b0110;
																assign node47337 = (inp[2]) ? 4'b0110 : 4'b0111;
															assign node47340 = (inp[0]) ? node47344 : node47341;
																assign node47341 = (inp[2]) ? 4'b0111 : 4'b0110;
																assign node47344 = (inp[2]) ? 4'b0110 : 4'b0111;
														assign node47347 = (inp[2]) ? node47355 : node47348;
															assign node47348 = (inp[5]) ? node47352 : node47349;
																assign node47349 = (inp[0]) ? 4'b0111 : 4'b0110;
																assign node47352 = (inp[0]) ? 4'b0110 : 4'b0111;
															assign node47355 = (inp[5]) ? node47359 : node47356;
																assign node47356 = (inp[0]) ? 4'b0110 : 4'b0111;
																assign node47359 = (inp[0]) ? 4'b0111 : 4'b0110;
												assign node47362 = (inp[1]) ? node47378 : node47363;
													assign node47363 = (inp[5]) ? node47371 : node47364;
														assign node47364 = (inp[0]) ? node47368 : node47365;
															assign node47365 = (inp[2]) ? 4'b0111 : 4'b0110;
															assign node47368 = (inp[2]) ? 4'b0110 : 4'b0111;
														assign node47371 = (inp[2]) ? node47375 : node47372;
															assign node47372 = (inp[0]) ? 4'b0111 : 4'b0110;
															assign node47375 = (inp[0]) ? 4'b0110 : 4'b0111;
													assign node47378 = (inp[15]) ? node47388 : node47379;
														assign node47379 = (inp[5]) ? node47381 : 4'b0010;
															assign node47381 = (inp[0]) ? node47385 : node47382;
																assign node47382 = (inp[2]) ? 4'b0011 : 4'b0010;
																assign node47385 = (inp[2]) ? 4'b0010 : 4'b0011;
														assign node47388 = (inp[5]) ? 4'b0011 : node47389;
															assign node47389 = (inp[2]) ? node47393 : node47390;
																assign node47390 = (inp[0]) ? 4'b0011 : 4'b0010;
																assign node47393 = (inp[0]) ? 4'b0010 : 4'b0011;
										assign node47397 = (inp[5]) ? node47455 : node47398;
											assign node47398 = (inp[0]) ? node47428 : node47399;
												assign node47399 = (inp[2]) ? node47413 : node47400;
													assign node47400 = (inp[15]) ? node47408 : node47401;
														assign node47401 = (inp[1]) ? node47405 : node47402;
															assign node47402 = (inp[12]) ? 4'b0110 : 4'b0010;
															assign node47405 = (inp[12]) ? 4'b0010 : 4'b0110;
														assign node47408 = (inp[12]) ? 4'b0011 : node47409;
															assign node47409 = (inp[1]) ? 4'b0110 : 4'b0011;
													assign node47413 = (inp[15]) ? node47421 : node47414;
														assign node47414 = (inp[12]) ? node47418 : node47415;
															assign node47415 = (inp[1]) ? 4'b0111 : 4'b0011;
															assign node47418 = (inp[1]) ? 4'b0011 : 4'b0111;
														assign node47421 = (inp[1]) ? node47425 : node47422;
															assign node47422 = (inp[12]) ? 4'b0110 : 4'b0010;
															assign node47425 = (inp[12]) ? 4'b0010 : 4'b0111;
												assign node47428 = (inp[2]) ? node47442 : node47429;
													assign node47429 = (inp[15]) ? node47435 : node47430;
														assign node47430 = (inp[1]) ? 4'b0111 : node47431;
															assign node47431 = (inp[12]) ? 4'b0111 : 4'b0011;
														assign node47435 = (inp[12]) ? node47439 : node47436;
															assign node47436 = (inp[1]) ? 4'b0111 : 4'b0010;
															assign node47439 = (inp[1]) ? 4'b0010 : 4'b0110;
													assign node47442 = (inp[15]) ? node47450 : node47443;
														assign node47443 = (inp[12]) ? node47447 : node47444;
															assign node47444 = (inp[1]) ? 4'b0110 : 4'b0010;
															assign node47447 = (inp[1]) ? 4'b0010 : 4'b0110;
														assign node47450 = (inp[12]) ? node47452 : 4'b0110;
															assign node47452 = (inp[1]) ? 4'b0011 : 4'b0111;
											assign node47455 = (inp[2]) ? node47487 : node47456;
												assign node47456 = (inp[0]) ? node47472 : node47457;
													assign node47457 = (inp[15]) ? node47465 : node47458;
														assign node47458 = (inp[12]) ? node47462 : node47459;
															assign node47459 = (inp[1]) ? 4'b0111 : 4'b0011;
															assign node47462 = (inp[1]) ? 4'b0010 : 4'b0111;
														assign node47465 = (inp[1]) ? node47469 : node47466;
															assign node47466 = (inp[12]) ? 4'b0110 : 4'b0010;
															assign node47469 = (inp[12]) ? 4'b0010 : 4'b0110;
													assign node47472 = (inp[15]) ? node47480 : node47473;
														assign node47473 = (inp[1]) ? node47477 : node47474;
															assign node47474 = (inp[12]) ? 4'b0110 : 4'b0010;
															assign node47477 = (inp[12]) ? 4'b0011 : 4'b0110;
														assign node47480 = (inp[1]) ? node47484 : node47481;
															assign node47481 = (inp[12]) ? 4'b0111 : 4'b0011;
															assign node47484 = (inp[12]) ? 4'b0011 : 4'b0111;
												assign node47487 = (inp[0]) ? node47503 : node47488;
													assign node47488 = (inp[15]) ? node47496 : node47489;
														assign node47489 = (inp[1]) ? node47493 : node47490;
															assign node47490 = (inp[12]) ? 4'b0110 : 4'b0010;
															assign node47493 = (inp[12]) ? 4'b0011 : 4'b0110;
														assign node47496 = (inp[12]) ? node47500 : node47497;
															assign node47497 = (inp[1]) ? 4'b0111 : 4'b0011;
															assign node47500 = (inp[1]) ? 4'b0011 : 4'b0111;
													assign node47503 = (inp[15]) ? node47511 : node47504;
														assign node47504 = (inp[12]) ? node47508 : node47505;
															assign node47505 = (inp[1]) ? 4'b0111 : 4'b0011;
															assign node47508 = (inp[1]) ? 4'b0010 : 4'b0111;
														assign node47511 = (inp[12]) ? node47515 : node47512;
															assign node47512 = (inp[1]) ? 4'b0110 : 4'b0010;
															assign node47515 = (inp[1]) ? 4'b0010 : 4'b0110;
						assign node47518 = (inp[13]) ? node48298 : node47519;
							assign node47519 = (inp[12]) ? node47957 : node47520;
								assign node47520 = (inp[8]) ? node47680 : node47521;
									assign node47521 = (inp[1]) ? node47633 : node47522;
										assign node47522 = (inp[15]) ? node47596 : node47523;
											assign node47523 = (inp[10]) ? node47547 : node47524;
												assign node47524 = (inp[9]) ? node47536 : node47525;
													assign node47525 = (inp[2]) ? node47531 : node47526;
														assign node47526 = (inp[0]) ? 4'b0010 : node47527;
															assign node47527 = (inp[5]) ? 4'b0011 : 4'b0010;
														assign node47531 = (inp[0]) ? 4'b0011 : node47532;
															assign node47532 = (inp[5]) ? 4'b0010 : 4'b0011;
													assign node47536 = (inp[2]) ? node47542 : node47537;
														assign node47537 = (inp[5]) ? node47539 : 4'b0011;
															assign node47539 = (inp[0]) ? 4'b0011 : 4'b0010;
														assign node47542 = (inp[5]) ? node47544 : 4'b0010;
															assign node47544 = (inp[0]) ? 4'b0010 : 4'b0011;
												assign node47547 = (inp[0]) ? node47577 : node47548;
													assign node47548 = (inp[11]) ? node47564 : node47549;
														assign node47549 = (inp[2]) ? node47557 : node47550;
															assign node47550 = (inp[9]) ? node47554 : node47551;
																assign node47551 = (inp[5]) ? 4'b0011 : 4'b0010;
																assign node47554 = (inp[5]) ? 4'b0010 : 4'b0011;
															assign node47557 = (inp[5]) ? node47561 : node47558;
																assign node47558 = (inp[9]) ? 4'b0010 : 4'b0011;
																assign node47561 = (inp[9]) ? 4'b0011 : 4'b0010;
														assign node47564 = (inp[5]) ? node47570 : node47565;
															assign node47565 = (inp[9]) ? node47567 : 4'b0011;
																assign node47567 = (inp[2]) ? 4'b0010 : 4'b0011;
															assign node47570 = (inp[9]) ? node47574 : node47571;
																assign node47571 = (inp[2]) ? 4'b0010 : 4'b0011;
																assign node47574 = (inp[2]) ? 4'b0011 : 4'b0010;
													assign node47577 = (inp[5]) ? node47589 : node47578;
														assign node47578 = (inp[11]) ? node47584 : node47579;
															assign node47579 = (inp[9]) ? 4'b0010 : node47580;
																assign node47580 = (inp[2]) ? 4'b0011 : 4'b0010;
															assign node47584 = (inp[2]) ? 4'b0010 : node47585;
																assign node47585 = (inp[9]) ? 4'b0011 : 4'b0010;
														assign node47589 = (inp[2]) ? node47593 : node47590;
															assign node47590 = (inp[9]) ? 4'b0011 : 4'b0010;
															assign node47593 = (inp[9]) ? 4'b0010 : 4'b0011;
											assign node47596 = (inp[5]) ? node47604 : node47597;
												assign node47597 = (inp[2]) ? node47601 : node47598;
													assign node47598 = (inp[9]) ? 4'b0111 : 4'b0110;
													assign node47601 = (inp[9]) ? 4'b0110 : 4'b0111;
												assign node47604 = (inp[9]) ? node47612 : node47605;
													assign node47605 = (inp[2]) ? node47609 : node47606;
														assign node47606 = (inp[0]) ? 4'b0110 : 4'b0111;
														assign node47609 = (inp[0]) ? 4'b0111 : 4'b0110;
													assign node47612 = (inp[10]) ? node47620 : node47613;
														assign node47613 = (inp[0]) ? node47617 : node47614;
															assign node47614 = (inp[2]) ? 4'b0111 : 4'b0110;
															assign node47617 = (inp[2]) ? 4'b0110 : 4'b0111;
														assign node47620 = (inp[11]) ? node47626 : node47621;
															assign node47621 = (inp[2]) ? 4'b0110 : node47622;
																assign node47622 = (inp[0]) ? 4'b0111 : 4'b0110;
															assign node47626 = (inp[2]) ? node47630 : node47627;
																assign node47627 = (inp[0]) ? 4'b0111 : 4'b0110;
																assign node47630 = (inp[0]) ? 4'b0110 : 4'b0111;
										assign node47633 = (inp[9]) ? node47657 : node47634;
											assign node47634 = (inp[15]) ? node47646 : node47635;
												assign node47635 = (inp[2]) ? node47641 : node47636;
													assign node47636 = (inp[5]) ? node47638 : 4'b0010;
														assign node47638 = (inp[0]) ? 4'b0010 : 4'b0011;
													assign node47641 = (inp[0]) ? 4'b0011 : node47642;
														assign node47642 = (inp[5]) ? 4'b0010 : 4'b0011;
												assign node47646 = (inp[2]) ? node47652 : node47647;
													assign node47647 = (inp[5]) ? node47649 : 4'b0011;
														assign node47649 = (inp[0]) ? 4'b0011 : 4'b0010;
													assign node47652 = (inp[5]) ? node47654 : 4'b0010;
														assign node47654 = (inp[0]) ? 4'b0010 : 4'b0011;
											assign node47657 = (inp[15]) ? node47669 : node47658;
												assign node47658 = (inp[2]) ? node47664 : node47659;
													assign node47659 = (inp[0]) ? 4'b0011 : node47660;
														assign node47660 = (inp[5]) ? 4'b0010 : 4'b0011;
													assign node47664 = (inp[5]) ? node47666 : 4'b0010;
														assign node47666 = (inp[0]) ? 4'b0010 : 4'b0011;
												assign node47669 = (inp[2]) ? node47675 : node47670;
													assign node47670 = (inp[5]) ? node47672 : 4'b0010;
														assign node47672 = (inp[0]) ? 4'b0010 : 4'b0011;
													assign node47675 = (inp[0]) ? 4'b0011 : node47676;
														assign node47676 = (inp[5]) ? 4'b0010 : 4'b0011;
									assign node47680 = (inp[1]) ? node47758 : node47681;
										assign node47681 = (inp[9]) ? node47735 : node47682;
											assign node47682 = (inp[11]) ? node47706 : node47683;
												assign node47683 = (inp[2]) ? node47695 : node47684;
													assign node47684 = (inp[0]) ? node47690 : node47685;
														assign node47685 = (inp[15]) ? 4'b0010 : node47686;
															assign node47686 = (inp[5]) ? 4'b0011 : 4'b0010;
														assign node47690 = (inp[15]) ? 4'b0011 : node47691;
															assign node47691 = (inp[5]) ? 4'b0010 : 4'b0011;
													assign node47695 = (inp[0]) ? node47701 : node47696;
														assign node47696 = (inp[5]) ? node47698 : 4'b0011;
															assign node47698 = (inp[15]) ? 4'b0011 : 4'b0010;
														assign node47701 = (inp[5]) ? node47703 : 4'b0010;
															assign node47703 = (inp[15]) ? 4'b0010 : 4'b0011;
												assign node47706 = (inp[5]) ? node47722 : node47707;
													assign node47707 = (inp[15]) ? node47715 : node47708;
														assign node47708 = (inp[2]) ? node47712 : node47709;
															assign node47709 = (inp[0]) ? 4'b0011 : 4'b0010;
															assign node47712 = (inp[0]) ? 4'b0010 : 4'b0011;
														assign node47715 = (inp[2]) ? node47719 : node47716;
															assign node47716 = (inp[0]) ? 4'b0011 : 4'b0010;
															assign node47719 = (inp[0]) ? 4'b0010 : 4'b0011;
													assign node47722 = (inp[15]) ? node47730 : node47723;
														assign node47723 = (inp[2]) ? node47727 : node47724;
															assign node47724 = (inp[0]) ? 4'b0010 : 4'b0011;
															assign node47727 = (inp[0]) ? 4'b0011 : 4'b0010;
														assign node47730 = (inp[2]) ? node47732 : 4'b0010;
															assign node47732 = (inp[0]) ? 4'b0010 : 4'b0011;
											assign node47735 = (inp[2]) ? node47747 : node47736;
												assign node47736 = (inp[0]) ? node47742 : node47737;
													assign node47737 = (inp[5]) ? node47739 : 4'b0010;
														assign node47739 = (inp[15]) ? 4'b0010 : 4'b0011;
													assign node47742 = (inp[15]) ? 4'b0011 : node47743;
														assign node47743 = (inp[5]) ? 4'b0010 : 4'b0011;
												assign node47747 = (inp[0]) ? node47753 : node47748;
													assign node47748 = (inp[15]) ? 4'b0011 : node47749;
														assign node47749 = (inp[5]) ? 4'b0010 : 4'b0011;
													assign node47753 = (inp[5]) ? node47755 : 4'b0010;
														assign node47755 = (inp[15]) ? 4'b0010 : 4'b0011;
										assign node47758 = (inp[10]) ? node47860 : node47759;
											assign node47759 = (inp[11]) ? node47803 : node47760;
												assign node47760 = (inp[5]) ? node47790 : node47761;
													assign node47761 = (inp[9]) ? node47777 : node47762;
														assign node47762 = (inp[2]) ? node47770 : node47763;
															assign node47763 = (inp[15]) ? node47767 : node47764;
																assign node47764 = (inp[0]) ? 4'b0111 : 4'b0110;
																assign node47767 = (inp[0]) ? 4'b0110 : 4'b0111;
															assign node47770 = (inp[0]) ? node47774 : node47771;
																assign node47771 = (inp[15]) ? 4'b0110 : 4'b0111;
																assign node47774 = (inp[15]) ? 4'b0111 : 4'b0110;
														assign node47777 = (inp[2]) ? node47783 : node47778;
															assign node47778 = (inp[15]) ? 4'b0110 : node47779;
																assign node47779 = (inp[0]) ? 4'b0111 : 4'b0110;
															assign node47783 = (inp[0]) ? node47787 : node47784;
																assign node47784 = (inp[15]) ? 4'b0110 : 4'b0111;
																assign node47787 = (inp[15]) ? 4'b0111 : 4'b0110;
													assign node47790 = (inp[0]) ? node47798 : node47791;
														assign node47791 = (inp[2]) ? node47795 : node47792;
															assign node47792 = (inp[15]) ? 4'b0110 : 4'b0111;
															assign node47795 = (inp[15]) ? 4'b0111 : 4'b0110;
														assign node47798 = (inp[15]) ? node47800 : 4'b0110;
															assign node47800 = (inp[2]) ? 4'b0110 : 4'b0111;
												assign node47803 = (inp[5]) ? node47829 : node47804;
													assign node47804 = (inp[15]) ? node47820 : node47805;
														assign node47805 = (inp[9]) ? node47813 : node47806;
															assign node47806 = (inp[0]) ? node47810 : node47807;
																assign node47807 = (inp[2]) ? 4'b0111 : 4'b0110;
																assign node47810 = (inp[2]) ? 4'b0110 : 4'b0111;
															assign node47813 = (inp[0]) ? node47817 : node47814;
																assign node47814 = (inp[2]) ? 4'b0111 : 4'b0110;
																assign node47817 = (inp[2]) ? 4'b0110 : 4'b0111;
														assign node47820 = (inp[9]) ? node47826 : node47821;
															assign node47821 = (inp[2]) ? node47823 : 4'b0111;
																assign node47823 = (inp[0]) ? 4'b0111 : 4'b0110;
															assign node47826 = (inp[0]) ? 4'b0110 : 4'b0111;
													assign node47829 = (inp[9]) ? node47845 : node47830;
														assign node47830 = (inp[0]) ? node47838 : node47831;
															assign node47831 = (inp[15]) ? node47835 : node47832;
																assign node47832 = (inp[2]) ? 4'b0110 : 4'b0111;
																assign node47835 = (inp[2]) ? 4'b0111 : 4'b0110;
															assign node47838 = (inp[2]) ? node47842 : node47839;
																assign node47839 = (inp[15]) ? 4'b0111 : 4'b0110;
																assign node47842 = (inp[15]) ? 4'b0110 : 4'b0111;
														assign node47845 = (inp[0]) ? node47853 : node47846;
															assign node47846 = (inp[2]) ? node47850 : node47847;
																assign node47847 = (inp[15]) ? 4'b0110 : 4'b0111;
																assign node47850 = (inp[15]) ? 4'b0111 : 4'b0110;
															assign node47853 = (inp[15]) ? node47857 : node47854;
																assign node47854 = (inp[2]) ? 4'b0111 : 4'b0110;
																assign node47857 = (inp[2]) ? 4'b0110 : 4'b0111;
											assign node47860 = (inp[11]) ? node47910 : node47861;
												assign node47861 = (inp[9]) ? node47887 : node47862;
													assign node47862 = (inp[15]) ? node47878 : node47863;
														assign node47863 = (inp[0]) ? node47871 : node47864;
															assign node47864 = (inp[5]) ? node47868 : node47865;
																assign node47865 = (inp[2]) ? 4'b0111 : 4'b0110;
																assign node47868 = (inp[2]) ? 4'b0110 : 4'b0111;
															assign node47871 = (inp[2]) ? node47875 : node47872;
																assign node47872 = (inp[5]) ? 4'b0110 : 4'b0111;
																assign node47875 = (inp[5]) ? 4'b0111 : 4'b0110;
														assign node47878 = (inp[5]) ? node47880 : 4'b0111;
															assign node47880 = (inp[2]) ? node47884 : node47881;
																assign node47881 = (inp[0]) ? 4'b0111 : 4'b0110;
																assign node47884 = (inp[0]) ? 4'b0110 : 4'b0111;
													assign node47887 = (inp[0]) ? node47897 : node47888;
														assign node47888 = (inp[15]) ? node47890 : 4'b0111;
															assign node47890 = (inp[2]) ? node47894 : node47891;
																assign node47891 = (inp[5]) ? 4'b0110 : 4'b0111;
																assign node47894 = (inp[5]) ? 4'b0111 : 4'b0110;
														assign node47897 = (inp[15]) ? node47905 : node47898;
															assign node47898 = (inp[2]) ? node47902 : node47899;
																assign node47899 = (inp[5]) ? 4'b0110 : 4'b0111;
																assign node47902 = (inp[5]) ? 4'b0111 : 4'b0110;
															assign node47905 = (inp[5]) ? 4'b0111 : node47906;
																assign node47906 = (inp[2]) ? 4'b0111 : 4'b0110;
												assign node47910 = (inp[5]) ? node47926 : node47911;
													assign node47911 = (inp[0]) ? node47919 : node47912;
														assign node47912 = (inp[2]) ? node47916 : node47913;
															assign node47913 = (inp[15]) ? 4'b0111 : 4'b0110;
															assign node47916 = (inp[15]) ? 4'b0110 : 4'b0111;
														assign node47919 = (inp[2]) ? node47923 : node47920;
															assign node47920 = (inp[15]) ? 4'b0110 : 4'b0111;
															assign node47923 = (inp[15]) ? 4'b0111 : 4'b0110;
													assign node47926 = (inp[9]) ? node47942 : node47927;
														assign node47927 = (inp[0]) ? node47935 : node47928;
															assign node47928 = (inp[15]) ? node47932 : node47929;
																assign node47929 = (inp[2]) ? 4'b0110 : 4'b0111;
																assign node47932 = (inp[2]) ? 4'b0111 : 4'b0110;
															assign node47935 = (inp[15]) ? node47939 : node47936;
																assign node47936 = (inp[2]) ? 4'b0111 : 4'b0110;
																assign node47939 = (inp[2]) ? 4'b0110 : 4'b0111;
														assign node47942 = (inp[0]) ? node47950 : node47943;
															assign node47943 = (inp[2]) ? node47947 : node47944;
																assign node47944 = (inp[15]) ? 4'b0110 : 4'b0111;
																assign node47947 = (inp[15]) ? 4'b0111 : 4'b0110;
															assign node47950 = (inp[15]) ? node47954 : node47951;
																assign node47951 = (inp[2]) ? 4'b0111 : 4'b0110;
																assign node47954 = (inp[2]) ? 4'b0110 : 4'b0111;
								assign node47957 = (inp[15]) ? node48143 : node47958;
									assign node47958 = (inp[8]) ? node48064 : node47959;
										assign node47959 = (inp[5]) ? node48021 : node47960;
											assign node47960 = (inp[0]) ? node47984 : node47961;
												assign node47961 = (inp[1]) ? node47969 : node47962;
													assign node47962 = (inp[2]) ? node47966 : node47963;
														assign node47963 = (inp[9]) ? 4'b0111 : 4'b0110;
														assign node47966 = (inp[9]) ? 4'b0110 : 4'b0111;
													assign node47969 = (inp[11]) ? node47977 : node47970;
														assign node47970 = (inp[2]) ? node47974 : node47971;
															assign node47971 = (inp[9]) ? 4'b0110 : 4'b0111;
															assign node47974 = (inp[9]) ? 4'b0111 : 4'b0110;
														assign node47977 = (inp[9]) ? node47981 : node47978;
															assign node47978 = (inp[2]) ? 4'b0110 : 4'b0111;
															assign node47981 = (inp[2]) ? 4'b0111 : 4'b0110;
												assign node47984 = (inp[10]) ? node48000 : node47985;
													assign node47985 = (inp[2]) ? node47993 : node47986;
														assign node47986 = (inp[1]) ? node47990 : node47987;
															assign node47987 = (inp[9]) ? 4'b0110 : 4'b0111;
															assign node47990 = (inp[9]) ? 4'b0111 : 4'b0110;
														assign node47993 = (inp[9]) ? node47997 : node47994;
															assign node47994 = (inp[1]) ? 4'b0111 : 4'b0110;
															assign node47997 = (inp[1]) ? 4'b0110 : 4'b0111;
													assign node48000 = (inp[9]) ? node48014 : node48001;
														assign node48001 = (inp[11]) ? node48009 : node48002;
															assign node48002 = (inp[2]) ? node48006 : node48003;
																assign node48003 = (inp[1]) ? 4'b0110 : 4'b0111;
																assign node48006 = (inp[1]) ? 4'b0111 : 4'b0110;
															assign node48009 = (inp[1]) ? node48011 : 4'b0110;
																assign node48011 = (inp[2]) ? 4'b0111 : 4'b0110;
														assign node48014 = (inp[1]) ? node48018 : node48015;
															assign node48015 = (inp[2]) ? 4'b0111 : 4'b0110;
															assign node48018 = (inp[2]) ? 4'b0110 : 4'b0111;
											assign node48021 = (inp[2]) ? node48057 : node48022;
												assign node48022 = (inp[11]) ? node48038 : node48023;
													assign node48023 = (inp[0]) ? node48031 : node48024;
														assign node48024 = (inp[9]) ? node48028 : node48025;
															assign node48025 = (inp[1]) ? 4'b0111 : 4'b0110;
															assign node48028 = (inp[1]) ? 4'b0110 : 4'b0111;
														assign node48031 = (inp[9]) ? node48035 : node48032;
															assign node48032 = (inp[1]) ? 4'b0111 : 4'b0110;
															assign node48035 = (inp[1]) ? 4'b0110 : 4'b0111;
													assign node48038 = (inp[10]) ? node48050 : node48039;
														assign node48039 = (inp[0]) ? node48045 : node48040;
															assign node48040 = (inp[1]) ? 4'b0111 : node48041;
																assign node48041 = (inp[9]) ? 4'b0111 : 4'b0110;
															assign node48045 = (inp[1]) ? node48047 : 4'b0111;
																assign node48047 = (inp[9]) ? 4'b0110 : 4'b0111;
														assign node48050 = (inp[9]) ? node48054 : node48051;
															assign node48051 = (inp[1]) ? 4'b0111 : 4'b0110;
															assign node48054 = (inp[1]) ? 4'b0110 : 4'b0111;
												assign node48057 = (inp[1]) ? node48061 : node48058;
													assign node48058 = (inp[9]) ? 4'b0110 : 4'b0111;
													assign node48061 = (inp[9]) ? 4'b0111 : 4'b0110;
										assign node48064 = (inp[1]) ? node48080 : node48065;
											assign node48065 = (inp[5]) ? node48073 : node48066;
												assign node48066 = (inp[2]) ? node48070 : node48067;
													assign node48067 = (inp[0]) ? 4'b0111 : 4'b0110;
													assign node48070 = (inp[0]) ? 4'b0110 : 4'b0111;
												assign node48073 = (inp[2]) ? node48077 : node48074;
													assign node48074 = (inp[0]) ? 4'b0111 : 4'b0110;
													assign node48077 = (inp[0]) ? 4'b0110 : 4'b0111;
											assign node48080 = (inp[10]) ? node48096 : node48081;
												assign node48081 = (inp[0]) ? node48089 : node48082;
													assign node48082 = (inp[2]) ? node48086 : node48083;
														assign node48083 = (inp[5]) ? 4'b0011 : 4'b0010;
														assign node48086 = (inp[5]) ? 4'b0010 : 4'b0011;
													assign node48089 = (inp[5]) ? node48093 : node48090;
														assign node48090 = (inp[2]) ? 4'b0010 : 4'b0011;
														assign node48093 = (inp[2]) ? 4'b0011 : 4'b0010;
												assign node48096 = (inp[9]) ? node48122 : node48097;
													assign node48097 = (inp[11]) ? node48107 : node48098;
														assign node48098 = (inp[2]) ? node48100 : 4'b0011;
															assign node48100 = (inp[5]) ? node48104 : node48101;
																assign node48101 = (inp[0]) ? 4'b0010 : 4'b0011;
																assign node48104 = (inp[0]) ? 4'b0011 : 4'b0010;
														assign node48107 = (inp[0]) ? node48115 : node48108;
															assign node48108 = (inp[2]) ? node48112 : node48109;
																assign node48109 = (inp[5]) ? 4'b0011 : 4'b0010;
																assign node48112 = (inp[5]) ? 4'b0010 : 4'b0011;
															assign node48115 = (inp[2]) ? node48119 : node48116;
																assign node48116 = (inp[5]) ? 4'b0010 : 4'b0011;
																assign node48119 = (inp[5]) ? 4'b0011 : 4'b0010;
													assign node48122 = (inp[5]) ? node48130 : node48123;
														assign node48123 = (inp[2]) ? node48127 : node48124;
															assign node48124 = (inp[0]) ? 4'b0011 : 4'b0010;
															assign node48127 = (inp[0]) ? 4'b0010 : 4'b0011;
														assign node48130 = (inp[11]) ? node48136 : node48131;
															assign node48131 = (inp[0]) ? node48133 : 4'b0010;
																assign node48133 = (inp[2]) ? 4'b0011 : 4'b0010;
															assign node48136 = (inp[2]) ? node48140 : node48137;
																assign node48137 = (inp[0]) ? 4'b0010 : 4'b0011;
																assign node48140 = (inp[0]) ? 4'b0011 : 4'b0010;
									assign node48143 = (inp[0]) ? node48215 : node48144;
										assign node48144 = (inp[2]) ? node48180 : node48145;
											assign node48145 = (inp[5]) ? node48157 : node48146;
												assign node48146 = (inp[8]) ? node48154 : node48147;
													assign node48147 = (inp[1]) ? node48151 : node48148;
														assign node48148 = (inp[9]) ? 4'b0010 : 4'b0011;
														assign node48151 = (inp[9]) ? 4'b0111 : 4'b0110;
													assign node48154 = (inp[1]) ? 4'b0011 : 4'b0111;
												assign node48157 = (inp[9]) ? node48173 : node48158;
													assign node48158 = (inp[11]) ? node48166 : node48159;
														assign node48159 = (inp[8]) ? node48163 : node48160;
															assign node48160 = (inp[1]) ? 4'b0110 : 4'b0010;
															assign node48163 = (inp[1]) ? 4'b0010 : 4'b0110;
														assign node48166 = (inp[1]) ? node48170 : node48167;
															assign node48167 = (inp[8]) ? 4'b0110 : 4'b0010;
															assign node48170 = (inp[8]) ? 4'b0010 : 4'b0110;
													assign node48173 = (inp[8]) ? node48177 : node48174;
														assign node48174 = (inp[1]) ? 4'b0111 : 4'b0011;
														assign node48177 = (inp[1]) ? 4'b0010 : 4'b0110;
											assign node48180 = (inp[5]) ? node48192 : node48181;
												assign node48181 = (inp[8]) ? node48189 : node48182;
													assign node48182 = (inp[1]) ? node48186 : node48183;
														assign node48183 = (inp[9]) ? 4'b0011 : 4'b0010;
														assign node48186 = (inp[9]) ? 4'b0110 : 4'b0111;
													assign node48189 = (inp[1]) ? 4'b0010 : 4'b0110;
												assign node48192 = (inp[9]) ? node48208 : node48193;
													assign node48193 = (inp[11]) ? node48201 : node48194;
														assign node48194 = (inp[8]) ? node48198 : node48195;
															assign node48195 = (inp[1]) ? 4'b0111 : 4'b0011;
															assign node48198 = (inp[1]) ? 4'b0011 : 4'b0111;
														assign node48201 = (inp[1]) ? node48205 : node48202;
															assign node48202 = (inp[8]) ? 4'b0111 : 4'b0011;
															assign node48205 = (inp[8]) ? 4'b0011 : 4'b0111;
													assign node48208 = (inp[8]) ? node48212 : node48209;
														assign node48209 = (inp[1]) ? 4'b0110 : 4'b0010;
														assign node48212 = (inp[1]) ? 4'b0011 : 4'b0111;
										assign node48215 = (inp[1]) ? node48239 : node48216;
											assign node48216 = (inp[8]) ? node48232 : node48217;
												assign node48217 = (inp[10]) ? node48225 : node48218;
													assign node48218 = (inp[2]) ? node48222 : node48219;
														assign node48219 = (inp[9]) ? 4'b0010 : 4'b0011;
														assign node48222 = (inp[9]) ? 4'b0011 : 4'b0010;
													assign node48225 = (inp[9]) ? node48229 : node48226;
														assign node48226 = (inp[2]) ? 4'b0010 : 4'b0011;
														assign node48229 = (inp[2]) ? 4'b0011 : 4'b0010;
												assign node48232 = (inp[2]) ? node48236 : node48233;
													assign node48233 = (inp[5]) ? 4'b0111 : 4'b0110;
													assign node48236 = (inp[5]) ? 4'b0110 : 4'b0111;
											assign node48239 = (inp[8]) ? node48291 : node48240;
												assign node48240 = (inp[11]) ? node48262 : node48241;
													assign node48241 = (inp[9]) ? node48255 : node48242;
														assign node48242 = (inp[10]) ? node48248 : node48243;
															assign node48243 = (inp[2]) ? 4'b0110 : node48244;
																assign node48244 = (inp[5]) ? 4'b0110 : 4'b0111;
															assign node48248 = (inp[2]) ? node48252 : node48249;
																assign node48249 = (inp[5]) ? 4'b0110 : 4'b0111;
																assign node48252 = (inp[5]) ? 4'b0111 : 4'b0110;
														assign node48255 = (inp[2]) ? node48259 : node48256;
															assign node48256 = (inp[5]) ? 4'b0111 : 4'b0110;
															assign node48259 = (inp[5]) ? 4'b0110 : 4'b0111;
													assign node48262 = (inp[5]) ? node48276 : node48263;
														assign node48263 = (inp[10]) ? node48271 : node48264;
															assign node48264 = (inp[9]) ? node48268 : node48265;
																assign node48265 = (inp[2]) ? 4'b0110 : 4'b0111;
																assign node48268 = (inp[2]) ? 4'b0111 : 4'b0110;
															assign node48271 = (inp[2]) ? 4'b0111 : node48272;
																assign node48272 = (inp[9]) ? 4'b0110 : 4'b0111;
														assign node48276 = (inp[10]) ? node48284 : node48277;
															assign node48277 = (inp[9]) ? node48281 : node48278;
																assign node48278 = (inp[2]) ? 4'b0111 : 4'b0110;
																assign node48281 = (inp[2]) ? 4'b0110 : 4'b0111;
															assign node48284 = (inp[2]) ? node48288 : node48285;
																assign node48285 = (inp[9]) ? 4'b0111 : 4'b0110;
																assign node48288 = (inp[9]) ? 4'b0110 : 4'b0111;
												assign node48291 = (inp[5]) ? node48295 : node48292;
													assign node48292 = (inp[2]) ? 4'b0011 : 4'b0010;
													assign node48295 = (inp[2]) ? 4'b0010 : 4'b0011;
							assign node48298 = (inp[12]) ? node48594 : node48299;
								assign node48299 = (inp[1]) ? node48493 : node48300;
									assign node48300 = (inp[15]) ? node48446 : node48301;
										assign node48301 = (inp[8]) ? node48407 : node48302;
											assign node48302 = (inp[0]) ? node48356 : node48303;
												assign node48303 = (inp[10]) ? node48327 : node48304;
													assign node48304 = (inp[5]) ? node48320 : node48305;
														assign node48305 = (inp[11]) ? node48313 : node48306;
															assign node48306 = (inp[9]) ? node48310 : node48307;
																assign node48307 = (inp[2]) ? 4'b0111 : 4'b0110;
																assign node48310 = (inp[2]) ? 4'b0110 : 4'b0111;
															assign node48313 = (inp[9]) ? node48317 : node48314;
																assign node48314 = (inp[2]) ? 4'b0111 : 4'b0110;
																assign node48317 = (inp[2]) ? 4'b0110 : 4'b0111;
														assign node48320 = (inp[11]) ? node48322 : 4'b0111;
															assign node48322 = (inp[2]) ? 4'b0111 : node48323;
																assign node48323 = (inp[9]) ? 4'b0110 : 4'b0111;
													assign node48327 = (inp[11]) ? node48341 : node48328;
														assign node48328 = (inp[5]) ? node48336 : node48329;
															assign node48329 = (inp[9]) ? node48333 : node48330;
																assign node48330 = (inp[2]) ? 4'b0111 : 4'b0110;
																assign node48333 = (inp[2]) ? 4'b0110 : 4'b0111;
															assign node48336 = (inp[2]) ? node48338 : 4'b0110;
																assign node48338 = (inp[9]) ? 4'b0111 : 4'b0110;
														assign node48341 = (inp[2]) ? node48349 : node48342;
															assign node48342 = (inp[9]) ? node48346 : node48343;
																assign node48343 = (inp[5]) ? 4'b0111 : 4'b0110;
																assign node48346 = (inp[5]) ? 4'b0110 : 4'b0111;
															assign node48349 = (inp[5]) ? node48353 : node48350;
																assign node48350 = (inp[9]) ? 4'b0110 : 4'b0111;
																assign node48353 = (inp[9]) ? 4'b0111 : 4'b0110;
												assign node48356 = (inp[5]) ? node48380 : node48357;
													assign node48357 = (inp[11]) ? node48373 : node48358;
														assign node48358 = (inp[10]) ? node48366 : node48359;
															assign node48359 = (inp[9]) ? node48363 : node48360;
																assign node48360 = (inp[2]) ? 4'b0111 : 4'b0110;
																assign node48363 = (inp[2]) ? 4'b0110 : 4'b0111;
															assign node48366 = (inp[9]) ? node48370 : node48367;
																assign node48367 = (inp[2]) ? 4'b0111 : 4'b0110;
																assign node48370 = (inp[2]) ? 4'b0110 : 4'b0111;
														assign node48373 = (inp[2]) ? node48377 : node48374;
															assign node48374 = (inp[9]) ? 4'b0111 : 4'b0110;
															assign node48377 = (inp[9]) ? 4'b0110 : 4'b0111;
													assign node48380 = (inp[11]) ? node48396 : node48381;
														assign node48381 = (inp[10]) ? node48389 : node48382;
															assign node48382 = (inp[2]) ? node48386 : node48383;
																assign node48383 = (inp[9]) ? 4'b0111 : 4'b0110;
																assign node48386 = (inp[9]) ? 4'b0110 : 4'b0111;
															assign node48389 = (inp[9]) ? node48393 : node48390;
																assign node48390 = (inp[2]) ? 4'b0111 : 4'b0110;
																assign node48393 = (inp[2]) ? 4'b0110 : 4'b0111;
														assign node48396 = (inp[10]) ? node48402 : node48397;
															assign node48397 = (inp[2]) ? node48399 : 4'b0110;
																assign node48399 = (inp[9]) ? 4'b0110 : 4'b0111;
															assign node48402 = (inp[9]) ? node48404 : 4'b0110;
																assign node48404 = (inp[2]) ? 4'b0110 : 4'b0111;
											assign node48407 = (inp[10]) ? node48415 : node48408;
												assign node48408 = (inp[2]) ? node48412 : node48409;
													assign node48409 = (inp[0]) ? 4'b0011 : 4'b0010;
													assign node48412 = (inp[0]) ? 4'b0010 : 4'b0011;
												assign node48415 = (inp[5]) ? node48439 : node48416;
													assign node48416 = (inp[9]) ? node48424 : node48417;
														assign node48417 = (inp[2]) ? node48421 : node48418;
															assign node48418 = (inp[0]) ? 4'b0011 : 4'b0010;
															assign node48421 = (inp[0]) ? 4'b0010 : 4'b0011;
														assign node48424 = (inp[11]) ? node48432 : node48425;
															assign node48425 = (inp[2]) ? node48429 : node48426;
																assign node48426 = (inp[0]) ? 4'b0011 : 4'b0010;
																assign node48429 = (inp[0]) ? 4'b0010 : 4'b0011;
															assign node48432 = (inp[0]) ? node48436 : node48433;
																assign node48433 = (inp[2]) ? 4'b0011 : 4'b0010;
																assign node48436 = (inp[2]) ? 4'b0010 : 4'b0011;
													assign node48439 = (inp[2]) ? node48443 : node48440;
														assign node48440 = (inp[0]) ? 4'b0011 : 4'b0010;
														assign node48443 = (inp[0]) ? 4'b0010 : 4'b0011;
										assign node48446 = (inp[0]) ? node48470 : node48447;
											assign node48447 = (inp[5]) ? node48459 : node48448;
												assign node48448 = (inp[2]) ? node48454 : node48449;
													assign node48449 = (inp[9]) ? 4'b0010 : node48450;
														assign node48450 = (inp[8]) ? 4'b0010 : 4'b0011;
													assign node48454 = (inp[9]) ? 4'b0011 : node48455;
														assign node48455 = (inp[8]) ? 4'b0011 : 4'b0010;
												assign node48459 = (inp[2]) ? node48465 : node48460;
													assign node48460 = (inp[8]) ? 4'b0011 : node48461;
														assign node48461 = (inp[9]) ? 4'b0010 : 4'b0011;
													assign node48465 = (inp[8]) ? 4'b0010 : node48466;
														assign node48466 = (inp[9]) ? 4'b0011 : 4'b0010;
											assign node48470 = (inp[5]) ? node48482 : node48471;
												assign node48471 = (inp[2]) ? node48477 : node48472;
													assign node48472 = (inp[9]) ? 4'b0011 : node48473;
														assign node48473 = (inp[8]) ? 4'b0011 : 4'b0010;
													assign node48477 = (inp[9]) ? 4'b0010 : node48478;
														assign node48478 = (inp[8]) ? 4'b0010 : 4'b0011;
												assign node48482 = (inp[2]) ? node48488 : node48483;
													assign node48483 = (inp[8]) ? 4'b0010 : node48484;
														assign node48484 = (inp[9]) ? 4'b0010 : 4'b0011;
													assign node48488 = (inp[8]) ? 4'b0011 : node48489;
														assign node48489 = (inp[9]) ? 4'b0011 : 4'b0010;
									assign node48493 = (inp[8]) ? node48533 : node48494;
										assign node48494 = (inp[0]) ? node48526 : node48495;
											assign node48495 = (inp[2]) ? node48519 : node48496;
												assign node48496 = (inp[15]) ? node48512 : node48497;
													assign node48497 = (inp[11]) ? node48505 : node48498;
														assign node48498 = (inp[5]) ? node48502 : node48499;
															assign node48499 = (inp[9]) ? 4'b0111 : 4'b0110;
															assign node48502 = (inp[9]) ? 4'b0110 : 4'b0111;
														assign node48505 = (inp[5]) ? node48509 : node48506;
															assign node48506 = (inp[9]) ? 4'b0111 : 4'b0110;
															assign node48509 = (inp[9]) ? 4'b0110 : 4'b0111;
													assign node48512 = (inp[9]) ? node48516 : node48513;
														assign node48513 = (inp[5]) ? 4'b0111 : 4'b0110;
														assign node48516 = (inp[5]) ? 4'b0110 : 4'b0111;
												assign node48519 = (inp[5]) ? node48523 : node48520;
													assign node48520 = (inp[9]) ? 4'b0110 : 4'b0111;
													assign node48523 = (inp[9]) ? 4'b0111 : 4'b0110;
											assign node48526 = (inp[2]) ? node48530 : node48527;
												assign node48527 = (inp[9]) ? 4'b0111 : 4'b0110;
												assign node48530 = (inp[9]) ? 4'b0110 : 4'b0111;
										assign node48533 = (inp[15]) ? node48565 : node48534;
											assign node48534 = (inp[9]) ? node48550 : node48535;
												assign node48535 = (inp[10]) ? node48543 : node48536;
													assign node48536 = (inp[0]) ? node48540 : node48537;
														assign node48537 = (inp[2]) ? 4'b0111 : 4'b0110;
														assign node48540 = (inp[2]) ? 4'b0110 : 4'b0111;
													assign node48543 = (inp[2]) ? node48547 : node48544;
														assign node48544 = (inp[0]) ? 4'b0111 : 4'b0110;
														assign node48547 = (inp[0]) ? 4'b0110 : 4'b0111;
												assign node48550 = (inp[10]) ? node48558 : node48551;
													assign node48551 = (inp[0]) ? node48555 : node48552;
														assign node48552 = (inp[2]) ? 4'b0111 : 4'b0110;
														assign node48555 = (inp[2]) ? 4'b0110 : 4'b0111;
													assign node48558 = (inp[2]) ? node48562 : node48559;
														assign node48559 = (inp[0]) ? 4'b0111 : 4'b0110;
														assign node48562 = (inp[0]) ? 4'b0110 : 4'b0111;
											assign node48565 = (inp[10]) ? node48573 : node48566;
												assign node48566 = (inp[0]) ? node48570 : node48567;
													assign node48567 = (inp[2]) ? 4'b0111 : 4'b0110;
													assign node48570 = (inp[2]) ? 4'b0110 : 4'b0111;
												assign node48573 = (inp[11]) ? node48587 : node48574;
													assign node48574 = (inp[5]) ? node48582 : node48575;
														assign node48575 = (inp[0]) ? node48579 : node48576;
															assign node48576 = (inp[2]) ? 4'b0111 : 4'b0110;
															assign node48579 = (inp[2]) ? 4'b0110 : 4'b0111;
														assign node48582 = (inp[0]) ? 4'b0111 : node48583;
															assign node48583 = (inp[2]) ? 4'b0111 : 4'b0110;
													assign node48587 = (inp[0]) ? node48591 : node48588;
														assign node48588 = (inp[2]) ? 4'b0111 : 4'b0110;
														assign node48591 = (inp[2]) ? 4'b0110 : 4'b0111;
								assign node48594 = (inp[1]) ? node48790 : node48595;
									assign node48595 = (inp[15]) ? node48737 : node48596;
										assign node48596 = (inp[8]) ? node48666 : node48597;
											assign node48597 = (inp[11]) ? node48639 : node48598;
												assign node48598 = (inp[10]) ? node48620 : node48599;
													assign node48599 = (inp[2]) ? node48609 : node48600;
														assign node48600 = (inp[9]) ? node48606 : node48601;
															assign node48601 = (inp[5]) ? node48603 : 4'b0011;
																assign node48603 = (inp[0]) ? 4'b0011 : 4'b0010;
															assign node48606 = (inp[0]) ? 4'b0010 : 4'b0011;
														assign node48609 = (inp[9]) ? node48615 : node48610;
															assign node48610 = (inp[0]) ? 4'b0010 : node48611;
																assign node48611 = (inp[5]) ? 4'b0011 : 4'b0010;
															assign node48615 = (inp[0]) ? 4'b0011 : node48616;
																assign node48616 = (inp[5]) ? 4'b0010 : 4'b0011;
													assign node48620 = (inp[9]) ? node48630 : node48621;
														assign node48621 = (inp[2]) ? node48625 : node48622;
															assign node48622 = (inp[5]) ? 4'b0010 : 4'b0011;
															assign node48625 = (inp[0]) ? 4'b0010 : node48626;
																assign node48626 = (inp[5]) ? 4'b0011 : 4'b0010;
														assign node48630 = (inp[2]) ? node48636 : node48631;
															assign node48631 = (inp[0]) ? 4'b0010 : node48632;
																assign node48632 = (inp[5]) ? 4'b0011 : 4'b0010;
															assign node48636 = (inp[5]) ? 4'b0010 : 4'b0011;
												assign node48639 = (inp[5]) ? node48647 : node48640;
													assign node48640 = (inp[9]) ? node48644 : node48641;
														assign node48641 = (inp[2]) ? 4'b0010 : 4'b0011;
														assign node48644 = (inp[2]) ? 4'b0011 : 4'b0010;
													assign node48647 = (inp[2]) ? node48655 : node48648;
														assign node48648 = (inp[9]) ? node48652 : node48649;
															assign node48649 = (inp[0]) ? 4'b0011 : 4'b0010;
															assign node48652 = (inp[0]) ? 4'b0010 : 4'b0011;
														assign node48655 = (inp[10]) ? node48661 : node48656;
															assign node48656 = (inp[9]) ? 4'b0011 : node48657;
																assign node48657 = (inp[0]) ? 4'b0010 : 4'b0011;
															assign node48661 = (inp[9]) ? node48663 : 4'b0011;
																assign node48663 = (inp[0]) ? 4'b0011 : 4'b0010;
											assign node48666 = (inp[10]) ? node48696 : node48667;
												assign node48667 = (inp[5]) ? node48683 : node48668;
													assign node48668 = (inp[11]) ? node48676 : node48669;
														assign node48669 = (inp[0]) ? node48673 : node48670;
															assign node48670 = (inp[2]) ? 4'b0110 : 4'b0111;
															assign node48673 = (inp[2]) ? 4'b0111 : 4'b0110;
														assign node48676 = (inp[2]) ? node48680 : node48677;
															assign node48677 = (inp[0]) ? 4'b0110 : 4'b0111;
															assign node48680 = (inp[0]) ? 4'b0111 : 4'b0110;
													assign node48683 = (inp[11]) ? node48691 : node48684;
														assign node48684 = (inp[2]) ? node48688 : node48685;
															assign node48685 = (inp[0]) ? 4'b0111 : 4'b0110;
															assign node48688 = (inp[0]) ? 4'b0110 : 4'b0111;
														assign node48691 = (inp[2]) ? node48693 : 4'b0110;
															assign node48693 = (inp[0]) ? 4'b0110 : 4'b0111;
												assign node48696 = (inp[11]) ? node48718 : node48697;
													assign node48697 = (inp[5]) ? node48705 : node48698;
														assign node48698 = (inp[0]) ? node48702 : node48699;
															assign node48699 = (inp[2]) ? 4'b0110 : 4'b0111;
															assign node48702 = (inp[2]) ? 4'b0111 : 4'b0110;
														assign node48705 = (inp[9]) ? node48711 : node48706;
															assign node48706 = (inp[2]) ? 4'b0111 : node48707;
																assign node48707 = (inp[0]) ? 4'b0111 : 4'b0110;
															assign node48711 = (inp[0]) ? node48715 : node48712;
																assign node48712 = (inp[2]) ? 4'b0111 : 4'b0110;
																assign node48715 = (inp[2]) ? 4'b0110 : 4'b0111;
													assign node48718 = (inp[9]) ? node48728 : node48719;
														assign node48719 = (inp[5]) ? 4'b0111 : node48720;
															assign node48720 = (inp[2]) ? node48724 : node48721;
																assign node48721 = (inp[0]) ? 4'b0110 : 4'b0111;
																assign node48724 = (inp[0]) ? 4'b0111 : 4'b0110;
														assign node48728 = (inp[5]) ? node48730 : 4'b0111;
															assign node48730 = (inp[2]) ? node48734 : node48731;
																assign node48731 = (inp[0]) ? 4'b0111 : 4'b0110;
																assign node48734 = (inp[0]) ? 4'b0110 : 4'b0111;
										assign node48737 = (inp[9]) ? node48775 : node48738;
											assign node48738 = (inp[2]) ? node48748 : node48739;
												assign node48739 = (inp[8]) ? node48745 : node48740;
													assign node48740 = (inp[0]) ? 4'b0110 : node48741;
														assign node48741 = (inp[5]) ? 4'b0111 : 4'b0110;
													assign node48745 = (inp[0]) ? 4'b0111 : 4'b0110;
												assign node48748 = (inp[5]) ? node48754 : node48749;
													assign node48749 = (inp[0]) ? node48751 : 4'b0111;
														assign node48751 = (inp[8]) ? 4'b0110 : 4'b0111;
													assign node48754 = (inp[10]) ? node48768 : node48755;
														assign node48755 = (inp[11]) ? node48761 : node48756;
															assign node48756 = (inp[8]) ? node48758 : 4'b0110;
																assign node48758 = (inp[0]) ? 4'b0110 : 4'b0111;
															assign node48761 = (inp[8]) ? node48765 : node48762;
																assign node48762 = (inp[0]) ? 4'b0111 : 4'b0110;
																assign node48765 = (inp[0]) ? 4'b0110 : 4'b0111;
														assign node48768 = (inp[8]) ? node48772 : node48769;
															assign node48769 = (inp[0]) ? 4'b0111 : 4'b0110;
															assign node48772 = (inp[0]) ? 4'b0110 : 4'b0111;
											assign node48775 = (inp[2]) ? node48783 : node48776;
												assign node48776 = (inp[0]) ? 4'b0111 : node48777;
													assign node48777 = (inp[8]) ? 4'b0110 : node48778;
														assign node48778 = (inp[5]) ? 4'b0110 : 4'b0111;
												assign node48783 = (inp[0]) ? 4'b0110 : node48784;
													assign node48784 = (inp[8]) ? 4'b0111 : node48785;
														assign node48785 = (inp[5]) ? 4'b0111 : 4'b0110;
									assign node48790 = (inp[10]) ? node48830 : node48791;
										assign node48791 = (inp[9]) ? node48815 : node48792;
											assign node48792 = (inp[2]) ? node48806 : node48793;
												assign node48793 = (inp[5]) ? node48799 : node48794;
													assign node48794 = (inp[0]) ? node48796 : 4'b0010;
														assign node48796 = (inp[8]) ? 4'b0011 : 4'b0010;
													assign node48799 = (inp[0]) ? node48803 : node48800;
														assign node48800 = (inp[8]) ? 4'b0010 : 4'b0011;
														assign node48803 = (inp[8]) ? 4'b0011 : 4'b0010;
												assign node48806 = (inp[8]) ? node48812 : node48807;
													assign node48807 = (inp[0]) ? 4'b0011 : node48808;
														assign node48808 = (inp[5]) ? 4'b0010 : 4'b0011;
													assign node48812 = (inp[0]) ? 4'b0010 : 4'b0011;
											assign node48815 = (inp[2]) ? node48823 : node48816;
												assign node48816 = (inp[0]) ? 4'b0011 : node48817;
													assign node48817 = (inp[8]) ? 4'b0010 : node48818;
														assign node48818 = (inp[5]) ? 4'b0010 : 4'b0011;
												assign node48823 = (inp[0]) ? 4'b0010 : node48824;
													assign node48824 = (inp[5]) ? 4'b0011 : node48825;
														assign node48825 = (inp[8]) ? 4'b0011 : 4'b0010;
										assign node48830 = (inp[8]) ? node48878 : node48831;
											assign node48831 = (inp[11]) ? node48855 : node48832;
												assign node48832 = (inp[2]) ? node48844 : node48833;
													assign node48833 = (inp[9]) ? node48839 : node48834;
														assign node48834 = (inp[5]) ? node48836 : 4'b0010;
															assign node48836 = (inp[0]) ? 4'b0010 : 4'b0011;
														assign node48839 = (inp[0]) ? 4'b0011 : node48840;
															assign node48840 = (inp[5]) ? 4'b0010 : 4'b0011;
													assign node48844 = (inp[9]) ? node48850 : node48845;
														assign node48845 = (inp[5]) ? node48847 : 4'b0011;
															assign node48847 = (inp[0]) ? 4'b0011 : 4'b0010;
														assign node48850 = (inp[0]) ? 4'b0010 : node48851;
															assign node48851 = (inp[5]) ? 4'b0011 : 4'b0010;
												assign node48855 = (inp[9]) ? node48867 : node48856;
													assign node48856 = (inp[2]) ? node48862 : node48857;
														assign node48857 = (inp[0]) ? 4'b0010 : node48858;
															assign node48858 = (inp[5]) ? 4'b0011 : 4'b0010;
														assign node48862 = (inp[5]) ? node48864 : 4'b0011;
															assign node48864 = (inp[0]) ? 4'b0011 : 4'b0010;
													assign node48867 = (inp[2]) ? node48873 : node48868;
														assign node48868 = (inp[5]) ? node48870 : 4'b0011;
															assign node48870 = (inp[0]) ? 4'b0011 : 4'b0010;
														assign node48873 = (inp[5]) ? node48875 : 4'b0010;
															assign node48875 = (inp[0]) ? 4'b0010 : 4'b0011;
											assign node48878 = (inp[15]) ? node48902 : node48879;
												assign node48879 = (inp[11]) ? node48895 : node48880;
													assign node48880 = (inp[9]) ? node48888 : node48881;
														assign node48881 = (inp[0]) ? node48885 : node48882;
															assign node48882 = (inp[2]) ? 4'b0011 : 4'b0010;
															assign node48885 = (inp[2]) ? 4'b0010 : 4'b0011;
														assign node48888 = (inp[0]) ? node48892 : node48889;
															assign node48889 = (inp[2]) ? 4'b0011 : 4'b0010;
															assign node48892 = (inp[2]) ? 4'b0010 : 4'b0011;
													assign node48895 = (inp[2]) ? node48899 : node48896;
														assign node48896 = (inp[0]) ? 4'b0011 : 4'b0010;
														assign node48899 = (inp[0]) ? 4'b0010 : 4'b0011;
												assign node48902 = (inp[2]) ? node48906 : node48903;
													assign node48903 = (inp[0]) ? 4'b0011 : 4'b0010;
													assign node48906 = (inp[0]) ? 4'b0010 : 4'b0011;
					assign node48909 = (inp[7]) ? node50083 : node48910;
						assign node48910 = (inp[8]) ? node49908 : node48911;
							assign node48911 = (inp[11]) ? node49539 : node48912;
								assign node48912 = (inp[10]) ? node49212 : node48913;
									assign node48913 = (inp[2]) ? node49061 : node48914;
										assign node48914 = (inp[9]) ? node48976 : node48915;
											assign node48915 = (inp[12]) ? node48951 : node48916;
												assign node48916 = (inp[13]) ? node48932 : node48917;
													assign node48917 = (inp[1]) ? node48923 : node48918;
														assign node48918 = (inp[5]) ? 4'b0010 : node48919;
															assign node48919 = (inp[0]) ? 4'b0011 : 4'b0010;
														assign node48923 = (inp[15]) ? node48927 : node48924;
															assign node48924 = (inp[0]) ? 4'b0111 : 4'b0110;
															assign node48927 = (inp[0]) ? node48929 : 4'b0011;
																assign node48929 = (inp[5]) ? 4'b0011 : 4'b0010;
													assign node48932 = (inp[5]) ? node48938 : node48933;
														assign node48933 = (inp[15]) ? node48935 : 4'b0110;
															assign node48935 = (inp[1]) ? 4'b0110 : 4'b0111;
														assign node48938 = (inp[15]) ? node48944 : node48939;
															assign node48939 = (inp[1]) ? 4'b0011 : node48940;
																assign node48940 = (inp[0]) ? 4'b0110 : 4'b0111;
															assign node48944 = (inp[0]) ? node48948 : node48945;
																assign node48945 = (inp[1]) ? 4'b0111 : 4'b0110;
																assign node48948 = (inp[1]) ? 4'b0110 : 4'b0111;
												assign node48951 = (inp[13]) ? node48963 : node48952;
													assign node48952 = (inp[5]) ? node48956 : node48953;
														assign node48953 = (inp[0]) ? 4'b0111 : 4'b0110;
														assign node48956 = (inp[0]) ? 4'b0110 : node48957;
															assign node48957 = (inp[1]) ? node48959 : 4'b0110;
																assign node48959 = (inp[15]) ? 4'b0110 : 4'b0010;
													assign node48963 = (inp[15]) ? node48971 : node48964;
														assign node48964 = (inp[1]) ? node48966 : 4'b0010;
															assign node48966 = (inp[5]) ? 4'b0110 : node48967;
																assign node48967 = (inp[0]) ? 4'b0111 : 4'b0110;
														assign node48971 = (inp[5]) ? 4'b0010 : node48972;
															assign node48972 = (inp[0]) ? 4'b0011 : 4'b0010;
											assign node48976 = (inp[5]) ? node49026 : node48977;
												assign node48977 = (inp[0]) ? node49003 : node48978;
													assign node48978 = (inp[1]) ? node48990 : node48979;
														assign node48979 = (inp[13]) ? node48983 : node48980;
															assign node48980 = (inp[12]) ? 4'b0111 : 4'b0011;
															assign node48983 = (inp[12]) ? node48987 : node48984;
																assign node48984 = (inp[15]) ? 4'b0110 : 4'b0111;
																assign node48987 = (inp[15]) ? 4'b0011 : 4'b0010;
														assign node48990 = (inp[13]) ? node48998 : node48991;
															assign node48991 = (inp[12]) ? node48995 : node48992;
																assign node48992 = (inp[15]) ? 4'b0010 : 4'b0111;
																assign node48995 = (inp[15]) ? 4'b0111 : 4'b0010;
															assign node48998 = (inp[12]) ? 4'b0111 : node48999;
																assign node48999 = (inp[15]) ? 4'b0111 : 4'b0010;
													assign node49003 = (inp[13]) ? node49015 : node49004;
														assign node49004 = (inp[12]) ? node49010 : node49005;
															assign node49005 = (inp[1]) ? node49007 : 4'b0010;
																assign node49007 = (inp[15]) ? 4'b0011 : 4'b0110;
															assign node49010 = (inp[1]) ? node49012 : 4'b0110;
																assign node49012 = (inp[15]) ? 4'b0110 : 4'b0010;
														assign node49015 = (inp[15]) ? node49021 : node49016;
															assign node49016 = (inp[12]) ? node49018 : 4'b0011;
																assign node49018 = (inp[1]) ? 4'b0110 : 4'b0011;
															assign node49021 = (inp[12]) ? 4'b0010 : node49022;
																assign node49022 = (inp[1]) ? 4'b0111 : 4'b0110;
												assign node49026 = (inp[12]) ? node49048 : node49027;
													assign node49027 = (inp[13]) ? node49035 : node49028;
														assign node49028 = (inp[15]) ? node49032 : node49029;
															assign node49029 = (inp[1]) ? 4'b0111 : 4'b0011;
															assign node49032 = (inp[1]) ? 4'b0010 : 4'b0011;
														assign node49035 = (inp[15]) ? node49041 : node49036;
															assign node49036 = (inp[1]) ? 4'b0010 : node49037;
																assign node49037 = (inp[0]) ? 4'b0111 : 4'b0110;
															assign node49041 = (inp[0]) ? node49045 : node49042;
																assign node49042 = (inp[1]) ? 4'b0110 : 4'b0111;
																assign node49045 = (inp[1]) ? 4'b0111 : 4'b0110;
													assign node49048 = (inp[13]) ? node49056 : node49049;
														assign node49049 = (inp[15]) ? 4'b0111 : node49050;
															assign node49050 = (inp[1]) ? node49052 : 4'b0111;
																assign node49052 = (inp[0]) ? 4'b0010 : 4'b0011;
														assign node49056 = (inp[15]) ? 4'b0011 : node49057;
															assign node49057 = (inp[1]) ? 4'b0111 : 4'b0010;
										assign node49061 = (inp[9]) ? node49137 : node49062;
											assign node49062 = (inp[13]) ? node49092 : node49063;
												assign node49063 = (inp[12]) ? node49079 : node49064;
													assign node49064 = (inp[1]) ? node49070 : node49065;
														assign node49065 = (inp[0]) ? node49067 : 4'b0011;
															assign node49067 = (inp[5]) ? 4'b0011 : 4'b0010;
														assign node49070 = (inp[15]) ? node49076 : node49071;
															assign node49071 = (inp[5]) ? 4'b0111 : node49072;
																assign node49072 = (inp[0]) ? 4'b0110 : 4'b0111;
															assign node49076 = (inp[5]) ? 4'b0010 : 4'b0011;
													assign node49079 = (inp[1]) ? node49085 : node49080;
														assign node49080 = (inp[5]) ? 4'b0111 : node49081;
															assign node49081 = (inp[0]) ? 4'b0110 : 4'b0111;
														assign node49085 = (inp[15]) ? node49087 : 4'b0010;
															assign node49087 = (inp[0]) ? node49089 : 4'b0111;
																assign node49089 = (inp[5]) ? 4'b0111 : 4'b0110;
												assign node49092 = (inp[12]) ? node49114 : node49093;
													assign node49093 = (inp[1]) ? node49105 : node49094;
														assign node49094 = (inp[15]) ? node49100 : node49095;
															assign node49095 = (inp[0]) ? 4'b0111 : node49096;
																assign node49096 = (inp[5]) ? 4'b0110 : 4'b0111;
															assign node49100 = (inp[0]) ? 4'b0110 : node49101;
																assign node49101 = (inp[5]) ? 4'b0111 : 4'b0110;
														assign node49105 = (inp[15]) ? node49111 : node49106;
															assign node49106 = (inp[5]) ? 4'b0010 : node49107;
																assign node49107 = (inp[0]) ? 4'b0011 : 4'b0010;
															assign node49111 = (inp[0]) ? 4'b0111 : 4'b0110;
													assign node49114 = (inp[1]) ? node49126 : node49115;
														assign node49115 = (inp[15]) ? node49121 : node49116;
															assign node49116 = (inp[0]) ? node49118 : 4'b0010;
																assign node49118 = (inp[5]) ? 4'b0010 : 4'b0011;
															assign node49121 = (inp[0]) ? node49123 : 4'b0011;
																assign node49123 = (inp[5]) ? 4'b0011 : 4'b0010;
														assign node49126 = (inp[15]) ? node49132 : node49127;
															assign node49127 = (inp[5]) ? 4'b0111 : node49128;
																assign node49128 = (inp[0]) ? 4'b0110 : 4'b0111;
															assign node49132 = (inp[5]) ? 4'b0011 : node49133;
																assign node49133 = (inp[0]) ? 4'b0010 : 4'b0011;
											assign node49137 = (inp[0]) ? node49169 : node49138;
												assign node49138 = (inp[13]) ? node49150 : node49139;
													assign node49139 = (inp[12]) ? node49145 : node49140;
														assign node49140 = (inp[1]) ? node49142 : 4'b0010;
															assign node49142 = (inp[15]) ? 4'b0011 : 4'b0110;
														assign node49145 = (inp[1]) ? node49147 : 4'b0110;
															assign node49147 = (inp[15]) ? 4'b0110 : 4'b0011;
													assign node49150 = (inp[12]) ? node49164 : node49151;
														assign node49151 = (inp[1]) ? node49159 : node49152;
															assign node49152 = (inp[5]) ? node49156 : node49153;
																assign node49153 = (inp[15]) ? 4'b0111 : 4'b0110;
																assign node49156 = (inp[15]) ? 4'b0110 : 4'b0111;
															assign node49159 = (inp[15]) ? node49161 : 4'b0011;
																assign node49161 = (inp[5]) ? 4'b0111 : 4'b0110;
														assign node49164 = (inp[15]) ? 4'b0010 : node49165;
															assign node49165 = (inp[1]) ? 4'b0110 : 4'b0011;
												assign node49169 = (inp[12]) ? node49195 : node49170;
													assign node49170 = (inp[13]) ? node49186 : node49171;
														assign node49171 = (inp[5]) ? node49179 : node49172;
															assign node49172 = (inp[15]) ? node49176 : node49173;
																assign node49173 = (inp[1]) ? 4'b0111 : 4'b0011;
																assign node49176 = (inp[1]) ? 4'b0010 : 4'b0011;
															assign node49179 = (inp[15]) ? node49183 : node49180;
																assign node49180 = (inp[1]) ? 4'b0110 : 4'b0010;
																assign node49183 = (inp[1]) ? 4'b0011 : 4'b0010;
														assign node49186 = (inp[1]) ? node49190 : node49187;
															assign node49187 = (inp[15]) ? 4'b0111 : 4'b0110;
															assign node49190 = (inp[15]) ? 4'b0110 : node49191;
																assign node49191 = (inp[5]) ? 4'b0011 : 4'b0010;
													assign node49195 = (inp[15]) ? node49209 : node49196;
														assign node49196 = (inp[13]) ? node49202 : node49197;
															assign node49197 = (inp[1]) ? 4'b0011 : node49198;
																assign node49198 = (inp[5]) ? 4'b0110 : 4'b0111;
															assign node49202 = (inp[1]) ? node49206 : node49203;
																assign node49203 = (inp[5]) ? 4'b0011 : 4'b0010;
																assign node49206 = (inp[5]) ? 4'b0110 : 4'b0111;
														assign node49209 = (inp[13]) ? 4'b0011 : 4'b0111;
									assign node49212 = (inp[9]) ? node49376 : node49213;
										assign node49213 = (inp[2]) ? node49295 : node49214;
											assign node49214 = (inp[0]) ? node49246 : node49215;
												assign node49215 = (inp[1]) ? node49229 : node49216;
													assign node49216 = (inp[13]) ? node49220 : node49217;
														assign node49217 = (inp[12]) ? 4'b0110 : 4'b0010;
														assign node49220 = (inp[12]) ? node49226 : node49221;
															assign node49221 = (inp[15]) ? node49223 : 4'b0110;
																assign node49223 = (inp[5]) ? 4'b0110 : 4'b0111;
															assign node49226 = (inp[15]) ? 4'b0010 : 4'b0011;
													assign node49229 = (inp[12]) ? node49239 : node49230;
														assign node49230 = (inp[15]) ? node49234 : node49231;
															assign node49231 = (inp[13]) ? 4'b0011 : 4'b0110;
															assign node49234 = (inp[13]) ? node49236 : 4'b0011;
																assign node49236 = (inp[5]) ? 4'b0111 : 4'b0110;
														assign node49239 = (inp[15]) ? node49243 : node49240;
															assign node49240 = (inp[5]) ? 4'b0010 : 4'b0011;
															assign node49243 = (inp[13]) ? 4'b0010 : 4'b0110;
												assign node49246 = (inp[5]) ? node49274 : node49247;
													assign node49247 = (inp[13]) ? node49261 : node49248;
														assign node49248 = (inp[12]) ? node49256 : node49249;
															assign node49249 = (inp[15]) ? node49253 : node49250;
																assign node49250 = (inp[1]) ? 4'b0111 : 4'b0011;
																assign node49253 = (inp[1]) ? 4'b0010 : 4'b0011;
															assign node49256 = (inp[15]) ? 4'b0111 : node49257;
																assign node49257 = (inp[1]) ? 4'b0011 : 4'b0111;
														assign node49261 = (inp[12]) ? node49269 : node49262;
															assign node49262 = (inp[15]) ? node49266 : node49263;
																assign node49263 = (inp[1]) ? 4'b0010 : 4'b0110;
																assign node49266 = (inp[1]) ? 4'b0110 : 4'b0111;
															assign node49269 = (inp[15]) ? 4'b0011 : node49270;
																assign node49270 = (inp[1]) ? 4'b0111 : 4'b0010;
													assign node49274 = (inp[15]) ? node49286 : node49275;
														assign node49275 = (inp[13]) ? node49279 : node49276;
															assign node49276 = (inp[12]) ? 4'b0011 : 4'b0010;
															assign node49279 = (inp[1]) ? node49283 : node49280;
																assign node49280 = (inp[12]) ? 4'b0011 : 4'b0110;
																assign node49283 = (inp[12]) ? 4'b0110 : 4'b0011;
														assign node49286 = (inp[12]) ? node49292 : node49287;
															assign node49287 = (inp[13]) ? node49289 : 4'b0011;
																assign node49289 = (inp[1]) ? 4'b0110 : 4'b0111;
															assign node49292 = (inp[13]) ? 4'b0010 : 4'b0110;
											assign node49295 = (inp[0]) ? node49331 : node49296;
												assign node49296 = (inp[1]) ? node49310 : node49297;
													assign node49297 = (inp[13]) ? node49301 : node49298;
														assign node49298 = (inp[12]) ? 4'b0111 : 4'b0011;
														assign node49301 = (inp[12]) ? node49307 : node49302;
															assign node49302 = (inp[5]) ? node49304 : 4'b0111;
																assign node49304 = (inp[15]) ? 4'b0111 : 4'b0110;
															assign node49307 = (inp[15]) ? 4'b0011 : 4'b0010;
													assign node49310 = (inp[12]) ? node49320 : node49311;
														assign node49311 = (inp[13]) ? node49315 : node49312;
															assign node49312 = (inp[15]) ? 4'b0010 : 4'b0111;
															assign node49315 = (inp[15]) ? node49317 : 4'b0010;
																assign node49317 = (inp[5]) ? 4'b0110 : 4'b0111;
														assign node49320 = (inp[5]) ? node49326 : node49321;
															assign node49321 = (inp[15]) ? 4'b0111 : node49322;
																assign node49322 = (inp[13]) ? 4'b0111 : 4'b0010;
															assign node49326 = (inp[13]) ? node49328 : 4'b0111;
																assign node49328 = (inp[15]) ? 4'b0011 : 4'b0111;
												assign node49331 = (inp[5]) ? node49353 : node49332;
													assign node49332 = (inp[13]) ? node49342 : node49333;
														assign node49333 = (inp[12]) ? node49339 : node49334;
															assign node49334 = (inp[1]) ? node49336 : 4'b0010;
																assign node49336 = (inp[15]) ? 4'b0011 : 4'b0110;
															assign node49339 = (inp[1]) ? 4'b0010 : 4'b0110;
														assign node49342 = (inp[12]) ? node49348 : node49343;
															assign node49343 = (inp[15]) ? node49345 : 4'b0011;
																assign node49345 = (inp[1]) ? 4'b0111 : 4'b0110;
															assign node49348 = (inp[15]) ? 4'b0010 : node49349;
																assign node49349 = (inp[1]) ? 4'b0110 : 4'b0011;
													assign node49353 = (inp[1]) ? node49365 : node49354;
														assign node49354 = (inp[13]) ? node49358 : node49355;
															assign node49355 = (inp[12]) ? 4'b0111 : 4'b0011;
															assign node49358 = (inp[12]) ? node49362 : node49359;
																assign node49359 = (inp[15]) ? 4'b0110 : 4'b0111;
																assign node49362 = (inp[15]) ? 4'b0011 : 4'b0010;
														assign node49365 = (inp[12]) ? node49373 : node49366;
															assign node49366 = (inp[13]) ? node49370 : node49367;
																assign node49367 = (inp[15]) ? 4'b0010 : 4'b0111;
																assign node49370 = (inp[15]) ? 4'b0111 : 4'b0010;
															assign node49373 = (inp[13]) ? 4'b0011 : 4'b0010;
										assign node49376 = (inp[2]) ? node49456 : node49377;
											assign node49377 = (inp[5]) ? node49425 : node49378;
												assign node49378 = (inp[0]) ? node49404 : node49379;
													assign node49379 = (inp[15]) ? node49393 : node49380;
														assign node49380 = (inp[12]) ? node49386 : node49381;
															assign node49381 = (inp[1]) ? node49383 : 4'b0111;
																assign node49383 = (inp[13]) ? 4'b0010 : 4'b0111;
															assign node49386 = (inp[1]) ? node49390 : node49387;
																assign node49387 = (inp[13]) ? 4'b0010 : 4'b0111;
																assign node49390 = (inp[13]) ? 4'b0111 : 4'b0010;
														assign node49393 = (inp[12]) ? node49401 : node49394;
															assign node49394 = (inp[13]) ? node49398 : node49395;
																assign node49395 = (inp[1]) ? 4'b0010 : 4'b0011;
																assign node49398 = (inp[1]) ? 4'b0111 : 4'b0110;
															assign node49401 = (inp[13]) ? 4'b0011 : 4'b0111;
													assign node49404 = (inp[12]) ? node49414 : node49405;
														assign node49405 = (inp[13]) ? 4'b0111 : node49406;
															assign node49406 = (inp[15]) ? node49410 : node49407;
																assign node49407 = (inp[1]) ? 4'b0110 : 4'b0010;
																assign node49410 = (inp[1]) ? 4'b0011 : 4'b0010;
														assign node49414 = (inp[13]) ? node49420 : node49415;
															assign node49415 = (inp[1]) ? node49417 : 4'b0110;
																assign node49417 = (inp[15]) ? 4'b0110 : 4'b0010;
															assign node49420 = (inp[15]) ? 4'b0010 : node49421;
																assign node49421 = (inp[1]) ? 4'b0110 : 4'b0011;
												assign node49425 = (inp[13]) ? node49439 : node49426;
													assign node49426 = (inp[12]) ? node49432 : node49427;
														assign node49427 = (inp[15]) ? 4'b0010 : node49428;
															assign node49428 = (inp[1]) ? 4'b0111 : 4'b0011;
														assign node49432 = (inp[1]) ? node49434 : 4'b0111;
															assign node49434 = (inp[15]) ? 4'b0111 : node49435;
																assign node49435 = (inp[0]) ? 4'b0010 : 4'b0011;
													assign node49439 = (inp[12]) ? node49451 : node49440;
														assign node49440 = (inp[0]) ? node49446 : node49441;
															assign node49441 = (inp[15]) ? 4'b0110 : node49442;
																assign node49442 = (inp[1]) ? 4'b0010 : 4'b0110;
															assign node49446 = (inp[15]) ? node49448 : 4'b0111;
																assign node49448 = (inp[1]) ? 4'b0111 : 4'b0110;
														assign node49451 = (inp[15]) ? 4'b0011 : node49452;
															assign node49452 = (inp[1]) ? 4'b0111 : 4'b0010;
											assign node49456 = (inp[1]) ? node49496 : node49457;
												assign node49457 = (inp[5]) ? node49483 : node49458;
													assign node49458 = (inp[0]) ? node49470 : node49459;
														assign node49459 = (inp[13]) ? node49463 : node49460;
															assign node49460 = (inp[12]) ? 4'b0110 : 4'b0010;
															assign node49463 = (inp[12]) ? node49467 : node49464;
																assign node49464 = (inp[15]) ? 4'b0111 : 4'b0110;
																assign node49467 = (inp[15]) ? 4'b0010 : 4'b0011;
														assign node49470 = (inp[15]) ? node49478 : node49471;
															assign node49471 = (inp[13]) ? node49475 : node49472;
																assign node49472 = (inp[12]) ? 4'b0111 : 4'b0011;
																assign node49475 = (inp[12]) ? 4'b0010 : 4'b0110;
															assign node49478 = (inp[12]) ? node49480 : 4'b0111;
																assign node49480 = (inp[13]) ? 4'b0011 : 4'b0111;
													assign node49483 = (inp[13]) ? node49487 : node49484;
														assign node49484 = (inp[12]) ? 4'b0110 : 4'b0010;
														assign node49487 = (inp[12]) ? 4'b0010 : node49488;
															assign node49488 = (inp[15]) ? node49492 : node49489;
																assign node49489 = (inp[0]) ? 4'b0110 : 4'b0111;
																assign node49492 = (inp[0]) ? 4'b0111 : 4'b0110;
												assign node49496 = (inp[15]) ? node49516 : node49497;
													assign node49497 = (inp[0]) ? node49507 : node49498;
														assign node49498 = (inp[13]) ? node49504 : node49499;
															assign node49499 = (inp[12]) ? node49501 : 4'b0110;
																assign node49501 = (inp[5]) ? 4'b0010 : 4'b0011;
															assign node49504 = (inp[12]) ? 4'b0110 : 4'b0011;
														assign node49507 = (inp[13]) ? node49509 : 4'b0011;
															assign node49509 = (inp[12]) ? node49513 : node49510;
																assign node49510 = (inp[5]) ? 4'b0011 : 4'b0010;
																assign node49513 = (inp[5]) ? 4'b0110 : 4'b0111;
													assign node49516 = (inp[12]) ? node49528 : node49517;
														assign node49517 = (inp[13]) ? node49523 : node49518;
															assign node49518 = (inp[5]) ? 4'b0011 : node49519;
																assign node49519 = (inp[0]) ? 4'b0010 : 4'b0011;
															assign node49523 = (inp[5]) ? node49525 : 4'b0110;
																assign node49525 = (inp[0]) ? 4'b0110 : 4'b0111;
														assign node49528 = (inp[13]) ? node49534 : node49529;
															assign node49529 = (inp[5]) ? 4'b0110 : node49530;
																assign node49530 = (inp[0]) ? 4'b0111 : 4'b0110;
															assign node49534 = (inp[5]) ? 4'b0010 : node49535;
																assign node49535 = (inp[0]) ? 4'b0011 : 4'b0010;
								assign node49539 = (inp[9]) ? node49723 : node49540;
									assign node49540 = (inp[2]) ? node49634 : node49541;
										assign node49541 = (inp[5]) ? node49599 : node49542;
											assign node49542 = (inp[0]) ? node49570 : node49543;
												assign node49543 = (inp[13]) ? node49557 : node49544;
													assign node49544 = (inp[12]) ? node49552 : node49545;
														assign node49545 = (inp[15]) ? node49549 : node49546;
															assign node49546 = (inp[1]) ? 4'b0110 : 4'b0010;
															assign node49549 = (inp[1]) ? 4'b0011 : 4'b0010;
														assign node49552 = (inp[1]) ? node49554 : 4'b0110;
															assign node49554 = (inp[15]) ? 4'b0110 : 4'b0011;
													assign node49557 = (inp[12]) ? node49565 : node49558;
														assign node49558 = (inp[1]) ? node49562 : node49559;
															assign node49559 = (inp[15]) ? 4'b0111 : 4'b0110;
															assign node49562 = (inp[15]) ? 4'b0110 : 4'b0011;
														assign node49565 = (inp[15]) ? 4'b0010 : node49566;
															assign node49566 = (inp[1]) ? 4'b0110 : 4'b0011;
												assign node49570 = (inp[12]) ? node49586 : node49571;
													assign node49571 = (inp[13]) ? node49579 : node49572;
														assign node49572 = (inp[15]) ? node49576 : node49573;
															assign node49573 = (inp[1]) ? 4'b0111 : 4'b0011;
															assign node49576 = (inp[1]) ? 4'b0010 : 4'b0011;
														assign node49579 = (inp[1]) ? node49583 : node49580;
															assign node49580 = (inp[15]) ? 4'b0111 : 4'b0110;
															assign node49583 = (inp[15]) ? 4'b0110 : 4'b0010;
													assign node49586 = (inp[1]) ? node49592 : node49587;
														assign node49587 = (inp[10]) ? 4'b0010 : node49588;
															assign node49588 = (inp[13]) ? 4'b0011 : 4'b0111;
														assign node49592 = (inp[13]) ? node49596 : node49593;
															assign node49593 = (inp[15]) ? 4'b0111 : 4'b0011;
															assign node49596 = (inp[15]) ? 4'b0011 : 4'b0111;
											assign node49599 = (inp[12]) ? node49621 : node49600;
												assign node49600 = (inp[13]) ? node49608 : node49601;
													assign node49601 = (inp[15]) ? node49605 : node49602;
														assign node49602 = (inp[1]) ? 4'b0110 : 4'b0010;
														assign node49605 = (inp[1]) ? 4'b0011 : 4'b0010;
													assign node49608 = (inp[15]) ? node49614 : node49609;
														assign node49609 = (inp[1]) ? 4'b0011 : node49610;
															assign node49610 = (inp[0]) ? 4'b0110 : 4'b0111;
														assign node49614 = (inp[0]) ? node49618 : node49615;
															assign node49615 = (inp[1]) ? 4'b0111 : 4'b0110;
															assign node49618 = (inp[1]) ? 4'b0110 : 4'b0111;
												assign node49621 = (inp[13]) ? node49629 : node49622;
													assign node49622 = (inp[1]) ? node49624 : 4'b0110;
														assign node49624 = (inp[15]) ? 4'b0110 : node49625;
															assign node49625 = (inp[0]) ? 4'b0011 : 4'b0010;
													assign node49629 = (inp[15]) ? 4'b0010 : node49630;
														assign node49630 = (inp[1]) ? 4'b0110 : 4'b0011;
										assign node49634 = (inp[0]) ? node49670 : node49635;
											assign node49635 = (inp[13]) ? node49649 : node49636;
												assign node49636 = (inp[12]) ? node49642 : node49637;
													assign node49637 = (inp[1]) ? node49639 : 4'b0011;
														assign node49639 = (inp[15]) ? 4'b0010 : 4'b0111;
													assign node49642 = (inp[1]) ? node49644 : 4'b0111;
														assign node49644 = (inp[15]) ? 4'b0111 : node49645;
															assign node49645 = (inp[5]) ? 4'b0011 : 4'b0010;
												assign node49649 = (inp[12]) ? node49663 : node49650;
													assign node49650 = (inp[1]) ? node49658 : node49651;
														assign node49651 = (inp[15]) ? node49655 : node49652;
															assign node49652 = (inp[5]) ? 4'b0110 : 4'b0111;
															assign node49655 = (inp[5]) ? 4'b0111 : 4'b0110;
														assign node49658 = (inp[15]) ? node49660 : 4'b0010;
															assign node49660 = (inp[5]) ? 4'b0110 : 4'b0111;
													assign node49663 = (inp[1]) ? node49667 : node49664;
														assign node49664 = (inp[15]) ? 4'b0011 : 4'b0010;
														assign node49667 = (inp[15]) ? 4'b0011 : 4'b0111;
											assign node49670 = (inp[5]) ? node49696 : node49671;
												assign node49671 = (inp[13]) ? node49683 : node49672;
													assign node49672 = (inp[12]) ? node49678 : node49673;
														assign node49673 = (inp[1]) ? node49675 : 4'b0010;
															assign node49675 = (inp[15]) ? 4'b0011 : 4'b0110;
														assign node49678 = (inp[1]) ? node49680 : 4'b0110;
															assign node49680 = (inp[15]) ? 4'b0110 : 4'b0010;
													assign node49683 = (inp[12]) ? node49691 : node49684;
														assign node49684 = (inp[15]) ? node49688 : node49685;
															assign node49685 = (inp[1]) ? 4'b0011 : 4'b0111;
															assign node49688 = (inp[1]) ? 4'b0111 : 4'b0110;
														assign node49691 = (inp[15]) ? 4'b0010 : node49692;
															assign node49692 = (inp[1]) ? 4'b0110 : 4'b0011;
												assign node49696 = (inp[13]) ? node49708 : node49697;
													assign node49697 = (inp[1]) ? node49701 : node49698;
														assign node49698 = (inp[12]) ? 4'b0111 : 4'b0011;
														assign node49701 = (inp[15]) ? node49705 : node49702;
															assign node49702 = (inp[12]) ? 4'b0010 : 4'b0111;
															assign node49705 = (inp[12]) ? 4'b0111 : 4'b0010;
													assign node49708 = (inp[12]) ? node49716 : node49709;
														assign node49709 = (inp[1]) ? node49713 : node49710;
															assign node49710 = (inp[15]) ? 4'b0110 : 4'b0111;
															assign node49713 = (inp[15]) ? 4'b0111 : 4'b0010;
														assign node49716 = (inp[1]) ? node49720 : node49717;
															assign node49717 = (inp[15]) ? 4'b0011 : 4'b0010;
															assign node49720 = (inp[15]) ? 4'b0011 : 4'b0111;
									assign node49723 = (inp[2]) ? node49823 : node49724;
										assign node49724 = (inp[0]) ? node49760 : node49725;
											assign node49725 = (inp[12]) ? node49745 : node49726;
												assign node49726 = (inp[13]) ? node49732 : node49727;
													assign node49727 = (inp[1]) ? node49729 : 4'b0011;
														assign node49729 = (inp[15]) ? 4'b0010 : 4'b0111;
													assign node49732 = (inp[5]) ? node49738 : node49733;
														assign node49733 = (inp[1]) ? 4'b0111 : node49734;
															assign node49734 = (inp[15]) ? 4'b0110 : 4'b0111;
														assign node49738 = (inp[15]) ? node49742 : node49739;
															assign node49739 = (inp[1]) ? 4'b0010 : 4'b0110;
															assign node49742 = (inp[1]) ? 4'b0110 : 4'b0111;
												assign node49745 = (inp[13]) ? node49753 : node49746;
													assign node49746 = (inp[15]) ? 4'b0111 : node49747;
														assign node49747 = (inp[1]) ? node49749 : 4'b0111;
															assign node49749 = (inp[5]) ? 4'b0011 : 4'b0010;
													assign node49753 = (inp[1]) ? node49757 : node49754;
														assign node49754 = (inp[15]) ? 4'b0011 : 4'b0010;
														assign node49757 = (inp[15]) ? 4'b0011 : 4'b0111;
											assign node49760 = (inp[5]) ? node49788 : node49761;
												assign node49761 = (inp[12]) ? node49775 : node49762;
													assign node49762 = (inp[1]) ? node49768 : node49763;
														assign node49763 = (inp[13]) ? node49765 : 4'b0010;
															assign node49765 = (inp[15]) ? 4'b0110 : 4'b0111;
														assign node49768 = (inp[13]) ? node49772 : node49769;
															assign node49769 = (inp[15]) ? 4'b0011 : 4'b0110;
															assign node49772 = (inp[15]) ? 4'b0111 : 4'b0011;
													assign node49775 = (inp[13]) ? node49781 : node49776;
														assign node49776 = (inp[1]) ? node49778 : 4'b0110;
															assign node49778 = (inp[15]) ? 4'b0110 : 4'b0010;
														assign node49781 = (inp[1]) ? node49785 : node49782;
															assign node49782 = (inp[15]) ? 4'b0010 : 4'b0011;
															assign node49785 = (inp[15]) ? 4'b0010 : 4'b0110;
												assign node49788 = (inp[15]) ? node49812 : node49789;
													assign node49789 = (inp[13]) ? node49797 : node49790;
														assign node49790 = (inp[12]) ? node49794 : node49791;
															assign node49791 = (inp[1]) ? 4'b0111 : 4'b0011;
															assign node49794 = (inp[1]) ? 4'b0010 : 4'b0111;
														assign node49797 = (inp[10]) ? node49805 : node49798;
															assign node49798 = (inp[1]) ? node49802 : node49799;
																assign node49799 = (inp[12]) ? 4'b0010 : 4'b0111;
																assign node49802 = (inp[12]) ? 4'b0111 : 4'b0010;
															assign node49805 = (inp[1]) ? node49809 : node49806;
																assign node49806 = (inp[12]) ? 4'b0010 : 4'b0111;
																assign node49809 = (inp[12]) ? 4'b0111 : 4'b0010;
													assign node49812 = (inp[12]) ? node49820 : node49813;
														assign node49813 = (inp[13]) ? node49817 : node49814;
															assign node49814 = (inp[1]) ? 4'b0010 : 4'b0011;
															assign node49817 = (inp[1]) ? 4'b0111 : 4'b0110;
														assign node49820 = (inp[13]) ? 4'b0011 : 4'b0111;
										assign node49823 = (inp[5]) ? node49875 : node49824;
											assign node49824 = (inp[0]) ? node49852 : node49825;
												assign node49825 = (inp[12]) ? node49841 : node49826;
													assign node49826 = (inp[13]) ? node49834 : node49827;
														assign node49827 = (inp[15]) ? node49831 : node49828;
															assign node49828 = (inp[1]) ? 4'b0110 : 4'b0010;
															assign node49831 = (inp[1]) ? 4'b0011 : 4'b0010;
														assign node49834 = (inp[1]) ? node49838 : node49835;
															assign node49835 = (inp[15]) ? 4'b0111 : 4'b0110;
															assign node49838 = (inp[15]) ? 4'b0110 : 4'b0011;
													assign node49841 = (inp[15]) ? node49849 : node49842;
														assign node49842 = (inp[1]) ? node49846 : node49843;
															assign node49843 = (inp[13]) ? 4'b0011 : 4'b0110;
															assign node49846 = (inp[13]) ? 4'b0110 : 4'b0011;
														assign node49849 = (inp[13]) ? 4'b0010 : 4'b0110;
												assign node49852 = (inp[13]) ? node49864 : node49853;
													assign node49853 = (inp[12]) ? node49859 : node49854;
														assign node49854 = (inp[1]) ? node49856 : 4'b0011;
															assign node49856 = (inp[15]) ? 4'b0010 : 4'b0111;
														assign node49859 = (inp[1]) ? node49861 : 4'b0111;
															assign node49861 = (inp[15]) ? 4'b0111 : 4'b0011;
													assign node49864 = (inp[12]) ? node49872 : node49865;
														assign node49865 = (inp[1]) ? node49869 : node49866;
															assign node49866 = (inp[15]) ? 4'b0111 : 4'b0110;
															assign node49869 = (inp[15]) ? 4'b0110 : 4'b0010;
														assign node49872 = (inp[15]) ? 4'b0011 : 4'b0010;
											assign node49875 = (inp[13]) ? node49889 : node49876;
												assign node49876 = (inp[12]) ? node49882 : node49877;
													assign node49877 = (inp[1]) ? node49879 : 4'b0010;
														assign node49879 = (inp[15]) ? 4'b0011 : 4'b0110;
													assign node49882 = (inp[1]) ? node49884 : 4'b0110;
														assign node49884 = (inp[15]) ? 4'b0110 : node49885;
															assign node49885 = (inp[0]) ? 4'b0011 : 4'b0010;
												assign node49889 = (inp[12]) ? node49903 : node49890;
													assign node49890 = (inp[1]) ? node49898 : node49891;
														assign node49891 = (inp[15]) ? node49895 : node49892;
															assign node49892 = (inp[0]) ? 4'b0110 : 4'b0111;
															assign node49895 = (inp[0]) ? 4'b0111 : 4'b0110;
														assign node49898 = (inp[15]) ? node49900 : 4'b0011;
															assign node49900 = (inp[0]) ? 4'b0110 : 4'b0111;
													assign node49903 = (inp[15]) ? 4'b0010 : node49904;
														assign node49904 = (inp[1]) ? 4'b0110 : 4'b0011;
							assign node49908 = (inp[12]) ? node49964 : node49909;
								assign node49909 = (inp[15]) ? node49957 : node49910;
									assign node49910 = (inp[10]) ? node49934 : node49911;
										assign node49911 = (inp[2]) ? node49923 : node49912;
											assign node49912 = (inp[13]) ? node49918 : node49913;
												assign node49913 = (inp[1]) ? node49915 : 4'b0000;
													assign node49915 = (inp[5]) ? 4'b0001 : 4'b0000;
												assign node49918 = (inp[5]) ? node49920 : 4'b0001;
													assign node49920 = (inp[1]) ? 4'b0000 : 4'b0001;
											assign node49923 = (inp[13]) ? node49929 : node49924;
												assign node49924 = (inp[5]) ? node49926 : 4'b0001;
													assign node49926 = (inp[1]) ? 4'b0000 : 4'b0001;
												assign node49929 = (inp[5]) ? node49931 : 4'b0000;
													assign node49931 = (inp[1]) ? 4'b0001 : 4'b0000;
										assign node49934 = (inp[2]) ? node49946 : node49935;
											assign node49935 = (inp[13]) ? node49941 : node49936;
												assign node49936 = (inp[1]) ? node49938 : 4'b0000;
													assign node49938 = (inp[5]) ? 4'b0001 : 4'b0000;
												assign node49941 = (inp[5]) ? node49943 : 4'b0001;
													assign node49943 = (inp[1]) ? 4'b0000 : 4'b0001;
											assign node49946 = (inp[13]) ? node49952 : node49947;
												assign node49947 = (inp[5]) ? node49949 : 4'b0001;
													assign node49949 = (inp[1]) ? 4'b0000 : 4'b0001;
												assign node49952 = (inp[1]) ? node49954 : 4'b0000;
													assign node49954 = (inp[5]) ? 4'b0001 : 4'b0000;
									assign node49957 = (inp[2]) ? node49961 : node49958;
										assign node49958 = (inp[1]) ? 4'b0101 : 4'b0100;
										assign node49961 = (inp[1]) ? 4'b0100 : 4'b0101;
								assign node49964 = (inp[15]) ? node50076 : node49965;
									assign node49965 = (inp[9]) ? node50029 : node49966;
										assign node49966 = (inp[1]) ? node49974 : node49967;
											assign node49967 = (inp[13]) ? node49971 : node49968;
												assign node49968 = (inp[2]) ? 4'b0101 : 4'b0100;
												assign node49971 = (inp[2]) ? 4'b0100 : 4'b0101;
											assign node49974 = (inp[10]) ? node49990 : node49975;
												assign node49975 = (inp[13]) ? node49983 : node49976;
													assign node49976 = (inp[2]) ? node49980 : node49977;
														assign node49977 = (inp[5]) ? 4'b0100 : 4'b0101;
														assign node49980 = (inp[5]) ? 4'b0101 : 4'b0100;
													assign node49983 = (inp[2]) ? node49987 : node49984;
														assign node49984 = (inp[5]) ? 4'b0101 : 4'b0100;
														assign node49987 = (inp[5]) ? 4'b0100 : 4'b0101;
												assign node49990 = (inp[0]) ? node50006 : node49991;
													assign node49991 = (inp[13]) ? node49999 : node49992;
														assign node49992 = (inp[2]) ? node49996 : node49993;
															assign node49993 = (inp[5]) ? 4'b0100 : 4'b0101;
															assign node49996 = (inp[5]) ? 4'b0101 : 4'b0100;
														assign node49999 = (inp[5]) ? node50003 : node50000;
															assign node50000 = (inp[2]) ? 4'b0101 : 4'b0100;
															assign node50003 = (inp[2]) ? 4'b0100 : 4'b0101;
													assign node50006 = (inp[2]) ? node50014 : node50007;
														assign node50007 = (inp[5]) ? node50011 : node50008;
															assign node50008 = (inp[13]) ? 4'b0100 : 4'b0101;
															assign node50011 = (inp[13]) ? 4'b0101 : 4'b0100;
														assign node50014 = (inp[11]) ? node50022 : node50015;
															assign node50015 = (inp[5]) ? node50019 : node50016;
																assign node50016 = (inp[13]) ? 4'b0101 : 4'b0100;
																assign node50019 = (inp[13]) ? 4'b0100 : 4'b0101;
															assign node50022 = (inp[5]) ? node50026 : node50023;
																assign node50023 = (inp[13]) ? 4'b0101 : 4'b0100;
																assign node50026 = (inp[13]) ? 4'b0100 : 4'b0101;
										assign node50029 = (inp[0]) ? node50053 : node50030;
											assign node50030 = (inp[13]) ? node50042 : node50031;
												assign node50031 = (inp[2]) ? node50037 : node50032;
													assign node50032 = (inp[5]) ? 4'b0100 : node50033;
														assign node50033 = (inp[1]) ? 4'b0101 : 4'b0100;
													assign node50037 = (inp[5]) ? 4'b0101 : node50038;
														assign node50038 = (inp[1]) ? 4'b0100 : 4'b0101;
												assign node50042 = (inp[2]) ? node50048 : node50043;
													assign node50043 = (inp[5]) ? 4'b0101 : node50044;
														assign node50044 = (inp[1]) ? 4'b0100 : 4'b0101;
													assign node50048 = (inp[1]) ? node50050 : 4'b0100;
														assign node50050 = (inp[5]) ? 4'b0100 : 4'b0101;
											assign node50053 = (inp[13]) ? node50065 : node50054;
												assign node50054 = (inp[2]) ? node50060 : node50055;
													assign node50055 = (inp[1]) ? node50057 : 4'b0100;
														assign node50057 = (inp[5]) ? 4'b0100 : 4'b0101;
													assign node50060 = (inp[1]) ? node50062 : 4'b0101;
														assign node50062 = (inp[5]) ? 4'b0101 : 4'b0100;
												assign node50065 = (inp[2]) ? node50071 : node50066;
													assign node50066 = (inp[5]) ? 4'b0101 : node50067;
														assign node50067 = (inp[1]) ? 4'b0100 : 4'b0101;
													assign node50071 = (inp[5]) ? 4'b0100 : node50072;
														assign node50072 = (inp[1]) ? 4'b0101 : 4'b0100;
									assign node50076 = (inp[5]) ? node50080 : node50077;
										assign node50077 = (inp[2]) ? 4'b0001 : 4'b0000;
										assign node50080 = (inp[2]) ? 4'b0000 : 4'b0001;
						assign node50083 = (inp[12]) ? node50769 : node50084;
							assign node50084 = (inp[8]) ? node50492 : node50085;
								assign node50085 = (inp[13]) ? node50307 : node50086;
									assign node50086 = (inp[1]) ? node50204 : node50087;
										assign node50087 = (inp[15]) ? node50181 : node50088;
											assign node50088 = (inp[11]) ? node50134 : node50089;
												assign node50089 = (inp[0]) ? node50113 : node50090;
													assign node50090 = (inp[10]) ? node50100 : node50091;
														assign node50091 = (inp[5]) ? 4'b0101 : node50092;
															assign node50092 = (inp[9]) ? node50096 : node50093;
																assign node50093 = (inp[2]) ? 4'b0101 : 4'b0100;
																assign node50096 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node50100 = (inp[9]) ? node50108 : node50101;
															assign node50101 = (inp[2]) ? node50105 : node50102;
																assign node50102 = (inp[5]) ? 4'b0101 : 4'b0100;
																assign node50105 = (inp[5]) ? 4'b0100 : 4'b0101;
															assign node50108 = (inp[2]) ? 4'b0101 : node50109;
																assign node50109 = (inp[5]) ? 4'b0100 : 4'b0101;
													assign node50113 = (inp[10]) ? node50127 : node50114;
														assign node50114 = (inp[5]) ? node50122 : node50115;
															assign node50115 = (inp[2]) ? node50119 : node50116;
																assign node50116 = (inp[9]) ? 4'b0100 : 4'b0101;
																assign node50119 = (inp[9]) ? 4'b0101 : 4'b0100;
															assign node50122 = (inp[2]) ? node50124 : 4'b0100;
																assign node50124 = (inp[9]) ? 4'b0101 : 4'b0100;
														assign node50127 = (inp[2]) ? node50131 : node50128;
															assign node50128 = (inp[9]) ? 4'b0100 : 4'b0101;
															assign node50131 = (inp[5]) ? 4'b0101 : 4'b0100;
												assign node50134 = (inp[10]) ? node50164 : node50135;
													assign node50135 = (inp[0]) ? node50149 : node50136;
														assign node50136 = (inp[2]) ? node50144 : node50137;
															assign node50137 = (inp[5]) ? node50141 : node50138;
																assign node50138 = (inp[9]) ? 4'b0101 : 4'b0100;
																assign node50141 = (inp[9]) ? 4'b0100 : 4'b0101;
															assign node50144 = (inp[5]) ? 4'b0101 : node50145;
																assign node50145 = (inp[9]) ? 4'b0100 : 4'b0101;
														assign node50149 = (inp[5]) ? node50157 : node50150;
															assign node50150 = (inp[2]) ? node50154 : node50151;
																assign node50151 = (inp[9]) ? 4'b0100 : 4'b0101;
																assign node50154 = (inp[9]) ? 4'b0101 : 4'b0100;
															assign node50157 = (inp[2]) ? node50161 : node50158;
																assign node50158 = (inp[9]) ? 4'b0100 : 4'b0101;
																assign node50161 = (inp[9]) ? 4'b0101 : 4'b0100;
													assign node50164 = (inp[9]) ? node50170 : node50165;
														assign node50165 = (inp[2]) ? 4'b0100 : node50166;
															assign node50166 = (inp[0]) ? 4'b0101 : 4'b0100;
														assign node50170 = (inp[2]) ? node50176 : node50171;
															assign node50171 = (inp[5]) ? 4'b0100 : node50172;
																assign node50172 = (inp[0]) ? 4'b0100 : 4'b0101;
															assign node50176 = (inp[0]) ? 4'b0101 : node50177;
																assign node50177 = (inp[5]) ? 4'b0101 : 4'b0100;
											assign node50181 = (inp[2]) ? node50193 : node50182;
												assign node50182 = (inp[9]) ? node50188 : node50183;
													assign node50183 = (inp[0]) ? node50185 : 4'b0000;
														assign node50185 = (inp[5]) ? 4'b0001 : 4'b0000;
													assign node50188 = (inp[0]) ? node50190 : 4'b0001;
														assign node50190 = (inp[5]) ? 4'b0000 : 4'b0001;
												assign node50193 = (inp[9]) ? node50199 : node50194;
													assign node50194 = (inp[5]) ? node50196 : 4'b0001;
														assign node50196 = (inp[0]) ? 4'b0000 : 4'b0001;
													assign node50199 = (inp[0]) ? node50201 : 4'b0000;
														assign node50201 = (inp[5]) ? 4'b0001 : 4'b0000;
										assign node50204 = (inp[11]) ? node50248 : node50205;
											assign node50205 = (inp[15]) ? node50227 : node50206;
												assign node50206 = (inp[9]) ? node50218 : node50207;
													assign node50207 = (inp[2]) ? node50213 : node50208;
														assign node50208 = (inp[5]) ? node50210 : 4'b0000;
															assign node50210 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node50213 = (inp[0]) ? node50215 : 4'b0001;
															assign node50215 = (inp[5]) ? 4'b0000 : 4'b0001;
													assign node50218 = (inp[2]) ? node50224 : node50219;
														assign node50219 = (inp[0]) ? node50221 : 4'b0001;
															assign node50221 = (inp[5]) ? 4'b0000 : 4'b0001;
														assign node50224 = (inp[0]) ? 4'b0001 : 4'b0000;
												assign node50227 = (inp[2]) ? node50237 : node50228;
													assign node50228 = (inp[9]) ? node50234 : node50229;
														assign node50229 = (inp[5]) ? node50231 : 4'b0001;
															assign node50231 = (inp[0]) ? 4'b0000 : 4'b0001;
														assign node50234 = (inp[0]) ? 4'b0001 : 4'b0000;
													assign node50237 = (inp[9]) ? node50243 : node50238;
														assign node50238 = (inp[5]) ? node50240 : 4'b0000;
															assign node50240 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node50243 = (inp[0]) ? node50245 : 4'b0001;
															assign node50245 = (inp[5]) ? 4'b0000 : 4'b0001;
											assign node50248 = (inp[5]) ? node50264 : node50249;
												assign node50249 = (inp[15]) ? node50257 : node50250;
													assign node50250 = (inp[9]) ? node50254 : node50251;
														assign node50251 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node50254 = (inp[2]) ? 4'b0000 : 4'b0001;
													assign node50257 = (inp[2]) ? node50261 : node50258;
														assign node50258 = (inp[9]) ? 4'b0000 : 4'b0001;
														assign node50261 = (inp[9]) ? 4'b0001 : 4'b0000;
												assign node50264 = (inp[9]) ? node50292 : node50265;
													assign node50265 = (inp[10]) ? node50279 : node50266;
														assign node50266 = (inp[0]) ? node50274 : node50267;
															assign node50267 = (inp[2]) ? node50271 : node50268;
																assign node50268 = (inp[15]) ? 4'b0001 : 4'b0000;
																assign node50271 = (inp[15]) ? 4'b0000 : 4'b0001;
															assign node50274 = (inp[15]) ? 4'b0000 : node50275;
																assign node50275 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node50279 = (inp[0]) ? node50287 : node50280;
															assign node50280 = (inp[2]) ? node50284 : node50281;
																assign node50281 = (inp[15]) ? 4'b0001 : 4'b0000;
																assign node50284 = (inp[15]) ? 4'b0000 : 4'b0001;
															assign node50287 = (inp[2]) ? node50289 : 4'b0001;
																assign node50289 = (inp[15]) ? 4'b0001 : 4'b0000;
													assign node50292 = (inp[2]) ? node50300 : node50293;
														assign node50293 = (inp[0]) ? node50297 : node50294;
															assign node50294 = (inp[15]) ? 4'b0000 : 4'b0001;
															assign node50297 = (inp[15]) ? 4'b0001 : 4'b0000;
														assign node50300 = (inp[15]) ? node50304 : node50301;
															assign node50301 = (inp[0]) ? 4'b0001 : 4'b0000;
															assign node50304 = (inp[0]) ? 4'b0000 : 4'b0001;
									assign node50307 = (inp[15]) ? node50355 : node50308;
										assign node50308 = (inp[1]) ? node50332 : node50309;
											assign node50309 = (inp[2]) ? node50321 : node50310;
												assign node50310 = (inp[9]) ? node50316 : node50311;
													assign node50311 = (inp[5]) ? 4'b0000 : node50312;
														assign node50312 = (inp[0]) ? 4'b0000 : 4'b0001;
													assign node50316 = (inp[0]) ? 4'b0001 : node50317;
														assign node50317 = (inp[5]) ? 4'b0001 : 4'b0000;
												assign node50321 = (inp[9]) ? node50327 : node50322;
													assign node50322 = (inp[0]) ? 4'b0001 : node50323;
														assign node50323 = (inp[5]) ? 4'b0001 : 4'b0000;
													assign node50327 = (inp[0]) ? 4'b0000 : node50328;
														assign node50328 = (inp[5]) ? 4'b0000 : 4'b0001;
											assign node50332 = (inp[9]) ? node50344 : node50333;
												assign node50333 = (inp[2]) ? node50339 : node50334;
													assign node50334 = (inp[5]) ? 4'b0100 : node50335;
														assign node50335 = (inp[0]) ? 4'b0100 : 4'b0101;
													assign node50339 = (inp[5]) ? 4'b0101 : node50340;
														assign node50340 = (inp[0]) ? 4'b0101 : 4'b0100;
												assign node50344 = (inp[2]) ? node50350 : node50345;
													assign node50345 = (inp[0]) ? 4'b0101 : node50346;
														assign node50346 = (inp[5]) ? 4'b0101 : 4'b0100;
													assign node50350 = (inp[5]) ? 4'b0100 : node50351;
														assign node50351 = (inp[0]) ? 4'b0100 : 4'b0101;
										assign node50355 = (inp[10]) ? node50435 : node50356;
											assign node50356 = (inp[0]) ? node50412 : node50357;
												assign node50357 = (inp[11]) ? node50383 : node50358;
													assign node50358 = (inp[1]) ? node50368 : node50359;
														assign node50359 = (inp[9]) ? node50361 : 4'b0101;
															assign node50361 = (inp[2]) ? node50365 : node50362;
																assign node50362 = (inp[5]) ? 4'b0100 : 4'b0101;
																assign node50365 = (inp[5]) ? 4'b0101 : 4'b0100;
														assign node50368 = (inp[2]) ? node50376 : node50369;
															assign node50369 = (inp[9]) ? node50373 : node50370;
																assign node50370 = (inp[5]) ? 4'b0100 : 4'b0101;
																assign node50373 = (inp[5]) ? 4'b0101 : 4'b0100;
															assign node50376 = (inp[5]) ? node50380 : node50377;
																assign node50377 = (inp[9]) ? 4'b0101 : 4'b0100;
																assign node50380 = (inp[9]) ? 4'b0100 : 4'b0101;
													assign node50383 = (inp[1]) ? node50397 : node50384;
														assign node50384 = (inp[2]) ? node50392 : node50385;
															assign node50385 = (inp[5]) ? node50389 : node50386;
																assign node50386 = (inp[9]) ? 4'b0101 : 4'b0100;
																assign node50389 = (inp[9]) ? 4'b0100 : 4'b0101;
															assign node50392 = (inp[9]) ? 4'b0100 : node50393;
																assign node50393 = (inp[5]) ? 4'b0100 : 4'b0101;
														assign node50397 = (inp[2]) ? node50405 : node50398;
															assign node50398 = (inp[9]) ? node50402 : node50399;
																assign node50399 = (inp[5]) ? 4'b0100 : 4'b0101;
																assign node50402 = (inp[5]) ? 4'b0101 : 4'b0100;
															assign node50405 = (inp[5]) ? node50409 : node50406;
																assign node50406 = (inp[9]) ? 4'b0101 : 4'b0100;
																assign node50409 = (inp[9]) ? 4'b0100 : 4'b0101;
												assign node50412 = (inp[9]) ? node50420 : node50413;
													assign node50413 = (inp[1]) ? node50417 : node50414;
														assign node50414 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node50417 = (inp[2]) ? 4'b0101 : 4'b0100;
													assign node50420 = (inp[11]) ? node50428 : node50421;
														assign node50421 = (inp[5]) ? node50423 : 4'b0101;
															assign node50423 = (inp[1]) ? 4'b0101 : node50424;
																assign node50424 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node50428 = (inp[1]) ? node50432 : node50429;
															assign node50429 = (inp[2]) ? 4'b0101 : 4'b0100;
															assign node50432 = (inp[2]) ? 4'b0100 : 4'b0101;
											assign node50435 = (inp[1]) ? node50469 : node50436;
												assign node50436 = (inp[0]) ? node50462 : node50437;
													assign node50437 = (inp[11]) ? node50447 : node50438;
														assign node50438 = (inp[9]) ? 4'b0101 : node50439;
															assign node50439 = (inp[5]) ? node50443 : node50440;
																assign node50440 = (inp[2]) ? 4'b0101 : 4'b0100;
																assign node50443 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node50447 = (inp[5]) ? node50455 : node50448;
															assign node50448 = (inp[2]) ? node50452 : node50449;
																assign node50449 = (inp[9]) ? 4'b0101 : 4'b0100;
																assign node50452 = (inp[9]) ? 4'b0100 : 4'b0101;
															assign node50455 = (inp[9]) ? node50459 : node50456;
																assign node50456 = (inp[2]) ? 4'b0100 : 4'b0101;
																assign node50459 = (inp[2]) ? 4'b0101 : 4'b0100;
													assign node50462 = (inp[2]) ? node50466 : node50463;
														assign node50463 = (inp[9]) ? 4'b0100 : 4'b0101;
														assign node50466 = (inp[9]) ? 4'b0101 : 4'b0100;
												assign node50469 = (inp[2]) ? node50481 : node50470;
													assign node50470 = (inp[9]) ? node50476 : node50471;
														assign node50471 = (inp[5]) ? 4'b0100 : node50472;
															assign node50472 = (inp[0]) ? 4'b0100 : 4'b0101;
														assign node50476 = (inp[0]) ? 4'b0101 : node50477;
															assign node50477 = (inp[5]) ? 4'b0101 : 4'b0100;
													assign node50481 = (inp[9]) ? node50487 : node50482;
														assign node50482 = (inp[0]) ? 4'b0101 : node50483;
															assign node50483 = (inp[5]) ? 4'b0101 : 4'b0100;
														assign node50487 = (inp[5]) ? 4'b0100 : node50488;
															assign node50488 = (inp[0]) ? 4'b0100 : 4'b0101;
								assign node50492 = (inp[9]) ? node50650 : node50493;
									assign node50493 = (inp[11]) ? node50611 : node50494;
										assign node50494 = (inp[15]) ? node50588 : node50495;
											assign node50495 = (inp[0]) ? node50537 : node50496;
												assign node50496 = (inp[10]) ? node50518 : node50497;
													assign node50497 = (inp[13]) ? node50507 : node50498;
														assign node50498 = (inp[1]) ? 4'b0101 : node50499;
															assign node50499 = (inp[2]) ? node50503 : node50500;
																assign node50500 = (inp[5]) ? 4'b0101 : 4'b0100;
																assign node50503 = (inp[5]) ? 4'b0100 : 4'b0101;
														assign node50507 = (inp[2]) ? node50513 : node50508;
															assign node50508 = (inp[1]) ? 4'b0101 : node50509;
																assign node50509 = (inp[5]) ? 4'b0100 : 4'b0101;
															assign node50513 = (inp[5]) ? node50515 : 4'b0100;
																assign node50515 = (inp[1]) ? 4'b0100 : 4'b0101;
													assign node50518 = (inp[2]) ? node50528 : node50519;
														assign node50519 = (inp[13]) ? node50525 : node50520;
															assign node50520 = (inp[5]) ? node50522 : 4'b0100;
																assign node50522 = (inp[1]) ? 4'b0100 : 4'b0101;
															assign node50525 = (inp[1]) ? 4'b0101 : 4'b0100;
														assign node50528 = (inp[13]) ? node50534 : node50529;
															assign node50529 = (inp[1]) ? 4'b0101 : node50530;
																assign node50530 = (inp[5]) ? 4'b0100 : 4'b0101;
															assign node50534 = (inp[1]) ? 4'b0100 : 4'b0101;
												assign node50537 = (inp[10]) ? node50561 : node50538;
													assign node50538 = (inp[5]) ? node50552 : node50539;
														assign node50539 = (inp[1]) ? node50545 : node50540;
															assign node50540 = (inp[2]) ? 4'b0100 : node50541;
																assign node50541 = (inp[13]) ? 4'b0101 : 4'b0100;
															assign node50545 = (inp[2]) ? node50549 : node50546;
																assign node50546 = (inp[13]) ? 4'b0101 : 4'b0100;
																assign node50549 = (inp[13]) ? 4'b0100 : 4'b0101;
														assign node50552 = (inp[2]) ? node50554 : 4'b0100;
															assign node50554 = (inp[1]) ? node50558 : node50555;
																assign node50555 = (inp[13]) ? 4'b0101 : 4'b0100;
																assign node50558 = (inp[13]) ? 4'b0100 : 4'b0101;
													assign node50561 = (inp[1]) ? node50575 : node50562;
														assign node50562 = (inp[13]) ? node50568 : node50563;
															assign node50563 = (inp[2]) ? 4'b0101 : node50564;
																assign node50564 = (inp[5]) ? 4'b0101 : 4'b0100;
															assign node50568 = (inp[2]) ? node50572 : node50569;
																assign node50569 = (inp[5]) ? 4'b0100 : 4'b0101;
																assign node50572 = (inp[5]) ? 4'b0101 : 4'b0100;
														assign node50575 = (inp[5]) ? node50583 : node50576;
															assign node50576 = (inp[13]) ? node50580 : node50577;
																assign node50577 = (inp[2]) ? 4'b0101 : 4'b0100;
																assign node50580 = (inp[2]) ? 4'b0100 : 4'b0101;
															assign node50583 = (inp[13]) ? node50585 : 4'b0100;
																assign node50585 = (inp[2]) ? 4'b0100 : 4'b0101;
											assign node50588 = (inp[5]) ? node50604 : node50589;
												assign node50589 = (inp[0]) ? node50597 : node50590;
													assign node50590 = (inp[2]) ? node50594 : node50591;
														assign node50591 = (inp[1]) ? 4'b0101 : 4'b0100;
														assign node50594 = (inp[1]) ? 4'b0100 : 4'b0101;
													assign node50597 = (inp[2]) ? node50601 : node50598;
														assign node50598 = (inp[1]) ? 4'b0101 : 4'b0100;
														assign node50601 = (inp[1]) ? 4'b0100 : 4'b0101;
												assign node50604 = (inp[2]) ? node50608 : node50605;
													assign node50605 = (inp[1]) ? 4'b0101 : 4'b0100;
													assign node50608 = (inp[1]) ? 4'b0100 : 4'b0101;
										assign node50611 = (inp[1]) ? node50639 : node50612;
											assign node50612 = (inp[2]) ? node50622 : node50613;
												assign node50613 = (inp[15]) ? 4'b0100 : node50614;
													assign node50614 = (inp[13]) ? node50618 : node50615;
														assign node50615 = (inp[5]) ? 4'b0101 : 4'b0100;
														assign node50618 = (inp[5]) ? 4'b0100 : 4'b0101;
												assign node50622 = (inp[15]) ? 4'b0101 : node50623;
													assign node50623 = (inp[0]) ? node50631 : node50624;
														assign node50624 = (inp[13]) ? node50628 : node50625;
															assign node50625 = (inp[5]) ? 4'b0100 : 4'b0101;
															assign node50628 = (inp[5]) ? 4'b0101 : 4'b0100;
														assign node50631 = (inp[5]) ? node50635 : node50632;
															assign node50632 = (inp[13]) ? 4'b0100 : 4'b0101;
															assign node50635 = (inp[13]) ? 4'b0101 : 4'b0100;
											assign node50639 = (inp[2]) ? node50645 : node50640;
												assign node50640 = (inp[13]) ? 4'b0101 : node50641;
													assign node50641 = (inp[15]) ? 4'b0101 : 4'b0100;
												assign node50645 = (inp[15]) ? 4'b0100 : node50646;
													assign node50646 = (inp[13]) ? 4'b0100 : 4'b0101;
									assign node50650 = (inp[5]) ? node50692 : node50651;
										assign node50651 = (inp[15]) ? node50659 : node50652;
											assign node50652 = (inp[2]) ? node50656 : node50653;
												assign node50653 = (inp[13]) ? 4'b0101 : 4'b0100;
												assign node50656 = (inp[13]) ? 4'b0100 : 4'b0101;
											assign node50659 = (inp[10]) ? node50667 : node50660;
												assign node50660 = (inp[2]) ? node50664 : node50661;
													assign node50661 = (inp[1]) ? 4'b0101 : 4'b0100;
													assign node50664 = (inp[1]) ? 4'b0100 : 4'b0101;
												assign node50667 = (inp[0]) ? node50685 : node50668;
													assign node50668 = (inp[13]) ? node50670 : 4'b0100;
														assign node50670 = (inp[11]) ? node50678 : node50671;
															assign node50671 = (inp[1]) ? node50675 : node50672;
																assign node50672 = (inp[2]) ? 4'b0101 : 4'b0100;
																assign node50675 = (inp[2]) ? 4'b0100 : 4'b0101;
															assign node50678 = (inp[1]) ? node50682 : node50679;
																assign node50679 = (inp[2]) ? 4'b0101 : 4'b0100;
																assign node50682 = (inp[2]) ? 4'b0100 : 4'b0101;
													assign node50685 = (inp[2]) ? node50689 : node50686;
														assign node50686 = (inp[1]) ? 4'b0101 : 4'b0100;
														assign node50689 = (inp[1]) ? 4'b0100 : 4'b0101;
										assign node50692 = (inp[11]) ? node50716 : node50693;
											assign node50693 = (inp[1]) ? node50705 : node50694;
												assign node50694 = (inp[2]) ? node50700 : node50695;
													assign node50695 = (inp[15]) ? 4'b0100 : node50696;
														assign node50696 = (inp[13]) ? 4'b0100 : 4'b0101;
													assign node50700 = (inp[13]) ? 4'b0101 : node50701;
														assign node50701 = (inp[15]) ? 4'b0101 : 4'b0100;
												assign node50705 = (inp[2]) ? node50711 : node50706;
													assign node50706 = (inp[13]) ? 4'b0101 : node50707;
														assign node50707 = (inp[15]) ? 4'b0101 : 4'b0100;
													assign node50711 = (inp[15]) ? 4'b0100 : node50712;
														assign node50712 = (inp[13]) ? 4'b0100 : 4'b0101;
											assign node50716 = (inp[15]) ? node50762 : node50717;
												assign node50717 = (inp[1]) ? node50733 : node50718;
													assign node50718 = (inp[0]) ? node50726 : node50719;
														assign node50719 = (inp[2]) ? node50723 : node50720;
															assign node50720 = (inp[13]) ? 4'b0100 : 4'b0101;
															assign node50723 = (inp[13]) ? 4'b0101 : 4'b0100;
														assign node50726 = (inp[2]) ? node50730 : node50727;
															assign node50727 = (inp[13]) ? 4'b0100 : 4'b0101;
															assign node50730 = (inp[13]) ? 4'b0101 : 4'b0100;
													assign node50733 = (inp[0]) ? node50747 : node50734;
														assign node50734 = (inp[10]) ? node50740 : node50735;
															assign node50735 = (inp[2]) ? 4'b0101 : node50736;
																assign node50736 = (inp[13]) ? 4'b0101 : 4'b0100;
															assign node50740 = (inp[2]) ? node50744 : node50741;
																assign node50741 = (inp[13]) ? 4'b0101 : 4'b0100;
																assign node50744 = (inp[13]) ? 4'b0100 : 4'b0101;
														assign node50747 = (inp[10]) ? node50755 : node50748;
															assign node50748 = (inp[2]) ? node50752 : node50749;
																assign node50749 = (inp[13]) ? 4'b0101 : 4'b0100;
																assign node50752 = (inp[13]) ? 4'b0100 : 4'b0101;
															assign node50755 = (inp[13]) ? node50759 : node50756;
																assign node50756 = (inp[2]) ? 4'b0101 : 4'b0100;
																assign node50759 = (inp[2]) ? 4'b0100 : 4'b0101;
												assign node50762 = (inp[1]) ? node50766 : node50763;
													assign node50763 = (inp[2]) ? 4'b0101 : 4'b0100;
													assign node50766 = (inp[2]) ? 4'b0100 : 4'b0101;
							assign node50769 = (inp[8]) ? node51049 : node50770;
								assign node50770 = (inp[13]) ? node50954 : node50771;
									assign node50771 = (inp[1]) ? node50875 : node50772;
										assign node50772 = (inp[15]) ? node50820 : node50773;
											assign node50773 = (inp[5]) ? node50813 : node50774;
												assign node50774 = (inp[10]) ? node50798 : node50775;
													assign node50775 = (inp[2]) ? node50791 : node50776;
														assign node50776 = (inp[11]) ? node50784 : node50777;
															assign node50777 = (inp[0]) ? node50781 : node50778;
																assign node50778 = (inp[9]) ? 4'b0000 : 4'b0001;
																assign node50781 = (inp[9]) ? 4'b0001 : 4'b0000;
															assign node50784 = (inp[9]) ? node50788 : node50785;
																assign node50785 = (inp[0]) ? 4'b0000 : 4'b0001;
																assign node50788 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node50791 = (inp[0]) ? node50795 : node50792;
															assign node50792 = (inp[9]) ? 4'b0001 : 4'b0000;
															assign node50795 = (inp[9]) ? 4'b0000 : 4'b0001;
													assign node50798 = (inp[2]) ? node50806 : node50799;
														assign node50799 = (inp[0]) ? node50803 : node50800;
															assign node50800 = (inp[9]) ? 4'b0000 : 4'b0001;
															assign node50803 = (inp[9]) ? 4'b0001 : 4'b0000;
														assign node50806 = (inp[0]) ? node50810 : node50807;
															assign node50807 = (inp[9]) ? 4'b0001 : 4'b0000;
															assign node50810 = (inp[9]) ? 4'b0000 : 4'b0001;
												assign node50813 = (inp[2]) ? node50817 : node50814;
													assign node50814 = (inp[9]) ? 4'b0001 : 4'b0000;
													assign node50817 = (inp[9]) ? 4'b0000 : 4'b0001;
											assign node50820 = (inp[11]) ? node50844 : node50821;
												assign node50821 = (inp[9]) ? node50833 : node50822;
													assign node50822 = (inp[2]) ? node50828 : node50823;
														assign node50823 = (inp[0]) ? 4'b0100 : node50824;
															assign node50824 = (inp[5]) ? 4'b0100 : 4'b0101;
														assign node50828 = (inp[5]) ? 4'b0101 : node50829;
															assign node50829 = (inp[0]) ? 4'b0101 : 4'b0100;
													assign node50833 = (inp[2]) ? node50839 : node50834;
														assign node50834 = (inp[5]) ? 4'b0101 : node50835;
															assign node50835 = (inp[0]) ? 4'b0101 : 4'b0100;
														assign node50839 = (inp[0]) ? 4'b0100 : node50840;
															assign node50840 = (inp[5]) ? 4'b0100 : 4'b0101;
												assign node50844 = (inp[10]) ? node50860 : node50845;
													assign node50845 = (inp[9]) ? node50853 : node50846;
														assign node50846 = (inp[2]) ? node50848 : 4'b0100;
															assign node50848 = (inp[5]) ? 4'b0101 : node50849;
																assign node50849 = (inp[0]) ? 4'b0101 : 4'b0100;
														assign node50853 = (inp[2]) ? node50855 : 4'b0101;
															assign node50855 = (inp[0]) ? 4'b0100 : node50856;
																assign node50856 = (inp[5]) ? 4'b0100 : 4'b0101;
													assign node50860 = (inp[2]) ? node50870 : node50861;
														assign node50861 = (inp[0]) ? node50867 : node50862;
															assign node50862 = (inp[9]) ? node50864 : 4'b0101;
																assign node50864 = (inp[5]) ? 4'b0101 : 4'b0100;
															assign node50867 = (inp[9]) ? 4'b0101 : 4'b0100;
														assign node50870 = (inp[9]) ? 4'b0100 : node50871;
															assign node50871 = (inp[5]) ? 4'b0101 : 4'b0100;
										assign node50875 = (inp[9]) ? node50931 : node50876;
											assign node50876 = (inp[11]) ? node50900 : node50877;
												assign node50877 = (inp[15]) ? node50889 : node50878;
													assign node50878 = (inp[2]) ? node50884 : node50879;
														assign node50879 = (inp[5]) ? 4'b0101 : node50880;
															assign node50880 = (inp[0]) ? 4'b0101 : 4'b0100;
														assign node50884 = (inp[5]) ? 4'b0100 : node50885;
															assign node50885 = (inp[0]) ? 4'b0100 : 4'b0101;
													assign node50889 = (inp[2]) ? node50895 : node50890;
														assign node50890 = (inp[0]) ? 4'b0100 : node50891;
															assign node50891 = (inp[5]) ? 4'b0100 : 4'b0101;
														assign node50895 = (inp[0]) ? 4'b0101 : node50896;
															assign node50896 = (inp[5]) ? 4'b0101 : 4'b0100;
												assign node50900 = (inp[5]) ? node50916 : node50901;
													assign node50901 = (inp[15]) ? node50909 : node50902;
														assign node50902 = (inp[0]) ? node50906 : node50903;
															assign node50903 = (inp[2]) ? 4'b0101 : 4'b0100;
															assign node50906 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node50909 = (inp[0]) ? node50913 : node50910;
															assign node50910 = (inp[2]) ? 4'b0100 : 4'b0101;
															assign node50913 = (inp[2]) ? 4'b0101 : 4'b0100;
													assign node50916 = (inp[0]) ? node50924 : node50917;
														assign node50917 = (inp[15]) ? node50921 : node50918;
															assign node50918 = (inp[2]) ? 4'b0100 : 4'b0101;
															assign node50921 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node50924 = (inp[2]) ? node50928 : node50925;
															assign node50925 = (inp[15]) ? 4'b0100 : 4'b0101;
															assign node50928 = (inp[15]) ? 4'b0101 : 4'b0100;
											assign node50931 = (inp[15]) ? node50943 : node50932;
												assign node50932 = (inp[2]) ? node50938 : node50933;
													assign node50933 = (inp[0]) ? 4'b0100 : node50934;
														assign node50934 = (inp[5]) ? 4'b0100 : 4'b0101;
													assign node50938 = (inp[0]) ? 4'b0101 : node50939;
														assign node50939 = (inp[5]) ? 4'b0101 : 4'b0100;
												assign node50943 = (inp[2]) ? node50949 : node50944;
													assign node50944 = (inp[5]) ? 4'b0101 : node50945;
														assign node50945 = (inp[0]) ? 4'b0101 : 4'b0100;
													assign node50949 = (inp[5]) ? 4'b0100 : node50950;
														assign node50950 = (inp[0]) ? 4'b0100 : 4'b0101;
									assign node50954 = (inp[1]) ? node51026 : node50955;
										assign node50955 = (inp[15]) ? node50979 : node50956;
											assign node50956 = (inp[9]) ? node50968 : node50957;
												assign node50957 = (inp[2]) ? node50963 : node50958;
													assign node50958 = (inp[5]) ? node50960 : 4'b0101;
														assign node50960 = (inp[0]) ? 4'b0100 : 4'b0101;
													assign node50963 = (inp[5]) ? node50965 : 4'b0100;
														assign node50965 = (inp[0]) ? 4'b0101 : 4'b0100;
												assign node50968 = (inp[2]) ? node50974 : node50969;
													assign node50969 = (inp[0]) ? node50971 : 4'b0100;
														assign node50971 = (inp[5]) ? 4'b0101 : 4'b0100;
													assign node50974 = (inp[5]) ? node50976 : 4'b0101;
														assign node50976 = (inp[0]) ? 4'b0100 : 4'b0101;
											assign node50979 = (inp[11]) ? node50999 : node50980;
												assign node50980 = (inp[2]) ? node50992 : node50981;
													assign node50981 = (inp[9]) ? node50987 : node50982;
														assign node50982 = (inp[5]) ? 4'b0000 : node50983;
															assign node50983 = (inp[0]) ? 4'b0000 : 4'b0001;
														assign node50987 = (inp[0]) ? 4'b0001 : node50988;
															assign node50988 = (inp[5]) ? 4'b0001 : 4'b0000;
													assign node50992 = (inp[9]) ? 4'b0000 : node50993;
														assign node50993 = (inp[5]) ? 4'b0001 : node50994;
															assign node50994 = (inp[0]) ? 4'b0001 : 4'b0000;
												assign node50999 = (inp[0]) ? node51019 : node51000;
													assign node51000 = (inp[5]) ? node51008 : node51001;
														assign node51001 = (inp[9]) ? node51005 : node51002;
															assign node51002 = (inp[2]) ? 4'b0000 : 4'b0001;
															assign node51005 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node51008 = (inp[10]) ? node51014 : node51009;
															assign node51009 = (inp[2]) ? 4'b0001 : node51010;
																assign node51010 = (inp[9]) ? 4'b0001 : 4'b0000;
															assign node51014 = (inp[9]) ? node51016 : 4'b0001;
																assign node51016 = (inp[2]) ? 4'b0000 : 4'b0001;
													assign node51019 = (inp[9]) ? node51023 : node51020;
														assign node51020 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node51023 = (inp[2]) ? 4'b0000 : 4'b0001;
										assign node51026 = (inp[2]) ? node51038 : node51027;
											assign node51027 = (inp[9]) ? node51033 : node51028;
												assign node51028 = (inp[0]) ? 4'b0000 : node51029;
													assign node51029 = (inp[5]) ? 4'b0000 : 4'b0001;
												assign node51033 = (inp[0]) ? 4'b0001 : node51034;
													assign node51034 = (inp[5]) ? 4'b0001 : 4'b0000;
											assign node51038 = (inp[9]) ? node51044 : node51039;
												assign node51039 = (inp[5]) ? 4'b0001 : node51040;
													assign node51040 = (inp[0]) ? 4'b0001 : 4'b0000;
												assign node51044 = (inp[5]) ? 4'b0000 : node51045;
													assign node51045 = (inp[0]) ? 4'b0000 : 4'b0001;
								assign node51049 = (inp[2]) ? node51063 : node51050;
									assign node51050 = (inp[15]) ? 4'b0001 : node51051;
										assign node51051 = (inp[13]) ? node51057 : node51052;
											assign node51052 = (inp[5]) ? 4'b0000 : node51053;
												assign node51053 = (inp[1]) ? 4'b0000 : 4'b0001;
											assign node51057 = (inp[1]) ? 4'b0001 : node51058;
												assign node51058 = (inp[5]) ? 4'b0001 : 4'b0000;
									assign node51063 = (inp[15]) ? 4'b0000 : node51064;
										assign node51064 = (inp[13]) ? node51070 : node51065;
											assign node51065 = (inp[1]) ? 4'b0001 : node51066;
												assign node51066 = (inp[5]) ? 4'b0001 : 4'b0000;
											assign node51070 = (inp[1]) ? 4'b0000 : node51071;
												assign node51071 = (inp[5]) ? 4'b0000 : 4'b0001;
				assign node51076 = (inp[7]) ? node53144 : node51077;
					assign node51077 = (inp[8]) ? node52781 : node51078;
						assign node51078 = (inp[11]) ? node51832 : node51079;
							assign node51079 = (inp[1]) ? node51411 : node51080;
								assign node51080 = (inp[13]) ? node51242 : node51081;
									assign node51081 = (inp[15]) ? node51165 : node51082;
										assign node51082 = (inp[3]) ? node51142 : node51083;
											assign node51083 = (inp[2]) ? node51121 : node51084;
												assign node51084 = (inp[10]) ? node51104 : node51085;
													assign node51085 = (inp[9]) ? node51093 : node51086;
														assign node51086 = (inp[5]) ? 4'b0011 : node51087;
															assign node51087 = (inp[12]) ? node51089 : 4'b0010;
																assign node51089 = (inp[0]) ? 4'b0011 : 4'b0010;
														assign node51093 = (inp[5]) ? node51099 : node51094;
															assign node51094 = (inp[12]) ? node51096 : 4'b0011;
																assign node51096 = (inp[0]) ? 4'b0010 : 4'b0011;
															assign node51099 = (inp[12]) ? node51101 : 4'b0010;
																assign node51101 = (inp[0]) ? 4'b0011 : 4'b0010;
													assign node51104 = (inp[0]) ? node51112 : node51105;
														assign node51105 = (inp[5]) ? node51109 : node51106;
															assign node51106 = (inp[9]) ? 4'b0011 : 4'b0010;
															assign node51109 = (inp[9]) ? 4'b0010 : 4'b0011;
														assign node51112 = (inp[12]) ? 4'b0010 : node51113;
															assign node51113 = (inp[9]) ? node51117 : node51114;
																assign node51114 = (inp[5]) ? 4'b0011 : 4'b0010;
																assign node51117 = (inp[5]) ? 4'b0010 : 4'b0011;
												assign node51121 = (inp[5]) ? node51133 : node51122;
													assign node51122 = (inp[9]) ? node51128 : node51123;
														assign node51123 = (inp[0]) ? node51125 : 4'b0010;
															assign node51125 = (inp[12]) ? 4'b0011 : 4'b0010;
														assign node51128 = (inp[0]) ? node51130 : 4'b0011;
															assign node51130 = (inp[12]) ? 4'b0010 : 4'b0011;
													assign node51133 = (inp[9]) ? node51139 : node51134;
														assign node51134 = (inp[0]) ? node51136 : 4'b0011;
															assign node51136 = (inp[12]) ? 4'b0010 : 4'b0011;
														assign node51139 = (inp[12]) ? 4'b0011 : 4'b0010;
											assign node51142 = (inp[0]) ? node51150 : node51143;
												assign node51143 = (inp[5]) ? node51147 : node51144;
													assign node51144 = (inp[9]) ? 4'b0011 : 4'b0010;
													assign node51147 = (inp[9]) ? 4'b0010 : 4'b0011;
												assign node51150 = (inp[5]) ? node51158 : node51151;
													assign node51151 = (inp[12]) ? node51155 : node51152;
														assign node51152 = (inp[9]) ? 4'b0010 : 4'b0011;
														assign node51155 = (inp[9]) ? 4'b0011 : 4'b0010;
													assign node51158 = (inp[9]) ? node51162 : node51159;
														assign node51159 = (inp[12]) ? 4'b0011 : 4'b0010;
														assign node51162 = (inp[12]) ? 4'b0010 : 4'b0011;
										assign node51165 = (inp[12]) ? node51189 : node51166;
											assign node51166 = (inp[9]) ? node51178 : node51167;
												assign node51167 = (inp[5]) ? node51173 : node51168;
													assign node51168 = (inp[0]) ? node51170 : 4'b0110;
														assign node51170 = (inp[3]) ? 4'b0111 : 4'b0110;
													assign node51173 = (inp[0]) ? node51175 : 4'b0111;
														assign node51175 = (inp[3]) ? 4'b0110 : 4'b0111;
												assign node51178 = (inp[5]) ? node51184 : node51179;
													assign node51179 = (inp[0]) ? node51181 : 4'b0111;
														assign node51181 = (inp[3]) ? 4'b0110 : 4'b0111;
													assign node51184 = (inp[3]) ? node51186 : 4'b0110;
														assign node51186 = (inp[0]) ? 4'b0111 : 4'b0110;
											assign node51189 = (inp[3]) ? node51219 : node51190;
												assign node51190 = (inp[5]) ? node51198 : node51191;
													assign node51191 = (inp[0]) ? node51195 : node51192;
														assign node51192 = (inp[9]) ? 4'b0111 : 4'b0110;
														assign node51195 = (inp[9]) ? 4'b0110 : 4'b0111;
													assign node51198 = (inp[10]) ? node51206 : node51199;
														assign node51199 = (inp[0]) ? node51203 : node51200;
															assign node51200 = (inp[9]) ? 4'b0110 : 4'b0111;
															assign node51203 = (inp[9]) ? 4'b0111 : 4'b0110;
														assign node51206 = (inp[2]) ? node51212 : node51207;
															assign node51207 = (inp[0]) ? 4'b0111 : node51208;
																assign node51208 = (inp[9]) ? 4'b0110 : 4'b0111;
															assign node51212 = (inp[9]) ? node51216 : node51213;
																assign node51213 = (inp[0]) ? 4'b0110 : 4'b0111;
																assign node51216 = (inp[0]) ? 4'b0111 : 4'b0110;
												assign node51219 = (inp[2]) ? node51227 : node51220;
													assign node51220 = (inp[5]) ? node51224 : node51221;
														assign node51221 = (inp[9]) ? 4'b0111 : 4'b0110;
														assign node51224 = (inp[9]) ? 4'b0110 : 4'b0111;
													assign node51227 = (inp[10]) ? node51235 : node51228;
														assign node51228 = (inp[5]) ? node51232 : node51229;
															assign node51229 = (inp[9]) ? 4'b0111 : 4'b0110;
															assign node51232 = (inp[9]) ? 4'b0110 : 4'b0111;
														assign node51235 = (inp[9]) ? node51239 : node51236;
															assign node51236 = (inp[5]) ? 4'b0111 : 4'b0110;
															assign node51239 = (inp[5]) ? 4'b0110 : 4'b0111;
									assign node51242 = (inp[15]) ? node51332 : node51243;
										assign node51243 = (inp[12]) ? node51251 : node51244;
											assign node51244 = (inp[5]) ? node51248 : node51245;
												assign node51245 = (inp[9]) ? 4'b0111 : 4'b0110;
												assign node51248 = (inp[9]) ? 4'b0110 : 4'b0111;
											assign node51251 = (inp[3]) ? node51305 : node51252;
												assign node51252 = (inp[2]) ? node51276 : node51253;
													assign node51253 = (inp[5]) ? node51269 : node51254;
														assign node51254 = (inp[10]) ? node51262 : node51255;
															assign node51255 = (inp[9]) ? node51259 : node51256;
																assign node51256 = (inp[0]) ? 4'b0111 : 4'b0110;
																assign node51259 = (inp[0]) ? 4'b0110 : 4'b0111;
															assign node51262 = (inp[9]) ? node51266 : node51263;
																assign node51263 = (inp[0]) ? 4'b0111 : 4'b0110;
																assign node51266 = (inp[0]) ? 4'b0110 : 4'b0111;
														assign node51269 = (inp[9]) ? node51273 : node51270;
															assign node51270 = (inp[0]) ? 4'b0110 : 4'b0111;
															assign node51273 = (inp[0]) ? 4'b0111 : 4'b0110;
													assign node51276 = (inp[10]) ? node51292 : node51277;
														assign node51277 = (inp[0]) ? node51285 : node51278;
															assign node51278 = (inp[5]) ? node51282 : node51279;
																assign node51279 = (inp[9]) ? 4'b0111 : 4'b0110;
																assign node51282 = (inp[9]) ? 4'b0110 : 4'b0111;
															assign node51285 = (inp[5]) ? node51289 : node51286;
																assign node51286 = (inp[9]) ? 4'b0110 : 4'b0111;
																assign node51289 = (inp[9]) ? 4'b0111 : 4'b0110;
														assign node51292 = (inp[9]) ? node51300 : node51293;
															assign node51293 = (inp[0]) ? node51297 : node51294;
																assign node51294 = (inp[5]) ? 4'b0111 : 4'b0110;
																assign node51297 = (inp[5]) ? 4'b0110 : 4'b0111;
															assign node51300 = (inp[0]) ? node51302 : 4'b0110;
																assign node51302 = (inp[5]) ? 4'b0111 : 4'b0110;
												assign node51305 = (inp[9]) ? node51325 : node51306;
													assign node51306 = (inp[2]) ? node51320 : node51307;
														assign node51307 = (inp[10]) ? node51313 : node51308;
															assign node51308 = (inp[5]) ? 4'b0110 : node51309;
																assign node51309 = (inp[0]) ? 4'b0110 : 4'b0111;
															assign node51313 = (inp[5]) ? node51317 : node51314;
																assign node51314 = (inp[0]) ? 4'b0110 : 4'b0111;
																assign node51317 = (inp[0]) ? 4'b0111 : 4'b0110;
														assign node51320 = (inp[10]) ? 4'b0110 : node51321;
															assign node51321 = (inp[0]) ? 4'b0111 : 4'b0110;
													assign node51325 = (inp[5]) ? node51329 : node51326;
														assign node51326 = (inp[0]) ? 4'b0111 : 4'b0110;
														assign node51329 = (inp[0]) ? 4'b0110 : 4'b0111;
										assign node51332 = (inp[12]) ? node51380 : node51333;
											assign node51333 = (inp[3]) ? node51365 : node51334;
												assign node51334 = (inp[10]) ? node51350 : node51335;
													assign node51335 = (inp[0]) ? node51343 : node51336;
														assign node51336 = (inp[9]) ? node51340 : node51337;
															assign node51337 = (inp[5]) ? 4'b0010 : 4'b0011;
															assign node51340 = (inp[5]) ? 4'b0011 : 4'b0010;
														assign node51343 = (inp[5]) ? node51347 : node51344;
															assign node51344 = (inp[9]) ? 4'b0011 : 4'b0010;
															assign node51347 = (inp[9]) ? 4'b0010 : 4'b0011;
													assign node51350 = (inp[9]) ? node51358 : node51351;
														assign node51351 = (inp[5]) ? node51355 : node51352;
															assign node51352 = (inp[0]) ? 4'b0010 : 4'b0011;
															assign node51355 = (inp[0]) ? 4'b0011 : 4'b0010;
														assign node51358 = (inp[0]) ? node51362 : node51359;
															assign node51359 = (inp[5]) ? 4'b0011 : 4'b0010;
															assign node51362 = (inp[5]) ? 4'b0010 : 4'b0011;
												assign node51365 = (inp[9]) ? node51373 : node51366;
													assign node51366 = (inp[0]) ? node51370 : node51367;
														assign node51367 = (inp[5]) ? 4'b0011 : 4'b0010;
														assign node51370 = (inp[5]) ? 4'b0010 : 4'b0011;
													assign node51373 = (inp[0]) ? node51377 : node51374;
														assign node51374 = (inp[5]) ? 4'b0010 : 4'b0011;
														assign node51377 = (inp[5]) ? 4'b0011 : 4'b0010;
											assign node51380 = (inp[2]) ? node51388 : node51381;
												assign node51381 = (inp[5]) ? node51385 : node51382;
													assign node51382 = (inp[9]) ? 4'b0011 : 4'b0010;
													assign node51385 = (inp[9]) ? 4'b0010 : 4'b0011;
												assign node51388 = (inp[0]) ? node51396 : node51389;
													assign node51389 = (inp[9]) ? node51393 : node51390;
														assign node51390 = (inp[5]) ? 4'b0011 : 4'b0010;
														assign node51393 = (inp[5]) ? 4'b0010 : 4'b0011;
													assign node51396 = (inp[3]) ? node51404 : node51397;
														assign node51397 = (inp[5]) ? node51401 : node51398;
															assign node51398 = (inp[9]) ? 4'b0011 : 4'b0010;
															assign node51401 = (inp[9]) ? 4'b0010 : 4'b0011;
														assign node51404 = (inp[9]) ? node51408 : node51405;
															assign node51405 = (inp[5]) ? 4'b0011 : 4'b0010;
															assign node51408 = (inp[5]) ? 4'b0010 : 4'b0011;
								assign node51411 = (inp[13]) ? node51647 : node51412;
									assign node51412 = (inp[15]) ? node51506 : node51413;
										assign node51413 = (inp[12]) ? node51421 : node51414;
											assign node51414 = (inp[9]) ? node51418 : node51415;
												assign node51415 = (inp[5]) ? 4'b0011 : 4'b0010;
												assign node51418 = (inp[5]) ? 4'b0010 : 4'b0011;
											assign node51421 = (inp[0]) ? node51461 : node51422;
												assign node51422 = (inp[3]) ? node51446 : node51423;
													assign node51423 = (inp[10]) ? node51431 : node51424;
														assign node51424 = (inp[5]) ? node51428 : node51425;
															assign node51425 = (inp[9]) ? 4'b0010 : 4'b0011;
															assign node51428 = (inp[9]) ? 4'b0011 : 4'b0010;
														assign node51431 = (inp[2]) ? node51439 : node51432;
															assign node51432 = (inp[5]) ? node51436 : node51433;
																assign node51433 = (inp[9]) ? 4'b0010 : 4'b0011;
																assign node51436 = (inp[9]) ? 4'b0011 : 4'b0010;
															assign node51439 = (inp[9]) ? node51443 : node51440;
																assign node51440 = (inp[5]) ? 4'b0010 : 4'b0011;
																assign node51443 = (inp[5]) ? 4'b0011 : 4'b0010;
													assign node51446 = (inp[2]) ? node51454 : node51447;
														assign node51447 = (inp[5]) ? node51451 : node51448;
															assign node51448 = (inp[9]) ? 4'b0011 : 4'b0010;
															assign node51451 = (inp[9]) ? 4'b0010 : 4'b0011;
														assign node51454 = (inp[9]) ? node51458 : node51455;
															assign node51455 = (inp[5]) ? 4'b0011 : 4'b0010;
															assign node51458 = (inp[5]) ? 4'b0010 : 4'b0011;
												assign node51461 = (inp[2]) ? node51489 : node51462;
													assign node51462 = (inp[10]) ? node51476 : node51463;
														assign node51463 = (inp[9]) ? node51469 : node51464;
															assign node51464 = (inp[3]) ? 4'b0010 : node51465;
																assign node51465 = (inp[5]) ? 4'b0011 : 4'b0010;
															assign node51469 = (inp[3]) ? node51473 : node51470;
																assign node51470 = (inp[5]) ? 4'b0010 : 4'b0011;
																assign node51473 = (inp[5]) ? 4'b0011 : 4'b0010;
														assign node51476 = (inp[9]) ? node51484 : node51477;
															assign node51477 = (inp[3]) ? node51481 : node51478;
																assign node51478 = (inp[5]) ? 4'b0011 : 4'b0010;
																assign node51481 = (inp[5]) ? 4'b0010 : 4'b0011;
															assign node51484 = (inp[5]) ? node51486 : 4'b0011;
																assign node51486 = (inp[3]) ? 4'b0011 : 4'b0010;
													assign node51489 = (inp[9]) ? node51497 : node51490;
														assign node51490 = (inp[5]) ? node51494 : node51491;
															assign node51491 = (inp[3]) ? 4'b0011 : 4'b0010;
															assign node51494 = (inp[3]) ? 4'b0010 : 4'b0011;
														assign node51497 = (inp[10]) ? 4'b0010 : node51498;
															assign node51498 = (inp[3]) ? node51502 : node51499;
																assign node51499 = (inp[5]) ? 4'b0010 : 4'b0011;
																assign node51502 = (inp[5]) ? 4'b0011 : 4'b0010;
										assign node51506 = (inp[2]) ? node51578 : node51507;
											assign node51507 = (inp[10]) ? node51543 : node51508;
												assign node51508 = (inp[9]) ? node51524 : node51509;
													assign node51509 = (inp[5]) ? node51515 : node51510;
														assign node51510 = (inp[12]) ? 4'b0110 : node51511;
															assign node51511 = (inp[0]) ? 4'b0111 : 4'b0110;
														assign node51515 = (inp[12]) ? 4'b0111 : node51516;
															assign node51516 = (inp[0]) ? node51520 : node51517;
																assign node51517 = (inp[3]) ? 4'b0110 : 4'b0111;
																assign node51520 = (inp[3]) ? 4'b0111 : 4'b0110;
													assign node51524 = (inp[5]) ? node51534 : node51525;
														assign node51525 = (inp[12]) ? 4'b0111 : node51526;
															assign node51526 = (inp[3]) ? node51530 : node51527;
																assign node51527 = (inp[0]) ? 4'b0110 : 4'b0111;
																assign node51530 = (inp[0]) ? 4'b0111 : 4'b0110;
														assign node51534 = (inp[12]) ? 4'b0110 : node51535;
															assign node51535 = (inp[0]) ? node51539 : node51536;
																assign node51536 = (inp[3]) ? 4'b0111 : 4'b0110;
																assign node51539 = (inp[3]) ? 4'b0110 : 4'b0111;
												assign node51543 = (inp[5]) ? node51561 : node51544;
													assign node51544 = (inp[9]) ? node51554 : node51545;
														assign node51545 = (inp[12]) ? 4'b0110 : node51546;
															assign node51546 = (inp[3]) ? node51550 : node51547;
																assign node51547 = (inp[0]) ? 4'b0111 : 4'b0110;
																assign node51550 = (inp[0]) ? 4'b0110 : 4'b0111;
														assign node51554 = (inp[12]) ? 4'b0111 : node51555;
															assign node51555 = (inp[0]) ? node51557 : 4'b0110;
																assign node51557 = (inp[3]) ? 4'b0111 : 4'b0110;
													assign node51561 = (inp[9]) ? node51569 : node51562;
														assign node51562 = (inp[12]) ? 4'b0111 : node51563;
															assign node51563 = (inp[0]) ? 4'b0110 : node51564;
																assign node51564 = (inp[3]) ? 4'b0110 : 4'b0111;
														assign node51569 = (inp[12]) ? 4'b0110 : node51570;
															assign node51570 = (inp[0]) ? node51574 : node51571;
																assign node51571 = (inp[3]) ? 4'b0111 : 4'b0110;
																assign node51574 = (inp[3]) ? 4'b0110 : 4'b0111;
											assign node51578 = (inp[12]) ? node51632 : node51579;
												assign node51579 = (inp[0]) ? node51605 : node51580;
													assign node51580 = (inp[10]) ? node51590 : node51581;
														assign node51581 = (inp[3]) ? node51583 : 4'b0111;
															assign node51583 = (inp[9]) ? node51587 : node51584;
																assign node51584 = (inp[5]) ? 4'b0110 : 4'b0111;
																assign node51587 = (inp[5]) ? 4'b0111 : 4'b0110;
														assign node51590 = (inp[5]) ? node51598 : node51591;
															assign node51591 = (inp[3]) ? node51595 : node51592;
																assign node51592 = (inp[9]) ? 4'b0111 : 4'b0110;
																assign node51595 = (inp[9]) ? 4'b0110 : 4'b0111;
															assign node51598 = (inp[3]) ? node51602 : node51599;
																assign node51599 = (inp[9]) ? 4'b0110 : 4'b0111;
																assign node51602 = (inp[9]) ? 4'b0111 : 4'b0110;
													assign node51605 = (inp[10]) ? node51619 : node51606;
														assign node51606 = (inp[3]) ? node51614 : node51607;
															assign node51607 = (inp[9]) ? node51611 : node51608;
																assign node51608 = (inp[5]) ? 4'b0110 : 4'b0111;
																assign node51611 = (inp[5]) ? 4'b0111 : 4'b0110;
															assign node51614 = (inp[5]) ? node51616 : 4'b0110;
																assign node51616 = (inp[9]) ? 4'b0110 : 4'b0111;
														assign node51619 = (inp[5]) ? node51625 : node51620;
															assign node51620 = (inp[3]) ? 4'b0111 : node51621;
																assign node51621 = (inp[9]) ? 4'b0110 : 4'b0111;
															assign node51625 = (inp[9]) ? node51629 : node51626;
																assign node51626 = (inp[3]) ? 4'b0111 : 4'b0110;
																assign node51629 = (inp[3]) ? 4'b0110 : 4'b0111;
												assign node51632 = (inp[0]) ? node51640 : node51633;
													assign node51633 = (inp[9]) ? node51637 : node51634;
														assign node51634 = (inp[5]) ? 4'b0111 : 4'b0110;
														assign node51637 = (inp[5]) ? 4'b0110 : 4'b0111;
													assign node51640 = (inp[5]) ? node51644 : node51641;
														assign node51641 = (inp[9]) ? 4'b0111 : 4'b0110;
														assign node51644 = (inp[9]) ? 4'b0110 : 4'b0111;
									assign node51647 = (inp[15]) ? node51709 : node51648;
										assign node51648 = (inp[5]) ? node51684 : node51649;
											assign node51649 = (inp[9]) ? node51667 : node51650;
												assign node51650 = (inp[0]) ? 4'b0110 : node51651;
													assign node51651 = (inp[10]) ? node51659 : node51652;
														assign node51652 = (inp[3]) ? node51656 : node51653;
															assign node51653 = (inp[12]) ? 4'b0111 : 4'b0110;
															assign node51656 = (inp[12]) ? 4'b0110 : 4'b0111;
														assign node51659 = (inp[12]) ? node51663 : node51660;
															assign node51660 = (inp[3]) ? 4'b0111 : 4'b0110;
															assign node51663 = (inp[3]) ? 4'b0110 : 4'b0111;
												assign node51667 = (inp[0]) ? 4'b0111 : node51668;
													assign node51668 = (inp[2]) ? node51676 : node51669;
														assign node51669 = (inp[3]) ? node51673 : node51670;
															assign node51670 = (inp[12]) ? 4'b0110 : 4'b0111;
															assign node51673 = (inp[12]) ? 4'b0111 : 4'b0110;
														assign node51676 = (inp[12]) ? node51680 : node51677;
															assign node51677 = (inp[3]) ? 4'b0110 : 4'b0111;
															assign node51680 = (inp[3]) ? 4'b0111 : 4'b0110;
											assign node51684 = (inp[9]) ? node51694 : node51685;
												assign node51685 = (inp[0]) ? 4'b0111 : node51686;
													assign node51686 = (inp[12]) ? node51690 : node51687;
														assign node51687 = (inp[3]) ? 4'b0110 : 4'b0111;
														assign node51690 = (inp[3]) ? 4'b0111 : 4'b0110;
												assign node51694 = (inp[0]) ? 4'b0110 : node51695;
													assign node51695 = (inp[10]) ? node51701 : node51696;
														assign node51696 = (inp[12]) ? node51698 : 4'b0111;
															assign node51698 = (inp[3]) ? 4'b0110 : 4'b0111;
														assign node51701 = (inp[12]) ? node51705 : node51702;
															assign node51702 = (inp[3]) ? 4'b0111 : 4'b0110;
															assign node51705 = (inp[3]) ? 4'b0110 : 4'b0111;
										assign node51709 = (inp[10]) ? node51781 : node51710;
											assign node51710 = (inp[0]) ? node51766 : node51711;
												assign node51711 = (inp[5]) ? node51735 : node51712;
													assign node51712 = (inp[12]) ? node51728 : node51713;
														assign node51713 = (inp[2]) ? node51721 : node51714;
															assign node51714 = (inp[9]) ? node51718 : node51715;
																assign node51715 = (inp[3]) ? 4'b0011 : 4'b0010;
																assign node51718 = (inp[3]) ? 4'b0010 : 4'b0011;
															assign node51721 = (inp[3]) ? node51725 : node51722;
																assign node51722 = (inp[9]) ? 4'b0011 : 4'b0010;
																assign node51725 = (inp[9]) ? 4'b0010 : 4'b0011;
														assign node51728 = (inp[3]) ? node51732 : node51729;
															assign node51729 = (inp[9]) ? 4'b0010 : 4'b0011;
															assign node51732 = (inp[9]) ? 4'b0011 : 4'b0010;
													assign node51735 = (inp[2]) ? node51751 : node51736;
														assign node51736 = (inp[3]) ? node51744 : node51737;
															assign node51737 = (inp[12]) ? node51741 : node51738;
																assign node51738 = (inp[9]) ? 4'b0010 : 4'b0011;
																assign node51741 = (inp[9]) ? 4'b0011 : 4'b0010;
															assign node51744 = (inp[9]) ? node51748 : node51745;
																assign node51745 = (inp[12]) ? 4'b0011 : 4'b0010;
																assign node51748 = (inp[12]) ? 4'b0010 : 4'b0011;
														assign node51751 = (inp[3]) ? node51759 : node51752;
															assign node51752 = (inp[9]) ? node51756 : node51753;
																assign node51753 = (inp[12]) ? 4'b0010 : 4'b0011;
																assign node51756 = (inp[12]) ? 4'b0011 : 4'b0010;
															assign node51759 = (inp[12]) ? node51763 : node51760;
																assign node51760 = (inp[9]) ? 4'b0011 : 4'b0010;
																assign node51763 = (inp[9]) ? 4'b0010 : 4'b0011;
												assign node51766 = (inp[3]) ? node51774 : node51767;
													assign node51767 = (inp[5]) ? node51771 : node51768;
														assign node51768 = (inp[9]) ? 4'b0011 : 4'b0010;
														assign node51771 = (inp[9]) ? 4'b0010 : 4'b0011;
													assign node51774 = (inp[5]) ? node51778 : node51775;
														assign node51775 = (inp[9]) ? 4'b0011 : 4'b0010;
														assign node51778 = (inp[9]) ? 4'b0010 : 4'b0011;
											assign node51781 = (inp[9]) ? node51801 : node51782;
												assign node51782 = (inp[5]) ? node51792 : node51783;
													assign node51783 = (inp[0]) ? 4'b0010 : node51784;
														assign node51784 = (inp[12]) ? node51788 : node51785;
															assign node51785 = (inp[3]) ? 4'b0011 : 4'b0010;
															assign node51788 = (inp[3]) ? 4'b0010 : 4'b0011;
													assign node51792 = (inp[0]) ? 4'b0011 : node51793;
														assign node51793 = (inp[12]) ? node51797 : node51794;
															assign node51794 = (inp[3]) ? 4'b0010 : 4'b0011;
															assign node51797 = (inp[3]) ? 4'b0011 : 4'b0010;
												assign node51801 = (inp[5]) ? node51817 : node51802;
													assign node51802 = (inp[0]) ? 4'b0011 : node51803;
														assign node51803 = (inp[2]) ? node51811 : node51804;
															assign node51804 = (inp[3]) ? node51808 : node51805;
																assign node51805 = (inp[12]) ? 4'b0010 : 4'b0011;
																assign node51808 = (inp[12]) ? 4'b0011 : 4'b0010;
															assign node51811 = (inp[12]) ? node51813 : 4'b0011;
																assign node51813 = (inp[3]) ? 4'b0011 : 4'b0010;
													assign node51817 = (inp[0]) ? 4'b0010 : node51818;
														assign node51818 = (inp[2]) ? node51824 : node51819;
															assign node51819 = (inp[3]) ? node51821 : 4'b0011;
																assign node51821 = (inp[12]) ? 4'b0010 : 4'b0011;
															assign node51824 = (inp[12]) ? node51828 : node51825;
																assign node51825 = (inp[3]) ? 4'b0011 : 4'b0010;
																assign node51828 = (inp[3]) ? 4'b0010 : 4'b0011;
							assign node51832 = (inp[15]) ? node52300 : node51833;
								assign node51833 = (inp[13]) ? node52117 : node51834;
									assign node51834 = (inp[10]) ? node52006 : node51835;
										assign node51835 = (inp[2]) ? node51909 : node51836;
											assign node51836 = (inp[12]) ? node51862 : node51837;
												assign node51837 = (inp[9]) ? node51847 : node51838;
													assign node51838 = (inp[5]) ? node51840 : 4'b0010;
														assign node51840 = (inp[3]) ? node51842 : 4'b0011;
															assign node51842 = (inp[0]) ? node51844 : 4'b0011;
																assign node51844 = (inp[1]) ? 4'b0011 : 4'b0010;
													assign node51847 = (inp[5]) ? node51855 : node51848;
														assign node51848 = (inp[1]) ? 4'b0011 : node51849;
															assign node51849 = (inp[0]) ? node51851 : 4'b0011;
																assign node51851 = (inp[3]) ? 4'b0010 : 4'b0011;
														assign node51855 = (inp[3]) ? node51857 : 4'b0010;
															assign node51857 = (inp[0]) ? node51859 : 4'b0010;
																assign node51859 = (inp[1]) ? 4'b0010 : 4'b0011;
												assign node51862 = (inp[3]) ? node51888 : node51863;
													assign node51863 = (inp[1]) ? node51879 : node51864;
														assign node51864 = (inp[9]) ? node51872 : node51865;
															assign node51865 = (inp[0]) ? node51869 : node51866;
																assign node51866 = (inp[5]) ? 4'b0011 : 4'b0010;
																assign node51869 = (inp[5]) ? 4'b0010 : 4'b0011;
															assign node51872 = (inp[5]) ? node51876 : node51873;
																assign node51873 = (inp[0]) ? 4'b0010 : 4'b0011;
																assign node51876 = (inp[0]) ? 4'b0011 : 4'b0010;
														assign node51879 = (inp[0]) ? 4'b0010 : node51880;
															assign node51880 = (inp[5]) ? node51884 : node51881;
																assign node51881 = (inp[9]) ? 4'b0010 : 4'b0011;
																assign node51884 = (inp[9]) ? 4'b0011 : 4'b0010;
													assign node51888 = (inp[1]) ? node51896 : node51889;
														assign node51889 = (inp[5]) ? node51893 : node51890;
															assign node51890 = (inp[9]) ? 4'b0011 : 4'b0010;
															assign node51893 = (inp[9]) ? 4'b0010 : 4'b0011;
														assign node51896 = (inp[9]) ? node51904 : node51897;
															assign node51897 = (inp[5]) ? node51901 : node51898;
																assign node51898 = (inp[0]) ? 4'b0011 : 4'b0010;
																assign node51901 = (inp[0]) ? 4'b0010 : 4'b0011;
															assign node51904 = (inp[0]) ? 4'b0011 : node51905;
																assign node51905 = (inp[5]) ? 4'b0010 : 4'b0011;
											assign node51909 = (inp[12]) ? node51951 : node51910;
												assign node51910 = (inp[0]) ? node51928 : node51911;
													assign node51911 = (inp[1]) ? node51919 : node51912;
														assign node51912 = (inp[9]) ? node51916 : node51913;
															assign node51913 = (inp[5]) ? 4'b0011 : 4'b0010;
															assign node51916 = (inp[5]) ? 4'b0010 : 4'b0011;
														assign node51919 = (inp[3]) ? 4'b0010 : node51920;
															assign node51920 = (inp[9]) ? node51924 : node51921;
																assign node51921 = (inp[5]) ? 4'b0011 : 4'b0010;
																assign node51924 = (inp[5]) ? 4'b0010 : 4'b0011;
													assign node51928 = (inp[3]) ? node51936 : node51929;
														assign node51929 = (inp[9]) ? node51933 : node51930;
															assign node51930 = (inp[5]) ? 4'b0011 : 4'b0010;
															assign node51933 = (inp[5]) ? 4'b0010 : 4'b0011;
														assign node51936 = (inp[9]) ? node51944 : node51937;
															assign node51937 = (inp[5]) ? node51941 : node51938;
																assign node51938 = (inp[1]) ? 4'b0010 : 4'b0011;
																assign node51941 = (inp[1]) ? 4'b0011 : 4'b0010;
															assign node51944 = (inp[5]) ? node51948 : node51945;
																assign node51945 = (inp[1]) ? 4'b0011 : 4'b0010;
																assign node51948 = (inp[1]) ? 4'b0010 : 4'b0011;
												assign node51951 = (inp[1]) ? node51975 : node51952;
													assign node51952 = (inp[5]) ? node51964 : node51953;
														assign node51953 = (inp[9]) ? node51959 : node51954;
															assign node51954 = (inp[0]) ? node51956 : 4'b0010;
																assign node51956 = (inp[3]) ? 4'b0010 : 4'b0011;
															assign node51959 = (inp[0]) ? node51961 : 4'b0011;
																assign node51961 = (inp[3]) ? 4'b0011 : 4'b0010;
														assign node51964 = (inp[9]) ? node51970 : node51965;
															assign node51965 = (inp[0]) ? node51967 : 4'b0011;
																assign node51967 = (inp[3]) ? 4'b0011 : 4'b0010;
															assign node51970 = (inp[3]) ? 4'b0010 : node51971;
																assign node51971 = (inp[0]) ? 4'b0011 : 4'b0010;
													assign node51975 = (inp[3]) ? node51991 : node51976;
														assign node51976 = (inp[0]) ? node51984 : node51977;
															assign node51977 = (inp[9]) ? node51981 : node51978;
																assign node51978 = (inp[5]) ? 4'b0010 : 4'b0011;
																assign node51981 = (inp[5]) ? 4'b0011 : 4'b0010;
															assign node51984 = (inp[9]) ? node51988 : node51985;
																assign node51985 = (inp[5]) ? 4'b0011 : 4'b0010;
																assign node51988 = (inp[5]) ? 4'b0010 : 4'b0011;
														assign node51991 = (inp[0]) ? node51999 : node51992;
															assign node51992 = (inp[9]) ? node51996 : node51993;
																assign node51993 = (inp[5]) ? 4'b0011 : 4'b0010;
																assign node51996 = (inp[5]) ? 4'b0010 : 4'b0011;
															assign node51999 = (inp[5]) ? node52003 : node52000;
																assign node52000 = (inp[9]) ? 4'b0010 : 4'b0011;
																assign node52003 = (inp[9]) ? 4'b0011 : 4'b0010;
										assign node52006 = (inp[3]) ? node52066 : node52007;
											assign node52007 = (inp[5]) ? node52041 : node52008;
												assign node52008 = (inp[9]) ? node52026 : node52009;
													assign node52009 = (inp[12]) ? node52011 : 4'b0010;
														assign node52011 = (inp[2]) ? node52019 : node52012;
															assign node52012 = (inp[0]) ? node52016 : node52013;
																assign node52013 = (inp[1]) ? 4'b0011 : 4'b0010;
																assign node52016 = (inp[1]) ? 4'b0010 : 4'b0011;
															assign node52019 = (inp[0]) ? node52023 : node52020;
																assign node52020 = (inp[1]) ? 4'b0011 : 4'b0010;
																assign node52023 = (inp[1]) ? 4'b0010 : 4'b0011;
													assign node52026 = (inp[12]) ? node52028 : 4'b0011;
														assign node52028 = (inp[2]) ? node52036 : node52029;
															assign node52029 = (inp[0]) ? node52033 : node52030;
																assign node52030 = (inp[1]) ? 4'b0010 : 4'b0011;
																assign node52033 = (inp[1]) ? 4'b0011 : 4'b0010;
															assign node52036 = (inp[0]) ? node52038 : 4'b0011;
																assign node52038 = (inp[1]) ? 4'b0011 : 4'b0010;
												assign node52041 = (inp[9]) ? node52057 : node52042;
													assign node52042 = (inp[12]) ? node52044 : 4'b0011;
														assign node52044 = (inp[2]) ? node52052 : node52045;
															assign node52045 = (inp[1]) ? node52049 : node52046;
																assign node52046 = (inp[0]) ? 4'b0010 : 4'b0011;
																assign node52049 = (inp[0]) ? 4'b0011 : 4'b0010;
															assign node52052 = (inp[1]) ? node52054 : 4'b0010;
																assign node52054 = (inp[0]) ? 4'b0011 : 4'b0010;
													assign node52057 = (inp[12]) ? node52059 : 4'b0010;
														assign node52059 = (inp[0]) ? node52063 : node52060;
															assign node52060 = (inp[1]) ? 4'b0011 : 4'b0010;
															assign node52063 = (inp[1]) ? 4'b0010 : 4'b0011;
											assign node52066 = (inp[0]) ? node52082 : node52067;
												assign node52067 = (inp[1]) ? node52075 : node52068;
													assign node52068 = (inp[9]) ? node52072 : node52069;
														assign node52069 = (inp[5]) ? 4'b0011 : 4'b0010;
														assign node52072 = (inp[5]) ? 4'b0010 : 4'b0011;
													assign node52075 = (inp[9]) ? node52079 : node52076;
														assign node52076 = (inp[5]) ? 4'b0011 : 4'b0010;
														assign node52079 = (inp[5]) ? 4'b0010 : 4'b0011;
												assign node52082 = (inp[12]) ? node52098 : node52083;
													assign node52083 = (inp[1]) ? node52091 : node52084;
														assign node52084 = (inp[9]) ? node52088 : node52085;
															assign node52085 = (inp[5]) ? 4'b0010 : 4'b0011;
															assign node52088 = (inp[5]) ? 4'b0011 : 4'b0010;
														assign node52091 = (inp[5]) ? node52095 : node52092;
															assign node52092 = (inp[9]) ? 4'b0011 : 4'b0010;
															assign node52095 = (inp[9]) ? 4'b0010 : 4'b0011;
													assign node52098 = (inp[2]) ? node52112 : node52099;
														assign node52099 = (inp[1]) ? node52105 : node52100;
															assign node52100 = (inp[5]) ? node52102 : 4'b0010;
																assign node52102 = (inp[9]) ? 4'b0010 : 4'b0011;
															assign node52105 = (inp[5]) ? node52109 : node52106;
																assign node52106 = (inp[9]) ? 4'b0010 : 4'b0011;
																assign node52109 = (inp[9]) ? 4'b0011 : 4'b0010;
														assign node52112 = (inp[5]) ? 4'b0010 : node52113;
															assign node52113 = (inp[1]) ? 4'b0010 : 4'b0011;
									assign node52117 = (inp[2]) ? node52211 : node52118;
										assign node52118 = (inp[9]) ? node52164 : node52119;
											assign node52119 = (inp[5]) ? node52141 : node52120;
												assign node52120 = (inp[12]) ? node52128 : node52121;
													assign node52121 = (inp[3]) ? node52123 : 4'b0110;
														assign node52123 = (inp[1]) ? node52125 : 4'b0110;
															assign node52125 = (inp[0]) ? 4'b0110 : 4'b0111;
													assign node52128 = (inp[3]) ? node52136 : node52129;
														assign node52129 = (inp[0]) ? node52133 : node52130;
															assign node52130 = (inp[1]) ? 4'b0111 : 4'b0110;
															assign node52133 = (inp[1]) ? 4'b0110 : 4'b0111;
														assign node52136 = (inp[0]) ? 4'b0110 : node52137;
															assign node52137 = (inp[1]) ? 4'b0110 : 4'b0111;
												assign node52141 = (inp[0]) ? node52155 : node52142;
													assign node52142 = (inp[12]) ? node52148 : node52143;
														assign node52143 = (inp[3]) ? node52145 : 4'b0111;
															assign node52145 = (inp[1]) ? 4'b0110 : 4'b0111;
														assign node52148 = (inp[1]) ? node52152 : node52149;
															assign node52149 = (inp[3]) ? 4'b0110 : 4'b0111;
															assign node52152 = (inp[3]) ? 4'b0111 : 4'b0110;
													assign node52155 = (inp[10]) ? 4'b0111 : node52156;
														assign node52156 = (inp[3]) ? 4'b0111 : node52157;
															assign node52157 = (inp[1]) ? 4'b0111 : node52158;
																assign node52158 = (inp[12]) ? 4'b0110 : 4'b0111;
											assign node52164 = (inp[5]) ? node52190 : node52165;
												assign node52165 = (inp[12]) ? node52173 : node52166;
													assign node52166 = (inp[1]) ? node52168 : 4'b0111;
														assign node52168 = (inp[3]) ? node52170 : 4'b0111;
															assign node52170 = (inp[0]) ? 4'b0111 : 4'b0110;
													assign node52173 = (inp[3]) ? node52185 : node52174;
														assign node52174 = (inp[10]) ? node52180 : node52175;
															assign node52175 = (inp[0]) ? node52177 : 4'b0110;
																assign node52177 = (inp[1]) ? 4'b0111 : 4'b0110;
															assign node52180 = (inp[1]) ? 4'b0110 : node52181;
																assign node52181 = (inp[0]) ? 4'b0110 : 4'b0111;
														assign node52185 = (inp[1]) ? 4'b0111 : node52186;
															assign node52186 = (inp[10]) ? 4'b0110 : 4'b0111;
												assign node52190 = (inp[0]) ? node52204 : node52191;
													assign node52191 = (inp[1]) ? node52197 : node52192;
														assign node52192 = (inp[12]) ? node52194 : 4'b0110;
															assign node52194 = (inp[3]) ? 4'b0111 : 4'b0110;
														assign node52197 = (inp[12]) ? node52201 : node52198;
															assign node52198 = (inp[3]) ? 4'b0111 : 4'b0110;
															assign node52201 = (inp[3]) ? 4'b0110 : 4'b0111;
													assign node52204 = (inp[12]) ? node52206 : 4'b0110;
														assign node52206 = (inp[1]) ? 4'b0110 : node52207;
															assign node52207 = (inp[3]) ? 4'b0110 : 4'b0111;
										assign node52211 = (inp[0]) ? node52269 : node52212;
											assign node52212 = (inp[12]) ? node52236 : node52213;
												assign node52213 = (inp[9]) ? node52225 : node52214;
													assign node52214 = (inp[5]) ? node52220 : node52215;
														assign node52215 = (inp[3]) ? node52217 : 4'b0110;
															assign node52217 = (inp[1]) ? 4'b0111 : 4'b0110;
														assign node52220 = (inp[3]) ? node52222 : 4'b0111;
															assign node52222 = (inp[1]) ? 4'b0110 : 4'b0111;
													assign node52225 = (inp[5]) ? node52231 : node52226;
														assign node52226 = (inp[1]) ? node52228 : 4'b0111;
															assign node52228 = (inp[3]) ? 4'b0110 : 4'b0111;
														assign node52231 = (inp[1]) ? node52233 : 4'b0110;
															assign node52233 = (inp[3]) ? 4'b0111 : 4'b0110;
												assign node52236 = (inp[9]) ? node52256 : node52237;
													assign node52237 = (inp[5]) ? node52249 : node52238;
														assign node52238 = (inp[10]) ? node52244 : node52239;
															assign node52239 = (inp[1]) ? 4'b0111 : node52240;
																assign node52240 = (inp[3]) ? 4'b0111 : 4'b0110;
															assign node52244 = (inp[1]) ? node52246 : 4'b0111;
																assign node52246 = (inp[3]) ? 4'b0110 : 4'b0111;
														assign node52249 = (inp[3]) ? node52253 : node52250;
															assign node52250 = (inp[1]) ? 4'b0110 : 4'b0111;
															assign node52253 = (inp[1]) ? 4'b0111 : 4'b0110;
													assign node52256 = (inp[5]) ? node52264 : node52257;
														assign node52257 = (inp[3]) ? node52261 : node52258;
															assign node52258 = (inp[1]) ? 4'b0110 : 4'b0111;
															assign node52261 = (inp[1]) ? 4'b0111 : 4'b0110;
														assign node52264 = (inp[1]) ? 4'b0111 : node52265;
															assign node52265 = (inp[3]) ? 4'b0111 : 4'b0110;
											assign node52269 = (inp[5]) ? node52285 : node52270;
												assign node52270 = (inp[9]) ? node52278 : node52271;
													assign node52271 = (inp[3]) ? 4'b0110 : node52272;
														assign node52272 = (inp[1]) ? 4'b0110 : node52273;
															assign node52273 = (inp[12]) ? 4'b0111 : 4'b0110;
													assign node52278 = (inp[1]) ? 4'b0111 : node52279;
														assign node52279 = (inp[10]) ? node52281 : 4'b0111;
															assign node52281 = (inp[3]) ? 4'b0111 : 4'b0110;
												assign node52285 = (inp[9]) ? node52293 : node52286;
													assign node52286 = (inp[1]) ? 4'b0111 : node52287;
														assign node52287 = (inp[12]) ? node52289 : 4'b0111;
															assign node52289 = (inp[3]) ? 4'b0111 : 4'b0110;
													assign node52293 = (inp[3]) ? 4'b0110 : node52294;
														assign node52294 = (inp[1]) ? 4'b0110 : node52295;
															assign node52295 = (inp[12]) ? 4'b0111 : 4'b0110;
								assign node52300 = (inp[13]) ? node52530 : node52301;
									assign node52301 = (inp[0]) ? node52399 : node52302;
										assign node52302 = (inp[3]) ? node52350 : node52303;
											assign node52303 = (inp[12]) ? node52311 : node52304;
												assign node52304 = (inp[9]) ? node52308 : node52305;
													assign node52305 = (inp[5]) ? 4'b0111 : 4'b0110;
													assign node52308 = (inp[5]) ? 4'b0110 : 4'b0111;
												assign node52311 = (inp[10]) ? node52343 : node52312;
													assign node52312 = (inp[1]) ? node52328 : node52313;
														assign node52313 = (inp[2]) ? node52321 : node52314;
															assign node52314 = (inp[9]) ? node52318 : node52315;
																assign node52315 = (inp[5]) ? 4'b0111 : 4'b0110;
																assign node52318 = (inp[5]) ? 4'b0110 : 4'b0111;
															assign node52321 = (inp[5]) ? node52325 : node52322;
																assign node52322 = (inp[9]) ? 4'b0111 : 4'b0110;
																assign node52325 = (inp[9]) ? 4'b0110 : 4'b0111;
														assign node52328 = (inp[2]) ? node52336 : node52329;
															assign node52329 = (inp[9]) ? node52333 : node52330;
																assign node52330 = (inp[5]) ? 4'b0111 : 4'b0110;
																assign node52333 = (inp[5]) ? 4'b0110 : 4'b0111;
															assign node52336 = (inp[5]) ? node52340 : node52337;
																assign node52337 = (inp[9]) ? 4'b0111 : 4'b0110;
																assign node52340 = (inp[9]) ? 4'b0110 : 4'b0111;
													assign node52343 = (inp[5]) ? node52347 : node52344;
														assign node52344 = (inp[9]) ? 4'b0111 : 4'b0110;
														assign node52347 = (inp[9]) ? 4'b0110 : 4'b0111;
											assign node52350 = (inp[2]) ? node52376 : node52351;
												assign node52351 = (inp[1]) ? node52361 : node52352;
													assign node52352 = (inp[10]) ? 4'b0110 : node52353;
														assign node52353 = (inp[9]) ? node52357 : node52354;
															assign node52354 = (inp[5]) ? 4'b0111 : 4'b0110;
															assign node52357 = (inp[5]) ? 4'b0110 : 4'b0111;
													assign node52361 = (inp[9]) ? node52369 : node52362;
														assign node52362 = (inp[12]) ? node52366 : node52363;
															assign node52363 = (inp[5]) ? 4'b0110 : 4'b0111;
															assign node52366 = (inp[5]) ? 4'b0111 : 4'b0110;
														assign node52369 = (inp[5]) ? node52373 : node52370;
															assign node52370 = (inp[12]) ? 4'b0111 : 4'b0110;
															assign node52373 = (inp[12]) ? 4'b0110 : 4'b0111;
												assign node52376 = (inp[9]) ? node52388 : node52377;
													assign node52377 = (inp[5]) ? node52383 : node52378;
														assign node52378 = (inp[12]) ? 4'b0110 : node52379;
															assign node52379 = (inp[1]) ? 4'b0111 : 4'b0110;
														assign node52383 = (inp[12]) ? 4'b0111 : node52384;
															assign node52384 = (inp[1]) ? 4'b0110 : 4'b0111;
													assign node52388 = (inp[5]) ? node52394 : node52389;
														assign node52389 = (inp[1]) ? node52391 : 4'b0111;
															assign node52391 = (inp[12]) ? 4'b0111 : 4'b0110;
														assign node52394 = (inp[1]) ? node52396 : 4'b0110;
															assign node52396 = (inp[12]) ? 4'b0110 : 4'b0111;
										assign node52399 = (inp[1]) ? node52473 : node52400;
											assign node52400 = (inp[9]) ? node52430 : node52401;
												assign node52401 = (inp[12]) ? node52423 : node52402;
													assign node52402 = (inp[2]) ? node52410 : node52403;
														assign node52403 = (inp[5]) ? node52407 : node52404;
															assign node52404 = (inp[3]) ? 4'b0111 : 4'b0110;
															assign node52407 = (inp[3]) ? 4'b0110 : 4'b0111;
														assign node52410 = (inp[10]) ? node52418 : node52411;
															assign node52411 = (inp[3]) ? node52415 : node52412;
																assign node52412 = (inp[5]) ? 4'b0111 : 4'b0110;
																assign node52415 = (inp[5]) ? 4'b0110 : 4'b0111;
															assign node52418 = (inp[5]) ? node52420 : 4'b0111;
																assign node52420 = (inp[3]) ? 4'b0110 : 4'b0111;
													assign node52423 = (inp[5]) ? node52427 : node52424;
														assign node52424 = (inp[3]) ? 4'b0110 : 4'b0111;
														assign node52427 = (inp[3]) ? 4'b0111 : 4'b0110;
												assign node52430 = (inp[2]) ? node52458 : node52431;
													assign node52431 = (inp[5]) ? node52447 : node52432;
														assign node52432 = (inp[10]) ? node52440 : node52433;
															assign node52433 = (inp[12]) ? node52437 : node52434;
																assign node52434 = (inp[3]) ? 4'b0110 : 4'b0111;
																assign node52437 = (inp[3]) ? 4'b0111 : 4'b0110;
															assign node52440 = (inp[12]) ? node52444 : node52441;
																assign node52441 = (inp[3]) ? 4'b0110 : 4'b0111;
																assign node52444 = (inp[3]) ? 4'b0111 : 4'b0110;
														assign node52447 = (inp[10]) ? node52453 : node52448;
															assign node52448 = (inp[12]) ? 4'b0111 : node52449;
																assign node52449 = (inp[3]) ? 4'b0111 : 4'b0110;
															assign node52453 = (inp[3]) ? node52455 : 4'b0111;
																assign node52455 = (inp[12]) ? 4'b0110 : 4'b0111;
													assign node52458 = (inp[5]) ? node52466 : node52459;
														assign node52459 = (inp[12]) ? node52463 : node52460;
															assign node52460 = (inp[3]) ? 4'b0110 : 4'b0111;
															assign node52463 = (inp[3]) ? 4'b0111 : 4'b0110;
														assign node52466 = (inp[3]) ? node52470 : node52467;
															assign node52467 = (inp[12]) ? 4'b0111 : 4'b0110;
															assign node52470 = (inp[12]) ? 4'b0110 : 4'b0111;
											assign node52473 = (inp[2]) ? node52505 : node52474;
												assign node52474 = (inp[3]) ? node52490 : node52475;
													assign node52475 = (inp[12]) ? node52483 : node52476;
														assign node52476 = (inp[5]) ? node52480 : node52477;
															assign node52477 = (inp[9]) ? 4'b0110 : 4'b0111;
															assign node52480 = (inp[9]) ? 4'b0111 : 4'b0110;
														assign node52483 = (inp[5]) ? node52487 : node52484;
															assign node52484 = (inp[9]) ? 4'b0111 : 4'b0110;
															assign node52487 = (inp[9]) ? 4'b0110 : 4'b0111;
													assign node52490 = (inp[12]) ? node52498 : node52491;
														assign node52491 = (inp[9]) ? node52495 : node52492;
															assign node52492 = (inp[5]) ? 4'b0111 : 4'b0110;
															assign node52495 = (inp[5]) ? 4'b0110 : 4'b0111;
														assign node52498 = (inp[9]) ? node52502 : node52499;
															assign node52499 = (inp[5]) ? 4'b0111 : 4'b0110;
															assign node52502 = (inp[5]) ? 4'b0110 : 4'b0111;
												assign node52505 = (inp[9]) ? node52519 : node52506;
													assign node52506 = (inp[5]) ? node52514 : node52507;
														assign node52507 = (inp[10]) ? node52509 : 4'b0111;
															assign node52509 = (inp[3]) ? 4'b0110 : node52510;
																assign node52510 = (inp[12]) ? 4'b0110 : 4'b0111;
														assign node52514 = (inp[3]) ? 4'b0111 : node52515;
															assign node52515 = (inp[12]) ? 4'b0111 : 4'b0110;
													assign node52519 = (inp[5]) ? node52525 : node52520;
														assign node52520 = (inp[3]) ? 4'b0111 : node52521;
															assign node52521 = (inp[12]) ? 4'b0111 : 4'b0110;
														assign node52525 = (inp[3]) ? 4'b0110 : node52526;
															assign node52526 = (inp[12]) ? 4'b0110 : 4'b0111;
									assign node52530 = (inp[2]) ? node52626 : node52531;
										assign node52531 = (inp[5]) ? node52583 : node52532;
											assign node52532 = (inp[9]) ? node52560 : node52533;
												assign node52533 = (inp[12]) ? node52553 : node52534;
													assign node52534 = (inp[1]) ? node52548 : node52535;
														assign node52535 = (inp[10]) ? node52543 : node52536;
															assign node52536 = (inp[3]) ? node52540 : node52537;
																assign node52537 = (inp[0]) ? 4'b0010 : 4'b0011;
																assign node52540 = (inp[0]) ? 4'b0011 : 4'b0010;
															assign node52543 = (inp[0]) ? 4'b0011 : node52544;
																assign node52544 = (inp[3]) ? 4'b0010 : 4'b0011;
														assign node52548 = (inp[0]) ? 4'b0010 : node52549;
															assign node52549 = (inp[3]) ? 4'b0011 : 4'b0010;
													assign node52553 = (inp[0]) ? 4'b0010 : node52554;
														assign node52554 = (inp[1]) ? node52556 : 4'b0010;
															assign node52556 = (inp[3]) ? 4'b0010 : 4'b0011;
												assign node52560 = (inp[0]) ? 4'b0011 : node52561;
													assign node52561 = (inp[1]) ? node52567 : node52562;
														assign node52562 = (inp[3]) ? 4'b0011 : node52563;
															assign node52563 = (inp[12]) ? 4'b0011 : 4'b0010;
														assign node52567 = (inp[10]) ? node52575 : node52568;
															assign node52568 = (inp[12]) ? node52572 : node52569;
																assign node52569 = (inp[3]) ? 4'b0010 : 4'b0011;
																assign node52572 = (inp[3]) ? 4'b0011 : 4'b0010;
															assign node52575 = (inp[12]) ? node52579 : node52576;
																assign node52576 = (inp[3]) ? 4'b0010 : 4'b0011;
																assign node52579 = (inp[3]) ? 4'b0011 : 4'b0010;
											assign node52583 = (inp[9]) ? node52605 : node52584;
												assign node52584 = (inp[0]) ? node52598 : node52585;
													assign node52585 = (inp[3]) ? node52593 : node52586;
														assign node52586 = (inp[1]) ? node52590 : node52587;
															assign node52587 = (inp[12]) ? 4'b0011 : 4'b0010;
															assign node52590 = (inp[12]) ? 4'b0010 : 4'b0011;
														assign node52593 = (inp[1]) ? node52595 : 4'b0011;
															assign node52595 = (inp[12]) ? 4'b0011 : 4'b0010;
													assign node52598 = (inp[3]) ? node52600 : 4'b0011;
														assign node52600 = (inp[12]) ? 4'b0011 : node52601;
															assign node52601 = (inp[10]) ? 4'b0010 : 4'b0011;
												assign node52605 = (inp[0]) ? node52619 : node52606;
													assign node52606 = (inp[1]) ? node52612 : node52607;
														assign node52607 = (inp[12]) ? 4'b0010 : node52608;
															assign node52608 = (inp[3]) ? 4'b0010 : 4'b0011;
														assign node52612 = (inp[3]) ? node52616 : node52613;
															assign node52613 = (inp[12]) ? 4'b0011 : 4'b0010;
															assign node52616 = (inp[12]) ? 4'b0010 : 4'b0011;
													assign node52619 = (inp[12]) ? 4'b0010 : node52620;
														assign node52620 = (inp[3]) ? node52622 : 4'b0010;
															assign node52622 = (inp[1]) ? 4'b0010 : 4'b0011;
										assign node52626 = (inp[1]) ? node52716 : node52627;
											assign node52627 = (inp[10]) ? node52667 : node52628;
												assign node52628 = (inp[0]) ? node52644 : node52629;
													assign node52629 = (inp[9]) ? node52635 : node52630;
														assign node52630 = (inp[5]) ? node52632 : 4'b0010;
															assign node52632 = (inp[3]) ? 4'b0011 : 4'b0010;
														assign node52635 = (inp[5]) ? node52639 : node52636;
															assign node52636 = (inp[12]) ? 4'b0011 : 4'b0010;
															assign node52639 = (inp[3]) ? 4'b0010 : node52640;
																assign node52640 = (inp[12]) ? 4'b0010 : 4'b0011;
													assign node52644 = (inp[5]) ? node52656 : node52645;
														assign node52645 = (inp[9]) ? node52651 : node52646;
															assign node52646 = (inp[3]) ? node52648 : 4'b0010;
																assign node52648 = (inp[12]) ? 4'b0010 : 4'b0011;
															assign node52651 = (inp[3]) ? node52653 : 4'b0011;
																assign node52653 = (inp[12]) ? 4'b0011 : 4'b0010;
														assign node52656 = (inp[9]) ? node52662 : node52657;
															assign node52657 = (inp[3]) ? node52659 : 4'b0011;
																assign node52659 = (inp[12]) ? 4'b0011 : 4'b0010;
															assign node52662 = (inp[12]) ? 4'b0010 : node52663;
																assign node52663 = (inp[3]) ? 4'b0011 : 4'b0010;
												assign node52667 = (inp[3]) ? node52687 : node52668;
													assign node52668 = (inp[9]) ? node52680 : node52669;
														assign node52669 = (inp[5]) ? node52675 : node52670;
															assign node52670 = (inp[0]) ? 4'b0010 : node52671;
																assign node52671 = (inp[12]) ? 4'b0010 : 4'b0011;
															assign node52675 = (inp[12]) ? 4'b0011 : node52676;
																assign node52676 = (inp[0]) ? 4'b0011 : 4'b0010;
														assign node52680 = (inp[5]) ? 4'b0010 : node52681;
															assign node52681 = (inp[12]) ? 4'b0011 : node52682;
																assign node52682 = (inp[0]) ? 4'b0011 : 4'b0010;
													assign node52687 = (inp[0]) ? node52701 : node52688;
														assign node52688 = (inp[12]) ? node52694 : node52689;
															assign node52689 = (inp[5]) ? 4'b0011 : node52690;
																assign node52690 = (inp[9]) ? 4'b0011 : 4'b0010;
															assign node52694 = (inp[9]) ? node52698 : node52695;
																assign node52695 = (inp[5]) ? 4'b0011 : 4'b0010;
																assign node52698 = (inp[5]) ? 4'b0010 : 4'b0011;
														assign node52701 = (inp[12]) ? node52709 : node52702;
															assign node52702 = (inp[5]) ? node52706 : node52703;
																assign node52703 = (inp[9]) ? 4'b0010 : 4'b0011;
																assign node52706 = (inp[9]) ? 4'b0011 : 4'b0010;
															assign node52709 = (inp[9]) ? node52713 : node52710;
																assign node52710 = (inp[5]) ? 4'b0011 : 4'b0010;
																assign node52713 = (inp[5]) ? 4'b0010 : 4'b0011;
											assign node52716 = (inp[12]) ? node52756 : node52717;
												assign node52717 = (inp[3]) ? node52733 : node52718;
													assign node52718 = (inp[10]) ? node52726 : node52719;
														assign node52719 = (inp[5]) ? node52723 : node52720;
															assign node52720 = (inp[9]) ? 4'b0011 : 4'b0010;
															assign node52723 = (inp[9]) ? 4'b0010 : 4'b0011;
														assign node52726 = (inp[9]) ? node52730 : node52727;
															assign node52727 = (inp[5]) ? 4'b0011 : 4'b0010;
															assign node52730 = (inp[5]) ? 4'b0010 : 4'b0011;
													assign node52733 = (inp[10]) ? node52749 : node52734;
														assign node52734 = (inp[0]) ? node52742 : node52735;
															assign node52735 = (inp[5]) ? node52739 : node52736;
																assign node52736 = (inp[9]) ? 4'b0010 : 4'b0011;
																assign node52739 = (inp[9]) ? 4'b0011 : 4'b0010;
															assign node52742 = (inp[5]) ? node52746 : node52743;
																assign node52743 = (inp[9]) ? 4'b0011 : 4'b0010;
																assign node52746 = (inp[9]) ? 4'b0010 : 4'b0011;
														assign node52749 = (inp[9]) ? node52751 : 4'b0010;
															assign node52751 = (inp[0]) ? 4'b0010 : node52752;
																assign node52752 = (inp[5]) ? 4'b0011 : 4'b0010;
												assign node52756 = (inp[5]) ? node52768 : node52757;
													assign node52757 = (inp[9]) ? node52763 : node52758;
														assign node52758 = (inp[0]) ? 4'b0010 : node52759;
															assign node52759 = (inp[3]) ? 4'b0010 : 4'b0011;
														assign node52763 = (inp[3]) ? 4'b0011 : node52764;
															assign node52764 = (inp[0]) ? 4'b0011 : 4'b0010;
													assign node52768 = (inp[9]) ? node52776 : node52769;
														assign node52769 = (inp[10]) ? 4'b0011 : node52770;
															assign node52770 = (inp[0]) ? 4'b0011 : node52771;
																assign node52771 = (inp[3]) ? 4'b0011 : 4'b0010;
														assign node52776 = (inp[3]) ? 4'b0010 : node52777;
															assign node52777 = (inp[0]) ? 4'b0010 : 4'b0011;
						assign node52781 = (inp[15]) ? node52979 : node52782;
							assign node52782 = (inp[1]) ? node52900 : node52783;
								assign node52783 = (inp[3]) ? node52893 : node52784;
									assign node52784 = (inp[12]) ? node52800 : node52785;
										assign node52785 = (inp[13]) ? node52793 : node52786;
											assign node52786 = (inp[5]) ? node52790 : node52787;
												assign node52787 = (inp[0]) ? 4'b0001 : 4'b0000;
												assign node52790 = (inp[0]) ? 4'b0000 : 4'b0001;
											assign node52793 = (inp[5]) ? node52797 : node52794;
												assign node52794 = (inp[0]) ? 4'b0001 : 4'b0000;
												assign node52797 = (inp[0]) ? 4'b0000 : 4'b0001;
										assign node52800 = (inp[11]) ? node52846 : node52801;
											assign node52801 = (inp[13]) ? node52809 : node52802;
												assign node52802 = (inp[5]) ? node52806 : node52803;
													assign node52803 = (inp[0]) ? 4'b0001 : 4'b0000;
													assign node52806 = (inp[0]) ? 4'b0000 : 4'b0001;
												assign node52809 = (inp[10]) ? node52823 : node52810;
													assign node52810 = (inp[9]) ? node52818 : node52811;
														assign node52811 = (inp[5]) ? node52815 : node52812;
															assign node52812 = (inp[0]) ? 4'b0000 : 4'b0001;
															assign node52815 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node52818 = (inp[5]) ? 4'b0001 : node52819;
															assign node52819 = (inp[0]) ? 4'b0000 : 4'b0001;
													assign node52823 = (inp[2]) ? node52831 : node52824;
														assign node52824 = (inp[5]) ? node52828 : node52825;
															assign node52825 = (inp[0]) ? 4'b0000 : 4'b0001;
															assign node52828 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node52831 = (inp[9]) ? node52839 : node52832;
															assign node52832 = (inp[0]) ? node52836 : node52833;
																assign node52833 = (inp[5]) ? 4'b0000 : 4'b0001;
																assign node52836 = (inp[5]) ? 4'b0001 : 4'b0000;
															assign node52839 = (inp[0]) ? node52843 : node52840;
																assign node52840 = (inp[5]) ? 4'b0000 : 4'b0001;
																assign node52843 = (inp[5]) ? 4'b0001 : 4'b0000;
											assign node52846 = (inp[5]) ? node52878 : node52847;
												assign node52847 = (inp[10]) ? node52871 : node52848;
													assign node52848 = (inp[2]) ? node52864 : node52849;
														assign node52849 = (inp[9]) ? node52857 : node52850;
															assign node52850 = (inp[0]) ? node52854 : node52851;
																assign node52851 = (inp[13]) ? 4'b0001 : 4'b0000;
																assign node52854 = (inp[13]) ? 4'b0000 : 4'b0001;
															assign node52857 = (inp[0]) ? node52861 : node52858;
																assign node52858 = (inp[13]) ? 4'b0001 : 4'b0000;
																assign node52861 = (inp[13]) ? 4'b0000 : 4'b0001;
														assign node52864 = (inp[0]) ? node52868 : node52865;
															assign node52865 = (inp[13]) ? 4'b0001 : 4'b0000;
															assign node52868 = (inp[13]) ? 4'b0000 : 4'b0001;
													assign node52871 = (inp[13]) ? node52875 : node52872;
														assign node52872 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node52875 = (inp[0]) ? 4'b0000 : 4'b0001;
												assign node52878 = (inp[9]) ? node52886 : node52879;
													assign node52879 = (inp[13]) ? node52883 : node52880;
														assign node52880 = (inp[0]) ? 4'b0000 : 4'b0001;
														assign node52883 = (inp[0]) ? 4'b0001 : 4'b0000;
													assign node52886 = (inp[13]) ? node52890 : node52887;
														assign node52887 = (inp[0]) ? 4'b0000 : 4'b0001;
														assign node52890 = (inp[0]) ? 4'b0001 : 4'b0000;
									assign node52893 = (inp[13]) ? node52897 : node52894;
										assign node52894 = (inp[5]) ? 4'b0101 : 4'b0100;
										assign node52897 = (inp[5]) ? 4'b0100 : 4'b0101;
								assign node52900 = (inp[13]) ? node52968 : node52901;
									assign node52901 = (inp[5]) ? node52943 : node52902;
										assign node52902 = (inp[3]) ? 4'b0100 : node52903;
											assign node52903 = (inp[2]) ? node52919 : node52904;
												assign node52904 = (inp[9]) ? node52912 : node52905;
													assign node52905 = (inp[12]) ? node52909 : node52906;
														assign node52906 = (inp[0]) ? 4'b0101 : 4'b0100;
														assign node52909 = (inp[0]) ? 4'b0100 : 4'b0101;
													assign node52912 = (inp[0]) ? node52916 : node52913;
														assign node52913 = (inp[12]) ? 4'b0101 : 4'b0100;
														assign node52916 = (inp[12]) ? 4'b0100 : 4'b0101;
												assign node52919 = (inp[10]) ? node52927 : node52920;
													assign node52920 = (inp[12]) ? node52924 : node52921;
														assign node52921 = (inp[0]) ? 4'b0101 : 4'b0100;
														assign node52924 = (inp[0]) ? 4'b0100 : 4'b0101;
													assign node52927 = (inp[11]) ? node52935 : node52928;
														assign node52928 = (inp[12]) ? node52932 : node52929;
															assign node52929 = (inp[9]) ? 4'b0101 : 4'b0100;
															assign node52932 = (inp[0]) ? 4'b0100 : 4'b0101;
														assign node52935 = (inp[0]) ? node52939 : node52936;
															assign node52936 = (inp[12]) ? 4'b0101 : 4'b0100;
															assign node52939 = (inp[12]) ? 4'b0100 : 4'b0101;
										assign node52943 = (inp[3]) ? 4'b0101 : node52944;
											assign node52944 = (inp[9]) ? node52952 : node52945;
												assign node52945 = (inp[12]) ? node52949 : node52946;
													assign node52946 = (inp[0]) ? 4'b0100 : 4'b0101;
													assign node52949 = (inp[0]) ? 4'b0101 : 4'b0100;
												assign node52952 = (inp[10]) ? node52960 : node52953;
													assign node52953 = (inp[12]) ? node52957 : node52954;
														assign node52954 = (inp[0]) ? 4'b0100 : 4'b0101;
														assign node52957 = (inp[0]) ? 4'b0101 : 4'b0100;
													assign node52960 = (inp[12]) ? node52964 : node52961;
														assign node52961 = (inp[0]) ? 4'b0100 : 4'b0101;
														assign node52964 = (inp[0]) ? 4'b0101 : 4'b0100;
									assign node52968 = (inp[5]) ? node52974 : node52969;
										assign node52969 = (inp[0]) ? 4'b0101 : node52970;
											assign node52970 = (inp[3]) ? 4'b0101 : 4'b0100;
										assign node52974 = (inp[0]) ? 4'b0100 : node52975;
											assign node52975 = (inp[3]) ? 4'b0100 : 4'b0101;
							assign node52979 = (inp[3]) ? node53133 : node52980;
								assign node52980 = (inp[1]) ? node53004 : node52981;
									assign node52981 = (inp[5]) ? node52993 : node52982;
										assign node52982 = (inp[0]) ? node52988 : node52983;
											assign node52983 = (inp[12]) ? 4'b0100 : node52984;
												assign node52984 = (inp[13]) ? 4'b0101 : 4'b0100;
											assign node52988 = (inp[13]) ? node52990 : 4'b0101;
												assign node52990 = (inp[12]) ? 4'b0101 : 4'b0100;
										assign node52993 = (inp[0]) ? node52999 : node52994;
											assign node52994 = (inp[13]) ? node52996 : 4'b0101;
												assign node52996 = (inp[12]) ? 4'b0101 : 4'b0100;
											assign node52999 = (inp[13]) ? node53001 : 4'b0100;
												assign node53001 = (inp[12]) ? 4'b0100 : 4'b0101;
									assign node53004 = (inp[13]) ? node53118 : node53005;
										assign node53005 = (inp[11]) ? node53059 : node53006;
											assign node53006 = (inp[2]) ? node53022 : node53007;
												assign node53007 = (inp[12]) ? node53015 : node53008;
													assign node53008 = (inp[0]) ? node53012 : node53009;
														assign node53009 = (inp[5]) ? 4'b0000 : 4'b0001;
														assign node53012 = (inp[5]) ? 4'b0001 : 4'b0000;
													assign node53015 = (inp[5]) ? node53019 : node53016;
														assign node53016 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node53019 = (inp[0]) ? 4'b0000 : 4'b0001;
												assign node53022 = (inp[10]) ? node53046 : node53023;
													assign node53023 = (inp[9]) ? node53033 : node53024;
														assign node53024 = (inp[0]) ? 4'b0000 : node53025;
															assign node53025 = (inp[12]) ? node53029 : node53026;
																assign node53026 = (inp[5]) ? 4'b0000 : 4'b0001;
																assign node53029 = (inp[5]) ? 4'b0001 : 4'b0000;
														assign node53033 = (inp[0]) ? node53041 : node53034;
															assign node53034 = (inp[5]) ? node53038 : node53035;
																assign node53035 = (inp[12]) ? 4'b0000 : 4'b0001;
																assign node53038 = (inp[12]) ? 4'b0001 : 4'b0000;
															assign node53041 = (inp[5]) ? node53043 : 4'b0001;
																assign node53043 = (inp[12]) ? 4'b0000 : 4'b0001;
													assign node53046 = (inp[0]) ? node53052 : node53047;
														assign node53047 = (inp[9]) ? 4'b0000 : node53048;
															assign node53048 = (inp[12]) ? 4'b0001 : 4'b0000;
														assign node53052 = (inp[5]) ? node53056 : node53053;
															assign node53053 = (inp[12]) ? 4'b0001 : 4'b0000;
															assign node53056 = (inp[12]) ? 4'b0000 : 4'b0001;
											assign node53059 = (inp[2]) ? node53103 : node53060;
												assign node53060 = (inp[10]) ? node53084 : node53061;
													assign node53061 = (inp[12]) ? node53069 : node53062;
														assign node53062 = (inp[0]) ? node53066 : node53063;
															assign node53063 = (inp[5]) ? 4'b0000 : 4'b0001;
															assign node53066 = (inp[5]) ? 4'b0001 : 4'b0000;
														assign node53069 = (inp[9]) ? node53077 : node53070;
															assign node53070 = (inp[5]) ? node53074 : node53071;
																assign node53071 = (inp[0]) ? 4'b0001 : 4'b0000;
																assign node53074 = (inp[0]) ? 4'b0000 : 4'b0001;
															assign node53077 = (inp[0]) ? node53081 : node53078;
																assign node53078 = (inp[5]) ? 4'b0001 : 4'b0000;
																assign node53081 = (inp[5]) ? 4'b0000 : 4'b0001;
													assign node53084 = (inp[0]) ? node53096 : node53085;
														assign node53085 = (inp[9]) ? node53091 : node53086;
															assign node53086 = (inp[5]) ? node53088 : 4'b0000;
																assign node53088 = (inp[12]) ? 4'b0001 : 4'b0000;
															assign node53091 = (inp[12]) ? 4'b0000 : node53092;
																assign node53092 = (inp[5]) ? 4'b0000 : 4'b0001;
														assign node53096 = (inp[5]) ? node53100 : node53097;
															assign node53097 = (inp[12]) ? 4'b0001 : 4'b0000;
															assign node53100 = (inp[12]) ? 4'b0000 : 4'b0001;
												assign node53103 = (inp[5]) ? node53111 : node53104;
													assign node53104 = (inp[12]) ? node53108 : node53105;
														assign node53105 = (inp[0]) ? 4'b0000 : 4'b0001;
														assign node53108 = (inp[0]) ? 4'b0001 : 4'b0000;
													assign node53111 = (inp[12]) ? node53115 : node53112;
														assign node53112 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node53115 = (inp[0]) ? 4'b0000 : 4'b0001;
										assign node53118 = (inp[12]) ? node53126 : node53119;
											assign node53119 = (inp[5]) ? node53123 : node53120;
												assign node53120 = (inp[0]) ? 4'b0001 : 4'b0000;
												assign node53123 = (inp[0]) ? 4'b0000 : 4'b0001;
											assign node53126 = (inp[0]) ? node53130 : node53127;
												assign node53127 = (inp[5]) ? 4'b0001 : 4'b0000;
												assign node53130 = (inp[5]) ? 4'b0000 : 4'b0001;
								assign node53133 = (inp[5]) ? node53139 : node53134;
									assign node53134 = (inp[12]) ? 4'b0001 : node53135;
										assign node53135 = (inp[1]) ? 4'b0001 : 4'b0000;
									assign node53139 = (inp[1]) ? 4'b0000 : node53140;
										assign node53140 = (inp[12]) ? 4'b0000 : 4'b0001;
					assign node53144 = (inp[13]) ? node53716 : node53145;
						assign node53145 = (inp[8]) ? node53467 : node53146;
							assign node53146 = (inp[1]) ? node53360 : node53147;
								assign node53147 = (inp[3]) ? node53337 : node53148;
									assign node53148 = (inp[15]) ? node53258 : node53149;
										assign node53149 = (inp[2]) ? node53201 : node53150;
											assign node53150 = (inp[5]) ? node53178 : node53151;
												assign node53151 = (inp[10]) ? node53159 : node53152;
													assign node53152 = (inp[9]) ? node53156 : node53153;
														assign node53153 = (inp[12]) ? 4'b0001 : 4'b0000;
														assign node53156 = (inp[12]) ? 4'b0000 : 4'b0001;
													assign node53159 = (inp[11]) ? node53167 : node53160;
														assign node53160 = (inp[9]) ? node53164 : node53161;
															assign node53161 = (inp[12]) ? 4'b0001 : 4'b0000;
															assign node53164 = (inp[12]) ? 4'b0000 : 4'b0001;
														assign node53167 = (inp[0]) ? node53173 : node53168;
															assign node53168 = (inp[9]) ? 4'b0001 : node53169;
																assign node53169 = (inp[12]) ? 4'b0001 : 4'b0000;
															assign node53173 = (inp[9]) ? node53175 : 4'b0001;
																assign node53175 = (inp[12]) ? 4'b0000 : 4'b0001;
												assign node53178 = (inp[0]) ? node53186 : node53179;
													assign node53179 = (inp[12]) ? node53183 : node53180;
														assign node53180 = (inp[9]) ? 4'b0001 : 4'b0000;
														assign node53183 = (inp[9]) ? 4'b0000 : 4'b0001;
													assign node53186 = (inp[11]) ? node53194 : node53187;
														assign node53187 = (inp[12]) ? node53191 : node53188;
															assign node53188 = (inp[9]) ? 4'b0001 : 4'b0000;
															assign node53191 = (inp[9]) ? 4'b0000 : 4'b0001;
														assign node53194 = (inp[9]) ? node53198 : node53195;
															assign node53195 = (inp[12]) ? 4'b0001 : 4'b0000;
															assign node53198 = (inp[12]) ? 4'b0000 : 4'b0001;
											assign node53201 = (inp[10]) ? node53233 : node53202;
												assign node53202 = (inp[11]) ? node53226 : node53203;
													assign node53203 = (inp[5]) ? node53211 : node53204;
														assign node53204 = (inp[9]) ? node53208 : node53205;
															assign node53205 = (inp[12]) ? 4'b0001 : 4'b0000;
															assign node53208 = (inp[12]) ? 4'b0000 : 4'b0001;
														assign node53211 = (inp[0]) ? node53219 : node53212;
															assign node53212 = (inp[9]) ? node53216 : node53213;
																assign node53213 = (inp[12]) ? 4'b0001 : 4'b0000;
																assign node53216 = (inp[12]) ? 4'b0000 : 4'b0001;
															assign node53219 = (inp[12]) ? node53223 : node53220;
																assign node53220 = (inp[9]) ? 4'b0001 : 4'b0000;
																assign node53223 = (inp[9]) ? 4'b0000 : 4'b0001;
													assign node53226 = (inp[12]) ? node53230 : node53227;
														assign node53227 = (inp[9]) ? 4'b0001 : 4'b0000;
														assign node53230 = (inp[9]) ? 4'b0000 : 4'b0001;
												assign node53233 = (inp[0]) ? node53251 : node53234;
													assign node53234 = (inp[5]) ? node53242 : node53235;
														assign node53235 = (inp[12]) ? node53239 : node53236;
															assign node53236 = (inp[9]) ? 4'b0001 : 4'b0000;
															assign node53239 = (inp[9]) ? 4'b0000 : 4'b0001;
														assign node53242 = (inp[11]) ? node53244 : 4'b0000;
															assign node53244 = (inp[9]) ? node53248 : node53245;
																assign node53245 = (inp[12]) ? 4'b0001 : 4'b0000;
																assign node53248 = (inp[12]) ? 4'b0000 : 4'b0001;
													assign node53251 = (inp[9]) ? node53255 : node53252;
														assign node53252 = (inp[12]) ? 4'b0001 : 4'b0000;
														assign node53255 = (inp[12]) ? 4'b0000 : 4'b0001;
										assign node53258 = (inp[11]) ? node53298 : node53259;
											assign node53259 = (inp[0]) ? node53283 : node53260;
												assign node53260 = (inp[5]) ? node53268 : node53261;
													assign node53261 = (inp[12]) ? node53265 : node53262;
														assign node53262 = (inp[9]) ? 4'b0001 : 4'b0000;
														assign node53265 = (inp[9]) ? 4'b0000 : 4'b0001;
													assign node53268 = (inp[2]) ? node53276 : node53269;
														assign node53269 = (inp[12]) ? node53273 : node53270;
															assign node53270 = (inp[9]) ? 4'b0001 : 4'b0000;
															assign node53273 = (inp[9]) ? 4'b0000 : 4'b0001;
														assign node53276 = (inp[9]) ? node53280 : node53277;
															assign node53277 = (inp[12]) ? 4'b0001 : 4'b0000;
															assign node53280 = (inp[12]) ? 4'b0000 : 4'b0001;
												assign node53283 = (inp[2]) ? node53291 : node53284;
													assign node53284 = (inp[12]) ? node53288 : node53285;
														assign node53285 = (inp[9]) ? 4'b0000 : 4'b0001;
														assign node53288 = (inp[9]) ? 4'b0001 : 4'b0000;
													assign node53291 = (inp[9]) ? node53295 : node53292;
														assign node53292 = (inp[12]) ? 4'b0000 : 4'b0001;
														assign node53295 = (inp[12]) ? 4'b0001 : 4'b0000;
											assign node53298 = (inp[12]) ? node53322 : node53299;
												assign node53299 = (inp[2]) ? node53307 : node53300;
													assign node53300 = (inp[9]) ? node53304 : node53301;
														assign node53301 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node53304 = (inp[0]) ? 4'b0000 : 4'b0001;
													assign node53307 = (inp[10]) ? node53315 : node53308;
														assign node53308 = (inp[0]) ? node53312 : node53309;
															assign node53309 = (inp[9]) ? 4'b0001 : 4'b0000;
															assign node53312 = (inp[9]) ? 4'b0000 : 4'b0001;
														assign node53315 = (inp[9]) ? node53319 : node53316;
															assign node53316 = (inp[0]) ? 4'b0001 : 4'b0000;
															assign node53319 = (inp[0]) ? 4'b0000 : 4'b0001;
												assign node53322 = (inp[2]) ? node53330 : node53323;
													assign node53323 = (inp[9]) ? node53327 : node53324;
														assign node53324 = (inp[0]) ? 4'b0000 : 4'b0001;
														assign node53327 = (inp[0]) ? 4'b0001 : 4'b0000;
													assign node53330 = (inp[0]) ? node53334 : node53331;
														assign node53331 = (inp[9]) ? 4'b0000 : 4'b0001;
														assign node53334 = (inp[9]) ? 4'b0001 : 4'b0000;
									assign node53337 = (inp[12]) ? node53349 : node53338;
										assign node53338 = (inp[9]) ? node53344 : node53339;
											assign node53339 = (inp[15]) ? 4'b0100 : node53340;
												assign node53340 = (inp[0]) ? 4'b0101 : 4'b0100;
											assign node53344 = (inp[15]) ? 4'b0101 : node53345;
												assign node53345 = (inp[0]) ? 4'b0100 : 4'b0101;
										assign node53349 = (inp[9]) ? node53355 : node53350;
											assign node53350 = (inp[15]) ? 4'b0101 : node53351;
												assign node53351 = (inp[0]) ? 4'b0100 : 4'b0101;
											assign node53355 = (inp[0]) ? node53357 : 4'b0100;
												assign node53357 = (inp[15]) ? 4'b0100 : 4'b0101;
								assign node53360 = (inp[12]) ? node53460 : node53361;
									assign node53361 = (inp[5]) ? node53405 : node53362;
										assign node53362 = (inp[0]) ? node53370 : node53363;
											assign node53363 = (inp[9]) ? node53367 : node53364;
												assign node53364 = (inp[15]) ? 4'b0101 : 4'b0100;
												assign node53367 = (inp[15]) ? 4'b0100 : 4'b0101;
											assign node53370 = (inp[10]) ? node53398 : node53371;
												assign node53371 = (inp[3]) ? node53391 : node53372;
													assign node53372 = (inp[11]) ? node53384 : node53373;
														assign node53373 = (inp[2]) ? node53379 : node53374;
															assign node53374 = (inp[15]) ? 4'b0100 : node53375;
																assign node53375 = (inp[9]) ? 4'b0101 : 4'b0100;
															assign node53379 = (inp[9]) ? 4'b0100 : node53380;
																assign node53380 = (inp[15]) ? 4'b0101 : 4'b0100;
														assign node53384 = (inp[15]) ? node53388 : node53385;
															assign node53385 = (inp[9]) ? 4'b0101 : 4'b0100;
															assign node53388 = (inp[9]) ? 4'b0100 : 4'b0101;
													assign node53391 = (inp[9]) ? node53395 : node53392;
														assign node53392 = (inp[15]) ? 4'b0101 : 4'b0100;
														assign node53395 = (inp[15]) ? 4'b0100 : 4'b0101;
												assign node53398 = (inp[9]) ? node53402 : node53399;
													assign node53399 = (inp[15]) ? 4'b0101 : 4'b0100;
													assign node53402 = (inp[15]) ? 4'b0100 : 4'b0101;
										assign node53405 = (inp[11]) ? node53413 : node53406;
											assign node53406 = (inp[15]) ? node53410 : node53407;
												assign node53407 = (inp[9]) ? 4'b0101 : 4'b0100;
												assign node53410 = (inp[9]) ? 4'b0100 : 4'b0101;
											assign node53413 = (inp[0]) ? node53437 : node53414;
												assign node53414 = (inp[2]) ? node53422 : node53415;
													assign node53415 = (inp[15]) ? node53419 : node53416;
														assign node53416 = (inp[9]) ? 4'b0101 : 4'b0100;
														assign node53419 = (inp[9]) ? 4'b0100 : 4'b0101;
													assign node53422 = (inp[10]) ? node53430 : node53423;
														assign node53423 = (inp[9]) ? node53427 : node53424;
															assign node53424 = (inp[15]) ? 4'b0101 : 4'b0100;
															assign node53427 = (inp[15]) ? 4'b0100 : 4'b0101;
														assign node53430 = (inp[9]) ? node53434 : node53431;
															assign node53431 = (inp[15]) ? 4'b0101 : 4'b0100;
															assign node53434 = (inp[15]) ? 4'b0100 : 4'b0101;
												assign node53437 = (inp[10]) ? node53445 : node53438;
													assign node53438 = (inp[9]) ? node53442 : node53439;
														assign node53439 = (inp[15]) ? 4'b0101 : 4'b0100;
														assign node53442 = (inp[15]) ? 4'b0100 : 4'b0101;
													assign node53445 = (inp[3]) ? node53453 : node53446;
														assign node53446 = (inp[15]) ? node53450 : node53447;
															assign node53447 = (inp[9]) ? 4'b0101 : 4'b0100;
															assign node53450 = (inp[9]) ? 4'b0100 : 4'b0101;
														assign node53453 = (inp[9]) ? node53457 : node53454;
															assign node53454 = (inp[15]) ? 4'b0101 : 4'b0100;
															assign node53457 = (inp[15]) ? 4'b0100 : 4'b0101;
									assign node53460 = (inp[9]) ? node53464 : node53461;
										assign node53461 = (inp[15]) ? 4'b0101 : 4'b0100;
										assign node53464 = (inp[15]) ? 4'b0100 : 4'b0101;
							assign node53467 = (inp[1]) ? node53705 : node53468;
								assign node53468 = (inp[3]) ? node53698 : node53469;
									assign node53469 = (inp[11]) ? node53577 : node53470;
										assign node53470 = (inp[2]) ? node53508 : node53471;
											assign node53471 = (inp[9]) ? node53501 : node53472;
												assign node53472 = (inp[10]) ? node53480 : node53473;
													assign node53473 = (inp[12]) ? node53477 : node53474;
														assign node53474 = (inp[0]) ? 4'b0101 : 4'b0100;
														assign node53477 = (inp[0]) ? 4'b0100 : 4'b0101;
													assign node53480 = (inp[5]) ? node53490 : node53481;
														assign node53481 = (inp[15]) ? 4'b0100 : node53482;
															assign node53482 = (inp[0]) ? node53486 : node53483;
																assign node53483 = (inp[12]) ? 4'b0101 : 4'b0100;
																assign node53486 = (inp[12]) ? 4'b0100 : 4'b0101;
														assign node53490 = (inp[15]) ? node53496 : node53491;
															assign node53491 = (inp[12]) ? 4'b0100 : node53492;
																assign node53492 = (inp[0]) ? 4'b0101 : 4'b0100;
															assign node53496 = (inp[12]) ? node53498 : 4'b0101;
																assign node53498 = (inp[0]) ? 4'b0100 : 4'b0101;
												assign node53501 = (inp[0]) ? node53505 : node53502;
													assign node53502 = (inp[12]) ? 4'b0101 : 4'b0100;
													assign node53505 = (inp[12]) ? 4'b0100 : 4'b0101;
											assign node53508 = (inp[15]) ? node53554 : node53509;
												assign node53509 = (inp[5]) ? node53531 : node53510;
													assign node53510 = (inp[10]) ? node53524 : node53511;
														assign node53511 = (inp[9]) ? node53517 : node53512;
															assign node53512 = (inp[12]) ? 4'b0100 : node53513;
																assign node53513 = (inp[0]) ? 4'b0101 : 4'b0100;
															assign node53517 = (inp[12]) ? node53521 : node53518;
																assign node53518 = (inp[0]) ? 4'b0101 : 4'b0100;
																assign node53521 = (inp[0]) ? 4'b0100 : 4'b0101;
														assign node53524 = (inp[0]) ? node53528 : node53525;
															assign node53525 = (inp[12]) ? 4'b0101 : 4'b0100;
															assign node53528 = (inp[12]) ? 4'b0100 : 4'b0101;
													assign node53531 = (inp[9]) ? node53539 : node53532;
														assign node53532 = (inp[0]) ? node53536 : node53533;
															assign node53533 = (inp[12]) ? 4'b0101 : 4'b0100;
															assign node53536 = (inp[12]) ? 4'b0100 : 4'b0101;
														assign node53539 = (inp[10]) ? node53547 : node53540;
															assign node53540 = (inp[12]) ? node53544 : node53541;
																assign node53541 = (inp[0]) ? 4'b0101 : 4'b0100;
																assign node53544 = (inp[0]) ? 4'b0100 : 4'b0101;
															assign node53547 = (inp[12]) ? node53551 : node53548;
																assign node53548 = (inp[0]) ? 4'b0101 : 4'b0100;
																assign node53551 = (inp[0]) ? 4'b0100 : 4'b0101;
												assign node53554 = (inp[5]) ? node53570 : node53555;
													assign node53555 = (inp[9]) ? node53563 : node53556;
														assign node53556 = (inp[0]) ? node53560 : node53557;
															assign node53557 = (inp[12]) ? 4'b0101 : 4'b0100;
															assign node53560 = (inp[12]) ? 4'b0100 : 4'b0101;
														assign node53563 = (inp[0]) ? node53567 : node53564;
															assign node53564 = (inp[12]) ? 4'b0101 : 4'b0100;
															assign node53567 = (inp[12]) ? 4'b0100 : 4'b0101;
													assign node53570 = (inp[0]) ? node53574 : node53571;
														assign node53571 = (inp[12]) ? 4'b0101 : 4'b0100;
														assign node53574 = (inp[12]) ? 4'b0100 : 4'b0101;
										assign node53577 = (inp[2]) ? node53633 : node53578;
											assign node53578 = (inp[15]) ? node53602 : node53579;
												assign node53579 = (inp[5]) ? node53587 : node53580;
													assign node53580 = (inp[0]) ? node53584 : node53581;
														assign node53581 = (inp[12]) ? 4'b0101 : 4'b0100;
														assign node53584 = (inp[12]) ? 4'b0100 : 4'b0101;
													assign node53587 = (inp[9]) ? node53595 : node53588;
														assign node53588 = (inp[12]) ? node53592 : node53589;
															assign node53589 = (inp[0]) ? 4'b0101 : 4'b0100;
															assign node53592 = (inp[0]) ? 4'b0100 : 4'b0101;
														assign node53595 = (inp[0]) ? node53599 : node53596;
															assign node53596 = (inp[12]) ? 4'b0101 : 4'b0100;
															assign node53599 = (inp[12]) ? 4'b0100 : 4'b0101;
												assign node53602 = (inp[9]) ? node53618 : node53603;
													assign node53603 = (inp[5]) ? node53611 : node53604;
														assign node53604 = (inp[0]) ? node53608 : node53605;
															assign node53605 = (inp[12]) ? 4'b0101 : 4'b0100;
															assign node53608 = (inp[12]) ? 4'b0100 : 4'b0101;
														assign node53611 = (inp[0]) ? node53615 : node53612;
															assign node53612 = (inp[12]) ? 4'b0101 : 4'b0100;
															assign node53615 = (inp[12]) ? 4'b0100 : 4'b0101;
													assign node53618 = (inp[10]) ? node53626 : node53619;
														assign node53619 = (inp[0]) ? node53623 : node53620;
															assign node53620 = (inp[12]) ? 4'b0101 : 4'b0100;
															assign node53623 = (inp[12]) ? 4'b0100 : 4'b0101;
														assign node53626 = (inp[0]) ? node53630 : node53627;
															assign node53627 = (inp[12]) ? 4'b0101 : 4'b0100;
															assign node53630 = (inp[12]) ? 4'b0100 : 4'b0101;
											assign node53633 = (inp[10]) ? node53641 : node53634;
												assign node53634 = (inp[12]) ? node53638 : node53635;
													assign node53635 = (inp[0]) ? 4'b0101 : 4'b0100;
													assign node53638 = (inp[0]) ? 4'b0100 : 4'b0101;
												assign node53641 = (inp[5]) ? node53667 : node53642;
													assign node53642 = (inp[15]) ? node53654 : node53643;
														assign node53643 = (inp[9]) ? node53649 : node53644;
															assign node53644 = (inp[12]) ? node53646 : 4'b0100;
																assign node53646 = (inp[0]) ? 4'b0100 : 4'b0101;
															assign node53649 = (inp[0]) ? 4'b0101 : node53650;
																assign node53650 = (inp[12]) ? 4'b0101 : 4'b0100;
														assign node53654 = (inp[9]) ? node53662 : node53655;
															assign node53655 = (inp[12]) ? node53659 : node53656;
																assign node53656 = (inp[0]) ? 4'b0101 : 4'b0100;
																assign node53659 = (inp[0]) ? 4'b0100 : 4'b0101;
															assign node53662 = (inp[12]) ? 4'b0100 : node53663;
																assign node53663 = (inp[0]) ? 4'b0101 : 4'b0100;
													assign node53667 = (inp[15]) ? node53683 : node53668;
														assign node53668 = (inp[9]) ? node53676 : node53669;
															assign node53669 = (inp[12]) ? node53673 : node53670;
																assign node53670 = (inp[0]) ? 4'b0101 : 4'b0100;
																assign node53673 = (inp[0]) ? 4'b0100 : 4'b0101;
															assign node53676 = (inp[0]) ? node53680 : node53677;
																assign node53677 = (inp[12]) ? 4'b0101 : 4'b0100;
																assign node53680 = (inp[12]) ? 4'b0100 : 4'b0101;
														assign node53683 = (inp[9]) ? node53691 : node53684;
															assign node53684 = (inp[0]) ? node53688 : node53685;
																assign node53685 = (inp[12]) ? 4'b0101 : 4'b0100;
																assign node53688 = (inp[12]) ? 4'b0100 : 4'b0101;
															assign node53691 = (inp[12]) ? node53695 : node53692;
																assign node53692 = (inp[0]) ? 4'b0101 : 4'b0100;
																assign node53695 = (inp[0]) ? 4'b0100 : 4'b0101;
									assign node53698 = (inp[15]) ? node53702 : node53699;
										assign node53699 = (inp[12]) ? 4'b0001 : 4'b0000;
										assign node53702 = (inp[12]) ? 4'b0000 : 4'b0001;
								assign node53705 = (inp[15]) ? node53711 : node53706;
									assign node53706 = (inp[3]) ? 4'b0001 : node53707;
										assign node53707 = (inp[0]) ? 4'b0001 : 4'b0000;
									assign node53711 = (inp[0]) ? 4'b0000 : node53712;
										assign node53712 = (inp[3]) ? 4'b0000 : 4'b0001;
						assign node53716 = (inp[1]) ? node53832 : node53717;
							assign node53717 = (inp[3]) ? node53805 : node53718;
								assign node53718 = (inp[0]) ? node53794 : node53719;
									assign node53719 = (inp[12]) ? node53777 : node53720;
										assign node53720 = (inp[8]) ? 4'b0100 : node53721;
											assign node53721 = (inp[10]) ? node53761 : node53722;
												assign node53722 = (inp[2]) ? node53746 : node53723;
													assign node53723 = (inp[11]) ? node53731 : node53724;
														assign node53724 = (inp[9]) ? node53728 : node53725;
															assign node53725 = (inp[15]) ? 4'b0101 : 4'b0100;
															assign node53728 = (inp[15]) ? 4'b0100 : 4'b0101;
														assign node53731 = (inp[5]) ? node53739 : node53732;
															assign node53732 = (inp[15]) ? node53736 : node53733;
																assign node53733 = (inp[9]) ? 4'b0101 : 4'b0100;
																assign node53736 = (inp[9]) ? 4'b0100 : 4'b0101;
															assign node53739 = (inp[15]) ? node53743 : node53740;
																assign node53740 = (inp[9]) ? 4'b0101 : 4'b0100;
																assign node53743 = (inp[9]) ? 4'b0100 : 4'b0101;
													assign node53746 = (inp[5]) ? node53754 : node53747;
														assign node53747 = (inp[9]) ? node53751 : node53748;
															assign node53748 = (inp[15]) ? 4'b0101 : 4'b0100;
															assign node53751 = (inp[15]) ? 4'b0100 : 4'b0101;
														assign node53754 = (inp[15]) ? node53758 : node53755;
															assign node53755 = (inp[9]) ? 4'b0101 : 4'b0100;
															assign node53758 = (inp[9]) ? 4'b0100 : 4'b0101;
												assign node53761 = (inp[2]) ? node53769 : node53762;
													assign node53762 = (inp[9]) ? node53766 : node53763;
														assign node53763 = (inp[15]) ? 4'b0101 : 4'b0100;
														assign node53766 = (inp[15]) ? 4'b0100 : 4'b0101;
													assign node53769 = (inp[9]) ? node53773 : node53770;
														assign node53770 = (inp[15]) ? 4'b0101 : 4'b0100;
														assign node53773 = (inp[15]) ? 4'b0100 : 4'b0101;
										assign node53777 = (inp[8]) ? 4'b0101 : node53778;
											assign node53778 = (inp[5]) ? node53786 : node53779;
												assign node53779 = (inp[15]) ? node53783 : node53780;
													assign node53780 = (inp[9]) ? 4'b0100 : 4'b0101;
													assign node53783 = (inp[9]) ? 4'b0101 : 4'b0100;
												assign node53786 = (inp[9]) ? node53790 : node53787;
													assign node53787 = (inp[15]) ? 4'b0100 : 4'b0101;
													assign node53790 = (inp[15]) ? 4'b0101 : 4'b0100;
									assign node53794 = (inp[12]) ? node53800 : node53795;
										assign node53795 = (inp[9]) ? 4'b0101 : node53796;
											assign node53796 = (inp[8]) ? 4'b0101 : 4'b0100;
										assign node53800 = (inp[8]) ? 4'b0100 : node53801;
											assign node53801 = (inp[9]) ? 4'b0100 : 4'b0101;
								assign node53805 = (inp[12]) ? node53819 : node53806;
									assign node53806 = (inp[8]) ? 4'b0001 : node53807;
										assign node53807 = (inp[9]) ? node53813 : node53808;
											assign node53808 = (inp[0]) ? 4'b0000 : node53809;
												assign node53809 = (inp[15]) ? 4'b0000 : 4'b0001;
											assign node53813 = (inp[15]) ? 4'b0001 : node53814;
												assign node53814 = (inp[0]) ? 4'b0001 : 4'b0000;
									assign node53819 = (inp[8]) ? 4'b0000 : node53820;
										assign node53820 = (inp[9]) ? node53826 : node53821;
											assign node53821 = (inp[15]) ? 4'b0001 : node53822;
												assign node53822 = (inp[0]) ? 4'b0001 : 4'b0000;
											assign node53826 = (inp[15]) ? 4'b0000 : node53827;
												assign node53827 = (inp[0]) ? 4'b0000 : 4'b0001;
							assign node53832 = (inp[0]) ? node53844 : node53833;
								assign node53833 = (inp[3]) ? node53839 : node53834;
									assign node53834 = (inp[8]) ? 4'b0001 : node53835;
										assign node53835 = (inp[9]) ? 4'b0001 : 4'b0000;
									assign node53839 = (inp[8]) ? 4'b0000 : node53840;
										assign node53840 = (inp[9]) ? 4'b0000 : 4'b0001;
								assign node53844 = (inp[8]) ? 4'b0000 : node53845;
									assign node53845 = (inp[9]) ? 4'b0000 : 4'b0001;

endmodule