module dtc_split33_bm14 (
	input  wire [13-1:0] inp,
	output wire [1-1:0] outp
);

	wire [1-1:0] node1;
	wire [1-1:0] node2;
	wire [1-1:0] node3;
	wire [1-1:0] node4;
	wire [1-1:0] node6;
	wire [1-1:0] node8;
	wire [1-1:0] node9;
	wire [1-1:0] node11;
	wire [1-1:0] node13;
	wire [1-1:0] node15;
	wire [1-1:0] node18;
	wire [1-1:0] node19;
	wire [1-1:0] node21;
	wire [1-1:0] node23;
	wire [1-1:0] node26;
	wire [1-1:0] node27;
	wire [1-1:0] node29;
	wire [1-1:0] node31;
	wire [1-1:0] node34;
	wire [1-1:0] node35;
	wire [1-1:0] node39;
	wire [1-1:0] node40;
	wire [1-1:0] node41;
	wire [1-1:0] node43;
	wire [1-1:0] node45;
	wire [1-1:0] node47;
	wire [1-1:0] node49;
	wire [1-1:0] node52;
	wire [1-1:0] node53;
	wire [1-1:0] node55;
	wire [1-1:0] node57;
	wire [1-1:0] node60;
	wire [1-1:0] node62;
	wire [1-1:0] node63;
	wire [1-1:0] node65;
	wire [1-1:0] node68;
	wire [1-1:0] node69;
	wire [1-1:0] node73;
	wire [1-1:0] node74;
	wire [1-1:0] node75;
	wire [1-1:0] node77;
	wire [1-1:0] node79;
	wire [1-1:0] node81;
	wire [1-1:0] node82;
	wire [1-1:0] node84;
	wire [1-1:0] node88;
	wire [1-1:0] node90;
	wire [1-1:0] node91;
	wire [1-1:0] node93;
	wire [1-1:0] node94;
	wire [1-1:0] node99;
	wire [1-1:0] node100;
	wire [1-1:0] node101;
	wire [1-1:0] node103;
	wire [1-1:0] node105;
	wire [1-1:0] node108;
	wire [1-1:0] node109;
	wire [1-1:0] node111;
	wire [1-1:0] node114;
	wire [1-1:0] node115;
	wire [1-1:0] node119;
	wire [1-1:0] node120;
	wire [1-1:0] node122;
	wire [1-1:0] node123;
	wire [1-1:0] node128;
	wire [1-1:0] node129;
	wire [1-1:0] node130;
	wire [1-1:0] node132;
	wire [1-1:0] node134;
	wire [1-1:0] node136;
	wire [1-1:0] node137;
	wire [1-1:0] node139;
	wire [1-1:0] node142;
	wire [1-1:0] node143;
	wire [1-1:0] node147;
	wire [1-1:0] node148;
	wire [1-1:0] node150;
	wire [1-1:0] node151;
	wire [1-1:0] node153;
	wire [1-1:0] node156;
	wire [1-1:0] node158;
	wire [1-1:0] node159;
	wire [1-1:0] node163;
	wire [1-1:0] node164;
	wire [1-1:0] node166;
	wire [1-1:0] node167;
	wire [1-1:0] node169;
	wire [1-1:0] node170;
	wire [1-1:0] node172;
	wire [1-1:0] node176;
	wire [1-1:0] node177;
	wire [1-1:0] node181;
	wire [1-1:0] node182;
	wire [1-1:0] node184;
	wire [1-1:0] node185;
	wire [1-1:0] node189;
	wire [1-1:0] node190;
	wire [1-1:0] node191;
	wire [1-1:0] node193;
	wire [1-1:0] node194;
	wire [1-1:0] node200;
	wire [1-1:0] node201;
	wire [1-1:0] node202;
	wire [1-1:0] node204;
	wire [1-1:0] node205;
	wire [1-1:0] node207;
	wire [1-1:0] node210;
	wire [1-1:0] node211;
	wire [1-1:0] node213;
	wire [1-1:0] node217;
	wire [1-1:0] node218;
	wire [1-1:0] node220;
	wire [1-1:0] node221;
	wire [1-1:0] node223;
	wire [1-1:0] node227;
	wire [1-1:0] node228;
	wire [1-1:0] node230;
	wire [1-1:0] node231;
	wire [1-1:0] node236;
	wire [1-1:0] node237;
	wire [1-1:0] node238;
	wire [1-1:0] node240;
	wire [1-1:0] node241;
	wire [1-1:0] node244;
	wire [1-1:0] node246;
	wire [1-1:0] node247;
	wire [1-1:0] node251;
	wire [1-1:0] node252;
	wire [1-1:0] node254;
	wire [1-1:0] node255;
	wire [1-1:0] node259;
	wire [1-1:0] node260;
	wire [1-1:0] node261;
	wire [1-1:0] node266;
	wire [1-1:0] node267;
	wire [1-1:0] node268;
	wire [1-1:0] node269;
	wire [1-1:0] node272;
	wire [1-1:0] node273;
	wire [1-1:0] node279;
	wire [1-1:0] node280;
	wire [1-1:0] node281;
	wire [1-1:0] node282;
	wire [1-1:0] node284;
	wire [1-1:0] node285;
	wire [1-1:0] node287;
	wire [1-1:0] node289;
	wire [1-1:0] node292;
	wire [1-1:0] node293;
	wire [1-1:0] node295;
	wire [1-1:0] node297;
	wire [1-1:0] node300;
	wire [1-1:0] node301;
	wire [1-1:0] node303;
	wire [1-1:0] node306;
	wire [1-1:0] node307;
	wire [1-1:0] node311;
	wire [1-1:0] node312;
	wire [1-1:0] node314;
	wire [1-1:0] node315;
	wire [1-1:0] node317;
	wire [1-1:0] node320;
	wire [1-1:0] node321;
	wire [1-1:0] node325;
	wire [1-1:0] node326;
	wire [1-1:0] node328;
	wire [1-1:0] node330;
	wire [1-1:0] node331;
	wire [1-1:0] node335;
	wire [1-1:0] node336;
	wire [1-1:0] node338;
	wire [1-1:0] node339;
	wire [1-1:0] node344;
	wire [1-1:0] node345;
	wire [1-1:0] node346;
	wire [1-1:0] node348;
	wire [1-1:0] node349;
	wire [1-1:0] node351;
	wire [1-1:0] node353;
	wire [1-1:0] node356;
	wire [1-1:0] node357;
	wire [1-1:0] node359;
	wire [1-1:0] node363;
	wire [1-1:0] node364;
	wire [1-1:0] node365;
	wire [1-1:0] node367;
	wire [1-1:0] node369;
	wire [1-1:0] node372;
	wire [1-1:0] node373;
	wire [1-1:0] node375;
	wire [1-1:0] node379;
	wire [1-1:0] node380;
	wire [1-1:0] node381;
	wire [1-1:0] node383;
	wire [1-1:0] node386;
	wire [1-1:0] node387;
	wire [1-1:0] node391;
	wire [1-1:0] node392;
	wire [1-1:0] node393;
	wire [1-1:0] node394;
	wire [1-1:0] node400;
	wire [1-1:0] node401;
	wire [1-1:0] node402;
	wire [1-1:0] node403;
	wire [1-1:0] node405;
	wire [1-1:0] node407;
	wire [1-1:0] node409;
	wire [1-1:0] node412;
	wire [1-1:0] node413;
	wire [1-1:0] node415;
	wire [1-1:0] node416;
	wire [1-1:0] node421;
	wire [1-1:0] node422;
	wire [1-1:0] node423;
	wire [1-1:0] node425;
	wire [1-1:0] node428;
	wire [1-1:0] node429;
	wire [1-1:0] node431;
	wire [1-1:0] node435;
	wire [1-1:0] node436;
	wire [1-1:0] node437;
	wire [1-1:0] node438;
	wire [1-1:0] node444;
	wire [1-1:0] node445;
	wire [1-1:0] node446;
	wire [1-1:0] node447;
	wire [1-1:0] node449;
	wire [1-1:0] node451;
	wire [1-1:0] node452;
	wire [1-1:0] node456;
	wire [1-1:0] node457;
	wire [1-1:0] node462;
	wire [1-1:0] node463;
	wire [1-1:0] node464;
	wire [1-1:0] node469;
	wire [1-1:0] node470;
	wire [1-1:0] node471;
	wire [1-1:0] node472;
	wire [1-1:0] node474;
	wire [1-1:0] node475;
	wire [1-1:0] node477;
	wire [1-1:0] node479;
	wire [1-1:0] node482;
	wire [1-1:0] node483;
	wire [1-1:0] node485;
	wire [1-1:0] node489;
	wire [1-1:0] node490;
	wire [1-1:0] node492;
	wire [1-1:0] node493;
	wire [1-1:0] node495;
	wire [1-1:0] node498;
	wire [1-1:0] node499;
	wire [1-1:0] node503;
	wire [1-1:0] node504;
	wire [1-1:0] node506;
	wire [1-1:0] node508;
	wire [1-1:0] node509;
	wire [1-1:0] node510;
	wire [1-1:0] node515;
	wire [1-1:0] node516;
	wire [1-1:0] node520;
	wire [1-1:0] node521;
	wire [1-1:0] node522;
	wire [1-1:0] node523;
	wire [1-1:0] node525;
	wire [1-1:0] node527;
	wire [1-1:0] node530;
	wire [1-1:0] node531;
	wire [1-1:0] node534;
	wire [1-1:0] node535;
	wire [1-1:0] node537;
	wire [1-1:0] node541;
	wire [1-1:0] node542;
	wire [1-1:0] node543;
	wire [1-1:0] node545;
	wire [1-1:0] node546;
	wire [1-1:0] node550;
	wire [1-1:0] node551;
	wire [1-1:0] node552;
	wire [1-1:0] node554;
	wire [1-1:0] node560;
	wire [1-1:0] node561;
	wire [1-1:0] node562;
	wire [1-1:0] node563;
	wire [1-1:0] node565;
	wire [1-1:0] node568;
	wire [1-1:0] node569;
	wire [1-1:0] node573;
	wire [1-1:0] node574;
	wire [1-1:0] node579;
	wire [1-1:0] node580;
	wire [1-1:0] node581;
	wire [1-1:0] node582;
	wire [1-1:0] node583;
	wire [1-1:0] node585;
	wire [1-1:0] node587;
	wire [1-1:0] node590;
	wire [1-1:0] node591;
	wire [1-1:0] node593;
	wire [1-1:0] node597;
	wire [1-1:0] node598;
	wire [1-1:0] node599;
	wire [1-1:0] node602;
	wire [1-1:0] node603;
	wire [1-1:0] node607;
	wire [1-1:0] node608;
	wire [1-1:0] node612;
	wire [1-1:0] node613;
	wire [1-1:0] node614;
	wire [1-1:0] node616;
	wire [1-1:0] node619;
	wire [1-1:0] node620;
	wire [1-1:0] node621;
	wire [1-1:0] node626;
	wire [1-1:0] node627;
	wire [1-1:0] node628;
	wire [1-1:0] node629;
	wire [1-1:0] node635;
	wire [1-1:0] node636;
	wire [1-1:0] node637;
	wire [1-1:0] node638;
	wire [1-1:0] node639;
	wire [1-1:0] node641;
	wire [1-1:0] node648;
	wire [1-1:0] node649;
	wire [1-1:0] node650;
	wire [1-1:0] node651;
	wire [1-1:0] node652;
	wire [1-1:0] node654;
	wire [1-1:0] node656;
	wire [1-1:0] node657;
	wire [1-1:0] node659;
	wire [1-1:0] node662;
	wire [1-1:0] node663;
	wire [1-1:0] node665;
	wire [1-1:0] node666;
	wire [1-1:0] node671;
	wire [1-1:0] node672;
	wire [1-1:0] node673;
	wire [1-1:0] node675;
	wire [1-1:0] node677;
	wire [1-1:0] node680;
	wire [1-1:0] node681;
	wire [1-1:0] node683;
	wire [1-1:0] node685;
	wire [1-1:0] node686;
	wire [1-1:0] node690;
	wire [1-1:0] node691;
	wire [1-1:0] node694;
	wire [1-1:0] node695;
	wire [1-1:0] node699;
	wire [1-1:0] node700;
	wire [1-1:0] node701;
	wire [1-1:0] node703;
	wire [1-1:0] node705;
	wire [1-1:0] node708;
	wire [1-1:0] node709;
	wire [1-1:0] node711;
	wire [1-1:0] node715;
	wire [1-1:0] node716;
	wire [1-1:0] node717;
	wire [1-1:0] node719;
	wire [1-1:0] node721;
	wire [1-1:0] node722;
	wire [1-1:0] node726;
	wire [1-1:0] node727;
	wire [1-1:0] node732;
	wire [1-1:0] node733;
	wire [1-1:0] node734;
	wire [1-1:0] node735;
	wire [1-1:0] node737;
	wire [1-1:0] node739;
	wire [1-1:0] node741;
	wire [1-1:0] node744;
	wire [1-1:0] node745;
	wire [1-1:0] node747;
	wire [1-1:0] node749;
	wire [1-1:0] node752;
	wire [1-1:0] node753;
	wire [1-1:0] node754;
	wire [1-1:0] node759;
	wire [1-1:0] node760;
	wire [1-1:0] node761;
	wire [1-1:0] node763;
	wire [1-1:0] node765;
	wire [1-1:0] node768;
	wire [1-1:0] node769;
	wire [1-1:0] node771;
	wire [1-1:0] node775;
	wire [1-1:0] node776;
	wire [1-1:0] node777;
	wire [1-1:0] node779;
	wire [1-1:0] node782;
	wire [1-1:0] node783;
	wire [1-1:0] node788;
	wire [1-1:0] node789;
	wire [1-1:0] node790;
	wire [1-1:0] node792;
	wire [1-1:0] node793;
	wire [1-1:0] node795;
	wire [1-1:0] node798;
	wire [1-1:0] node799;
	wire [1-1:0] node800;
	wire [1-1:0] node802;
	wire [1-1:0] node807;
	wire [1-1:0] node808;
	wire [1-1:0] node810;
	wire [1-1:0] node811;
	wire [1-1:0] node815;
	wire [1-1:0] node816;
	wire [1-1:0] node817;
	wire [1-1:0] node822;
	wire [1-1:0] node823;
	wire [1-1:0] node824;
	wire [1-1:0] node826;
	wire [1-1:0] node827;
	wire [1-1:0] node829;
	wire [1-1:0] node833;
	wire [1-1:0] node834;
	wire [1-1:0] node835;
	wire [1-1:0] node840;
	wire [1-1:0] node841;
	wire [1-1:0] node842;
	wire [1-1:0] node847;
	wire [1-1:0] node848;
	wire [1-1:0] node849;
	wire [1-1:0] node850;
	wire [1-1:0] node852;
	wire [1-1:0] node853;
	wire [1-1:0] node855;
	wire [1-1:0] node858;
	wire [1-1:0] node859;
	wire [1-1:0] node863;
	wire [1-1:0] node864;
	wire [1-1:0] node865;
	wire [1-1:0] node867;
	wire [1-1:0] node870;
	wire [1-1:0] node872;
	wire [1-1:0] node873;
	wire [1-1:0] node877;
	wire [1-1:0] node878;
	wire [1-1:0] node879;
	wire [1-1:0] node881;
	wire [1-1:0] node882;
	wire [1-1:0] node884;
	wire [1-1:0] node888;
	wire [1-1:0] node889;
	wire [1-1:0] node893;
	wire [1-1:0] node894;
	wire [1-1:0] node896;
	wire [1-1:0] node900;
	wire [1-1:0] node901;
	wire [1-1:0] node902;
	wire [1-1:0] node904;
	wire [1-1:0] node906;
	wire [1-1:0] node907;
	wire [1-1:0] node911;
	wire [1-1:0] node912;
	wire [1-1:0] node913;
	wire [1-1:0] node915;
	wire [1-1:0] node918;
	wire [1-1:0] node921;
	wire [1-1:0] node922;
	wire [1-1:0] node923;
	wire [1-1:0] node928;
	wire [1-1:0] node929;
	wire [1-1:0] node930;
	wire [1-1:0] node931;
	wire [1-1:0] node933;
	wire [1-1:0] node936;
	wire [1-1:0] node937;
	wire [1-1:0] node943;
	wire [1-1:0] node944;
	wire [1-1:0] node945;
	wire [1-1:0] node946;
	wire [1-1:0] node948;
	wire [1-1:0] node950;
	wire [1-1:0] node951;
	wire [1-1:0] node955;
	wire [1-1:0] node956;
	wire [1-1:0] node957;
	wire [1-1:0] node961;
	wire [1-1:0] node962;
	wire [1-1:0] node966;
	wire [1-1:0] node967;
	wire [1-1:0] node968;
	wire [1-1:0] node969;
	wire [1-1:0] node971;
	wire [1-1:0] node974;
	wire [1-1:0] node975;
	wire [1-1:0] node979;
	wire [1-1:0] node980;
	wire [1-1:0] node981;
	wire [1-1:0] node986;
	wire [1-1:0] node987;
	wire [1-1:0] node988;
	wire [1-1:0] node993;
	wire [1-1:0] node994;
	wire [1-1:0] node995;
	wire [1-1:0] node996;
	wire [1-1:0] node998;
	wire [1-1:0] node999;
	wire [1-1:0] node1003;
	wire [1-1:0] node1004;
	wire [1-1:0] node1005;
	wire [1-1:0] node1012;
	wire [1-1:0] node1013;
	wire [1-1:0] node1014;
	wire [1-1:0] node1015;
	wire [1-1:0] node1016;
	wire [1-1:0] node1017;
	wire [1-1:0] node1018;
	wire [1-1:0] node1020;
	wire [1-1:0] node1022;
	wire [1-1:0] node1024;
	wire [1-1:0] node1028;
	wire [1-1:0] node1029;
	wire [1-1:0] node1031;
	wire [1-1:0] node1033;
	wire [1-1:0] node1036;
	wire [1-1:0] node1037;
	wire [1-1:0] node1041;
	wire [1-1:0] node1042;
	wire [1-1:0] node1044;
	wire [1-1:0] node1045;
	wire [1-1:0] node1047;
	wire [1-1:0] node1051;
	wire [1-1:0] node1052;
	wire [1-1:0] node1054;
	wire [1-1:0] node1055;
	wire [1-1:0] node1060;
	wire [1-1:0] node1061;
	wire [1-1:0] node1062;
	wire [1-1:0] node1063;
	wire [1-1:0] node1065;
	wire [1-1:0] node1067;
	wire [1-1:0] node1070;
	wire [1-1:0] node1071;
	wire [1-1:0] node1073;
	wire [1-1:0] node1076;
	wire [1-1:0] node1077;
	wire [1-1:0] node1081;
	wire [1-1:0] node1082;
	wire [1-1:0] node1083;
	wire [1-1:0] node1085;
	wire [1-1:0] node1088;
	wire [1-1:0] node1089;
	wire [1-1:0] node1094;
	wire [1-1:0] node1095;
	wire [1-1:0] node1096;
	wire [1-1:0] node1097;
	wire [1-1:0] node1099;
	wire [1-1:0] node1102;
	wire [1-1:0] node1103;
	wire [1-1:0] node1104;
	wire [1-1:0] node1110;
	wire [1-1:0] node1111;
	wire [1-1:0] node1112;
	wire [1-1:0] node1113;
	wire [1-1:0] node1119;
	wire [1-1:0] node1120;
	wire [1-1:0] node1121;
	wire [1-1:0] node1122;
	wire [1-1:0] node1124;
	wire [1-1:0] node1126;
	wire [1-1:0] node1129;
	wire [1-1:0] node1130;
	wire [1-1:0] node1132;
	wire [1-1:0] node1133;
	wire [1-1:0] node1135;
	wire [1-1:0] node1139;
	wire [1-1:0] node1140;
	wire [1-1:0] node1144;
	wire [1-1:0] node1145;
	wire [1-1:0] node1146;
	wire [1-1:0] node1148;
	wire [1-1:0] node1149;
	wire [1-1:0] node1154;
	wire [1-1:0] node1155;
	wire [1-1:0] node1156;
	wire [1-1:0] node1161;
	wire [1-1:0] node1162;
	wire [1-1:0] node1163;
	wire [1-1:0] node1164;
	wire [1-1:0] node1165;
	wire [1-1:0] node1167;
	wire [1-1:0] node1170;
	wire [1-1:0] node1171;
	wire [1-1:0] node1175;
	wire [1-1:0] node1176;
	wire [1-1:0] node1177;
	wire [1-1:0] node1182;
	wire [1-1:0] node1183;
	wire [1-1:0] node1184;
	wire [1-1:0] node1189;
	wire [1-1:0] node1190;
	wire [1-1:0] node1191;
	wire [1-1:0] node1192;
	wire [1-1:0] node1198;
	wire [1-1:0] node1199;
	wire [1-1:0] node1200;
	wire [1-1:0] node1201;
	wire [1-1:0] node1202;
	wire [1-1:0] node1203;
	wire [1-1:0] node1205;
	wire [1-1:0] node1208;
	wire [1-1:0] node1209;
	wire [1-1:0] node1211;
	wire [1-1:0] node1212;
	wire [1-1:0] node1217;
	wire [1-1:0] node1218;
	wire [1-1:0] node1219;
	wire [1-1:0] node1221;
	wire [1-1:0] node1226;
	wire [1-1:0] node1227;
	wire [1-1:0] node1228;
	wire [1-1:0] node1229;
	wire [1-1:0] node1231;
	wire [1-1:0] node1234;
	wire [1-1:0] node1235;
	wire [1-1:0] node1237;
	wire [1-1:0] node1241;
	wire [1-1:0] node1242;
	wire [1-1:0] node1246;
	wire [1-1:0] node1248;
	wire [1-1:0] node1249;
	wire [1-1:0] node1250;
	wire [1-1:0] node1251;
	wire [1-1:0] node1257;
	wire [1-1:0] node1258;
	wire [1-1:0] node1259;
	wire [1-1:0] node1260;
	wire [1-1:0] node1261;
	wire [1-1:0] node1263;
	wire [1-1:0] node1266;
	wire [1-1:0] node1268;
	wire [1-1:0] node1269;
	wire [1-1:0] node1270;
	wire [1-1:0] node1275;
	wire [1-1:0] node1276;
	wire [1-1:0] node1277;
	wire [1-1:0] node1282;
	wire [1-1:0] node1283;
	wire [1-1:0] node1285;
	wire [1-1:0] node1286;
	wire [1-1:0] node1292;
	wire [1-1:0] node1293;
	wire [1-1:0] node1294;
	wire [1-1:0] node1295;
	wire [1-1:0] node1296;
	wire [1-1:0] node1298;
	wire [1-1:0] node1301;
	wire [1-1:0] node1302;
	wire [1-1:0] node1303;
	wire [1-1:0] node1308;
	wire [1-1:0] node1309;
	wire [1-1:0] node1310;
	wire [1-1:0] node1311;
	wire [1-1:0] node1313;
	wire [1-1:0] node1314;

	assign outp = (inp[10]) ? node648 : node1;
		assign node1 = (inp[9]) ? node279 : node2;
			assign node2 = (inp[8]) ? node128 : node3;
				assign node3 = (inp[7]) ? node39 : node4;
					assign node4 = (inp[4]) ? node6 : 1'b1;
						assign node6 = (inp[5]) ? node8 : 1'b1;
							assign node8 = (inp[3]) ? node18 : node9;
								assign node9 = (inp[2]) ? node11 : 1'b1;
									assign node11 = (inp[1]) ? node13 : 1'b1;
										assign node13 = (inp[6]) ? node15 : 1'b1;
											assign node15 = (inp[12]) ? 1'b0 : 1'b1;
								assign node18 = (inp[11]) ? node26 : node19;
									assign node19 = (inp[2]) ? node21 : 1'b1;
										assign node21 = (inp[0]) ? node23 : 1'b1;
											assign node23 = (inp[12]) ? 1'b0 : 1'b1;
									assign node26 = (inp[1]) ? node34 : node27;
										assign node27 = (inp[12]) ? node29 : 1'b1;
											assign node29 = (inp[2]) ? node31 : 1'b1;
												assign node31 = (inp[6]) ? 1'b0 : 1'b1;
										assign node34 = (inp[0]) ? 1'b0 : node35;
											assign node35 = (inp[6]) ? 1'b0 : 1'b1;
					assign node39 = (inp[1]) ? node73 : node40;
						assign node40 = (inp[2]) ? node52 : node41;
							assign node41 = (inp[3]) ? node43 : 1'b1;
								assign node43 = (inp[12]) ? node45 : 1'b1;
									assign node45 = (inp[4]) ? node47 : 1'b1;
										assign node47 = (inp[11]) ? node49 : 1'b1;
											assign node49 = (inp[5]) ? 1'b0 : 1'b1;
							assign node52 = (inp[0]) ? node60 : node53;
								assign node53 = (inp[6]) ? node55 : 1'b1;
									assign node55 = (inp[5]) ? node57 : 1'b1;
										assign node57 = (inp[4]) ? 1'b0 : 1'b1;
								assign node60 = (inp[12]) ? node62 : 1'b1;
									assign node62 = (inp[3]) ? node68 : node63;
										assign node63 = (inp[6]) ? node65 : 1'b1;
											assign node65 = (inp[4]) ? 1'b0 : 1'b1;
										assign node68 = (inp[5]) ? 1'b0 : node69;
											assign node69 = (inp[4]) ? 1'b0 : 1'b1;
						assign node73 = (inp[0]) ? node99 : node74;
							assign node74 = (inp[6]) ? node88 : node75;
								assign node75 = (inp[11]) ? node77 : 1'b1;
									assign node77 = (inp[4]) ? node79 : 1'b1;
										assign node79 = (inp[2]) ? node81 : 1'b1;
											assign node81 = (inp[3]) ? 1'b0 : node82;
												assign node82 = (inp[12]) ? node84 : 1'b1;
													assign node84 = (inp[5]) ? 1'b0 : 1'b1;
								assign node88 = (inp[5]) ? node90 : 1'b1;
									assign node90 = (inp[3]) ? 1'b0 : node91;
										assign node91 = (inp[4]) ? node93 : 1'b1;
											assign node93 = (inp[2]) ? 1'b0 : node94;
												assign node94 = (inp[11]) ? 1'b0 : 1'b1;
							assign node99 = (inp[5]) ? node119 : node100;
								assign node100 = (inp[4]) ? node108 : node101;
									assign node101 = (inp[6]) ? node103 : 1'b1;
										assign node103 = (inp[3]) ? node105 : 1'b1;
											assign node105 = (inp[2]) ? 1'b0 : 1'b1;
									assign node108 = (inp[6]) ? node114 : node109;
										assign node109 = (inp[2]) ? node111 : 1'b1;
											assign node111 = (inp[11]) ? 1'b0 : 1'b1;
										assign node114 = (inp[11]) ? 1'b0 : node115;
											assign node115 = (inp[12]) ? 1'b0 : 1'b1;
								assign node119 = (inp[3]) ? 1'b0 : node120;
									assign node120 = (inp[2]) ? node122 : 1'b1;
										assign node122 = (inp[4]) ? 1'b0 : node123;
											assign node123 = (inp[11]) ? 1'b0 : 1'b1;
				assign node128 = (inp[0]) ? node200 : node129;
					assign node129 = (inp[6]) ? node147 : node130;
						assign node130 = (inp[1]) ? node132 : 1'b1;
							assign node132 = (inp[12]) ? node134 : 1'b1;
								assign node134 = (inp[4]) ? node136 : 1'b1;
									assign node136 = (inp[2]) ? node142 : node137;
										assign node137 = (inp[3]) ? node139 : 1'b1;
											assign node139 = (inp[5]) ? 1'b0 : 1'b1;
										assign node142 = (inp[5]) ? 1'b0 : node143;
											assign node143 = (inp[7]) ? 1'b0 : 1'b1;
						assign node147 = (inp[3]) ? node163 : node148;
							assign node148 = (inp[7]) ? node150 : 1'b1;
								assign node150 = (inp[4]) ? node156 : node151;
									assign node151 = (inp[12]) ? node153 : 1'b1;
										assign node153 = (inp[1]) ? 1'b0 : 1'b1;
									assign node156 = (inp[2]) ? node158 : 1'b1;
										assign node158 = (inp[11]) ? 1'b0 : node159;
											assign node159 = (inp[5]) ? 1'b0 : 1'b1;
							assign node163 = (inp[2]) ? node181 : node164;
								assign node164 = (inp[4]) ? node166 : 1'b1;
									assign node166 = (inp[7]) ? node176 : node167;
										assign node167 = (inp[5]) ? node169 : 1'b1;
											assign node169 = (inp[1]) ? 1'b0 : node170;
												assign node170 = (inp[12]) ? node172 : 1'b1;
													assign node172 = (inp[11]) ? 1'b0 : 1'b1;
										assign node176 = (inp[5]) ? 1'b0 : node177;
											assign node177 = (inp[11]) ? 1'b0 : 1'b1;
								assign node181 = (inp[11]) ? node189 : node182;
									assign node182 = (inp[12]) ? node184 : 1'b1;
										assign node184 = (inp[5]) ? 1'b0 : node185;
											assign node185 = (inp[1]) ? 1'b0 : 1'b1;
									assign node189 = (inp[1]) ? 1'b0 : node190;
										assign node190 = (inp[4]) ? 1'b0 : node191;
											assign node191 = (inp[12]) ? node193 : 1'b1;
												assign node193 = (inp[5]) ? 1'b0 : node194;
													assign node194 = (inp[7]) ? 1'b0 : 1'b1;
					assign node200 = (inp[2]) ? node236 : node201;
						assign node201 = (inp[12]) ? node217 : node202;
							assign node202 = (inp[6]) ? node204 : 1'b1;
								assign node204 = (inp[11]) ? node210 : node205;
									assign node205 = (inp[1]) ? node207 : 1'b1;
										assign node207 = (inp[3]) ? 1'b0 : 1'b1;
									assign node210 = (inp[1]) ? 1'b0 : node211;
										assign node211 = (inp[5]) ? node213 : 1'b1;
											assign node213 = (inp[7]) ? 1'b0 : 1'b1;
							assign node217 = (inp[4]) ? node227 : node218;
								assign node218 = (inp[1]) ? node220 : 1'b1;
									assign node220 = (inp[7]) ? 1'b0 : node221;
										assign node221 = (inp[5]) ? node223 : 1'b1;
											assign node223 = (inp[11]) ? 1'b0 : 1'b1;
								assign node227 = (inp[11]) ? 1'b0 : node228;
									assign node228 = (inp[6]) ? node230 : 1'b1;
										assign node230 = (inp[7]) ? 1'b0 : node231;
											assign node231 = (inp[3]) ? 1'b0 : 1'b1;
						assign node236 = (inp[6]) ? node266 : node237;
							assign node237 = (inp[11]) ? node251 : node238;
								assign node238 = (inp[12]) ? node240 : 1'b1;
									assign node240 = (inp[4]) ? node244 : node241;
										assign node241 = (inp[3]) ? 1'b0 : 1'b1;
										assign node244 = (inp[3]) ? node246 : 1'b0;
											assign node246 = (inp[7]) ? 1'b0 : node247;
												assign node247 = (inp[1]) ? 1'b0 : 1'b1;
								assign node251 = (inp[7]) ? node259 : node252;
									assign node252 = (inp[12]) ? node254 : 1'b1;
										assign node254 = (inp[4]) ? 1'b0 : node255;
											assign node255 = (inp[5]) ? 1'b0 : 1'b1;
									assign node259 = (inp[1]) ? 1'b0 : node260;
										assign node260 = (inp[3]) ? 1'b0 : node261;
											assign node261 = (inp[5]) ? 1'b0 : 1'b1;
							assign node266 = (inp[11]) ? 1'b0 : node267;
								assign node267 = (inp[1]) ? 1'b0 : node268;
									assign node268 = (inp[3]) ? node272 : node269;
										assign node269 = (inp[12]) ? 1'b0 : 1'b1;
										assign node272 = (inp[4]) ? 1'b0 : node273;
											assign node273 = (inp[5]) ? 1'b0 : 1'b1;
			assign node279 = (inp[7]) ? node469 : node280;
				assign node280 = (inp[5]) ? node344 : node281;
					assign node281 = (inp[6]) ? node311 : node282;
						assign node282 = (inp[2]) ? node284 : 1'b1;
							assign node284 = (inp[0]) ? node292 : node285;
								assign node285 = (inp[1]) ? node287 : 1'b1;
									assign node287 = (inp[12]) ? node289 : 1'b1;
										assign node289 = (inp[4]) ? 1'b0 : 1'b1;
								assign node292 = (inp[8]) ? node300 : node293;
									assign node293 = (inp[4]) ? node295 : 1'b1;
										assign node295 = (inp[12]) ? node297 : 1'b1;
											assign node297 = (inp[3]) ? 1'b0 : 1'b1;
									assign node300 = (inp[3]) ? node306 : node301;
										assign node301 = (inp[12]) ? node303 : 1'b1;
											assign node303 = (inp[1]) ? 1'b0 : 1'b1;
										assign node306 = (inp[1]) ? 1'b0 : node307;
											assign node307 = (inp[11]) ? 1'b0 : 1'b1;
						assign node311 = (inp[2]) ? node325 : node312;
							assign node312 = (inp[11]) ? node314 : 1'b1;
								assign node314 = (inp[4]) ? node320 : node315;
									assign node315 = (inp[1]) ? node317 : 1'b1;
										assign node317 = (inp[8]) ? 1'b0 : 1'b1;
									assign node320 = (inp[8]) ? 1'b0 : node321;
										assign node321 = (inp[3]) ? 1'b0 : 1'b1;
							assign node325 = (inp[12]) ? node335 : node326;
								assign node326 = (inp[0]) ? node328 : 1'b1;
									assign node328 = (inp[1]) ? node330 : 1'b1;
										assign node330 = (inp[4]) ? 1'b0 : node331;
											assign node331 = (inp[8]) ? 1'b0 : 1'b1;
								assign node335 = (inp[0]) ? 1'b0 : node336;
									assign node336 = (inp[1]) ? node338 : 1'b1;
										assign node338 = (inp[3]) ? 1'b0 : node339;
											assign node339 = (inp[11]) ? 1'b0 : 1'b1;
					assign node344 = (inp[4]) ? node400 : node345;
						assign node345 = (inp[12]) ? node363 : node346;
							assign node346 = (inp[11]) ? node348 : 1'b1;
								assign node348 = (inp[1]) ? node356 : node349;
									assign node349 = (inp[0]) ? node351 : 1'b1;
										assign node351 = (inp[8]) ? node353 : 1'b1;
											assign node353 = (inp[6]) ? 1'b0 : 1'b1;
									assign node356 = (inp[2]) ? 1'b0 : node357;
										assign node357 = (inp[6]) ? node359 : 1'b1;
											assign node359 = (inp[3]) ? 1'b0 : 1'b1;
							assign node363 = (inp[1]) ? node379 : node364;
								assign node364 = (inp[8]) ? node372 : node365;
									assign node365 = (inp[2]) ? node367 : 1'b1;
										assign node367 = (inp[0]) ? node369 : 1'b1;
											assign node369 = (inp[3]) ? 1'b0 : 1'b1;
									assign node372 = (inp[3]) ? 1'b0 : node373;
										assign node373 = (inp[6]) ? node375 : 1'b1;
											assign node375 = (inp[0]) ? 1'b0 : 1'b1;
								assign node379 = (inp[6]) ? node391 : node380;
									assign node380 = (inp[0]) ? node386 : node381;
										assign node381 = (inp[3]) ? node383 : 1'b1;
											assign node383 = (inp[11]) ? 1'b1 : 1'b0;
										assign node386 = (inp[11]) ? 1'b0 : node387;
											assign node387 = (inp[8]) ? 1'b0 : 1'b1;
									assign node391 = (inp[8]) ? 1'b0 : node392;
										assign node392 = (inp[2]) ? 1'b0 : node393;
											assign node393 = (inp[11]) ? 1'b0 : node394;
												assign node394 = (inp[3]) ? 1'b0 : 1'b1;
						assign node400 = (inp[3]) ? node444 : node401;
							assign node401 = (inp[8]) ? node421 : node402;
								assign node402 = (inp[11]) ? node412 : node403;
									assign node403 = (inp[6]) ? node405 : 1'b1;
										assign node405 = (inp[2]) ? node407 : 1'b1;
											assign node407 = (inp[12]) ? node409 : 1'b1;
												assign node409 = (inp[0]) ? 1'b0 : 1'b1;
									assign node412 = (inp[6]) ? 1'b0 : node413;
										assign node413 = (inp[0]) ? node415 : 1'b1;
											assign node415 = (inp[1]) ? 1'b0 : node416;
												assign node416 = (inp[2]) ? 1'b0 : 1'b1;
								assign node421 = (inp[11]) ? node435 : node422;
									assign node422 = (inp[0]) ? node428 : node423;
										assign node423 = (inp[1]) ? node425 : 1'b1;
											assign node425 = (inp[2]) ? 1'b0 : 1'b1;
										assign node428 = (inp[2]) ? 1'b0 : node429;
											assign node429 = (inp[12]) ? node431 : 1'b1;
												assign node431 = (inp[6]) ? 1'b0 : 1'b1;
									assign node435 = (inp[0]) ? 1'b0 : node436;
										assign node436 = (inp[12]) ? 1'b0 : node437;
											assign node437 = (inp[6]) ? 1'b0 : node438;
												assign node438 = (inp[1]) ? 1'b0 : 1'b1;
							assign node444 = (inp[2]) ? node462 : node445;
								assign node445 = (inp[0]) ? 1'b0 : node446;
									assign node446 = (inp[11]) ? node456 : node447;
										assign node447 = (inp[12]) ? node449 : 1'b1;
											assign node449 = (inp[1]) ? node451 : 1'b1;
												assign node451 = (inp[6]) ? 1'b0 : node452;
													assign node452 = (inp[8]) ? 1'b0 : 1'b1;
										assign node456 = (inp[1]) ? 1'b0 : node457;
											assign node457 = (inp[6]) ? 1'b0 : 1'b1;
								assign node462 = (inp[12]) ? 1'b0 : node463;
									assign node463 = (inp[8]) ? 1'b0 : node464;
										assign node464 = (inp[1]) ? 1'b0 : 1'b1;
				assign node469 = (inp[0]) ? node579 : node470;
					assign node470 = (inp[11]) ? node520 : node471;
						assign node471 = (inp[3]) ? node489 : node472;
							assign node472 = (inp[1]) ? node474 : 1'b1;
								assign node474 = (inp[2]) ? node482 : node475;
									assign node475 = (inp[5]) ? node477 : 1'b1;
										assign node477 = (inp[6]) ? node479 : 1'b1;
											assign node479 = (inp[4]) ? 1'b1 : 1'b0;
									assign node482 = (inp[12]) ? 1'b0 : node483;
										assign node483 = (inp[5]) ? node485 : 1'b1;
											assign node485 = (inp[6]) ? 1'b0 : 1'b1;
							assign node489 = (inp[4]) ? node503 : node490;
								assign node490 = (inp[12]) ? node492 : 1'b1;
									assign node492 = (inp[8]) ? node498 : node493;
										assign node493 = (inp[5]) ? node495 : 1'b1;
											assign node495 = (inp[1]) ? 1'b0 : 1'b1;
										assign node498 = (inp[1]) ? 1'b0 : node499;
											assign node499 = (inp[2]) ? 1'b0 : 1'b1;
								assign node503 = (inp[6]) ? node515 : node504;
									assign node504 = (inp[2]) ? node506 : 1'b1;
										assign node506 = (inp[1]) ? node508 : 1'b1;
											assign node508 = (inp[8]) ? 1'b0 : node509;
												assign node509 = (inp[12]) ? 1'b0 : node510;
													assign node510 = (inp[5]) ? 1'b0 : 1'b1;
									assign node515 = (inp[1]) ? 1'b0 : node516;
										assign node516 = (inp[8]) ? 1'b0 : 1'b1;
						assign node520 = (inp[6]) ? node560 : node521;
							assign node521 = (inp[8]) ? node541 : node522;
								assign node522 = (inp[5]) ? node530 : node523;
									assign node523 = (inp[12]) ? node525 : 1'b1;
										assign node525 = (inp[3]) ? node527 : 1'b1;
											assign node527 = (inp[2]) ? 1'b0 : 1'b1;
									assign node530 = (inp[3]) ? node534 : node531;
										assign node531 = (inp[4]) ? 1'b0 : 1'b1;
										assign node534 = (inp[1]) ? 1'b0 : node535;
											assign node535 = (inp[2]) ? node537 : 1'b1;
												assign node537 = (inp[12]) ? 1'b0 : 1'b1;
								assign node541 = (inp[2]) ? 1'b0 : node542;
									assign node542 = (inp[4]) ? node550 : node543;
										assign node543 = (inp[5]) ? node545 : 1'b1;
											assign node545 = (inp[1]) ? 1'b0 : node546;
												assign node546 = (inp[12]) ? 1'b0 : 1'b1;
										assign node550 = (inp[1]) ? 1'b0 : node551;
											assign node551 = (inp[12]) ? 1'b0 : node552;
												assign node552 = (inp[5]) ? node554 : 1'b1;
													assign node554 = (inp[3]) ? 1'b0 : 1'b1;
							assign node560 = (inp[4]) ? 1'b0 : node561;
								assign node561 = (inp[8]) ? node573 : node562;
									assign node562 = (inp[2]) ? node568 : node563;
										assign node563 = (inp[5]) ? node565 : 1'b1;
											assign node565 = (inp[1]) ? 1'b0 : 1'b1;
										assign node568 = (inp[1]) ? 1'b0 : node569;
											assign node569 = (inp[12]) ? 1'b0 : 1'b1;
									assign node573 = (inp[1]) ? 1'b0 : node574;
										assign node574 = (inp[5]) ? 1'b0 : 1'b1;
					assign node579 = (inp[4]) ? node635 : node580;
						assign node580 = (inp[1]) ? node612 : node581;
							assign node581 = (inp[5]) ? node597 : node582;
								assign node582 = (inp[8]) ? node590 : node583;
									assign node583 = (inp[12]) ? node585 : 1'b1;
										assign node585 = (inp[6]) ? node587 : 1'b1;
											assign node587 = (inp[3]) ? 1'b0 : 1'b1;
									assign node590 = (inp[11]) ? 1'b0 : node591;
										assign node591 = (inp[6]) ? node593 : 1'b1;
											assign node593 = (inp[12]) ? 1'b0 : 1'b1;
								assign node597 = (inp[11]) ? node607 : node598;
									assign node598 = (inp[2]) ? node602 : node599;
										assign node599 = (inp[8]) ? 1'b0 : 1'b1;
										assign node602 = (inp[6]) ? 1'b0 : node603;
											assign node603 = (inp[3]) ? 1'b0 : 1'b1;
									assign node607 = (inp[12]) ? 1'b0 : node608;
										assign node608 = (inp[6]) ? 1'b0 : 1'b1;
							assign node612 = (inp[3]) ? node626 : node613;
								assign node613 = (inp[2]) ? node619 : node614;
									assign node614 = (inp[11]) ? node616 : 1'b1;
										assign node616 = (inp[8]) ? 1'b0 : 1'b1;
									assign node619 = (inp[12]) ? 1'b0 : node620;
										assign node620 = (inp[11]) ? 1'b0 : node621;
											assign node621 = (inp[5]) ? 1'b0 : 1'b1;
								assign node626 = (inp[6]) ? 1'b0 : node627;
									assign node627 = (inp[2]) ? 1'b0 : node628;
										assign node628 = (inp[8]) ? 1'b0 : node629;
											assign node629 = (inp[5]) ? 1'b0 : 1'b1;
						assign node635 = (inp[8]) ? 1'b0 : node636;
							assign node636 = (inp[12]) ? 1'b0 : node637;
								assign node637 = (inp[2]) ? 1'b0 : node638;
									assign node638 = (inp[1]) ? 1'b0 : node639;
										assign node639 = (inp[3]) ? node641 : 1'b1;
											assign node641 = (inp[6]) ? 1'b0 : 1'b1;
		assign node648 = (inp[2]) ? node1012 : node649;
			assign node649 = (inp[4]) ? node847 : node650;
				assign node650 = (inp[1]) ? node732 : node651;
					assign node651 = (inp[3]) ? node671 : node652;
						assign node652 = (inp[5]) ? node654 : 1'b1;
							assign node654 = (inp[8]) ? node656 : 1'b1;
								assign node656 = (inp[9]) ? node662 : node657;
									assign node657 = (inp[11]) ? node659 : 1'b1;
										assign node659 = (inp[6]) ? 1'b0 : 1'b1;
									assign node662 = (inp[6]) ? 1'b0 : node663;
										assign node663 = (inp[0]) ? node665 : 1'b1;
											assign node665 = (inp[12]) ? 1'b0 : node666;
												assign node666 = (inp[7]) ? 1'b0 : 1'b1;
						assign node671 = (inp[0]) ? node699 : node672;
							assign node672 = (inp[12]) ? node680 : node673;
								assign node673 = (inp[9]) ? node675 : 1'b1;
									assign node675 = (inp[7]) ? node677 : 1'b1;
										assign node677 = (inp[5]) ? 1'b0 : 1'b1;
								assign node680 = (inp[7]) ? node690 : node681;
									assign node681 = (inp[8]) ? node683 : 1'b1;
										assign node683 = (inp[9]) ? node685 : 1'b1;
											assign node685 = (inp[5]) ? 1'b0 : node686;
												assign node686 = (inp[6]) ? 1'b0 : 1'b1;
									assign node690 = (inp[5]) ? node694 : node691;
										assign node691 = (inp[11]) ? 1'b0 : 1'b1;
										assign node694 = (inp[6]) ? 1'b0 : node695;
											assign node695 = (inp[9]) ? 1'b0 : 1'b1;
							assign node699 = (inp[5]) ? node715 : node700;
								assign node700 = (inp[6]) ? node708 : node701;
									assign node701 = (inp[11]) ? node703 : 1'b1;
										assign node703 = (inp[8]) ? node705 : 1'b1;
											assign node705 = (inp[12]) ? 1'b0 : 1'b1;
									assign node708 = (inp[9]) ? 1'b0 : node709;
										assign node709 = (inp[8]) ? node711 : 1'b1;
											assign node711 = (inp[12]) ? 1'b0 : 1'b1;
								assign node715 = (inp[9]) ? 1'b0 : node716;
									assign node716 = (inp[6]) ? node726 : node717;
										assign node717 = (inp[12]) ? node719 : 1'b1;
											assign node719 = (inp[8]) ? node721 : 1'b1;
												assign node721 = (inp[11]) ? 1'b0 : node722;
													assign node722 = (inp[7]) ? 1'b0 : 1'b1;
										assign node726 = (inp[8]) ? 1'b0 : node727;
											assign node727 = (inp[12]) ? 1'b0 : 1'b1;
					assign node732 = (inp[5]) ? node788 : node733;
						assign node733 = (inp[6]) ? node759 : node734;
							assign node734 = (inp[11]) ? node744 : node735;
								assign node735 = (inp[7]) ? node737 : 1'b1;
									assign node737 = (inp[0]) ? node739 : 1'b1;
										assign node739 = (inp[9]) ? node741 : 1'b1;
											assign node741 = (inp[3]) ? 1'b0 : 1'b1;
								assign node744 = (inp[9]) ? node752 : node745;
									assign node745 = (inp[7]) ? node747 : 1'b1;
										assign node747 = (inp[0]) ? node749 : 1'b1;
											assign node749 = (inp[12]) ? 1'b0 : 1'b1;
									assign node752 = (inp[3]) ? 1'b0 : node753;
										assign node753 = (inp[8]) ? 1'b1 : node754;
											assign node754 = (inp[12]) ? 1'b0 : 1'b1;
							assign node759 = (inp[8]) ? node775 : node760;
								assign node760 = (inp[12]) ? node768 : node761;
									assign node761 = (inp[3]) ? node763 : 1'b1;
										assign node763 = (inp[9]) ? node765 : 1'b1;
											assign node765 = (inp[11]) ? 1'b0 : 1'b1;
									assign node768 = (inp[0]) ? 1'b0 : node769;
										assign node769 = (inp[7]) ? node771 : 1'b1;
											assign node771 = (inp[3]) ? 1'b0 : 1'b1;
								assign node775 = (inp[3]) ? 1'b0 : node776;
									assign node776 = (inp[11]) ? node782 : node777;
										assign node777 = (inp[0]) ? node779 : 1'b1;
											assign node779 = (inp[12]) ? 1'b0 : 1'b1;
										assign node782 = (inp[9]) ? 1'b0 : node783;
											assign node783 = (inp[0]) ? 1'b0 : 1'b1;
						assign node788 = (inp[12]) ? node822 : node789;
							assign node789 = (inp[0]) ? node807 : node790;
								assign node790 = (inp[11]) ? node792 : 1'b1;
									assign node792 = (inp[9]) ? node798 : node793;
										assign node793 = (inp[7]) ? node795 : 1'b1;
											assign node795 = (inp[6]) ? 1'b0 : 1'b1;
										assign node798 = (inp[3]) ? 1'b0 : node799;
											assign node799 = (inp[8]) ? 1'b0 : node800;
												assign node800 = (inp[7]) ? node802 : 1'b1;
													assign node802 = (inp[6]) ? 1'b0 : 1'b1;
								assign node807 = (inp[3]) ? node815 : node808;
									assign node808 = (inp[9]) ? node810 : 1'b1;
										assign node810 = (inp[8]) ? 1'b0 : node811;
											assign node811 = (inp[7]) ? 1'b0 : 1'b1;
									assign node815 = (inp[11]) ? 1'b0 : node816;
										assign node816 = (inp[7]) ? 1'b0 : node817;
											assign node817 = (inp[6]) ? 1'b1 : 1'b0;
							assign node822 = (inp[9]) ? node840 : node823;
								assign node823 = (inp[7]) ? node833 : node824;
									assign node824 = (inp[8]) ? node826 : 1'b1;
										assign node826 = (inp[11]) ? 1'b0 : node827;
											assign node827 = (inp[3]) ? node829 : 1'b1;
												assign node829 = (inp[6]) ? 1'b0 : 1'b1;
									assign node833 = (inp[3]) ? 1'b0 : node834;
										assign node834 = (inp[8]) ? 1'b0 : node835;
											assign node835 = (inp[6]) ? 1'b0 : 1'b1;
								assign node840 = (inp[8]) ? 1'b0 : node841;
									assign node841 = (inp[7]) ? 1'b0 : node842;
										assign node842 = (inp[11]) ? 1'b0 : 1'b1;
				assign node847 = (inp[8]) ? node943 : node848;
					assign node848 = (inp[12]) ? node900 : node849;
						assign node849 = (inp[7]) ? node863 : node850;
							assign node850 = (inp[11]) ? node852 : 1'b1;
								assign node852 = (inp[6]) ? node858 : node853;
									assign node853 = (inp[3]) ? node855 : 1'b1;
										assign node855 = (inp[5]) ? 1'b0 : 1'b1;
									assign node858 = (inp[0]) ? 1'b0 : node859;
										assign node859 = (inp[3]) ? 1'b0 : 1'b1;
							assign node863 = (inp[9]) ? node877 : node864;
								assign node864 = (inp[0]) ? node870 : node865;
									assign node865 = (inp[5]) ? node867 : 1'b1;
										assign node867 = (inp[6]) ? 1'b0 : 1'b1;
									assign node870 = (inp[3]) ? node872 : 1'b1;
										assign node872 = (inp[1]) ? 1'b0 : node873;
											assign node873 = (inp[5]) ? 1'b0 : 1'b1;
								assign node877 = (inp[5]) ? node893 : node878;
									assign node878 = (inp[3]) ? node888 : node879;
										assign node879 = (inp[6]) ? node881 : 1'b1;
											assign node881 = (inp[0]) ? 1'b0 : node882;
												assign node882 = (inp[1]) ? node884 : 1'b1;
													assign node884 = (inp[11]) ? 1'b0 : 1'b1;
										assign node888 = (inp[11]) ? 1'b0 : node889;
											assign node889 = (inp[0]) ? 1'b0 : 1'b1;
									assign node893 = (inp[11]) ? 1'b0 : node894;
										assign node894 = (inp[3]) ? node896 : 1'b0;
											assign node896 = (inp[6]) ? 1'b0 : 1'b1;
						assign node900 = (inp[11]) ? node928 : node901;
							assign node901 = (inp[1]) ? node911 : node902;
								assign node902 = (inp[7]) ? node904 : 1'b1;
									assign node904 = (inp[3]) ? node906 : 1'b1;
										assign node906 = (inp[0]) ? 1'b0 : node907;
											assign node907 = (inp[5]) ? 1'b0 : 1'b1;
								assign node911 = (inp[3]) ? node921 : node912;
									assign node912 = (inp[5]) ? node918 : node913;
										assign node913 = (inp[7]) ? node915 : 1'b1;
											assign node915 = (inp[6]) ? 1'b0 : 1'b1;
										assign node918 = (inp[0]) ? 1'b0 : 1'b1;
									assign node921 = (inp[9]) ? 1'b0 : node922;
										assign node922 = (inp[0]) ? 1'b0 : node923;
											assign node923 = (inp[7]) ? 1'b0 : 1'b1;
							assign node928 = (inp[1]) ? 1'b0 : node929;
								assign node929 = (inp[0]) ? 1'b0 : node930;
									assign node930 = (inp[9]) ? node936 : node931;
										assign node931 = (inp[5]) ? node933 : 1'b1;
											assign node933 = (inp[6]) ? 1'b0 : 1'b1;
										assign node936 = (inp[5]) ? 1'b0 : node937;
											assign node937 = (inp[6]) ? 1'b0 : 1'b1;
					assign node943 = (inp[12]) ? node993 : node944;
						assign node944 = (inp[3]) ? node966 : node945;
							assign node945 = (inp[6]) ? node955 : node946;
								assign node946 = (inp[9]) ? node948 : 1'b1;
									assign node948 = (inp[5]) ? node950 : 1'b1;
										assign node950 = (inp[7]) ? 1'b0 : node951;
											assign node951 = (inp[0]) ? 1'b0 : 1'b1;
								assign node955 = (inp[5]) ? node961 : node956;
									assign node956 = (inp[11]) ? 1'b0 : node957;
										assign node957 = (inp[0]) ? 1'b0 : 1'b1;
									assign node961 = (inp[7]) ? 1'b0 : node962;
										assign node962 = (inp[1]) ? 1'b0 : 1'b1;
							assign node966 = (inp[1]) ? node986 : node967;
								assign node967 = (inp[9]) ? node979 : node968;
									assign node968 = (inp[11]) ? node974 : node969;
										assign node969 = (inp[0]) ? node971 : 1'b1;
											assign node971 = (inp[5]) ? 1'b0 : 1'b1;
										assign node974 = (inp[7]) ? 1'b0 : node975;
											assign node975 = (inp[6]) ? 1'b0 : 1'b1;
									assign node979 = (inp[0]) ? 1'b0 : node980;
										assign node980 = (inp[11]) ? 1'b0 : node981;
											assign node981 = (inp[6]) ? 1'b0 : 1'b1;
								assign node986 = (inp[11]) ? 1'b0 : node987;
									assign node987 = (inp[7]) ? 1'b0 : node988;
										assign node988 = (inp[5]) ? 1'b0 : 1'b1;
						assign node993 = (inp[6]) ? 1'b0 : node994;
							assign node994 = (inp[0]) ? 1'b0 : node995;
								assign node995 = (inp[11]) ? node1003 : node996;
									assign node996 = (inp[1]) ? node998 : 1'b1;
										assign node998 = (inp[9]) ? 1'b0 : node999;
											assign node999 = (inp[3]) ? 1'b0 : 1'b1;
									assign node1003 = (inp[7]) ? 1'b0 : node1004;
										assign node1004 = (inp[9]) ? 1'b0 : node1005;
											assign node1005 = (inp[5]) ? 1'b1 : 1'b0;
			assign node1012 = (inp[3]) ? node1198 : node1013;
				assign node1013 = (inp[4]) ? node1119 : node1014;
					assign node1014 = (inp[7]) ? node1060 : node1015;
						assign node1015 = (inp[6]) ? node1041 : node1016;
							assign node1016 = (inp[12]) ? node1028 : node1017;
								assign node1017 = (inp[1]) ? 1'b1 : node1018;
									assign node1018 = (inp[5]) ? node1020 : 1'b1;
										assign node1020 = (inp[9]) ? node1022 : 1'b1;
											assign node1022 = (inp[8]) ? node1024 : 1'b1;
												assign node1024 = (inp[0]) ? 1'b0 : 1'b1;
								assign node1028 = (inp[8]) ? node1036 : node1029;
									assign node1029 = (inp[9]) ? node1031 : 1'b1;
										assign node1031 = (inp[11]) ? node1033 : 1'b1;
											assign node1033 = (inp[5]) ? 1'b0 : 1'b1;
									assign node1036 = (inp[0]) ? 1'b0 : node1037;
										assign node1037 = (inp[1]) ? 1'b0 : 1'b1;
							assign node1041 = (inp[1]) ? node1051 : node1042;
								assign node1042 = (inp[9]) ? node1044 : 1'b1;
									assign node1044 = (inp[8]) ? 1'b0 : node1045;
										assign node1045 = (inp[5]) ? node1047 : 1'b1;
											assign node1047 = (inp[0]) ? 1'b0 : 1'b1;
								assign node1051 = (inp[0]) ? 1'b0 : node1052;
									assign node1052 = (inp[8]) ? node1054 : 1'b1;
										assign node1054 = (inp[5]) ? 1'b0 : node1055;
											assign node1055 = (inp[12]) ? 1'b0 : 1'b1;
						assign node1060 = (inp[12]) ? node1094 : node1061;
							assign node1061 = (inp[6]) ? node1081 : node1062;
								assign node1062 = (inp[0]) ? node1070 : node1063;
									assign node1063 = (inp[9]) ? node1065 : 1'b1;
										assign node1065 = (inp[11]) ? node1067 : 1'b1;
											assign node1067 = (inp[5]) ? 1'b0 : 1'b1;
									assign node1070 = (inp[11]) ? node1076 : node1071;
										assign node1071 = (inp[9]) ? node1073 : 1'b1;
											assign node1073 = (inp[8]) ? 1'b0 : 1'b1;
										assign node1076 = (inp[1]) ? 1'b0 : node1077;
											assign node1077 = (inp[5]) ? 1'b0 : 1'b1;
								assign node1081 = (inp[8]) ? 1'b0 : node1082;
									assign node1082 = (inp[0]) ? node1088 : node1083;
										assign node1083 = (inp[5]) ? node1085 : 1'b1;
											assign node1085 = (inp[11]) ? 1'b0 : 1'b1;
										assign node1088 = (inp[11]) ? 1'b0 : node1089;
											assign node1089 = (inp[1]) ? 1'b0 : 1'b1;
							assign node1094 = (inp[5]) ? node1110 : node1095;
								assign node1095 = (inp[11]) ? 1'b0 : node1096;
									assign node1096 = (inp[0]) ? node1102 : node1097;
										assign node1097 = (inp[1]) ? node1099 : 1'b1;
											assign node1099 = (inp[9]) ? 1'b0 : 1'b1;
										assign node1102 = (inp[9]) ? 1'b0 : node1103;
											assign node1103 = (inp[1]) ? 1'b0 : node1104;
												assign node1104 = (inp[8]) ? 1'b0 : 1'b1;
								assign node1110 = (inp[8]) ? 1'b0 : node1111;
									assign node1111 = (inp[6]) ? 1'b0 : node1112;
										assign node1112 = (inp[0]) ? 1'b0 : node1113;
											assign node1113 = (inp[9]) ? 1'b0 : 1'b1;
					assign node1119 = (inp[0]) ? node1161 : node1120;
						assign node1120 = (inp[5]) ? node1144 : node1121;
							assign node1121 = (inp[11]) ? node1129 : node1122;
								assign node1122 = (inp[9]) ? node1124 : 1'b1;
									assign node1124 = (inp[7]) ? node1126 : 1'b1;
										assign node1126 = (inp[8]) ? 1'b0 : 1'b1;
								assign node1129 = (inp[8]) ? node1139 : node1130;
									assign node1130 = (inp[6]) ? node1132 : 1'b1;
										assign node1132 = (inp[7]) ? 1'b0 : node1133;
											assign node1133 = (inp[1]) ? node1135 : 1'b1;
												assign node1135 = (inp[9]) ? 1'b0 : 1'b1;
									assign node1139 = (inp[1]) ? 1'b0 : node1140;
										assign node1140 = (inp[12]) ? 1'b0 : 1'b1;
							assign node1144 = (inp[8]) ? node1154 : node1145;
								assign node1145 = (inp[7]) ? 1'b0 : node1146;
									assign node1146 = (inp[12]) ? node1148 : 1'b1;
										assign node1148 = (inp[1]) ? 1'b0 : node1149;
											assign node1149 = (inp[6]) ? 1'b0 : 1'b1;
								assign node1154 = (inp[12]) ? 1'b0 : node1155;
									assign node1155 = (inp[1]) ? 1'b0 : node1156;
										assign node1156 = (inp[11]) ? 1'b0 : 1'b1;
						assign node1161 = (inp[9]) ? node1189 : node1162;
							assign node1162 = (inp[8]) ? node1182 : node1163;
								assign node1163 = (inp[5]) ? node1175 : node1164;
									assign node1164 = (inp[6]) ? node1170 : node1165;
										assign node1165 = (inp[11]) ? node1167 : 1'b1;
											assign node1167 = (inp[1]) ? 1'b0 : 1'b1;
										assign node1170 = (inp[1]) ? 1'b0 : node1171;
											assign node1171 = (inp[11]) ? 1'b0 : 1'b1;
									assign node1175 = (inp[12]) ? 1'b0 : node1176;
										assign node1176 = (inp[1]) ? 1'b0 : node1177;
											assign node1177 = (inp[7]) ? 1'b0 : 1'b1;
								assign node1182 = (inp[12]) ? 1'b0 : node1183;
									assign node1183 = (inp[7]) ? 1'b0 : node1184;
										assign node1184 = (inp[11]) ? 1'b0 : 1'b1;
							assign node1189 = (inp[12]) ? 1'b0 : node1190;
								assign node1190 = (inp[11]) ? 1'b0 : node1191;
									assign node1191 = (inp[1]) ? 1'b0 : node1192;
										assign node1192 = (inp[7]) ? 1'b0 : 1'b1;
				assign node1198 = (inp[11]) ? node1292 : node1199;
					assign node1199 = (inp[12]) ? node1257 : node1200;
						assign node1200 = (inp[6]) ? node1226 : node1201;
							assign node1201 = (inp[4]) ? node1217 : node1202;
								assign node1202 = (inp[8]) ? node1208 : node1203;
									assign node1203 = (inp[0]) ? node1205 : 1'b1;
										assign node1205 = (inp[1]) ? 1'b0 : 1'b1;
									assign node1208 = (inp[9]) ? 1'b0 : node1209;
										assign node1209 = (inp[1]) ? node1211 : 1'b1;
											assign node1211 = (inp[5]) ? 1'b0 : node1212;
												assign node1212 = (inp[7]) ? 1'b0 : 1'b1;
								assign node1217 = (inp[5]) ? 1'b0 : node1218;
									assign node1218 = (inp[1]) ? 1'b0 : node1219;
										assign node1219 = (inp[9]) ? node1221 : 1'b1;
											assign node1221 = (inp[0]) ? 1'b0 : 1'b1;
							assign node1226 = (inp[8]) ? node1246 : node1227;
								assign node1227 = (inp[7]) ? node1241 : node1228;
									assign node1228 = (inp[1]) ? node1234 : node1229;
										assign node1229 = (inp[4]) ? node1231 : 1'b1;
											assign node1231 = (inp[9]) ? 1'b0 : 1'b1;
										assign node1234 = (inp[9]) ? 1'b0 : node1235;
											assign node1235 = (inp[0]) ? node1237 : 1'b1;
												assign node1237 = (inp[5]) ? 1'b0 : 1'b1;
									assign node1241 = (inp[9]) ? 1'b0 : node1242;
										assign node1242 = (inp[1]) ? 1'b0 : 1'b1;
								assign node1246 = (inp[4]) ? node1248 : 1'b0;
									assign node1248 = (inp[1]) ? 1'b0 : node1249;
										assign node1249 = (inp[0]) ? 1'b0 : node1250;
											assign node1250 = (inp[9]) ? 1'b0 : node1251;
												assign node1251 = (inp[7]) ? 1'b0 : 1'b1;
						assign node1257 = (inp[5]) ? 1'b0 : node1258;
							assign node1258 = (inp[8]) ? node1282 : node1259;
								assign node1259 = (inp[6]) ? node1275 : node1260;
									assign node1260 = (inp[4]) ? node1266 : node1261;
										assign node1261 = (inp[0]) ? node1263 : 1'b1;
											assign node1263 = (inp[7]) ? 1'b0 : 1'b1;
										assign node1266 = (inp[1]) ? node1268 : 1'b1;
											assign node1268 = (inp[0]) ? 1'b0 : node1269;
												assign node1269 = (inp[9]) ? 1'b0 : node1270;
													assign node1270 = (inp[7]) ? 1'b0 : 1'b1;
									assign node1275 = (inp[1]) ? 1'b0 : node1276;
										assign node1276 = (inp[0]) ? 1'b0 : node1277;
											assign node1277 = (inp[9]) ? 1'b0 : 1'b1;
								assign node1282 = (inp[7]) ? 1'b0 : node1283;
									assign node1283 = (inp[0]) ? node1285 : 1'b0;
										assign node1285 = (inp[9]) ? 1'b0 : node1286;
											assign node1286 = (inp[1]) ? 1'b0 : 1'b1;
					assign node1292 = (inp[1]) ? 1'b0 : node1293;
						assign node1293 = (inp[4]) ? 1'b0 : node1294;
							assign node1294 = (inp[9]) ? node1308 : node1295;
								assign node1295 = (inp[8]) ? node1301 : node1296;
									assign node1296 = (inp[5]) ? node1298 : 1'b1;
										assign node1298 = (inp[7]) ? 1'b1 : 1'b0;
									assign node1301 = (inp[6]) ? 1'b0 : node1302;
										assign node1302 = (inp[7]) ? 1'b0 : node1303;
											assign node1303 = (inp[0]) ? 1'b0 : 1'b1;
								assign node1308 = (inp[5]) ? 1'b0 : node1309;
									assign node1309 = (inp[12]) ? 1'b0 : node1310;
										assign node1310 = (inp[6]) ? 1'b0 : node1311;
											assign node1311 = (inp[0]) ? node1313 : 1'b1;
												assign node1313 = (inp[8]) ? 1'b0 : node1314;
													assign node1314 = (inp[7]) ? 1'b0 : 1'b1;

endmodule