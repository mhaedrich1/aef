module dtc_split875_bm60 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node6;
	wire [3-1:0] node8;
	wire [3-1:0] node10;
	wire [3-1:0] node12;
	wire [3-1:0] node14;
	wire [3-1:0] node17;
	wire [3-1:0] node18;
	wire [3-1:0] node20;
	wire [3-1:0] node22;
	wire [3-1:0] node26;
	wire [3-1:0] node27;
	wire [3-1:0] node29;
	wire [3-1:0] node31;
	wire [3-1:0] node33;
	wire [3-1:0] node36;
	wire [3-1:0] node37;
	wire [3-1:0] node38;
	wire [3-1:0] node39;
	wire [3-1:0] node41;
	wire [3-1:0] node43;
	wire [3-1:0] node48;
	wire [3-1:0] node51;
	wire [3-1:0] node52;
	wire [3-1:0] node53;
	wire [3-1:0] node55;
	wire [3-1:0] node57;
	wire [3-1:0] node58;
	wire [3-1:0] node60;
	wire [3-1:0] node62;
	wire [3-1:0] node66;
	wire [3-1:0] node68;
	wire [3-1:0] node71;
	wire [3-1:0] node72;
	wire [3-1:0] node74;
	wire [3-1:0] node75;
	wire [3-1:0] node77;
	wire [3-1:0] node79;
	wire [3-1:0] node81;
	wire [3-1:0] node84;
	wire [3-1:0] node86;
	wire [3-1:0] node88;
	wire [3-1:0] node90;
	wire [3-1:0] node93;
	wire [3-1:0] node94;
	wire [3-1:0] node96;
	wire [3-1:0] node98;
	wire [3-1:0] node102;
	wire [3-1:0] node103;
	wire [3-1:0] node104;
	wire [3-1:0] node105;
	wire [3-1:0] node107;
	wire [3-1:0] node108;
	wire [3-1:0] node110;
	wire [3-1:0] node112;
	wire [3-1:0] node114;
	wire [3-1:0] node118;
	wire [3-1:0] node119;
	wire [3-1:0] node120;
	wire [3-1:0] node121;
	wire [3-1:0] node123;
	wire [3-1:0] node125;
	wire [3-1:0] node131;
	wire [3-1:0] node132;
	wire [3-1:0] node133;
	wire [3-1:0] node135;
	wire [3-1:0] node137;
	wire [3-1:0] node141;
	wire [3-1:0] node143;
	wire [3-1:0] node144;
	wire [3-1:0] node146;
	wire [3-1:0] node148;
	wire [3-1:0] node150;
	wire [3-1:0] node154;
	wire [3-1:0] node155;
	wire [3-1:0] node156;
	wire [3-1:0] node158;
	wire [3-1:0] node159;
	wire [3-1:0] node161;
	wire [3-1:0] node163;
	wire [3-1:0] node165;
	wire [3-1:0] node168;
	wire [3-1:0] node169;
	wire [3-1:0] node171;
	wire [3-1:0] node173;
	wire [3-1:0] node177;
	wire [3-1:0] node179;
	wire [3-1:0] node180;
	wire [3-1:0] node182;
	wire [3-1:0] node186;
	wire [3-1:0] node187;
	wire [3-1:0] node188;
	wire [3-1:0] node189;
	wire [3-1:0] node190;
	wire [3-1:0] node192;
	wire [3-1:0] node194;
	wire [3-1:0] node198;
	wire [3-1:0] node200;
	wire [3-1:0] node202;
	wire [3-1:0] node204;
	wire [3-1:0] node207;
	wire [3-1:0] node209;
	wire [3-1:0] node210;
	wire [3-1:0] node214;
	wire [3-1:0] node215;
	wire [3-1:0] node216;
	wire [3-1:0] node218;
	wire [3-1:0] node220;
	wire [3-1:0] node222;
	wire [3-1:0] node225;
	wire [3-1:0] node226;
	wire [3-1:0] node228;
	wire [3-1:0] node230;
	wire [3-1:0] node234;
	wire [3-1:0] node235;
	wire [3-1:0] node237;
	wire [3-1:0] node240;
	wire [3-1:0] node241;
	wire [3-1:0] node243;
	wire [3-1:0] node245;
	wire [3-1:0] node248;
	wire [3-1:0] node250;
	wire [3-1:0] node252;

	assign outp = (inp[2]) ? node102 : node1;
		assign node1 = (inp[3]) ? node51 : node2;
			assign node2 = (inp[10]) ? node26 : node3;
				assign node3 = (inp[4]) ? node17 : node4;
					assign node4 = (inp[11]) ? node6 : 3'b111;
						assign node6 = (inp[5]) ? node8 : 3'b111;
							assign node8 = (inp[7]) ? node10 : 3'b111;
								assign node10 = (inp[6]) ? node12 : 3'b111;
									assign node12 = (inp[9]) ? node14 : 3'b111;
										assign node14 = (inp[8]) ? 3'b110 : 3'b111;
					assign node17 = (inp[5]) ? 3'b111 : node18;
						assign node18 = (inp[7]) ? node20 : 3'b110;
							assign node20 = (inp[9]) ? node22 : 3'b110;
								assign node22 = (inp[8]) ? 3'b111 : 3'b110;
				assign node26 = (inp[4]) ? node36 : node27;
					assign node27 = (inp[7]) ? node29 : 3'b110;
						assign node29 = (inp[8]) ? node31 : 3'b110;
							assign node31 = (inp[5]) ? node33 : 3'b110;
								assign node33 = (inp[9]) ? 3'b111 : 3'b110;
					assign node36 = (inp[9]) ? node48 : node37;
						assign node37 = (inp[5]) ? 3'b110 : node38;
							assign node38 = (inp[7]) ? 3'b110 : node39;
								assign node39 = (inp[8]) ? node41 : 3'b111;
									assign node41 = (inp[6]) ? node43 : 3'b111;
										assign node43 = (inp[11]) ? 3'b110 : 3'b111;
						assign node48 = (inp[5]) ? 3'b011 : 3'b110;
			assign node51 = (inp[4]) ? node71 : node52;
				assign node52 = (inp[10]) ? node66 : node53;
					assign node53 = (inp[9]) ? node55 : 3'b111;
						assign node55 = (inp[5]) ? node57 : 3'b111;
							assign node57 = (inp[7]) ? 3'b110 : node58;
								assign node58 = (inp[6]) ? node60 : 3'b111;
									assign node60 = (inp[8]) ? node62 : 3'b111;
										assign node62 = (inp[11]) ? 3'b110 : 3'b111;
					assign node66 = (inp[5]) ? node68 : 3'b110;
						assign node68 = (inp[9]) ? 3'b011 : 3'b110;
				assign node71 = (inp[5]) ? node93 : node72;
					assign node72 = (inp[9]) ? node74 : 3'b011;
						assign node74 = (inp[7]) ? node84 : node75;
							assign node75 = (inp[8]) ? node77 : 3'b011;
								assign node77 = (inp[6]) ? node79 : 3'b011;
									assign node79 = (inp[11]) ? node81 : 3'b011;
										assign node81 = (inp[10]) ? 3'b011 : 3'b010;
							assign node84 = (inp[10]) ? node86 : 3'b010;
								assign node86 = (inp[11]) ? node88 : 3'b011;
									assign node88 = (inp[6]) ? node90 : 3'b011;
										assign node90 = (inp[8]) ? 3'b010 : 3'b011;
					assign node93 = (inp[10]) ? 3'b010 : node94;
						assign node94 = (inp[9]) ? node96 : 3'b010;
							assign node96 = (inp[7]) ? node98 : 3'b010;
								assign node98 = (inp[8]) ? 3'b011 : 3'b010;
		assign node102 = (inp[4]) ? node154 : node103;
			assign node103 = (inp[10]) ? node131 : node104;
				assign node104 = (inp[5]) ? node118 : node105;
					assign node105 = (inp[3]) ? node107 : 3'b011;
						assign node107 = (inp[9]) ? 3'b010 : node108;
							assign node108 = (inp[7]) ? node110 : 3'b011;
								assign node110 = (inp[6]) ? node112 : 3'b011;
									assign node112 = (inp[8]) ? node114 : 3'b011;
										assign node114 = (inp[11]) ? 3'b010 : 3'b011;
					assign node118 = (inp[7]) ? 3'b010 : node119;
						assign node119 = (inp[3]) ? 3'b010 : node120;
							assign node120 = (inp[9]) ? 3'b010 : node121;
								assign node121 = (inp[6]) ? node123 : 3'b011;
									assign node123 = (inp[11]) ? node125 : 3'b011;
										assign node125 = (inp[8]) ? 3'b010 : 3'b011;
				assign node131 = (inp[3]) ? node141 : node132;
					assign node132 = (inp[5]) ? 3'b011 : node133;
						assign node133 = (inp[8]) ? node135 : 3'b010;
							assign node135 = (inp[9]) ? node137 : 3'b010;
								assign node137 = (inp[7]) ? 3'b011 : 3'b010;
					assign node141 = (inp[5]) ? node143 : 3'b111;
						assign node143 = (inp[9]) ? 3'b110 : node144;
							assign node144 = (inp[8]) ? node146 : 3'b111;
								assign node146 = (inp[7]) ? node148 : 3'b111;
									assign node148 = (inp[11]) ? node150 : 3'b111;
										assign node150 = (inp[6]) ? 3'b110 : 3'b111;
			assign node154 = (inp[3]) ? node186 : node155;
				assign node155 = (inp[5]) ? node177 : node156;
					assign node156 = (inp[9]) ? node158 : 3'b101;
						assign node158 = (inp[10]) ? node168 : node159;
							assign node159 = (inp[6]) ? node161 : 3'b101;
								assign node161 = (inp[11]) ? node163 : 3'b101;
									assign node163 = (inp[8]) ? node165 : 3'b101;
										assign node165 = (inp[7]) ? 3'b100 : 3'b101;
							assign node168 = (inp[7]) ? 3'b100 : node169;
								assign node169 = (inp[8]) ? node171 : 3'b101;
									assign node171 = (inp[11]) ? node173 : 3'b101;
										assign node173 = (inp[6]) ? 3'b100 : 3'b101;
					assign node177 = (inp[9]) ? node179 : 3'b100;
						assign node179 = (inp[10]) ? 3'b001 : node180;
							assign node180 = (inp[8]) ? node182 : 3'b100;
								assign node182 = (inp[7]) ? 3'b101 : 3'b100;
				assign node186 = (inp[10]) ? node214 : node187;
					assign node187 = (inp[9]) ? node207 : node188;
						assign node188 = (inp[5]) ? node198 : node189;
							assign node189 = (inp[7]) ? 3'b000 : node190;
								assign node190 = (inp[8]) ? node192 : 3'b001;
									assign node192 = (inp[11]) ? node194 : 3'b001;
										assign node194 = (inp[6]) ? 3'b000 : 3'b001;
							assign node198 = (inp[6]) ? node200 : 3'b001;
								assign node200 = (inp[7]) ? node202 : 3'b001;
									assign node202 = (inp[11]) ? node204 : 3'b001;
										assign node204 = (inp[8]) ? 3'b000 : 3'b001;
						assign node207 = (inp[7]) ? node209 : 3'b000;
							assign node209 = (inp[5]) ? 3'b000 : node210;
								assign node210 = (inp[8]) ? 3'b001 : 3'b000;
					assign node214 = (inp[9]) ? node234 : node215;
						assign node215 = (inp[7]) ? node225 : node216;
							assign node216 = (inp[6]) ? node218 : 3'b101;
								assign node218 = (inp[5]) ? node220 : 3'b101;
									assign node220 = (inp[11]) ? node222 : 3'b101;
										assign node222 = (inp[8]) ? 3'b100 : 3'b101;
							assign node225 = (inp[5]) ? 3'b100 : node226;
								assign node226 = (inp[11]) ? node228 : 3'b101;
									assign node228 = (inp[8]) ? node230 : 3'b101;
										assign node230 = (inp[6]) ? 3'b100 : 3'b101;
						assign node234 = (inp[5]) ? node240 : node235;
							assign node235 = (inp[8]) ? node237 : 3'b100;
								assign node237 = (inp[7]) ? 3'b101 : 3'b100;
							assign node240 = (inp[7]) ? node248 : node241;
								assign node241 = (inp[8]) ? node243 : 3'b001;
									assign node243 = (inp[11]) ? node245 : 3'b001;
										assign node245 = (inp[6]) ? 3'b000 : 3'b001;
								assign node248 = (inp[8]) ? node250 : 3'b000;
									assign node250 = (inp[11]) ? node252 : 3'b001;
										assign node252 = (inp[6]) ? 3'b000 : 3'b001;

endmodule