module dtc_split66_bm76 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node6;
	wire [3-1:0] node8;
	wire [3-1:0] node10;
	wire [3-1:0] node11;
	wire [3-1:0] node15;
	wire [3-1:0] node16;
	wire [3-1:0] node17;
	wire [3-1:0] node19;
	wire [3-1:0] node21;
	wire [3-1:0] node22;
	wire [3-1:0] node24;
	wire [3-1:0] node28;
	wire [3-1:0] node29;
	wire [3-1:0] node31;
	wire [3-1:0] node32;
	wire [3-1:0] node34;
	wire [3-1:0] node37;
	wire [3-1:0] node38;
	wire [3-1:0] node43;
	wire [3-1:0] node44;
	wire [3-1:0] node45;
	wire [3-1:0] node46;
	wire [3-1:0] node48;
	wire [3-1:0] node52;
	wire [3-1:0] node54;
	wire [3-1:0] node55;
	wire [3-1:0] node57;
	wire [3-1:0] node58;
	wire [3-1:0] node62;
	wire [3-1:0] node63;
	wire [3-1:0] node67;
	wire [3-1:0] node68;
	wire [3-1:0] node70;
	wire [3-1:0] node71;
	wire [3-1:0] node76;
	wire [3-1:0] node77;
	wire [3-1:0] node78;
	wire [3-1:0] node79;
	wire [3-1:0] node81;
	wire [3-1:0] node82;
	wire [3-1:0] node83;
	wire [3-1:0] node88;
	wire [3-1:0] node90;
	wire [3-1:0] node91;
	wire [3-1:0] node95;
	wire [3-1:0] node96;
	wire [3-1:0] node97;
	wire [3-1:0] node99;
	wire [3-1:0] node101;
	wire [3-1:0] node105;
	wire [3-1:0] node107;
	wire [3-1:0] node108;
	wire [3-1:0] node109;
	wire [3-1:0] node111;
	wire [3-1:0] node114;
	wire [3-1:0] node115;
	wire [3-1:0] node120;
	wire [3-1:0] node121;
	wire [3-1:0] node122;
	wire [3-1:0] node123;
	wire [3-1:0] node124;
	wire [3-1:0] node126;
	wire [3-1:0] node128;
	wire [3-1:0] node132;
	wire [3-1:0] node134;
	wire [3-1:0] node135;
	wire [3-1:0] node139;
	wire [3-1:0] node140;
	wire [3-1:0] node141;
	wire [3-1:0] node143;
	wire [3-1:0] node145;
	wire [3-1:0] node148;
	wire [3-1:0] node149;
	wire [3-1:0] node150;
	wire [3-1:0] node155;
	wire [3-1:0] node157;
	wire [3-1:0] node159;
	wire [3-1:0] node161;
	wire [3-1:0] node164;
	wire [3-1:0] node165;
	wire [3-1:0] node166;
	wire [3-1:0] node167;
	wire [3-1:0] node168;
	wire [3-1:0] node173;
	wire [3-1:0] node174;
	wire [3-1:0] node176;
	wire [3-1:0] node178;
	wire [3-1:0] node182;
	wire [3-1:0] node183;
	wire [3-1:0] node184;
	wire [3-1:0] node186;
	wire [3-1:0] node188;
	wire [3-1:0] node192;
	wire [3-1:0] node194;
	wire [3-1:0] node196;
	wire [3-1:0] node199;
	wire [3-1:0] node200;
	wire [3-1:0] node201;
	wire [3-1:0] node202;
	wire [3-1:0] node203;
	wire [3-1:0] node204;
	wire [3-1:0] node205;
	wire [3-1:0] node209;
	wire [3-1:0] node210;
	wire [3-1:0] node211;
	wire [3-1:0] node216;
	wire [3-1:0] node217;
	wire [3-1:0] node218;
	wire [3-1:0] node219;
	wire [3-1:0] node220;
	wire [3-1:0] node226;
	wire [3-1:0] node227;
	wire [3-1:0] node229;
	wire [3-1:0] node233;
	wire [3-1:0] node234;
	wire [3-1:0] node235;
	wire [3-1:0] node237;
	wire [3-1:0] node239;
	wire [3-1:0] node243;
	wire [3-1:0] node245;
	wire [3-1:0] node246;
	wire [3-1:0] node247;
	wire [3-1:0] node249;
	wire [3-1:0] node250;
	wire [3-1:0] node256;
	wire [3-1:0] node257;
	wire [3-1:0] node258;
	wire [3-1:0] node259;
	wire [3-1:0] node260;
	wire [3-1:0] node261;
	wire [3-1:0] node263;
	wire [3-1:0] node266;
	wire [3-1:0] node267;
	wire [3-1:0] node272;
	wire [3-1:0] node274;
	wire [3-1:0] node275;
	wire [3-1:0] node277;
	wire [3-1:0] node280;
	wire [3-1:0] node281;
	wire [3-1:0] node285;
	wire [3-1:0] node286;
	wire [3-1:0] node288;
	wire [3-1:0] node289;
	wire [3-1:0] node293;
	wire [3-1:0] node295;
	wire [3-1:0] node297;
	wire [3-1:0] node298;
	wire [3-1:0] node300;
	wire [3-1:0] node304;
	wire [3-1:0] node305;
	wire [3-1:0] node306;
	wire [3-1:0] node307;
	wire [3-1:0] node308;
	wire [3-1:0] node310;
	wire [3-1:0] node314;
	wire [3-1:0] node316;
	wire [3-1:0] node317;
	wire [3-1:0] node321;
	wire [3-1:0] node323;
	wire [3-1:0] node325;
	wire [3-1:0] node326;
	wire [3-1:0] node330;
	wire [3-1:0] node331;
	wire [3-1:0] node332;
	wire [3-1:0] node333;
	wire [3-1:0] node337;
	wire [3-1:0] node338;
	wire [3-1:0] node342;
	wire [3-1:0] node344;
	wire [3-1:0] node346;
	wire [3-1:0] node348;
	wire [3-1:0] node351;
	wire [3-1:0] node352;
	wire [3-1:0] node353;
	wire [3-1:0] node354;
	wire [3-1:0] node355;
	wire [3-1:0] node357;
	wire [3-1:0] node359;
	wire [3-1:0] node363;
	wire [3-1:0] node365;
	wire [3-1:0] node366;
	wire [3-1:0] node368;
	wire [3-1:0] node369;
	wire [3-1:0] node374;
	wire [3-1:0] node375;
	wire [3-1:0] node376;
	wire [3-1:0] node378;
	wire [3-1:0] node382;
	wire [3-1:0] node384;
	wire [3-1:0] node385;
	wire [3-1:0] node386;
	wire [3-1:0] node391;
	wire [3-1:0] node392;
	wire [3-1:0] node393;
	wire [3-1:0] node394;
	wire [3-1:0] node395;
	wire [3-1:0] node396;
	wire [3-1:0] node401;
	wire [3-1:0] node402;
	wire [3-1:0] node404;
	wire [3-1:0] node406;
	wire [3-1:0] node409;
	wire [3-1:0] node410;
	wire [3-1:0] node411;
	wire [3-1:0] node416;
	wire [3-1:0] node417;
	wire [3-1:0] node418;
	wire [3-1:0] node419;
	wire [3-1:0] node421;
	wire [3-1:0] node425;
	wire [3-1:0] node426;
	wire [3-1:0] node430;
	wire [3-1:0] node432;
	wire [3-1:0] node434;
	wire [3-1:0] node437;
	wire [3-1:0] node438;
	wire [3-1:0] node439;
	wire [3-1:0] node440;
	wire [3-1:0] node441;
	wire [3-1:0] node445;
	wire [3-1:0] node447;
	wire [3-1:0] node449;
	wire [3-1:0] node452;
	wire [3-1:0] node454;
	wire [3-1:0] node455;
	wire [3-1:0] node456;
	wire [3-1:0] node461;
	wire [3-1:0] node462;
	wire [3-1:0] node466;
	wire [3-1:0] node467;
	wire [3-1:0] node468;
	wire [3-1:0] node469;
	wire [3-1:0] node470;
	wire [3-1:0] node471;
	wire [3-1:0] node472;
	wire [3-1:0] node474;
	wire [3-1:0] node476;
	wire [3-1:0] node477;
	wire [3-1:0] node482;
	wire [3-1:0] node484;
	wire [3-1:0] node485;
	wire [3-1:0] node486;
	wire [3-1:0] node491;
	wire [3-1:0] node492;
	wire [3-1:0] node493;
	wire [3-1:0] node495;
	wire [3-1:0] node496;
	wire [3-1:0] node501;
	wire [3-1:0] node503;
	wire [3-1:0] node504;
	wire [3-1:0] node505;
	wire [3-1:0] node510;
	wire [3-1:0] node511;
	wire [3-1:0] node512;
	wire [3-1:0] node513;
	wire [3-1:0] node514;
	wire [3-1:0] node515;
	wire [3-1:0] node520;
	wire [3-1:0] node521;
	wire [3-1:0] node523;
	wire [3-1:0] node525;
	wire [3-1:0] node528;
	wire [3-1:0] node529;
	wire [3-1:0] node533;
	wire [3-1:0] node534;
	wire [3-1:0] node535;
	wire [3-1:0] node537;
	wire [3-1:0] node541;
	wire [3-1:0] node543;
	wire [3-1:0] node544;
	wire [3-1:0] node548;
	wire [3-1:0] node549;
	wire [3-1:0] node550;
	wire [3-1:0] node553;
	wire [3-1:0] node554;
	wire [3-1:0] node556;
	wire [3-1:0] node558;
	wire [3-1:0] node562;
	wire [3-1:0] node563;
	wire [3-1:0] node564;
	wire [3-1:0] node566;
	wire [3-1:0] node570;
	wire [3-1:0] node572;
	wire [3-1:0] node573;
	wire [3-1:0] node576;
	wire [3-1:0] node577;
	wire [3-1:0] node581;
	wire [3-1:0] node582;
	wire [3-1:0] node583;
	wire [3-1:0] node584;
	wire [3-1:0] node585;
	wire [3-1:0] node587;
	wire [3-1:0] node591;
	wire [3-1:0] node592;
	wire [3-1:0] node594;
	wire [3-1:0] node597;
	wire [3-1:0] node598;
	wire [3-1:0] node599;
	wire [3-1:0] node600;
	wire [3-1:0] node606;
	wire [3-1:0] node607;
	wire [3-1:0] node608;
	wire [3-1:0] node609;
	wire [3-1:0] node611;
	wire [3-1:0] node613;
	wire [3-1:0] node616;
	wire [3-1:0] node617;
	wire [3-1:0] node621;
	wire [3-1:0] node623;
	wire [3-1:0] node625;
	wire [3-1:0] node628;
	wire [3-1:0] node629;
	wire [3-1:0] node631;
	wire [3-1:0] node633;
	wire [3-1:0] node635;
	wire [3-1:0] node638;
	wire [3-1:0] node639;
	wire [3-1:0] node640;
	wire [3-1:0] node641;
	wire [3-1:0] node647;
	wire [3-1:0] node648;
	wire [3-1:0] node649;
	wire [3-1:0] node650;
	wire [3-1:0] node651;
	wire [3-1:0] node655;
	wire [3-1:0] node656;
	wire [3-1:0] node658;
	wire [3-1:0] node662;
	wire [3-1:0] node663;
	wire [3-1:0] node664;
	wire [3-1:0] node670;
	wire [3-1:0] node671;
	wire [3-1:0] node672;
	wire [3-1:0] node673;
	wire [3-1:0] node674;
	wire [3-1:0] node675;
	wire [3-1:0] node677;
	wire [3-1:0] node681;
	wire [3-1:0] node682;
	wire [3-1:0] node684;
	wire [3-1:0] node686;
	wire [3-1:0] node688;
	wire [3-1:0] node691;
	wire [3-1:0] node692;
	wire [3-1:0] node694;
	wire [3-1:0] node695;
	wire [3-1:0] node700;
	wire [3-1:0] node701;
	wire [3-1:0] node702;
	wire [3-1:0] node704;

	assign outp = (inp[9]) ? node466 : node1;
		assign node1 = (inp[6]) ? node199 : node2;
			assign node2 = (inp[10]) ? node76 : node3;
				assign node3 = (inp[7]) ? node15 : node4;
					assign node4 = (inp[11]) ? node6 : 3'b111;
						assign node6 = (inp[3]) ? node8 : 3'b111;
							assign node8 = (inp[8]) ? node10 : 3'b111;
								assign node10 = (inp[4]) ? 3'b011 : node11;
									assign node11 = (inp[0]) ? 3'b011 : 3'b111;
					assign node15 = (inp[11]) ? node43 : node16;
						assign node16 = (inp[8]) ? node28 : node17;
							assign node17 = (inp[3]) ? node19 : 3'b111;
								assign node19 = (inp[4]) ? node21 : 3'b111;
									assign node21 = (inp[1]) ? 3'b011 : node22;
										assign node22 = (inp[0]) ? node24 : 3'b111;
											assign node24 = (inp[5]) ? 3'b011 : 3'b111;
							assign node28 = (inp[3]) ? 3'b011 : node29;
								assign node29 = (inp[4]) ? node31 : 3'b111;
									assign node31 = (inp[0]) ? node37 : node32;
										assign node32 = (inp[5]) ? node34 : 3'b111;
											assign node34 = (inp[2]) ? 3'b011 : 3'b111;
										assign node37 = (inp[2]) ? 3'b011 : node38;
											assign node38 = (inp[1]) ? 3'b011 : 3'b111;
						assign node43 = (inp[8]) ? node67 : node44;
							assign node44 = (inp[4]) ? node52 : node45;
								assign node45 = (inp[3]) ? 3'b011 : node46;
									assign node46 = (inp[0]) ? node48 : 3'b111;
										assign node48 = (inp[5]) ? 3'b011 : 3'b111;
								assign node52 = (inp[3]) ? node54 : 3'b011;
									assign node54 = (inp[0]) ? node62 : node55;
										assign node55 = (inp[5]) ? node57 : 3'b011;
											assign node57 = (inp[2]) ? 3'b101 : node58;
												assign node58 = (inp[1]) ? 3'b101 : 3'b011;
										assign node62 = (inp[2]) ? 3'b101 : node63;
											assign node63 = (inp[5]) ? 3'b101 : 3'b011;
							assign node67 = (inp[3]) ? 3'b101 : node68;
								assign node68 = (inp[4]) ? node70 : 3'b011;
									assign node70 = (inp[5]) ? 3'b101 : node71;
										assign node71 = (inp[0]) ? 3'b101 : 3'b011;
				assign node76 = (inp[7]) ? node120 : node77;
					assign node77 = (inp[11]) ? node95 : node78;
						assign node78 = (inp[8]) ? node88 : node79;
							assign node79 = (inp[3]) ? node81 : 3'b111;
								assign node81 = (inp[5]) ? 3'b011 : node82;
									assign node82 = (inp[2]) ? 3'b011 : node83;
										assign node83 = (inp[4]) ? 3'b011 : 3'b111;
							assign node88 = (inp[3]) ? node90 : 3'b011;
								assign node90 = (inp[4]) ? 3'b101 : node91;
									assign node91 = (inp[5]) ? 3'b101 : 3'b011;
						assign node95 = (inp[3]) ? node105 : node96;
							assign node96 = (inp[8]) ? 3'b101 : node97;
								assign node97 = (inp[0]) ? node99 : 3'b011;
									assign node99 = (inp[4]) ? node101 : 3'b011;
										assign node101 = (inp[5]) ? 3'b101 : 3'b011;
							assign node105 = (inp[8]) ? node107 : 3'b101;
								assign node107 = (inp[4]) ? 3'b001 : node108;
									assign node108 = (inp[1]) ? node114 : node109;
										assign node109 = (inp[0]) ? node111 : 3'b101;
											assign node111 = (inp[5]) ? 3'b001 : 3'b101;
										assign node114 = (inp[5]) ? 3'b001 : node115;
											assign node115 = (inp[0]) ? 3'b001 : 3'b101;
					assign node120 = (inp[11]) ? node164 : node121;
						assign node121 = (inp[8]) ? node139 : node122;
							assign node122 = (inp[3]) ? node132 : node123;
								assign node123 = (inp[4]) ? 3'b101 : node124;
									assign node124 = (inp[5]) ? node126 : 3'b011;
										assign node126 = (inp[1]) ? node128 : 3'b011;
											assign node128 = (inp[0]) ? 3'b101 : 3'b111;
								assign node132 = (inp[4]) ? node134 : 3'b101;
									assign node134 = (inp[5]) ? 3'b001 : node135;
										assign node135 = (inp[0]) ? 3'b001 : 3'b101;
							assign node139 = (inp[3]) ? node155 : node140;
								assign node140 = (inp[4]) ? node148 : node141;
									assign node141 = (inp[2]) ? node143 : 3'b101;
										assign node143 = (inp[5]) ? node145 : 3'b101;
											assign node145 = (inp[0]) ? 3'b001 : 3'b101;
									assign node148 = (inp[5]) ? 3'b001 : node149;
										assign node149 = (inp[2]) ? 3'b001 : node150;
											assign node150 = (inp[0]) ? 3'b001 : 3'b101;
								assign node155 = (inp[0]) ? node157 : 3'b001;
									assign node157 = (inp[5]) ? node159 : 3'b001;
										assign node159 = (inp[4]) ? node161 : 3'b001;
											assign node161 = (inp[1]) ? 3'b110 : 3'b001;
						assign node164 = (inp[8]) ? node182 : node165;
							assign node165 = (inp[3]) ? node173 : node166;
								assign node166 = (inp[5]) ? 3'b001 : node167;
									assign node167 = (inp[0]) ? 3'b001 : node168;
										assign node168 = (inp[4]) ? 3'b001 : 3'b101;
								assign node173 = (inp[4]) ? 3'b110 : node174;
									assign node174 = (inp[5]) ? node176 : 3'b001;
										assign node176 = (inp[2]) ? node178 : 3'b001;
											assign node178 = (inp[0]) ? 3'b110 : 3'b001;
							assign node182 = (inp[4]) ? node192 : node183;
								assign node183 = (inp[3]) ? 3'b110 : node184;
									assign node184 = (inp[2]) ? node186 : 3'b001;
										assign node186 = (inp[0]) ? node188 : 3'b001;
											assign node188 = (inp[5]) ? 3'b110 : 3'b001;
								assign node192 = (inp[3]) ? node194 : 3'b110;
									assign node194 = (inp[0]) ? node196 : 3'b110;
										assign node196 = (inp[5]) ? 3'b010 : 3'b110;
			assign node199 = (inp[10]) ? node351 : node200;
				assign node200 = (inp[7]) ? node256 : node201;
					assign node201 = (inp[11]) ? node233 : node202;
						assign node202 = (inp[3]) ? node216 : node203;
							assign node203 = (inp[8]) ? node209 : node204;
								assign node204 = (inp[1]) ? 3'b011 : node205;
									assign node205 = (inp[2]) ? 3'b101 : 3'b011;
								assign node209 = (inp[0]) ? 3'b101 : node210;
									assign node210 = (inp[4]) ? 3'b101 : node211;
										assign node211 = (inp[5]) ? 3'b101 : 3'b011;
							assign node216 = (inp[8]) ? node226 : node217;
								assign node217 = (inp[1]) ? 3'b101 : node218;
									assign node218 = (inp[4]) ? 3'b101 : node219;
										assign node219 = (inp[5]) ? 3'b101 : node220;
											assign node220 = (inp[0]) ? 3'b101 : 3'b011;
								assign node226 = (inp[4]) ? 3'b001 : node227;
									assign node227 = (inp[0]) ? node229 : 3'b101;
										assign node229 = (inp[5]) ? 3'b001 : 3'b101;
						assign node233 = (inp[3]) ? node243 : node234;
							assign node234 = (inp[8]) ? 3'b001 : node235;
								assign node235 = (inp[0]) ? node237 : 3'b101;
									assign node237 = (inp[4]) ? node239 : 3'b101;
										assign node239 = (inp[5]) ? 3'b001 : 3'b101;
							assign node243 = (inp[8]) ? node245 : 3'b001;
								assign node245 = (inp[4]) ? 3'b110 : node246;
									assign node246 = (inp[0]) ? 3'b110 : node247;
										assign node247 = (inp[5]) ? node249 : 3'b001;
											assign node249 = (inp[2]) ? 3'b110 : node250;
												assign node250 = (inp[1]) ? 3'b110 : 3'b001;
					assign node256 = (inp[11]) ? node304 : node257;
						assign node257 = (inp[8]) ? node285 : node258;
							assign node258 = (inp[3]) ? node272 : node259;
								assign node259 = (inp[4]) ? 3'b001 : node260;
									assign node260 = (inp[1]) ? node266 : node261;
										assign node261 = (inp[5]) ? node263 : 3'b101;
											assign node263 = (inp[0]) ? 3'b001 : 3'b101;
										assign node266 = (inp[0]) ? 3'b001 : node267;
											assign node267 = (inp[5]) ? 3'b001 : 3'b101;
								assign node272 = (inp[4]) ? node274 : 3'b001;
									assign node274 = (inp[5]) ? node280 : node275;
										assign node275 = (inp[0]) ? node277 : 3'b001;
											assign node277 = (inp[1]) ? 3'b110 : 3'b111;
										assign node280 = (inp[2]) ? 3'b110 : node281;
											assign node281 = (inp[1]) ? 3'b110 : 3'b111;
							assign node285 = (inp[3]) ? node293 : node286;
								assign node286 = (inp[4]) ? node288 : 3'b001;
									assign node288 = (inp[0]) ? 3'b110 : node289;
										assign node289 = (inp[5]) ? 3'b110 : 3'b001;
								assign node293 = (inp[5]) ? node295 : 3'b110;
									assign node295 = (inp[0]) ? node297 : 3'b110;
										assign node297 = (inp[1]) ? 3'b010 : node298;
											assign node298 = (inp[2]) ? node300 : 3'b110;
												assign node300 = (inp[4]) ? 3'b010 : 3'b110;
						assign node304 = (inp[8]) ? node330 : node305;
							assign node305 = (inp[1]) ? node321 : node306;
								assign node306 = (inp[3]) ? node314 : node307;
									assign node307 = (inp[4]) ? 3'b110 : node308;
										assign node308 = (inp[5]) ? node310 : 3'b001;
											assign node310 = (inp[0]) ? 3'b110 : 3'b001;
									assign node314 = (inp[4]) ? node316 : 3'b110;
										assign node316 = (inp[0]) ? 3'b010 : node317;
											assign node317 = (inp[5]) ? 3'b010 : 3'b110;
								assign node321 = (inp[4]) ? node323 : 3'b110;
									assign node323 = (inp[3]) ? node325 : 3'b110;
										assign node325 = (inp[5]) ? 3'b010 : node326;
											assign node326 = (inp[0]) ? 3'b010 : 3'b110;
							assign node330 = (inp[3]) ? node342 : node331;
								assign node331 = (inp[1]) ? node337 : node332;
									assign node332 = (inp[2]) ? 3'b110 : node333;
										assign node333 = (inp[5]) ? 3'b010 : 3'b110;
									assign node337 = (inp[2]) ? 3'b010 : node338;
										assign node338 = (inp[5]) ? 3'b010 : 3'b110;
								assign node342 = (inp[0]) ? node344 : 3'b010;
									assign node344 = (inp[1]) ? node346 : 3'b010;
										assign node346 = (inp[2]) ? node348 : 3'b100;
											assign node348 = (inp[4]) ? 3'b100 : 3'b010;
				assign node351 = (inp[7]) ? node391 : node352;
					assign node352 = (inp[11]) ? node374 : node353;
						assign node353 = (inp[8]) ? node363 : node354;
							assign node354 = (inp[3]) ? 3'b110 : node355;
								assign node355 = (inp[0]) ? node357 : 3'b001;
									assign node357 = (inp[5]) ? node359 : 3'b001;
										assign node359 = (inp[4]) ? 3'b110 : 3'b001;
							assign node363 = (inp[3]) ? node365 : 3'b110;
								assign node365 = (inp[4]) ? 3'b010 : node366;
									assign node366 = (inp[1]) ? node368 : 3'b110;
										assign node368 = (inp[0]) ? 3'b010 : node369;
											assign node369 = (inp[5]) ? 3'b010 : 3'b110;
						assign node374 = (inp[8]) ? node382 : node375;
							assign node375 = (inp[3]) ? 3'b010 : node376;
								assign node376 = (inp[2]) ? node378 : 3'b110;
									assign node378 = (inp[4]) ? 3'b010 : 3'b110;
							assign node382 = (inp[3]) ? node384 : 3'b010;
								assign node384 = (inp[4]) ? 3'b100 : node385;
									assign node385 = (inp[5]) ? 3'b100 : node386;
										assign node386 = (inp[0]) ? 3'b100 : 3'b010;
					assign node391 = (inp[11]) ? node437 : node392;
						assign node392 = (inp[3]) ? node416 : node393;
							assign node393 = (inp[8]) ? node401 : node394;
								assign node394 = (inp[0]) ? 3'b010 : node395;
									assign node395 = (inp[4]) ? 3'b010 : node396;
										assign node396 = (inp[5]) ? 3'b010 : 3'b110;
								assign node401 = (inp[4]) ? node409 : node402;
									assign node402 = (inp[0]) ? node404 : 3'b010;
										assign node404 = (inp[5]) ? node406 : 3'b010;
											assign node406 = (inp[2]) ? 3'b100 : 3'b010;
									assign node409 = (inp[1]) ? 3'b100 : node410;
										assign node410 = (inp[2]) ? 3'b100 : node411;
											assign node411 = (inp[5]) ? 3'b100 : 3'b010;
							assign node416 = (inp[8]) ? node430 : node417;
								assign node417 = (inp[4]) ? node425 : node418;
									assign node418 = (inp[1]) ? 3'b010 : node419;
										assign node419 = (inp[0]) ? node421 : 3'b010;
											assign node421 = (inp[2]) ? 3'b100 : 3'b010;
									assign node425 = (inp[0]) ? 3'b100 : node426;
										assign node426 = (inp[5]) ? 3'b100 : 3'b010;
								assign node430 = (inp[5]) ? node432 : 3'b100;
									assign node432 = (inp[4]) ? node434 : 3'b100;
										assign node434 = (inp[0]) ? 3'b000 : 3'b100;
						assign node437 = (inp[8]) ? node461 : node438;
							assign node438 = (inp[4]) ? node452 : node439;
								assign node439 = (inp[5]) ? node445 : node440;
									assign node440 = (inp[3]) ? 3'b100 : node441;
										assign node441 = (inp[0]) ? 3'b100 : 3'b010;
									assign node445 = (inp[2]) ? node447 : 3'b100;
										assign node447 = (inp[0]) ? node449 : 3'b100;
											assign node449 = (inp[3]) ? 3'b000 : 3'b100;
								assign node452 = (inp[3]) ? node454 : 3'b100;
									assign node454 = (inp[5]) ? 3'b000 : node455;
										assign node455 = (inp[2]) ? 3'b000 : node456;
											assign node456 = (inp[1]) ? 3'b000 : 3'b100;
							assign node461 = (inp[4]) ? 3'b000 : node462;
								assign node462 = (inp[3]) ? 3'b000 : 3'b100;
		assign node466 = (inp[6]) ? node670 : node467;
			assign node467 = (inp[10]) ? node581 : node468;
				assign node468 = (inp[7]) ? node510 : node469;
					assign node469 = (inp[11]) ? node491 : node470;
						assign node470 = (inp[3]) ? node482 : node471;
							assign node471 = (inp[8]) ? 3'b001 : node472;
								assign node472 = (inp[5]) ? node474 : 3'b101;
									assign node474 = (inp[4]) ? node476 : 3'b101;
										assign node476 = (inp[0]) ? 3'b001 : node477;
											assign node477 = (inp[1]) ? 3'b001 : 3'b101;
							assign node482 = (inp[8]) ? node484 : 3'b001;
								assign node484 = (inp[5]) ? 3'b110 : node485;
									assign node485 = (inp[4]) ? 3'b110 : node486;
										assign node486 = (inp[0]) ? 3'b110 : 3'b001;
						assign node491 = (inp[8]) ? node501 : node492;
							assign node492 = (inp[3]) ? 3'b110 : node493;
								assign node493 = (inp[4]) ? node495 : 3'b001;
									assign node495 = (inp[5]) ? 3'b110 : node496;
										assign node496 = (inp[0]) ? 3'b110 : 3'b001;
							assign node501 = (inp[3]) ? node503 : 3'b110;
								assign node503 = (inp[5]) ? 3'b010 : node504;
									assign node504 = (inp[4]) ? 3'b010 : node505;
										assign node505 = (inp[0]) ? 3'b010 : 3'b110;
					assign node510 = (inp[11]) ? node548 : node511;
						assign node511 = (inp[8]) ? node533 : node512;
							assign node512 = (inp[3]) ? node520 : node513;
								assign node513 = (inp[5]) ? 3'b110 : node514;
									assign node514 = (inp[4]) ? 3'b110 : node515;
										assign node515 = (inp[0]) ? 3'b110 : 3'b001;
								assign node520 = (inp[4]) ? node528 : node521;
									assign node521 = (inp[1]) ? node523 : 3'b110;
										assign node523 = (inp[5]) ? node525 : 3'b110;
											assign node525 = (inp[0]) ? 3'b010 : 3'b110;
									assign node528 = (inp[5]) ? 3'b010 : node529;
										assign node529 = (inp[0]) ? 3'b010 : 3'b110;
							assign node533 = (inp[4]) ? node541 : node534;
								assign node534 = (inp[3]) ? 3'b010 : node535;
									assign node535 = (inp[0]) ? node537 : 3'b110;
										assign node537 = (inp[5]) ? 3'b010 : 3'b110;
								assign node541 = (inp[3]) ? node543 : 3'b010;
									assign node543 = (inp[0]) ? 3'b100 : node544;
										assign node544 = (inp[1]) ? 3'b010 : 3'b100;
						assign node548 = (inp[8]) ? node562 : node549;
							assign node549 = (inp[3]) ? node553 : node550;
								assign node550 = (inp[4]) ? 3'b010 : 3'b110;
								assign node553 = (inp[4]) ? 3'b100 : node554;
									assign node554 = (inp[5]) ? node556 : 3'b010;
										assign node556 = (inp[2]) ? node558 : 3'b010;
											assign node558 = (inp[0]) ? 3'b100 : 3'b010;
							assign node562 = (inp[4]) ? node570 : node563;
								assign node563 = (inp[3]) ? 3'b100 : node564;
									assign node564 = (inp[0]) ? node566 : 3'b010;
										assign node566 = (inp[5]) ? 3'b100 : 3'b010;
								assign node570 = (inp[3]) ? node572 : 3'b100;
									assign node572 = (inp[1]) ? node576 : node573;
										assign node573 = (inp[2]) ? 3'b000 : 3'b100;
										assign node576 = (inp[0]) ? 3'b000 : node577;
											assign node577 = (inp[5]) ? 3'b000 : 3'b100;
				assign node581 = (inp[7]) ? node647 : node582;
					assign node582 = (inp[11]) ? node606 : node583;
						assign node583 = (inp[8]) ? node591 : node584;
							assign node584 = (inp[3]) ? 3'b010 : node585;
								assign node585 = (inp[1]) ? node587 : 3'b110;
									assign node587 = (inp[4]) ? 3'b010 : 3'b110;
							assign node591 = (inp[3]) ? node597 : node592;
								assign node592 = (inp[2]) ? node594 : 3'b010;
									assign node594 = (inp[1]) ? 3'b010 : 3'b100;
								assign node597 = (inp[0]) ? 3'b100 : node598;
									assign node598 = (inp[5]) ? 3'b100 : node599;
										assign node599 = (inp[4]) ? 3'b100 : node600;
											assign node600 = (inp[2]) ? 3'b100 : 3'b010;
						assign node606 = (inp[8]) ? node628 : node607;
							assign node607 = (inp[3]) ? node621 : node608;
								assign node608 = (inp[4]) ? node616 : node609;
									assign node609 = (inp[0]) ? node611 : 3'b000;
										assign node611 = (inp[2]) ? node613 : 3'b000;
											assign node613 = (inp[5]) ? 3'b100 : 3'b000;
									assign node616 = (inp[5]) ? 3'b100 : node617;
										assign node617 = (inp[2]) ? 3'b100 : 3'b000;
								assign node621 = (inp[4]) ? node623 : 3'b100;
									assign node623 = (inp[5]) ? node625 : 3'b100;
										assign node625 = (inp[0]) ? 3'b000 : 3'b100;
							assign node628 = (inp[3]) ? node638 : node629;
								assign node629 = (inp[2]) ? node631 : 3'b100;
									assign node631 = (inp[1]) ? node633 : 3'b000;
										assign node633 = (inp[0]) ? node635 : 3'b100;
											assign node635 = (inp[4]) ? 3'b000 : 3'b100;
								assign node638 = (inp[2]) ? 3'b000 : node639;
									assign node639 = (inp[4]) ? 3'b000 : node640;
										assign node640 = (inp[5]) ? 3'b000 : node641;
											assign node641 = (inp[0]) ? 3'b000 : 3'b100;
					assign node647 = (inp[11]) ? 3'b000 : node648;
						assign node648 = (inp[8]) ? node662 : node649;
							assign node649 = (inp[3]) ? node655 : node650;
								assign node650 = (inp[4]) ? 3'b100 : node651;
									assign node651 = (inp[0]) ? 3'b100 : 3'b000;
								assign node655 = (inp[4]) ? 3'b000 : node656;
									assign node656 = (inp[5]) ? node658 : 3'b100;
										assign node658 = (inp[0]) ? 3'b000 : 3'b100;
							assign node662 = (inp[4]) ? 3'b000 : node663;
								assign node663 = (inp[5]) ? 3'b000 : node664;
									assign node664 = (inp[0]) ? 3'b000 : 3'b100;
			assign node670 = (inp[7]) ? 3'b000 : node671;
				assign node671 = (inp[10]) ? 3'b000 : node672;
					assign node672 = (inp[11]) ? node700 : node673;
						assign node673 = (inp[8]) ? node681 : node674;
							assign node674 = (inp[3]) ? 3'b100 : node675;
								assign node675 = (inp[4]) ? node677 : 3'b010;
									assign node677 = (inp[1]) ? 3'b100 : 3'b010;
							assign node681 = (inp[3]) ? node691 : node682;
								assign node682 = (inp[2]) ? node684 : 3'b100;
									assign node684 = (inp[1]) ? node686 : 3'b000;
										assign node686 = (inp[5]) ? node688 : 3'b100;
											assign node688 = (inp[0]) ? 3'b000 : 3'b100;
								assign node691 = (inp[2]) ? 3'b000 : node692;
									assign node692 = (inp[1]) ? node694 : 3'b000;
										assign node694 = (inp[4]) ? 3'b000 : node695;
											assign node695 = (inp[5]) ? 3'b000 : 3'b100;
						assign node700 = (inp[3]) ? 3'b000 : node701;
							assign node701 = (inp[8]) ? 3'b000 : node702;
								assign node702 = (inp[2]) ? node704 : 3'b100;
									assign node704 = (inp[4]) ? 3'b000 : 3'b100;

endmodule