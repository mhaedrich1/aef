module dtc_split66_bm96 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node5;
	wire [3-1:0] node7;
	wire [3-1:0] node8;
	wire [3-1:0] node9;
	wire [3-1:0] node11;
	wire [3-1:0] node13;
	wire [3-1:0] node18;
	wire [3-1:0] node19;
	wire [3-1:0] node20;
	wire [3-1:0] node21;
	wire [3-1:0] node23;
	wire [3-1:0] node24;
	wire [3-1:0] node27;
	wire [3-1:0] node31;
	wire [3-1:0] node32;
	wire [3-1:0] node33;
	wire [3-1:0] node34;
	wire [3-1:0] node35;
	wire [3-1:0] node36;
	wire [3-1:0] node39;
	wire [3-1:0] node42;
	wire [3-1:0] node43;
	wire [3-1:0] node45;
	wire [3-1:0] node49;
	wire [3-1:0] node50;
	wire [3-1:0] node53;
	wire [3-1:0] node55;
	wire [3-1:0] node58;
	wire [3-1:0] node59;
	wire [3-1:0] node61;
	wire [3-1:0] node63;
	wire [3-1:0] node65;
	wire [3-1:0] node68;
	wire [3-1:0] node69;
	wire [3-1:0] node70;
	wire [3-1:0] node73;
	wire [3-1:0] node74;
	wire [3-1:0] node76;
	wire [3-1:0] node79;
	wire [3-1:0] node82;
	wire [3-1:0] node83;
	wire [3-1:0] node85;
	wire [3-1:0] node88;
	wire [3-1:0] node89;
	wire [3-1:0] node93;
	wire [3-1:0] node94;
	wire [3-1:0] node96;
	wire [3-1:0] node98;
	wire [3-1:0] node100;
	wire [3-1:0] node102;
	wire [3-1:0] node105;
	wire [3-1:0] node106;
	wire [3-1:0] node107;
	wire [3-1:0] node108;
	wire [3-1:0] node109;
	wire [3-1:0] node112;
	wire [3-1:0] node116;
	wire [3-1:0] node118;
	wire [3-1:0] node121;
	wire [3-1:0] node122;
	wire [3-1:0] node124;
	wire [3-1:0] node128;
	wire [3-1:0] node129;
	wire [3-1:0] node130;
	wire [3-1:0] node131;
	wire [3-1:0] node133;
	wire [3-1:0] node134;
	wire [3-1:0] node137;
	wire [3-1:0] node140;
	wire [3-1:0] node141;
	wire [3-1:0] node144;
	wire [3-1:0] node145;
	wire [3-1:0] node148;
	wire [3-1:0] node151;
	wire [3-1:0] node152;
	wire [3-1:0] node153;
	wire [3-1:0] node154;
	wire [3-1:0] node155;
	wire [3-1:0] node158;
	wire [3-1:0] node160;
	wire [3-1:0] node163;
	wire [3-1:0] node165;
	wire [3-1:0] node168;
	wire [3-1:0] node169;
	wire [3-1:0] node172;
	wire [3-1:0] node174;
	wire [3-1:0] node177;
	wire [3-1:0] node178;
	wire [3-1:0] node180;
	wire [3-1:0] node182;
	wire [3-1:0] node184;
	wire [3-1:0] node187;
	wire [3-1:0] node188;
	wire [3-1:0] node189;
	wire [3-1:0] node193;
	wire [3-1:0] node194;
	wire [3-1:0] node197;
	wire [3-1:0] node200;
	wire [3-1:0] node201;
	wire [3-1:0] node202;
	wire [3-1:0] node204;
	wire [3-1:0] node206;
	wire [3-1:0] node208;
	wire [3-1:0] node211;
	wire [3-1:0] node212;
	wire [3-1:0] node213;
	wire [3-1:0] node215;
	wire [3-1:0] node217;
	wire [3-1:0] node220;
	wire [3-1:0] node222;
	wire [3-1:0] node226;
	wire [3-1:0] node227;
	wire [3-1:0] node228;
	wire [3-1:0] node230;
	wire [3-1:0] node232;
	wire [3-1:0] node234;
	wire [3-1:0] node237;
	wire [3-1:0] node239;
	wire [3-1:0] node241;
	wire [3-1:0] node244;
	wire [3-1:0] node245;
	wire [3-1:0] node246;
	wire [3-1:0] node247;
	wire [3-1:0] node250;
	wire [3-1:0] node253;
	wire [3-1:0] node255;
	wire [3-1:0] node257;
	wire [3-1:0] node260;
	wire [3-1:0] node261;
	wire [3-1:0] node263;
	wire [3-1:0] node264;

	assign outp = (inp[6]) ? node2 : 3'b000;
		assign node2 = (inp[7]) ? node18 : node3;
			assign node3 = (inp[8]) ? node5 : 3'b000;
				assign node5 = (inp[4]) ? node7 : 3'b000;
					assign node7 = (inp[10]) ? 3'b000 : node8;
						assign node8 = (inp[9]) ? 3'b000 : node9;
							assign node9 = (inp[3]) ? node11 : 3'b000;
								assign node11 = (inp[1]) ? node13 : 3'b000;
									assign node13 = (inp[2]) ? 3'b100 : 3'b000;
			assign node18 = (inp[3]) ? node128 : node19;
				assign node19 = (inp[4]) ? node31 : node20;
					assign node20 = (inp[1]) ? 3'b011 : node21;
						assign node21 = (inp[9]) ? node23 : 3'b011;
							assign node23 = (inp[5]) ? node27 : node24;
								assign node24 = (inp[10]) ? 3'b011 : 3'b111;
								assign node27 = (inp[10]) ? 3'b101 : 3'b011;
					assign node31 = (inp[1]) ? node93 : node32;
						assign node32 = (inp[0]) ? node58 : node33;
							assign node33 = (inp[9]) ? node49 : node34;
								assign node34 = (inp[11]) ? node42 : node35;
									assign node35 = (inp[8]) ? node39 : node36;
										assign node36 = (inp[10]) ? 3'b010 : 3'b001;
										assign node39 = (inp[10]) ? 3'b001 : 3'b010;
									assign node42 = (inp[10]) ? 3'b010 : node43;
										assign node43 = (inp[2]) ? node45 : 3'b010;
											assign node45 = (inp[8]) ? 3'b001 : 3'b010;
								assign node49 = (inp[10]) ? node53 : node50;
									assign node50 = (inp[11]) ? 3'b001 : 3'b010;
									assign node53 = (inp[5]) ? node55 : 3'b001;
										assign node55 = (inp[11]) ? 3'b010 : 3'b001;
							assign node58 = (inp[9]) ? node68 : node59;
								assign node59 = (inp[11]) ? node61 : 3'b001;
									assign node61 = (inp[10]) ? node63 : 3'b001;
										assign node63 = (inp[5]) ? node65 : 3'b001;
											assign node65 = (inp[8]) ? 3'b010 : 3'b001;
								assign node68 = (inp[2]) ? node82 : node69;
									assign node69 = (inp[11]) ? node73 : node70;
										assign node70 = (inp[10]) ? 3'b001 : 3'b110;
										assign node73 = (inp[10]) ? node79 : node74;
											assign node74 = (inp[8]) ? node76 : 3'b001;
												assign node76 = (inp[5]) ? 3'b001 : 3'b101;
											assign node79 = (inp[5]) ? 3'b010 : 3'b001;
									assign node82 = (inp[10]) ? node88 : node83;
										assign node83 = (inp[11]) ? node85 : 3'b110;
											assign node85 = (inp[5]) ? 3'b001 : 3'b101;
										assign node88 = (inp[11]) ? 3'b110 : node89;
											assign node89 = (inp[5]) ? 3'b001 : 3'b101;
						assign node93 = (inp[0]) ? node105 : node94;
							assign node94 = (inp[9]) ? node96 : 3'b010;
								assign node96 = (inp[5]) ? node98 : 3'b010;
									assign node98 = (inp[10]) ? node100 : 3'b010;
										assign node100 = (inp[8]) ? node102 : 3'b010;
											assign node102 = (inp[11]) ? 3'b001 : 3'b010;
							assign node105 = (inp[9]) ? node121 : node106;
								assign node106 = (inp[11]) ? node116 : node107;
									assign node107 = (inp[5]) ? 3'b010 : node108;
										assign node108 = (inp[8]) ? node112 : node109;
											assign node109 = (inp[10]) ? 3'b001 : 3'b010;
											assign node112 = (inp[10]) ? 3'b010 : 3'b001;
									assign node116 = (inp[8]) ? node118 : 3'b001;
										assign node118 = (inp[2]) ? 3'b010 : 3'b001;
								assign node121 = (inp[11]) ? 3'b010 : node122;
									assign node122 = (inp[8]) ? node124 : 3'b010;
										assign node124 = (inp[2]) ? 3'b001 : 3'b010;
				assign node128 = (inp[1]) ? node200 : node129;
					assign node129 = (inp[4]) ? node151 : node130;
						assign node130 = (inp[10]) ? node140 : node131;
							assign node131 = (inp[9]) ? node133 : 3'b111;
								assign node133 = (inp[11]) ? node137 : node134;
									assign node134 = (inp[0]) ? 3'b111 : 3'b110;
									assign node137 = (inp[0]) ? 3'b110 : 3'b111;
							assign node140 = (inp[9]) ? node144 : node141;
								assign node141 = (inp[0]) ? 3'b111 : 3'b110;
								assign node144 = (inp[0]) ? node148 : node145;
									assign node145 = (inp[5]) ? 3'b011 : 3'b111;
									assign node148 = (inp[5]) ? 3'b010 : 3'b110;
						assign node151 = (inp[0]) ? node177 : node152;
							assign node152 = (inp[9]) ? node168 : node153;
								assign node153 = (inp[10]) ? node163 : node154;
									assign node154 = (inp[8]) ? node158 : node155;
										assign node155 = (inp[11]) ? 3'b011 : 3'b111;
										assign node158 = (inp[2]) ? node160 : 3'b011;
											assign node160 = (inp[11]) ? 3'b111 : 3'b011;
									assign node163 = (inp[8]) ? node165 : 3'b001;
										assign node165 = (inp[11]) ? 3'b001 : 3'b101;
								assign node168 = (inp[11]) ? node172 : node169;
									assign node169 = (inp[10]) ? 3'b110 : 3'b001;
									assign node172 = (inp[10]) ? node174 : 3'b110;
										assign node174 = (inp[5]) ? 3'b010 : 3'b110;
							assign node177 = (inp[9]) ? node187 : node178;
								assign node178 = (inp[11]) ? node180 : 3'b110;
									assign node180 = (inp[5]) ? node182 : 3'b110;
										assign node182 = (inp[10]) ? node184 : 3'b110;
											assign node184 = (inp[8]) ? 3'b010 : 3'b110;
								assign node187 = (inp[5]) ? node193 : node188;
									assign node188 = (inp[11]) ? 3'b100 : node189;
										assign node189 = (inp[10]) ? 3'b100 : 3'b010;
									assign node193 = (inp[10]) ? node197 : node194;
										assign node194 = (inp[11]) ? 3'b100 : 3'b010;
										assign node197 = (inp[11]) ? 3'b000 : 3'b100;
					assign node200 = (inp[4]) ? node226 : node201;
						assign node201 = (inp[0]) ? node211 : node202;
							assign node202 = (inp[9]) ? node204 : 3'b100;
								assign node204 = (inp[5]) ? node206 : 3'b101;
									assign node206 = (inp[10]) ? node208 : 3'b101;
										assign node208 = (inp[11]) ? 3'b100 : 3'b101;
							assign node211 = (inp[9]) ? 3'b100 : node212;
								assign node212 = (inp[10]) ? node220 : node213;
									assign node213 = (inp[11]) ? node215 : 3'b101;
										assign node215 = (inp[8]) ? node217 : 3'b100;
											assign node217 = (inp[2]) ? 3'b101 : 3'b100;
									assign node220 = (inp[8]) ? node222 : 3'b100;
										assign node222 = (inp[11]) ? 3'b100 : 3'b101;
						assign node226 = (inp[0]) ? node244 : node227;
							assign node227 = (inp[9]) ? node237 : node228;
								assign node228 = (inp[8]) ? node230 : 3'b001;
									assign node230 = (inp[11]) ? node232 : 3'b001;
										assign node232 = (inp[5]) ? node234 : 3'b001;
											assign node234 = (inp[2]) ? 3'b001 : 3'b000;
								assign node237 = (inp[5]) ? node239 : 3'b010;
									assign node239 = (inp[8]) ? node241 : 3'b010;
										assign node241 = (inp[11]) ? 3'b100 : 3'b010;
							assign node244 = (inp[9]) ? node260 : node245;
								assign node245 = (inp[11]) ? node253 : node246;
									assign node246 = (inp[10]) ? node250 : node247;
										assign node247 = (inp[8]) ? 3'b110 : 3'b010;
										assign node250 = (inp[8]) ? 3'b010 : 3'b100;
									assign node253 = (inp[2]) ? node255 : 3'b100;
										assign node255 = (inp[8]) ? node257 : 3'b100;
											assign node257 = (inp[10]) ? 3'b100 : 3'b010;
								assign node260 = (inp[10]) ? 3'b000 : node261;
									assign node261 = (inp[8]) ? node263 : 3'b000;
										assign node263 = (inp[11]) ? 3'b000 : node264;
											assign node264 = (inp[2]) ? 3'b100 : 3'b000;

endmodule